2SAM|1|1|After the death of Saul, when David had returned from striking down the Amalekites, David remained two days in Ziklag.
2SAM|1|2|And on the third day, behold, a man came from Saul's camp, with his clothes torn and dirt on his head. And when he came to David, he fell to the ground and paid homage.
2SAM|1|3|David said to him, "Where do you come from?" And he said to him, "I have escaped from the camp of Israel."
2SAM|1|4|And David said to him, "How did it go? Tell me." And he answered, "The people fled from the battle, and also many of the people have fallen and are dead, and Saul and his son Jonathan are also dead."
2SAM|1|5|Then David said to the young man who told him, "How do you know that Saul and his son Jonathan are dead?"
2SAM|1|6|And the young man who told him said, "By chance I happened to be on Mount Gilboa, and there was Saul leaning on his spear, and behold, the chariots and the horsemen were close upon him.
2SAM|1|7|And when he looked behind him, he saw me, and called to me. And I answered, 'Here I am.'
2SAM|1|8|And he said to me, 'Who are you?' I answered him, 'I am an Amalekite.'
2SAM|1|9|And he said to me 'Stand beside me and kill me, for anguish has seized me, and yet my life still lingers.'
2SAM|1|10|So I stood beside him and killed him, because I was sure that he could not live after he had fallen. And I took the crown that was on his head and the armlet that was on his arm, and I have brought them here to my lord."
2SAM|1|11|Then David took hold of his clothes and tore them, and so did all the men who were with him.
2SAM|1|12|And they mourned and wept and fasted until evening for Saul and for Jonathan his son and for the people of the LORD and for the house of Israel, because they had fallen by the sword.
2SAM|1|13|And David said to the young man who told him, "Where do you come from?" And he answered, "I am the son of a sojourner, an Amalekite."
2SAM|1|14|David said to him, "How is it you were not afraid to put out your hand to destroy the LORD's anointed?"
2SAM|1|15|Then David called one of the young men and said, "Go, execute him." And he struck him down so that he died.
2SAM|1|16|And David said to him, "Your blood be on your head, for your own mouth has testified against you, saying, 'I have killed the LORD's anointed.'"
2SAM|1|17|And David lamented with this lamentation over Saul and Jonathan his son,
2SAM|1|18|and he said it should be taught to the people of Judah; behold, it is written in the Book of Jashar. He said:
2SAM|1|19|"Your glory, O Israel, is slain on your high places! How the mighty have fallen!
2SAM|1|20|Tell it not in Gath, publish it not in the streets of Ashkelon, lest the daughters of the Philistines rejoice, lest the daughters of the uncircumcised exult.
2SAM|1|21|"You mountains of Gilboa, let there be no dew or rain upon you, nor fields of offerings! For there the shield of the mighty was defiled, the shield of Saul, not anointed with oil.
2SAM|1|22|"From the blood of the slain, from the fat of the mighty, the bow of Jonathan turned not back, and the sword of Saul returned not empty.
2SAM|1|23|"Saul and Jonathan, beloved and lovely! In life and in death they were not divided; they were swifter than eagles; they were stronger than lions.
2SAM|1|24|"You daughters of Israel, weep over Saul, who clothed you luxuriously in scarlet, who put ornaments of gold on your apparel.
2SAM|1|25|"How the mighty have fallen in the midst of the battle! "Jonathan lies slain on your high places.
2SAM|1|26|I am distressed for you, my brother Jonathan; very pleasant have you been to me; your love to me was extraordinary, surpassing the love of women.
2SAM|1|27|"How the mighty have fallen, and the weapons of war perished!"
2SAM|2|1|After this David inquired of the LORD, "Shall I go up into any of the cities of Judah?" And the LORD said to him, "Go up." David said, "To which shall I go up?" And he said, "To Hebron."
2SAM|2|2|So David went up there, and his two wives also, Ahinoam of Jezreel and Abigail the widow of Nabal of Carmel.
2SAM|2|3|And David brought up his men who were with him, everyone with his household, and they lived in the towns of Hebron.
2SAM|2|4|And the men of Judah came, and there they anointed David king over the house of Judah. When they told David, "It was the men of Jabesh-gilead who buried Saul,"
2SAM|2|5|David sent messengers to the men of Jabesh-gilead and said to them, "May you be blessed by the LORD, because you showed this loyalty to Saul your lord and buried him.
2SAM|2|6|Now may the LORD show steadfast love and faithfulness to you. And I will do good to you because you have done this thing.
2SAM|2|7|Now therefore let your hands be strong, and be valiant, for Saul your lord is dead, and the house of Judah has anointed me king over them."
2SAM|2|8|But Abner the son of Ner, commander of Saul's army, took Ish-bosheth the son of Saul and brought him over to Mahanaim,
2SAM|2|9|and he made him king over Gilead and the Ashurites and Jezreel and Ephraim and Benjamin and all Israel.
2SAM|2|10|Ish-bosheth, Saul's son, was forty years old when he began to reign over Israel, and he reigned two years. But the house of Judah followed David.
2SAM|2|11|And the time that David was king in Hebron over the house of Judah was seven years and six months.
2SAM|2|12|Abner the son of Ner, and the servants of Ish-bosheth the son of Saul, went out from Mahanaim to Gibeon.
2SAM|2|13|And Joab the son of Zeruiah and the servants of David went out and met them at the pool of Gibeon. And they sat down, the one on the one side of the pool, and the other on the other side of the pool.
2SAM|2|14|And Abner said to Joab, "Let the young men arise and compete before us." And Joab said, "Let them arise."
2SAM|2|15|Then they arose and passed over by number, twelve for Benjamin and Ish-bosheth the son of Saul, and twelve of the servants of David.
2SAM|2|16|And each caught his opponent by the head and thrust his sword in his opponent's side, so they fell down together. Therefore that place was called Helkath-hazzurim, which is at Gibeon.
2SAM|2|17|And the battle was very fierce that day. And Abner and the men of Israel were beaten before the servants of David.
2SAM|2|18|And the three sons of Zeruiah were there, Joab, Abishai, and Asahel. Now Asahel was as swift of foot as a wild gazelle.
2SAM|2|19|And Asahel pursued Abner, and as he went, he turned neither to the right hand nor to the left from following Abner.
2SAM|2|20|Then Abner looked behind him and said, "Is it you, Asahel?" And he answered, "It is I."
2SAM|2|21|Abner said to him, "Turn aside to your right hand or to your left, and seize one of the young men and take his spoil." But Asahel would not turn aside from following him.
2SAM|2|22|And Abner said again to Asahel, "Turn aside from following me. Why should I strike you to the ground? How then could I lift up my face to your brother Joab?"
2SAM|2|23|But he refused to turn aside. Therefore Abner struck him in the stomach with the butt of his spear, so that the spear came out at his back. And he fell there and died where he was. And all who came to the place where Asahel had fallen and died, stood still.
2SAM|2|24|But Joab and Abishai pursued Abner. And as the sun was going down they came to the hill of Ammah, which lies before Giah on the way to the wilderness of Gibeon.
2SAM|2|25|And the people of Benjamin gathered themselves together behind Abner and became one group and took their stand on the top of a hill.
2SAM|2|26|Then Abner called to Joab, "Shall the sword devour forever? Do you not know that the end will be bitter? How long will it be before you tell your people to turn from the pursuit of their brothers?"
2SAM|2|27|And Joab said, "As God lives, if you had not spoken, surely the men would not have given up the pursuit of their brothers until the morning."
2SAM|2|28|So Joab blew the trumpet, and all the men stopped and pursued Israel no more, nor did they fight anymore.
2SAM|2|29|And Abner and his men went all that night through the Arabah. They crossed the Jordan, and marching the whole morning, they came to Mahanaim.
2SAM|2|30|Joab returned from the pursuit of Abner. And when he had gathered all the people together, there were missing from David's servants nineteen men besides Asahel.
2SAM|2|31|But the servants of David had struck down of Benjamin 360 of Abner's men.
2SAM|2|32|And they took up Asahel and buried him in the tomb of his father, which was at Bethlehem. And Joab and his men marched all night, and the day broke upon them at Hebron.
2SAM|3|1|There was a long war between the house of Saul and the house of David. And David grew stronger and stronger, while the house of Saul became weaker and weaker.
2SAM|3|2|And sons were born to David at Hebron: his firstborn was Amnon, of Ahinoam of Jezreel;
2SAM|3|3|and his second, Chileab, of Abigail the widow of Nabal of Carmel; and the third, Absalom the son of Maacah the daughter of Talmai king of Geshur;
2SAM|3|4|and the fourth, Adonijah the son of Haggith; and the fifth, Shephatiah the son of Abital;
2SAM|3|5|and the sixth, Ithream, of Eglah, David's wife. These were born to David in Hebron.
2SAM|3|6|While there was war between the house of Saul and the house of David, Abner was making himself strong in the house of Saul.
2SAM|3|7|Now Saul had a concubine whose name was Rizpah, the daughter of Aiah. And Ish-bosheth said to Abner, "Why have you gone in to my father's concubine?"
2SAM|3|8|Then Abner was very angry over the words of Ish-bosheth and said, "Am I a dog's head of Judah? To this day I keep showing steadfast love to the house of Saul your father, to his brothers, and to his friends, and have not given you into the hand of David. And yet you charge me today with a fault concerning a woman.
2SAM|3|9|God do so to Abner and more also, if I do not accomplish for David what the LORD has sworn to him,
2SAM|3|10|to transfer the kingdom from the house of Saul and set up the throne of David over Israel and over Judah, from Dan to Beersheba."
2SAM|3|11|And Ish-bosheth could not answer Abner another word, because he feared him.
2SAM|3|12|And Abner sent messengers to David on his behalf, saying, "To whom does the land belong? Make your covenant with me, and behold, my hand shall be with you to bring over all Israel to you."
2SAM|3|13|And he said, "Good; I will make a covenant with you. But one thing I require of you; that is, you shall not see my face unless you first bring Michal, Saul's daughter, when you come to see my face."
2SAM|3|14|Then David sent messengers to Ish-bosheth, Saul's son, saying, "Give me my wife Michal, for whom I paid the bridal price of a hundred foreskins of the Philistines."
2SAM|3|15|And Ish-bosheth sent and took her from her husband Paltiel the son of Laish.
2SAM|3|16|But her husband went with her, weeping after her all the way to Bahurim. Then Abner said to him, "Go, return." And he returned.
2SAM|3|17|And Abner conferred with the elders of Israel, saying, "For some time past you have been seeking David as king over you.
2SAM|3|18|Now then bring it about, for the LORD has promised David, saying, 'By the hand of my servant David I will save my people Israel from the hand of the Philistines, and from the hand of all their enemies.'"
2SAM|3|19|Abner also spoke to Benjamin. And then Abner went to tell David at Hebron all that Israel and the whole house of Benjamin thought good to do.
2SAM|3|20|When Abner came with twenty men to David at Hebron, David made a feast for Abner and the men who were with him.
2SAM|3|21|And Abner said to David, "I will arise and go and will gather all Israel to my lord the king, that they may make a covenant with you, and that you may reign over all that your heart desires." So David sent Abner away, and he went in peace.
2SAM|3|22|Just then the servants of David arrived with Joab from a raid, bringing much spoil with them. But Abner was not with David at Hebron, for he had sent him away, and he had gone in peace.
2SAM|3|23|When Joab and all the army that was with him came, it was told Joab, "Abner the son of Ner came to the king, and he has let him go, and he has gone in peace."
2SAM|3|24|Then Joab went to the king and said, "What have you done? Behold, Abner came to you. Why is it that you have sent him away, so that he is gone?
2SAM|3|25|You know that Abner the son of Ner came to deceive you and to know your going out and your coming in, and to know all that you are doing."
2SAM|3|26|When Joab came out from David's presence, he sent messengers after Abner, and they brought him back from the cistern of Sirah. But David did not know about it.
2SAM|3|27|And when Abner returned to Hebron, Joab took him aside into the midst of the gate to speak with him privately, and there he struck him in the stomach, so that he died, for the blood of Asahel his brother.
2SAM|3|28|Afterward, when David heard of it, he said, "I and my kingdom are forever guiltless before the LORD for the blood of Abner the son of Ner.
2SAM|3|29|May it fall upon the head of Joab and upon all his father's house, and may the house of Joab never be without one who has a discharge or who is leprous or who holds a spindle or who falls by the sword or who lacks bread!"
2SAM|3|30|So Joab and Abishai his brother killed Abner, because he had put their brother Asahel to death in the battle at Gibeon.
2SAM|3|31|Then David said to Joab and to all the people who were with him, "Tear your clothes and put on sackcloth and mourn before Abner." And King David followed the bier.
2SAM|3|32|They buried Abner at Hebron. And the king lifted up his voice and wept at the grave of Abner, and all the people wept.
2SAM|3|33|And the king lamented for Abner, saying, "Should Abner die as a fool dies?
2SAM|3|34|Your hands were not bound; your feet were not fettered; as one falls before the wicked you have fallen." And all the people wept again over him.
2SAM|3|35|Then all the people came to persuade David to eat bread while it was yet day. But David swore, saying, "God do so to me and more also, if I taste bread or anything else till the sun goes down!"
2SAM|3|36|And all the people took notice of it, and it pleased them, as everything that the king did pleased all the people.
2SAM|3|37|So all the people and all Israel understood that day that it had not been the king's will to put to death Abner the son of Ner.
2SAM|3|38|And the king said to his servants, "Do you not know that a prince and a great man has fallen this day in Israel?
2SAM|3|39|And I was gentle today, though anointed king. These men, the sons of Zeruiah, are more severe than I. The LORD repay the evildoer according to his wickedness!"
2SAM|4|1|When Ish-bosheth, Saul's son, heard that Abner had died at Hebron, his courage failed, and all Israel was dismayed.
2SAM|4|2|Now Saul's son had two men who were captains of raiding bands; the name of the one was Baanah, and the name of the other Rechab, sons of Rimmon a man of Benjamin from Beeroth (for Beeroth also is counted part of Benjamin;
2SAM|4|3|the Beerothites fled to Gittaim and have been sojourners there to this day).
2SAM|4|4|Jonathan, the son of Saul, had a son who was crippled in his feet. He was five years old when the news about Saul and Jonathan came from Jezreel, and his nurse took him up and fled, and as she fled in her haste, he fell and became lame. And his name was Mephibosheth.
2SAM|4|5|Now the sons of Rimmon the Beerothite, Rechab and Baanah, set out, and about the heat of the day they came to the house of Ish-bosheth as he was taking his noonday rest.
2SAM|4|6|And they came into the midst of the house as if to get wheat, and they stabbed him in the stomach. Then Rechab and Baanah his brother escaped.
2SAM|4|7|When they came into the house, as he lay on his bed in his bedroom, they struck him and put him to death and beheaded him. They took his head and went by the way of the Arabah all night,
2SAM|4|8|and brought the head of Ish-bosheth to David at Hebron. And they said to the king, "Here is the head of Ish-bosheth, the son of Saul, your enemy, who sought your life. The LORD has avenged my lord the king this day on Saul and on his offspring."
2SAM|4|9|But David answered Rechab and Baanah his brother, the sons of Rimmon the Beerothite, "As the LORD lives, who has redeemed my life out of every adversity,
2SAM|4|10|when one told me, 'Behold, Saul is dead,' and thought he was bringing good news, I seized him and killed him at Ziklag, which was the reward I gave him for his news.
2SAM|4|11|How much more, when wicked men have killed a righteous man in his own house on his bed, shall I not now require his blood at your hand and destroy you from the earth?"
2SAM|4|12|And David commanded his young men, and they killed them and cut off their hands and feet and hanged them beside the pool at Hebron. But they took the head of Ish-bosheth and buried it in the tomb of Abner at Hebron.
2SAM|5|1|Then all the tribes of Israel came to David at Hebron and said, "Behold, we are your bone and flesh.
2SAM|5|2|In times past, when Saul was king over us, it was you who led out and brought in Israel. And the LORD said to you, 'You shall be shepherd of my people Israel, and you shall be prince over Israel.'"
2SAM|5|3|So all the elders of Israel came to the king at Hebron, and King David made a covenant with them at Hebron before the LORD, and they anointed David king over Israel.
2SAM|5|4|David was thirty years old when he began to reign, and he reigned forty years.
2SAM|5|5|At Hebron he reigned over Judah seven years and six months, and at Jerusalem he reigned over all Israel and Judah thirty-three years.
2SAM|5|6|And the king and his men went to Jerusalem against the Jebusites, the inhabitants of the land, who said to David, "You will not come in here, but the blind and the lame will ward you off"- thinking, "David cannot come in here."
2SAM|5|7|Nevertheless, David took the stronghold of Zion, that is, the city of David.
2SAM|5|8|And David said on that day, "Whoever would strike the Jebusites, let him get up the water shaft to attack 'the lame and the blind,' who are hated by David's soul." Therefore it is said, "The blind and the lame shall not come into the house."
2SAM|5|9|And David lived in the stronghold and called it the city of David. And David built the city all around from the Millo inward.
2SAM|5|10|And David became greater and greater, for the LORD, the God of hosts, was with him.
2SAM|5|11|And Hiram king of Tyre sent messengers to David, and cedar trees, also carpenters and masons who built David a house.
2SAM|5|12|And David knew that the LORD had established him king over Israel, and that he had exalted his kingdom for the sake of his people Israel.
2SAM|5|13|And David took more concubines and wives from Jerusalem, after he came from Hebron, and more sons and daughters were born to David.
2SAM|5|14|And these are the names of those who were born to him in Jerusalem: Shammua, Shobab, Nathan, Solomon,
2SAM|5|15|Ibhar, Elishua, Nepheg, Japhia,
2SAM|5|16|Elishama, Eliada, and Eliphelet.
2SAM|5|17|When the Philistines heard that David had been anointed king over Israel, all the Philistines went up to search for David. But David heard of it and went down to the stronghold.
2SAM|5|18|Now the Philistines had come and spread out in the Valley of Rephaim.
2SAM|5|19|And David inquired of the LORD, "Shall I go up against the Philistines? Will you give them into my hand?" And the LORD said to David, "Go up, for I will certainly give the Philistines into your hand."
2SAM|5|20|And David came to Baal-perazim, and David defeated them there. And he said, "The LORD has burst through my enemies before me like a bursting flood." Therefore the name of that place is called Baal-perazim.
2SAM|5|21|And the Philistines left their idols there, and David and his men carried them away.
2SAM|5|22|And the Philistines came up yet again and spread out in the Valley of Rephaim.
2SAM|5|23|And when David inquired of the LORD, he said, "You shall not go up; go around to their rear, and come against them opposite the balsam trees.
2SAM|5|24|And when you hear the sound of marching in the tops of the balsam trees, then rouse yourself, for then the LORD has gone out before you to strike down the army of the Philistines."
2SAM|5|25|And David did as the LORD commanded him, and struck down the Philistines from Geba to Gezer.
2SAM|6|1|David again gathered all the chosen men of Israel, thirty thousand.
2SAM|6|2|And David arose and went with all the people who were with him from Baale-judah to bring up from there the ark of God, which is called by the name of the LORD of hosts who sits enthroned on the cherubim.
2SAM|6|3|And they carried the ark of God on a new cart and brought it out of the house of Abinadab, which was on the hill. And Uzzah and Ahio, the sons of Abinadab, were driving the new cart,
2SAM|6|4|with the ark of God, and Ahio went before the ark.
2SAM|6|5|And David and all the house of Israel were making merry before the LORD, with songs and lyres and harps and tambourines and castanets and cymbals.
2SAM|6|6|And when they came to the threshing floor of Nacon, Uzzah put out his hand to the ark of God and took hold of it, for the oxen stumbled.
2SAM|6|7|And the anger of the LORD was kindled against Uzzah, and God struck him down there because of his error, and he died there beside the ark of God.
2SAM|6|8|And David was angry because the LORD had burst forth against Uzzah. And that place is called Perez-uzzah, to this day.
2SAM|6|9|And David was afraid of the LORD that day, and he said, "How can the ark of the LORD come to me?"
2SAM|6|10|So David was not willing to take the ark of the LORD into the city of David. But David took it aside to the house of Obed-edom the Gittite.
2SAM|6|11|And the ark of the LORD remained in the house of Obed-edom the Gittite three months, and the LORD blessed Obed-edom and all his household.
2SAM|6|12|And it was told King David, "The LORD has blessed the household of Obed-edom and all that belongs to him, because of the ark of God." So David went and brought up the ark of God from the house of Obed-edom to the city of David with rejoicing.
2SAM|6|13|And when those who bore the ark of the LORD had gone six steps, he sacrificed an ox and a fattened animal.
2SAM|6|14|And David danced before the LORD with all his might. And David was wearing a linen ephod.
2SAM|6|15|So David and all the house of Israel brought up the ark of the LORD with shouting and with the sound of the horn.
2SAM|6|16|As the ark of the LORD came into the city of David, Michal the daughter of Saul looked out of the window and saw King David leaping and dancing before the LORD, and she despised him in her heart.
2SAM|6|17|And they brought in the ark of the LORD and set it in its place, inside the tent that David had pitched for it. And David offered burnt offerings and peace offerings before the LORD.
2SAM|6|18|And when David had finished offering the burnt offerings and the peace offerings, he blessed the people in the name of the LORD of hosts
2SAM|6|19|and distributed among all the people, the whole multitude of Israel, both men and women, a cake of bread, a portion of meat, and a cake of raisins to each one. Then all the people departed, each to his house.
2SAM|6|20|And David returned to bless his household. But Michal the daughter of Saul came out to meet David and said, "How the king of Israel honored himself today, uncovering himself today before the eyes of his servants' female servants, as one of the vulgar fellows shamelessly uncovers himself!"
2SAM|6|21|And David said to Michal, "It was before the LORD, who chose me above your father and above all his house, to appoint me as prince over Israel, the people of the LORD- and I will make merry before the LORD.
2SAM|6|22|I will make myself yet more contemptible than this, and I will be abased in your eyes. But by the female servants of whom you have spoken, by them I shall be held in honor."
2SAM|6|23|And Michal the daughter of Saul had no child to the day of her death.
2SAM|7|1|Now when the king lived in his house and the LORD had given him rest from all his surrounding enemies,
2SAM|7|2|the king said to Nathan the prophet, "See now, I dwell in a house of cedar, but the ark of God dwells in a tent."
2SAM|7|3|And Nathan said to the king, "Go, do all that is in your heart, for the LORD is with you."
2SAM|7|4|But that same night the word of the LORD came to Nathan,
2SAM|7|5|"Go and tell my servant David, 'Thus says the LORD: Would you build me a house to dwell in?
2SAM|7|6|I have not lived in a house since the day I brought up the people of Israel from Egypt to this day, but I have been moving about in a tent for my dwelling.
2SAM|7|7|In all places where I have moved with all the people of Israel, did I speak a word with any of the judges of Israel, whom I commanded to shepherd my people Israel, saying, "Why have you not built me a house of cedar?"'
2SAM|7|8|Now, therefore, thus you shall say to my servant David, 'Thus says the LORD of hosts, I took you from the pasture, from following the sheep, that you should be prince over my people Israel.
2SAM|7|9|And I have been with you wherever you went and have cut off all your enemies from before you. And I will make for you a great name, like the name of the great ones of the earth.
2SAM|7|10|And I will appoint a place for my people Israel and will plant them, so that they may dwell in their own place and be disturbed no more. And violent men shall afflict them no more, as formerly,
2SAM|7|11|from the time that I appointed judges over my people Israel. And I will give you rest from all your enemies. Moreover, the LORD declares to you that the LORD will make you a house.
2SAM|7|12|When your days are fulfilled and you lie down with your fathers, I will raise up your offspring after you, who shall come from your body, and I will establish his kingdom.
2SAM|7|13|He shall build a house for my name, and I will establish the throne of his kingdom forever.
2SAM|7|14|I will be to him a father, and he shall be to me a son. When he commits iniquity, I will discipline him with the rod of men, with the stripes of the sons of men,
2SAM|7|15|but my steadfast love will not depart from him, as I took it from Saul, whom I put away from before you.
2SAM|7|16|And your house and your kingdom shall be made sure forever before me. Your throne shall be established forever.'"
2SAM|7|17|In accordance with all these words, and in accordance with all this vision, Nathan spoke to David.
2SAM|7|18|Then King David went in and sat before the LORD and said, "Who am I, O Lord GOD, and what is my house, that you have brought me thus far?
2SAM|7|19|And yet this was a small thing in your eyes, O Lord GOD. You have spoken also of your servant's house for a great while to come, and this is instruction for mankind, O Lord GOD!
2SAM|7|20|And what more can David say to you? For you know your servant, O Lord GOD!
2SAM|7|21|Because of your promise, and according to your own heart, you have brought about all this greatness, to make your servant know it.
2SAM|7|22|Therefore you are great, O LORD God. For there is none like you, and there is no God besides you, according to all that we have heard with our ears.
2SAM|7|23|And who is like your people Israel, the one nation on earth whom God went to redeem to be his people, making himself a name and doing for them great and awesome things by driving out before your people, whom you redeemed for yourself from Egypt, a nation and its gods?
2SAM|7|24|And you established for yourself your people Israel to be your people forever. And you, O LORD, became their God.
2SAM|7|25|And now, O LORD God, confirm forever the word that you have spoken concerning your servant and concerning his house, and do as you have spoken.
2SAM|7|26|And your name will be magnified forever, saying, 'The LORD of hosts is God over Israel,' and the house of your servant David will be established before you.
2SAM|7|27|For you, O LORD of hosts, the God of Israel, have made this revelation to your servant, saying, 'I will build you a house.' Therefore your servant has found courage to pray this prayer to you.
2SAM|7|28|And now, O Lord GOD, you are God, and your words are true, and you have promised this good thing to your servant.
2SAM|7|29|Now therefore may it please you to bless the house of your servant, so that it may continue forever before you. For you, O Lord GOD, have spoken, and with your blessing shall the house of your servant be blessed forever."
2SAM|8|1|After this David defeated the Philistines and subdued them, and David took Metheg-ammah out of the hand of the Philistines.
2SAM|8|2|And he defeated Moab and he measured them with a line, making them lie down on the ground. Two lines he measured to be put to death, and one full line to be spared. And the Moabites became servants to David and brought tribute.
2SAM|8|3|David also defeated Hadadezer the son of Rehob, king of Zobah, as he went to restore his power at the river Euphrates.
2SAM|8|4|And David took from him 1,700 horsemen, and 20,000 foot soldiers. And David hamstrung all the chariot horses but left enough for a hundred chariots.
2SAM|8|5|And when the Syrians of Damascus came to help Hadadezer king of Zobah, David struck down 22,000 men of the Syrians.
2SAM|8|6|Then David put garrisons in Aram of Damascus, and the Syrians became servants to David and brought tribute. And the LORD gave victory to David wherever he went.
2SAM|8|7|And David took the shields of gold that were carried by the servants of Hadadezer and brought them to Jerusalem.
2SAM|8|8|And from Betah and from Berothai, cities of Hadadezer, King David took very much bronze.
2SAM|8|9|When Toi king of Hamath heard that David had defeated the whole army of Hadadezer,
2SAM|8|10|Toi sent his son Joram to King David, to ask about his health and to bless him because he had fought against Hadadezer and defeated him, for Hadadezer had often been at war with Toi. And Joram brought with him articles of silver, of gold, and of bronze.
2SAM|8|11|These also King David dedicated to the LORD, together with the silver and gold that he dedicated from all the nations he subdued,
2SAM|8|12|from Edom, Moab, the Ammonites, the Philistines, Amalek, and from the spoil of Hadadezer the son of Rehob, king of Zobah.
2SAM|8|13|And David made a name for himself when he returned from striking down 18,000 Edomites in the Valley of Salt.
2SAM|8|14|Then he put garrisons in Edom; throughout all Edom he put garrisons, and all the Edomites became David's servants. And the LORD gave victory to David wherever he went.
2SAM|8|15|So David reigned over all Israel. And David administered justice and equity to all his people.
2SAM|8|16|Joab the son of Zeruiah was over the army, and Jehoshaphat the son of Ahilud was recorder,
2SAM|8|17|and Zadok the son of Ahitub and Ahimelech the son of Abiathar were priests, and Seraiah was secretary,
2SAM|8|18|and Benaiah the son of Jehoiada was over the Cherethites and the Pelethites, and David's sons were priests.
2SAM|9|1|And David said, "Is there still anyone left of the house of Saul, that I may show him kindness for Jonathan's sake?"
2SAM|9|2|Now there was a servant of the house of Saul whose name was Ziba, and they called him to David. And the king said to him, "Are you Ziba?" And he said, "I am your servant."
2SAM|9|3|And the king said, "Is there not still someone of the house of Saul, that I may show the kindness of God to him?" Ziba said to the king, "There is still a son of Jonathan; he is crippled in his feet."
2SAM|9|4|The king said to him, "Where is he?" And Ziba said to the king, "He is in the house of Machir the son of Ammiel, at Lo-debar."
2SAM|9|5|Then King David sent and brought him from the house of Machir the son of Ammiel, at Lo-debar.
2SAM|9|6|And Mephibosheth the son of Jonathan, son of Saul, came to David and fell on his face and paid homage. And David said, "Mephibosheth!" And he answered, "Behold, I am your servant."
2SAM|9|7|And David said to him, "Do not fear, for I will show you kindness for the sake of your father Jonathan, and I will restore to you all the land of Saul your father, and you shall eat at my table always."
2SAM|9|8|And he paid homage and said, "What is your servant, that you should show regard for a dead dog such as I?"
2SAM|9|9|Then the king called Ziba, Saul's servant, and said to him, "All that belonged to Saul and to all his house I have given to your master's grandson.
2SAM|9|10|And you and your sons and your servants shall till the land for him and shall bring in the produce, that your master's grandson may have bread to eat. But Mephibosheth your master's grandson shall always eat at my table." Now Ziba had fifteen sons and twenty servants.
2SAM|9|11|Then Ziba said to the king, "According to all that my lord the king commands his servant, so will your servant do." So Mephibosheth ate at David's table, like one of the king's sons.
2SAM|9|12|And Mephibosheth had a young son, whose name was Mica. And all who lived in Ziba's house became Mephibosheth's servants.
2SAM|9|13|So Mephibosheth lived in Jerusalem, for he ate always at the king's table. Now he was lame in both his feet.
2SAM|10|1|After this the king of the Ammonites died, and Hanun his son reigned in his place.
2SAM|10|2|And David said, "I will deal loyally with Hanun the son of Nahash, as his father dealt loyally with me." So David sent by his servants to console him concerning his father. And David's servants came into the land of the Ammonites.
2SAM|10|3|But the princes of the Ammonites said to Hanun their lord, "Do you think, because David has sent comforters to you, that he is honoring your father? Has not David sent his servants to you to search the city and to spy it out and to overthrow it?"
2SAM|10|4|So Hanun took David's servants and shaved off half the beard of each and cut off their garments in the middle, at their hips, and sent them away.
2SAM|10|5|When it was told David, he sent to meet them, for the men were greatly ashamed. And the king said, "Remain at Jericho until your beards have grown and then return."
2SAM|10|6|When the Ammonites saw that they had become a stench to David, the Ammonites sent and hired the Syrians of Beth-rehob, and the Syrians of Zobah, 20,000 foot soldiers, and the king of Maacah with 1,000 men, and the men of Tob, 12,000 men.
2SAM|10|7|And when David heard of it, he sent Joab and all the host of the mighty men.
2SAM|10|8|And the Ammonites came out and drew up in battle array at the entrance of the gate, and the Syrians of Zobah and of Rehob and the men of Tob and Maacah were by themselves in the open country.
2SAM|10|9|When Joab saw that the battle was set against him both in front and in the rear, he chose some of the best men of Israel and arrayed them against the Syrians.
2SAM|10|10|The rest of his men he put in the charge of Abishai his brother, and he arrayed them against the Ammonites.
2SAM|10|11|And he said, "If the Syrians are too strong for me, then you shall help me, but if the Ammonites are too strong for you, then I will come and help you.
2SAM|10|12|Be of good courage, and let us be courageous for our people, and for the cities of our God, and may the LORD do what seems good to him."
2SAM|10|13|So Joab and the people who were with him drew near to battle against the Syrians, and they fled before him.
2SAM|10|14|And when the Ammonites saw that the Syrians fled, they likewise fled before Abishai and entered the city. Then Joab returned from fighting against the Ammonites and came to Jerusalem.
2SAM|10|15|But when the Syrians saw that they had been defeated by Israel, they gathered themselves together.
2SAM|10|16|And Hadadezer sent and brought out the Syrians who were beyond the Euphrates. They came to Helam, with Shobach the commander of the army of Hadadezer at their head.
2SAM|10|17|And when it was told David, he gathered all Israel together and crossed the Jordan and came to Helam. The Syrians arrayed themselves against David and fought with him.
2SAM|10|18|And the Syrians fled before Israel, and David killed of the Syrians the men of 700 chariots, and 40,000 horsemen, and wounded Shobach the commander of their army, so that he died there.
2SAM|10|19|And when all the kings who were servants of Hadadezer saw that they had been defeated by Israel, they made peace with Israel and became subject to them. So the Syrians were afraid to save the Ammonites anymore.
2SAM|11|1|In the spring of the year, the time when kings go out to battle, David sent Joab, and his servants with him, and all Israel. And they ravaged the Ammonites and besieged Rabbah. But David remained at Jerusalem.
2SAM|11|2|It happened, late one afternoon, when David arose from his couch and was walking on the roof of the king's house, that he saw from the roof a woman bathing; and the woman was very beautiful.
2SAM|11|3|And David sent and inquired about the woman. And one said, "Is not this Bathsheba, the daughter of Eliam, the wife of Uriah the Hittite?"
2SAM|11|4|So David sent messengers and took her, and she came to him, and he lay with her. (Now she had been purifying herself from her uncleanness.) Then she returned to her house.
2SAM|11|5|And the woman conceived, and she sent and told David, "I am pregnant."
2SAM|11|6|So David sent word to Joab, "Send me Uriah the Hittite." And Joab sent Uriah to David.
2SAM|11|7|When Uriah came to him, David asked how Joab was doing and how the people were doing and how the war was going.
2SAM|11|8|Then David said to Uriah, "Go down to your house and wash your feet." And Uriah went out of the king's house, and there followed him a present from the king.
2SAM|11|9|But Uriah slept at the door of the king's house with all the servants of his lord, and did not go down to his house.
2SAM|11|10|When they told David, "Uriah did not go down to his house," David said to Uriah, "Have you not come from a journey? Why did you not go down to your house?"
2SAM|11|11|Uriah said to David, "The ark and Israel and Judah dwell in booths, and my lord Joab and the servants of my lord are camping in the open field. Shall I then go to my house, to eat and to drink and to lie with my wife? As you live, and as your soul lives, I will not do this thing."
2SAM|11|12|Then David said to Uriah, "Remain here today also, and tomorrow I will send you back." So Uriah remained in Jerusalem that day and the next.
2SAM|11|13|And David invited him, and he ate in his presence and drank, so that he made him drunk. And in the evening he went out to lie on his couch with the servants of his lord, but he did not go down to his house.
2SAM|11|14|In the morning David wrote a letter to Joab and sent it by the hand of Uriah.
2SAM|11|15|In the letter he wrote, "Set Uriah in the forefront of the hardest fighting, and then draw back from him, that he may be struck down, and die."
2SAM|11|16|And as Joab was besieging the city, he assigned Uriah to the place where he knew there were valiant men.
2SAM|11|17|And the men of the city came out and fought with Joab, and some of the servants of David among the people fell. Uriah the Hittite also died.
2SAM|11|18|Then Joab sent and told David all the news about the fighting.
2SAM|11|19|And he instructed the messenger, "When you have finished telling all the news about the fighting to the king,
2SAM|11|20|then, if the king's anger rises, and if he says to you, 'Why did you go so near the city to fight? Did you not know that they would shoot from the wall?
2SAM|11|21|Who killed Abimelech the son of Jerubbesheth? Did not a woman cast an upper millstone on him from the wall, so that he died at Thebez? Why did you go so near the wall?' then you shall say, 'Your servant Uriah the Hittite is dead also.'"
2SAM|11|22|So the messenger went and came and told David all that Joab had sent him to tell.
2SAM|11|23|The messenger said to David, "The men gained an advantage over us and came out against us in the field, but we drove them back to the entrance of the gate.
2SAM|11|24|Then the archers shot at your servants from the wall. Some of the king's servants are dead, and your servant Uriah the Hittite is dead also."
2SAM|11|25|David said to the messenger, "Thus shall you say to Joab, 'Do not let this matter trouble you, for the sword devours now one and now another. Strengthen your attack against the city and overthrow it.' And encourage him."
2SAM|11|26|When the wife of Uriah heard that Uriah her husband was dead, she lamented over her husband.
2SAM|11|27|And when the mourning was over, David sent and brought her to his house, and she became his wife and bore him a son. But the thing that David had done displeased the LORD.
2SAM|12|1|And the LORD sent Nathan to David. He came to him and said to him, "There were two men in a certain city, the one rich and the other poor.
2SAM|12|2|The rich man had very many flocks and herds,
2SAM|12|3|but the poor man had nothing but one little ewe lamb, which he had bought. And he brought it up, and it grew up with him and with his children. It used to eat of his morsel and drink from his cup and lie in his arms, and it was like a daughter to him.
2SAM|12|4|Now there came a traveler to the rich man, and he was unwilling to take one of his own flock or herd to prepare for the guest who had come to him, but he took the poor man's lamb and prepared it for the man who had come to him."
2SAM|12|5|Then David's anger was greatly kindled against the man, and he said to Nathan, "As the LORD lives, the man who has done this deserves to die,
2SAM|12|6|and he shall restore the lamb fourfold, because he did this thing, and because he had no pity."
2SAM|12|7|Nathan said to David, "You are the man! Thus says the LORD, the God of Israel, 'I anointed you king over Israel, and I delivered you out of the hand of Saul.
2SAM|12|8|And I gave you your master's house and your master's wives into your arms and gave you the house of Israel and of Judah. And if this were too little, I would add to you as much more.
2SAM|12|9|Why have you despised the word of the LORD, to do what is evil in his sight? You have struck down Uriah the Hittite with the sword and have taken his wife to be your wife and have killed him with the sword of the Ammonites.
2SAM|12|10|Now therefore the sword shall never depart from your house, because you have despised me and have taken the wife of Uriah the Hittite to be your wife.'
2SAM|12|11|Thus says the LORD, 'Behold, I will raise up evil against you out of your own house. And I will take your wives before your eyes and give them to your neighbor, and he shall lie with your wives in the sight of this sun.
2SAM|12|12|For you did it secretly, but I will do this thing before all Israel and before the sun.'"
2SAM|12|13|David said to Nathan, "I have sinned against the LORD." And Nathan said to David, "The LORD also has put away your sin; you shall not die.
2SAM|12|14|Nevertheless, because by this deed you have utterly scorned the LORD, the child who is born to you shall die."
2SAM|12|15|Then Nathan went to his house. And the LORD afflicted the child that Uriah's wife bore to David, and he became sick.
2SAM|12|16|David therefore sought God on behalf of the child. And David fasted and went in and lay all night on the ground.
2SAM|12|17|And the elders of his house stood beside him, to raise him from the ground, but he would not, nor did he eat food with them.
2SAM|12|18|On the seventh day the child died. And the servants of David were afraid to tell him that the child was dead, for they said, "Behold, while the child was yet alive, we spoke to him, and he did not listen to us. How then can we say to him the child is dead? He may do himself some harm."
2SAM|12|19|But when David saw that his servants were whispering together, David understood that the child was dead. And David said to his servants, "Is the child dead?" They said, "He is dead."
2SAM|12|20|Then David arose from the earth and washed and anointed himself and changed his clothes. And he went into the house of the LORD and worshiped. He then went to his own house. And when he asked, they set food before him, and he ate.
2SAM|12|21|Then his servants said to him, "What is this thing that you have done? You fasted and wept for the child while he was alive; but when the child died, you arose and ate food."
2SAM|12|22|He said, "While the child was still alive, I fasted and wept, for I said, 'Who knows whether the LORD will be gracious to me, that the child may live?'
2SAM|12|23|But now he is dead. Why should I fast? Can I bring him back again? I shall go to him, but he will not return to me."
2SAM|12|24|Then David comforted his wife, Bathsheba, and went in to her and lay with her, and she bore a son, and he called his name Solomon. And the LORD loved him
2SAM|12|25|and sent a message by Nathan the prophet. So he called his name Jedidiah, because of the LORD.
2SAM|12|26|Now Joab fought against Rabbah of the Ammonites and took the royal city.
2SAM|12|27|And Joab sent messengers to David and said, "I have fought against Rabbah; moreover, I have taken the city of waters.
2SAM|12|28|Now then gather the rest of the people together and encamp against the city and take it, lest I take the city and it be called by my name."
2SAM|12|29|So David gathered all the people together and went to Rabbah and fought against it and took it.
2SAM|12|30|And he took the crown of their king from his head. The weight of it was a talent of gold, and in it was a precious stone, and it was placed on David's head. And he brought out the spoil of the city, a very great amount.
2SAM|12|31|And he brought out the people who were in it and set them to labor with saws and iron picks and iron axes and made them toil at the brick kilns. And thus he did to all the cities of the Ammonites. Then David and all the people returned to Jerusalem.
2SAM|13|1|Now Absalom, David's son, had a beautiful sister, whose name was Tamar. And after a time Amnon, David's son, loved her.
2SAM|13|2|And Amnon was so tormented that he made himself ill because of his sister Tamar, for she was a virgin, and it seemed impossible to Amnon to do anything to her.
2SAM|13|3|But Amnon had a friend, whose name was Jonadab, the son of Shimeah, David's brother. And Jonadab was a very crafty man.
2SAM|13|4|And he said to him, "O son of the king, why are you so haggard morning after morning? Will you not tell me?" Amnon said to him, "I love Tamar, my brother Absalom's sister."
2SAM|13|5|Jonadab said to him, "Lie down on your bed and pretend to be ill. And when your father comes to see you, say to him, 'Let my sister Tamar come and give me bread to eat, and prepare the food in my sight, that I may see it and eat it from her hand.'"
2SAM|13|6|So Amnon lay down and pretended to be ill. And when the king came to see him, Amnon said to the king, "Please let my sister Tamar come and make a couple of cakes in my sight, that I may eat from her hand."
2SAM|13|7|Then David sent home to Tamar, saying, "Go to your brother Amnon's house and prepare food for him."
2SAM|13|8|So Tamar went to her brother Amnon's house, where he was lying down. And she took dough and kneaded it and made cakes in his sight and baked the cakes.
2SAM|13|9|And she took the pan and emptied it out before him, but he refused to eat. And Amnon said, "Send out everyone from me." So everyone went out from him.
2SAM|13|10|Then Amnon said to Tamar, "Bring the food into the chamber, that I may eat from your hand." And Tamar took the cakes she had made and brought them into the chamber to Amnon her brother.
2SAM|13|11|But when she brought them near him to eat, he took hold of her and said to her, "Come, lie with me, my sister."
2SAM|13|12|She answered him, "No, my brother, do not violate me, for such a thing is not done in Israel; do not do this outrageous thing.
2SAM|13|13|As for me, where could I carry my shame? And as for you, you would be as one of the outrageous fools in Israel. Now therefore, please speak to the king, for he will not withhold me from you."
2SAM|13|14|But he would not listen to her, and being stronger than she, he violated her and lay with her.
2SAM|13|15|Then Amnon hated her with very great hatred, so that the hatred with which he hated her was greater than the love with which he had loved her. And Amnon said to her, "Get up! Go!"
2SAM|13|16|But she said to him, "No, my brother, for this wrong in sending me away is greater than the other that you did to me." But he would not listen to her.
2SAM|13|17|He called the young man who served him and said, "Put this woman out of my presence and bolt the door after her."
2SAM|13|18|Now she was wearing a long robe with sleeves, for thus were the virgin daughters of the king dressed. So his servant put her out and bolted the door after her.
2SAM|13|19|And Tamar put ashes on her head and tore the long robe that she wore. And she laid her hand on her head and went away, crying aloud as she went.
2SAM|13|20|And her brother Absalom said to her, "Has Amnon your brother been with you? Now hold your peace, my sister. He is your brother; do not take this to heart." So Tamar lived, a desolate woman, in her brother Absalom's house.
2SAM|13|21|When King David heard of all these things, he was very angry.
2SAM|13|22|But Absalom spoke to Amnon neither good nor bad, for Absalom hated Amnon, because he had violated his sister Tamar.
2SAM|13|23|After two full years Absalom had sheepshearers at Baal-hazor, which is near Ephraim, and Absalom invited all the king's sons.
2SAM|13|24|And Absalom came to the king and said, "Behold, your servant has sheepshearers. Please let the king and his servants go with your servant."
2SAM|13|25|But the king said to Absalom, "No, my son, let us not all go, lest we be burdensome to you." He pressed him, but he would not go but gave him his blessing.
2SAM|13|26|Then Absalom said, "If not, please let my brother Amnon go with us." And the king said to him, "Why should he go with you?"
2SAM|13|27|But Absalom pressed him until he let Amnon and all the king's sons go with him.
2SAM|13|28|Then Absalom commanded his servants, "Mark when Amnon's heart is merry with wine, and when I say to you, 'Strike Amnon,' then kill him. Do not fear; have I not commanded you? Be courageous and be valiant."
2SAM|13|29|So the servants of Absalom did to Amnon as Absalom had commanded. Then all the king's sons arose, and each mounted his mule and fled.
2SAM|13|30|While they were on the way, news came to David, "Absalom has struck down all the king's sons, and not one of them is left."
2SAM|13|31|Then the king arose and tore his garments and lay on the earth. And all his servants who were standing by tore their garments.
2SAM|13|32|But Jonadab the son of Shimeah, David's brother, said, "Let not my lord suppose that they have killed all the young men the king's sons, for Amnon alone is dead. For by the command of Absalom this has been determined from the day he violated his sister Tamar.
2SAM|13|33|Now therefore let not my lord the king so take it to heart as to suppose that all the king's sons are dead, for Amnon alone is dead."
2SAM|13|34|But Absalom fled. And the young man who kept the watch lifted up his eyes and looked, and behold, many people were coming from the road behind him by the side of the mountain.
2SAM|13|35|And Jonadab said to the king, "Behold, the king's sons have come; as your servant said, so it has come about."
2SAM|13|36|And as soon as he had finished speaking, behold, the king's sons came and lifted up their voice and wept. And the king also and all his servants wept very bitterly.
2SAM|13|37|But Absalom fled and went to Talmai the son of Ammihud, king of Geshur. And David mourned for his son day after day.
2SAM|13|38|So Absalom fled and went to Geshur, and was there three years.
2SAM|13|39|And the spirit of the king longed to go out to Absalom, because he was comforted about Amnon, since he was dead.
2SAM|14|1|Now Joab the son of Zeruiah knew that the king's heart went out to Absalom.
2SAM|14|2|And Joab sent to Tekoa and brought from there a wise woman and said to her, "Pretend to be a mourner and put on mourning garments. Do not anoint yourself with oil, but behave like a woman who has been mourning many days for the dead.
2SAM|14|3|Go to the king and speak thus to him." So Joab put the words in her mouth.
2SAM|14|4|When the woman of Tekoa came to the king, she fell on her face to the ground and paid homage and said, "Save me, O king."
2SAM|14|5|And the king said to her, "What is your trouble?" She answered, "Alas, I am a widow; my husband is dead.
2SAM|14|6|And your servant had two sons, and they quarreled with one another in the field. There was no one to separate them, and one struck the other and killed him.
2SAM|14|7|And now the whole clan has risen against your servant, and they say, 'Give up the man who struck his brother, that we may put him to death for the life of his brother whom he killed.' And so they would destroy the heir also. Thus they would quench my coal that is left and leave to my husband neither name nor remnant on the face of the earth."
2SAM|14|8|Then the king said to the woman, "Go to your house, and I will give orders concerning you."
2SAM|14|9|And the woman of Tekoa said to the king, "On me be the guilt, my lord the king, and on my father's house; let the king and his throne be guiltless."
2SAM|14|10|The king said, "If anyone says anything to you, bring him to me, and he shall never touch you again."
2SAM|14|11|Then she said, "Please let the king invoke the LORD your God, that the avenger of blood kill no more, and my son be not destroyed." He said, "As the LORD lives, not one hair of your son shall fall to the ground."
2SAM|14|12|Then the woman said, "Please let your servant speak a word to my lord the king." He said, "Speak."
2SAM|14|13|And the woman said, "Why then have you planned such a thing against the people of God? For in giving this decision the king convicts himself, inasmuch as the king does not bring his banished one home again.
2SAM|14|14|We must all die; we are like water spilled on the ground, which cannot be gathered up again. But God will not take away life, and he devises means so that the banished one will not remain an outcast.
2SAM|14|15|Now I have come to say this to my lord the king because the people have made me afraid, and your servant thought, 'I will speak to the king; it may be that the king will perform the request of his servant.
2SAM|14|16|For the king will hear and deliver his servant from the hand of the man who would destroy me and my son together from the heritage of God.'
2SAM|14|17|And your servant thought, 'The word of my lord the king will set me at rest,' for my lord the king is like the angel of God to discern good and evil. The LORD your God be with you!"
2SAM|14|18|Then the king answered the woman, "Do not hide from me anything I ask you." And the woman said, "Let my lord the king speak."
2SAM|14|19|The king said, "Is the hand of Joab with you in all this?" The woman answered and said, "As surely as you live, my lord the king, one cannot turn to the right hand or to the left from anything that my lord the king has said. It was your servant Joab who commanded me; it was he who put all these words in the mouth of your servant.
2SAM|14|20|In order to change the course of things your servant Joab did this. But my lord has wisdom like the wisdom of the angel of God to know all things that are on the earth."
2SAM|14|21|Then the king said to Joab, "Behold now, I grant this; go, bring back the young man Absalom."
2SAM|14|22|And Joab fell on his face to the ground and paid homage and blessed the king. And Joab said, "Today your servant knows that I have found favor in your sight, my lord the king, in that the king has granted the request of his servant."
2SAM|14|23|So Joab arose and went to Geshur and brought Absalom to Jerusalem.
2SAM|14|24|And the king said, "Let him dwell apart in his own house; he is not to come into my presence." So Absalom lived apart in his own house and did not come into the king's presence.
2SAM|14|25|Now in all Israel there was no one so much to be praised for his handsome appearance as Absalom. From the sole of his foot to the crown of his head there was no blemish in him.
2SAM|14|26|And when he cut the hair of his head (for at the end of every year he used to cut it; when it was heavy on him, he cut it), he weighed the hair of his head, two hundred shekels by the king's weight.
2SAM|14|27|There were born to Absalom three sons, and one daughter whose name was Tamar. She was a beautiful woman.
2SAM|14|28|So Absalom lived two full years in Jerusalem, without coming into the king's presence.
2SAM|14|29|Then Absalom sent for Joab, to send him to the king, but Joab would not come to him. And he sent a second time, but Joab would not come.
2SAM|14|30|Then he said to his servants, "See, Joab's field is next to mine, and he has barley there; go and set it on fire." So Absalom's servants set the field on fire.
2SAM|14|31|Then Joab arose and went to Absalom at his house and said to him, "Why have your servants set my field on fire?"
2SAM|14|32|Absalom answered Joab, "Behold, I sent word to you, 'Come here, that I may send you to the king, to ask, "Why have I come from Geshur? It would be better for me to be there still." Now therefore let me go into the presence of the king, and if there is guilt in me, let him put me to death.'"
2SAM|14|33|Then Joab went to the king and told him, and he summoned Absalom. So he came to the king and bowed himself on his face to the ground before the king, and the king kissed Absalom.
2SAM|15|1|After this Absalom got himself a chariot and horses, and fifty men to run before him.
2SAM|15|2|And Absalom used to rise early and stand beside the way of the gate. And when any man had a dispute to come before the king for judgment, Absalom would call to him and say, "From what city are you?" And when he said, "Your servant is of such and such a tribe in Israel,"
2SAM|15|3|Absalom would say to him, "See, your claims are good and right, but there is no man designated by the king to hear you."
2SAM|15|4|Then Absalom would say, "Oh that I were judge in the land! Then every man with a dispute or cause might come to me, and I would give him justice."
2SAM|15|5|And whenever a man came near to pay homage to him, he would put out his hand and take hold of him and kiss him.
2SAM|15|6|Thus Absalom did to all of Israel who came to the king for judgment. So Absalom stole the hearts of the men of Israel.
2SAM|15|7|And at the end of four years Absalom said to the king, "Please let me go and pay my vow, which I have vowed to the LORD, in Hebron.
2SAM|15|8|For your servant vowed a vow while I lived at Geshur in Aram, saying, 'If the LORD will indeed bring me back to Jerusalem, then I will offer worship to the LORD.'"
2SAM|15|9|The king said to him, "Go in peace." So he arose and went to Hebron.
2SAM|15|10|But Absalom sent secret messengers throughout all the tribes of Israel, saying, "As soon as you hear the sound of the trumpet, then say, 'Absalom is king at Hebron!'"
2SAM|15|11|With Absalom went two hundred men from Jerusalem who were invited guests, and they went in their innocence and knew nothing.
2SAM|15|12|And while Absalom was offering the sacrifices, he sent for Ahithophel the Gilonite, David's counselor, from his city Giloh. And the conspiracy grew strong, and the people with Absalom kept increasing.
2SAM|15|13|And a messenger came to David, saying, "The hearts of the men of Israel have gone after Absalom."
2SAM|15|14|Then David said to all his servants who were with him at Jerusalem, "Arise, and let us flee, or else there will be no escape for us from Absalom. Go quickly, lest he overtake us quickly and bring down ruin on us and strike the city with the edge of the sword."
2SAM|15|15|And the king's servants said to the king, "Behold, your servants are ready to do whatever my lord the king decides."
2SAM|15|16|So the king went out, and all his household after him. And the king left ten concubines to keep the house.
2SAM|15|17|And the king went out, and all the people after him. And they halted at the last house.
2SAM|15|18|And all his servants passed by him, and all the Cherethites, and all the Pelethites, and all the six hundred Gittites who had followed him from Gath, passed on before the king.
2SAM|15|19|Then the king said to Ittai the Gittite, "Why do you also go with us? Go back and stay with the king, for you are a foreigner and also an exile from your home.
2SAM|15|20|You came only yesterday, and shall I today make you wander about with us, since I go I know not where? Go back and take your brothers with you, and may the LORD show steadfast love and faithfulness to you."
2SAM|15|21|But Ittai answered the king, "As the LORD lives, and as my lord the king lives, wherever my lord the king shall be, whether for death or for life, there also will your servant be."
2SAM|15|22|And David said to Ittai, "Go then, pass on." So Ittai the Gittite passed on with all his men and all the little ones who were with him.
2SAM|15|23|And all the land wept aloud as all the people passed by, and the king crossed the brook Kidron, and all the people passed on toward the wilderness.
2SAM|15|24|And Abiathar came up, and behold, Zadok came also with all the Levites, bearing the ark of the covenant of God. And they set down the ark of God until the people had all passed out of the city.
2SAM|15|25|Then the king said to Zadok, "Carry the ark of God back into the city. If I find favor in the eyes of the LORD, he will bring me back and let me see both it and his dwelling place.
2SAM|15|26|But if he says, 'I have no pleasure in you,' behold, here I am, let him do to me what seems good to him."
2SAM|15|27|The king also said to Zadok the priest, "Are you not a seer? Go back to the city in peace, with your two sons, Ahimaaz your son, and Jonathan the son of Abiathar.
2SAM|15|28|See, I will wait at the fords of the wilderness until word comes from you to inform me."
2SAM|15|29|So Zadok and Abiathar carried the ark of God back to Jerusalem, and they remained there.
2SAM|15|30|But David went up the ascent of the Mount of Olives, weeping as he went, barefoot and with his head covered. And all the people who were with him covered their heads, and they went up, weeping as they went.
2SAM|15|31|And it was told David, "Ahithophel is among the conspirators with Absalom." And David said, "O LORD, please turn the counsel of Ahithophel into foolishness."
2SAM|15|32|While David was coming to the summit, where God was worshiped, behold, Hushai the Archite came to meet him with his coat torn and dirt on his head.
2SAM|15|33|David said to him, "If you go on with me, you will be a burden to me.
2SAM|15|34|But if you return to the city and say to Absalom, 'I will be your servant, O king; as I have been your father's servant in time past, so now I will be your servant,' then you will defeat for me the counsel of Ahithophel.
2SAM|15|35|Are not Zadok and Abiathar the priests with you there? So whatever you hear from the king's house, tell it to Zadok and Abiathar the priests.
2SAM|15|36|Behold, their two sons are with them there, Ahimaaz, Zadok's son, and Jonathan, Abiathar's son, and by them you shall send to me everything you hear."
2SAM|15|37|So Hushai, David's friend, came into the city, just as Absalom was entering Jerusalem.
2SAM|16|1|When David had passed a little beyond the summit, Ziba the servant of Mephibosheth met him, with a couple of donkeys saddled, bearing two hundred loaves of bread, a hundred bunches of raisins, a hundred of summer fruits, and a skin of wine.
2SAM|16|2|And the king said to Ziba, "Why have you brought these?" Ziba answered, "The donkeys are for the king's household to ride on, the bread and summer fruit for the young men to eat, and the wine for those who faint in the wilderness to drink."
2SAM|16|3|And the king said, "And where is your master's son?" Ziba said to the king, "Behold, he remains in Jerusalem, for he said, 'Today the house of Israel will give me back the kingdom of my father.'"
2SAM|16|4|Then the king said to Ziba, "Behold, all that belonged to Mephibosheth is now yours." And Ziba said, "I pay homage; let me ever find favor in your sight, my lord the king."
2SAM|16|5|When King David came to Bahurim, there came out a man of the family of the house of Saul, whose name was Shimei, the son of Gera, and as he came he cursed continually.
2SAM|16|6|And he threw stones at David and at all the servants of King David, and all the people and all the mighty men were on his right hand and on his left.
2SAM|16|7|And Shimei said as he cursed, "Get out, get out, you man of blood, you worthless man!
2SAM|16|8|The LORD has avenged on you all the blood of the house of Saul, in whose place you have reigned, and the LORD has given the kingdom into the hand of your son Absalom. See, your evil is on you, for you are a man of blood."
2SAM|16|9|Then Abishai the son of Zeruiah said to the king, "Why should this dead dog curse my lord the king? Let me go over and take off his head."
2SAM|16|10|But the king said, "What have I to do with you, you sons of Zeruiah? If he is cursing because the LORD has said to him, 'Curse David,' who then shall say, 'Why have you done so?'"
2SAM|16|11|And David said to Abishai and to all his servants, "Behold, my own son seeks my life; how much more now may this Benjaminite! Leave him alone, and let him curse, for the LORD has told him to.
2SAM|16|12|It may be that the LORD will look on the wrong done to me, and that the LORD will repay me with good for his cursing today."
2SAM|16|13|So David and his men went on the road, while Shimei went along on the hillside opposite him and cursed as he went and threw stones at him and flung dust.
2SAM|16|14|And the king, and all the people who were with him, arrived weary at the Jordan. And there he refreshed himself.
2SAM|16|15|Now Absalom and all the people, the men of Israel, came to Jerusalem, and Ahithophel with him.
2SAM|16|16|And when Hushai the Archite, David's friend, came to Absalom, Hushai said to Absalom, "Long live the king! Long live the king!"
2SAM|16|17|And Absalom said to Hushai, "Is this your loyalty to your friend? Why did you not go with your friend?"
2SAM|16|18|And Hushai said to Absalom, "No, for whom the LORD and this people and all the men of Israel have chosen, his I will be, and with him I will remain.
2SAM|16|19|And again, whom should I serve? Should it not be his son? As I have served your father, so I will serve you."
2SAM|16|20|Then Absalom said to Ahithophel, "Give your counsel. What shall we do?"
2SAM|16|21|Ahithophel said to Absalom, "Go in to your father's concubines, whom he has left to keep the house, and all Israel will hear that you have made yourself a stench to your father, and the hands of all who are with you will be strengthened."
2SAM|16|22|So they pitched a tent for Absalom on the roof. And Absalom went in to his father's concubines in the sight of all Israel.
2SAM|16|23|Now in those days the counsel that Ahithophel gave was as if one consulted the word of God; so was all the counsel of Ahithophel esteemed, both by David and by Absalom.
2SAM|17|1|Moreover, Ahithophel said to Absalom, "Let me choose twelve thousand men, and I will arise and pursue David tonight.
2SAM|17|2|I will come upon him while he is weary and discouraged and throw him into a panic, and all the people who are with him will flee. I will strike down only the king,
2SAM|17|3|and I will bring all the people back to you as a bride comes home to her husband. You seek the life of only one man, and all the people will be at peace."
2SAM|17|4|And the advice seemed right in the eyes of Absalom and all the elders of Israel.
2SAM|17|5|Then Absalom said, "Call Hushai the Archite also, and let us hear what he has to say."
2SAM|17|6|And when Hushai came to Absalom, Absalom said to him, "Thus has Ahithophel spoken; shall we do as he says? If not, you speak."
2SAM|17|7|Then Hushai said to Absalom, "This time the counsel that Ahithophel has given is not good."
2SAM|17|8|Hushai said, "You know that your father and his men are mighty men, and that they are enraged, like a bear robbed of her cubs in the field. Besides, your father is expert in war; he will not spend the night with the people.
2SAM|17|9|Behold, even now he has hidden himself in one of the pits or in some other place. And as soon as some of the people fall at the first attack, whoever hears it will say, 'There has been a slaughter among the people who follow Absalom.'
2SAM|17|10|Then even the valiant man, whose heart is like the heart of a lion, will utterly melt with fear, for all Israel knows that your father is a mighty man, and that those who are with him are valiant men.
2SAM|17|11|But my counsel is that all Israel be gathered to you, from Dan to Beersheba, as the sand by the sea for multitude, and that you go to battle in person.
2SAM|17|12|So we shall come upon him in some place where he is to be found, and we shall light upon him as the dew falls on the ground, and of him and all the men with him not one will be left.
2SAM|17|13|If he withdraws into a city, then all Israel will bring ropes to that city, and we shall drag it into the valley, until not even a pebble is to be found there."
2SAM|17|14|And Absalom and all the men of Israel said, "The counsel of Hushai the Archite is better than the counsel of Ahithophel." For the LORD had ordained to defeat the good counsel of Ahithophel, so that the LORD might bring harm upon Absalom.
2SAM|17|15|Then Hushai said to Zadok and Abiathar the priests, "Thus and so did Ahithophel counsel Absalom and the elders of Israel, and thus and so have I counseled.
2SAM|17|16|Now therefore send quickly and tell David, 'Do not stay tonight at the fords of the wilderness, but by all means pass over, lest the king and all the people who are with him be swallowed up.'"
2SAM|17|17|Now Jonathan and Ahimaaz were waiting at En-rogel. A female servant was to go and tell them, and they were to go and tell King David, for they were not to be seen entering the city.
2SAM|17|18|But a young man saw them and told Absalom. So both of them went away quickly and came to the house of a man at Bahurim, who had a well in his courtyard. And they went down into it.
2SAM|17|19|And the woman took and spread a covering over the well's mouth and scattered grain on it, and nothing was known of it.
2SAM|17|20|When Absalom's servants came to the woman at the house, they said, "Where are Ahimaaz and Jonathan?" And the woman said to them, "They have gone over the brook of water." And when they had sought and could not find them, they returned to Jerusalem.
2SAM|17|21|After they had gone, the men came up out of the well, and went and told King David. They said to David, "Arise, and go quickly over the water, for thus and so has Ahithophel counseled against you."
2SAM|17|22|Then David arose, and all the people who were with him, and they crossed the Jordan. By daybreak not one was left who had not crossed the Jordan.
2SAM|17|23|When Ahithophel saw that his counsel was not followed, he saddled his donkey and went off home to his own city. He set his house in order and hanged himself, and he died and was buried in the tomb of his father.
2SAM|17|24|Then David came to Mahanaim. And Absalom crossed the Jordan with all the men of Israel.
2SAM|17|25|Now Absalom had set Amasa over the army instead of Joab. Amasa was the son of a man named Ithra the Ishmaelite, who had married Abigal the daughter of Nahash, sister of Zeruiah, Joab's mother.
2SAM|17|26|And Israel and Absalom encamped in the land of Gilead.
2SAM|17|27|When David came to Mahanaim, Shobi the son of Nahash from Rabbah of the Ammonites, and Machir the son of Ammiel from Lo-debar, and Barzillai the Gileadite from Rogelim,
2SAM|17|28|brought beds, basins, and earthen vessels, wheat, barley, flour, parched grain, beans and lentils,
2SAM|17|29|honey and curds and sheep and cheese from the herd, for David and the people with him to eat, for they said, "The people are hungry and weary and thirsty in the wilderness."
2SAM|18|1|Then David mustered the men who were with him and set over them commanders of thousands and commanders of hundreds.
2SAM|18|2|And David sent out the army, one third under the command of Joab, one third under the command of Abishai the son of Zeruiah, Joab's brother, and one third under the command of Ittai the Gittite. And the king said to the men, "I myself will also go out with you."
2SAM|18|3|But the men said, "You shall not go out. For if we flee, they will not care about us. If half of us die, they will not care about us. But you are worth ten thousand of us. Therefore it is better that you send us help from the city."
2SAM|18|4|The king said to them, "Whatever seems best to you I will do." So the king stood at the side of the gate, while all the army marched out by hundreds and by thousands.
2SAM|18|5|And the king ordered Joab and Abishai and Ittai, "Deal gently for my sake with the young man Absalom." And all the people heard when the king gave orders to all the commanders about Absalom.
2SAM|18|6|So the army went out into the field against Israel, and the battle was fought in the forest of Ephraim.
2SAM|18|7|And the men of Israel were defeated there by the servants of David, and the loss there was great on that day, twenty thousand men.
2SAM|18|8|The battle spread over the face of all the country, and the forest devoured more people that day than the sword.
2SAM|18|9|And Absalom happened to meet the servants of David. Absalom was riding on his mule, and the mule went under the thick branches of a great terebinth, and his head caught fast in the oak, and he was suspended between heaven and earth, while the mule that was under him went on.
2SAM|18|10|And a certain man saw it and told Joab, "Behold, I saw Absalom hanging in an oak."
2SAM|18|11|Joab said to the man who told him, "What, you saw him! Why then did you not strike him there to the ground? I would have been glad to give you ten pieces of silver and a belt."
2SAM|18|12|But the man said to Joab, "Even if I felt in my hand the weight of a thousand pieces of silver, I would not reach out my hand against the king's son, for in our hearing the king commanded you and Abishai and Ittai, 'For my sake protect the young man Absalom.'
2SAM|18|13|On the other hand, if I had dealt treacherously against his life (and there is nothing hidden from the king), then you yourself would have stood aloof."
2SAM|18|14|Joab said, "I will not waste time like this with you." And he took three javelins in his hand and thrust them into the heart of Absalom while he was still alive in the oak.
2SAM|18|15|And ten young men, Joab's armor-bearers, surrounded Absalom and struck him and killed him.
2SAM|18|16|Then Joab blew the trumpet, and the troops came back from pursuing Israel, for Joab restrained them.
2SAM|18|17|And they took Absalom and threw him into a great pit in the forest and raised over him a very great heap of stones. And all Israel fled every one to his own home.
2SAM|18|18|Now Absalom in his lifetime had taken and set up for himself the pillar that is in the King's Valley, for he said, "I have no son to keep my name in remembrance." He called the pillar after his own name, and it is called Absalom's monument to this day.
2SAM|18|19|Then Ahimaaz the son of Zadok said, "Let me run and carry news to the king that the LORD has delivered him from the hand of his enemies."
2SAM|18|20|And Joab said to him, "You are not to carry news today. You may carry news another day, but today you shall carry no news, because the king's son is dead."
2SAM|18|21|Then Joab said to the Cushite, "Go, tell the king what you have seen." The Cushite bowed before Joab, and ran.
2SAM|18|22|Then Ahimaaz the son of Zadok said again to Joab, "Come what may, let me also run after the Cushite." And Joab said, "Why will you run, my son, seeing that you will have no reward for the news?"
2SAM|18|23|"Come what may," he said, "I will run." So he said to him, "Run." Then Ahimaaz ran by the way of the plain, and outran the Cushite.
2SAM|18|24|Now David was sitting between the two gates, and the watchman went up to the roof of the gate by the wall, and when he lifted up his eyes and looked, he saw a man running alone.
2SAM|18|25|The watchman called out and told the king. And the king said, "If he is alone, there is news in his mouth." And he drew nearer and nearer.
2SAM|18|26|The watchman saw another man running. And the watchman called to the gate and said, "See, another man running alone!" The king said, "He also brings news."
2SAM|18|27|The watchman said, "I think the running of the first is like the running of Ahimaaz the son of Zadok." And the king said, "He is a good man and comes with good news."
2SAM|18|28|Then Ahimaaz cried out to the king, "All is well." And he bowed before the king with his face to the earth and said, "Blessed be the LORD your God, who has delivered up the men who raised their hand against my lord the king."
2SAM|18|29|And the king said, "Is it well with the young man Absalom?" Ahimaaz answered, "When Joab sent the king's servant, your servant, I saw a great commotion, but I do not know what it was."
2SAM|18|30|And the king said, "Turn aside and stand here." So he turned aside and stood still.
2SAM|18|31|And behold, the Cushite came, and the Cushite said, "Good news for my lord the king! For the LORD has delivered you this day from the hand of all who rose up against you."
2SAM|18|32|The king said to the Cushite, "Is it well with the young man Absalom?" And the Cushite answered, "May the enemies of my lord the king and all who rise up against you for evil be like that young man."
2SAM|18|33|And the king was deeply moved and went up to the chamber over the gate and wept. And as he went, he said, "O my son Absalom, my son, my son Absalom! Would I had died instead of you, O Absalom, my son, my son!"
2SAM|19|1|It was told Joab, "Behold, the king is weeping and mourning for Absalom."
2SAM|19|2|So the victory that day was turned into mourning for all the people, for the people heard that day, "The king is grieving for his son."
2SAM|19|3|And the people stole into the city that day as people steal in who are ashamed when they flee in battle.
2SAM|19|4|The king covered his face, and the king cried with a loud voice, "O my son Absalom, O Absalom, my son, my son!"
2SAM|19|5|Then Joab came into the house to the king and said, "You have today covered with shame the faces of all your servants, who have this day saved your life and the lives of your sons and your daughters and the lives of your wives and your concubines,
2SAM|19|6|because you love those who hate you and hate those who love you. For you have made it clear today that commanders and servants are nothing to you, for today I know that if Absalom were alive and all of us were dead today, then you would be pleased.
2SAM|19|7|Now therefore arise, go out and speak kindly to your servants, for I swear by the LORD, if you do not go, not a man will stay with you this night, and this will be worse for you than all the evil that has come upon you from your youth until now."
2SAM|19|8|Then the king arose and took his seat in the gate. And the people were all told, "Behold, the king is sitting in the gate." And all the people came before the king. Now Israel had fled every man to his own home.
2SAM|19|9|And all the people were arguing throughout all the tribes of Israel, saying, "The king delivered us from the hand of our enemies and saved us from the hand of the Philistines, and now he has fled out of the land from Absalom.
2SAM|19|10|But Absalom, whom we anointed over us, is dead in battle. Now therefore why do you say nothing about bringing the king back?"
2SAM|19|11|And King David sent this message to Zadok and Abiathar the priests, "Say to the elders of Judah, 'Why should you be the last to bring the king back to his house, when the word of all Israel has come to the king?
2SAM|19|12|You are my brothers; you are my bone and my flesh. Why then should you be the last to bring back the king?'
2SAM|19|13|And say to Amasa, 'Are you not my bone and my flesh? God do so to me and more also, if you are not commander of my army from now on in place of Joab.'"
2SAM|19|14|And he swayed the heart of all the men of Judah as one man, so that they sent word to the king, "Return, both you and all your servants."
2SAM|19|15|So the king came back to the Jordan, and Judah came to Gilgal to meet the king and to bring the king over the Jordan.
2SAM|19|16|And Shimei the son of Gera, the Benjaminite, from Bahurim, hurried to come down with the men of Judah to meet King David.
2SAM|19|17|And with him were a thousand men from Benjamin. And Ziba the servant of the house of Saul, with his fifteen sons and his twenty servants, rushed down to the Jordan before the king,
2SAM|19|18|and they crossed the ford to bring over the king's household and to do his pleasure. And Shimei the son of Gera fell down before the king, as he was about to cross the Jordan,
2SAM|19|19|and said to the king, "Let not my lord hold me guilty or remember how your servant did wrong on the day my lord the king left Jerusalem. Do not let the king take it to heart.
2SAM|19|20|For your servant knows that I have sinned. Therefore, behold, I have come this day, the first of all the house of Joseph to come down to meet my lord the king."
2SAM|19|21|Abishai the son of Zeruiah answered, "Shall not Shimei be put to death for this, because he cursed the LORD's anointed?"
2SAM|19|22|But David said, "What have I to do with you, you sons of Zeruiah, that you should this day be as an adversary to me? Shall anyone be put to death in Israel this day? For do I not know that I am this day king over Israel?"
2SAM|19|23|And the king said to Shimei, "You shall not die." And the king gave him his oath.
2SAM|19|24|And Mephibosheth the son of Saul came down to meet the king. He had neither taken care of his feet nor trimmed his beard nor washed his clothes, from the day the king departed until the day he came back in safety.
2SAM|19|25|And when he came to Jerusalem to meet the king, the king said to him, "Why did you not go with me, Mephibosheth?"
2SAM|19|26|He answered, "My lord, O king, my servant deceived me, for your servant said to him, 'I will saddle a donkey for myself, that I may ride on it and go with the king.' For your servant is lame.
2SAM|19|27|He has slandered your servant to my lord the king. But my lord the king is like the angel of God; do therefore what seems good to you.
2SAM|19|28|For all my father's house were but men doomed to death before my lord the king, but you set your servant among those who eat at your table. What further right have I, then, to cry to the king?"
2SAM|19|29|And the king said to him, "Why speak any more of your affairs? I have decided: you and Ziba shall divide the land."
2SAM|19|30|And Mephibosheth said to the king, "Oh, let him take it all, since my lord the king has come safely home."
2SAM|19|31|Now Barzillai the Gileadite had come down from Rogelim, and he went on with the king to the Jordan, to escort him over the Jordan.
2SAM|19|32|Barzillai was a very aged man, eighty years old. He had provided the king with food while he stayed at Mahanaim, for he was a very wealthy man.
2SAM|19|33|And the king said to Barzillai, "Come over with me, and I will provide for you with me in Jerusalem."
2SAM|19|34|But Barzillai said to the king, "How many years have I still to live, that I should go up with the king to Jerusalem?
2SAM|19|35|I am this day eighty years old. Can I discern what is pleasant and what is not? Can your servant taste what he eats or what he drinks? Can I still listen to the voice of singing men and singing women? Why then should your servant be an added burden to my lord the king?
2SAM|19|36|Your servant will go a little way over the Jordan with the king. Why should the king repay me with such a reward?
2SAM|19|37|Please let your servant return, that I may die in my own city near the grave of my father and my mother. But here is your servant Chimham. Let him go over with my lord the king, and do for him whatever seems good to you."
2SAM|19|38|And the king answered, "Chimham shall go over with me, and I will do for him whatever seems good to you, and all that you desire of me I will do for you."
2SAM|19|39|Then all the people went over the Jordan, and the king went over. And the king kissed Barzillai and blessed him, and he returned to his own home.
2SAM|19|40|The king went on to Gilgal, and Chimham went on with him. All the people of Judah, and also half the people of Israel, brought the king on his way.
2SAM|19|41|Then all the men of Israel came to the king and said to the king, "Why have our brothers the men of Judah stolen you away and brought the king and his household over the Jordan, and all David's men with him?"
2SAM|19|42|All the men of Judah answered the men of Israel, "Because the king is our close relative. Why then are you angry over this matter? Have we eaten at all at the king's expense? Or has he given us any gift?"
2SAM|19|43|And the men of Israel answered the men of Judah, "We have ten shares in the king, and in David also we have more than you. Why then did you despise us? Were we not the first to speak of bringing back our king?" But the words of the men of Judah were fiercer than the words of the men of Israel.
2SAM|20|1|Now there happened to be there a worthless man, whose name was Sheba, the son of Bichri, a Benjaminite. And he blew the trumpet and said, "We have no portion in David, and we have no inheritance in the son of Jesse; every man to his tents, O Israel!"
2SAM|20|2|So all the men of Israel withdrew from David and followed Sheba the son of Bichri. But the men of Judah followed their king steadfastly from the Jordan to Jerusalem.
2SAM|20|3|And David came to his house at Jerusalem. And the king took the ten concubines whom he had left to care for the house and put them in a house under guard and provided for them, but did not go in to them. So they were shut up until the day of their death, living as if in widowhood.
2SAM|20|4|Then the king said to Amasa, "Call the men of Judah together to me within three days, and be here yourself."
2SAM|20|5|So Amasa went to summon Judah, but he delayed beyond the set time that had been appointed him.
2SAM|20|6|And David said to Abishai, "Now Sheba the son of Bichri will do us more harm than Absalom. Take your lord's servants and pursue him, lest he get himself to fortified cities and escape from us."
2SAM|20|7|And there went out after him Joab's men and the Cherethites and the Pelethites, and all the mighty men. They went out from Jerusalem to pursue Sheba the son of Bichri.
2SAM|20|8|When they were at the great stone that is in Gibeon, Amasa came to meet them. Now Joab was wearing a soldier's garment, and over it was a belt with a sword in its sheath fastened on his thigh, and as he went forward it fell out.
2SAM|20|9|And Joab said to Amasa, "Is it well with you, my brother?" And Joab took Amasa by the beard with his right hand to kiss him.
2SAM|20|10|But Amasa did not observe the sword that was in Joab's hand. So Joab struck him with it in the stomach and spilled his entrails to the ground without striking a second blow, and he died. Then Joab and Abishai his brother pursued Sheba the son of Bichri.
2SAM|20|11|And one of Joab's young men took his stand by Amasa and said, "Whoever favors Joab, and whoever is for David, let him follow Joab."
2SAM|20|12|And Amasa lay wallowing in his blood in the highway. And anyone who came by, seeing him, stopped. And when the man saw that all the people stopped, he carried Amasa out of the highway into the field and threw a garment over him.
2SAM|20|13|When he was taken out of the highway, all the people went on after Joab to pursue Sheba the son of Bichri.
2SAM|20|14|And Sheba passed through all the tribes of Israel to Abel of Beth-maacah, and all the Bichrites assembled and followed him in.
2SAM|20|15|And all the men who were with Joab came and besieged him in Abel of Beth-maacah. They cast up a mound against the city, and it stood against the rampart, and they were battering the wall to throw it down.
2SAM|20|16|Then a wise woman called from the city, "Listen! Listen! Tell Joab, 'Come here, that I may speak to you.'"
2SAM|20|17|And he came near her, and the woman said, "Are you Joab?" He answered, "I am." Then she said to him, "Listen to the words of your servant." And he answered, "I am listening."
2SAM|20|18|Then she said, "They used to say in former times, 'Let them but ask counsel at Abel,' and so they settled a matter.
2SAM|20|19|I am one of those who are peaceable and faithful in Israel. You seek to destroy a city that is a mother in Israel. Why will you swallow up the heritage of the LORD?"
2SAM|20|20|Joab answered, "Far be it from me, far be it, that I should swallow up or destroy!
2SAM|20|21|That is not true. But a man of the hill country of Ephraim, called Sheba the son of Bichri, has lifted up his hand against King David. Give up him alone, and I will withdraw from the city." And the woman said to Joab, "Behold, his head shall be thrown to you over the wall."
2SAM|20|22|Then the woman went to all the people in her wisdom. And they cut off the head of Sheba the son of Bichri and threw it out to Joab. So he blew the trumpet, and they dispersed from the city, every man to his home. And Joab returned to Jerusalem to the king.
2SAM|20|23|Now Joab was in command of all the army of Israel; and Benaiah the son of Jehoiada was in command of the Cherethites and the Pelethites;
2SAM|20|24|and Adoram was in charge of the forced labor; and Jehoshaphat the son of Ahilud was the recorder;
2SAM|20|25|and Sheva was secretary; and Zadok and Abiathar were priests;
2SAM|20|26|and Ira the Jairite was also David's priest.
2SAM|21|1|Now there was a famine in the days of David for three years, year after year. And David sought the face of the LORD. And the LORD said, "There is bloodguilt on Saul and on his house, because he put the Gibeonites to death."
2SAM|21|2|So the king called the Gibeonites and spoke to them. Now the Gibeonites were not of the people of Israel but of the remnant of the Amorites. Although the people of Israel had sworn to spare them, Saul had sought to strike them down in his zeal for the people of Israel and Judah.
2SAM|21|3|And David said to the Gibeonites, "What shall I do for you? And how shall I make atonement, that you may bless the heritage of the LORD?"
2SAM|21|4|The Gibeonites said to him, "It is not a matter of silver or gold between us and Saul or his house; neither is it for us to put any man to death in Israel." And he said, "What do you say that I shall do for you?"
2SAM|21|5|They said to the king, "The man who consumed us and planned to destroy us, so that we should have no place in all the territory of Israel,
2SAM|21|6|let seven of his sons be given to us, so that we may hang them before the LORD at Gibeah of Saul, the chosen of the LORD." And the king said, "I will give them."
2SAM|21|7|But the king spared Mephibosheth, the son of Saul's son Jonathan, because of the oath of the LORD that was between them, between David and Jonathan the son of Saul.
2SAM|21|8|The king took the two sons of Rizpah the daughter of Aiah, whom she bore to Saul, Armoni and Mephibosheth; and the five sons of Merab the daughter of Saul, whom she bore to Adriel the son of Barzillai the Meholathite;
2SAM|21|9|and he gave them into the hands of the Gibeonites, and they hanged them on the mountain before the LORD, and the seven of them perished together. They were put to death in the first days of harvest, at the beginning of barley harvest.
2SAM|21|10|Then Rizpah the daughter of Aiah took sackcloth and spread it for herself on the rock, from the beginning of harvest until rain fell upon them from the heavens. And she did not allow the birds of the air to come upon them by day, or the beasts of the field by night.
2SAM|21|11|When David was told what Rizpah the daughter of Aiah, the concubine of Saul, had done,
2SAM|21|12|David went and took the bones of Saul and the bones of his son Jonathan from the men of Jabesh-gilead, who had stolen them from the public square of Beth-shan, where the Philistines had hanged them, on the day the Philistines killed Saul on Gilboa.
2SAM|21|13|And he brought up from there the bones of Saul and the bones of his son Jonathan; and they gathered the bones of those who were hanged.
2SAM|21|14|And they buried the bones of Saul and his son Jonathan in the land of Benjamin in Zela, in the tomb of Kish his father. And they did all that the king commanded. And after that God responded to the plea for the land.
2SAM|21|15|There was war again between the Philistines and Israel, and David went down together with his servants, and they fought against the Philistines. And David grew weary.
2SAM|21|16|And Ishbi-benob, one of the descendants of the giants, whose spear weighed three hundred shekels of bronze, and who was armed with a new sword, thought to kill David.
2SAM|21|17|But Abishai the son of Zeruiah came to his aid and attacked the Philistine and killed him. Then David's men swore to him, "You shall no longer go out with us to battle, lest you quench the lamp of Israel."
2SAM|21|18|After this there was again war with the Philistines at Gob. Then Sibbecai the Hushathite struck down Saph, who was one of the descendants of the giants.
2SAM|21|19|And there was again war with the Philistines at Gob, and Elhanan the son of Jaare-oregim, the Bethlehemite, struck down Goliath the Gittite, the shaft of whose spear was like a weaver's beam.
2SAM|21|20|And there was again war at Gath, where there was a man of great stature, who had six fingers on each hand, and six toes on each foot, twenty-four in number, and he also was descended from the giants.
2SAM|21|21|And when he taunted Israel, Jonathan the son of Shimei, David's brother, struck him down.
2SAM|21|22|These four were descended from the giants in Gath, and they fell by the hand of David and by the hand of his servants.
2SAM|22|1|And David spoke to the LORD the words of this song on the day when the LORD delivered him from the hand of all his enemies, and from the hand of Saul.
2SAM|22|2|He said, "The LORD is my rock and my fortress and my deliverer,
2SAM|22|3|my God, my rock, in whom I take refuge, my shield, and the horn of my salvation, my stronghold and my refuge, my savior; you save me from violence.
2SAM|22|4|I call upon the LORD, who is worthy to be praised, and I am saved from my enemies.
2SAM|22|5|"For the waves of death encompassed me, the torrents of destruction assailed me;
2SAM|22|6|the cords of Sheol entangled me; the snares of death confronted me.
2SAM|22|7|"In my distress I called upon the LORD; to my God I called. From his temple he heard my voice, and my cry came to his ears.
2SAM|22|8|"Then the earth reeled and rocked; the foundations of the heavens trembled and quaked, because he was angry.
2SAM|22|9|Smoke went up from his nostrils, and devouring fire from his mouth; glowing coals flamed forth from him.
2SAM|22|10|He bowed the heavens and came down; thick darkness was under his feet.
2SAM|22|11|He rode on a cherub and flew; he was seen on the wings of the wind.
2SAM|22|12|He made darkness around him his canopy, thick clouds, a gathering of water.
2SAM|22|13|Out of the brightness before him coals of fire flamed forth.
2SAM|22|14|The LORD thundered from heaven, and the Most High uttered his voice.
2SAM|22|15|And he sent out arrows and scattered them; lightning, and routed them.
2SAM|22|16|Then the channels of the sea were seen; the foundations of the world were laid bare, at the rebuke of the LORD, at the blast of the breath of his nostrils.
2SAM|22|17|"He sent from on high, he took me; he drew me out of many waters.
2SAM|22|18|He rescued me from my strong enemy, from those who hated me, for they were too mighty for me.
2SAM|22|19|They confronted me in the day of my calamity, but the LORD was my support.
2SAM|22|20|He brought me out into a broad place; he rescued me, because he delighted in me.
2SAM|22|21|"The LORD dealt with me according to my righteousness; according to the cleanness of my hands he rewarded me.
2SAM|22|22|For I have kept the ways of the LORD and have not wickedly departed from my God.
2SAM|22|23|For all his rules were before me, and from his statutes I did not turn aside.
2SAM|22|24|I was blameless before him, and I kept myself from guilt.
2SAM|22|25|And the LORD has rewarded me according to my righteousness, according to my cleanness in his sight.
2SAM|22|26|"With the merciful you show yourself merciful; with the blameless man you show yourself blameless;
2SAM|22|27|with the purified you deal purely, and with the crooked you make yourself seem tortuous.
2SAM|22|28|You save a humble people, but your eyes are on the haughty to bring them down.
2SAM|22|29|For you are my lamp, O LORD, and my God lightens my darkness.
2SAM|22|30|For by you I can run against a troop, and by my God I can leap over a wall.
2SAM|22|31|This God- his way is perfect; the word of the LORD proves true; he is a shield for all those who take refuge in him.
2SAM|22|32|"For who is God, but the LORD? And who is a rock, except our God?
2SAM|22|33|This God is my strong refuge and has made my way blameless.
2SAM|22|34|He made my feet like the feet of a deer and set me secure on the heights.
2SAM|22|35|He trains my hands for war, so that my arms can bend a bow of bronze.
2SAM|22|36|You have given me the shield of your salvation, and your gentleness made me great.
2SAM|22|37|You gave a wide place for my steps under me, and my feet did not slip;
2SAM|22|38|I pursued my enemies and destroyed them, and did not turn back until they were consumed.
2SAM|22|39|I consumed them; I thrust them through, so that they did not rise; they fell under my feet.
2SAM|22|40|For you equipped me with strength for the battle; you made those who rise against me sink under me.
2SAM|22|41|You made my enemies turn their backs to me, those who hated me, and I destroyed them.
2SAM|22|42|They looked, but there was none to save; they cried to the LORD, but he did not answer them.
2SAM|22|43|I beat them fine as the dust of the earth; I crushed them and stamped them down like the mire of the streets.
2SAM|22|44|"You delivered me from strife with my people; you kept me as the head of the nations; people whom I had not known served me.
2SAM|22|45|Foreigners came cringing to me; as soon as they heard of me, they obeyed me.
2SAM|22|46|Foreigners lost heart and came trembling out of their fortresses.
2SAM|22|47|"The LORD lives, and blessed be my rock, and exalted be my God, the rock of my salvation,
2SAM|22|48|the God who gave me vengeance and brought down peoples under me,
2SAM|22|49|who brought me out from my enemies; you exalted me above those who rose against me; you delivered me from men of violence.
2SAM|22|50|"For this I will praise you, O LORD, among the nations, and sing praises to your name.
2SAM|22|51|Great salvation he brings to his king, and shows steadfast love to his anointed, to David and his offspring forever."
2SAM|23|1|Now these are the last words of David: The oracle of David, the son of Jesse, the oracle of the man who was raised on high, the anointed of the God of Jacob, the sweet psalmist of Israel:
2SAM|23|2|"The Spirit of the LORD speaks by me; his word is on my tongue.
2SAM|23|3|The God of Israel has spoken; the Rock of Israel has said to me: When one rules justly over men, ruling in the fear of God,
2SAM|23|4|he dawns on them like the morning light, like the sun shining forth on a cloudless morning, like rain that makes grass to sprout from the earth.
2SAM|23|5|For does not my house stand so with God? For he has made with me an everlasting covenant, ordered in all things and secure. For will he not cause to prosper all my help and my desire?
2SAM|23|6|But worthless men are all like thorns that are thrown away, for they cannot be taken with the hand;
2SAM|23|7|but the man who touches them arms himself with iron and the shaft of a spear, and they are utterly consumed with fire."
2SAM|23|8|These are the names of the mighty men whom David had: Josheb-basshebeth a Tahchemonite; he was chief of the three. He wielded his spear against eight hundred whom he killed at one time.
2SAM|23|9|And next to him among the three mighty men was Eleazar the son of Dodo, son of Ahohi. He was with David when they defied the Philistines who were gathered there for battle, and the men of Israel withdrew.
2SAM|23|10|He rose and struck down the Philistines until his hand was weary, and his hand clung to the sword. And the LORD brought about a great victory that day, and the men returned after him only to strip the slain.
2SAM|23|11|And next to him was Shammah, the son of Agee the Hararite. The Philistines gathered together at Lehi, where there was a plot of ground full of lentils, and the men fled from the Philistines.
2SAM|23|12|But he took his stand in the midst of the plot and defended it and struck down the Philistines, and the LORD worked a great victory.
2SAM|23|13|And three of the thirty chief men went down and came about harvest time to David at the cave of Adullam, when a band of Philistines was encamped in the Valley of Rephaim.
2SAM|23|14|David was then in the stronghold, and the garrison of the Philistines was then at Bethlehem.
2SAM|23|15|And David said longingly, "Oh, that someone would give me water to drink from the well of Bethlehem that is by the gate!"
2SAM|23|16|Then the three mighty men broke through the camp of the Philistines and drew water out of the well of Bethlehem that was by the gate and carried and brought it to David. But he would not drink of it. He poured it out to the LORD
2SAM|23|17|and said, "Far be it from me, O LORD, that I should do this. Shall I drink the blood of the men who went at the risk of their lives?" Therefore he would not drink it. These things the three mighty men did.
2SAM|23|18|Now Abishai, the brother of Joab, the son of Zeruiah, was chief of the thirty. And he wielded his spear against three hundred men and killed them and won a name beside the three.
2SAM|23|19|He was the most renowned of the thirty and became their commander, but he did not attain to the three.
2SAM|23|20|And Benaiah the son of Jehoiada was a valiant man of Kabzeel, a doer of great deeds. He struck down two ariels of Moab. He also went down and struck down a lion in a pit on a day when snow had fallen.
2SAM|23|21|And he struck down an Egyptian, a handsome man. The Egyptian had a spear in his hand, but Benaiah went down to him with a staff and snatched the spear out of the Egyptian's hand and killed him with his own spear.
2SAM|23|22|These things did Benaiah the son of Jehoiada, and won a name beside the three mighty men.
2SAM|23|23|He was renowned among the thirty, but he did not attain to the three. And David set him over his bodyguard.
2SAM|23|24|Asahel the brother of Joab was one of the thirty; Elhanan the son of Dodo of Bethlehem,
2SAM|23|25|Shammah of Harod, Elika of Harod,
2SAM|23|26|Helez the Paltite, Ira the son of Ikkesh of Tekoa,
2SAM|23|27|Abiezer of Anathoth, Mebunnai the Hushathite,
2SAM|23|28|Zalmon the Ahohite, Maharai of Netophah,
2SAM|23|29|Heleb the son of Baanah of Netophah, Ittai the son of Ribai of Gibeah of the people of Benjamin,
2SAM|23|30|Benaiah of Pirathon, Hiddai of the brooks of Gaash,
2SAM|23|31|Abi-albon the Arbathite, Azmaveth of Bahurim,
2SAM|23|32|Eliahba the Shaalbonite, the sons of Jashen, Jonathan,
2SAM|23|33|Shammah the Hararite, Ahiam the son of Sharar the Hararite,
2SAM|23|34|Eliphelet the son of Ahasbai of Maacah, Eliam the son of Ahithophel of Gilo,
2SAM|23|35|Hezro of Carmel, Paarai the Arbite,
2SAM|23|36|Igal the son of Nathan of Zobah, Bani the Gadite,
2SAM|23|37|Zelek the Ammonite, Naharai of Beeroth, the armor-bearer of Joab the son of Zeruiah,
2SAM|23|38|Ira the Ithrite, Gareb the Ithrite,
2SAM|23|39|Uriah the Hittite: thirty-seven in all.
2SAM|24|1|Again the anger of the LORD was kindled against Israel, and he incited David against them, saying, "Go, number Israel and Judah."
2SAM|24|2|So the king said to Joab, the commander of the army, who was with him, "Go through all the tribes of Israel, from Dan to Beersheba, and number the people, that I may know the number of the people."
2SAM|24|3|But Joab said to the king, "May the LORD your God add to the people a hundred times as many as they are, while the eyes of my lord the king still see it, but why does my lord the king delight in this thing?"
2SAM|24|4|But the king's word prevailed against Joab and the commanders of the army. So Joab and the commanders of the army went out from the presence of the king to number the people of Israel.
2SAM|24|5|They crossed the Jordan and began from Aroer, and from the city that is in the middle of the valley, toward Gad and on to Jazer.
2SAM|24|6|Then they came to Gilead, and to Kadesh in the land of the Hittites; and they came to Dan, and from Dan they went around to Sidon,
2SAM|24|7|and came to the fortress of Tyre and to all the cities of the Hivites and Canaanites; and they went out to the Negeb of Judah at Beersheba.
2SAM|24|8|So when they had gone through all the land, they came to Jerusalem at the end of nine months and twenty days.
2SAM|24|9|And Joab gave the sum of the numbering of the people to the king: in Israel there were 800,000 valiant men who drew the sword, and the men of Judah were 500,000.
2SAM|24|10|But David's heart struck him after he had numbered the people. And David said to the LORD, "I have sinned greatly in what I have done. But now, O LORD, please take away the iniquity of your servant, for I have done very foolishly."
2SAM|24|11|And when David arose in the morning, the word of the LORD came to the prophet Gad, David's seer, saying,
2SAM|24|12|"Go and say to David, 'Thus says the LORD, Three things I offer you. Choose one of them, that I may do it to you.'"
2SAM|24|13|So Gad came to David and told him, and said to him, "Shall three years of famine come to you in your land? Or will you flee three months before your foes while they pursue you? Or shall there be three days' pestilence in your land? Now consider, and decide what answer I shall return to him who sent me."
2SAM|24|14|Then David said to Gad, "I am in great distress. Let us fall into the hand of the LORD, for his mercy is great; but let me not fall into the hand of man."
2SAM|24|15|So the LORD sent a pestilence on Israel from the morning until the appointed time. And there died of the people from Dan to Beersheba 70,000 men.
2SAM|24|16|And when the angel stretched out his hand toward Jerusalem to destroy it, the LORD relented from the calamity and said to the angel who was working destruction among the people, "It is enough; now stay your hand." And the angel of the LORD was by the threshing floor of Araunah the Jebusite.
2SAM|24|17|Then David spoke to the LORD when he saw the angel who was striking the people, and said, "Behold, I have sinned, and I have done wickedly. But these sheep, what have they done? Please let your hand be against me and against my father's house."
2SAM|24|18|And Gad came that day to David and said to him, "Go up, raise an altar to the LORD on the threshing floor of Araunah the Jebusite."
2SAM|24|19|So David went up at Gad's word, as the LORD commanded.
2SAM|24|20|And when Araunah looked down, he saw the king and his servants coming on toward him. And Araunah went out and paid homage to the king with his face to the ground.
2SAM|24|21|And Araunah said, "Why has my lord the king come to his servant?" David said, "To buy the threshing floor from you, in order to build an altar to the LORD, that the plague may be averted from the people."
2SAM|24|22|Then Araunah said to David, "Let my lord the king take and offer up what seems good to him. Here are the oxen for the burnt offering and the threshing sledges and the yokes of the oxen for the wood.
2SAM|24|23|All this, O king, Araunah gives to the king." And Araunah said to the king, "The LORD your God accept you."
2SAM|24|24|But the king said to Araunah, "No, but I will buy it from you for a price. I will not offer burnt offerings to the LORD my God that cost me nothing." So David bought the threshing floor and the oxen for fifty shekels of silver.
2SAM|24|25|And David built there an altar to the LORD and offered burnt offerings and peace offerings. So the LORD responded to the plea for the land, and the plague was averted from Israel.
