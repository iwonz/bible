MARK|1|1|Initium evangelii Iesu Christi Filii Dei.
MARK|1|2|Sicut scriptum est in Isaia propheta: Ecce mitto angelum meum ante faciem tuam,qui praeparabit viam tuam;
MARK|1|3|vox clamantis in deserto:Parate viam Domini, rectas facite semitas eius" ",
MARK|1|4|fuit Ioannes Baptista in deserto praedicans baptismum paenitentiae in remissionem peccatorum.
MARK|1|5|Et egrediebatur ad illum omnis Iudaeae regio et Hierosolymitae universi et baptizabantur ab illo in Iordane flumine confitentes peccata sua.
MARK|1|6|Et erat Ioannes vestitus pilis cameli, et zona pellicea circa lumbos eius, et locustas et mel silvestre edebat.
MARK|1|7|Et praedicabat dicens: " Venit fortior me post me, cuius non sum dignus procumbens solvere corrigiam calceamentorum eius.
MARK|1|8|Ego baptizavi vos aqua; ille vero baptizabit vos in Spiritu Sancto ".
MARK|1|9|Et factum est in diebus illis, venit Iesus a Nazareth Galilaeae et baptizatus est in Iordane ab Ioanne.
MARK|1|10|Et statim ascendens de aqua vidit apertos caelos et Spiritum tamquam columbam descendentem in ipsum;
MARK|1|11|et vox facta est de caelis: " Tu es Filius meus dilectus; in te complacui ".
MARK|1|12|Et statim Spiritus expellit eum in desertum.
MARK|1|13|Et erat in deserto quadraginta diebus et tentabatur a Satana; eratque cum bestiis, et angeli ministrabant illi.
MARK|1|14|Postquam autem traditus est Ioannes, venit Iesus in Galilaeam praedicans evangelium Dei
MARK|1|15|et dicens: " Impletum est tempus, et appropinquavit regnum Dei; paenitemini et credite evangelio ".
MARK|1|16|Et praeteriens secus mare Galilaeae vidit Simonem et Andream fratrem Simonis mittentes in mare; erant enim piscatores.
MARK|1|17|Et dixit eis Iesus: " Venite post me, et faciam vos fieri piscatores hominum ".
MARK|1|18|Et protinus, relictis retibus, secuti sunt eum.
MARK|1|19|Et progressus pusillum vidit Iacobum Zebedaei et Ioannem fratrem eius, et ipsos in navi componentes retia,
MARK|1|20|et statim vocavit illos. Et, relicto patre suo Zebedaeo in navi cum mercennariis, abierunt post eum.
MARK|1|21|Et ingrediuntur Capharnaum. Et statim sabbatis ingressus synagogam docebat.
MARK|1|22|Et stupebant super doctrina eius: erat enim docens eos quasi potestatem habens et non sicut scribae.
MARK|1|23|Et statim erat in synagoga eorum homo in spiritu immundo; et exclamavit
MARK|1|24|dicens: " Quid nobis et tibi, Iesu Nazarene? Venisti perdere nos? Scio qui sis: Sanctus Dei ".
MARK|1|25|Et comminatus est ei Iesus dicens: " Obmutesce et exi de homine! ".
MARK|1|26|Et discerpens eum spiritus immundus et exclamans voce magna exivit ab eo.
MARK|1|27|Et mirati sunt omnes, ita ut conquirerent inter se dicentes: " Quidnam est hoc? Doctrina nova cum potestate; et spiritibus immundis imperat, et oboediunt ei ".
MARK|1|28|Et processit rumor eius statim ubique in omnem regionem Galilaeae.
MARK|1|29|Et protinus egredientes de synagoga venerunt in domum Simonis et Andreae cum Iacobo et Ioanne.
MARK|1|30|Socrus autem Simonis decumbebat febricitans; et statim dicunt ei de illa.
MARK|1|31|Et accedens elevavit eam apprehensa manu; et dimisit eam febris, et ministrabat eis.
MARK|1|32|Vespere autem facto, cum occidisset sol, afferebant ad eum omnes male habentes et daemonia habentes;
MARK|1|33|et erat omnis civitas congregata ad ianuam.
MARK|1|34|Et curavit multos, qui vexabantur variis languoribus, et daemonia multa eiecit et non sinebat loqui daemonia, quoniam sciebant eum.
MARK|1|35|Et diluculo valde mane surgens egressus est et abiit in desertum locum ibique orabat.
MARK|1|36|Et persecutus est eum Simon et qui cum illo erant;
MARK|1|37|et cum invenissent eum, dixerunt ei: " Omnes quaerunt te! ".
MARK|1|38|Et ait illis: " Eamus alibi in proximos vicos, ut et ibi praedicem: ad hoc enim veni ".
MARK|1|39|Et venit praedicans in synagogis eorum per omnem Galilaeam et daemonia eiciens.
MARK|1|40|Et venit ad eum leprosus deprecans eum et genu flectens et dicens ei: " Si vis, potes me mundare ".
MARK|1|41|Et misertus extendens manum suam tetigit eum et ait illi: " Volo, mundare! ";
MARK|1|42|et statim discessit ab eo lepra, et mundatus est.
MARK|1|43|Et infremuit in eum statimque eiecit illum
MARK|1|44|et dicit ei: "Vide, nemini quidquam dixeris; sed vade, ostende te sacerdoti et offer pro emundatione tua, quae praecepit Moyses, in testimonium illis ".
MARK|1|45|At ille egressus coepit praedicare multum et diffamare sermonem, ita ut iam non posset manifesto in civitatem introire, sed foris in desertis locis erat; et conveniebant ad eum undique.
MARK|2|1|Et iterum intravit Capharnaum post dies, et auditum est quod in domo esset.
MARK|2|2|Et convenerunt multi, ita ut non amplius caperentur neque ad ianuam, et loquebatur eis verbum.
MARK|2|3|Et veniunt ferentes ad eum paralyticum, qui a quattuor portabatur.
MARK|2|4|Et cum non possent offerre eum illi prae turba, nudaverunt tectum, ubi erat, et perfodientes summittunt grabatum, in quo paralyticus iacebat.
MARK|2|5|Cum vidisset autem Iesus fidem illorum, ait paralytico: " Fili, dimittuntur peccata tua ".
MARK|2|6|Erant autem illic quidam de scribis sedentes et cogitantes in cordibus suis:
MARK|2|7|" Quid hic sic loquitur? Blasphemat! Quis potest dimittere peccata nisi solus Deus? ".
MARK|2|8|Quo statim cognito Iesus spiritu suo quia sic cogitarent intra se, dicit illis: " Quid ista cogitatis in cordibus vestris?
MARK|2|9|Quid est facilius, dicere paralytico: "Dimittuntur peccata tua", an dicere: "Surge et tolle grabatum tuum et ambula"?
MARK|2|10|Ut autem sciatis quia potestatem habet Filius hominis interra dimittendi peccata - ait paralytico -:
MARK|2|11|Tibi dico: Surge, tolle grabatum tuum et vade in domum tuam ".
MARK|2|12|Et surrexit et protinus sublato grabato abiit coram omnibus, ita ut admirarentur omnes et glorificarent Deum dicentes: " Numquam sic vidimus!.
MARK|2|13|Et egressus est rursus ad mare; omnisque turba veniebat ad eum, et docebat eos.
MARK|2|14|Et cum praeteriret, vidit Levin Alphaei sedentem ad teloneum et ait illi: " Sequere me ". Et surgens secutus est eum.
MARK|2|15|Et factum est, cum accumberet in domo illius, et multi publicani et peccatores simul discumbebant cum Iesu et discipulis eius; erant enim multi et sequebantur eum.
MARK|2|16|Et scribae pharisaeorum, videntes quia manducaret cum peccatoribus et publicanis, dicebant discipulis eius: " Quare cum publicanis et peccatoribus manducat? ".
MARK|2|17|Et Iesus hoc audito ait illis: " Non necesse habent sani medicum, sed qui male habent; non veni vocare iustos sed peccatores ".
MARK|2|18|Et erant discipuli Ioannis et pharisaei ieiunantes. Et veniunt et dicunt illi: " Cur discipuli Ioannis et discipuli pharisaeorum ieiunant, tui autem discipuli non ieiunant? ".
MARK|2|19|Et ait illis Iesus: " Numquid possunt convivae nuptiarum, quamdiu sponsus cum illis est, ieiunare? Quanto tempore habent secum sponsum, non possunt ieiunare;
MARK|2|20|venient autem dies, cum auferetur ab eis sponsus, et tunc ieiunabunt in illa die.
MARK|2|21|Nemo assumentum panni rudis assuit vestimento veteri; alioquin supplementum aufert aliquid ab eo, novum a veteri, et peior scissura fit.
MARK|2|22|Et nemo mittit vinum novellum in utres veteres, alioquin dirumpet vinum utres et vinum perit et utres; sed vinum novum in utres novos ".
MARK|2|23|Et factum est, cum ipse sabbatis ambularet per sata, discipuli eius coeperunt praegredi vellentes spicas.
MARK|2|24|Pharisaei autem dicebant ei: " Ecce, quid faciunt sabbatis, quod non licet? ".
MARK|2|25|Et ait illis: " Numquam legistis quid fecerit David, quando necessitatem habuit et esuriit ipse et qui cum eo erant?
MARK|2|26|Quomodo introivit in domum Dei sub Abiathar principe sacerdotum et panes propositionis manducavit, quos non licet manducare nisi sacerdotibus, et dedit etiam eis, qui cum eo erant? ".
MARK|2|27|Et dicebat eis: " Sabbatum propter hominem factum est, et non homo propter sabbatum;
MARK|2|28|itaque dominus est Filius hominis etiam sabbati ".
MARK|3|1|Et introivit iterum in synago gam. Et erat ibi homo habens manum aridam;
MARK|3|2|et observabant eum, si sabbatis curaret illum, ut accusarent eum.
MARK|3|3|Et ait homini habenti manum aridam: " Surge in medium ".
MARK|3|4|Et dicit eis: " Licet sabbatis bene facere an male? Animam salvam facere an perdere? ". At illi tacebant.
MARK|3|5|Et circumspiciens eos cum ira, contristatus super caecitate cordis eorum, dicit homini: " Extende manum ". Et extendit, et restituta est manus eius.
MARK|3|6|Et exeuntes pharisaei statim cum herodianis consilium faciebant adversus eum quomodo eum perderent.
MARK|3|7|Et Iesus cum discipulis suis secessit ad mare. Et multa turba a Galilaea secuta est et a Iudaea
MARK|3|8|et ab Hierosolymis et ab Idumaea; et, qui trans Iordanem et circa Tyrum et Sidonem, multitudo magna, audientes, quae faciebat, venerunt ad eum.
MARK|3|9|Et dixit discipulis suis, ut navicula sibi praesto esset propter turbam, ne comprimerent eum.
MARK|3|10|Multos enim sanavit, ita ut irruerent in eum, ut illum tangerent, quotquot habebant plagas.
MARK|3|11|Et spiritus immundi, cum illum videbant, procidebant ei et clamabant dicentes: " Tu es Filius Dei! ".
MARK|3|12|Et vehementer comminabatur eis, ne manifestarent illum.
MARK|3|13|Et ascendit in montem et vocat ad se, quos voluit ipse, et venerunt ad eum.
MARK|3|14|Et fecit Duodecim, ut essent cum illo, et ut mitteret eos praedicare
MARK|3|15|habentes potestatem eiciendi daemonia:
MARK|3|16|et imposuit Simoni nomen Petrum;
MARK|3|17|et Iacobum Zebedaei et Ioannem fratrem Iacobi, et imposuit eis nomina Boanerges, quod est Filii tonitrui;
MARK|3|18|et Andream et Philippum et Bartholomaeum et Matthaeum et Thomam et Iacobum Alphaei et Thaddaeum et Simonem Chananaeum
MARK|3|19|et Iudam Iscarioth, qui et tradidit illum.
MARK|3|20|Et venit ad domum; et convenit iterum turba, ita ut non possent neque panem manducare.
MARK|3|21|Et cum audissent sui, exierunt tenere eum; dicebant enim: " In furorem versus est ".
MARK|3|22|Et scribae, qui ab Hierosolymis descenderant, dicebant: " Beelzebul habet " et: " In principe daemonum eicit daemonia ".
MARK|3|23|Et convocatis eis, in parabolis dicebat illis: " Quomodo potest Satanas Satanam eicere?
MARK|3|24|Et si regnum in se dividatur, non potest stare regnum illud;
MARK|3|25|et si domus in semetipsam dispertiatur, non poterit domus illa stare.
MARK|3|26|Et si Satanas consurrexit in semetipsum et dispertitus est, non potest stare, sed finem habet.
MARK|3|27|Nemo autem potest in domum fortis ingressus vasa eius diripere, nisi prius fortem alliget; et tunc domum eius diripiet.
MARK|3|28|Amen dico vobis: Omnia dimittentur filiis hominum peccata et blasphemiae, quibus blasphemaverint;
MARK|3|29|qui autem blasphemaverit in Spiritum Sanctum, non habet remissionem in aeternum, sed reus est aeterni delicti ".
MARK|3|30|Quoniam dicebant: " Spiritum immundum habet ".
MARK|3|31|Et venit mater eius et fratres eius, et foris stantes miserunt ad eum vocantes eum.
MARK|3|32|Et sedebat circa eum turba, et dicunt ei: " Ecce mater tua et fratres tui et sorores tuae foris quaerunt te ".
MARK|3|33|Et respondens eis ait: " Quae est mater mea et fratres mei? ".
MARK|3|34|Et circumspiciens eos, qui in circuitu eius sedebant, ait: " Ecce mater mea et fratres mei.
MARK|3|35|Qui enim fecerit voluntatem Dei, hic frater meus et soror mea et mater est ".
MARK|4|1|Et iterum coepit docere ad ma re. Et congregatur ad eum tur ba plurima, ita ut in navem ascendens sederet in mari, et omnis turba circa mare super terram erant.
MARK|4|2|Et docebat eos in parabolis multa et dicebat illis in doctrina sua:
MARK|4|3|" Audite. Ecce exiit seminans ad seminandum.
MARK|4|4|Et factum est, dum seminat, aliud cecidit circa viam, et venerunt volucres et comederunt illud.
MARK|4|5|Aliud cecidit super petrosa, ubi non habebat terram multam, et statim exortum est, quoniam non habebat altitudinem terrae;
MARK|4|6|et quando exortus est sol, exaestuavit et, eo quod non haberet radicem, exaruit.
MARK|4|7|Et aliud cecidit in spinas, et ascenderunt spinae et suffocaverunt illud, et fructum non dedit.
MARK|4|8|Et alia ceciderunt in terram bonam et dabant fructum: ascendebant et crescebant et afferebant unum triginta et unum sexaginta et unum centum ".
MARK|4|9|Et dicebat: " Qui habet aures audiendi, audiat ".
MARK|4|10|Et cum esset singularis, interrogaverunt eum hi, qui circa eum erant cum Duodecim, parabolas.
MARK|4|11|Et dicebat eis: " Vobis datum est mysterium regni Dei; illis autem, qui foris sunt, in parabolis omnia fiunt,
MARK|4|12|ut videntes videant et non videant,et audientes audiant et non intellegant,ne quando convertantur,et dimittatur eis ".
MARK|4|13|Et ait illis: " Nescitis parabolam hanc, et quomodo omnes parabolas cognoscetis?
MARK|4|14|Qui seminat, verbum seminat.
MARK|4|15|Hi autem sunt, qui circa viam, ubi seminatur verbum: et cum audierint, confestim venit Satanas et aufert verbum, quod seminatum est in eos.
MARK|4|16|Et hi sunt, qui super petrosa seminantur: qui cum audierint verbum, statim cum gaudio accipiunt illud
MARK|4|17|et non habent radicem in se, sed temporales sunt; deinde orta tribulatione vel persecutione propter verbum, confestim scandalizantur.
MARK|4|18|Et alii sunt, qui in spinis seminantur: hi sunt, qui verbum audierunt,
MARK|4|19|et aerumnae saeculi et deceptio divitiarum et circa reliqua concupiscentiae introeuntes suffocant verbum, et sine fructu efficitur.
MARK|4|20|Et hi sunt, qui super terram bonam seminati sunt: qui audiunt verbum et suscipiunt et fructificant unum triginta et unum sexaginta et unum centum.
MARK|4|21|Et dicebat illis: " Numquid venit lucerna, ut sub modio ponatur aut sub lecto? Nonne ut super candelabrum ponatur?
MARK|4|22|Non enim est aliquid absconditum, nisi ut manifestetur, nec factum est occultum, nisi ut in palam veniat.
MARK|4|23|Si quis habet aures audiendi, audiat ".
MARK|4|24|Et dicebat illis: " Videte quid audiatis. In qua mensura mensi fueritis, remetietur vobis et adicietur vobis.
MARK|4|25|Qui enim habet, dabitur illi; et, qui non habet, etiam quod habet, auferetur ab illo ".
MARK|4|26|Et dicebat: " Sic est regnum Dei, quemadmodum si homo iaciat sementem in terram
MARK|4|27|et dormiat et exsurgat nocte ac die, et semen germinet et increscat, dum nescit ille.
MARK|4|28|Ultro terra fructificat primum herbam, deinde spicam, deinde plenum frumentum in spica.
MARK|4|29|Et cum se produxerit fructus, statim mittit falcem, quoniam adest messis ".
MARK|4|30|Et dicebat: " Quomodo assimilabimus regnum Dei aut in qua parabola ponemus illud?
MARK|4|31|Sicut granum sinapis, quod cum seminatum fuerit in terra, minus est omnibus seminibus, quae sunt in terra;
MARK|4|32|et cum seminatum fuerit, ascendit et fit maius omnibus holeribus et facit ramos magnos, ita ut possint sub umbra eius aves caeli habitare ".
MARK|4|33|Et talibus multis parabolis loquebatur eis verbum, prout poterant audire;
MARK|4|34|sine parabola autem non loquebatur eis. Seorsum autem discipulis suis disserebat omnia.
MARK|4|35|Et ait illis illa die, cum sero esset factum: " Transeamus contra ".
MARK|4|36|Et dimittentes turbam, assumunt eum, ut erat in navi; et aliae naves erant cum illo.
MARK|4|37|Et exoritur procella magna venti, et fluctus se mittebant in navem, ita ut iam impleretur navis.
MARK|4|38|Et erat ipse in puppi supra cervical dormiens; et excitant eum et dicunt ei: " Magister, non ad te pertinet quia perimus? ".
MARK|4|39|Et exsurgens comminatus est vento et dixit mari: " Tace, obmutesce! ". Et cessavit ventus, et facta est tranquillitas magna.
MARK|4|40|Et ait illis: " Quid timidi estis? Necdum habetis fidem? ".
MARK|4|41|Et timuerunt magno timore et dicebant ad alterutrum: " Quis putas est iste, quia et ventus et mare oboediunt ei? ".
MARK|5|1|Et venerunt trans fretum maris in regionem Gerasenorum.
MARK|5|2|Et exeunte eo de navi, statim occurrit ei de monumentis homo in spiritu immundo,
MARK|5|3|qui domicilium habebat in monumentis; et neque catenis iam quisquam eum poterat ligare,
MARK|5|4|quoniam saepe compedibus et catenis vinctus dirupisset catenas et compedes comminuisset, et nemo poterat eum domare;
MARK|5|5|et semper nocte ac die in monumentis et in montibus erat clamans et concidens se lapidibus.
MARK|5|6|Et videns Iesum a longe cucurrit et adoravit eum
MARK|5|7|et clamans voce magna dicit: " Quid mihi et tibi, Iesu, fili Dei Altissimi? Adiuro te per Deum, ne me torqueas ".
MARK|5|8|Dicebat enim illi: " Exi, spiritus immunde, ab homine ".
MARK|5|9|Et interrogabat eum: " Quod tibi nomen est? ". Et dicit ei: " Legio nomen mihi est, quia multi sumus ".
MARK|5|10|Et deprecabatur eum multum, ne se expelleret extra regionem.
MARK|5|11|Erat autem ibi circa montem grex porcorum magnus pascens;
MARK|5|12|et deprecati sunt eum dicentes: " Mitte nos in porcos, ut in eos introeamus ".
MARK|5|13|Et concessit eis. Et exeuntes spiritus immundi introierunt in porcos. Et magno impetu grex ruit per praecipitium in mare, ad duo milia, et suffocabantur in mari.
MARK|5|14|Qui autem pascebant eos, fugerunt et nuntiaverunt in civitatem et in agros; et egressi sunt videre quid esset facti.
MARK|5|15|Et veniunt ad Iesum; et vident illum, qui a daemonio vexabatur, sedentem, vestitum et sanae mentis, eum qui legionem habuerat, et timuerunt.
MARK|5|16|Et qui viderant, narraverunt illis qualiter factum esset ei, qui daemonium habuerat, et de porcis.
MARK|5|17|Et rogare eum coeperunt, ut discederet a finibus eorum.
MARK|5|18|Cumque ascenderet navem, qui daemonio vexatus fuerat, deprecabatur eum, ut esset cum illo.
MARK|5|19|Et non admisit eum, sed ait illi: " Vade in domum tuam ad tuos et annuntia illis quanta tibi Dominus fecerit et misertus sit tui ".
MARK|5|20|Et abiit et coepit praedicare in Decapoli quanta sibi fecisset Iesus, et omnes mirabantur.
MARK|5|21|Et cum transcendisset Iesus in navi rursus trans fretum, convenit turba multa ad illum, et erat circa mare.
MARK|5|22|Et venit quidam de archisynagogis nomine Iairus et videns eum procidit ad pedes eius
MARK|5|23|et deprecatur eum multum dicens: " Filiola mea in extremis est; veni, impone manus super eam, ut salva sit et vivat ".
MARK|5|24|Et abiit cum illo. Et sequebatur eum turba multa et comprimebant illum.
MARK|5|25|Et mulier, quae erat in profluvio sanguinis annis duodecim
MARK|5|26|et fuerat multa perpessa a compluribus medicis et erogaverat omnia sua nec quidquam profecerat, sed magis deterius habebat,
MARK|5|27|cum audisset de Iesu, venit in turba retro et tetigit vestimentum eius;
MARK|5|28|dicebat enim: " Si vel vestimenta eius tetigero, salva ero ".
MARK|5|29|Et confestim siccatus est fons sanguinis eius, et sensit corpore quod sanata esset a plaga.
MARK|5|30|Et statim Iesus cognoscens in semetipso virtutem, quae exierat de eo, conversus ad turbam aiebat: " Quis tetigit vestimenta mea? ".
MARK|5|31|Et dicebant ei discipuli sui: " Vides turbam comprimentem te et dicis: Quis me tetigit?" ".
MARK|5|32|Et circumspiciebat videre eam, quae hoc fecerat.
MARK|5|33|Mulier autem timens et tremens, sciens quod factum esset in se, venit et procidit ante eum et dixit ei omnem veritatem.
MARK|5|34|Ille autem dixit ei: " Filia, fides tua te salvam fecit. Vade in pace et esto sana a plaga tua ".
MARK|5|35|Adhuc eo loquente, veniunt ab archisynagogo dicentes: " Filia tua mortua est; quid ultra vexas magistrum? ".
MARK|5|36|Iesus autem, verbo, quod dicebatur, audito, ait archisynagogo: " Noli timere; tantummodo crede! ".
MARK|5|37|Et non admisit quemquam sequi se nisi Petrum et Iacobum et Ioannem fratrem Iacobi.
MARK|5|38|Et veniunt ad domum archisynagogi; et videt tumultum et flentes et eiulantes multum,
MARK|5|39|et ingressus ait eis: " Quid turbamini et ploratis? Puella non est mortua, sed dormit ".
MARK|5|40|Et irridebant eum. Ipse vero, eiectis omnibus, assumit patrem puellae et matrem et, qui secum erant, et ingreditur, ubi erat puella;
MARK|5|41|et tenens manum puellae ait illi: " Talitha, qum! " - quod est interpretatum: " Puella, tibi dico: Surge! " -.
MARK|5|42|Et confestim surrexit puella et ambulabat; erat enim annorum duodecim. Et obstupuerunt continuo stupore magno.
MARK|5|43|Et praecepit illis vehementer, ut nemo id sciret, et dixit dari illi manducare.
MARK|6|1|Et egressus est inde et venit in patriam suam, et sequuntur il lum discipuli sui.
MARK|6|2|Et facto sabbato, coepit in synagoga docere; et multi audientes admirabantur dicentes: " Unde huic haec, et quae est sapientia, quae data est illi, et virtutes tales, quae per manus eius efficiuntur?
MARK|6|3|Nonne iste est faber, filius Mariae et frater Iacobi et Iosetis et Iudae et Simonis? Et nonne sorores eius hic nobiscum sunt? ". Et scandalizabantur in illo.
MARK|6|4|Et dicebat eis Iesus: " Non est propheta sine honore nisi in patria sua et in cognatione sua et in domo sua ".
MARK|6|5|Et non poterat ibi virtutem ullam facere, nisi paucos infirmos impositis manibus curavit;
MARK|6|6|et mirabatur propter incredulitatem eorum.Et circumibat castella in circuitu docens.
MARK|6|7|Et convocat Duodecim et coepit eos mittere binos et dabat illis potestatem in spiritus immundos;
MARK|6|8|et praecepit eis, ne quid tollerent in via nisi virgam tantum: non panem, non peram neque in zona aes,
MARK|6|9|sed ut calcearentur sandaliis et ne induerentur duabus tunicis.
MARK|6|10|Et dicebat eis: " Quocumque introieritis in domum, illic manete, donec exeatis inde.
MARK|6|11|Et quicumque locus non receperit vos nec audierint vos, exeuntes inde excutite pulverem de pedibus vestris in testimonium illis ".
MARK|6|12|Et exeuntes praedicaverunt, ut paenitentiam agerent;
MARK|6|13|et daemonia multa eiciebant et ungebant oleo multos aegrotos et sanabant.
MARK|6|14|Et audivit Herodes rex; manifestum enim factum est nomen eius. Et dicebant: " Ioannes Baptista resurrexit a mortuis, et propterea inoperantur virtutes in illo ".
MARK|6|15|Alii autem dicebant: " Elias est ". Alii vero dicebant: " Propheta est, quasi unus ex prophetis ".
MARK|6|16|Quo audito, Herodes aiebat: " Quem ego decollavi Ioannem, hic resurrexit! ".
MARK|6|17|Ipse enim Herodes misit ac tenuit Ioannem et vinxit eum in carcere propter Herodiadem uxorem Philippi fratris sui, quia duxerat eam.
MARK|6|18|Dicebat enim Ioannes Herodi: " Non licet tibi habere uxorem fratris tui.
MARK|6|19|Herodias autem insidiabatur illi et volebat occidere eum nec poterat:
MARK|6|20|Herodes enim metuebat Ioannem, sciens eum virum iustum et sanctum, et custodiebat eum, et, audito eo, multum haesitabat et libenter eum audiebat.
MARK|6|21|Et cum dies opportunus accidisset, quo Herodes natali suo cenam fecit principibus suis et tribunis et primis Galilaeae,
MARK|6|22|cumque introisset filia ipsius Herodiadis et saltasset, placuit Herodi simulque recumbentibus. Rex ait puellae: " Pete a me, quod vis, et dabo tibi ".
MARK|6|23|Et iuravit illi multum: " Quidquid petieris a me, dabo tibi, usque ad dimidium regni mei ".
MARK|6|24|Quae cum exisset, dixit matri suae: " Quid petam? ". At illa dixit: " Caput Ioannis Baptistae ".
MARK|6|25|Cumque introisset statim cum festinatione ad regem, petivit dicens: " Volo ut protinus des mihi in disco caput Ioannis Baptistae ".
MARK|6|26|Et contristatus rex, propter iusiurandum et propter recumbentes noluit eam decipere;
MARK|6|27|et statim misso spiculatore rex praecepit afferri caput eius. Et abiens decollavit eum in carcere
MARK|6|28|et attulit caput eius in disco; et dedit illud puellae, et puella dedit illud matri suae.
MARK|6|29|Quo audito, discipuli eius venerunt et tulerunt corpus eius et posuerunt illud in monumento.
MARK|6|30|Et convenientes apostoli ad Iesum renuntiaverunt illi omnia, quae egerant et docuerant.
MARK|6|31|Et ait illis: " Venite vos ipsi seorsum in desertum locum et requiescite pusillum ". Erant enim, qui veniebant et redibant, multi, et nec manducandi spatium habebant.
MARK|6|32|Et abierunt in navi in desertum locum seorsum.
MARK|6|33|Et viderunt eos abeuntes et cognoverunt multi; et pedestre de omnibus civitatibus concurrerunt illuc et praevenerunt eos.
MARK|6|34|Et exiens vidit multam turbam et misertus est super eos, quia erant sicut oves non habentes pastorem, et coepit docere illos multa.
MARK|6|35|Et cum iam hora multa facta esset, accesserunt discipuli eius dicentes: Desertus est locus hic, et hora iam est multa;
MARK|6|36|dimitte illos, ut euntes in villas et vicos in circuitu emant sibi, quod manducent ".
MARK|6|37|Respondens autem ait illis: " Date illis vos manducare ". Et dicunt ei: Euntes emamus denariis ducentis panes et dabimus eis manducare? ".
MARK|6|38|Et dicit eis: " Quot panes habetis? Ite, videte ". Et cum cognovissent, dicunt: " Quinque et duos pisces ".
MARK|6|39|Et praecepit illis, ut accumbere facerent omnes secundum contubernia super viride fenum.
MARK|6|40|Et discubuerunt secundum areas per centenos et per quinquagenos.
MARK|6|41|Et acceptis quinque panibus et duobus piscibus, intuens in caelum benedixit et fregit panes et dabat discipulis suis, ut ponerent ante eos; et duos pisces divisit omnibus.
MARK|6|42|Et manducaverunt omnes et saturati sunt;
MARK|6|43|et sustulerunt fragmenta duodecim cophinos plenos, et de piscibus.
MARK|6|44|Et erant, qui manducaverunt panes, quinque milia virorum.
MARK|6|45|Et statim coegit discipulos suos ascendere navem, ut praecederent trans fretum ad Bethsaidam, dum ipse dimitteret populum.
MARK|6|46|Et cum dimisisset eos, abiit in montem orare.
MARK|6|47|Et cum sero factum esset, erat navis in medio mari, et ipse solus in terra.
MARK|6|48|Et videns eos laborantes in remigando, erat enim ventus contrarius eis, circa quartam vigiliam noctis venit ad eos ambulans super mare et volebat praeterire eos.
MARK|6|49|At illi, ut viderunt eum ambulantem super mare, putaverunt phantasma esse et exclamaverunt;
MARK|6|50|omnes enim eum viderunt et conturbati sunt. Statim autem locutus est cum eis et dicit illis: " Confidite, ego sum; nolite timere! ".
MARK|6|51|Et ascendit ad illos in navem, et cessavit ventus. Et valde nimis intra se stupebant;
MARK|6|52|non enim intellexerant de panibus, sed erat cor illorum obcaecatum.
MARK|6|53|Et cum transfretassent in terram, pervenerunt Gennesaret et applicuerunt.
MARK|6|54|Cumque egressi essent de navi, continuo cognoverunt eum
MARK|6|55|et percurrentes universam regionem illam coeperunt in grabatis eos, qui se male habebant, circumferre, ubi audiebant eum esse.
MARK|6|56|Et quocumque introibat in vicos aut in civitates vel in villas, in plateis ponebant infirmos; et deprecabantur eum, ut vel fimbriam vestimenti eius tangerent; et, quotquot tangebant eum, salvi fiebant.
MARK|7|1|Et conveniunt ad eum pharisaei et quidam de scribis venientes ab Hierosolymis;
MARK|7|2|et cum vidissent quosdam ex discipulis eius communibus manibus, id est non lotis, manducare panes
MARK|7|3|- pharisaei enim et omnes Iudaei, nisi pugillo lavent manus, non manducant, tenentes traditionem seniorum;
MARK|7|4|et a foro nisi baptizentur, non comedunt; et alia multa sunt, quae acceperunt servanda: baptismata calicum et urceorum et aeramentorum et lectorum -
MARK|7|5|et interrogant eum pharisaei et scribae: " Quare discipuli tui non ambulant iuxta traditionem seniorum, sed communibus manibus manducant panem? ".
MARK|7|6|At ille dixit eis: " Bene prophetavit Isaias de vobis hypocritis, sicut scriptum est:Populus hic labiis me honorat,cor autem eorum longe est a me;
MARK|7|7|in vanum autem me coluntdocentes doctrinas praecepta hominum".
MARK|7|8|Relinquentes mandatum Dei tenetis traditionem hominum ".
MARK|7|9|Et dicebat illis: " Bene irritum facitis praeceptum Dei, ut traditionem vestram servetis.
MARK|7|10|Moyses enim dixit: "Honora patrem tuum et matrem tuam" et: "Qui maledixerit patri aut matri, morte moriatur";
MARK|7|11|vos autem dicitis: "Si dixerit homo patri aut matri: Corban, quod est donum, quodcumque ex me tibi profuerit",
MARK|7|12|ultra non permittitis ei facere quidquam patri aut matri
MARK|7|13|rescindentes verbum Dei per traditionem vestram, quam tradidistis; et similia huiusmodi multa facitis ".
MARK|7|14|Et advocata iterum turba, dicebat illis: " Audite me, omnes, et intellegite:
MARK|7|15|Nihil est extra hominem introiens in eum, quod possiteum coinquinare; sed quae de homine procedunt, illa sunt, quae coinquinant hominem! ".
MARK|7|16|()
MARK|7|17|Et cum introisset in domum a turba, interrogabant eum discipuli eius parabolam.
MARK|7|18|Et ait illis: " Sic et vos imprudentes estis? Non intellegitis quia omne extrinsecus introiens in hominem non potest eum coinquinare,
MARK|7|19|quia non introit in cor eius sed in ventrem et in secessum exit? ", purgans omnes escas.
MARK|7|20|Dicebat autem: " Quod de homine exit, illud coinquinat hominem;
MARK|7|21|ab intus enim de corde hominum cogitationes malae procedunt, fornicationes, furta, homicidia,
MARK|7|22|adulteria, avaritiae, nequitiae, dolus, impudicitia, oculus malus, blasphemia, superbia, stultitia:
MARK|7|23|omnia haec mala ab intus procedunt et coinquinant hominem ".
MARK|7|24|Inde autem surgens abiit in fines Tyri et Sidonis. Et ingressus domum neminem voluit scire et non potuit latere.
MARK|7|25|Sed statim ut audivit de eo mulier, cuius habebat filia spiritum immundum, veniens procidit ad pedes eius.
MARK|7|26|Erat autem mulier Graeca, Syrophoenissa genere. Et rogabat eum, ut daemonium eiceret de filia eius.
MARK|7|27|Et dicebat illi: " Sine prius saturari filios; non est enim bonum sumere panem filiorum et mittere catellis ".
MARK|7|28|At illa respondit et dicit ei: " Domine, etiam catelli sub mensa comedunt de micis puerorum ".
MARK|7|29|Et ait illi: " Propter hunc sermonem vade; exiit daemonium de filia tua.
MARK|7|30|Et cum abisset domum suam, invenit puellam iacentem supra lectum et daemonium exisse.
MARK|7|31|Et iterum exiens de finibus Tyri venit per Sidonem ad mare Galilaeae inter medios fines Decapoleos.
MARK|7|32|Et adducunt ei surdum et mutum et deprecantur eum, ut imponat illi manum.
MARK|7|33|Et apprehendens eum de turba seorsum misit digitos suos in auriculas eius et exspuens tetigit linguam eius
MARK|7|34|et suspiciens in caelum ingemuit et ait illi: " Effetha ", quod est: " Adaperire ".
MARK|7|35|Et statim apertae sunt aures eius, et solutum est vinculum linguae eius, et loquebatur recte.
MARK|7|36|Et praecepit illis, ne cui dicerent; quanto autem eis praecipiebat, tanto magis plus praedicabant.
MARK|7|37|Et eo amplius admirabantur dicentes: " Bene omnia fecit, et surdos facit audire et mutos loqui! ".
MARK|8|1|In illis diebus iterum cum turba multa esset nec haberent, quod manducarent, convocatis discipulis, ait illis:
MARK|8|2|" Misereor super turbam, quia iam triduo sustinent me nec habent, quod manducent;
MARK|8|3|et si dimisero eos ieiunos in domum suam, deficient in via; et quidam ex eis de longe venerunt ".
MARK|8|4|Et responderunt ei discipuli sui: " Unde istos poterit quis hic saturare panibus in solitudine? ".
MARK|8|5|Et interrogabat eos: " Quot panes habetis? ". Qui dixerunt: " Septem ".
MARK|8|6|Et praecipit turbae discumbere supra terram; et accipiens septem panes, gratias agens fregit et dabat discipulis suis, ut apponerent; et apposuerunt turbae.
MARK|8|7|Et habebant pisciculos paucos; et benedicens eos, iussit hos quoque apponi.
MARK|8|8|Et manducaverunt et saturati sunt; et sustulerunt, quod superaverat de fragmentis, septem sportas.
MARK|8|9|Erant autem quasi quattuor milia. Et dimisit eos.
MARK|8|10|Et statim ascendens navem cum discipulis suis venit in partes Dalmanutha.
MARK|8|11|Et exierunt pharisaei et coeperunt conquirere cum eo quaerentes ab illo signum de caelo, tentantes eum.
MARK|8|12|Et ingemiscens spiritu suo ait: " Quid generatio ista quaerit signum? Amen dico vobis: Non dabitur generationi isti signum ".
MARK|8|13|Et dimittens eos, iterum ascendens abiit trans fretum.
MARK|8|14|Et obliti sunt sumere panes et nisi unum panem non habebant secum in navi.
MARK|8|15|Et praecipiebat eis dicens: " Videte, cavete a fermento pharisaeorum et fermento Herodis! ".
MARK|8|16|Et disputabant ad invicem, quia panes non haberent.
MARK|8|17|Quo cognito, ait illis: " Quid disputatis, quia panes non habetis? Nondum cognoscitis nec intellegitis? Caecatum habetis cor vestrum?
MARK|8|18|Oculos habentes non videtis, et aures habentes non auditis? Nec recordamini,
MARK|8|19|quando quinque panes fregi in quinque milia, quot cophinos fragmentorum plenos sustulistis? ". Dicunt ei: " Duodecim ".
MARK|8|20|" Quando illos septem in quattuor milia, quot sportas plenas fragmentorum tulistis? ". Et dicunt ei: " Septem ".
MARK|8|21|Et dicebat eis: " Nondum intellegitis? ".
MARK|8|22|Et veniunt Bethsaida. Et adducunt ei caecum et rogant eum, ut illum tangat.
MARK|8|23|Et apprehendens manum caeci eduxit eum extra vicum; et exspuens in oculos eius, impositis manibus ei, interrogabat eum: " Vides aliquid? ".
MARK|8|24|Et aspiciens dicebat: " Video homines, quia velut arbores video ambulantes ".
MARK|8|25|Deinde iterum imposuit manus super oculos eius; et coepit videre et restitutus est et videbat clare omnia.
MARK|8|26|Et misit illum in domum suam dicens: " Nec in vicum introieris ".
MARK|8|27|Et egressus est Iesus et discipuli eius in castella Caesareae Philippi; et in via interrogabat discipulos suos dicens eis: " Quem me dicunt esse homines? ".
MARK|8|28|Qui responderunt illi dicentcs: " Ioannem Baptistam, alii Eliam, alii vero unum de prophetis ".
MARK|8|29|Et ipse interrogabat eos: " Vos vero quem me dicitis esse? ". Respondens Petrus ait ei: " Tu es Christus ".
MARK|8|30|Et comminatus est eis, ne cui dicerent de illo.
MARK|8|31|Et coepit docere illos: " Oportet Filium hominis multa pati et reprobari a senioribus et a summis sacerdotibus et scribis et occidi et post tres dies resurgere ";
MARK|8|32|et palam verbum loquebatur. Et apprehendens eum Petrus coepit increpare eum.
MARK|8|33|Qui conversus et videns discipulos suos comminatus est Petro et dicit: Vade retro me, Satana, quoniam non sapis, quae Dei sunt, sed quae sunt hominum ".
MARK|8|34|Et convocata turba cum discipulis suis, dixit eis: " Si quis vult post me sequi, deneget semetipsum et tollat crucem suam et sequatur me.
MARK|8|35|Qui enim voluerit animam suam salvam facere, perdet eam; qui autem perdiderit animam suam propter me et evangelium, salvam eam faciet.
MARK|8|36|Quid enim prodest homini, si lucretur mundum totum et detrimentum faciat animae suae?
MARK|8|37|Quid enim dabit homo commutationem pro anima sua?
MARK|8|38|Qui enim me confusus fuerit et mea verba in generatione ista adultera et peccatrice, et Filius hominis confundetur eum, cum venerit in gloria Patris sui cum angelis sanctis ".
MARK|9|1|Et dicebat illis: " Amen dico vobis: Sunt quidam de hic stan tibus, qui non gustabunt mortem, donec videant regnum Dei venisse in virtute ".
MARK|9|2|Et post dies sex assumit Iesus Petrum et Iacobum et Ioannem, et ducit illos in montem excelsum seorsum solos. Et transfiguratus est coram ipsis;
MARK|9|3|et vestimenta eius facta sunt splendentia, candida nimis, qualia fullo super terram non potest tam candida facere.
MARK|9|4|Et apparuit illis Elias cum Moyse, et erant loquentes cum Iesu.
MARK|9|5|Et respondens Petrus ait Iesu: " Rabbi, bonum est nos hic esse; et faciamus tria tabernacula: tibi unum et Moysi unum et Eliae unum ".
MARK|9|6|Non enim sciebat quid responderet; erant enim exterriti.
MARK|9|7|Et facta est nubes obumbrans eos, et venit vox de nube: " Hic est Filius meus dilectus; audite illum ".
MARK|9|8|Et statim circumspicientes neminem amplius viderunt nisi Iesum tantum secum.
MARK|9|9|Et descendentibus illis de monte, praecepit illis, ne cui, quae vidissent, narrarent, nisi cum Filius hominis a mortuis resurrexerit.
MARK|9|10|Et verbum continuerunt apud se, conquirentes quid esset illud: " a mortuis resurgere ".
MARK|9|11|Et interrogabant eum dicentes: " Quid ergo dicunt scribae quia Eliam oporteat venire primum? ".
MARK|9|12|Qui ait illis: " Elias veniens primo, restituit omnia; et quomodo scriptum est super Filio hominis, ut multa patiatur et contemnatur?
MARK|9|13|Sed dico vobis: Et Elias venit; et fecerunt illi, quaecumque volebant, sicut scriptum est de eo ".
MARK|9|14|Et venientes ad discipulos viderunt turbam magnam circa eos et scribas conquirentes cum illis.
MARK|9|15|Et confestim omnis populus videns eum stupefactus est, et accurrentes salutabant eum.
MARK|9|16|Et interrogavit eos: " Quid inter vos conquiritis? ".
MARK|9|17|Et respondit ei unus de turba: " Magister, attuli filium meum ad te habentem spiritum mutum;
MARK|9|18|et ubicumque eum apprehenderit, allidit eum, et spumat et stridet dentibus et arescit. Et dixi discipulis tuis, ut eicerent illum, et non potuerunt ".
MARK|9|19|Qui respondens eis dicit: " O generatio incredula, quamdiu apud vos ero? Quamdiu vos patiar? Afferte illum ad me ".
MARK|9|20|Et attulerunt illum ad eum. Et cum vidisset illum, spiritus statim conturbavit eum; et corruens in terram volutabatur spumans.
MARK|9|21|Et interrogavit patrem eius: " Quantum temporis est, ex quo hoc ei accidit? ". At ille ait: " Ab infantia;
MARK|9|22|et frequenter eum etiam in ignem et in aquas misit, ut eum perderet; sed si quid potes, adiuva nos, misertus nostri ".
MARK|9|23|Iesus autem ait illi: " "Si potes!". Omnia possibilia credenti ".
MARK|9|24|Et continuo exclamans pater pueri aiebat: " Credo; adiuva incredulitatem meam ".
MARK|9|25|Et cum videret Iesus concurrentem turbam, comminatus est spiritui immundo dicens illi: " Mute et surde spiritus, ego tibi praecipio: Exi ab eo et amplius ne introeas in eum ".
MARK|9|26|Et clamans et multum discerpens eum exiit; et factus est sicut mortuus, ita ut multi dicerent: " Mortuus est! ".
MARK|9|27|Iesus autem tenens manum eius elevavit illum, et surrexit.
MARK|9|28|Et cum introisset in domum, discipuli eius secreto interrogabant eum: " Quare nos non potuimus eicere eum? ".
MARK|9|29|Et dixit illis: " Hoc genus in nullo potest exire nisi in oratione ".
MARK|9|30|Et inde profecti peragrabant Galilaeam; nec volebat quemquam scire.
MARK|9|31|Docebat enim discipulos suos et dicebat illis: " Filius hominis traditur in manus hominum, et occident eum, et occisus post tres dies resurget ".
MARK|9|32|At illi ignorabant verbum et timebant eum interrogare.
MARK|9|33|Et venerunt Capharnaum. Qui cum domi esset, interrogabat eos: " Quid in via tractabatis? ".
MARK|9|34|At illi tacebant. Siquidem inter se in via disputaverant, quis esset maior.
MARK|9|35|Et residens vocavit Duodecim et ait illis: " Si quis vult primus esse, erit omnium novissimus et omnium minister ".
MARK|9|36|Et accipiens puerum, statuit eum in medio eorum; quem ut complexus esset, ait illis:
MARK|9|37|" Quisquis unum ex huiusmodi pueris receperit in nomine meo, me recipit; et, quicumque me susceperit, non me suscipit, sed eum qui me misit ".
MARK|9|38|Dixit illi Ioannes: " Magister, vidimus quendam in nomine tuo eicientem daemonia, et prohibebamus eum, quia non sequebatur nos ".
MARK|9|39|Iesus autem ait: " Nolite prohibere eum. Nemo est enim, qui faciat virtutem in nomine meo et possit cito male loqui de me;
MARK|9|40|qui enim non est adversum nos, pro nobis est.
MARK|9|41|Quisquis enim potum dederit vobis calicem aquae in nomine, quia Christi estis, amen dico vobis: Non perdet mercedem suam.
MARK|9|42|Et quisquis scandalizaverit unum ex his pusillis credentibus in me, bonum est ei magis, ut circumdetur mola asinaria collo eius, et in mare mittatur.
MARK|9|43|Et si scandalizaverit te manus tua, abscide illam: bonum est tibi debilem introire in vitam, quam duas manus habentem ire ingehennam, in ignem inexstinguibilem.
MARK|9|44|()
MARK|9|45|Et si pes tuus te scandalizat, amputa illum: bonum est tibi claudum introire in vitam,quam duos pedes habentem mitti in gehennam.
MARK|9|46|()
MARK|9|47|Et si oculus tuus scandalizat te, eice eum: bonum est tibi luscum introire in regnum Dei, quam duos oculos habentem mitti in gehennam,
MARK|9|48|ubi vermis eorum non moritur, et ignis non exstinguitur;
MARK|9|49|omnis enim igne salietur.
MARK|9|50|Bonum est sal; quod si sal insulsum fuerit, in quo illud condietis? Habete in vobis sal et pacem habete inter vos ".
MARK|10|1|Et inde exsurgens venit in fines Iudaeae ultra Iorda nem; et conveniunt iterum turbae ad eum, et, sicut consueverat, iterum docebat illos.
MARK|10|2|Et accedentes pharisaei interrogabant eum, si licet viro uxorem dimittere, tentantes eum.
MARK|10|3|At ille respondens dixit eis: " Quid vobis praecepit Moyses? ".
MARK|10|4|Qui dixerunt: " Moyses permisit libellum repudii scribere et dimittere.
MARK|10|5|Iesus autem ait eis: " Ad duritiam cordis vestri scripsit vobis praeceptum istud.
MARK|10|6|Ab initio autem creaturae masculum et feminam fecit eos.
MARK|10|7|Propter hoc relinquet homo patrem suum et matrem et adhaerebit ad uxorern suam,
MARK|10|8|et erunt duo in carne una; itaque iam non sunt duo sed una caro.
MARK|10|9|Quod ergo Deus coniunxit, homo non separet ".
MARK|10|10|Et domo iterum discipuli de hoc interrogabant eum.
MARK|10|11|Et dicit illis: " Quicumque dimiserit uxorem suam et aliam duxerit, adulterium committit in eam;
MARK|10|12|et si ipsa dimiserit virum suum et alii nupserit, moechatur ".
MARK|10|13|Et offerebant illi parvulos, ut tangeret illos; discipuli autem comminabantur eis.
MARK|10|14|At videns Iesus, indigne tulit et ait illis: " Sinite parvulos venire ad me. Ne prohibueritis eos; talium est enim regnum Dei.
MARK|10|15|Amen dico vobis: Quisquis non receperit regnum Dei velut parvulus, non intrabit in illud ".
MARK|10|16|Et complexans eos benedicebat imponens manus super illos.
MARK|10|17|Et cum egrederetur in viam, accurrens quidam et, genu flexo ante eum, rogabat eum: " Magister bone, quid faciam ut vitam aeternam percipiam? ".
MARK|10|18|Iesus autem dixit ei: " Quid me dicis bonum? Nemo bonus, nisi unus Deus.
MARK|10|19|Praecepta nosti: ne occidas, ne adulteres, ne fureris, ne falsum testimonium dixeris, ne fraudem feceris, honora patrem tuum et matrem ".
MARK|10|20|Ille autem dixit ei: " Magister, haec omnia conservavi a iuventute mea.
MARK|10|21|Iesus autem intuitus eum dilexit eum et dixit illi: " Unum tibi deest: vade, quaecumque habes, vende et da pauperibus et habebis thesaurum in caelo; et veni, sequere me ".
MARK|10|22|Qui contristatus in hoc verbo, abiit maerens: erat enim habens possessiones multas.
MARK|10|23|Et circumspiciens Iesus ait discipulis suis: " Quam difficile, qui pecunias habent, in regnum Dei introibunt ".
MARK|10|24|Discipuli autem obstupescebant in verbis eius. At Iesus rursus respondens ait illis: " Filii, quam diffficile est in regnum Dei introire.
MARK|10|25|Facilius est camelum per foramen acus transire quam divitem intrare in regnum Dei ".
MARK|10|26|Qui magis admirabantur dicentes ad semetipsos: " Et quis potest salvus fieri? ".
MARK|10|27|Intuens illos Iesus ait: " Apud homines impossibile est sed non apud Deum: omnia enim possibilia sunt apud Deum ".
MARK|10|28|Coepit Petrus ei dicere: " Ecce nos dimisimus omnia et secuti sumus te.
MARK|10|29|Ait Iesus: " Amen dico vobis: Nemo est, qui reliquerit domum aut fratres aut sorores aut matrem aut patrem aut filios aut agros propter me et propter evangelium,
MARK|10|30|qui non accipiat centies tantum nunc in tempore hoc, domos et fratres et sorores et matres et filios et agros cum persecutionibus, et in saeculo futuro vitam aeternam.
MARK|10|31|Multi autem erunt primi novissimi, et novissimi primi ".
MARK|10|32|Erant autem in via ascendentes in Hierosolymam, et praecedebat illos Iesus, et stupebant; illi autem sequentes timebant. Et assumens iterum Duodecim coepit illis dicere, quae essent ei eventura:
MARK|10|33|" Ecce ascendimus in Hierosolymam; et Filius hominis tradetur principibus sacerdotum et scribis, et damnabunt eum morte et tradent eum gentibus
MARK|10|34|et illudent ei et conspuent eum et flagellabunt eum et interficient eum, et post tres dies resurget ".
MARK|10|35|Et accedunt ad eum Iacobus et Ioannes filii Zebedaei dicentes ei: " Magister, volumus, ut quodcumque petierimus a te, facias nobis ".
MARK|10|36|At ille dixit eis: " Quid vultis, ut faciam vobis? ".
MARK|10|37|Illi autem dixerunt ei: " Da nobis, ut unus ad dexteram tuam et alius ad sinistram sedeamus in gloria tua ".
MARK|10|38|Iesus autem ait eis: " Nescitis quid petatis. Potestis bibere calicem, quem ego bibo, aut baptismum, quo ego baptizor, baptizari? ".
MARK|10|39|At illi dixerunt ei: " Possumus ". Iesus autem ait eis: " Calicem quidem, quem ego bibo, bibetis et baptismum, quo ego baptizor, baptizabimini;
MARK|10|40|sedere autem ad dexteram meam vel ad sinistram non est meum dare, sed quibus paratum est ".
MARK|10|41|Et audientes decem coeperunt indignari de Iacobo et Ioanne.
MARK|10|42|Et vocans eos Iesus ait illis: " Scitis quia hi, qui videntur principari gentibus, dominantur eis, et principes eorum potestatem habent ipsorum.
MARK|10|43|Non ita est autem in vobis, sed quicumque voluerit fieri maior inter vos, erit vester minister;
MARK|10|44|et, quicumque voluerit in vobis primus esse, erit omnium servus;
MARK|10|45|nam et Filius hominis non venit, ut ministraretur ei, sed ut ministraret et daret animam suam redemptionem pro multis ".
MARK|10|46|Et veniunt Ierichum. Et proficiscente eo de Iericho et discipulis eius et plurima multitudine, filius Timaei Bartimaeus caecus sedebat iuxta viam mendicans.
MARK|10|47|Qui cum audisset quia Iesus Nazarenus est, coepit clamare et dicere: " Fili David Iesu, miserere mei! ".
MARK|10|48|Et comminabantur ei multi, ut taceret; at ille multo magis clamabat: " Fili David, miserere mei! ".
MARK|10|49|Et stans Iesus dixit: " Vocate illum ". Et vocant caecum dicentes ei: " Animaequior esto. Surge, vocat te ".
MARK|10|50|Qui, proiecto vestimento suo, exsiliens venit ad Iesum.
MARK|10|51|Et respondens ei Iesus dixit: " Quid vis tibi faciam? ". Caecus autem dixit ei: " Rabboni, ut videam ".
MARK|10|52|Et Iesus ait illi: " Vade; fides tua te salvum fecit ". Et confestim vidit et sequebatur eum in via.
MARK|11|1|Et cum appropinquarent Hierosolymae, Bethphage et Bethaniae ad montem Olivarum, mittit duos ex discipulis suis
MARK|11|2|et ait illis: " Ite in castellum, quod est contra vos, et statim introeuntes illud invenietis pullum ligatum, super quem nemo adhuc hominum sedit; solvite illum et adducite.
MARK|11|3|Et si quis vobis dixerit: "Quid facitis hoc?", dicite: "Domino necessarius est, et continuo illum remittit iterum huc" ".
MARK|11|4|Et abeuntes invenerunt pullum ligatum ante ianuam foris in bivio et solvunt eum.
MARK|11|5|Et quidam de illic stantibus dicebant illis: " Quid facitis solventes pullum? ".
MARK|11|6|Qui dixerunt eis, sicut dixerat Iesus; et dimiserunt eis.
MARK|11|7|Et ducunt pullum ad Iesum et imponunt illi vestimenta sua; et sedit super eum.
MARK|11|8|Et multi vestimenta sua straverunt in via, alii autem frondes, quas exciderant in agris.
MARK|11|9|Et qui praeibant et qui sequebantur, clamabant: " Hosanna! Benedictus, qui venit in nomine Domini!
MARK|11|10|Benedictum, quod venit regnum patris nostri David! Hosanna in excelsis!.
MARK|11|11|Et introivit Hierosolymam in templum; et circumspectis omnibus, cum iam vespera esset hora, exivit in Bethaniam cum Duodecim.
MARK|11|12|Et altera die cum exirent a Bethania, esuriit.
MARK|11|13|Cumque vidisset a longe ficum habentem folia, venit si quid forte inveniret in ea; et cum venisset ad eam, nihil invenit praeter folia: non enim erat tempus ficorum.
MARK|11|14|Et respondens dixit ei: " Iam non amplius in aeternum quisquam fructum ex te manducet ". Et audiebant discipuli eius.
MARK|11|15|Et veniunt Hierosolymam. Et cum introisset in templum, coepit eicere vendentes et ementes in templo et mensas nummulariorum et cathedras vendentium columbas evertit;
MARK|11|16|et non sinebat, ut quisquam vas transferret per templum.
MARK|11|17|Et docebat dicens eis: " Non scriptum est: "Domus mea domus orationis vocabitur omnibus gentibus"? Vos autem fecistis eam speluncam latronum ".
MARK|11|18|Quo audito, principes sacerdotum et scribae quaerebant quomodo eum perderent; timebant enim eum, quoniam universa turba admirabatur super doctrina eius.
MARK|11|19|Et cum vespera facta esset, egrediebantur de civitate.
MARK|11|20|Et cum mane transirent, viderunt ficum aridam factam a radicibus.
MARK|11|21|Et recordatus Petrus dicit ei: " Rabbi, ecce ficus, cui maledixisti, aruit ".
MARK|11|22|Et respondens Iesus ait illis: " Habete fidem Dei!
MARK|11|23|Amen dico vobis: Quicumque dixerit huic monti: "Tollere et mittere in mare", et non haesitaverit in corde suo, sed crediderit quia, quod dixerit, fiat, fiet ei.
MARK|11|24|Propterea dico vobis: Omnia, quaecumque orantes petitis, credite quia iam accepistis, et erunt vobis.
MARK|11|25|Et cum statis in oratione, dimittite, si quid habetis adversus aliquem, ut etPater vester, qui in caelis est, dimittat vobis peccata vestra ".
MARK|11|26|()
MARK|11|27|Et veniunt rursus Hierosolymam. Et cum ambularet in templo, accedunt ad eum summi sacerdotes et scribae et seniores
MARK|11|28|et dicebant illi: " In qua potestate haec facis? Vel quis tibi dedit hanc potestatem, ut ista facias? ".
MARK|11|29|Iesus autem ait illis: " Interrogabo vos unum verbum, et respondete mihi; et dicam vobis, in qua potestate haec faciam:
MARK|11|30|Baptismum Ioannis de caelo erat an ex hominibus? Respondete mihi ".
MARK|11|31|At illi cogitabant secum dicentes: " Si dixerimus: "De caelo", dicet: Quare ergo non credidistis ei?";
MARK|11|32|si autem dixerimus: "Ex hominibus?" ". Timebant populum: omnes enim habebant Ioannem quia vere propheta esset.
MARK|11|33|Et respondentes dicunt Iesu: " Nescimus ". Et Iesus ait illis: " Neque ego dico vobis in qua potestate haec faciam ".
MARK|12|1|Et coepit illis in parabolis loqui: " Vineam pastinavit ho mo et circumdedit saepem et fodit lacum et aedificavit turrim et locavit eam agricolis et peregre profectus est.
MARK|12|2|Et misit ad agricolas in tempore servum, ut ab agricolis acciperet de fructu vineae;
MARK|12|3|qui apprehensum eum caeciderunt et dimiserunt vacuum.
MARK|12|4|Et iterum misit ad illos alium servum; et illum in capite vulneraverunt et contumeliis affecerunt.
MARK|12|5|Et alium misit, et illum occiderunt, et plures alios, quosdam caedentes, alios vero occidentes.
MARK|12|6|Adhuc unum habebat, filium dilectum. Misit illum ad eos novissimum dicens: "Reverebuntur filium meum".
MARK|12|7|Coloni autem illi dixerunt ad invicem: "Hic est heres. Venite, occidamus eum, et nostra erit hereditas".
MARK|12|8|Et apprehendentes eum occiderunt et eiecerunt extra vineam.
MARK|12|9|Quid ergo faciet dominus vineae? Veniet et perdet colonos et dabit vineam aliis.
MARK|12|10|Nec Scripturam hanc legistis: "Lapidem quem reprobaverunt aedificantes,hic factus est in caput anguli;
MARK|12|11|a Domino factum est istudet est mirabile in oculis nostris"? ".
MARK|12|12|Et quaerebant eum tenere et timuerunt turbam; cognoverunt enim quoniam ad eos parabolam hanc dixerit. Et relicto eo abierunt.
MARK|12|13|Et mittunt ad eum quosdam ex pharisaeis et herodianis, ut eum caperent in verbo.
MARK|12|14|Qui venientes dicunt ei: " Magister, scimus quia verax es et non curas quemquam; nec enim vides in faciem hominum, sed in veritate viam Dei doces. Licet dare tributum Caesari an non? Dabimus an non dabimus? ".
MARK|12|15|Qui sciens versutiam eorum ait illis: " Quid me tentatis? Afferte mihi denarium, ut videam ".
MARK|12|16|At illi attulerunt. Et ait illis: " Cuius est imago haec et inscriptio?. Illi autem dixerunt ei: " Caesaris ".
MARK|12|17|Iesus autem dixit illis: " Quae sunt Caesaris, reddite Caesari et, quae sunt Dei, Deo ". Et mirabantur super eo.
MARK|12|18|Et veniunt ad eum sadducaei, qui dicunt resurrectionem non esse, et interrogabant eum dicentes:
MARK|12|19|" Magister, Moyses nobis scripsit, ut si cuius frater mortuus fuerit et reliquerit uxorem et filium non reliquerit, accipiat frater eius uxorem et resuscitet semen fratri suo.
MARK|12|20|Septem fratres erant: et primus accepit uxorem et moriens non reliquit semen;
MARK|12|21|et secundus accepit eam et mortuus est, non relicto semine; et tertius similiter;
MARK|12|22|et septem non reliquerunt semen. Novissima omnium defuncta est et mulier.
MARK|12|23|In resurrectione, cum resurrexerint, cuius de his erit uxor? Septem enim habuerunt eam uxorem ".
MARK|12|24|Ait illis Iesus: " Non ideo erratis, quia non scitis Scripturas neque virtutem Dei?
MARK|12|25|Cum enim a mortuis resurrexerint, neque nubent neque nubentur, sed sunt sicut angeli in caelis.
MARK|12|26|De mortuis autem quod resurgant, non legistis in libro Moysis super rubum, quomodo dixerit illi Deus inquiens: "Ego sum Deus Abraham et Deus Isaac et Deus Iacob"?
MARK|12|27|Non est Deus mortuorum sed vivorum! Multum erratis ".
MARK|12|28|Et accessit unus de scribis, qui audierat illos conquirentes, videns quoniam bene illis responderit, interrogavit eum: " Quod est primum omnium mandatum? ".
MARK|12|29|Iesus respondit: " Primum est: "Audi, Israel: Dominus Deus noster Dominus unus est,
MARK|12|30|et diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex tota mente tua et ex tota virtute tua".
MARK|12|31|Secundum est illud: "Diliges proximum tuum tamquam teipsum". Maius horum aliud mandatum non est ".
MARK|12|32|Et ait illi scriba: " Bene, Magister, in veritate dixisti: "Unus est, et non est alius praeter eum;
MARK|12|33|et diligere eum ex toto corde et ex toto intellectu et ex tota fortitudine" et: "Diligere proximum tamquam seipsum" maius est omnibus holocautomatibus et sacrificiis ".
MARK|12|34|Et Iesus videns quod sapienter respondisset, dixit illi: " Non es longe a regno Dei ". Et nemo iam audebat eum interrogare.
MARK|12|35|Et respondens Iesus dicebat docens in templo: " Quomodo dicunt scribae Christum filium esse David?
MARK|12|36|Ipse David dixit in Spiritu Sancto:Dixit Dominus Domino meo: Sede a dextris meis,donec ponam inimicos tuos sub pedibus tuis".
MARK|12|37|Ipse David dicit eum Dominum, et unde est filius eius? ". Et multa turba eum libenter audiebat.
MARK|12|38|Et dicebat in doctrina sua: " Cavete a scribis, qui volunt in stolis ambulare et salutari in foro
MARK|12|39|et in primis cathedris sedere in synagogis et primos discubitus in cenis;
MARK|12|40|qui devorant domos viduarum et ostentant prolixas orationes. Hi accipient amplius iudicium ".
MARK|12|41|Et sedens contra gazophylacium aspiciebat quomodo turba iactaret aes in gazophylacium; et multi divites iactabant multa.
MARK|12|42|Et cum venisset una vidua pauper, misit duo minuta, quod est quadrans.
MARK|12|43|Et convocans discipulos suos ait illis: " Amen dico vobis: Vidua haec pauper plus omnibus misit, qui miserunt in gazophylacium:
MARK|12|44|Omnes enim ex eo, quod abundabat illis, miserunt; haec vero de penuria sua omnia, quae habuit, misit, totum victum suum ".
MARK|13|1|Et cum egrederetur de tem plo, ait illi unus ex discipulis suis: " Magister, aspice quales lapides et quales structurae ".
MARK|13|2|Et Iesus ait illi: " Vides has magnas aedificationes? Hic non relinquetur lapis super lapidem, qui non destruatur ".
MARK|13|3|Et cum sederet in montem Olivarum contra templum, interrogabat eum separatim Petrus et Iacobus et Ioannes et Andreas:
MARK|13|4|" Dic nobis: Quando ista erunt, et quod signum erit, quando haec omnia incipient consummari? ".
MARK|13|5|Iesus autem coepit dicere illis: " Videte, ne quis vos seducat.
MARK|13|6|Multi venient in nomine meo dicentes: "Ego sum", et multos seducent.
MARK|13|7|Cum audieritis autem bella et opiniones bellorum, ne timueritis; oportet fieri sed nondum finis.
MARK|13|8|Exsurget enim gens super gentem, et regnum super regnum, erunt terrae motus per loca, erunt fames; initium dolorum haec.
MARK|13|9|Videte autem vosmetipsos. Tradent vos conciliis, et in synagogis vapulabitis et ante praesides et reges stabitis propter me in testimonium illis.
MARK|13|10|Et in omnes gentes primum oportet praedicari evangelium.
MARK|13|11|Et cum duxerint vos tradentes, nolite praecogitare quid loquamini, sed, quod datum vobis fuerit in illa hora, id loquimini: non enim estis vos loquentes sed Spiritus Sanctus.
MARK|13|12|Et tradet frater fratrem in mortem, et pater filium; et consurgent filii in parentes et morte afficient eos;
MARK|13|13|et eritis odio omnibus propter nomen meum. Qui autem sustinuerit in finem, hic salvus erit.
MARK|13|14|Cum autem videritis abominationem desolationis stantem, ubi non debet, qui legit, intellegat: tunc, qui in Iudaea sunt, fugiant in montes;
MARK|13|15|qui autem super tectum, ne descendat nec introeat, ut tollat quid de domo sua;
MARK|13|16|et, qui in agro erit, non revertatur retro tollere vestimentum suum.
MARK|13|17|Vae autem praegnantibus et nutrientibus in illis diebus!
MARK|13|18|Orate vero, ut hieme non fiat:
MARK|13|19|erunt enim dies illi tribulatio talis, qualis non fuit ab initio creaturae, quam condidit Deus, usque nunc, neque fiet.
MARK|13|20|Et nisi breviasset Dominus dies, non fuisset salva omnis caro. Sed propter electos, quos elegit, breviavit dies.
MARK|13|21|Et tunc, si quis vobis dixerit: "Ecce hic est Christus, ecce illic", ne credideritis.
MARK|13|22|Exsurgent enim pseudochristi et pseudoprophetae et dabunt signa et portenta ad seducendos, si potest fieri, electos.
MARK|13|23|Vos autem videte; praedixi vobis omnia.
MARK|13|24|Sed in illis diebus post tribulationem illam sol contenebrabitur, et luna non dabit splendorem suum,
MARK|13|25|et erunt stellae de caelo decidentes, et virtutes, quae sunt in caelis, movebuntur.
MARK|13|26|Et tunc videbunt Filium hominis venientem in nubibus cum virtute multa et gloria.
MARK|13|27|Et tunc mittet angelos et congregabit electos suos a quattuor ventis, a summo terrae usque ad summum caeli.
MARK|13|28|A ficu autem discite parabolam: cum iam ramus eius tener fuerit et germinaverit folia, cognoscitis quia in proximo sit aestas.
MARK|13|29|Sic et vos, cum videritis haec fieri, scitote quod in proximo sit in ostiis.
MARK|13|30|Amen dico vobis: Non transiet generatio haec, donec omnia ista fiant.
MARK|13|31|Caelum et terra transibunt, verba autem mea non transibunt.
MARK|13|32|De die autem illo vel hora nemo scit, neque angeli in caelo neque Filius, nisi Pater.
MARK|13|33|Videte, vigilate; nescitis enim, quando tempus sit.
MARK|13|34|Sicut homo, qui peregre profectus reliquit domum suam et dedit servis suis potestatem, unicuique opus suum, ianitori quoque praecepit, ut vigilaret.
MARK|13|35|Vigilate ergo; nescitis enim quando dominus domus veniat, sero an media nocte an galli cantu an mane;
MARK|13|36|ne, cum venerit repente, inveniat vos dormientes.
MARK|13|37|Quod autem vobis dico, omnibus dico: Vigilate! ".
MARK|14|1|Erat autem Pascha et Azy ma post biduum. Et quaerebant summi sacerdotes et scribae, quomodo eum dolo tenerent et occiderent;
MARK|14|2|dicebant enim: " Non in die festo, ne forte tumultus fieret populi ".
MARK|14|3|Et cum esset Bethaniae in domo Simonis leprosi et recumberet, venit mulier habens alabastrum unguenti nardi puri pretiosi; fracto alabastro, effudit super caput eius.
MARK|14|4|Erant autem quidam indigne ferentes intra semetipsos: " Ut quid perditio ista unguenti facta est?
MARK|14|5|Poterat enim unguentum istud veniri plus quam trecentis denariis et dari pauperibus ". Et fremebant in eam.
MARK|14|6|Iesus autem dixit: " Sinite eam; quid illi molesti estis? Bonum opus operata est in me.
MARK|14|7|Semper enim pauperes habetis vobiscum et, cum volueritis, potestis illis bene facere; me autem non semper habetis.
MARK|14|8|Quod habuit, operata est: praevenit ungere corpus meum in sepulturam.
MARK|14|9|Amen autem dico vobis: Ubicumque praedicatum fuerit evangelium in universum mundum, et, quod fecit haec, narrabitur in memoriam eius ".
MARK|14|10|Et Iudas Iscarioth, unus de Duodecim, abiit ad summos sacerdotes, ut proderet eum illis.
MARK|14|11|Qui audientes gavisi sunt et promiserunt ei pecuniam se daturos. Et quaerebat quomodo illum opportune traderet.
MARK|14|12|Et primo die Azymorum, quando Pascha immolabant, dicunt ei discipuli eius: " Quo vis eamus et paremus, ut manduces Pascha? ".
MARK|14|13|Et mittit duos ex discipulis suis et dicit eis: " Ite in civitatem, et occurret vobis homo lagoenam aquae baiulans; sequimini eum
MARK|14|14|et, quocumque introierit, dicite domino domus: "Magister dicit: Ubi est refectio mea, ubi Pascha cum discipulis meis manducem?".
MARK|14|15|Et ipse vobis demonstrabit cenaculum grande stratum paratum; et illic parate nobis ".
MARK|14|16|Et abierunt discipuli et venerunt in civitatem et invenerunt, sicut dixerat illis, et paraverunt Pascha.
MARK|14|17|Et vespere facto, venit cum Duodecim.
MARK|14|18|Et discumbentibus eis et manducantibus, ait Iesus: " Amen dico vobis: Unus ex vobis me tradet, qui manducat mecum ".
MARK|14|19|Coeperunt contristari et dicere ei singillatim: " Numquid ego? ".
MARK|14|20|Qui ait illis: " Unus ex Duodecim, qui intingit mecum in catino.
MARK|14|21|Nam Filius quidem hominis vadit, sicut scriptum est de eo. Vae autem homini illi, per quem Filius hominis traditur! Bonum est ei, si non esset natus homo ille ".
MARK|14|22|Et manducantibus illis, accepit panem et benedicens fregit et dedit eis et ait: " Sumite: hoc est corpus meum ".
MARK|14|23|Et accepto calice, gratias agens dedit eis; et biberunt ex illo omnes.
MARK|14|24|Et ait illis: " Hic est sanguis meus novi testamenti, qui pro multis effunditur.
MARK|14|25|Amen dico vobis: Iam non bibam de genimine vitis usque in diem illum, cum illud bibam novum in regno Dei ".
MARK|14|26|Et hymno dicto, exierunt in montem Olivarum.
MARK|14|27|Et ait eis Iesus: " Omnes scandalizabimini, quia scriptum est: Percutiam pastorem, et dispergentur oves".
MARK|14|28|Sed posteaquam resurrexero, praecedam vos in Galilaeam ".
MARK|14|29|Petrus autem ait ei: " Et si omnes scandalizati fuerint, sed non ego ".
MARK|14|30|Et ait illi Iesus: " Amen dico tibi: Tu hodie, in nocte hac, priusquam bis gallus vocem dederit, ter me es negaturus ".
MARK|14|31|At ille amplius loquebatur: " Et si oportuerit me commori tibi, non te negabo ". Similiter autem et omnes dicebant.
MARK|14|32|Et veniunt in praedium, cui nomen Gethsemani; et ait discipulis suis: " Sedete hic, donec orem ".
MARK|14|33|Et assumit Petrum et Iacobum et Ioannem secum et coepit pavere et taedere;
MARK|14|34|et ait illis: " Tristis est anima mea usque ad mortem; sustinete hic et vigilate ".
MARK|14|35|Et cum processisset paululum, procidebat super terram et orabat, ut, si fieri posset, transiret ab eo hora;
MARK|14|36|et dicebat: " Abba, Pater! Omnia tibi possibilia sunt. Transfer calicem hunc a me; sed non quod ego volo, sed quod tu ".
MARK|14|37|Et venit et invenit eos dormientes; et ait Petro: " Simon, dormis? Non potuisti una hora vigilare?
MARK|14|38|Vigilate et orate, ut non intretis in tentationem; spiritus quidem promptus, caro vero infirma ".
MARK|14|39|Et iterum abiens oravit, eundem sermonem dicens.
MARK|14|40|Et veniens denuo invenit eos dormientes; erant enim oculi illorum ingravati, et ignorabant quid responderent ei.
MARK|14|41|Et venit tertio et ait illis: " Dormite iam et requiescite? Sufficit, venit hora: ecce traditur Filius hominis in manus peccatorum.
MARK|14|42|Surgite, eamus; ecce, qui me tradit, prope est ".
MARK|14|43|Et confestim, adhuc eo loquente, venit Iudas unus ex Duodecim, et cum illo turba cum gladiis et lignis a summis sacerdotibus et scribis et senioribus.
MARK|14|44|Dederat autem traditor eius signum eis dicens: " Quemcumque osculatus fuero, ipse est; tenete eum et ducite caute ".
MARK|14|45|Et cum venisset, statim accedens ad eum ait: " Rabbi "; et osculatus est eum.
MARK|14|46|At illi manus iniecerunt in eum et tenuerunt eum.
MARK|14|47|Unus autem quidam de circumstantibus educens gladium percussit servum summi sacerdotis et amputavit illi auriculam.
MARK|14|48|Et respondens Iesus ait illis: " Tamquam ad latronem existis cum gladiis et lignis comprehendere me?
MARK|14|49|Cotidie eram apud vos in templo docens, et non me tenuistis; sed adimpleantur Scripturae ".
MARK|14|50|Et relinquentes eum omnes fugerunt.
MARK|14|51|Et adulescens quidam sequebatur eum amictus sindone super nudo, et tenent eum;
MARK|14|52|at ille, reiecta sindone, nudus profugit.
MARK|14|53|Et adduxerunt Iesum ad summum sacerdotem; et conveniunt omnes summi sacerdotes et seniores et scribae.
MARK|14|54|Et Petrus a longe secutus est eum usque intro in atrium summi sacerdotis et sedebat cum ministris et calefaciebat se ad ignem.
MARK|14|55|Summi vero sacerdotes et omne concilium quaerebant adversus Iesum testimonium, ut eum morte afficerent, nec inveniebant.
MARK|14|56|Multi enim testimonium falsum dicebant adversus eum, et convenientia testimonia non erant.
MARK|14|57|Et quidam surgentes falsum testimonium ferebant adversus eum dicentes:
MARK|14|58|" Nos audivimus eum dicentem: "Ego dissolvam templum hoc manu factum et intra triduum aliud non manu factum aedificabo" ".
MARK|14|59|Et ne ita quidem conveniens erat testimonium illorum.
MARK|14|60|Et exsurgens summus sacerdos in medium interrogavit Iesum dicens: " Non respondes quidquam ad ea, quae isti testantur adversum te? ".
MARK|14|61|Ille autem tacebat et nihil respondit. Rursum summus sacerdos interrogabat eum et dicit ei: " Tu es Christus filius Benedicti? ".
MARK|14|62|Iesus autem dixit: " Ego sum, et videbitis Filium hominis a dextris sedentem Virtutis et venientem cum nubibus caeli ".
MARK|14|63|Summus autem sacerdos scindens vestimenta sua ait: " Quid adhuc necessarii sunt nobis testes?
MARK|14|64|Audistis blasphemiam. Quid vobis videtur? ". Qui omnes condemnaverunt eum esse reum mortis.
MARK|14|65|Et coeperunt quidam conspuere eum et velare faciem eius et colaphis eum caedere et dicere ei: " Prophetiza "; et ministri alapis eum caedebant.
MARK|14|66|Et cum esset Petrus in atrio deorsum, venit una ex ancillis summi sacerdotis
MARK|14|67|et, cum vidisset Petrum calefacientem se, aspiciens illum ait: " Et tu cum hoc Nazareno, Iesu, eras! ".
MARK|14|68|At ille negavit dicens: " Neque scio neque novi quid tu dicas! ". Et exiit foras ante atrium, et gallus cantavit.
MARK|14|69|Et ancilla, cum vidisset illum, rursus coepit dicere circumstantibus: " Hic ex illis est! ".
MARK|14|70|At ille iterum negabat. Et post pusillum rursus, qui astabant, dicebant Petro: " Vere ex illis es, nam et Galilaeus es ".
MARK|14|71|Ille autem coepit anathematizare et iurare: " Nescio hominem istum, quem dicitis! ".
MARK|14|72|Et statim iterum gallus cantavit; et recordatus est Petrus verbi, sicut dixerat ei Iesus: " Priusquam gallus cantet bis, ter me negabis ". Et coepit flere.
MARK|15|1|Et confestim mane consilium facientes summi sacerdotes cum senioribus et scribis, id est universum concilium, vincientes Iesum duxerunt et tradiderunt Pilato.
MARK|15|2|Et interrogavit eum Pilatus: " Tu es rex Iudaeorum? ". At ille respondens ait illi: " Tu dicis ".
MARK|15|3|Et accusabant eum summi sacerdotes in multis.
MARK|15|4|Pilatus autem rursum interrogabat eum dicens: " Non respondes quidquam? Vide in quantis te accusant ".
MARK|15|5|Iesus autem amplius nihil respondit, ita ut miraretur Pilatus.
MARK|15|6|Per diem autem festum dimittere solebat illis unum ex vinctis, quem peterent.
MARK|15|7|Erat autem qui dicebatur Barabbas, vinctus cum seditiosis, qui in seditione fecerant homicidium.
MARK|15|8|Et cum ascendisset turba, coepit rogare, sicut faciebat illis.
MARK|15|9|Pilatus autem respondit eis et dixit: " Vultis dimittam vobis regem Iudaeorum? ".
MARK|15|10|Sciebat enim quod per invidiam tradidissent eum summi sacerdotes.
MARK|15|11|Pontifices autem concitaverunt turbam, ut magis Barabbam dimitteret eis.
MARK|15|12|Pilatus autem iterum respondens aiebat illis: " Quid ergo vultis faciam regi Iudaeorum? ".
MARK|15|13|At illi iterum clamaverunt: " Crucifige eum! ".
MARK|15|14|Pilatus vero dicebat eis: " Quid enim mali fecit? ". At illi magis clamaverunt: " Crucifige eum! ".
MARK|15|15|Pilatus autem, volens populo satisfacere, dimisit illis Barabbam et tradidit Iesum flagellis caesum, ut crucifigeretur.
MARK|15|16|Milites autem duxerunt eum intro in atrium, quod est praetorium, et convocant totam cohortem.
MARK|15|17|Et induunt eum purpuram et imponunt ei plectentes spineam coronam;
MARK|15|18|et coeperunt salutare eum: " Ave, rex Iudaeorum! ",
MARK|15|19|et percutiebant caput eius arundine et conspuebant eum et ponentes genua adorabant eum.
MARK|15|20|Et postquam illuserunt ei, exuerunt illum purpuram et induerunt eum vestimentis suis. Et educunt illum, ut crucifigerent eum.
MARK|15|21|Et angariant praetereuntem quempiam Simonem Cyrenaeum venientem de villa, patrem Alexandri et Rufi, ut tolleret crucem eius.
MARK|15|22|Et perducunt illum in Golgotha locum, quod est interpretatum Calvariae locus.
MARK|15|23|Et dabant ei myrrhatum vinum; ille autem non accepit.
MARK|15|24|Et crucifigunt eum et dividunt vestimenta eius, mittentes sortem super eis, quis quid tolleret.
MARK|15|25|Erat autem hora tertia, et crucifixerunt eum.
MARK|15|26|Et erat titulus causae eius inscriptus: " Rex Iudaeorum ".
MARK|15|27|Et cum eo crucifigunt duos latrones, unum a dextris et alium asinistris eius.
MARK|15|28|()
MARK|15|29|Et praetereuntes blasphemabant eum moventes capita sua et dicentes: " Vah, qui destruit templum et in tribus diebus aedificat;
MARK|15|30|salvum fac temetipsum descendens de cruce! ".
MARK|15|31|Similiter et summi sacerdotes ludentes ad alterutrum cum scribis dicebant: " Alios salvos fecit, seipsum non potest salvum facere.
MARK|15|32|Christus rex Israel descendat nunc de cruce, ut videamus et credamus ". Etiam qui cum eo crucifixi erant, conviciabantur ei.
MARK|15|33|Et, facta hora sexta, tenebrae factae sunt per totam terram usque in horam nonam.
MARK|15|34|Et hora nona exclamavit Iesus voce magna: " Heloi, Heloi, lema sabacthani? ", quod est interpretatum: " Deus meus, Deus meus, ut quid dereliquisti me? ".
MARK|15|35|Et quidam de circumstantibus audientes dicebant: " Ecce, Eliam vocat ".
MARK|15|36|Currens autem unus et implens spongiam aceto circumponensque calamo potum dabat ei dicens: " Sinite, videamus, si veniat Elias ad deponendum eum ".
MARK|15|37|Iesus autem, emissa voce magna, exspiravit.
MARK|15|38|Et velum templi scissum est in duo a sursum usque deorsum.
MARK|15|39|Videns autem centurio, qui ex adverso stabat, quia sic clamans exspirasset, ait: " Vere homo hic Filius Dei erat ".
MARK|15|40|Erant autem et mulieres de longe aspicientes, inter quas et Maria Magdalene et Maria Iacobi minoris et Iosetis mater et Salome,
MARK|15|41|quae, cum esset in Galilaea, sequebantur eum et ministrabant ei, et aliae multae, quae simul cum eo ascenderant Hierosolymam.
MARK|15|42|Et cum iam sero esset factum, quia erat Parasceve, quod est ante sabbatum,
MARK|15|43|venit Ioseph ab Arimathaea nobilis decurio, qui et ipse erat exspectans regnum Dei, et audacter introivit ad Pilatum et petiit corpus Iesu.
MARK|15|44|Pilatus autem miratus est si iam obisset, et, accersito centurione, interrogavit eum si iam mortuus esset,
MARK|15|45|et, cum cognovisset a centurione, donavit corpus Ioseph.
MARK|15|46|Is autem mercatus sindonem et deponens eum involvit sindone et posuit eum in monumento, quod erat excisum de petra, et advolvit lapidem ad ostium monumenti.
MARK|15|47|Maria autem Magdalene et Maria Iosetis aspiciebant, ubi positus esset.
MARK|16|1|Et cum transisset sabbatum, Maria Magdalene et Maria Iacobi et Salome emerunt aromata, ut venientes ungerent eum.
MARK|16|2|Et valde mane, prima sabbatorum, veniunt ad monumentum, orto iam sole.
MARK|16|3|Et dicebant ad invicem: " Quis revolvet nobis lapidem ab ostio monumenti? ".
MARK|16|4|Et respicientes vident revolutum lapidem; erat quippe magnus valde.
MARK|16|5|Et introeuntes in monumentum viderunt iuvenem sedentem in dextris, coopertum stola candida, et obstupuerunt.
MARK|16|6|Qui dicit illis: " Nolite expavescere! Iesum quaeritis Nazarenum crucifixum. Surrexit, non est hic; ecce locus, ubi posuerunt eum.
MARK|16|7|Sed ite, dicite discipulis eius et Petro: "Praecedit vos in Galilaeam. Ibi eum videbitis, sicut dixit vobis" ".
MARK|16|8|Et exeuntes fugerunt de monumento; invaserat enim eas tremor et pavor, et nemini quidquam dixerunt, timebant enim.
MARK|16|9|Surgens autem mane, prima sabbati, apparuit primo Mariae Magdalenae, de qua eiecerat septem daemonia.
MARK|16|10|Illa vadens nuntiavit his, qui cum eo fuerant, lugentibus et flentibus;
MARK|16|11|et illi audientes quia viveret et visus esset ab ea, non crediderunt.
MARK|16|12|Post haec autem duobus ex eis ambulantibus ostensus est in alia effigie euntibus in villam;
MARK|16|13|et illi euntes nuntiaverunt ceteris, nec illis crediderunt.
MARK|16|14|Novissime recumbentibus illis Undecim apparuit, et exprobravit incredulitatem illorum et duritiam cordis, quia his, qui viderant eum resuscitatum, non crediderant.
MARK|16|15|Et dixit eis: " Euntes in mundum universum praedicate evangelium omni creaturae.
MARK|16|16|Qui crediderit et baptizatus fuerit, salvus erit; qui vero non crediderit, condemnabitur.
MARK|16|17|Signa autem eos, qui crediderint, haec sequentur: in nomine meo daemonia eicient, linguis loquentur novis,
MARK|16|18|serpentes tollent, et, si mortiferum quid biberint, non eos nocebit, super aegrotos manus imponent, et bene habebunt ".
MARK|16|19|Et Dominus quidem Iesus, postquam locutus est eis, assumptus est in caelum et sedit a dextris Dei.
MARK|16|20|Illi autem profecti praedicaverunt ubique, Domino cooperante et sermonem confirmante, sequentibus signis.
