1CHR|1|1|Adam, Seth, Enos,
1CHR|1|2|Cainan, Malaleel, Iared,
1CHR|1|3|Henoch, Ma thusala, Lamech,
1CHR|1|4|Noe, Sem, Cham et Iapheth.
1CHR|1|5|Filii Iapheth: Gomer, Magog, Madai et Iavan, Thubal, Mosoch, Thiras.
1CHR|1|6|Porro filii Gomer: Aschenez et Riphath et Thogorma.
1CHR|1|7|Filii autem Iavan: Elisa et Tharsis, Getthim et Rodanim.
1CHR|1|8|Filii Cham: Chus et Mesraim, Phut et Chanaan.
1CHR|1|9|Filii autem Chus: Saba et Hevila, Sabatha et Regma et Sabathacha. Porro filii Regma: Saba et Dedan.
1CHR|1|10|Chus autem genuit Nemrod; iste coepit esse potens in terra.
1CHR|1|11|Mesraim vero genuit Ludim et Anamim et Laabim et Nephthuim,
1CHR|1|12|Phetrusim quoque et Chasluim, de quibus egressi sunt Philisthim e Caphtorim.
1CHR|1|13|Chanaan vero genuit Sidonem primogenitum, Heth,
1CHR|1|14|Iebusaeum quoque et Amorraeum et Gergesaeum
1CHR|1|15|Hevaeumque et Aracaeum et Sinaeum,
1CHR|1|16|Aradium quoque et Samaraeum et Emathaeum.
1CHR|1|17|Filii Sem: Elam et Assur et Arphaxad et Lud et Aram. Filii autem Aram: Us et Hul et Gether et Mes.
1CHR|1|18|Arphaxad autem genuit Sala, qui et ipse genuit Heber.
1CHR|1|19|Porro Heber nati sunt duo filii: nomen uni Phaleg, quia in diebus eius divisa est terra, et nomen fratris eius Iectan.
1CHR|1|20|Iectan autem genuit Elmodad et Saleph et Asarmoth et Iare,
1CHR|1|21|Adoram quoque et Uzal et Decla,
1CHR|1|22|Ebal etiam et Abimael et Saba necnon
1CHR|1|23|et Ophir et Hevila et Iobab; omnes isti filii Iectan.
1CHR|1|24|Sem, Arphaxad, Sala,
1CHR|1|25|Heber, Phaleg, Reu,
1CHR|1|26|Seruch, Nachor, Thare,
1CHR|1|27|Abram: iste est Abraham.
1CHR|1|28|Filii autem Abraham: Isaac et Ismael.
1CHR|1|29|Et hae generationes eorum: primogenitus Ismaelis Nabaioth et Cedar et Adbeel et Mabsam,
1CHR|1|30|Masma et Duma, Massa, Hadad et Thema,
1CHR|1|31|Iethur, Naphis, Cedma; hi sunt filii Ismaelis.
1CHR|1|32|Filii autem Ceturae concubinae Abraham, quos genuit: Zamran, Iecsan, Madan, Madian, Iesboc, Sue. Porro filii Iecsan: Saba et Dedan. Filii autem Dedan: Assurim et Latusim et Loommim.
1CHR|1|33|Filii autem Madian: Epha et Opher et Henoch et Abida et Eldaa. Omnes hi filii Ceturae.
1CHR|1|34|Generavit autem Abraham Isaac, cuius fuerunt filii Esau et Israel.
1CHR|1|35|Filii Esau: Eliphaz, Rahuel, Iehus, Ialam, Core.
1CHR|1|36|Filii Eliphaz: Theman, Omar, Sepho, Gatham, Cenez, Thamna, Amalec.
1CHR|1|37|Filii Rahuel: Nahath, Zara, Samma, Meza.
1CHR|1|38|Filii Seir: Lotan, Sobal, Sebeon, Ana, Dison, Eser, Disan.
1CHR|1|39|Filii Lotan: Hori, Hemam; soror autem Lotan fuit Thamna.
1CHR|1|40|Filii Sobal: Alvan et Manahath et Ebal et Sepho et Onam. Filii Sebeon: Aia et Ana.
1CHR|1|41|Filii Ana: Dison. Filii Dison: Hemdan et Eseban et Iethran et Charran.
1CHR|1|42|Filii Eser: Bilhan et Zavan et Iacan. Filii Disan: Us et Aran.
1CHR|1|43|Isti sunt reges, qui imperaverunt in terra Edom, antequam esset rex super filios Israel: Bela filius Beor, et nomen civitatis eius Denaba.
1CHR|1|44|Mortuus est autem Bela, et regnavit pro eo Iobab filius Zarae de Bosra.
1CHR|1|45|Cumque et Iobab fuisset mortuus, regnavit pro eo Husam de terra Themanorum.
1CHR|1|46|Obiit quoque et Husam, et regnavit pro eo Adad filius Badad, qui percussit Madian in terra Moab; et nomen civitatis eius Avith.
1CHR|1|47|Cumque et Adad fuisset mortuus, regnavit pro eo Semla de Masreca.
1CHR|1|48|Sed et Semla mortuus est; et regnavit pro eo Saul de Rohoboth, quae iuxta amnem sita est.
1CHR|1|49|Mortuo quoque Saul, regnavit pro eo Baalhanan filius Achobor.
1CHR|1|50|Sed et hic mortuus est, et regnavit pro eo Adad, cuius urbis fuit nomen Phau; et appellata est uxor eius Meetabel filia Matred filiae Mezaab.
1CHR|1|51|Adad autem mortuo, duces pro regibus in Edom esse coeperunt: dux Thamna, dux Alva, dux Ietheth,
1CHR|1|52|dux Oolibama, dux Ela, dux Phinon,
1CHR|1|53|dux Cenez, dux Theman, dux Mabsar,
1CHR|1|54|dux Magdiel, dux Iram. Hi duces Edom.
1CHR|2|1|Filii autem Israel: Ruben, Simeon, Levi, Iuda, Issachar et Zabulon,
1CHR|2|2|Dan, Ioseph, Beniamin, Nephthali, Gad, Aser.
1CHR|2|3|Filii Iudae: Her, Onan et Sela; hi tres nati sunt ei de filia Sue Chananitide. Fuit autem Her primogenitus Iudae malus coram Domino, et occidit eum.
1CHR|2|4|Thamar autem nurus eius peperit ei Phares et Zara; omnes ergo filii Iudae quinque.
1CHR|2|5|Filii autem Phares: Esrom et Hamul.
1CHR|2|6|Filii quoque Zarae: Zamri et Ethan et Heman, Chalchol quoque et Darda; simul quinque.
1CHR|2|7|Filii Charmi: Achar, qui turbavit Israel et peccavit in furto anathematis.
1CHR|2|8|Filii Ethan: Azarias.
1CHR|2|9|Filii autem Esrom, qui nati sunt ei: Ierameel et Aram et Chaleb.
1CHR|2|10|Porro Aram genuit Aminadab, Aminadab autem genuit Naasson principem filiorum Iudae,
1CHR|2|11|Naasson quoque genuit Salmon, de quo ortus est Booz.
1CHR|2|12|Booz vero genuit Obed, qui et ipse genuit Isai.
1CHR|2|13|Isai autem genuit primogenitum Eliab, secundum Abinadab, tertium Samma,
1CHR|2|14|quartum Nathanael, quintum Raddai,
1CHR|2|15|sextum Asom, septimum David.
1CHR|2|16|Quorum sorores fuerunt: Sarvia et Abigail; filii Sarviae: Abisai, Ioab et Asael, tres.
1CHR|2|17|Abigail autem genuit Amasa, cuius pater fuit Iether Ismaelites.
1CHR|2|18|Chaleb vero filius Esrom genuit de uxore sua nomine Azuba, de qua nati sunt Ierioth, Ieser et Sobab et Ardon.
1CHR|2|19|Cumque mortua fuisset Azuba, accepit uxorem Chaleb Ephratha, quae peperit ei Hur.
1CHR|2|20|Porro Hur genuit Uri, et Uri genuit Beseleel.
1CHR|2|21|Post haec ingressus est Esrom ad filiam Machir patris Galaad et accepit eam, cum ipse esset annorum sexaginta; quae peperit ei Segub.
1CHR|2|22|Sed et Segub genuit Iair, qui possedit viginti tres civitates in terra Galaad.
1CHR|2|23|Cepitque Gesur et Aram oppida Iair ipsis et Canath et viculos eius sexaginta civitates. Omnes isti filii Machir patris Galaad.
1CHR|2|24|Cum autem mortuus esset Esrom, ingressus est Chaleb ad Ephratha uxorem Esrom patris sui. Habuit quoque Esrom uxorem Abia, quae peperit ei Ashur patrem Thecue.
1CHR|2|25|Nati sunt autem filii Ierameel primogeniti Esrom: Ram primogenitus eius et Buna et Aran et Asom et Ahia.
1CHR|2|26|Duxit quoque uxorem alteram Ierameel nomine Atara, quae fuit mater Onam.
1CHR|2|27|Sed et filii Ram primogeniti Ierameel fuerunt: Moos et Iamin et Acar.
1CHR|2|28|Onam autem habuit filios: Sammai et Iada. Filii autem Sammai: Nadab et Abisur.
1CHR|2|29|Nomen vero uxoris Abisur Abiail, quae peperit ei Ahobban et Molid.
1CHR|2|30|Filii autem Nadab fuerunt Saled et Apphaim; mortuus est autem Saled absque liberis.
1CHR|2|31|Filius vero Apphaim: Iesi, qui Iesi genuit Sesan; porro Sesan genuit Oholai.
1CHR|2|32|Filii autem Iada fratris Semmei: Iether et Ionathan; sed et Iether mortuus est absque liberis.
1CHR|2|33|Porro Ionathan genuit Phaleth et Ziza. Isti fuerunt filii Ierameel.
1CHR|2|34|Sesan autem non habuit filios sed filias et servum Aegyptium nomine Ieraa;
1CHR|2|35|deditque ei filiam suam uxorem, quae peperit ei Eththei.
1CHR|2|36|Eththei autem genuit Nathan, et Nathan genuit Zabad;
1CHR|2|37|Zabad quoque genuit Ophlal, et Ophlal genuit Obed.
1CHR|2|38|Obed genuit Iehu, Iehu genuit Azariam;
1CHR|2|39|Azarias genuit Helles, Helles genuit Elasa.
1CHR|2|40|Elasa genuit Sisamoi, Sisamoi genuit Sellum;
1CHR|2|41|Sellum genuit Iecemiam, Iecemias genuit Elisama.
1CHR|2|42|Filii autem Chaleb fratris Ierameel: Mesa primogenitus eius, ipse est pater Ziph; et filius eius Maresa pater Hebron.
1CHR|2|43|Porro filii Hebron: Core et Thapphua et Recem et Samma;
1CHR|2|44|Samma autem genuit Raham patrem Iercaam, et Recem genuit Sammai.
1CHR|2|45|Filius Sammai: Maon, et Maon pater Bethsur.
1CHR|2|46|Epha autem concubina Chaleb peperit Charran et Mosa et Gezez; porro Charran genuit Gezez.
1CHR|2|47|Filii Iahaddai: Regem et Iotham et Gesan et Phalet et Epha et Saaph.
1CHR|2|48|Concubina Chaleb Maacha peperit Saber et Tharana.
1CHR|2|49|Genuit autem Saaph pater Madmena Sue patrem Machbena et patrem Gabaa. Filia vero Chaleb fuit Achsa.
1CHR|2|50|Hi erant filii Chaleb.Filii Hur primogeniti Ephratha: Sobal pater Cariathiarim,
1CHR|2|51|Salmon pater Bethlehem, Hariph pater Bethgader.
1CHR|2|52|Fuerunt autem filii Sobal patris Cariathiarim Raaia, dimidium Manahat
1CHR|2|53|et cognationes Cariathiarim: Iethraei et Phutaei et Sumathaei et Maseraei. Ex his egressi sunt Saraitae et Esthaolitae.
1CHR|2|54|Filii Salmon: Bethlehem et Netophathitae, Atarothbethioab et dimidium Manahat de Saraa,
1CHR|2|55|cognationes quoque de Cariathsepher habitantes in Iabes: Therathaei, Semathaei et Suchathaei. Hi sunt Cinaei, qui orti sunt de Ammath patre domus Rechab.
1CHR|3|1|David vero hos habuit filios, qui ei nati sunt in Hebron: primoge nitum Amnon ex Achinoam Iezrahelitide, secundum Daniel de Abigail de Carmel,
1CHR|3|2|tertium Absalom filium Maacha filiae Tholmai regis Gesur, quartum Adoniam filium Haggith,
1CHR|3|3|quintum Saphatiam ex Abital, sextum Iethraam de Egla uxore sua.
1CHR|3|4|Sex ergo nati sunt ei in Hebron, ubi regnavit septem annis et sex mensibus. Triginta autem et tribus annis regnavit in Ierusalem.
1CHR|3|5|Porro in Ierusalem nati sunt ei filii: Samua et Sobab et Nathan et Salomon, quattuor de Bethsabee filia Ammiel;
1CHR|3|6|Iebahar quoque et Elisama et Eliphalet
1CHR|3|7|et Noga et Napheg et Iaphia
1CHR|3|8|necnon Elisama et Eliada et Eliphalet, novem.
1CHR|3|9|Omnes hi filii David absque filiis concubinarum; habueruntque sororem Thamar.
1CHR|3|10|Filius autem Salomonis Roboam, cuius Abia filius genuit Asa; de hoc quoque natus est Iosaphat
1CHR|3|11|pater Ioram; qui Ioram genuit Ochoziam, ex quo ortus est Ioas.
1CHR|3|12|Et huius Amasias filius genuit Azariam, porro Azariae filius Ioatham
1CHR|3|13|procreavit Achaz patrem Ezechiae, de quo natus est Manasses.
1CHR|3|14|Sed et Manasses genuit Amon patrem Iosiae;
1CHR|3|15|filii autem Iosiae fuerunt: primogenitus Iohanan, secundus Ioachim, tertius Sedecias, quartus Sellum.
1CHR|3|16|Filii Ioachim: Iechonias filius eius, Sedecias filius eius.
1CHR|3|17|Filii Iechoniae captivi fuerunt: Salathiel filius eius,
1CHR|3|18|Melchiram, Phadaia, Senasser et Iecemias, Hosama et Nadabias.
1CHR|3|19|De Phadaia orti sunt Zorobabel et Semei. Zorobabel genuit Mosollam, Hananiam et Salomith sororem eorum
1CHR|3|20|Hasabamque et Ohol et Barachiam et Hasadiam, Iosabhesed, quinque.
1CHR|3|21|Filii autem Hananiae: Pheltias, Iesaias, Raphaia, Arnan, Abdia et Sechenias.
1CHR|3|22|Filii Secheniae: Semeia et Hattus et Igal et Baria et Naaria et Saphat, sex numero.
1CHR|3|23|Filii Naariae: Elioenai et Ezechias et Ezricam, tres.
1CHR|3|24|Filii Elioenai: Odovia et Eliasib et Pheleia et Accub et Iohanan et Dalaia et Anani, septem.
1CHR|4|1|Filii Iudae: Phares, Esrom et Charmi et Hur et Sobal.
1CHR|4|2|Reaia vero filius Sobal genuit Iahath, de quo nati sunt Ahumai et Laad; hae cognationes Saraitarum.
1CHR|4|3|Et ista stirps Etam: Iezrahel et Iesema et Iedebos, nomenque sororis eorum Asalelphuni.
1CHR|4|4|Phanuel autem pater Gedor et Ezer pater Hosa; isti sunt filii Hur primogeniti Ephratha patris Bethlehem.
1CHR|4|5|Ashur vero patris Thecue erant duae uxores: Halaa et Naara.
1CHR|4|6|Peperit autem ei Naara Oozam et Hepher et Themani et Ahasthari; isti sunt filii Naara.
1CHR|4|7|Porro filii Halaa: Sereth et Sohar et Ethnan.
1CHR|4|8|Cos autem genuit Anob et Sobeba et cognationes Aharehel filii Arum.
1CHR|4|9|Fuit autem Iabes inclitus prae fratribus suis; et mater eius vocavit nomen illius Iabes dicens: " Quia peperi eum in dolore ".
1CHR|4|10|Invocavit vero Iabes Deum Israel dicens: " Si benedicens benedixeris mihi et dilataveris terminos meos, et fuerit manus tua mecum, et feceris me a malitia non opprimi! ". Et praestitit Deus quae precatus est.
1CHR|4|11|Chelub autem frater Suaa genuit Mahir, qui fuit pater Esthon.
1CHR|4|12|Porro Esthon genuit Bethrapha et Phasea et Tehinna patrem Hirnaas (id est urbis Naas); hi sunt viri Recha.
1CHR|4|13|Filii autem Cenez: Othoniel et Saraia; porro filii Othoniel: Hathath et Maonathi.
1CHR|4|14|Maonathi genuit Ophra, Saraia autem genuit Ioab patrem Geharasim (id est vallis Artificum); ibi quippe artifices erant.
1CHR|4|15|Filii vero Chaleb filii Iephonne: Hir et Ela et Naham; filius quoque Ela: Cenez.
1CHR|4|16|Filii quoque Iallelel: Ziph et Zipha, Thiria et Asarel.
1CHR|4|17|Et filii Ezra: Iether et Mered et Epher et Ialon. Et genuit Iether Mariam et Sammai et Iesba patrem Esthemo.
1CHR|4|18|Hi autem sunt filii Bethiae filiae pharaonis, quam accepit Mered.
1CHR|4|19|Filii autem uxoris eius Iudaicae sororis Naham patris Ceilae: Dalaia et Simeon pater Ioman. Filii autem Naham patris Ceilae: Garmitae et Esthemo Maachathitarum.
1CHR|4|20|Filii quoque Simon: Ammon et Rinna, Benhanan et Thilon. Et filii Iesi: Zoheth et Benzoheth.
1CHR|4|21|Filii Sela filii Iudae: Her pater Lecha et Laada pater Maresa et cognationes domus operantium byssum in Bethasbea
1CHR|4|22|et Iochim virique Chozeba et Ioas et Saraph, qui principes fuerunt in Moab et qui reversi sunt in Bethlehem; hae autem sunt res veteres.
1CHR|4|23|Hi sunt figuli habitantes Netaim et Gedera; apud regem in operibus eius commorati sunt ibi.
1CHR|4|24|Filii Simeon: Namuel et Iamin, Iarib, Zara, Saul;
1CHR|4|25|Sellum filius eius, Mabsam filius eius, Masma filius eius.
1CHR|4|26|Filii Masma: Hamuel filius eius, Zacchur filius eius, Semei filius eius.
1CHR|4|27|Filii Semei sedecim et filiae sex; fratres autem eius non habuerunt filios multos, et universa cognatio eorum non potuit adaequare summam filiorum Iudae.
1CHR|4|28|Habitaverunt autem in Bersabee et Molada et Asarsual
1CHR|4|29|et in Bilha et in Esem et in Tholad
1CHR|4|30|et in Bathuel et in Horma et in Siceleg
1CHR|4|31|et in Bethmarchaboth et in Asarsusim et in Bethberai et in Saarim; hae civitates eorum usque ad regem David.
1CHR|4|32|Villae quoque eorum: Etam et Ain, Remmon et Thochen et Asan, civitates quinque.
1CHR|4|33|Et universi viculi eorum per circuitum civitatum istarum usque ad Baal; haec est habitatio eorum et genealogia.
1CHR|4|34|Masobab quoque et Iemlech et Iosa filius Amasiae
1CHR|4|35|et Ioel et Iehu filius Iosabiae filii Saraiae filii Asiel
1CHR|4|36|et Elioenai et Iacoba et Isuhaia et Asaia et Adiel et Isimiel et Banaia,
1CHR|4|37|Ziza quoque filius Sephei filii Allon filii Iedaia filii Semri filii Samaia.
1CHR|4|38|Isti nominatim inscripti erant principes in cognationibus suis; et familiae eorum expansae sunt vehementer,
1CHR|4|39|et profecti sunt ad introitum Gedor usque ad orientem vallis, ut quaererent pascua gregibus suis.
1CHR|4|40|Inveneruntque pascuas uberes et valde bonas et terram latissimam et quietam et fertilem, in qua ante habitaverunt de stirpe Cham.
1CHR|4|41|Hi ergo venerunt, qui inscripti erant nominatim, in diebus Ezechiae regis Iudae, et percusserunt tabernacula eorum et Meunitas, qui inventi fuerunt ibi, et deleverunt eos usque in praesentem diem habitaveruntque pro eis, quoniam uberrimas ibidem pascuas reppererunt.
1CHR|4|42|De filiis quoque Simeon abierunt in montem Seir viri quingenti habentes principes Pheltiam et Naariam et Raphaiam et Oziel filios Iesi
1CHR|4|43|et percusserunt reliquias, quae evadere potuerant Amalecitarum, et habitaverunt ibi pro eis usque ad diem hanc.
1CHR|5|1|Filii quoque Ruben primogeniti Israel: ipse quippe fuit primoge nitus eius, sed, cum violasset torum patris sui, data sunt primogenita eius filiis Ioseph filii Israel, ut non computaretur in primogenitum,
1CHR|5|2|quia Iuda erat quidem fortissimus inter fratres suos et de stirpe eius principes germinati sunt, primogenita autem reputata sunt Ioseph.
1CHR|5|3|Filii ergo Ruben primogeniti Israel: Henoch et Phallu, Hesron et Charmi.
1CHR|5|4|Filii Ioel: Semeia filius eius, Gog filius eius, Semei filius eius,
1CHR|5|5|Micha filius eius, Reaia filius eius, Baal filius eius,
1CHR|5|6|Beera filius eius, quem captivum duxit Theglathphalasar rex Assyriorum, et fuit princeps in tribu Ruben.
1CHR|5|7|Fratres autem eius in cognationibus eius, quando numerabantur in genealogiis suis, erant: caput Iehiel, deinde Zacharias;
1CHR|5|8|porro Bela filius Azaz filii Samma filii Ioel, ipse habitavit in Aroer usque ad Nabo et Baalmeon.
1CHR|5|9|Contra orientalem quoque plagam habitavit usque ad introitum eremi, quae est inde a flumine Euphrate; multum quippe gregum eorum numerus creverat in terra Galaad.
1CHR|5|10|In diebus autem Saul proeliati sunt contra Agarenos et interfecerunt illos; habitaveruntque pro eis in tabernaculis eorum in omni plaga, quae respicit ad orientem Galaad.
1CHR|5|11|Filii vero Gad e regione eorum habitaverunt in terra Basan usque Salcha:
1CHR|5|12|Ioel in capite et Sapham secundus, porro Ianai et Saphat in Basan;
1CHR|5|13|fratres vero eorum secundum familias suas: Michael et Mosollam et Seba et Iorai et Iachan et Zie et Heber, septem.
1CHR|5|14|Hi filii Abihail filii Huri filii Iaroe filii Galaad filii Michael filii Iesesi filii Ieddo filii Buz.
1CHR|5|15|Ahi filius Abdiel filii Guni princeps familiarum eorum.
1CHR|5|16|Et habitaverunt in Galaad et in Basan et in viculis eius et in cunctis suburbanis Saron usque ad terminos.
1CHR|5|17|Omnes hi numerati sunt in diebus Ioatham regis Iudae et in diebus Ieroboam regis Israel.
1CHR|5|18|Filii Ruben et Gad et dimidiae tribus Manasse viri bellatores scuta portantes et gladios et tendentes arcum eruditique ad proelia, quadraginta quattuor milia et septingenti sexaginta procedentes ad pugnam;
1CHR|5|19|dimicaverunt contra Agarenos et Ituraeos et Naphisaeos et Nodabaeos.
1CHR|5|20|Et datum est eis auxilium, traditique sunt in manus eorum Agareni et universi, qui fuerant cum eis, quia Deum invocaverunt cum proeliarentur, et exaudivit eos, eo quod credidissent in eum.
1CHR|5|21|Ceperuntque omnia, quae possederant, camelorum quinquaginta milia et ovium ducenta quinquaginta milia, asinos duo milia et animas hominum centum milia;
1CHR|5|22|vulnerati autem multi corruerunt; fuit enim bellum Domini. Habitaveruntque pro eis usque ad transmigrationem.
1CHR|5|23|Filii quoque dimidiae tribus Manasse possederunt terram a Basan usque Baalhermon et Sanir et montem Hermon; ingens quippe numerus erat.
1CHR|5|24|Et hi fuerunt principes familiarum eorum: Epher et Iesi et Eliel et Azriel et Ieremia et Odovia et Iediel; viri bellatores fortissimi et nominati, duces in familiis suis.
1CHR|5|25|Reliquerunt autem Deum patrum suorum et fornicati sunt post deos populorum terrae, quos abstulit Deus coram eis.
1CHR|5|26|Et suscitavit Deus Israel spiritum Phul regis Assyriorum et spiritum Theglathphalasar regis Assur; et transtulit Ruben et Gad et dimidium tribus Manasse et adduxit eos in Hala et Habor et Ara et fluvium Gozan usque ad diem hanc.
1CHR|5|27|Filii Levi: Gerson, Caath, Merari.
1CHR|5|28|Filii Caath: Amram, Isaar, Hebron et Oziel.
1CHR|5|29|Filii Amram: Aaron, Moyses et Maria. Filii Aaron: Nadab et Abiu, Eleazar et Ithamar.
1CHR|5|30|Eleazar genuit Phinees, et Phinees genuit Abisue;
1CHR|5|31|Abisue vero genuit Bocci, et Bocci genuit Ozi.
1CHR|5|32|Ozi genuit Zaraiam, et Zaraias genuit Meraioth,
1CHR|5|33|porro Meraioth genuit Amariam, et Amarias genuit Achitob;
1CHR|5|34|Achitob genuit Sadoc, Sadoc genuit Achimaas,
1CHR|5|35|Achimaas genuit Azariam, Azarias genuit Iohanan;
1CHR|5|36|Iohanan genuit Azariam: ipse est qui sacerdotio functus est in domo, quam aedificavit Salomon in Ierusalem.
1CHR|5|37|Genuit autem Azarias Amariam, et Amarias genuit Achitob,
1CHR|5|38|Achitob genuit Sadoc, et Sadoc genuit Sellum;
1CHR|5|39|Sellum genuit Helciam, et Helcias genuit Azariam.
1CHR|5|40|Azarias genuit Saraiam, et Saraias genuit Iosedec;
1CHR|5|41|porro Iosedec egressus est, quando transtulit Dominus Iudam et Ierusalem per manus Nabuchodonosor.
1CHR|6|1|Filii ergo Levi: Gerson, Caath et Merari.
1CHR|6|2|Et haec nomina filio rum Gerson: Lobni et Semei.
1CHR|6|3|Filii Caath: Amram et Isaar et Hebron et Oziel.
1CHR|6|4|Filii Merari: Moholi et Musi.Hae autem cognationes Levi secundum familias eorum:
1CHR|6|5|Gerson, Lobni filius eius, Iahath filius eius, Zimma filius eius,
1CHR|6|6|Ioah filius eius, Addo filius eius, Zara filius eius, Iethrai filius eius.
1CHR|6|7|Filii Caath: Aminadab filius eius, Core filius eius, Asir filius eius,
1CHR|6|8|Elcana filius eius, Abiasaph filius eius, Asir filius eius,
1CHR|6|9|Thahath filius eius, Uriel filius eius, Ozias filius eius, Saul filius eius.
1CHR|6|10|Filii Elcana: Amasai et Achimoth,
1CHR|6|11|Elcana filius eius, Sophai filius eius, Nahath filius eius,
1CHR|6|12|Eliab filius eius, Ieroham filius eius, Elcana filius eius, Samuel filius eius.
1CHR|6|13|Filii Samuel: primogenitus Ioel et secundus Abia.
1CHR|6|14|Filii autem Merari: Moholi, Lobni filius eius, Semei filius eius, Oza filius eius,
1CHR|6|15|Samaa filius eius, Haggia filius eius, Asaia filius eius.
1CHR|6|16|Isti sunt, quos constituit David super cantum domus Domini, ex quo collocata est arca;
1CHR|6|17|et ministrabant coram habitatione tabernaculi conventus canentes, donec aedificaret Salomon domum Domini in Ierusalem; stabant autem iuxta ordinem suum in ministerio.
1CHR|6|18|Hi vero sunt, qui assistebant cum filiis suis. De filiis Caath: Heman cantor filius Ioel filii Samuel
1CHR|6|19|filii Elcana filii Ieroham filii Eliel filii Thohu
1CHR|6|20|filii Suph filii Elcana filii Mahath filii Amasai
1CHR|6|21|filii Elcana filii Ioel filii Azariae filii Sophoniae
1CHR|6|22|filii Thahath filii Asir filii Abiasaph filii Core
1CHR|6|23|filii Isaar filii Caath filii Levi filii Israel.
1CHR|6|24|Et frater eius Asaph, qui stabat a dextris eius, Asaph filius Barachiae filii Samaa
1CHR|6|25|filii Michael filii Basaiae filii Melchiae
1CHR|6|26|filii Athnai filii Zara filii Adaia
1CHR|6|27|filii Ethan filii Zimma filii Semei
1CHR|6|28|filii Iahath filii Gerson filii Levi.
1CHR|6|29|Filii autem Merari fratres eorum ad sinistram: Ethan filius Cusi filii Abdi filii Melluch
1CHR|6|30|filii Hasabiae filii Amasiae filii Helciae
1CHR|6|31|filii Amsi filii Bani filii Somer
1CHR|6|32|filii Moholi filii Musi filii Merari filii Levi.
1CHR|6|33|Fratres quoque eorum Levitae, qui ordinati sunt in cunctum ministerium habitaculi domus Domini;
1CHR|6|34|Aaron vero et filii eius adolebant super altare holocausti et super altare thymiamatis in omne opus sancti sanctorum, et ut expiarent pro Israel, iuxta omnia quae praecepit Moyses servus Dei.
1CHR|6|35|Hi sunt autem filii Aaron: Eleazar filius eius, Phinees filius eius, Abisue filius eius,
1CHR|6|36|Bocci filius eius, Ozi filius eius, Zaraia filius eius,
1CHR|6|37|Meraioth filius eius, Amarias filius eius, Achitob filius eius,
1CHR|6|38|Sadoc filius eius, Achimaas filius eius.
1CHR|6|39|Et haec habitacula eorum per castra atque confinia, filiorum scilicet Aaron ex cognatione Caathitarum; ipsis enim sorte contigerat.
1CHR|6|40|Dederunt igitur eis Hebron in terra Iudae et suburbana eius per circuitum;
1CHR|6|41|agros autem civitatis et villas Chaleb filio Iephonne.
1CHR|6|42|Porro filiis Aaron dederunt civitatem ad confugiendum: Hebron et Lobna et suburbana eius,
1CHR|6|43|Iether quoque et Esthemo cum suburbanis eius, sed et Helon et Dabir cum suburbanis suis,
1CHR|6|44|Asan quoque et Iutta et Bethsames et suburbana earum;
1CHR|6|45|de tribu autem Beniamin: Gabaon et Gabaa et suburbana earum et Almath cum suburbanis suis, Anathoth quoque cum suburbanis suis: omnes civitates tredecim, singulae per cognationes suas.
1CHR|6|46|Filiis autem Caath residuis de cognatione sua dederunt ex tribu Ephraim et ex tribu Dan et ex dimidia tribu Manasse in possessionem urbes decem.
1CHR|6|47|Porro filiis Gerson per cognationes suas de tribu Issachar et de tribu Aser et de tribu Nephthali et de tribu Manasse in Basan urbes tredecim.
1CHR|6|48|Filiis autem Merari per cognationes suas de tribu Ruben et de tribu Gad et de tribu Zabulon dederunt sorte civitates duodecim.
1CHR|6|49|Dederunt quoque filii Israel Levitis civitates et suburbana earum;
1CHR|6|50|dederuntque per sortem ex tribu filiorum Iudae et ex tribu filiorum Simeon et ex tribu filiorum Beniamin urbes has, quas vocaverunt nominibus suis.
1CHR|6|51|Et his, qui erant ex cognationibus filiorum Caath, fuerunt civitates in terminis eorum de tribu Ephraim.
1CHR|6|52|Dederunt ergo eis urbem ad confugiendum: Sichem cum suburbanis suis in monte Ephraim et Gazer cum suburbanis suis,
1CHR|6|53|Iecmaam quoque cum suburbanis suis et Bethoron similiter;
1CHR|6|54|necnon et Aialon cum suburbanis suis et Gethremmon in eundem modum.
1CHR|6|55|Porro ex dimidia tribu Manasse Thanach et suburbana eius, Ieblaam et suburbana eius, his videlicet qui de cognationibus filiorum Caath reliqui erant.
1CHR|6|56|Filiis autem Gerson de cognationibus dimidiae tribus Manasse: Golan in Basan et suburbana eius et Astharoth cum suburbanis suis.
1CHR|6|57|De tribu Issachar Cedes et suburbana illius et Dabereth cum suburbanis suis,
1CHR|6|58|Ramoth quoque et suburbana illius et Anem cum suburbanis suis.
1CHR|6|59|De tribu vero Aser: Masal cum suburbanis suis et Abdon similiter,
1CHR|6|60|Hucoc quoque et suburbana eius et Rohob cum suburbanis suis.
1CHR|6|61|Porro de tribu Nephthali: Cedes in Galilaea et suburbana eius, Hamon cum suburbanis suis et Cariathaim et suburbana eius.
1CHR|6|62|Filiis autem Merari residuis de tribu Zabulon: Remmon et suburbana eius et Thabor cum suburbanis suis.
1CHR|6|63|Trans Iordanem quoque ex adverso Iericho, contra orientem Iordanis de tribu Ruben: Bosor in solitudine cum suburbanis suis et Iasa cum suburbanis suis,
1CHR|6|64|Cademoth quoque et suburbana eius et Mephaath cum suburbanis suis.
1CHR|6|65|Necnon et de tribu Gad: Ramoth in Galaad et suburbana eius et Mahanaim cum suburbanis suis,
1CHR|6|66|sed et Hesebon cum suburbanis eius, et Iazer cum suburbanis suis.
1CHR|7|1|Porro filii Issachar: Thola et Phua, Iasub et Semron, quat tuor.
1CHR|7|2|Filii Thola: Ozi et Raphaia et Ieriel et Iemai et Iebsem et Samuel, principes familiarum suarum; de stirpe Thola viri fortissimi numerati sunt iuxta genealogias suas in diebus David viginti duo milia sescenti.
1CHR|7|3|Filii Ozi: Izrahia, de quo nati sunt Michael et Obadia et Ioel et Iesia, quinque principes omnes.
1CHR|7|4|Cumque eis erant secundum genealogias familiarum suarum turmae accinctae ad proelium, viri fortissimi, triginta sex milia; multas enim habuere uxores et filios.
1CHR|7|5|Fratresque eorum per omnes cognationes Issachar robustissimi ad pugnandum octoginta septem milia numerati sunt.
1CHR|7|6|Filii Beniamin: Bela et Bochor et Iedihel, tres.
1CHR|7|7|Filii Bela: Esebon et Ozi et Oziel et Ierimoth et Urai, quinque principes familiarum et ad pugnandum robustissimi; numerus autem eorum viginti duo milia et triginta quattuor.
1CHR|7|8|Porro filii Bochor: Zamira et Ioas et Eliezer et Elioenai et Amri et Ierimoth et Abia et Anathoth et Almath; omnes hi filii Bochor.
1CHR|7|9|Numerati sunt autem in genealogiis suis principes familiarum suarum ad bella fortissimi viginti milia et ducenti.
1CHR|7|10|Porro filii Iedihel: Bilhan; filii autem Bilhan: Iehus et Beniamin et Aod et Chanaana et Zethan et Tharsis et Ahisahar;
1CHR|7|11|omnes hi filii Iedihel principes familiarum suarum viri fortissimi decem et septem milia et ducenti ad proelium procedentes.
1CHR|7|12|Suphim quoque et Huphim filii Hir et Husim filii Aher.
1CHR|7|13|Filii autem Nephthali: Iasiel et Guni et Ieser et Sellum, filii Bilhae.
1CHR|7|14|Porro filius Manasse: Asriel, quem peperit concubina eius Syra; peperit quoque Machir patrem Galaad.
1CHR|7|15|Machir autem accepit uxorem de Huphim et Suphim et habuit sororem nomine Maacha; nomen autem secundi Salphaad, nataeque sunt Salphaad filiae.
1CHR|7|16|Et peperit Maacha uxor Machir filium vocavitque nomen eius Phares; porro nomen fratris eius Sares et filii eius Ulam et Recem.
1CHR|7|17|Filius autem Ulam: Badan; hi sunt filii Galaad filii Machir filii Manasse.
1CHR|7|18|Soror autem eius Ammalecheth peperit Isod et Abiezer et Maala.
1CHR|7|19|Erant autem filii Semida: Ahin et Sechem et Leci et Aniam.
1CHR|7|20|Filii autem Ephraim: Suthala, Bared filius eius, Thahath filius eius, Elada filius eius, Thahath filius eius,
1CHR|7|21|et huius filius Zabad et huius filius Suthala et huius filius Ezer et Elad. Occiderunt autem eos viri Geth indigenae, quia descenderant, ut invaderent possessiones eorum.
1CHR|7|22|Luxit igitur Ephraim pater eorum multis diebus, et venerunt fratres eius, ut consolarentur eum;
1CHR|7|23|ingressusque est ad uxorem suam, quae concepit et peperit filium, et vocavit nomen eius Beria, eo quod in malis domus eius ortus esset.
1CHR|7|24|Filia autem eius fuit Sara, quae aedificavit Bethoron inferiorem et superiorem et Ozensara.
1CHR|7|25|Porro filius eius Rapha et Reseph et Thale filius eius, de quo natus est Thaan,
1CHR|7|26|qui genuit Laadan; huius quoque filius Ammiud genuit Elisama,
1CHR|7|27|de quo ortus est Nun, qui habuit filium Iosue.
1CHR|7|28|Possessio autem eorum et habitationes: Bethel cum filiabus suis et contra orientem Noran, ad occidentalem plagam Gazer et filiae eius, Sichem quoque cum filiabus suis usque Hai et filias eius.
1CHR|7|29|Iuxta filios quoque Manasse: Bethsan et filias eius, Thanach et filias eius, Mageddo et filias eius, Dor et filias eius. In his habitaverunt filii Ioseph filii Israel.
1CHR|7|30|Filii Aser: Iemna et Iesua et Isui et Beria et Sara soror eorum.
1CHR|7|31|Filii autem Beria: Heber et Melchiel, ipse est pater Barzaith.
1CHR|7|32|Heber autem genuit Iephlat et Somer et Hotham et Suaa sororem eorum.
1CHR|7|33|Filii Iephlat: Phosech et Bamaal et Asoth; hi filii Iephlat.
1CHR|7|34|Porro filii Somer fratris sui: Roaga et Haba et Aram.
1CHR|7|35|Filii autem Hotham fratris eius: Supha et Iemna et Selles et Amal.
1CHR|7|36|Filii Supha: Sue, Hamapher et Sual et Beri et Iamra,
1CHR|7|37|Bosor et Od et Samma et Salusa et Iethran et Beera.
1CHR|7|38|Filii Iether: Iephonne et Phaspha et Ara.
1CHR|7|39|Filii autem Olla: Area et Hanniel et Resia.
1CHR|7|40|Omnes hi filii Aser, principes familiarum electi atque fortissimi, capita principum; numerus autem eorum, qui inscripti erant in exercitu ad bellum, viginti sex milia.
1CHR|8|1|Beniamin autem genuit Bela primogenitum suum, Asbel se cundum, Ahara tertium,
1CHR|8|2|Nohaa quartum et Rapha quintum.
1CHR|8|3|Fueruntque filii Bela: Addar et Gera pater Aod,
1CHR|8|4|Abisue quoque et Naaman et Ahoe,
1CHR|8|5|sed et Gera et Sephuphan et Huram.
1CHR|8|6|Hi sunt filii Aod principes familiarum habitantium in Gabaa, qui translati sunt in Manahath;
1CHR|8|7|Naaman autem et Ahia et Gera: ipse transtulit eos et genuit Oza et Ahiud.
1CHR|8|8|Porro Saharaim genuit in regione Moab, postquam dimisit Husim et Bara uxores suas;
1CHR|8|9|genuit autem de Hodes uxore sua Iobab et Sebia et Mesa et Melcham,
1CHR|8|10|Iehus quoque et Sechia et Marma; hi sunt filii eius principes in familiis suis.
1CHR|8|11|De Husim vero genuit Abitob et Elphaal;
1CHR|8|12|porro filii Elphaal Heber et Misaam et Samad; hic aedificavit Ono et Lod et filias eius.
1CHR|8|13|Beria autem et Samma principes familiarum habitantium in Aialon; hi fugaverunt habitatores Geth.
1CHR|8|14|Et Ahi et Sesac et Ierimoth
1CHR|8|15|et Zabadia et Arad et Eder,
1CHR|8|16|Michael quoque et Iespha et Ioha filii Beria.
1CHR|8|17|Et Zabadia et Mosollam et Hezeci et Heber
1CHR|8|18|et Iesamari et Iezlia et Iobab filii Elphaal
1CHR|8|19|et Iacim et Zechri et Zabdi
1CHR|8|20|et Elioenai et Selethai et Eliel
1CHR|8|21|et Adaia et Baraia et Samarath filii Semei
1CHR|8|22|et Iesphan et Heber et Eliel
1CHR|8|23|et Abdon et Zechri et Hanan
1CHR|8|24|et Hanania et Elam et Anathothia
1CHR|8|25|et Iephdaia et Phanuel filii Sesac.
1CHR|8|26|Et Samsari et Sohoria et Otholia
1CHR|8|27|et Iersia et Elia et Zechri filii Ieroham.
1CHR|8|28|Hi capita familiarum secundum genealogias, principes qui habitaverunt in Ierusalem.
1CHR|8|29|In Gabaon autem habitaverunt Iehiel pater Gabaon, et nomen uxoris eius Maacha,
1CHR|8|30|filiusque eius primogenitus Abdon et Sur et Cis et Baal et Ner et Nadab,
1CHR|8|31|Gedor quoque et Ahio et Zacher et Macelloth;
1CHR|8|32|et Macelloth genuit Samaa. Habitaveruntque ex adverso fratrum suorum in Ierusalem cum fratribus suis.
1CHR|8|33|Ner autem genuit Cis, et Cis genuit Saul. Porro Saul genuit Ionathan et Melchisua et Abinadab et Isbaal.
1CHR|8|34|Filius autem Ionathan Meribbaal, et Meribbaal genuit Micha;
1CHR|8|35|filii Micha Phithon et Melech et Tharaa et Ahaz.
1CHR|8|36|Et Ahaz genuit Ioada, et Ioada genuit Almath et Azmaveth et Zamri; porro Zamri genuit Mosa.
1CHR|8|37|Et Mosa genuit Banaa, cuius filius fuit Raphaia, de quo ortus est Elasa, qui genuit Asel.
1CHR|8|38|Porro Asel sex filii fuere his nominibus: Ezricam primogenitus eius, Ismael, Saria, Azarias, Obdia et Hanan; omnes hi filii Asel.
1CHR|8|39|Filii autem Esec fratris eius: Ulam primogenitus et Iehus secundus et Eliphalet tertius.
1CHR|8|40|Fueruntque filii Ulam viri robustissimi ad bellum et magno robore tendentes arcum et multos habentes filios ac nepotes usque ad centum quinquaginta. Omnes hi filii Beniamin.
1CHR|9|1|Universus ergo Israel dinume ratus est, et summa eorum scrip ta est in libro regum Israel et Iudae. Translatique sunt in Babylonem propter delictum suum.
1CHR|9|2|Qui autem habitaverunt primi in possessionibus et in urbibus suis: Israel et sacerdotes et Levitae et Nathinaei.
1CHR|9|3|Commorati sunt in Ierusalem de filiis Iudae et de filiis Beniamin, de filiis quoque Ephraim et Manasse.
1CHR|9|4|Uthai filius Ammiud filii Amri filii Imri filii Bani: de filiis Phares filii Iudae;
1CHR|9|5|et de Selanitis: Asaia primogenitus et filii eius;
1CHR|9|6|de filiis autem Zara: Iehuel et fratres eorum sescenti nonaginta.
1CHR|9|7|Porro de filiis Beniamin: Sallu filius Mosollam filii Odovia filii Asana
1CHR|9|8|et Iobania filius Ieroham et Ela filius Ozi filii Mochori et Mosollam filius Saphatiae filii Rahuel filii Iebaniae
1CHR|9|9|et fratres eorum secundum genealogias suas nongenti quinquaginta sex; omnes hi principes familiarum secundum familias suas.
1CHR|9|10|De sacerdotibus autem: Iedaia, Ioiarib et Iachin,
1CHR|9|11|Azarias quoque filius Helciae filii Mosollam filii Sadoc filii Meraioth filii Achitob principes domus Dei.
1CHR|9|12|Porro Adaias filius Ieroham filii Phassur filii Melchiae et Maasai filius Adiel filii Iezra filii Mosollam filii Mosollamoth filii Emmer,
1CHR|9|13|fratres quoque eorum principes per familias suas mille septingenti sexaginta, fortissimi robore ad faciendum opus ministerii in domo Dei.
1CHR|9|14|De Levitis autem: Semeia filius Hassub filii Ezricam filii Hasabia de filiis Merari;
1CHR|9|15|Bacbacar quoque, Hares et Galal et Matthania filius Micha filii Zechri filii Asaph
1CHR|9|16|et Abdia filius Semeiae filii Galal filii Idithun et Barachia filius Asa filii Elcana, qui habitavit in atriis Netophathitarum.
1CHR|9|17|Ianitores autem: Sellum et Accub et Telmon et Ahiman; et frater eorum Sellum princeps
1CHR|9|18|et usque ad hoc tempus est in porta regis ad orientem. Hi erant ianitores castris filiorum Levi.
1CHR|9|19|Sellum vero filius Core filii Abiasaph filii Core cum fratribus suis de domo patris sui: hi Coritae erant super opera ministerii custodes liminum tabernaculi; patres autem eorum super castra Domini custodiebant introitum,
1CHR|9|20|et Phinees filius Eleazari princeps erat super eos olim - Dominus sit cum eo! -
1CHR|9|21|Zacharias filius Mosollamia ianitor portae tabernaculi conventus.
1CHR|9|22|Omnes hi electi in ostiarios liminum ducenti duodecim, et descripti in villis propriis, quos constituerunt David et Samuel videns in munus perpetuum,
1CHR|9|23|tam ipsos quam filios eorum in ostiis domus Domini, domus tabernaculi, in custodias.
1CHR|9|24|Per quattuor ventos erant ostiarii, id est ad orientem et ad occidentem, ad aquilonem et ad austrum.
1CHR|9|25|Fratres autem eorum in viculis suis morabantur et veniebant per septem dies de tempore usque ad tempus, ut essent cum illis.
1CHR|9|26|Nam munus habebant perpetuum hi quattuor principes ianitorum. Hi scilicet Levitae erant super exedras et thesauros domus Domini;
1CHR|9|27|per gyrum quoque templi Domini pernoctabant in custodiis suis, ut et ipsi mane aperirent fores.
1CHR|9|28|De horum genere erant et super vasa ministerii, ad numerum enim et inferebantur vasa et efferebantur;
1CHR|9|29|de ipsis et, qui credita habebant utensilia et omnia utensilia sancta, praeerant similae et vino et oleo et turi et aromatibus.
1CHR|9|30|Filii quidam autem sacerdotum unguenta ex aromatibus conficiebant;
1CHR|9|31|et Matthathias Levites, primogenitus Sellum Coritae, munere perpetuo praefectus erat eorum, quae in sartagine frigebantur.
1CHR|9|32|Porro de filiis Caath fratribus eorum super panes erant propositionis, ut semper novos per singula sabbata praepararent.
1CHR|9|33|Hi sunt cantores, principes per familias Levitarum, qui in exedris vacantes morabantur, ita ut die et nocte iugiter suo ministerio deservirent.
1CHR|9|34|Hi sunt capita Levitarum per familias suas secundum genealogias suas principes; hi habitaverunt in Ierusalem.
1CHR|9|35|In Gabaon autem commorati sunt pater Gabaon Iehiel, et nomen uxoris eius Maacha.
1CHR|9|36|Filius primogenitus eius Abdon et Sur et Cis et Baal et Ner et Nadab,
1CHR|9|37|Gedor quoque et Ahio et Zacharias et Macelloth.
1CHR|9|38|Porro Macelloth genuit Samaam; isti habitaverunt e regione fratrum suorum in Ierusalem cum fratribus suis.
1CHR|9|39|Ner autem genuit Cis, et Cis genuit Saul. Et Saul genuit Ionathan et Melchisua et Abinadab et Isbaal.
1CHR|9|40|Filius autem Ionathan Meribbaal, et Meribbaal genuit Micha;
1CHR|9|41|porro filii Micha: Phithon et Melech et Tharaa et Ahaz.
1CHR|9|42|Ahaz autem genuit Iara, et Iara genuit Almath et Azmaveth et Zamri; Zamri autem genuit Mosa.
1CHR|9|43|Mosa vero genuit Banaa, cuius filius Raphaia genuit Elasa, de quo ortus est Asel.
1CHR|9|44|Porro Asel sex filios habuit his nominibus: Ezricam primogenitus eius, Ismael, Saria, Azarias, Obdia, Hanan; hi filii Asel.
1CHR|10|1|Philisthim autem pugnabant contra Israel, fugeruntque viri Israel a facie Philisthim et ceciderunt vulnerati in monte Gelboe;
1CHR|10|2|cumque appropinquassent Philisthaei persequentes Saul et filios eius, percusserunt Ionathan et Abinadab et Melchisua filios Saul.
1CHR|10|3|Et aggravatum est proelium contra Saul, inveneruntque eum sagittarii et vulneraverunt iaculis;
1CHR|10|4|et dixit Saul ad armigerum suum: " Evagina gladium tuum et interfice me, ne forte veniant incircumcisi isti et illudant mihi ". Noluit autem armiger eius hoc facere timore perterritus. Arripuit igitur Saul ensem et irruit in eum;
1CHR|10|5|quod cum vidisset armiger eius, videlicet mortuum esse Saul, irruit etiam ipse in gladium suum et mortuus est.
1CHR|10|6|Interiit ergo Saul et tres filii eius; omnis domus illius pariter concidit.
1CHR|10|7|Quod cum vidissent omnes viri Israel, qui habitabant in campestribus, quod fugissent, et mortui essent Saul et filii eius, dereliquerunt urbes suas et huc illucque dispersi sunt; veneruntque Philisthim et habitaverunt in eis.
1CHR|10|8|Die igitur altero venerunt Philisthim, ut spoliarent interfectos, et invenerunt Saul et filios eius iacentes in monte Gelboe;
1CHR|10|9|cumque spoliassent eum et amputassent caput armisque nudassent, miserunt in terram suam per circuitum, ut annuntiaretur in idolorum templis et in populis.
1CHR|10|10|Arma autem eius consecraverunt in fano Astharoth et caput affixerunt in templo Dagon.
1CHR|10|11|Hoc cum audissent viri Iabes Galaad, omnia scilicet quae Philisthim fecerunt super Saul,
1CHR|10|12|consurrexerunt omnes viri fortes et tulerunt cadavera Saul et filiorum eius attuleruntque ea in Iabes et sepelierunt ossa eorum subter quercum, quae erat in Iabes, et ieiunaverunt septem diebus.
1CHR|10|13|Mortuus est ergo Saul propter iniquitatem suam, eo quod praevaricatus sit mandatum Domini, quod praeceperat, et non custodierit illud, sed insuper etiam pythonissam consuluerit
1CHR|10|14|nec quaesierit Dominum; propter quod et interfecit eum et transtulit regnum eius ad David filium Isai.
1CHR|11|1|Congregatus est igitur omnis Israel ad David in Hebron dicens: " Os tuum sumus et caro tua.
1CHR|11|2|Heri quoque et nudiustertius, cum adhuc regnaret Saul, tu eras qui educebas et introducebas Israel; tibi enim dixit Dominus Deus tuus: "Tu pasces populum meum Israel et tu eris princeps super eum" ".
1CHR|11|3|Venerunt ergo omnes maiores natu Israel ad regem in Hebron, et iniit David cum eis foedus in Hebron coram Domino; unxeruntque eum regem super Israel iuxta sermonem Domini, quem locutus est in manu Samuel.
1CHR|11|4|Abiit quoque David et omnis Israel in Ierusalem, haec est Iebus, ubi erant Iebusaei habitatores terrae.
1CHR|11|5|Dixeruntque, qui habitabant in Iebus, ad David: " Non ingredieris huc ". Porro David cepit arcem Sion, quae est civitas David;
1CHR|11|6|dixitque: " Omnis, qui percusserit Iebusaeum, in primis erit princeps et dux ". Ascendit igitur primus Ioab filius Sarviae et factus est princeps.
1CHR|11|7|Habitavit autem David in arce, et idcirco appellata est civitas David.
1CHR|11|8|Aedificavitque urbem in circuitu a Mello usque ad gyrum; Ioab autem reliqua urbis instauravit.
1CHR|11|9|Proficiebatque David vadens et crescens, et Dominus exercituum erat cum eo.
1CHR|11|10|Hi principes virorum fortium David, qui adiuverunt eum, ut rex fieret super omnem Israel iuxta verbum Domini, quod locutus est ad Israel;
1CHR|11|11|et iste numerus robustorum David: Iesbaam filius Hachamon filius Hachamonitis princeps inter triginta; iste levavit hastam suam super trecentos, quos occidit impetu uno.
1CHR|11|12|Et post eum Eleazar filius Dodo Ahohites, qui erat inter tres potentes;
1CHR|11|13|iste fuit cum David in Aphesdommim, quando Philisthim congregati sunt ad locum illum in proelium. Et erat ager regionis illius plenus hordeo, fugeratque populus a facie Philisthinorum.
1CHR|11|14|Hic stetit in medio agri et defendit eum; cumque percussisset Philisthaeos, dedit Dominus salutem magnam populo suo.
1CHR|11|15|Descenderunt autem tres de triginta principibus ad petram, in qua erat David, ad speluncam Odollam, quando Philisthim fuerant castrametati in valle Raphaim.
1CHR|11|16|Porro David erat in praesidio, et statio Philisthinorum in Bethlehem;
1CHR|11|17|desideravit igitur David et dixit: " O si quis daret mihi aquam de cisterna Bethlehem, quae est in porta! ".
1CHR|11|18|Tres ergo isti per media castra Philisthinorum perrexerunt et hauserunt aquam de cisterna Bethlehem, quae erat in porta, et attulerunt ad David, ut biberet. Qui noluit, sed magis libavit illam Domino
1CHR|11|19|dicens: " Avertat a me Deus meus, ut hoc faciam et sanguinem virorum istorum bibam, quia in periculo animarum suarum attulerunt mihi aquam ". Et ob hanc causam noluit bibere. Haec fecerunt tres robustissimi.
1CHR|11|20|Abisai quoque frater Ioab; ipse erat princeps inter triginta et ipse levavit hastam suam contra trecentos, quos interfecit, et ipse erat inter tres nominatus,
1CHR|11|21|inter triginta duplici honore eminens et princeps eorum; verumtamen usque ad tres non pervenerat.
1CHR|11|22|Banaias filius Ioiadae vir robustissimus, qui multa opera perpetrarat, de Cabseel; ipse percussit duos Ariel de Moab et ipse descendit et interfecit leonem in media cisterna tempore nivis.
1CHR|11|23|Et ipse percussit virum Aegyptium, cuius statura erat quinque cubitorum, et habebat lanceam ut liciatorium texentium; descendit ergo ad eum cum virga et rapuit hastam, quam tenebat manu, et interfecit eum hasta sua.
1CHR|11|24|Haec fecit Banaias filius Ioiadae, qui erat inter tres robustos nominatus,
1CHR|11|25|inter triginta primus; verumtamen ad tres usque non pervenerat, posuit autem eum David super satellites suos.
1CHR|11|26|Porro fortissimi in exercitu: Asael frater Ioab et Elchanan filius Dodo de Bethlehem,
1CHR|11|27|Sammoth Harodites, Elica Harodites, Heles Phalonites,
1CHR|11|28|Hira filius Acces Thecuites, Abiezer Anathothites,
1CHR|11|29|Sobbochai Husathites, Ilai Ahohites,
1CHR|11|30|Maharai Netophathites, Heled filius Baana Netophathites,
1CHR|11|31|Ithai filius Ribai de Gabaa filiorum Beniamin, Banaia Pharathonites,
1CHR|11|32|Hurai de tor rentibus Gaas, Abiel Arbathites,
1CHR|11|33|Azmaveth Bahurimites, Eliaba Saalbonites,
1CHR|11|34|Asem Gezonites, Ionathan filius Sage Ararites,
1CHR|11|35|Ahiam filius Sachar Ararites, Eliphal filius Ur,
1CHR|11|36|Hepher Mecherathites, Ahia Phelonites,
1CHR|11|37|Hesro de Carmel, Naarai filius Azbai,
1CHR|11|38|Ioel frater Nathan, Mibahar filius Agarai,
1CHR|11|39|Selec Ammonites, Naharai Berothites armiger Ioab filii Sarviae,
1CHR|11|40|Hira Iethraeus, Gareb Iethraeus,
1CHR|11|41|Urias Hetthaeus, Zabad filius Oholai,
1CHR|11|42|Adina filius Siza Rubenites princeps Rubenitarum, et cum eo triginta;
1CHR|11|43|Hanan filius Maacha et Iosaphat Matthanites,
1CHR|11|44|Ozia Astharothites, Sama et Iehiel filii Hotham Aroerites,
1CHR|11|45|Iedihel filius Semri et Ioha frater eius Thosaites,
1CHR|11|46|Eliel Mahumites et Ieribai et Iosaia filii Elnaem et Iethma Moabites,
1CHR|11|47|Eliel et Obed et Iasiel de Soba.
1CHR|12|1|Hi quoque venerunt ad Da vid in Siceleg, cum adhuc fu geret Saul filium Cis; qui erant fortissimi et egregii pugnatores
1CHR|12|2|tendentes arcum et utraque manu fundis saxa iacientes et dirigentes sagittas. De fratribus Saul ex Beniamin:
1CHR|12|3|princeps Ahiezer et Ioas filii Samaa Gabaathites et Iaziel et Phalet filii Azmaveth et Baracha et Iehu Anathothites;
1CHR|12|4|Iesmaias quoque Gabaonites fortissimus inter triginta et super triginta,
1CHR|12|5|Ieremias et Iahaziel et Iohanan et Iozabad Gederothites,
1CHR|12|6|Eluzai et Ierimoth et Baalia et Samaria et Saphatia Haruphites,
1CHR|12|7|Elcana et Iesia et Azareel et Ioezer et Iesbaam Coritae,
1CHR|12|8|Ioela quoque et Zabadia filii Ieroham de Gedor.
1CHR|12|9|Sed et de Gad transfugerunt ad David, cum lateret in deserto, viri robustissimi et pugnatores optimi tenentes clipeum et hastam; facies eorum quasi facies leonis et veloces quasi capreae in montibus:
1CHR|12|10|Ezer princeps, Abdias secundus, Eliab tertius,
1CHR|12|11|Masmana quartus, Ieremias quintus,
1CHR|12|12|Etthei sextus, Eliel septimus,
1CHR|12|13|Iohanan octavus, Elzebad nonus,
1CHR|12|14|Ieremias decimus, Machbanai undecimus.
1CHR|12|15|Hi de filiis Gad principes exercitus, minimus contra centum praevalebat et maximus contra mille.
1CHR|12|16|Isti sunt qui transierunt Iordanem mense primo, quando inundare consuevit super ripas suas, et omnes fugaverunt, qui morabantur in vallibus ad orientalem plagam et occidentalem.
1CHR|12|17|Venerunt autem et de Beniamin et de Iuda ad praesidium, in quo morabatur David.
1CHR|12|18|Egressusque est David obviam eis et ait: " Si pacifice venistis ad me, ut auxiliemini mihi, cor meum iungatur vobis; si autem insidiamini mihi pro adversariis meis, cum ego iniquitatem in manibus non habeam, videat Deus patrum nostrorum et iudicet ".
1CHR|12|19|Spiritus vero induit Amasai principem inter triginta, et ait: Tui sumus, o David,et tecum, fili Isai!Pax, pax tibiet pax adiutoribus tuis;te enim adiuvat Deus tuus ".Suscepit ergo eos David et constituit principes turmae.
1CHR|12|20|Porro de Manasse transfugerunt ad David, quando veniebat cum Philisthim adversus Saul, ut pugnaret; et non dimicavit cum eis, quia inito consilio remiserunt eum principes Philisthinorum dicentes: " Periculo capitis nostri revertetur ad dominum suum Saul ".
1CHR|12|21|Quando igitur reversus est in Siceleg, transfugerunt ad eum de Manasse Ednas et Iozabad et Iedihel et Michael et Iozabad et Eliu et Selathai principes milium in Manasse:
1CHR|12|22|hi praebuerunt auxilium David adversus latrunculos; omnes enim erant viri fortissimi et facti sunt principes in exercitu.
1CHR|12|23|Sed et per singulos dies veniebant ad David ad auxiliandum ei, usque dum fieret grandis numerus quasi exercitus Dei.
1CHR|12|24|Iste quoque est numerus principum exercitus, qui venerunt ad David, cum esset in Hebron, ut transferrent regnum Saul ad eum iuxta verbum Domini.
1CHR|12|25|Filii Iudae portantes clipeum et hastam sex milia octingenti expediti ad proelium.
1CHR|12|26|De filiis Simeon virorum fortissimorum ad pugnandum septem milia centum.
1CHR|12|27|De filiis Levi quattuor milia sescenti;
1CHR|12|28|Ioiada quoque princeps de stirpe Aaron et cum eo tria milia septingenti;
1CHR|12|29|Sadoc etiam iuvenis fortissimus et familia eius principes viginti duo.
1CHR|12|30|De filiis autem Beniamin fratribus Saul tria milia; magna enim pars eorum adhuc sequebatur domum Saul.
1CHR|12|31|Porro de filiis Ephraim viginti milia octingenti, fortissimi robore viri nominati in familiis suis.
1CHR|12|32|Et ex dimidia parte tribus Manasse decem et octo milia; singuli per nomina sua destinati, ut venirent et constituerent regem David.
1CHR|12|33|De filiis quoque Issachar viri eruditi, qui norant singula tempora ad sciendum quid facere deberet Israel, principes ducenti et omnes fratres eorum ad iussa eorum.
1CHR|12|34|Porro de Zabulon, qui egrediebantur ad proelium et stabant in acie instructi omnibus armis bellicis, quinquaginta milia venerunt, ut congregarentur non in corde duplici.
1CHR|12|35|Et de Nephthali principes mille; et cum eis instructa clipeo et hasta triginta septem milia.
1CHR|12|36|De Dan etiam praeparata ad proelium viginti octo milia sescenti.
1CHR|12|37|Et de Aser egredientes ad pugnam et in acie procedentes quadraginta milia.
1CHR|12|38|Trans Iordanem autem de filiis Ruben et de Gad et dimidia parte tribus Manasse, instructi omnibus armis bellicis, centum viginti milia.
1CHR|12|39|Omnes isti viri bellatores expediti ad pugnandum corde perfecto venerunt in Hebron, ut constituerent regem David super universum Israel; sed et omnes reliqui ex Israel uno corde erant, ut rex fieret David.
1CHR|12|40|Fueruntque ibi apud David tribus diebus comedentes et bibentes; praeparaverunt enim eis fratres sui.
1CHR|12|41|Sed et qui iuxta eos erant, usque ad Issachar et Zabulon et Nephthali, afferebant panes in asinis et camelis et mulis et bobus, escam farinae, palathas, uvam passam, vinum, oleum, boves, oves ad omnem copiam; gaudium quippe erat in Israel.
1CHR|13|1|Iniit autem consilium David cum tribunis et centurionibus et universis principibus
1CHR|13|2|et ait ad omnem coetum Israel: " Si placet vobis, et a Domino Deo nostro egreditur sermo, quem loquor, mittamus ad fratres nostros reliquos in universas regiones Israel et ad sacerdotes et Levitas, qui habitant in suburbanis urbium, ut congregentur ad nos,
1CHR|13|3|et reducamus arcam Dei nostri ad nos; non enim requisivimus eam in diebus Saul ".
1CHR|13|4|Et respondit universa multitudo, ut ita fieret; placuerat enim sermo omni populo.
1CHR|13|5|Congregavit ergo David cunctum Israel a Sihor Aegypti usque ad introitum dum ingrediaris Emath, ut adduceret arcam Dei de Cariathiarim.
1CHR|13|6|Et ascendit David et omnis Israel in Baala, in Cariathiarim, quae est in Iuda, ut afferrent inde arcam Dei Domini sedentis super cherubim, ubi invocatum est nomen eius.
1CHR|13|7|Imposueruntque arcam Dei super plaustrum novum de domo Abinadab. Oza autem et Ahio minabant plaustrum.
1CHR|13|8|Porro David et universus Israel ludebant coram Deo omni virtute in canticis et in citharis et psalteriis et tympanis et cymbalis et tubis.
1CHR|13|9|Cum autem pervenissent ad aream Chidon, tetendit Oza manum suam, ut sustentaret arcam; boves quippe lascivientes proruperunt.
1CHR|13|10|Iratus est itaque Dominus contra Ozam et percussit eum, eo quod contigisset arcam; et mortuus est ibi coram Deo.
1CHR|13|11|Contristatusque est David, eo quod dirupisset Dominus Ozam; et vocatus est locus ille Pharesoza (id est Diruptio Ozae) usque in praesentem diem.
1CHR|13|12|Et timuit Deum tunc temporis dicens: " Quomodo possum ad me introducere arcam Dei? ".
1CHR|13|13|Et ob hanc causam non eam adduxit ad se, hoc est in civitatem David, sed avertit in domum Obededom Getthaei.
1CHR|13|14|Mansit ergo arca Dei apud domum Obededom tribus mensibus; et benedixit Dominus domui eius et omnibus quae habebat.
1CHR|14|1|Misit quoque Hiram rex Tyri nuntios ad David et ligna cedrina et artifices parietum lignorumque, ut aedificarent ei domum.
1CHR|14|2|Cognovitque David quod confirmasset eum Dominus in regem super Israel et sublevatum esset regnum suum propter populum eius Israel.
1CHR|14|3|Accepit quoque David alias uxores in Ierusalem genuitque filios et filias;
1CHR|14|4|et haec nomina eorum, qui nati sunt ei in Ierusalem: Samua et Sobab, Nathan et Salomon,
1CHR|14|5|Iebahar et Elisua et Eliphalet,
1CHR|14|6|Noga quoque et Napheg et Iaphia,
1CHR|14|7|Elisama et Beeliada et Eliphalet.
1CHR|14|8|Audientes autem Philisthim quod unctus esset David in regem super universum Israel, ascenderunt omnes, ut quaererent eum; quod cum audisset David, egressus est obviam eis.
1CHR|14|9|Porro Philisthim venientes diffusi sunt in valle Raphaim.
1CHR|14|10|Consuluitque David Deum dicens: " Si ascendam contra Philisthaeos, et si trades eos in manu mea? ". Et dixit ei Dominus: " Ascende, et tradam eos in manu tua ".
1CHR|14|11|Cumque illi ascendissent in Baalpharasim, percussit eos ibi David et dixit: " Dirupit Deus inimicos meos per manum meam sicut dirumpuntur aquae. Et idcirco vocatum est nomen loci illius Baalpharasim (id est Dominus diruptionum).
1CHR|14|12|Dereliqueruntque ibi deos suos, quos David iussit exuri.
1CHR|14|13|Alia etiam vice Philisthim irruerunt et diffusi sunt in valle;
1CHR|14|14|consuluitque rursum David Deum, et dixit ei Deus: " Non ascendas post eos; circumdabis eos et venies contra illos ex adverso arborum celthium;
1CHR|14|15|cumque audieris sonitum gradientis in cacumine arborum celthium, tunc egredieris ad bellum; egressus est enim Deus ante te, ut percutias castra Philisthim ".
1CHR|14|16|Fecit ergo David, sicut praeceperat ei Deus, et percussit castra Philisthinorum de Gabaon usque Gazer.
1CHR|14|17|Divulgatumque est nomen David in universis regionibus, et Dominus dedit pavorem eius super omnes gentes.
1CHR|15|1|Fecit quoque sibi domos in civitate David et praeparavit locum arcae Dei tetenditque ei tabernaculum.
1CHR|15|2|Tunc dixit David: " Illicitum est, ut a quocumque portetur arca Dei, nisi a Levitis, quos elegit Dominus ad portandum eam et ad ministrandum sibi usque in aeternum ".
1CHR|15|3|Congregavitque David universum Israel in Ierusalem, ut afferretur arca Domini in locum suum, quem praeparaverat ei;
1CHR|15|4|necnon et filios Aaron et Levitas.
1CHR|15|5|De filiis Caath Uriel princeps fuit et fratres eius centum viginti;
1CHR|15|6|de filiis Merari Asaia princeps et fratres eius ducenti viginti;
1CHR|15|7|de filiis Gerson Ioel princeps et fratres eius centum triginta;
1CHR|15|8|de filiis Elisaphan Semeias princeps et fratres eius ducenti;
1CHR|15|9|de filiis Hebron Eliel princeps et fratres eius octoginta;
1CHR|15|10|de filiis Oziel Aminadab princeps et fratres eius centum duodecim.
1CHR|15|11|Vocavitque David Sadoc et Abiathar sacerdotes et Levitas Uriel, Asaiam, Ioel, Semeiam, Eliel et Aminadab
1CHR|15|12|et dixit ad eos: " Vos, qui estis principes familiarum Leviticarum, sanctificamini cum fratribus vestris et afferte arcam Domini, Dei Israel, ad locum, quem praeparavi.
1CHR|15|13|Quia a principio non eratis praesentes, fecit Dominus, Deus Israel, diruptionem in nobis; non enim quaesivimus eum, sicut fas erat ".
1CHR|15|14|Sanctificati sunt ergo sacerdotes et Levitae, ut portarent arcam Domini, Dei Israel;
1CHR|15|15|et tulerunt filii Levi arcam Dei, sicut praeceperat Moyses iuxta verbum Domini, umeris suis in vectibus.
1CHR|15|16|Dixitque David principibus Levitarum, ut constituerent de fratribus suis cantores in organis musicorum, nablis videlicet et lyris et cymbalis, ut resonaret fortiter sonitus laetitiae.
1CHR|15|17|Constitueruntque Levitae Heman filium Ioel et de fratribus eius Asaph filium Barachiae, de filiis vero Merari fratribus eorum Ethan filium Casaiae
1CHR|15|18|et cum eis fratres eorum in secundo ordine Zachariam et Bani et Iaziel et Semiramoth et Iahiel et Ani, Eliab et Banaiam et Maasiam et Matthathiam et Eliphalu et Maceniam et Obededom et Iehiel ianitores.
1CHR|15|19|Porro cantores Heman, Asaph et Ethan in cymbalis aeneis bene sonantibus,
1CHR|15|20|Zacharias autem et Oziel et Semiramoth et Iahiel et Ani et Eliab et Maasias et Banaias in nablis secundum " Virgines ".
1CHR|15|21|Porro Matthathias et Eliphalu et Macenias et Obededom et Iehiel et Ozaziu in citharis super octavam, ut dirigerent;
1CHR|15|22|Chonenias autem princeps Levitarum portantium arcam praeerat ad portandum, erat quippe valde sapiens.
1CHR|15|23|Et Barachias et Elcana ianitores pro arca.
1CHR|15|24|Porro Sebania et Iosaphat et Nathanael et Amasai et Zacharias et Banaias et Eliezer sacerdotes clangebant tubis coram arca Dei, et Obededom et Iehias erant ianitores pro arca.
1CHR|15|25|Igitur David et maiores natu Israel et tribuni ierunt ad deportandam arcam foederis Domini de domo Obededom cum laetitia.
1CHR|15|26|Cumque adiuvisset Deus Levitas, qui portabant arcam foederis Domini, immolati sunt septem tauri et septem arietes.
1CHR|15|27|Porro David indutus pallio byssino et universi Levitae, qui portabant arcam, cantoresque et Chonenias princeps pro portanda arca - David autem indutus erat etiam ephod lineo -
1CHR|15|28|universusque Israel deducebant arcam foederis Domini in iubilo et sonitu bucinae et tubis et cymbalis bene sonantibus et nablis et citharis.
1CHR|15|29|Cumque pervenisset arca foederis Domini usque ad civitatem David, Michol filia Saul prospiciens per fenestram vidit regem David saltantem atque ludentem et despexit eum in corde suo.
1CHR|16|1|Attulerunt igitur arcam Dei et constituerunt eam in me dio tabernaculi, quod tetenderat ei David, et obtulerunt holocausta et pacifica coram Deo.
1CHR|16|2|Cumque complesset David offerens holocausta et pacifica, benedixit populo in nomine Domini.
1CHR|16|3|Et divisit unicuique de Israel a viro usque ad mulierem tortam panis et laganum palmarum et palatham.
1CHR|16|4|Constituitque coram arca Domini de Levitis ministros, qui recordarentur operum eius et glorificarent atque laudarent Dominum, Deum Israel:
1CHR|16|5|Asaph principem et secundum eius Zachariam, porro Iehiel et Semiramoth et Iahiel et Matthathiam et Eliab et Banaiam et Obededom et Iehiel in organis psalterii et citharis, Asaph autem, ut cymbalis personaret,
1CHR|16|6|Banaiam vero et Iahaziel sacerdotes, ut canerent tubis iugiter coram arca foederis Dei.
1CHR|16|7|In illo die, tunc fecit David prima vice confiteri Domino per manum Asaph et fratrum eius:
1CHR|16|8|" Confitemini Domino, invocate nomen eius,notas facite in populis opera eius.
1CHR|16|9|Canite ei et psalliteet narrate omnia mirabilia eius.
1CHR|16|10|Laudate nomen sanctum eius,laetetur cor quaerentium Dominum.
1CHR|16|11|Quaerite Dominum et virtutem eius,quaerite faciem eius semper.
1CHR|16|12|Recordamini mirabilium eius, quae fecit,signorum illius et iudiciorum oris eius,
1CHR|16|13|semen Israel, servi eius,filii Iacob, electi illius.
1CHR|16|14|Ipse Dominus Deus noster;in universa terra iudicia eius.
1CHR|16|15|Recordamini in sempiternum pacti eius,sermonis, quem praecepit in mille generationes,
1CHR|16|16|pacti, quod pepigit cum Abraham,et iuramenti illius cum Isaac.
1CHR|16|17|Et constituit illud Iacob in praeceptumet Israel in pactum sempiternum
1CHR|16|18|dicens: "Tibi dabo terram Chanaanfuniculum hereditatis vestrae",
1CHR|16|19|cum essent pauci numero,parvi et coloni in ea.
1CHR|16|20|Et transierunt de gente in gentemet de regno ad populum alterum;
1CHR|16|21|non dimisit quemquam calumniari eos,sed increpuit pro eis reges:
1CHR|16|22|"Nolite tangere christos meoset in prophetis meis nolite malignari".
1CHR|16|23|Canite Domino, omnis terra,annuntiate ex die in diem salutare eius.
1CHR|16|24|Narrate in gentibus gloriam eius,in cunctis populis mirabilia illius.
1CHR|16|25|Quia magnus Dominus et laudabilis nimiset horribilis super omnes deos;
1CHR|16|26|omnes enim dii populorum inania,Dominus autem caelos fecit.
1CHR|16|27|Magnificentia et pulchritudo coram eo,fortitudo et gaudium in loco eius.
1CHR|16|28|Afferte Domino, familiae populorumafferte Domino gloriam et imperium;
1CHR|16|29|date Domino gloriam nominis eius,levate oblationem et venite in conspectu eiuset adorate Dominum in decore sancto.
1CHR|16|30|Commoveatur a facie illius omnis terra;ipse enim fundavit orbem immobilem.
1CHR|16|31|Laetentur caeli, et exsultet terra,et dicant in nationibus: "Dominus regnat!".
1CHR|16|32|Tonet mare et plenitudo eius,exsultent agri et omnia, quae in eis sunt.
1CHR|16|33|Tunc laudabunt ligna saltus coram Domino,quia venit iudicare terram.
1CHR|16|34|Confitemini Domino, quoniam bonus,quoniam in aeternum misericordia eius.
1CHR|16|35|Et dicite: "Salva nos, Deus salvator noster,et congrega nos et erue de gentibus, ut confiteamur nomini sancto tuoet exsultemus in carminibus tuis.
1CHR|16|36|Benedictus Dominus, Deus Israel,ab aeterno usque in aeternum" ".Et dixit omnis populus: " Amen! " et " Laus Domino! ".
1CHR|16|37|Dereliquit itaque ibi coram arca foederis Domini Asaph et fratres eius, ut ministrarent in conspectu arcae iugiter secundum ritum singulorum dierum.
1CHR|16|38|Porro Obededom et fratres eius sexaginta octo et Obededom filium Idithun et Hosa constituit ianitores.
1CHR|16|39|Sadoc autem sacerdotem et fratres illius sacerdotes coram habitaculo Domini in excelso, quod erat in Gabaon,
1CHR|16|40|ut offerrent holocausta Domino super altare holocautomatis iugiter, mane et vespere, iuxta omnia, quae scripta sunt in lege Domini, quam praecepit Israeli.
1CHR|16|41|Et cum eis Heman et Idithun et reliquos electos, qui nominatim memorati sunt ad confitendum Domino: " Quoniam in aeternum misericordia eius ".
1CHR|16|42|Et cum eis Heman et Idithun canentes tuba et quatientes cymbala bene sonantia et omnia musicorum organa ad canendum Deo; filios autem Idithun fecit esse portarios.
1CHR|16|43|Reversusque est omnis populus unusquisque in domum suam et David, ut benediceret etiam domui suae.
1CHR|17|1|Cum autem habitaret David in domo sua, dixit ad Nathan prophetam: " Ecce ego habito in domo cedrina, arca autem foederis Domini sub pellibus est ".
1CHR|17|2|Et ait Nathan ad David: " Omnia, quae in corde tuo sunt, fac; Deus enim tecum est ".
1CHR|17|3|Igitur nocte illa factus est sermo Dei ad Nathan dicens:
1CHR|17|4|" Vade et loquere David servo meo: Haec dicit Dominus: Non aedificabis tu mihi domum ad habitandum;
1CHR|17|5|neque enim mansi in domo ex eo tempore, quo eduxi Israel usque ad hanc diem, sed fui semper migrans de tabernaculo in tabernaculum et de habitatione in habitationem.
1CHR|17|6|Ubicumque ambulabam in omni Israel, numquid locutus sum uni iudicum Israel, quibus praeceperam, ut pascerent populum meum, et dixi: Quare non aedificastis mihi domum cedrinam?
1CHR|17|7|Nunc itaque, sic loqueris ad servum meum David: Haec dicit Dominus exercituum: Ego tuli te, cum in pascuis sequereris gregem, ut esses dux populi mei Israel;
1CHR|17|8|et fui tecum, quocumque perrexisti, et interfeci omnes inimicos tuos coram te fecique tibi nomen quasi unius magnorum, qui celebrantur in terra.
1CHR|17|9|Et dedi locum populo meo Israel et plantavi eum, ut habitaret in eo, et ultra non commovebitur, nec filii iniquitatis atterent eos sicut in principio
1CHR|17|10|et ex diebus, quibus dedi iudices populo meo Israel et humiliavi universos inimicos tuos. Annuntio ergo tibi quod aedificaturus sit domum tibi Dominus.
1CHR|17|11|Cumque impleveris dies tuos, ut vadas ad patres tuos, suscitabo semen tuum post te, quod erit de filiis tuis, et stabiliam regnum eius.
1CHR|17|12|Ipse aedificabit mihi domum, et firmabo solium eius usque in aeternum.
1CHR|17|13|Ego ero ei in patrem, et ipse erit mihi in filium; et misericordiam meam non auferam ab eo, sicut abstuli ab eo, qui ante te fuit.
1CHR|17|14|Et statuam eum in domo mea et in regno meo usque in sempiternum, et thronus eius erit firmissimus in perpetuum ".
1CHR|17|15|Iuxta omnia verba haec et iuxta universam visionem istam, sic locutus est Nathan ad David.
1CHR|17|16|Cumque venisset rex David et sedisset coram Domino, dixit: " Quis ego sum, Domine Deus, et quae domus mea, quia adduxisti me hucusque?
1CHR|17|17|Sed hoc parum visum est in conspectu tuo, Deus; ideoque locutus es super domum servi tui etiam in futurum et aspexisti me excelsum super ordinem hominum, Domine Deus.
1CHR|17|18|Quid ultra addere potest David, cum ita glorificaveris servum tuum et cognoveris eum?
1CHR|17|19|Domine, propter famulum tuum iuxta cor tuum fecisti omnem magnificentiam hanc; et nota esse voluisti universa magnalia.
1CHR|17|20|Domine, non est similis tui, et non est alius deus absque te secundum omnia, quae audivimus auribus nostris.
1CHR|17|21|Quis autem est alius ut populus tuus Israel, gens una in terra, ad quam perrexit Deus, ut liberaret sibi populum, ut faceres tibi nomen magnum et terribile eiciens nationes a facie populi tui, quem de Aegypto liberasti?
1CHR|17|22|Et posuisti populum tuum Israel tibi in populum usque in aeternum; et tu, Domine, factus es Deus eius.
1CHR|17|23|Nunc igitur, Domine, sermo, quem locutus es super famulum tuum et super domum eius, confirmetur in perpetuum; et fac, sicut locutus es.
1CHR|17|24|Permaneatque et magnificetur nomen tuum usque in sempiternum, et dicatur: "Dominus exercituum, Deus Israel, est Deus pro Israel, et domus David servi tui permanens coram te".
1CHR|17|25|Tu enim, Deus meus, revelasti auriculam servi tui, ut aedificares ei domum; et idcirco invenit servus tuus fiduciam, ut oret coram te.
1CHR|17|26|Nunc ergo, Domine, tu es Deus; et locutus es super servum tuum tanta beneficia
1CHR|17|27|et coepisti benedicere domui servi tui, ut sit semper coram te: te enim, Domine, benedicente, benedicta erit in perpetuum ".
1CHR|18|1|Factum est autem post haec, ut percuteret David Phili sthim et humiliaret eos et tolleret Geth et filias eius de manu Philisthim
1CHR|18|2|percuteretque Moab, et fierent Moabitae servi David offerentes ei tributum.
1CHR|18|3|Et percussit David etiam Adadezer regem Soba in regione ad Emath, quando perrexit, ut dilataret imperium suum usque ad flumen Euphraten.
1CHR|18|4|Cepit ergo David mille quadrigas eius et septem milia equites ac viginti milia virorum peditum; subnervavitque omnes equos curruum, exceptis centum quadrigis, quas reservavit sibi.
1CHR|18|5|Supervenit autem et Syrus Damascenus, ut auxilium praeberet Adadezer regi Soba; sed et huius percussit David viginti duo milia virorum
1CHR|18|6|et posuit praesidium in Syria Damasci, ut Syria quoque serviret sibi et offerret tributum. Adiuvitque eum Dominus in cunctis, ad quae perrexerat.
1CHR|18|7|Tulit quoque David arma aurea, quae habuerant servi Adadezer, et attulit ea in Ierusalem;
1CHR|18|8|necnon de Tebah et Chun urbibus Adadezer aeris plurimum, de quo fecit Salomon mare aeneum et columnas et vasa aenea.
1CHR|18|9|Quod cum audisset Thou rex Emath, percussisse videlicet David omnem exercitum Adadezer regis Soba,
1CHR|18|10|misit Adoram filium suum ad regem David, ut salutaret eum et congratularetur, eo quod pugnasset cum Adadezer et percussisset eum; adversarius quippe erat Thou Adadezer.
1CHR|18|11|Sed et omnia vasa aurea et argentea et aenea consecravit rex David Domino cum argento et auro, quod tulerat ex universis gentibus, tam de Idumaea et Moab et filiis Ammon, quam de Philisthim et Amalec.
1CHR|18|12|Abisai vero filius Sarviae percussit Edom in valle Salis decem et octo milia
1CHR|18|13|et constituit in Edom praesidium, ut serviret Idumaea David. Salvavitque Dominus David in cunctis, ad quae perrexerat.
1CHR|18|14|Regnavit ergo David super universum Israel et faciebat iudicium atque iustitiam cuncto populo suo.
1CHR|18|15|Porro Ioab filius Sarviae erat super exercitum, et Iosaphat filius Ahilud a commentariis.
1CHR|18|16|Sadoc autem filius Achitob et Achimelech filius Abiathar sacerdotes et Susa scriba.
1CHR|18|17|Banaias vero filius Ioiadae super legiones Cherethi et Phelethi; porro filii David primi ad manum regis.
1CHR|19|1|Accidit autem post haec, ut moreretur Naas rex filiorum Ammon, et regnaret filius eius pro eo.
1CHR|19|2|Dixitque David: " Faciam misericordiam cum Hanon filio Naas; praestitit enim pater eius mihi gratiam ". Misitque David nuntios ad consolandum eum super morte patris sui. Qui cum pervenissent in terram filiorum Ammon, ut consolarentur Hanon,
1CHR|19|3|dixerunt principes filiorum Ammon ad Hanon: " Tu forsitan putas quod David honoris causa in patrem tuum miserit, qui consolentur te; nec animadvertis quod, ut explorent et investigent et evertant terram tuam, venerint ad te servi eius ".
1CHR|19|4|Igitur Hanon pueros David tulit et rasit et praecidit tunicas eorum a natibus usque ad pedes et dimisit eos.
1CHR|19|5|Qui cum abissent et hoc mandassent David, misit in occursum eorum - grandem enim contumeliam sustinuerant - et praecepit, ut manerent in Iericho, donec cresceret barba eorum, et tunc reverterentur.
1CHR|19|6|Videntes autem filii Ammon quod odiosos se fecissent David, tam Hanon quam reliquus populus miserunt mille talenta argenti, ut conducerent sibi de Mesopotamia et de Syria Maacha et de Soba currus et equites;
1CHR|19|7|conduxeruntque sibi triginta duo milia curruum et regem Maacha cum populo eius. Qui cum venissent, castrametati sunt e regione Medaba; filii quoque Ammon congregati de urbibus suis venerunt ad bellum.
1CHR|19|8|Quod cum audisset David, misit Ioab et omnem exercitum virorum fortium.
1CHR|19|9|Egressique filii Ammon direxerunt aciem iuxta portam civitatis; reges autem, qui ad auxilium venerant, separatim in agro steterunt.
1CHR|19|10|Igitur Ioab intellegens bellum et ex adverso et post tergum contra se fieri elegit viros fortissimos de universo Israel et perrexit contra Syrum;
1CHR|19|11|reliquam autem partem populi dedit sub manu Abisai fratris sui, et perrexerunt contra filios Ammon.
1CHR|19|12|Dixitque: " Si vicerit me Syrus, auxilio eris mihi; si autem superaverint te filii Ammon, ero tibi in praesidium.
1CHR|19|13|Confortare et agamus viriliter pro populo nostro et pro urbibus Dei nostri; Dominus autem, quod in conspectu suo bonum est, faciet ".
1CHR|19|14|Appropinquavit ergo Ioab et populus, qui cum eo erat, contra Syrum ad proelium, et fugerunt a facie eorum.
1CHR|19|15|Porro filii Ammon videntes quod fugisset Syrus, ipsi quoque fugerunt Abisai fratrem eius et ingressi sunt civitatem. Reversusque est etiam Ioab in Ierusalem.
1CHR|19|16|Videns autem Syrus quod cecidisset coram Israel, misit nuntios et adduxit Syrum, qui erat trans fluvium; Sophach autem princeps militiae Adadezer erat dux eorum.
1CHR|19|17|Quod cum nuntiatum esset David, congregavit universum Israel et transivit Iordanem venitque ad eos et direxit ex adverso aciem et pugnavit cum eis.
1CHR|19|18|Fugit autem Syrus Israel, et interfecit David de Syris septem milia curruum et quadraginta milia peditum et Sophach exercitus principem.
1CHR|19|19|Videntes autem servi Adadezer se ab Israel esse superatos, fecerunt pacem cum David et servierunt ei; noluitque ultra Syria auxilium praebere filiis Ammon.
1CHR|20|1|Factum est autem post anni circulum, eo tempore, quo solent reges ad bella procedere, eduxit Ioab robur exercitus et vastavit terram filiorum Ammon; perrexitque et obsedit Rabba. Porro David manebat in Ierusalem, quando Ioab percussit Rabba et destruxit eam.
1CHR|20|2|Tulit autem David coronam Melchom de capite eius et invenit in ea auri pondo talentum et pretiosissimam gemmam, venitque super caput David; manubias quoque urbis plurimas tulit.
1CHR|20|3|Populum autem, qui erat in ea, eduxit et condemnavit ad operam lapicidinarum et ad secures et dolabras ferreas. Sic fecit David cunctis urbibus filiorum Ammon et reversus est cum omni populo suo in Ierusalem.
1CHR|20|4|Post haec initum est bellum in Gazer adversum Philisthaeos, in quo percussit Sobbochai Husathites Saphai de genere Raphaim, et humiliavit eos.
1CHR|20|5|Aliud quoque bellum gestum est adversus Philisthaeos, in quo percussit Elchanan filius Iair Lahmi fratrem Goliath Getthaeum, cuius hastae lignum erat quasi liciatorium texentium.
1CHR|20|6|Sed et aliud bellum accidit in Geth, in quo fuit homo longissimus senos habens digitos, id est simul viginti quattuor, qui et ipse de Rapha fuerat stirpe generatus;
1CHR|20|7|hic blasphemavit Israel, et percussit eum Ionathan filius Samma fratris David. Hi sunt filii Rapha in Geth, qui ceciderunt in manu David et servorum eius.
1CHR|21|1|Consurrexit autem Satan contra Israel et incitavit Da vid, ut numeraret Israel.
1CHR|21|2|Dixitque David ad Ioab et ad principes populi: " Ite et numerate Israel a Bersabee usque Dan et afferte mihi numerum, ut sciam ".
1CHR|21|3|Responditque Ioab: " Augeat Dominus populum suum centuplum quam sunt. Nonne, domine mi rex, omnes servi tui sunt? Quare hoc quaerit dominus meus, quod in peccatum reputetur Israeli? ".
1CHR|21|4|Sed sermo regis magis praevaluit; egressusque est Ioab et circuivit universum Israel et reversus est Ierusalem.
1CHR|21|5|Deditque David numerum census, et inventus est omnis Israel numerus mille milia et centum milia virorum educentium gladium; de Iuda autem quadringenta septuaginta milia bellatorum;
1CHR|21|6|nam Levi et Beniamin non numeravit in medio eorum, eo quod invitus exequeretur regis imperium.
1CHR|21|7|Displicuit autem Deo, quod iussum erat, et percussit Israel.
1CHR|21|8|Dixitque David ad Deum: " Peccavi nimis, ut hoc facerem; obsecro, aufer iniquitatem servi tui, quia valde insipienter egi ".
1CHR|21|9|Et locutus est Dominus ad Gad videntem David dicens:
1CHR|21|10|" Vade et loquere ad David et dic: Haec dicit Dominus: Trium tibi optionem do: unum, quod volueris, elige, et faciam tibi ".
1CHR|21|11|Cumque venisset Gad ad David, dixit ei: " Haec dicit Dominus: Elige, quod volueris:
1CHR|21|12|aut tribus annis famem aut tribus mensibus fugere te hostes tuos et gladium eorum non posse evadere aut tribus diebus gladium Domini et pestilentiam versari in terra et angelum Domini interficere in universis finibus Israel. Nunc igitur vide quid respondeam ei, qui misit me ".
1CHR|21|13|Et dixit David ad Gad: " Ex omni parte me angustiae premunt, sed melius mihi est, ut incidam in manus Domini, quia multae sunt miserationes eius, quam in manus hominum ".
1CHR|21|14|Misit ergo Dominus pestilentiam in Israel, et ceciderunt de Israel septuaginta milia virorum.
1CHR|21|15|Misit quoque Deus angelum in Ierusalem, ut percuteret eam. Cumque percuteretur, vidit Dominus et misertus est super magnitudinem mali et imperavit angelo, qui percutiebat: " Sufficit, iam cesset manus tua ".Porro angelus Domini stabat iuxta aream Ornan Iebusaei.
1CHR|21|16|Levansque David oculos suos vidit angelum Domini stantem inter terram et caelum et evaginatum gladium in manu eius et versum contra Ierusalem; et ceciderunt tam ipse quam maiores natu vestiti ciliciis proni in terram.
1CHR|21|17|Dixitque David ad Deum: " Nonne ego sum, qui iussi, ut numeraretur populus? Ego qui peccavi, ego qui malum feci; iste grex quid commeruit? Domine Deus meus, vertatur, obsecro, manus tua in me et in domum patris mei; populus autem tuus non percutiatur ".
1CHR|21|18|Angelus autem Domini praecepit Gad dicere David, ut ascenderet exstrueretque altare Domino in area Ornan Iebusaei.
1CHR|21|19|Ascendit ergo David iuxta sermonem Gad, quem locutus fuerat ex nomine Domini.
1CHR|21|20|Porro Ornan, cum conversus vidisset angelum, quattuorque filii eius cum eo absconderunt se; nam eo tempore terebat in area triticum.
1CHR|21|21|Igitur, cum veniret David ad Ornan, conspexit eum Ornan et processit ei obviam de area et adoravit illum pronus in terram.
1CHR|21|22|Dixitque ei David: " Da mihi locum areae tuae, ut aedificem in ea altare Domino, ita ut quantum valet argenti accipias, et cesset plaga a populo ".
1CHR|21|23|Dixit autem Ornan ad David: " Tolle, et faciat dominus meus rex, quodcumque ei placet; sed et boves do in holocaustum et tribulas in ligna et triticum in sacrificium; omnia libens praebebo ".
1CHR|21|24|Dixitque ei rex David: " Nequaquam ita fiet, sed argentum dabo quantum valet; neque enim tibi auferre debeo et sic offerre Domino holocausta gratuita ".
1CHR|21|25|Dedit ergo David Ornan pro loco siclos auri iustissimi ponderis sescentos
1CHR|21|26|et aedificavit ibi altare Domino obtulitque holocausta et pacifica et invocavit Dominum. Et exaudivit eum in igne de caelo super altare holocausti,
1CHR|21|27|praecepitque Dominus angelo, et convertit gladium suum in vaginam.
1CHR|21|28|In illo ergo tempore David videns quod exaudisset eum Dominus in area Ornan Iebusaei immolavit ibi victimas.
1CHR|21|29|Tabernaculum autem Domini, quod fecerat Moyses in deserto, et altare holocaustorum ea tempestate erat in excelso Gabaon;
1CHR|21|30|et non praevaluit David ire, ut ibi obsecraret Deum; nimio enim fuerat timore perterritus videns gladium angeli Domini.
1CHR|22|1|Dixitque David: " Haec est domus Domini Dei, et hoc est altare holocausti pro Israel ".
1CHR|22|2|Et praecepit, ut congregarentur omnes advenae de terra Israel, et constituit ex eis latomos ad caedendos lapides et poliendos, ut aedificaretur domus Dei.
1CHR|22|3|Ferrum quoque plurimum ad clavos ianuarum et ad commissuras atque iuncturas praeparavit David et aeris pondus innumerabile.
1CHR|22|4|Ligna quoque cedrina non poterant aestimari, quae Sidonii et Tyrii deportaverant ad David.
1CHR|22|5|Et dixit David: " Salomon filius meus puer parvulus est et tener; domus autem, quae aedificanda est Domino, talis esse debet, ut in cunctis regionibus nominetur et glorificetur. Praeparabo ergo ei necessaria ". Et ob hanc causam ante mortem suam omnes paravit impensas.
1CHR|22|6|Vocavitque Salomonem filium suum et praecepit ei, ut aedificaret domum Domino, Deo Israel;
1CHR|22|7|dixitque David ad Salomonem: " Fili mi, voluntatis meae fuit, ut aedificarem domum nomini Domini Dei mei,
1CHR|22|8|sed factus est ad me sermo Domini dicens: "Multum sanguinem effudisti et magna bella bellasti. Non poteris aedificare domum nomini meo, tanto effuso sanguine coram me.
1CHR|22|9|Filius, qui nascetur tibi, erit vir quietissimus; faciam enim eum requiescere ab omnibus inimicis suis per circuitum et ob hanc causam Salomon vocabitur, et pacem et otium dabo in Israel cunctis diebus eius.
1CHR|22|10|Ipse aedificabit domum nomini meo, et ipse erit mihi in filium, et ego ero ei in patrem; firmaboque solium regni eius super Israel in aeternum".
1CHR|22|11|Nunc ergo, fili mi, sit Dominus tecum; et prosperare et aedifica domum Domino Deo tuo, sicut locutus est de te.
1CHR|22|12|Tantum det tibi Dominus prudentiam et sensum, ut regere possis Israel et custodire legem Domini Dei tui;
1CHR|22|13|tunc enim proficere poteris, si custodieris mandata et iudicia, quae praecepit Dominus Moysi super Israel. Confortare et viriliter age; ne timeas neque paveas.
1CHR|22|14|Ecce ego in labore meo praeparavi impensas domus Domini: auri talenta centum milia et argenti mille milia talentorum, aeris vero et ferri non est pondus, vincitur enim numerus magnitudine. Ligna et lapides praeparavi; tu autem ad ea adicies.
1CHR|22|15|Habes quoque plurimos artifices latomos et caementarios artificesque lignorum et omnium artium ad faciendum opus prudentissimos
1CHR|22|16|in auro et argento et aere et ferro, cuius non est numerus. Surge igitur et fac, et erit Dominus tecum ".
1CHR|22|17|Praecepit quoque David cunctis principibus Israel, ut adiuvarent Salomonem filium suum: "
1CHR|22|18|Cernitis, inquiens, quod Dominus Deus vester vobiscum sit et dederit vobis requiem per circuitum et tradiderit habitatores terrae in manu vestra, et subiecta sit terra coram Domino et coram populo eius.
1CHR|22|19|Praebete igitur corda vestra et animas vestras, ut quaeratis Dominum Deum vestrum; et consurgite et aedificate sanctuarium Domini Dei, ut introducatur arca foederis Domini et vasa Deo consecrata in domum, quae aedificatur nomini Domini ".
1CHR|23|1|Igitur David senex et plenus dierum regem constituit Sa lomonem filium suum super Israel
1CHR|23|2|et congregavit omnes principes Israel et sacerdotes atque Levitas.
1CHR|23|3|Numeratique sunt Levitae a triginta annis et supra, et inventa sunt triginta octo milia virorum.
1CHR|23|4|" Ex his, inquit, praesint ministerio domus Domini viginti quattuor milia, praepositi autem et iudices sex milia;
1CHR|23|5|porro quattuor milia ianitores et totidem psaltae canentes Domino in organis, quae feci ad canendum ".
1CHR|23|6|Et distribuit eos David per vices filiorum Levi Gerson videlicet et Caath et Merari.
1CHR|23|7|Filii Gerson: Ladan et Semei.
1CHR|23|8|Filii Ladan: princeps Iahiel et Zetham et Ioel, tres.
1CHR|23|9|Filii Semei: Salomith et Hoziel et Aran, tres; isti principes familiarum Ladan.
1CHR|23|10|Porro filii Semei: Iahath et Ziza et Iehus et Beria; isti filii Semei, quattuor.
1CHR|23|11|Erat autem Iahath prior, Ziza secundus; porro Iehus et Beria non habuerunt plurimos filios, et idcirco in una familia unaque domo computati sunt.
1CHR|23|12|Filii Caath: Amram et Isaar, Hebron et Oziel, quattuor.
1CHR|23|13|Filii Amram: Aaron et Moyses. Separatusque est Aaron, ut sanctificaret sanctissima, ipse et filii eius in sempiternum, et adoleret Domino et serviret ei ac benediceret in nomine eius in perpetuum.
1CHR|23|14|Moysi quoque hominis Dei filii annumerati sunt in tribu Levi.
1CHR|23|15|Filii Moysi: Gersam et Eliezer.
1CHR|23|16|Filii Gersam: Subael primus.
1CHR|23|17|Fuerunt autem filii Eliezer: Rohobia primus, et non erant Eliezer filii alii; porro filii Rohobia multiplicati sunt nimis.
1CHR|23|18|Filii Isaar: Salomoth primus.
1CHR|23|19|Filii Hebron: Ieriau primus, Amarias secundus, Iahaziel tertius, Iecmaam quartus.
1CHR|23|20|Filii Oziel: Micha primus, Iesia secundus.
1CHR|23|21|Filii Merari: Moholi et Musi. Filii Moholi: Eleazar et Cis;
1CHR|23|22|mortuus est autem Eleazar et non habuit filios sed filias acceperuntque eas filii Cis fratres earum.
1CHR|23|23|Filii Musi: Moholi et Eder et Ierimoth, tres.
1CHR|23|24|Hi filii Levi in familiis suis, principes familiarum per vices et numerum capitum singulorum, qui faciebant opera ministerii domus Domini a viginti annis et supra.
1CHR|23|25|Dixit enim David: " Requiem dedit Dominus, Deus Israel, populo suo et habitat in Ierusalem usque in aeternum;
1CHR|23|26|nec erit officii Levitarum, ut ultra portent tabernaculum et omnia vasa eius ad ministrandum.
1CHR|23|27|Iuxta praecepta igitur David novissima, supputabitur numerus filiorum Levi a viginti annis et supra,
1CHR|23|28|et erunt sub manu filiorum Aaron in cultum domus Domini pro atriis et exedris et in purificationem omnis rei sacrae et in ministerium templi Dei,
1CHR|23|29|pro panibus propositionis et farina oblationis et laganis azymorum et pro sartagine et ad torrendum et super omne pondus atque mensuram.
1CHR|23|30|Et stent mane ad confitendum et canendum Domino similiterque ad vesperam,
1CHR|23|31|tam in oblatione holocaustorum Domini quam in sabbatis et calendis et sollemnitatibus reliquis, iuxta numerum et caeremonias uniuscuiusque rei iugiter coram Domino.
1CHR|23|32|Et custodiant observationes tabernaculi conventus et ritum sanctuarii et observationem filiorum Aaron fratrum suorum, ut ministrent in domo Domini ".
1CHR|24|1|Porro filiis Aaron hae partiones erant.Filii Aaron: Nadab et Abiu et Eleazar et Ithamar.
1CHR|24|2|Mortui sunt autem Nadab et Abiu ante patrem suum absque liberis; sacerdotioque functus est Eleazar et Ithamar.
1CHR|24|3|Et divisit eos David cum Sadoc de filiis Eleazari et cum Achimelech de filiis Ithamar, secundum vices suas et ministerium.
1CHR|24|4|Inventique sunt multo plures filii Eleazar secundum capita virorum quam filii Ithamar; divisit igitur eis, hoc est filiis Eleazar principes per familias sedecim, et filiis Ithamar per familias et domos suas octo.
1CHR|24|5|Porro divisit utrasque inter se familias sortibus; erant enim principes sanctuarii et principes Dei tam de filiis Eleazar quam de filiis Ithamar.
1CHR|24|6|Descripsitque eos Semeias filius Nathanael scriba Levites coram rege et principibus et Sadoc sacerdote et Achimelech filio Abiathar, principibus quoque familiarum sacerdotalium et leviticarum: unam familiam pro Eleazar et unam pro Ithamar.
1CHR|24|7|Exivit autem sors prima Ioiarib, secunda Iedaiae,
1CHR|24|8|tertia Harim, quarta Seorim,
1CHR|24|9|quinta Melchia, sexta Miamin,
1CHR|24|10|septima Accos, octava Abia,
1CHR|24|11|nona Iesua, decima Sechenia,
1CHR|24|12|undecima Eliasib, duodecima Iacim,
1CHR|24|13|tertia decima Hoppha, quarta decima Isbaab,
1CHR|24|14|quinta decima Belga, sexta decima Emmer,
1CHR|24|15|septima decima Hezir, octava decima Aphses,
1CHR|24|16|nona decima Phethahia, vicesima Hezechiel,
1CHR|24|17|vicesima prima Iachin, vicesima secunda Gamul,
1CHR|24|18|vicesima tertia Dalaiau, vicesima quarta Maaziau.
1CHR|24|19|Hae vices eorum secundum ministeria sua, ut ingrediantur domum Domini, et iuxta ritum suum sub manu Aaron patris eorum, sicut praecepit Dominus, Deus Israel.
1CHR|24|20|Porro filiorum Levi, qui reliqui fuerant: de filiis Amram Subael et de filiis Subael Iehedeia.
1CHR|24|21|De filiis quoque Rohobiae princeps Iesias.
1CHR|24|22|De Isaaritis vero Salomoth; de filiis Salomoth Iahath.
1CHR|24|23|De Hebronitis: Ieriau, Amarias secundus, Iahaziel tertius, Iecmaam quartus.
1CHR|24|24|Filius Oziel Micha; de filiis Micha Samir;
1CHR|24|25|frater Micha Iesia; de filiis Iesiae Zacharias.
1CHR|24|26|Filii Merari: Moholi et Musi. Filii eius: Iaziau et Bani.
1CHR|24|27|Filius Merari: de Iaziau filio suo Soam et Zacchur et Hebri.
1CHR|24|28|Porro de Moholi filius Eleazar, qui non habebat liberos.
1CHR|24|29|Filius vero Cis Ierameel;
1CHR|24|30|filii Musi: Moholi, Eder et Ierimoth.Isti filii Levi secundum familias suas.
1CHR|24|31|Ipsi quoque miserunt sortes sicut fratres sui, filii Aaron coram David rege et Sadoc et Achimelech et principibus familiarum sacerdotalium et leviticarum tam maiores quam minores; omnes sors aequaliter dividebat.
1CHR|25|1|Igitur David et magistratus exercitus segregaverunt in ministerium filios Asaph et Heman et Idithun, qui prophetarent in citharis et psalteriis et cymbalis, secundum numerum suum dedicato sibi officio servientes.
1CHR|25|2|De filiis Asaph: Zacchur et Ioseph et Nathania et Asarela filii Asaph erant sub manu Asaph prophetantis sub manu regis.
1CHR|25|3|De Idithun; filii Idithun: Godolias, Sori, Iesaias et Hasabias et Matthathias, sex, sub manu patris sui Idithun, qui in cithara prophetabat ad confitendum et laudandum Dominum.
1CHR|25|4|De Heman quoque; filii Heman: Bocciau, Matthaniau, Oziel, Subael et Ierimoth, Hananias, Hanani, Eliatha, Geddelthi et Romemthiezer et Iesbacasa, Mellothi, Othir, Mahazioth;
1CHR|25|5|omnes isti filii Heman videntis regis iuxta sermones Dei, quod exaltaret cornu eius; deditque Deus Heman filios quattuordecim et filias tres.
1CHR|25|6|Universi sub manu patris sui ad cantandum in templo Domini distributi erant in cymbalis et psalteriis et citharis, in ministeria domus Dei sub manu regis: Asaph et Idithun et Heman.
1CHR|25|7|Fuit autem numerus eorum cum fratribus suis eruditis in cantando Domino, cuncti magistri, ducenti octoginta octo.
1CHR|25|8|Miseruntque sortes pro ministerio ex aequo, tam maior quam minor, magister pariter et discipulus.
1CHR|25|9|Egressaque est sors prima Ioseph, qui erat de Asaph. Secunda Godoliae, ipsi et fratribus eius et filiis eius, duodecim.
1CHR|25|10|Tertia Zacchur, filiis et fratribus eius, duodecim.
1CHR|25|11|Quarta Isari, filiis et fratribus eius, duodecim.
1CHR|25|12|Quinta Nathaniau, filiis et fratribus eius, duodecim.
1CHR|25|13|Sexta Bocciau, filiis et fratribus eius, duodecim.
1CHR|25|14|Septima Isreela, filiis et fratribus eius, duodecim.
1CHR|25|15|Octava Iesaiae, filiis et fratribus eius, duodecim.
1CHR|25|16|Nona Matthaniau, filiis et fratribus eius, duodecim.
1CHR|25|17|Decima Semei, filiis et fratribus eius, duodecim.
1CHR|25|18|Undecima Azareel, filiis et fratribus eius, duodecim.
1CHR|25|19|Duodecima Hasabiae, filiis et fratribus eius, duodecim.
1CHR|25|20|Tertia decima Subael, filiis et fratribus eius, duodecim.
1CHR|25|21|Quarta decima Matthathiae, filiis et fratribus eius, duodecim.
1CHR|25|22|Quinta decima Ierimoth, filiis et fratribus eius, duodecim.
1CHR|25|23|Sexta decima Hananiae, filiis et fratribus eius, duodecim.
1CHR|25|24|Septima decima Iesbacasae, filiis et fratribus eius, duodecim.
1CHR|25|25|Octava decima Hanani, filiis et fratribus eius, duodecim.
1CHR|25|26|Nona decima Mellothi, filiis et fratribus eius, duodecim.
1CHR|25|27|Vicesima Eliatha, filiis et fratribus eius, duodecim.
1CHR|25|28|Vicesima prima Othir, filiis et fratribus eius, duodecim.
1CHR|25|29|Vicesima secunda Geddelthi, filiis et fratribus eius, duodecim.
1CHR|25|30|Vicesima tertia Mahazioth, filiis et fratribus eius, duodecim.
1CHR|25|31|Vicesima quarta Romemthiezer, filiis et fratribus eius, duodecim.
1CHR|26|1|Divisiones autem ianitorum.De Coritis: Meselemia filius Core de filiis Abiasaph.
1CHR|26|2|Filii Meselemiae: Zacharias primogenitus, Iedihel secundus, Zabadias tertius, Iathanael quartus,
1CHR|26|3|Elam quintus, Iohanan sextus, Elioenai septimus.
1CHR|26|4|Filii autem Obededom: Semeias primogenitus, Iozabad secundus, Ioah tertius, Sachar quartus, Nathanael quintus,
1CHR|26|5|Ammiel sextus, Issachar septimus, Phollathi octavus, quia benedixit illi Deus.
1CHR|26|6|Semeiae autem filio eius nati sunt filii praefecti familiarum suarum, erant enim viri fortissimi;
1CHR|26|7|filii ergo Semeiae: Othni et Raphael et Obed, Elzabad, fratres eius viri fortissimi, Eliu quoque et Samachias;
1CHR|26|8|omnes hi de filiis Obededom, ipsi et filii et fratres eorum fortissimi ad ministrandum sexaginta duo de Obededom.
1CHR|26|9|Porro Meselemiae filii et fratres eorum robustissimi decem et octo.
1CHR|26|10|De Hosa autem, de filiis Merari, erant filii: Semri princeps - non enim fuerat primogenitus, et idcirco posuerat eum pater eius in principem -
1CHR|26|11|Helcias secundus, Tabelias tertius, Zacharias quartus; omnes hi filii et fratres Hosa tredecim.
1CHR|26|12|Hae divisiones ianitorum: secundum capita virorum habebant ministeria sicut et fratres eorum ad ministrandum in domo Domini.
1CHR|26|13|Missae sunt ergo sortes ex aequo et parvis et magnis per familias suas in unamquamque portarum.
1CHR|26|14|Cecidit igitur sors orientalis Selemiae; porro Zachariae filio eius consiliario prudentissimo et erudito sortito obtigit plaga septentrionalis;
1CHR|26|15|Obededom vero australis, et filiis eius horreum;
1CHR|26|16|Sephim et Hosa occidentalis iuxta portam Sallecheth apud viam ascensionis. Custodia iuxta custodiam:
1CHR|26|17|ad orientem per diem sex et ad aquilonem quattuor per diem, atque ad meridiem similiter in die quattuor et pro horreo bini et bini,
1CHR|26|18|pro Parbar quoque ad occidentem quattuor in via, duo pro Parbar.
1CHR|26|19|Hae sunt divisiones ianitorum filiorum Core et Merari.
1CHR|26|20|Porro Levitae fratres eorum super thesauros domus Dei ac thesauros rerum consecratarum.
1CHR|26|21|De filiis Ladan Gersonitae principes familiarum Ladan Gersonitae erant Iahielitae.
1CHR|26|22|Filii Iahiel et Zetham et Ioel fratrum eius erant super thesauros domus Domini.
1CHR|26|23|De Amramitis et Isaaritis et Hebronitis et Ozielitis:
1CHR|26|24|Subael filius Gersam filii Moysi praepositus thesauris.
1CHR|26|25|Fratres quoque eius Eliezer, cuius filius Rohobia et huius filius Iesaias; et huius filius Ioram, huius quoque filius Zechri et huius filius Selemith.
1CHR|26|26|Ipse Selemith et fratres eius super omnes thesauros rerum consecratarum, quas sanctificavit David rex et principes familiarum et tribuni et centuriones et duces exercitus
1CHR|26|27|de bellis et manubiis proeliorum, quas consecraverant ad sustentandum templum Domini.
1CHR|26|28|Et universa, quae consecraverant Samuel videns et Saul filius Cis et Abner filius Ner et Ioab filius Sarviae, omnia donaria sacra erant sub manu Selemith et fratrum eius.
1CHR|26|29|De Isaaritis vero erant Chonenias et filii eius ad opera forinsecus super Israel praefecti et iudices.
1CHR|26|30|Porro de Hebronitis Hasabias et fratres eius viri strenui mille septingenti erant magistratus Israel trans Iordanem contra occidentem in cunctis operibus Domini et in ministerium regis;
1CHR|26|31|Hebronitarum autem princeps fuit Ieria secundum cognationes et familias eorum. Quadragesimo anno regni David recensiti sunt et inventi viri fortes in Iazer Galaad
1CHR|26|32|fratresque eius viri strenui duo milia septingenti principes familiarum; praeposuit autem eos David rex Rubenitis et Gadditis et dimidio tribus Manasse in omne ministerium Dei et regis.
1CHR|27|1|Filii autem Israel secundum numerum suum, principes fa miliarum, tribuni et centuriones et praefecti, qui ministrabant regi iuxta turmas suas ingredientes et egredientes per singulos menses in anno, unaquaeque turma viginti quattuor milia.
1CHR|27|2|Primae turmae in primo mense Iesbaam praeerat filius Zabdiel, et sub eo viginti quattuor milia;
1CHR|27|3|erat de filiis Phares princeps cunctorum principum in exercitu mense primo.
1CHR|27|4|Secundi mensis habebat turmam Dudi Ahohites, et sub eo viginti quattuor milia.
1CHR|27|5|Dux quoque turmae tertiae in mense tertio erat Banaias filius Ioiadae sacerdotis, et in divisione sua viginti quattuor milia;
1CHR|27|6|ipse est Banaias fortissimus inter triginta et super triginta; praeerat autem turmae ipsius Amizabad filius eius.
1CHR|27|7|Quartus, mense quarto, Asael frater Ioab et Zabadias filius eius post eum, et in turma eius viginti quattuor milia.
1CHR|27|8|Quintus, mense quinto, princeps Samaoth Zaraita, et in turma eius viginti quattuor milia.
1CHR|27|9|Sextus, mense sexto, Hira filius Acces Thecuites, et in turma eius viginti quattuor milia.
1CHR|27|10|Septimus, mense septimo, Helles Phalonites de filiis Ephraim, et in turma eius viginti quattuor milia.
1CHR|27|11|Octavus, mense octavo, Sobbochai Husathites de stirpe Zara, et in turma eius viginti quattuor milia.
1CHR|27|12|Nonus, mense nono, Abiezer Anathothites de filiis Beniamin, et in turma eius viginti quattuor milia.
1CHR|27|13|Decimus, mense decimo, Maharai Netophathites de stirpe Zara, et in turma eius viginti quattuor milia.
1CHR|27|14|Undecimus, mense undecimo, Banaias Pharathonites de filiis Ephraim, et in turma eius viginti quattuor milia.
1CHR|27|15|Duodecimus, mense duodecimo, Holdai Netophathites de stirpe Othoniel, et in turma eius viginti quattuor milia.
1CHR|27|16|Porro tribubus praeerant Israel: Rubenitis dux Eliezer filius Zechri; Simeonitis Saphatia filius Maacha;
1CHR|27|17|Levitis Hasabias filius Camuel; Aaronitis Sadoc;
1CHR|27|18|Iudae Eliu de fratribus David; Issachar Amri filius Michael;
1CHR|27|19|Zabulon Iesmaias filius Abdiae; Nephthali Ierimoth filius Azriel;
1CHR|27|20|filiis Ephraim Osee filius Ozaziu; dimidio tribus Manasse Ioel filius Phadaiae;
1CHR|27|21|et dimidio tribus Manasse in Galaad Iaddo filius Zachariae; Beniamin autem Iasiel filius Abner;
1CHR|27|22|Dan vero Azareel filius Ieroham: hi principes tribuum Israel.
1CHR|27|23|Noluit autem David numerare eos a viginti annis inferius, quia dixerat Dominus ut multiplicaret Israel quasi stellas caeli.
1CHR|27|24|Ioab filius Sarviae coeperat numerare nec complevit, quia super hoc ira irruerat in Israel, et idcirco numerus non est relatus in librum annalium regis David.
1CHR|27|25|Super thesauros autem regis fuit Azmaveth filius Adiel; his autem thesauris, qui erant in regione, in urbibus et in vicis et in turribus praesidebat Ionathan filius Oziae.
1CHR|27|26|Operi autem rustico et agricolis, qui exercebant terram, praeerat Ezri filius Chelub.
1CHR|27|27|Vinearumque cultoribus Semei Ramathites; cellis autem vinariis in vineis Zabdi Sephamatites.
1CHR|27|28|Nam super oliveta et ficeta, quae erant in Sephela, Baalhanan Gederites; super apothecas autem olei Ioas.
1CHR|27|29|Porro armentis, quae pascebantur in Saron, praepositus fuit Setrai Saronites, et super boves in vallibus Saphat filius Adli.
1CHR|27|30|Super camelos vero Ubil Ismaelites, et super asinas Iehedeia Meronathites;
1CHR|27|31|super oves quoque Iaziz Agarenus: omnes hi principes substantiae regis David.
1CHR|27|32|Ionathan autem patruus David consiliarius, vir prudens et litteratus, ipse et Iahiel filius Hachamonitis erant cum filiis regis.
1CHR|27|33|Achitophel etiam consiliarius regis, et Chusai Arachites amicus regis;
1CHR|27|34|post Achitophel fuit Ioiada filius Banaiae et Abiathar. Princeps autem exercitus regis erat Ioab.
1CHR|28|1|Convocavit igitur David om nes principes Israel, duces tri buum et praepositos turmarum, qui ministrabant regi, tribunos quoque et centuriones et, qui praeerant substantiae et gregibus regis filiorumque suorum, cum eunuchis et fortibus et robustissimis quibusque in exercitu Ierusalem.
1CHR|28|2|Cumque surrexisset rex et stetisset, ait: " Audite me, fratres mei et populus meus. Cogitavi ut aedificarem domum, in qua requiesceret arca foederis Domini et scabellum pedum Dei nostri, et ad aedificandum omnia praeparavi;
1CHR|28|3|Deus autem dixit mihi: "Non aedificabis domum nomini meo, eo quod sis vir bellator et sanguinem fuderis".
1CHR|28|4|Sed elegit Dominus, Deus Israel, me de universa domo patris mei, ut essem rex super Israel in sempiternum; Iudam enim elegit principem, porro in domo Iudae domum patris mei, et in filiis patris mei placuit ei, ut me eligeret regem super cunctum Israel.
1CHR|28|5|Sed et de filiis meis - filios enim multos dedit mihi Dominus - elegit Salomonem filium meum, ut sederet in throno regni Domini super Israel.
1CHR|28|6|Dixitque mihi: "Salomon filius tuus aedificabit domum meam et atria mea; ipsum enim elegi mihi in filium, et ego ero ei in patrem.
1CHR|28|7|Et firmabo regnum eius usque in aeternum, si perseveraverit facere praecepta mea et iudicia, sicut et hodie".
1CHR|28|8|Nunc igitur coram universo Israel coetu Domini, audiente Deo nostro, custodite et perquirite cuncta mandata Domini Dei vestri, ut possideatis terram bonam et relinquatis eam in hereditatem filiis vestris post vos usque in sempiternum.
1CHR|28|9|Tu autem, Salomon, fili mi, scito Deum patris tui et servi ei corde perfecto et animo voluntario; omnia enim corda scrutatur Dominus et universas mentium cogitationes intellegit. Si quaesieris eum, invenies; si autem dereliqueris illum, proiciet te in aeternum.
1CHR|28|10|Nunc ergo vide quia elegit te Dominus, ut aedificares domum sanctuarii; confortare et perfice ".
1CHR|28|11|Dedit autem David Salomoni filio suo descriptionem porticus et templi et cellariorum et cenaculorum et cubiculorum interiorum et domus propitiatorii
1CHR|28|12|necnon et omnium, quae per Spiritum cum eo erant, de atriis domus Domini et de omnibus exedris per circuitum, de thesauris domus Dei et de thesauris rerum consecratarum
1CHR|28|13|et de divisionibus sacerdotalibus et leviticis, de omni opere ministerii domus Domini et de universis vasis ministerii templi Domini,
1CHR|28|14|de auro in pondere per singula vasa ministerii, de omnibus vasis argenteis in pondere per omnia vasa pro operum diversitate;
1CHR|28|15|sed et ad candelabra aurea et ad lucernas eorum aurum pro mensura uniuscuiusque candelabri et lucernarum, similiter et in candelabris argenteis et in lucernis eorum pro diversitate mensurae, pondus argenti indicavit.
1CHR|28|16|Aurum quoque in mensas propositionis pro diversitate mensarum, similiter et argentum in alias mensas argenteas;
1CHR|28|17|ad fuscinulas quoque et phialas et crateras ex auro purissimo et scyphos aureos pro qualitate mensurae pondus distribuit in scyphum et scyphum; similiter et in scyphos argenteos diversum argenti pondus constituit,
1CHR|28|18|altari autem, in quo adoletur incensum, aurum purissimum, et aurum pro structura quadrigae cherubim extendentium alas et velantium arcam foederis Domini.
1CHR|28|19|" Omnia, inquit, venerunt scripta manu Domini ad me, ut intellegerem universa opera exemplaris ".
1CHR|28|20|Dixit quoque David Salomoni filio suo: " Viriliter age et confortare et fac, ne timeas et ne paveas; Dominus enim Deus meus tecum erit et non dimittet te nec derelinquet, donec perficias omne opus ministerii domus Domini.
1CHR|28|21|Ecce divisiones sacerdotum et Levitarum: parati erunt in omne ministerium domus Dei; et assistet tibi in omni opere quisquis in sapientia ad omne ministerium promptus fuerit, principes quoque et universus populus in negotiis tuis ".
1CHR|29|1|Locutusque est David rex ad omnem ecclesiam: " Salomo nem filium meum unum elegit Deus adhuc puerum et tenellum; opus autem grande est: neque enim homini praeparatur habitatio sed Domino Deo.
1CHR|29|2|Ego autem totis viribus meis praeparavi impensas domus Dei mei: aurum ad vasa aurea et argentum in argentea, aes in aenea, ferrum in ferrea, ligna ad lignea, lapides onychinos et ad inserendum, durum caementum et lapides diversorum colorum omnemque pretiosum lapidem et marmor Parium abundantissime.
1CHR|29|3|Et super haec, cum delectarer super domo Dei mei, de peculio meo aurum et argentum do in templum Dei mei, exceptis his, quae paravi in aedem sanctam:
1CHR|29|4|tria milia talenta auri de auro Ophir et septem milia talentorum argenti probatissimi ad operiendos parietes templi;
1CHR|29|5|et ubicumque opus est aurum pro aureis, et ubicumque opus est argentum pro argenteis et pro quolibet opere per manus artificum; et si quis sponte offert, impleat manum suam hodie et offerat, quod voluerit, Domino ".
1CHR|29|6|Sponte obtulerunt itaque principes familiarum et proceres tribuum Israel, tribuni quoque et centuriones et principes operis regis;
1CHR|29|7|dederuntque in opera domus Dei auri talenta quinque milia et solidos decem milia, argenti talenta decem milia et aeris talenta decem et octo milia, ferri quoque centum milia talentorum.
1CHR|29|8|Et apud quemcumque inventi sunt lapides, dederunt in thesaurum domus Domini in manum Iahiel Gersonitis.
1CHR|29|9|Laetatusque est populus super prompto animo eorum, quia corde toto offerebant ea Domino; sed et David rex laetatus est gaudio magno.
1CHR|29|10|Et benedixit Domino coram universa multitudine et ait: Benedictus es, Domine, Deus Israel patris nostri,ab aeterno in aeternum.
1CHR|29|11|Tua est, Domine, magnificentia et potentia,gloria, splendor atque maiestas.Cuncta enim, quae in caelo sunt et in terra, tua sunt.Tuum, Domine, regnum, et tu elevaris ut caput super omnia.
1CHR|29|12|De te sunt divitiae et gloria,tu dominaris omnium.In manu tua virtus et potentia,in manu tua est magnificare et firmare omnia.
1CHR|29|13|Nunc igitur, Deus noster, confitemur tibiet laudamus nomen tuum inclitum.
1CHR|29|14|Quis ego, et quis populus meus, ut possimus haec tibi universa offerre? Tua sunt haec omnia; et, quae de manu tua accepimus, dedimus tibi.
1CHR|29|15|Peregrini enim sumus coram te et advenae, sicut omnes patres nostri; dies nostri quasi umbra super terram, et nulla est spes.
1CHR|29|16|Domine Deus noster, omnis haec copia, quam paravimus, ut aedificaretur domus nomini sancto tuo, de manu tua est, et tua sunt omnia.
1CHR|29|17|Scio, Deus meus, quod probes corda et simplicitatem diligas; unde et ego in simplicitate cordis mei laetus obtuli universa haec et populum tuum, qui hic repertus est, vidi cum ingenti gaudio sponte tibi offerre donaria.
1CHR|29|18|Domine, Deus Abraham et Isaac et Israel patrum nostrorum, custodi in aeternum hanc voluntatem cordis eorum; et semper in venerationem tui mens ista permaneat.
1CHR|29|19|Salomoni quoque filio meo da cor perfectum, ut custodiat mandata tua, testimonia tua et legitima tua et faciat universa et aedificet aedem, cuius impensas paravi ".
1CHR|29|20|Praecepit autem David universae ecclesiae: " Benedicite Domino Deo vestro! ". Et benedixit omnis ecclesia Domino, Deo patrum suorum; et inclinaverunt se et adoraverunt Deum et deinde regem.
1CHR|29|21|Immolaveruntque victimas Domino et obtulerunt holocausta die sequenti, tauros mille, arietes mille, agnos mille cum libaminibus suis et sacrificia abundantissime in omnem Israel.
1CHR|29|22|Et comederunt et biberunt coram Domino in die illo cum grandi laetitia; et fecerunt regem secundo Salomonem filium David atque unxerunt Domino in principem et Sadoc in pontificem.
1CHR|29|23|Seditque Salomon super solium Domini, ut esset rex pro David patre suo, et prosperatus est, et paruit illi omnis Israel.
1CHR|29|24|Sed et universi principes et fortes et cuncti filii regis David dederunt manum subicientes se Salomoni regi.
1CHR|29|25|Magnificavit ergo Dominus Salomonem in excelsum in conspectu omnis Israel et dedit illi gloriam regni, qualem nullus habuit ante eum rex Israel.
1CHR|29|26|Igitur David filius Isai regnavit super universum Israel;
1CHR|29|27|et dies, quibus regnavit super Israel, fuerunt quadraginta anni: in Hebron regnavit septem annis et in Ierusalem annis triginta tribus.
1CHR|29|28|Et mortuus est in senectute bona plenus dierum et divitiis et gloria; et regnavit Salomon filius eius pro eo.
1CHR|29|29|Gesta autem David regis priora et novissima scripta sunt in libro Samuel videntis et in libro Nathan prophetae atque in volumine Gad videntis,
1CHR|29|30|universique regni eius et fortitudinis et temporum, quae transierunt sub eo sive in Israel sive in cunctis regnis terrarum.
