JONAH|1|1|et factum est verbum Domini ad Ionam filium Amathi dicens
JONAH|1|2|surge vade in Nineven civitatem grandem et praedica in ea quia ascendit malitia eius coram me
JONAH|1|3|et surrexit Iona ut fugeret in Tharsis a facie Domini et descendit Ioppen et invenit navem euntem in Tharsis et dedit naulum eius et descendit in eam ut iret cum eis in Tharsis a facie Domini
JONAH|1|4|Dominus autem misit ventum magnum in mari et facta est tempestas magna in mari et navis periclitabatur conteri
JONAH|1|5|et timuerunt nautae et clamaverunt viri ad deum suum et miserunt vasa quae erant in navi in mare ut adleviaretur ab eis et Iona descendit ad interiora navis et dormiebat sopore gravi
JONAH|1|6|et accessit ad eum gubernator et dixit ei quid tu sopore deprimeris surge invoca Deum tuum si forte recogitet Deus de nobis et non pereamus
JONAH|1|7|et dixit vir ad collegam suum venite et mittamus sortes et sciamus quare hoc malum sit nobis et miserunt sortes et cecidit sors super Ionam
JONAH|1|8|et dixerunt ad eum indica nobis cuius causa malum istud sit nobis quod est opus tuum quae terra tua et quo vel ex quo populo es tu
JONAH|1|9|et dixit ad eos Hebraeus ego sum et Dominum Deum caeli ego timeo qui fecit mare et aridam
JONAH|1|10|et timuerunt viri timore magno et dixerunt ad eum quid hoc fecisti cognoverunt enim viri quod a facie Domini fugeret quia indicaverat eis
JONAH|1|11|et dixerunt ad eum quid faciemus tibi et cessabit mare a nobis quia mare ibat et intumescebat
JONAH|1|12|et dixit ad eos tollite me et mittite in mare et cessabit mare a vobis scio enim ego quoniam propter me tempestas grandis haec super vos
JONAH|1|13|et remigabant viri ut reverterentur ad aridam et non valebant quia mare ibat et intumescebat super eos
JONAH|1|14|et clamaverunt ad Dominum et dixerunt quaesumus Domine ne pereamus in anima viri istius et ne des super nos sanguinem innocentem quia tu Domine sicut voluisti fecisti
JONAH|1|15|et tulerunt Ionam et miserunt in mare et stetit mare a fervore suo
JONAH|1|16|et timuerunt viri timore magno Dominum et immolaverunt hostias Domino et voverunt vota
JONAH|2|1|et praeparavit Dominus piscem grandem ut degluttiret Ionam et erat Iona in ventre piscis tribus diebus et tribus noctibus
JONAH|2|2|et oravit Iona ad Dominum Deum suum de utero piscis
JONAH|2|3|et dixit clamavi de tribulatione mea ad Dominum et exaudivit me de ventre inferni clamavi et exaudisti vocem meam
JONAH|2|4|et proiecisti me in profundum in corde maris et flumen circumdedit me omnes gurgites tui et fluctus tui super me transierunt
JONAH|2|5|et ego dixi abiectus sum a conspectu oculorum tuorum verumtamen rursus videbo templum sanctum tuum
JONAH|2|6|circumdederunt me aquae usque ad animam abyssus vallavit me pelagus operuit caput meum
JONAH|2|7|ad extrema montium descendi terrae vectes concluserunt me in aeternum et sublevabis de corruptione vitam meam Domine Deus meus
JONAH|2|8|cum angustiaretur in me anima mea Domini recordatus sum ut veniat ad te oratio mea ad templum sanctum tuum
JONAH|2|9|qui custodiunt vanitates frustra misericordiam suam derelinquunt
JONAH|2|10|ego autem in voce laudis immolabo tibi quaecumque vovi reddam pro salute Domino
JONAH|2|11|et dixit Dominus pisci et evomuit Ionam in aridam
JONAH|3|1|et factum est verbum Domini ad Ionam secundo dicens
JONAH|3|2|surge vade ad Nineven civitatem magnam et praedica in ea praedicationem quam ego loquor ad te
JONAH|3|3|et surrexit Iona et abiit in Nineven iuxta verbum Domini et Nineve erat civitas magna Dei itinere dierum trium
JONAH|3|4|et coepit Iona introire in civitatem itinere diei unius et clamavit et dixit adhuc quadraginta dies et Nineve subvertetur
JONAH|3|5|et crediderunt viri ninevitae in Deo et praedicaverunt ieiunium et vestiti sunt saccis a maiore usque ad minorem
JONAH|3|6|et pervenit verbum ad regem Nineve et surrexit de solio suo et abiecit vestimentum suum a se et indutus est sacco et sedit in cinere
JONAH|3|7|et clamavit et dixit in Nineve ex ore regis et principum eius dicens homines et iumenta et boves et pecora non gustent quicquam nec pascantur et aquam non bibant
JONAH|3|8|et operiantur saccis homines et iumenta et clament ad Dominum in fortitudine et convertatur vir a via sua mala et ab iniquitate quae est in manibus eorum
JONAH|3|9|quis scit si convertatur et ignoscat Deus et revertatur a furore irae suae et non peribimus
JONAH|3|10|et vidit Deus opera eorum quia conversi sunt a via sua mala et misertus est Deus super malitiam quam locutus fuerat ut faceret eis et non fecit
JONAH|4|1|et adflictus est Iona adflictione magna et iratus est
JONAH|4|2|et oravit ad Dominum et dixit obsecro Domine numquid non hoc est verbum meum cum adhuc essem in terra mea propter hoc praeoccupavi ut fugerem in Tharsis scio enim quia tu Deus clemens et misericors es patiens et multae miserationis et ignoscens super malitia
JONAH|4|3|et nunc Domine tolle quaeso animam meam a me quia melior est mihi mors quam vita
JONAH|4|4|et dixit Dominus putasne bene irasceris tu
JONAH|4|5|et egressus est Iona de civitate et sedit contra orientem civitatis et fecit sibimet ibi umbraculum et sedebat subter eum in umbra donec videret quid accideret civitati
JONAH|4|6|et praeparavit Dominus Deus hederam et ascendit super caput Ionae ut esset umbra super caput eius et protegeret eum laboraverat enim et laetatus est Iona super hedera laetitia magna
JONAH|4|7|et paravit Deus vermem ascensu diluculo in crastinum et percussit hederam et exaruit
JONAH|4|8|et cum ortus fuisset sol praecepit Dominus vento calido et urenti et percussit sol super caput Ionae et aestuabat et petivit animae suae ut moreretur et dixit melius est mihi mori quam vivere
JONAH|4|9|et dixit Dominus ad Ionam putasne bene irasceris tu super hederam et dixit bene irascor ego usque ad mortem
JONAH|4|10|et dixit Dominus tu doles super hederam in qua non laborasti neque fecisti ut cresceret quae sub una nocte nata est et una nocte periit
JONAH|4|11|et ego non parcam Nineve civitati magnae in qua sunt plus quam centum viginti milia hominum qui nesciunt quid sit inter dexteram et sinistram suam et iumenta multa
