OBAD|1|1|Видение Авдия. Так говорит Господь Бог об Едоме: весть услышали мы от Господа, и посол послан [объявить] народам: "вставайте, и выступим против него войною!"
OBAD|1|2|Вот, Я сделал тебя малым между народами, и ты в большом презрении.
OBAD|1|3|Гордость сердца твоего обольстила тебя; ты живешь в расселинах скал, на возвышенном месте, и говоришь в сердце твоем: "кто низринет меня на землю?"
OBAD|1|4|Но хотя бы ты, как орел, поднялся высоко и среди звезд устроил гнездо твое, то и оттуда Я низрину тебя, говорит Господь.
OBAD|1|5|Не воры ли приходили к тебе? не ночные ли грабители, что ты так разорен? Но они украли бы столько, сколько надобно им. Если бы проникли к тебе обиратели винограда, то и они разве не оставили бы несколько ягод?
OBAD|1|6|Как обобрано все у Исава и обысканы тайники его!
OBAD|1|7|До границы выпроводят тебя все союзники твои, обманут тебя, одолеют тебя живущие с тобою в мире, ядущие хлеб твой нанесут тебе удар. Нет в нем смысла!
OBAD|1|8|Не в тот ли день это будет, говорит Господь, когда Я истреблю мудрых в Едоме и благоразумных на горе Исава?
OBAD|1|9|Поражены будут страхом храбрецы твои, Феман, дабы все на горе Исава истреблены были убийством.
OBAD|1|10|За притеснение брата твоего, Иакова, покроет тебя стыд и ты истреблен будешь навсегда.
OBAD|1|11|В тот день, когда ты стоял напротив, в тот день, когда чужие уводили войско его в плен и иноплеменники вошли в ворота его и бросали жребий о Иерусалиме, ты был как один из них.
OBAD|1|12|Не следовало бы тебе злорадно смотреть на день брата твоего, на день отчуждения его; не следовало бы радоваться о сынах Иуды в день гибели их и расширять рот в день бедствия.
OBAD|1|13|Не следовало бы тебе входить в ворота народа Моего в день несчастья его и даже смотреть на злополучие его в день погибели его, ни касаться имущества его в день бедствия его,
OBAD|1|14|ни стоять на перекрестках для убивания бежавших его, ни выдавать уцелевших из него в день бедствия.
OBAD|1|15|Ибо близок день Господень на все народы: как ты поступал, так поступлено будет и с тобою; воздаяние твое обратится на голову твою.
OBAD|1|16|Ибо, как вы пили на святой горе Моей, так все народы всегда будут пить, будут пить, проглотят и будут, как бы их не было.
OBAD|1|17|А на горе Сионе будет спасение, и будет она святынею; и дом Иакова получит во владение наследие свое.
OBAD|1|18|И дом Иакова будет огнем, и дом Иосифа – пламенем, а дом Исавов – соломою: зажгут его, и истребят его, и никого не останется из дома Исава: ибо Господь сказал это.
OBAD|1|19|И завладеют те, которые к югу, горою Исава, а которые в долине, – Филистимлянами; и завладеют полем Ефрема и полем Самарии, а Вениамин завладеет Галаадом.
OBAD|1|20|И переселенные из войска сынов Израилевых завладеют землею Ханаанскою до Сарепты, а переселенные из Иерусалима, находящиеся в Сефараде, получат во владение города южные.
OBAD|1|21|И придут спасители на гору Сион, чтобы судить гору Исава, и будет царство Господа.
