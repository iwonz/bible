NUM|1|1|The LORD spoke to Moses in the Tent of Meeting in the Desert of Sinai on the first day of the second month of the second year after the Israelites came out of Egypt. He said:
NUM|1|2|"Take a census of the whole Israelite community by their clans and families, listing every man by name, one by one.
NUM|1|3|You and Aaron are to number by their divisions all the men in Israel twenty years old or more who are able to serve in the army.
NUM|1|4|One man from each tribe, each the head of his family, is to help you.
NUM|1|5|These are the names of the men who are to assist you: from Reuben, Elizur son of Shedeur;
NUM|1|6|from Simeon, Shelumiel son of Zurishaddai;
NUM|1|7|from Judah, Nahshon son of Amminadab;
NUM|1|8|from Issachar, Nethanel son of Zuar;
NUM|1|9|from Zebulun, Eliab son of Helon;
NUM|1|10|from the sons of Joseph: from Ephraim, Elishama son of Ammihud; from Manasseh, Gamaliel son of Pedahzur;
NUM|1|11|from Benjamin, Abidan son of Gideoni;
NUM|1|12|from Dan, Ahiezer son of Ammishaddai;
NUM|1|13|from Asher, Pagiel son of Ocran;
NUM|1|14|from Gad, Eliasaph son of Deuel;
NUM|1|15|from Naphtali, Ahira son of Enan."
NUM|1|16|These were the men appointed from the community, the leaders of their ancestral tribes. They were the heads of the clans of Israel.
NUM|1|17|Moses and Aaron took these men whose names had been given,
NUM|1|18|and they called the whole community together on the first day of the second month. The people indicated their ancestry by their clans and families, and the men twenty years old or more were listed by name, one by one,
NUM|1|19|as the LORD commanded Moses. And so he counted them in the Desert of Sinai:
NUM|1|20|From the descendants of Reuben the firstborn son of Israel: All the men twenty years old or more who were able to serve in the army were listed by name, one by one, according to the records of their clans and families.
NUM|1|21|The number from the tribe of Reuben was 46,500.
NUM|1|22|From the descendants of Simeon: All the men twenty years old or more who were able to serve in the army were counted and listed by name, one by one, according to the records of their clans and families.
NUM|1|23|The number from the tribe of Simeon was 59,300.
NUM|1|24|From the descendants of Gad: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|25|The number from the tribe of Gad was 45,650.
NUM|1|26|From the descendants of Judah: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|27|The number from the tribe of Judah was 74,600.
NUM|1|28|From the descendants of Issachar: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|29|The number from the tribe of Issachar was 54,400.
NUM|1|30|From the descendants of Zebulun: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|31|The number from the tribe of Zebulun was 57,400.
NUM|1|32|From the sons of Joseph: From the descendants of Ephraim: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|33|The number from the tribe of Ephraim was 40,500.
NUM|1|34|From the descendants of Manasseh: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|35|The number from the tribe of Manasseh was 32,200.
NUM|1|36|From the descendants of Benjamin: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|37|The number from the tribe of Benjamin was 35,400.
NUM|1|38|From the descendants of Dan: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|39|The number from the tribe of Dan was 62,700.
NUM|1|40|From the descendants of Asher: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|41|The number from the tribe of Asher was 41,500.
NUM|1|42|From the descendants of Naphtali: All the men twenty years old or more who were able to serve in the army were listed by name, according to the records of their clans and families.
NUM|1|43|The number from the tribe of Naphtali was 53,400.
NUM|1|44|These were the men counted by Moses and Aaron and the twelve leaders of Israel, each one representing his family.
NUM|1|45|All the Israelites twenty years old or more who were able to serve in Israel's army were counted according to their families.
NUM|1|46|The total number was 603,550.
NUM|1|47|The families of the tribe of Levi, however, were not counted along with the others.
NUM|1|48|The LORD had said to Moses:
NUM|1|49|"You must not count the tribe of Levi or include them in the census of the other Israelites.
NUM|1|50|Instead, appoint the Levites to be in charge of the tabernacle of the Testimony-over all its furnishings and everything belonging to it. They are to carry the tabernacle and all its furnishings; they are to take care of it and encamp around it.
NUM|1|51|Whenever the tabernacle is to move, the Levites are to take it down, and whenever the tabernacle is to be set up, the Levites shall do it. Anyone else who goes near it shall be put to death.
NUM|1|52|The Israelites are to set up their tents by divisions, each man in his own camp under his own standard.
NUM|1|53|The Levites, however, are to set up their tents around the tabernacle of the Testimony so that wrath will not fall on the Israelite community. The Levites are to be responsible for the care of the tabernacle of the Testimony."
NUM|1|54|The Israelites did all this just as the LORD commanded Moses.
NUM|2|1|The LORD said to Moses and Aaron:
NUM|2|2|"The Israelites are to camp around the Tent of Meeting some distance from it, each man under his standard with the banners of his family."
NUM|2|3|On the east, toward the sunrise, the divisions of the camp of Judah are to encamp under their standard. The leader of the people of Judah is Nahshon son of Amminadab.
NUM|2|4|His division numbers 74,600.
NUM|2|5|The tribe of Issachar will camp next to them. The leader of the people of Issachar is Nethanel son of Zuar.
NUM|2|6|His division numbers 54,400.
NUM|2|7|The tribe of Zebulun will be next. The leader of the people of Zebulun is Eliab son of Helon.
NUM|2|8|His division numbers 57,400.
NUM|2|9|All the men assigned to the camp of Judah, according to their divisions, number 186,400. They will set out first.
NUM|2|10|On the south will be the divisions of the camp of Reuben under their standard. The leader of the people of Reuben is Elizur son of Shedeur.
NUM|2|11|His division numbers 46,500.
NUM|2|12|The tribe of Simeon will camp next to them. The leader of the people of Simeon is Shelumiel son of Zurishaddai.
NUM|2|13|His division numbers 59,300.
NUM|2|14|The tribe of Gad will be next. The leader of the people of Gad is Eliasaph son of Deuel.
NUM|2|15|His division numbers 45,650.
NUM|2|16|All the men assigned to the camp of Reuben, according to their divisions, number 151,450. They will set out second.
NUM|2|17|Then the Tent of Meeting and the camp of the Levites will set out in the middle of the camps. They will set out in the same order as they encamp, each in his own place under his standard.
NUM|2|18|On the west will be the divisions of the camp of Ephraim under their standard. The leader of the people of Ephraim is Elishama son of Ammihud.
NUM|2|19|His division numbers 40,500.
NUM|2|20|The tribe of Manasseh will be next to them. The leader of the people of Manasseh is Gamaliel son of Pedahzur.
NUM|2|21|His division numbers 32,200.
NUM|2|22|The tribe of Benjamin will be next. The leader of the people of Benjamin is Abidan son of Gideoni.
NUM|2|23|His division numbers 35,400.
NUM|2|24|All the men assigned to the camp of Ephraim, according to their divisions, number 108,100. They will set out third.
NUM|2|25|On the north will be the divisions of the camp of Dan, under their standard. The leader of the people of Dan is Ahiezer son of Ammishaddai.
NUM|2|26|His division numbers 62,700.
NUM|2|27|The tribe of Asher will camp next to them. The leader of the people of Asher is Pagiel son of Ocran.
NUM|2|28|His division numbers 41,500.
NUM|2|29|The tribe of Naphtali will be next. The leader of the people of Naphtali is Ahira son of Enan.
NUM|2|30|His division numbers 53,400.
NUM|2|31|All the men assigned to the camp of Dan number 157,600. They will set out last, under their standards.
NUM|2|32|These are the Israelites, counted according to their families. All those in the camps, by their divisions, number 603,550.
NUM|2|33|The Levites, however, were not counted along with the other Israelites, as the LORD commanded Moses.
NUM|2|34|So the Israelites did everything the LORD commanded Moses; that is the way they encamped under their standards, and that is the way they set out, each with his clan and family.
NUM|3|1|This is the account of the family of Aaron and Moses at the time the LORD talked with Moses on Mount Sinai.
NUM|3|2|The names of the sons of Aaron were Nadab the firstborn and Abihu, Eleazar and Ithamar.
NUM|3|3|Those were the names of Aaron's sons, the anointed priests, who were ordained to serve as priests.
NUM|3|4|Nadab and Abihu, however, fell dead before the LORD when they made an offering with unauthorized fire before him in the Desert of Sinai. They had no sons; so only Eleazar and Ithamar served as priests during the lifetime of their father Aaron.
NUM|3|5|The LORD said to Moses,
NUM|3|6|"Bring the tribe of Levi and present them to Aaron the priest to assist him.
NUM|3|7|They are to perform duties for him and for the whole community at the Tent of Meeting by doing the work of the tabernacle.
NUM|3|8|They are to take care of all the furnishings of the Tent of Meeting, fulfilling the obligations of the Israelites by doing the work of the tabernacle.
NUM|3|9|Give the Levites to Aaron and his sons; they are the Israelites who are to be given wholly to him.
NUM|3|10|Appoint Aaron and his sons to serve as priests; anyone else who approaches the sanctuary must be put to death."
NUM|3|11|The LORD also said to Moses,
NUM|3|12|"I have taken the Levites from among the Israelites in place of the first male offspring of every Israelite woman. The Levites are mine,
NUM|3|13|for all the firstborn are mine. When I struck down all the firstborn in Egypt, I set apart for myself every firstborn in Israel, whether man or animal. They are to be mine. I am the LORD."
NUM|3|14|The LORD said to Moses in the Desert of Sinai,
NUM|3|15|"Count the Levites by their families and clans. Count every male a month old or more."
NUM|3|16|So Moses counted them, as he was commanded by the word of the LORD.
NUM|3|17|These were the names of the sons of Levi: Gershon, Kohath and Merari.
NUM|3|18|These were the names of the Gershonite clans: Libni and Shimei.
NUM|3|19|The Kohathite clans: Amram, Izhar, Hebron and Uzziel.
NUM|3|20|The Merarite clans: Mahli and Mushi. These were the Levite clans, according to their families.
NUM|3|21|To Gershon belonged the clans of the Libnites and Shimeites; these were the Gershonite clans.
NUM|3|22|The number of all the males a month old or more who were counted was 7,500.
NUM|3|23|The Gershonite clans were to camp on the west, behind the tabernacle.
NUM|3|24|The leader of the families of the Gershonites was Eliasaph son of Lael.
NUM|3|25|At the Tent of Meeting the Gershonites were responsible for the care of the tabernacle and tent, its coverings, the curtain at the entrance to the Tent of Meeting,
NUM|3|26|the curtains of the courtyard, the curtain at the entrance to the courtyard surrounding the tabernacle and altar, and the ropes-and everything related to their use.
NUM|3|27|To Kohath belonged the clans of the Amramites, Izharites, Hebronites and Uzzielites; these were the Kohathite clans.
NUM|3|28|The number of all the males a month old or more was 8,600. The Kohathites were responsible for the care of the sanctuary.
NUM|3|29|The Kohathite clans were to camp on the south side of the tabernacle.
NUM|3|30|The leader of the families of the Kohathite clans was Elizaphan son of Uzziel.
NUM|3|31|They were responsible for the care of the ark, the table, the lampstand, the altars, the articles of the sanctuary used in ministering, the curtain, and everything related to their use.
NUM|3|32|The chief leader of the Levites was Eleazar son of Aaron, the priest. He was appointed over those who were responsible for the care of the sanctuary.
NUM|3|33|To Merari belonged the clans of the Mahlites and the Mushites; these were the Merarite clans.
NUM|3|34|The number of all the males a month old or more who were counted was 6,200.
NUM|3|35|The leader of the families of the Merarite clans was Zuriel son of Abihail; they were to camp on the north side of the tabernacle.
NUM|3|36|The Merarites were appointed to take care of the frames of the tabernacle, its crossbars, posts, bases, all its equipment, and everything related to their use,
NUM|3|37|as well as the posts of the surrounding courtyard with their bases, tent pegs and ropes.
NUM|3|38|Moses and Aaron and his sons were to camp to the east of the tabernacle, toward the sunrise, in front of the Tent of Meeting. They were responsible for the care of the sanctuary on behalf of the Israelites. Anyone else who approached the sanctuary was to be put to death.
NUM|3|39|The total number of Levites counted at the LORD's command by Moses and Aaron according to their clans, including every male a month old or more, was 22,000.
NUM|3|40|The LORD said to Moses, "Count all the firstborn Israelite males who are a month old or more and make a list of their names.
NUM|3|41|Take the Levites for me in place of all the firstborn of the Israelites, and the livestock of the Levites in place of all the firstborn of the livestock of the Israelites. I am the LORD."
NUM|3|42|So Moses counted all the firstborn of the Israelites, as the LORD commanded him.
NUM|3|43|The total number of firstborn males a month old or more, listed by name, was 22,273.
NUM|3|44|The LORD also said to Moses,
NUM|3|45|"Take the Levites in place of all the firstborn of Israel, and the livestock of the Levites in place of their livestock. The Levites are to be mine. I am the LORD.
NUM|3|46|To redeem the 273 firstborn Israelites who exceed the number of the Levites,
NUM|3|47|collect five shekels for each one, according to the sanctuary shekel, which weighs twenty gerahs.
NUM|3|48|Give the money for the redemption of the additional Israelites to Aaron and his sons."
NUM|3|49|So Moses collected the redemption money from those who exceeded the number redeemed by the Levites.
NUM|3|50|From the firstborn of the Israelites he collected silver weighing 1,365 shekels, according to the sanctuary shekel.
NUM|3|51|Moses gave the redemption money to Aaron and his sons, as he was commanded by the word of the LORD.
NUM|4|1|The LORD said to Moses and Aaron:
NUM|4|2|"Take a census of the Kohathite branch of the Levites by their clans and families.
NUM|4|3|Count all the men from thirty to fifty years of age who come to serve in the work in the Tent of Meeting.
NUM|4|4|"This is the work of the Kohathites in the Tent of Meeting: the care of the most holy things.
NUM|4|5|When the camp is to move, Aaron and his sons are to go in and take down the shielding curtain and cover the ark of the Testimony with it.
NUM|4|6|Then they are to cover this with hides of sea cows, spread a cloth of solid blue over that and put the poles in place.
NUM|4|7|"Over the table of the Presence they are to spread a blue cloth and put on it the plates, dishes and bowls, and the jars for drink offerings; the bread that is continually there is to remain on it.
NUM|4|8|Over these they are to spread a scarlet cloth, cover that with hides of sea cows and put its poles in place.
NUM|4|9|"They are to take a blue cloth and cover the lampstand that is for light, together with its lamps, its wick trimmers and trays, and all its jars for the oil used to supply it.
NUM|4|10|Then they are to wrap it and all its accessories in a covering of hides of sea cows and put it on a carrying frame.
NUM|4|11|"Over the gold altar they are to spread a blue cloth and cover that with hides of sea cows and put its poles in place.
NUM|4|12|"They are to take all the articles used for ministering in the sanctuary, wrap them in a blue cloth, cover that with hides of sea cows and put them on a carrying frame.
NUM|4|13|"They are to remove the ashes from the bronze altar and spread a purple cloth over it.
NUM|4|14|Then they are to place on it all the utensils used for ministering at the altar, including the firepans, meat forks, shovels and sprinkling bowls. Over it they are to spread a covering of hides of sea cows and put its poles in place.
NUM|4|15|"After Aaron and his sons have finished covering the holy furnishings and all the holy articles, and when the camp is ready to move, the Kohathites are to come to do the carrying. But they must not touch the holy things or they will die. The Kohathites are to carry those things that are in the Tent of Meeting.
NUM|4|16|"Eleazar son of Aaron, the priest, is to have charge of the oil for the light, the fragrant incense, the regular grain offering and the anointing oil. He is to be in charge of the entire tabernacle and everything in it, including its holy furnishings and articles."
NUM|4|17|The LORD said to Moses and Aaron,
NUM|4|18|"See that the Kohathite tribal clans are not cut off from the Levites.
NUM|4|19|So that they may live and not die when they come near the most holy things, do this for them: Aaron and his sons are to go into the sanctuary and assign to each man his work and what he is to carry.
NUM|4|20|But the Kohathites must not go in to look at the holy things, even for a moment, or they will die."
NUM|4|21|The LORD said to Moses,
NUM|4|22|"Take a census also of the Gershonites by their families and clans.
NUM|4|23|Count all the men from thirty to fifty years of age who come to serve in the work at the Tent of Meeting.
NUM|4|24|"This is the service of the Gershonite clans as they work and carry burdens:
NUM|4|25|They are to carry the curtains of the tabernacle, the Tent of Meeting, its covering and the outer covering of hides of sea cows, the curtains for the entrance to the Tent of Meeting,
NUM|4|26|the curtains of the courtyard surrounding the tabernacle and altar, the curtain for the entrance, the ropes and all the equipment used in its service. The Gershonites are to do all that needs to be done with these things.
NUM|4|27|All their service, whether carrying or doing other work, is to be done under the direction of Aaron and his sons. You shall assign to them as their responsibility all they are to carry.
NUM|4|28|This is the service of the Gershonite clans at the Tent of Meeting. Their duties are to be under the direction of Ithamar son of Aaron, the priest.
NUM|4|29|"Count the Merarites by their clans and families.
NUM|4|30|Count all the men from thirty to fifty years of age who come to serve in the work at the Tent of Meeting.
NUM|4|31|This is their duty as they perform service at the Tent of Meeting: to carry the frames of the tabernacle, its crossbars, posts and bases,
NUM|4|32|as well as the posts of the surrounding courtyard with their bases, tent pegs, ropes, all their equipment and everything related to their use. Assign to each man the specific things he is to carry.
NUM|4|33|This is the service of the Merarite clans as they work at the Tent of Meeting under the direction of Ithamar son of Aaron, the priest."
NUM|4|34|Moses, Aaron and the leaders of the community counted the Kohathites by their clans and families.
NUM|4|35|All the men from thirty to fifty years of age who came to serve in the work in the Tent of Meeting,
NUM|4|36|counted by clans, were 2,750.
NUM|4|37|This was the total of all those in the Kohathite clans who served in the Tent of Meeting. Moses and Aaron counted them according to the LORD's command through Moses.
NUM|4|38|The Gershonites were counted by their clans and families.
NUM|4|39|All the men from thirty to fifty years of age who came to serve in the work at the Tent of Meeting,
NUM|4|40|counted by their clans and families, were 2,630.
NUM|4|41|This was the total of those in the Gershonite clans who served at the Tent of Meeting. Moses and Aaron counted them according to the LORD's command.
NUM|4|42|The Merarites were counted by their clans and families.
NUM|4|43|All the men from thirty to fifty years of age who came to serve in the work at the Tent of Meeting,
NUM|4|44|counted by their clans, were 3,200.
NUM|4|45|This was the total of those in the Merarite clans. Moses and Aaron counted them according to the LORD's command through Moses.
NUM|4|46|So Moses, Aaron and the leaders of Israel counted all the Levites by their clans and families.
NUM|4|47|All the men from thirty to fifty years of age who came to do the work of serving and carrying the Tent of Meeting
NUM|4|48|numbered 8,580.
NUM|4|49|At the LORD's command through Moses, each was assigned his work and told what to carry. Thus they were counted, as the LORD commanded Moses.
NUM|5|1|The LORD said to Moses,
NUM|5|2|"Command the Israelites to send away from the camp anyone who has an infectious skin disease or a discharge of any kind, or who is ceremonially unclean because of a dead body.
NUM|5|3|Send away male and female alike; send them outside the camp so they will not defile their camp, where I dwell among them."
NUM|5|4|The Israelites did this; they sent them outside the camp. They did just as the LORD had instructed Moses.
NUM|5|5|The LORD said to Moses,
NUM|5|6|"Say to the Israelites: 'When a man or woman wrongs another in any way and so is unfaithful to the LORD, that person is guilty
NUM|5|7|and must confess the sin he has committed. He must make full restitution for his wrong, add one fifth to it and give it all to the person he has wronged.
NUM|5|8|But if that person has no close relative to whom restitution can be made for the wrong, the restitution belongs to the LORD and must be given to the priest, along with the ram with which atonement is made for him.
NUM|5|9|All the sacred contributions the Israelites bring to a priest will belong to him.
NUM|5|10|Each man's sacred gifts are his own, but what he gives to the priest will belong to the priest.'"
NUM|5|11|Then the LORD said to Moses,
NUM|5|12|"Speak to the Israelites and say to them: 'If a man's wife goes astray and is unfaithful to him
NUM|5|13|by sleeping with another man, and this is hidden from her husband and her impurity is undetected (since there is no witness against her and she has not been caught in the act),
NUM|5|14|and if feelings of jealousy come over her husband and he suspects his wife and she is impure-or if he is jealous and suspects her even though she is not impure-
NUM|5|15|then he is to take his wife to the priest. He must also take an offering of a tenth of an ephah of barley flour on her behalf. He must not pour oil on it or put incense on it, because it is a grain offering for jealousy, a reminder offering to draw attention to guilt.
NUM|5|16|"'The priest shall bring her and have her stand before the LORD.
NUM|5|17|Then he shall take some holy water in a clay jar and put some dust from the tabernacle floor into the water.
NUM|5|18|After the priest has had the woman stand before the LORD, he shall loosen her hair and place in her hands the reminder offering, the grain offering for jealousy, while he himself holds the bitter water that brings a curse.
NUM|5|19|Then the priest shall put the woman under oath and say to her, "If no other man has slept with you and you have not gone astray and become impure while married to your husband, may this bitter water that brings a curse not harm you.
NUM|5|20|But if you have gone astray while married to your husband and you have defiled yourself by sleeping with a man other than your husband"-
NUM|5|21|here the priest is to put the woman under this curse of the oath-"may the LORD cause your people to curse and denounce you when he causes your thigh to waste away and your abdomen to swell.
NUM|5|22|May this water that brings a curse enter your body so that your abdomen swells and your thigh wastes away.  'Then the woman is to say, "Amen. So be it."
NUM|5|23|"'The priest is to write these curses on a scroll and then wash them off into the bitter water.
NUM|5|24|He shall have the woman drink the bitter water that brings a curse, and this water will enter her and cause bitter suffering.
NUM|5|25|The priest is to take from her hands the grain offering for jealousy, wave it before the LORD and bring it to the altar.
NUM|5|26|The priest is then to take a handful of the grain offering as a memorial offering and burn it on the altar; after that, he is to have the woman drink the water.
NUM|5|27|If she has defiled herself and been unfaithful to her husband, then when she is made to drink the water that brings a curse, it will go into her and cause bitter suffering; her abdomen will swell and her thigh waste away, and she will become accursed among her people.
NUM|5|28|If, however, the woman has not defiled herself and is free from impurity, she will be cleared of guilt and will be able to have children.
NUM|5|29|"'This, then, is the law of jealousy when a woman goes astray and defiles herself while married to her husband,
NUM|5|30|or when feelings of jealousy come over a man because he suspects his wife. The priest is to have her stand before the LORD and is to apply this entire law to her.
NUM|5|31|The husband will be innocent of any wrongdoing, but the woman will bear the consequences of her sin.'"
NUM|6|1|The LORD said to Moses,
NUM|6|2|"Speak to the Israelites and say to them: 'If a man or woman wants to make a special vow, a vow of separation to the LORD as a Nazirite,
NUM|6|3|he must abstain from wine and other fermented drink and must not drink vinegar made from wine or from other fermented drink. He must not drink grape juice or eat grapes or raisins.
NUM|6|4|As long as he is a Nazirite, he must not eat anything that comes from the grapevine, not even the seeds or skins.
NUM|6|5|"'During the entire period of his vow of separation no razor may be used on his head. He must be holy until the period of his separation to the LORD is over; he must let the hair of his head grow long.
NUM|6|6|Throughout the period of his separation to the LORD he must not go near a dead body.
NUM|6|7|Even if his own father or mother or brother or sister dies, he must not make himself ceremonially unclean on account of them, because the symbol of his separation to God is on his head.
NUM|6|8|Throughout the period of his separation he is consecrated to the LORD.
NUM|6|9|"'If someone dies suddenly in his presence, thus defiling the hair he has dedicated, he must shave his head on the day of his cleansing-the seventh day.
NUM|6|10|Then on the eighth day he must bring two doves or two young pigeons to the priest at the entrance to the Tent of Meeting.
NUM|6|11|The priest is to offer one as a sin offering and the other as a burnt offering to make atonement for him because he sinned by being in the presence of the dead body. That same day he is to consecrate his head.
NUM|6|12|He must dedicate himself to the LORD for the period of his separation and must bring a year-old male lamb as a guilt offering. The previous days do not count, because he became defiled during his separation.
NUM|6|13|"'Now this is the law for the Nazirite when the period of his separation is over. He is to be brought to the entrance to the Tent of Meeting.
NUM|6|14|There he is to present his offerings to the LORD: a year-old male lamb without defect for a burnt offering, a year-old ewe lamb without defect for a sin offering, a ram without defect for a fellowship offering,
NUM|6|15|together with their grain offerings and drink offerings, and a basket of bread made without yeast-cakes made of fine flour mixed with oil, and wafers spread with oil.
NUM|6|16|"'The priest is to present them before the LORD and make the sin offering and the burnt offering.
NUM|6|17|He is to present the basket of unleavened bread and is to sacrifice the ram as a fellowship offering to the LORD, together with its grain offering and drink offering.
NUM|6|18|"'Then at the entrance to the Tent of Meeting, the Nazirite must shave off the hair that he dedicated. He is to take the hair and put it in the fire that is under the sacrifice of the fellowship offering.
NUM|6|19|"'After the Nazirite has shaved off the hair of his dedication, the priest is to place in his hands a boiled shoulder of the ram, and a cake and a wafer from the basket, both made without yeast.
NUM|6|20|The priest shall then wave them before the LORD as a wave offering; they are holy and belong to the priest, together with the breast that was waved and the thigh that was presented. After that, the Nazirite may drink wine.
NUM|6|21|"'This is the law of the Nazirite who vows his offering to the LORD in accordance with his separation, in addition to whatever else he can afford. He must fulfill the vow he has made, according to the law of the Nazirite.'"
NUM|6|22|The LORD said to Moses,
NUM|6|23|"Tell Aaron and his sons, 'This is how you are to bless the Israelites. Say to them:
NUM|6|24|"'"The LORD bless you and keep you;
NUM|6|25|the LORD make his face shine upon you and be gracious to you;
NUM|6|26|the LORD turn his face toward you and give you peace."'
NUM|6|27|"So they will put my name on the Israelites, and I will bless them."
NUM|7|1|When Moses finished setting up the tabernacle, he anointed it and consecrated it and all its furnishings. He also anointed and consecrated the altar and all its utensils.
NUM|7|2|Then the leaders of Israel, the heads of families who were the tribal leaders in charge of those who were counted, made offerings.
NUM|7|3|They brought as their gifts before the LORD six covered carts and twelve oxen-an ox from each leader and a cart from every two. These they presented before the tabernacle.
NUM|7|4|The LORD said to Moses,
NUM|7|5|"Accept these from them, that they may be used in the work at the Tent of Meeting. Give them to the Levites as each man's work requires."
NUM|7|6|So Moses took the carts and oxen and gave them to the Levites.
NUM|7|7|He gave two carts and four oxen to the Gershonites, as their work required,
NUM|7|8|and he gave four carts and eight oxen to the Merarites, as their work required. They were all under the direction of Ithamar son of Aaron, the priest.
NUM|7|9|But Moses did not give any to the Kohathites, because they were to carry on their shoulders the holy things, for which they were responsible.
NUM|7|10|When the altar was anointed, the leaders brought their offerings for its dedication and presented them before the altar.
NUM|7|11|For the LORD had said to Moses, "Each day one leader is to bring his offering for the dedication of the altar."
NUM|7|12|The one who brought his offering on the first day was Nahshon son of Amminadab of the tribe of Judah.
NUM|7|13|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|14|one gold dish weighing ten shekels, filled with incense;
NUM|7|15|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|16|one male goat for a sin offering;
NUM|7|17|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Nahshon son of Amminadab.
NUM|7|18|On the second day Nethanel son of Zuar, the leader of Issachar, brought his offering.
NUM|7|19|The offering he brought was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|20|one gold dish weighing ten shekels, filled with incense;
NUM|7|21|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|22|one male goat for a sin offering;
NUM|7|23|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Nethanel son of Zuar.
NUM|7|24|On the third day, Eliab son of Helon, the leader of the people of Zebulun, brought his offering.
NUM|7|25|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|26|one gold dish weighing ten shekels, filled with incense;
NUM|7|27|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|28|one male goat for a sin offering;
NUM|7|29|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Eliab son of Helon.
NUM|7|30|On the fourth day Elizur son of Shedeur, the leader of the people of Reuben, brought his offering.
NUM|7|31|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|32|one gold dish weighing ten shekels, filled with incense;
NUM|7|33|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|34|one male goat for a sin offering;
NUM|7|35|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Elizur son of Shedeur.
NUM|7|36|On the fifth day Shelumiel son of Zurishaddai, the leader of the people of Simeon, brought his offering.
NUM|7|37|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|38|one gold dish weighing ten shekels, filled with incense;
NUM|7|39|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|40|one male goat for a sin offering;
NUM|7|41|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Shelumiel son of Zurishaddai.
NUM|7|42|On the sixth day Eliasaph son of Deuel, the leader of the people of Gad, brought his offering.
NUM|7|43|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|44|one gold dish weighing ten shekels, filled with incense;
NUM|7|45|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|46|one male goat for a sin offering;
NUM|7|47|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Eliasaph son of Deuel.
NUM|7|48|On the seventh day Elishama son of Ammihud, the leader of the people of Ephraim, brought his offering.
NUM|7|49|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|50|one gold dish weighing ten shekels, filled with incense;
NUM|7|51|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|52|one male goat for a sin offering;
NUM|7|53|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Elishama son of Ammihud.
NUM|7|54|On the eighth day Gamaliel son of Pedahzur, the leader of the people of Manasseh, brought his offering.
NUM|7|55|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|56|one gold dish weighing ten shekels, filled with incense;
NUM|7|57|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|58|one male goat for a sin offering;
NUM|7|59|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Gamaliel son of Pedahzur.
NUM|7|60|On the ninth day Abidan son of Gideoni, the leader of the people of Benjamin, brought his offering.
NUM|7|61|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|62|one gold dish weighing ten shekels, filled with incense;
NUM|7|63|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|64|one male goat for a sin offering;
NUM|7|65|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Abidan son of Gideoni.
NUM|7|66|On the tenth day Ahiezer son of Ammishaddai, the leader of the people of Dan, brought his offering.
NUM|7|67|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|68|one gold dish weighing ten shekels, filled with incense;
NUM|7|69|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|70|one male goat for a sin offering;
NUM|7|71|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Ahiezer son of Ammishaddai.
NUM|7|72|On the eleventh day Pagiel son of Ocran, the leader of the people of Asher, brought his offering.
NUM|7|73|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|74|one gold dish weighing ten shekels, filled with incense;
NUM|7|75|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|76|one male goat for a sin offering;
NUM|7|77|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Pagiel son of Ocran.
NUM|7|78|On the twelfth day Ahira son of Enan, the leader of the people of Naphtali, brought his offering.
NUM|7|79|His offering was one silver plate weighing a hundred and thirty shekels, and one silver sprinkling bowl weighing seventy shekels, both according to the sanctuary shekel, each filled with fine flour mixed with oil as a grain offering;
NUM|7|80|one gold dish weighing ten shekels, filled with incense;
NUM|7|81|one young bull, one ram and one male lamb a year old, for a burnt offering;
NUM|7|82|one male goat for a sin offering;
NUM|7|83|and two oxen, five rams, five male goats and five male lambs a year old, to be sacrificed as a fellowship offering. This was the offering of Ahira son of Enan.
NUM|7|84|These were the offerings of the Israelite leaders for the dedication of the altar when it was anointed: twelve silver plates, twelve silver sprinkling bowls and twelve gold dishes.
NUM|7|85|Each silver plate weighed a hundred and thirty shekels, and each sprinkling bowl seventy shekels. Altogether, the silver dishes weighed two thousand four hundred shekels, according to the sanctuary shekel.
NUM|7|86|The twelve gold dishes filled with incense weighed ten shekels each, according to the sanctuary shekel. Altogether, the gold dishes weighed a hundred and twenty shekels.
NUM|7|87|The total number of animals for the burnt offering came to twelve young bulls, twelve rams and twelve male lambs a year old, together with their grain offering. Twelve male goats were used for the sin offering.
NUM|7|88|The total number of animals for the sacrifice of the fellowship offering came to twenty-four oxen, sixty rams, sixty male goats and sixty male lambs a year old. These were the offerings for the dedication of the altar after it was anointed.
NUM|7|89|When Moses entered the Tent of Meeting to speak with the LORD, he heard the voice speaking to him from between the two cherubim above the atonement cover on the ark of the Testimony. And he spoke with him.
NUM|8|1|The LORD said to Moses,
NUM|8|2|"Speak to Aaron and say to him, 'When you set up the seven lamps, they are to light the area in front of the lampstand.'"
NUM|8|3|Aaron did so; he set up the lamps so that they faced forward on the lampstand, just as the LORD commanded Moses.
NUM|8|4|This is how the lampstand was made: It was made of hammered gold-from its base to its blossoms. The lampstand was made exactly like the pattern the LORD had shown Moses.
NUM|8|5|The LORD said to Moses:
NUM|8|6|"Take the Levites from among the other Israelites and make them ceremonially clean.
NUM|8|7|To purify them, do this: Sprinkle the water of cleansing on them; then have them shave their whole bodies and wash their clothes, and so purify themselves.
NUM|8|8|Have them take a young bull with its grain offering of fine flour mixed with oil; then you are to take a second young bull for a sin offering.
NUM|8|9|Bring the Levites to the front of the Tent of Meeting and assemble the whole Israelite community.
NUM|8|10|You are to bring the Levites before the LORD, and the Israelites are to lay their hands on them.
NUM|8|11|Aaron is to present the Levites before the LORD as a wave offering from the Israelites, so that they may be ready to do the work of the LORD.
NUM|8|12|"After the Levites lay their hands on the heads of the bulls, use the one for a sin offering to the LORD and the other for a burnt offering, to make atonement for the Levites.
NUM|8|13|Have the Levites stand in front of Aaron and his sons and then present them as a wave offering to the LORD.
NUM|8|14|In this way you are to set the Levites apart from the other Israelites, and the Levites will be mine.
NUM|8|15|"After you have purified the Levites and presented them as a wave offering, they are to come to do their work at the Tent of Meeting.
NUM|8|16|They are the Israelites who are to be given wholly to me. I have taken them as my own in place of the firstborn, the first male offspring from every Israelite woman.
NUM|8|17|Every firstborn male in Israel, whether man or animal, is mine. When I struck down all the firstborn in Egypt, I set them apart for myself.
NUM|8|18|And I have taken the Levites in place of all the firstborn sons in Israel.
NUM|8|19|Of all the Israelites, I have given the Levites as gifts to Aaron and his sons to do the work at the Tent of Meeting on behalf of the Israelites and to make atonement for them so that no plague will strike the Israelites when they go near the sanctuary."
NUM|8|20|Moses, Aaron and the whole Israelite community did with the Levites just as the LORD commanded Moses.
NUM|8|21|The Levites purified themselves and washed their clothes. Then Aaron presented them as a wave offering before the LORD and made atonement for them to purify them.
NUM|8|22|After that, the Levites came to do their work at the Tent of Meeting under the supervision of Aaron and his sons. They did with the Levites just as the LORD commanded Moses.
NUM|8|23|The LORD said to Moses,
NUM|8|24|"This applies to the Levites: Men twenty-five years old or more shall come to take part in the work at the Tent of Meeting,
NUM|8|25|but at the age of fifty, they must retire from their regular service and work no longer.
NUM|8|26|They may assist their brothers in performing their duties at the Tent of Meeting, but they themselves must not do the work. This, then, is how you are to assign the responsibilities of the Levites."
NUM|9|1|The LORD spoke to Moses in the Desert of Sinai in the first month of the second year after they came out of Egypt. He said,
NUM|9|2|"Have the Israelites celebrate the Passover at the appointed time.
NUM|9|3|Celebrate it at the appointed time, at twilight on the fourteenth day of this month, in accordance with all its rules and regulations."
NUM|9|4|So Moses told the Israelites to celebrate the Passover,
NUM|9|5|and they did so in the Desert of Sinai at twilight on the fourteenth day of the first month. The Israelites did everything just as the LORD commanded Moses.
NUM|9|6|But some of them could not celebrate the Passover on that day because they were ceremonially unclean on account of a dead body. So they came to Moses and Aaron that same day
NUM|9|7|and said to Moses, "We have become unclean because of a dead body, but why should we be kept from presenting the LORD's offering with the other Israelites at the appointed time?"
NUM|9|8|Moses answered them, "Wait until I find out what the LORD commands concerning you."
NUM|9|9|Then the LORD said to Moses,
NUM|9|10|"Tell the Israelites: 'When any of you or your descendants are unclean because of a dead body or are away on a journey, they may still celebrate the LORD's Passover.
NUM|9|11|They are to celebrate it on the fourteenth day of the second month at twilight. They are to eat the lamb, together with unleavened bread and bitter herbs.
NUM|9|12|They must not leave any of it till morning or break any of its bones. When they celebrate the Passover, they must follow all the regulations.
NUM|9|13|But if a man who is ceremonially clean and not on a journey fails to celebrate the Passover, that person must be cut off from his people because he did not present the LORD's offering at the appointed time. That man will bear the consequences of his sin.
NUM|9|14|"'An alien living among you who wants to celebrate the LORD's Passover must do so in accordance with its rules and regulations. You must have the same regulations for the alien and the native-born.'"
NUM|9|15|On the day the tabernacle, the Tent of the Testimony, was set up, the cloud covered it. From evening till morning the cloud above the tabernacle looked like fire.
NUM|9|16|That is how it continued to be; the cloud covered it, and at night it looked like fire.
NUM|9|17|Whenever the cloud lifted from above the Tent, the Israelites set out; wherever the cloud settled, the Israelites encamped.
NUM|9|18|At the LORD's command the Israelites set out, and at his command they encamped. As long as the cloud stayed over the tabernacle, they remained in camp.
NUM|9|19|When the cloud remained over the tabernacle a long time, the Israelites obeyed the LORD's order and did not set out.
NUM|9|20|Sometimes the cloud was over the tabernacle only a few days; at the LORD's command they would encamp, and then at his command they would set out.
NUM|9|21|Sometimes the cloud stayed only from evening till morning, and when it lifted in the morning, they set out. Whether by day or by night, whenever the cloud lifted, they set out.
NUM|9|22|Whether the cloud stayed over the tabernacle for two days or a month or a year, the Israelites would remain in camp and not set out; but when it lifted, they would set out.
NUM|9|23|At the LORD's command they encamped, and at the LORD's command they set out. They obeyed the LORD's order, in accordance with his command through Moses.
NUM|10|1|The LORD said to Moses:
NUM|10|2|"Make two trumpets of hammered silver, and use them for calling the community together and for having the camps set out.
NUM|10|3|When both are sounded, the whole community is to assemble before you at the entrance to the Tent of Meeting.
NUM|10|4|If only one is sounded, the leaders-the heads of the clans of Israel-are to assemble before you.
NUM|10|5|When a trumpet blast is sounded, the tribes camping on the east are to set out.
NUM|10|6|At the sounding of a second blast, the camps on the south are to set out. The blast will be the signal for setting out.
NUM|10|7|To gather the assembly, blow the trumpets, but not with the same signal.
NUM|10|8|"The sons of Aaron, the priests, are to blow the trumpets. This is to be a lasting ordinance for you and the generations to come.
NUM|10|9|When you go into battle in your own land against an enemy who is oppressing you, sound a blast on the trumpets. Then you will be remembered by the LORD your God and rescued from your enemies.
NUM|10|10|Also at your times of rejoicing-your appointed feasts and New Moon festivals-you are to sound the trumpets over your burnt offerings and fellowship offerings, and they will be a memorial for you before your God. I am the LORD your God."
NUM|10|11|On the twentieth day of the second month of the second year, the cloud lifted from above the tabernacle of the Testimony.
NUM|10|12|Then the Israelites set out from the Desert of Sinai and traveled from place to place until the cloud came to rest in the Desert of Paran.
NUM|10|13|They set out, this first time, at the LORD's command through Moses.
NUM|10|14|The divisions of the camp of Judah went first, under their standard. Nahshon son of Amminadab was in command.
NUM|10|15|Nethanel son of Zuar was over the division of the tribe of Issachar,
NUM|10|16|and Eliab son of Helon was over the division of the tribe of Zebulun.
NUM|10|17|Then the tabernacle was taken down, and the Gershonites and Merarites, who carried it, set out.
NUM|10|18|The divisions of the camp of Reuben went next, under their standard. Elizur son of Shedeur was in command.
NUM|10|19|Shelumiel son of Zurishaddai was over the division of the tribe of Simeon,
NUM|10|20|and Eliasaph son of Deuel was over the division of the tribe of Gad.
NUM|10|21|Then the Kohathites set out, carrying the holy things. The tabernacle was to be set up before they arrived.
NUM|10|22|The divisions of the camp of Ephraim went next, under their standard. Elishama son of Ammihud was in command.
NUM|10|23|Gamaliel son of Pedahzur was over the division of the tribe of Manasseh,
NUM|10|24|and Abidan son of Gideoni was over the division of the tribe of Benjamin.
NUM|10|25|Finally, as the rear guard for all the units, the divisions of the camp of Dan set out, under their standard. Ahiezer son of Ammishaddai was in command.
NUM|10|26|Pagiel son of Ocran was over the division of the tribe of Asher,
NUM|10|27|and Ahira son of Enan was over the division of the tribe of Naphtali.
NUM|10|28|This was the order of march for the Israelite divisions as they set out.
NUM|10|29|Now Moses said to Hobab son of Reuel the Midianite, Moses' father-in-law, "We are setting out for the place about which the LORD said, 'I will give it to you.' Come with us and we will treat you well, for the LORD has promised good things to Israel."
NUM|10|30|He answered, "No, I will not go; I am going back to my own land and my own people."
NUM|10|31|But Moses said, "Please do not leave us. You know where we should camp in the desert, and you can be our eyes.
NUM|10|32|If you come with us, we will share with you whatever good things the LORD gives us."
NUM|10|33|So they set out from the mountain of the LORD and traveled for three days. The ark of the covenant of the LORD went before them during those three days to find them a place to rest.
NUM|10|34|The cloud of the LORD was over them by day when they set out from the camp.
NUM|10|35|Whenever the ark set out, Moses said, "Rise up, O LORD! May your enemies be scattered; may your foes flee before you."
NUM|10|36|Whenever it came to rest, he said, "Return, O LORD, to the countless thousands of Israel."
NUM|11|1|Now the people complained about their hardships in the hearing of the LORD, and when he heard them his anger was aroused. Then fire from the LORD burned among them and consumed some of the outskirts of the camp.
NUM|11|2|When the people cried out to Moses, he prayed to the LORD and the fire died down.
NUM|11|3|So that place was called Taberah, because fire from the LORD had burned among them. Quail From the LORD
NUM|11|4|The rabble with them began to crave other food, and again the Israelites started wailing and said, "If only we had meat to eat!
NUM|11|5|We remember the fish we ate in Egypt at no cost-also the cucumbers, melons, leeks, onions and garlic.
NUM|11|6|But now we have lost our appetite; we never see anything but this manna!"
NUM|11|7|The manna was like coriander seed and looked like resin.
NUM|11|8|The people went around gathering it, and then ground it in a handmill or crushed it in a mortar. They cooked it in a pot or made it into cakes. And it tasted like something made with olive oil.
NUM|11|9|When the dew settled on the camp at night, the manna also came down.
NUM|11|10|Moses heard the people of every family wailing, each at the entrance to his tent. The LORD became exceedingly angry, and Moses was troubled.
NUM|11|11|He asked the LORD, "Why have you brought this trouble on your servant? What have I done to displease you that you put the burden of all these people on me?
NUM|11|12|Did I conceive all these people? Did I give them birth? Why do you tell me to carry them in my arms, as a nurse carries an infant, to the land you promised on oath to their forefathers?
NUM|11|13|Where can I get meat for all these people? They keep wailing to me, 'Give us meat to eat!'
NUM|11|14|I cannot carry all these people by myself; the burden is too heavy for me.
NUM|11|15|If this is how you are going to treat me, put me to death right now-if I have found favor in your eyes-and do not let me face my own ruin."
NUM|11|16|The LORD said to Moses: "Bring me seventy of Israel's elders who are known to you as leaders and officials among the people. Have them come to the Tent of Meeting, that they may stand there with you.
NUM|11|17|I will come down and speak with you there, and I will take of the Spirit that is on you and put the Spirit on them. They will help you carry the burden of the people so that you will not have to carry it alone.
NUM|11|18|"Tell the people: 'Consecrate yourselves in preparation for tomorrow, when you will eat meat. The LORD heard you when you wailed, "If only we had meat to eat! We were better off in Egypt!" Now the LORD will give you meat, and you will eat it.
NUM|11|19|You will not eat it for just one day, or two days, or five, ten or twenty days,
NUM|11|20|but for a whole month-until it comes out of your nostrils and you loathe it-because you have rejected the LORD, who is among you, and have wailed before him, saying, "Why did we ever leave Egypt?"'"
NUM|11|21|But Moses said, "Here I am among six hundred thousand men on foot, and you say, 'I will give them meat to eat for a whole month!'
NUM|11|22|Would they have enough if flocks and herds were slaughtered for them? Would they have enough if all the fish in the sea were caught for them?"
NUM|11|23|The LORD answered Moses, "Is the LORD's arm too short? You will now see whether or not what I say will come true for you."
NUM|11|24|So Moses went out and told the people what the LORD had said. He brought together seventy of their elders and had them stand around the Tent.
NUM|11|25|Then the LORD came down in the cloud and spoke with him, and he took of the Spirit that was on him and put the Spirit on the seventy elders. When the Spirit rested on them, they prophesied, but they did not do so again.
NUM|11|26|However, two men, whose names were Eldad and Medad, had remained in the camp. They were listed among the elders, but did not go out to the Tent. Yet the Spirit also rested on them, and they prophesied in the camp.
NUM|11|27|A young man ran and told Moses, "Eldad and Medad are prophesying in the camp."
NUM|11|28|Joshua son of Nun, who had been Moses' aide since youth, spoke up and said, "Moses, my lord, stop them!"
NUM|11|29|But Moses replied, "Are you jealous for my sake? I wish that all the LORD's people were prophets and that the LORD would put his Spirit on them!"
NUM|11|30|Then Moses and the elders of Israel returned to the camp.
NUM|11|31|Now a wind went out from the LORD and drove quail in from the sea. It brought them down all around the camp to about three feet above the ground, as far as a day's walk in any direction.
NUM|11|32|All that day and night and all the next day the people went out and gathered quail. No one gathered less than ten homers. Then they spread them out all around the camp.
NUM|11|33|But while the meat was still between their teeth and before it could be consumed, the anger of the LORD burned against the people, and he struck them with a severe plague.
NUM|11|34|Therefore the place was named Kibroth Hattaavah, because there they buried the people who had craved other food.
NUM|11|35|From Kibroth Hattaavah the people traveled to Hazeroth and stayed there.
NUM|12|1|Miriam and Aaron began to talk against Moses because of his Cushite wife, for he had married a Cushite.
NUM|12|2|"Has the LORD spoken only through Moses?" they asked. "Hasn't he also spoken through us?" And the LORD heard this.
NUM|12|3|(Now Moses was a very humble man, more humble than anyone else on the face of the earth.)
NUM|12|4|At once the LORD said to Moses, Aaron and Miriam, "Come out to the Tent of Meeting, all three of you." So the three of them came out.
NUM|12|5|Then the LORD came down in a pillar of cloud; he stood at the entrance to the Tent and summoned Aaron and Miriam. When both of them stepped forward,
NUM|12|6|he said, "Listen to my words: "When a prophet of the LORD is among you, I reveal myself to him in visions, I speak to him in dreams.
NUM|12|7|But this is not true of my servant Moses; he is faithful in all my house.
NUM|12|8|With him I speak face to face, clearly and not in riddles; he sees the form of the LORD. Why then were you not afraid to speak against my servant Moses?"
NUM|12|9|The anger of the LORD burned against them, and he left them.
NUM|12|10|When the cloud lifted from above the Tent, there stood Miriam-leprous, like snow. Aaron turned toward her and saw that she had leprosy;
NUM|12|11|and he said to Moses, "Please, my lord, do not hold against us the sin we have so foolishly committed.
NUM|12|12|Do not let her be like a stillborn infant coming from its mother's womb with its flesh half eaten away."
NUM|12|13|So Moses cried out to the LORD, "O God, please heal her!"
NUM|12|14|The LORD replied to Moses, "If her father had spit in her face, would she not have been in disgrace for seven days? Confine her outside the camp for seven days; after that she can be brought back."
NUM|12|15|So Miriam was confined outside the camp for seven days, and the people did not move on till she was brought back.
NUM|12|16|After that, the people left Hazeroth and encamped in the Desert of Paran.
NUM|13|1|The LORD said to Moses,
NUM|13|2|"Send some men to explore the land of Canaan, which I am giving to the Israelites. From each ancestral tribe send one of its leaders."
NUM|13|3|So at the LORD's command Moses sent them out from the Desert of Paran. All of them were leaders of the Israelites.
NUM|13|4|These are their names: from the tribe of Reuben, Shammua son of Zaccur;
NUM|13|5|from the tribe of Simeon, Shaphat son of Hori;
NUM|13|6|from the tribe of Judah, Caleb son of Jephunneh;
NUM|13|7|from the tribe of Issachar, Igal son of Joseph;
NUM|13|8|from the tribe of Ephraim, Hoshea son of Nun;
NUM|13|9|from the tribe of Benjamin, Palti son of Raphu;
NUM|13|10|from the tribe of Zebulun, Gaddiel son of Sodi;
NUM|13|11|from the tribe of Manasseh (a tribe of Joseph), Gaddi son of Susi;
NUM|13|12|from the tribe of Dan, Ammiel son of Gemalli;
NUM|13|13|from the tribe of Asher, Sethur son of Michael;
NUM|13|14|from the tribe of Naphtali, Nahbi son of Vophsi;
NUM|13|15|from the tribe of Gad, Geuel son of Maki.
NUM|13|16|These are the names of the men Moses sent to explore the land. (Moses gave Hoshea son of Nun the name Joshua.)
NUM|13|17|When Moses sent them to explore Canaan, he said, "Go up through the Negev and on into the hill country.
NUM|13|18|See what the land is like and whether the people who live there are strong or weak, few or many.
NUM|13|19|What kind of land do they live in? Is it good or bad? What kind of towns do they live in? Are they unwalled or fortified?
NUM|13|20|How is the soil? Is it fertile or poor? Are there trees on it or not? Do your best to bring back some of the fruit of the land." (It was the season for the first ripe grapes.)
NUM|13|21|So they went up and explored the land from the Desert of Zin as far as Rehob, toward Lebo Hamath.
NUM|13|22|They went up through the Negev and came to Hebron, where Ahiman, Sheshai and Talmai, the descendants of Anak, lived. (Hebron had been built seven years before Zoan in Egypt.)
NUM|13|23|When they reached the Valley of Eshcol, they cut off a branch bearing a single cluster of grapes. Two of them carried it on a pole between them, along with some pomegranates and figs.
NUM|13|24|That place was called the Valley of Eshcol because of the cluster of grapes the Israelites cut off there.
NUM|13|25|At the end of forty days they returned from exploring the land.
NUM|13|26|They came back to Moses and Aaron and the whole Israelite community at Kadesh in the Desert of Paran. There they reported to them and to the whole assembly and showed them the fruit of the land.
NUM|13|27|They gave Moses this account: "We went into the land to which you sent us, and it does flow with milk and honey! Here is its fruit.
NUM|13|28|But the people who live there are powerful, and the cities are fortified and very large. We even saw descendants of Anak there.
NUM|13|29|The Amalekites live in the Negev; the Hittites, Jebusites and Amorites live in the hill country; and the Canaanites live near the sea and along the Jordan."
NUM|13|30|Then Caleb silenced the people before Moses and said, "We should go up and take possession of the land, for we can certainly do it."
NUM|13|31|But the men who had gone up with him said, "We can't attack those people; they are stronger than we are."
NUM|13|32|And they spread among the Israelites a bad report about the land they had explored. They said, "The land we explored devours those living in it. All the people we saw there are of great size.
NUM|13|33|We saw the Nephilim there (the descendants of Anak come from the Nephilim). We seemed like grasshoppers in our own eyes, and we looked the same to them."
NUM|14|1|That night all the people of the community raised their voices and wept aloud.
NUM|14|2|All the Israelites grumbled against Moses and Aaron, and the whole assembly said to them, "If only we had died in Egypt! Or in this desert!
NUM|14|3|Why is the LORD bringing us to this land only to let us fall by the sword? Our wives and children will be taken as plunder. Wouldn't it be better for us to go back to Egypt?"
NUM|14|4|And they said to each other, "We should choose a leader and go back to Egypt."
NUM|14|5|Then Moses and Aaron fell facedown in front of the whole Israelite assembly gathered there.
NUM|14|6|Joshua son of Nun and Caleb son of Jephunneh, who were among those who had explored the land, tore their clothes
NUM|14|7|and said to the entire Israelite assembly, "The land we passed through and explored is exceedingly good.
NUM|14|8|If the LORD is pleased with us, he will lead us into that land, a land flowing with milk and honey, and will give it to us.
NUM|14|9|Only do not rebel against the LORD. And do not be afraid of the people of the land, because we will swallow them up. Their protection is gone, but the LORD is with us. Do not be afraid of them."
NUM|14|10|But the whole assembly talked about stoning them. Then the glory of the LORD appeared at the Tent of Meeting to all the Israelites.
NUM|14|11|The LORD said to Moses, "How long will these people treat me with contempt? How long will they refuse to believe in me, in spite of all the miraculous signs I have performed among them?
NUM|14|12|I will strike them down with a plague and destroy them, but I will make you into a nation greater and stronger than they."
NUM|14|13|Moses said to the LORD, "Then the Egyptians will hear about it! By your power you brought these people up from among them.
NUM|14|14|And they will tell the inhabitants of this land about it. They have already heard that you, O LORD, are with these people and that you, O LORD, have been seen face to face, that your cloud stays over them, and that you go before them in a pillar of cloud by day and a pillar of fire by night.
NUM|14|15|If you put these people to death all at one time, the nations who have heard this report about you will say,
NUM|14|16|'The LORD was not able to bring these people into the land he promised them on oath; so he slaughtered them in the desert.'
NUM|14|17|"Now may the Lord's strength be displayed, just as you have declared:
NUM|14|18|'The LORD is slow to anger, abounding in love and forgiving sin and rebellion. Yet he does not leave the guilty unpunished; he punishes the children for the sin of the fathers to the third and fourth generation.'
NUM|14|19|In accordance with your great love, forgive the sin of these people, just as you have pardoned them from the time they left Egypt until now."
NUM|14|20|The LORD replied, "I have forgiven them, as you asked.
NUM|14|21|Nevertheless, as surely as I live and as surely as the glory of the LORD fills the whole earth,
NUM|14|22|not one of the men who saw my glory and the miraculous signs I performed in Egypt and in the desert but who disobeyed me and tested me ten times-
NUM|14|23|not one of them will ever see the land I promised on oath to their forefathers. No one who has treated me with contempt will ever see it.
NUM|14|24|But because my servant Caleb has a different spirit and follows me wholeheartedly, I will bring him into the land he went to, and his descendants will inherit it.
NUM|14|25|Since the Amalekites and Canaanites are living in the valleys, turn back tomorrow and set out toward the desert along the route to the Red Sea. "
NUM|14|26|The LORD said to Moses and Aaron:
NUM|14|27|"How long will this wicked community grumble against me? I have heard the complaints of these grumbling Israelites.
NUM|14|28|So tell them, 'As surely as I live, declares the LORD, I will do to you the very things I heard you say:
NUM|14|29|In this desert your bodies will fall-every one of you twenty years old or more who was counted in the census and who has grumbled against me.
NUM|14|30|Not one of you will enter the land I swore with uplifted hand to make your home, except Caleb son of Jephunneh and Joshua son of Nun.
NUM|14|31|As for your children that you said would be taken as plunder, I will bring them in to enjoy the land you have rejected.
NUM|14|32|But you-your bodies will fall in this desert.
NUM|14|33|Your children will be shepherds here for forty years, suffering for your unfaithfulness, until the last of your bodies lies in the desert.
NUM|14|34|For forty years-one year for each of the forty days you explored the land-you will suffer for your sins and know what it is like to have me against you.'
NUM|14|35|I, the LORD, have spoken, and I will surely do these things to this whole wicked community, which has banded together against me. They will meet their end in this desert; here they will die."
NUM|14|36|So the men Moses had sent to explore the land, who returned and made the whole community grumble against him by spreading a bad report about it-
NUM|14|37|these men responsible for spreading the bad report about the land were struck down and died of a plague before the LORD.
NUM|14|38|Of the men who went to explore the land, only Joshua son of Nun and Caleb son of Jephunneh survived.
NUM|14|39|When Moses reported this to all the Israelites, they mourned bitterly.
NUM|14|40|Early the next morning they went up toward the high hill country. "We have sinned," they said. "We will go up to the place the LORD promised."
NUM|14|41|But Moses said, "Why are you disobeying the LORD's command? This will not succeed!
NUM|14|42|Do not go up, because the LORD is not with you. You will be defeated by your enemies,
NUM|14|43|for the Amalekites and Canaanites will face you there. Because you have turned away from the LORD, he will not be with you and you will fall by the sword."
NUM|14|44|Nevertheless, in their presumption they went up toward the high hill country, though neither Moses nor the ark of the LORD's covenant moved from the camp.
NUM|14|45|Then the Amalekites and Canaanites who lived in that hill country came down and attacked them and beat them down all the way to Hormah.
NUM|15|1|The LORD said to Moses,
NUM|15|2|"Speak to the Israelites and say to them: 'After you enter the land I am giving you as a home
NUM|15|3|and you present to the LORD offerings made by fire, from the herd or the flock, as an aroma pleasing to the LORD -whether burnt offerings or sacrifices, for special vows or freewill offerings or festival offerings-
NUM|15|4|then the one who brings his offering shall present to the LORD a grain offering of a tenth of an ephah of fine flour mixed with a quarter of a hin of oil.
NUM|15|5|With each lamb for the burnt offering or the sacrifice, prepare a quarter of a hin of wine as a drink offering.
NUM|15|6|"'With a ram prepare a grain offering of two-tenths of an ephah of fine flour mixed with a third of a hin of oil,
NUM|15|7|and a third of a hin of wine as a drink offering. Offer it as an aroma pleasing to the LORD.
NUM|15|8|"'When you prepare a young bull as a burnt offering or sacrifice, for a special vow or a fellowship offering to the LORD,
NUM|15|9|bring with the bull a grain offering of three-tenths of an ephah of fine flour mixed with half a hin of oil.
NUM|15|10|Also bring half a hin of wine as a drink offering. It will be an offering made by fire, an aroma pleasing to the LORD.
NUM|15|11|Each bull or ram, each lamb or young goat, is to be prepared in this manner.
NUM|15|12|Do this for each one, for as many as you prepare.
NUM|15|13|"'Everyone who is native-born must do these things in this way when he brings an offering made by fire as an aroma pleasing to the LORD.
NUM|15|14|For the generations to come, whenever an alien or anyone else living among you presents an offering made by fire as an aroma pleasing to the LORD, he must do exactly as you do.
NUM|15|15|The community is to have the same rules for you and for the alien living among you; this is a lasting ordinance for the generations to come. You and the alien shall be the same before the LORD:
NUM|15|16|The same laws and regulations will apply both to you and to the alien living among you.'"
NUM|15|17|The LORD said to Moses,
NUM|15|18|"Speak to the Israelites and say to them: 'When you enter the land to which I am taking you
NUM|15|19|and you eat the food of the land, present a portion as an offering to the LORD.
NUM|15|20|Present a cake from the first of your ground meal and present it as an offering from the threshing floor.
NUM|15|21|Throughout the generations to come you are to give this offering to the LORD from the first of your ground meal.
NUM|15|22|"'Now if you unintentionally fail to keep any of these commands the LORD gave Moses-
NUM|15|23|any of the LORD's commands to you through him, from the day the LORD gave them and continuing through the generations to come-
NUM|15|24|and if this is done unintentionally without the community being aware of it, then the whole community is to offer a young bull for a burnt offering as an aroma pleasing to the LORD, along with its prescribed grain offering and drink offering, and a male goat for a sin offering.
NUM|15|25|The priest is to make atonement for the whole Israelite community, and they will be forgiven, for it was not intentional and they have brought to the LORD for their wrong an offering made by fire and a sin offering.
NUM|15|26|The whole Israelite community and the aliens living among them will be forgiven, because all the people were involved in the unintentional wrong.
NUM|15|27|"'But if just one person sins unintentionally, he must bring a year-old female goat for a sin offering.
NUM|15|28|The priest is to make atonement before the LORD for the one who erred by sinning unintentionally, and when atonement has been made for him, he will be forgiven.
NUM|15|29|One and the same law applies to everyone who sins unintentionally, whether he is a native-born Israelite or an alien.
NUM|15|30|"'But anyone who sins defiantly, whether native-born or alien, blasphemes the LORD, and that person must be cut off from his people.
NUM|15|31|Because he has despised the LORD's word and broken his commands, that person must surely be cut off; his guilt remains on him.'"
NUM|15|32|While the Israelites were in the desert, a man was found gathering wood on the Sabbath day.
NUM|15|33|Those who found him gathering wood brought him to Moses and Aaron and the whole assembly,
NUM|15|34|and they kept him in custody, because it was not clear what should be done to him.
NUM|15|35|Then the LORD said to Moses, "The man must die. The whole assembly must stone him outside the camp."
NUM|15|36|So the assembly took him outside the camp and stoned him to death, as the LORD commanded Moses.
NUM|15|37|The LORD said to Moses,
NUM|15|38|"Speak to the Israelites and say to them: 'Throughout the generations to come you are to make tassels on the corners of your garments, with a blue cord on each tassel.
NUM|15|39|You will have these tassels to look at and so you will remember all the commands of the LORD, that you may obey them and not prostitute yourselves by going after the lusts of your own hearts and eyes.
NUM|15|40|Then you will remember to obey all my commands and will be consecrated to your God.
NUM|15|41|I am the LORD your God, who brought you out of Egypt to be your God. I am the LORD your God.'"
NUM|16|1|Korah son of Izhar, the son of Kohath, the son of Levi, and certain Reubenites-Dathan and Abiram, sons of Eliab, and On son of Peleth-became insolent
NUM|16|2|and rose up against Moses. With them were 250 Israelite men, well-known community leaders who had been appointed members of the council.
NUM|16|3|They came as a group to oppose Moses and Aaron and said to them, "You have gone too far! The whole community is holy, every one of them, and the LORD is with them. Why then do you set yourselves above the LORD's assembly?"
NUM|16|4|When Moses heard this, he fell facedown.
NUM|16|5|Then he said to Korah and all his followers: "In the morning the LORD will show who belongs to him and who is holy, and he will have that person come near him. The man he chooses he will cause to come near him.
NUM|16|6|You, Korah, and all your followers are to do this: Take censers
NUM|16|7|and tomorrow put fire and incense in them before the LORD. The man the LORD chooses will be the one who is holy. You Levites have gone too far!"
NUM|16|8|Moses also said to Korah, "Now listen, you Levites!
NUM|16|9|Isn't it enough for you that the God of Israel has separated you from the rest of the Israelite community and brought you near himself to do the work at the LORD's tabernacle and to stand before the community and minister to them?
NUM|16|10|He has brought you and all your fellow Levites near himself, but now you are trying to get the priesthood too.
NUM|16|11|It is against the LORD that you and all your followers have banded together. Who is Aaron that you should grumble against him?"
NUM|16|12|Then Moses summoned Dathan and Abiram, the sons of Eliab. But they said, "We will not come!
NUM|16|13|Isn't it enough that you have brought us up out of a land flowing with milk and honey to kill us in the desert? And now you also want to lord it over us?
NUM|16|14|Moreover, you haven't brought us into a land flowing with milk and honey or given us an inheritance of fields and vineyards. Will you gouge out the eyes of these men? No, we will not come!"
NUM|16|15|Then Moses became very angry and said to the LORD, "Do not accept their offering. I have not taken so much as a donkey from them, nor have I wronged any of them."
NUM|16|16|Moses said to Korah, "You and all your followers are to appear before the LORD tomorrow-you and they and Aaron.
NUM|16|17|Each man is to take his censer and put incense in it-250 censers in all-and present it before the LORD. You and Aaron are to present your censers also."
NUM|16|18|So each man took his censer, put fire and incense in it, and stood with Moses and Aaron at the entrance to the Tent of Meeting.
NUM|16|19|When Korah had gathered all his followers in opposition to them at the entrance to the Tent of Meeting, the glory of the LORD appeared to the entire assembly.
NUM|16|20|The LORD said to Moses and Aaron,
NUM|16|21|"Separate yourselves from this assembly so I can put an end to them at once."
NUM|16|22|But Moses and Aaron fell facedown and cried out, "O God, God of the spirits of all mankind, will you be angry with the entire assembly when only one man sins?"
NUM|16|23|Then the LORD said to Moses,
NUM|16|24|"Say to the assembly, 'Move away from the tents of Korah, Dathan and Abiram.'"
NUM|16|25|Moses got up and went to Dathan and Abiram, and the elders of Israel followed him.
NUM|16|26|He warned the assembly, "Move back from the tents of these wicked men! Do not touch anything belonging to them, or you will be swept away because of all their sins."
NUM|16|27|So they moved away from the tents of Korah, Dathan and Abiram. Dathan and Abiram had come out and were standing with their wives, children and little ones at the entrances to their tents.
NUM|16|28|Then Moses said, "This is how you will know that the LORD has sent me to do all these things and that it was not my idea:
NUM|16|29|If these men die a natural death and experience only what usually happens to men, then the LORD has not sent me.
NUM|16|30|But if the LORD brings about something totally new, and the earth opens its mouth and swallows them, with everything that belongs to them, and they go down alive into the grave, then you will know that these men have treated the LORD with contempt."
NUM|16|31|As soon as he finished saying all this, the ground under them split apart
NUM|16|32|and the earth opened its mouth and swallowed them, with their households and all Korah's men and all their possessions.
NUM|16|33|They went down alive into the grave, with everything they owned; the earth closed over them, and they perished and were gone from the community.
NUM|16|34|At their cries, all the Israelites around them fled, shouting, "The earth is going to swallow us too!"
NUM|16|35|And fire came out from the LORD and consumed the 250 men who were offering the incense.
NUM|16|36|The LORD said to Moses,
NUM|16|37|"Tell Eleazar son of Aaron, the priest, to take the censers out of the smoldering remains and scatter the coals some distance away, for the censers are holy-
NUM|16|38|the censers of the men who sinned at the cost of their lives. Hammer the censers into sheets to overlay the altar, for they were presented before the LORD and have become holy. Let them be a sign to the Israelites."
NUM|16|39|So Eleazar the priest collected the bronze censers brought by those who had been burned up, and he had them hammered out to overlay the altar,
NUM|16|40|as the LORD directed him through Moses. This was to remind the Israelites that no one except a descendant of Aaron should come to burn incense before the LORD, or he would become like Korah and his followers.
NUM|16|41|The next day the whole Israelite community grumbled against Moses and Aaron. "You have killed the LORD's people," they said.
NUM|16|42|But when the assembly gathered in opposition to Moses and Aaron and turned toward the Tent of Meeting, suddenly the cloud covered it and the glory of the LORD appeared.
NUM|16|43|Then Moses and Aaron went to the front of the Tent of Meeting,
NUM|16|44|and the LORD said to Moses,
NUM|16|45|"Get away from this assembly so I can put an end to them at once." And they fell facedown.
NUM|16|46|Then Moses said to Aaron, "Take your censer and put incense in it, along with fire from the altar, and hurry to the assembly to make atonement for them. Wrath has come out from the LORD; the plague has started."
NUM|16|47|So Aaron did as Moses said, and ran into the midst of the assembly. The plague had already started among the people, but Aaron offered the incense and made atonement for them.
NUM|16|48|He stood between the living and the dead, and the plague stopped.
NUM|16|49|But 14,700 people died from the plague, in addition to those who had died because of Korah.
NUM|16|50|Then Aaron returned to Moses at the entrance to the Tent of Meeting, for the plague had stopped.
NUM|17|1|The LORD said to Moses,
NUM|17|2|"Speak to the Israelites and get twelve staffs from them, one from the leader of each of their ancestral tribes. Write the name of each man on his staff.
NUM|17|3|On the staff of Levi write Aaron's name, for there must be one staff for the head of each ancestral tribe.
NUM|17|4|Place them in the Tent of Meeting in front of the Testimony, where I meet with you.
NUM|17|5|The staff belonging to the man I choose will sprout, and I will rid myself of this constant grumbling against you by the Israelites."
NUM|17|6|So Moses spoke to the Israelites, and their leaders gave him twelve staffs, one for the leader of each of their ancestral tribes, and Aaron's staff was among them.
NUM|17|7|Moses placed the staffs before the LORD in the Tent of the Testimony.
NUM|17|8|The next day Moses entered the Tent of the Testimony and saw that Aaron's staff, which represented the house of Levi, had not only sprouted but had budded, blossomed and produced almonds.
NUM|17|9|Then Moses brought out all the staffs from the LORD's presence to all the Israelites. They looked at them, and each man took his own staff.
NUM|17|10|The LORD said to Moses, "Put back Aaron's staff in front of the Testimony, to be kept as a sign to the rebellious. This will put an end to their grumbling against me, so that they will not die."
NUM|17|11|Moses did just as the LORD commanded him.
NUM|17|12|The Israelites said to Moses, "We will die! We are lost, we are all lost!
NUM|17|13|Anyone who even comes near the tabernacle of the LORD will die. Are we all going to die?"
NUM|18|1|The LORD said to Aaron, "You, your sons and your father's family are to bear the responsibility for offenses against the sanctuary, and you and your sons alone are to bear the responsibility for offenses against the priesthood.
NUM|18|2|Bring your fellow Levites from your ancestral tribe to join you and assist you when you and your sons minister before the Tent of the Testimony.
NUM|18|3|They are to be responsible to you and are to perform all the duties of the Tent, but they must not go near the furnishings of the sanctuary or the altar, or both they and you will die.
NUM|18|4|They are to join you and be responsible for the care of the Tent of Meeting-all the work at the Tent-and no one else may come near where you are.
NUM|18|5|"You are to be responsible for the care of the sanctuary and the altar, so that wrath will not fall on the Israelites again.
NUM|18|6|I myself have selected your fellow Levites from among the Israelites as a gift to you, dedicated to the LORD to do the work at the Tent of Meeting.
NUM|18|7|But only you and your sons may serve as priests in connection with everything at the altar and inside the curtain. I am giving you the service of the priesthood as a gift. Anyone else who comes near the sanctuary must be put to death."
NUM|18|8|Then the LORD said to Aaron, "I myself have put you in charge of the offerings presented to me; all the holy offerings the Israelites give me I give to you and your sons as your portion and regular share.
NUM|18|9|You are to have the part of the most holy offerings that is kept from the fire. From all the gifts they bring me as most holy offerings, whether grain or sin or guilt offerings, that part belongs to you and your sons.
NUM|18|10|Eat it as something most holy; every male shall eat it. You must regard it as holy.
NUM|18|11|"This also is yours: whatever is set aside from the gifts of all the wave offerings of the Israelites. I give this to you and your sons and daughters as your regular share. Everyone in your household who is ceremonially clean may eat it.
NUM|18|12|"I give you all the finest olive oil and all the finest new wine and grain they give the LORD as the firstfruits of their harvest.
NUM|18|13|All the land's firstfruits that they bring to the LORD will be yours. Everyone in your household who is ceremonially clean may eat it.
NUM|18|14|"Everything in Israel that is devoted to the LORD is yours.
NUM|18|15|The first offspring of every womb, both man and animal, that is offered to the LORD is yours. But you must redeem every firstborn son and every firstborn male of unclean animals.
NUM|18|16|When they are a month old, you must redeem them at the redemption price set at five shekels of silver, according to the sanctuary shekel, which weighs twenty gerahs.
NUM|18|17|"But you must not redeem the firstborn of an ox, a sheep or a goat; they are holy. Sprinkle their blood on the altar and burn their fat as an offering made by fire, an aroma pleasing to the LORD.
NUM|18|18|Their meat is to be yours, just as the breast of the wave offering and the right thigh are yours.
NUM|18|19|Whatever is set aside from the holy offerings the Israelites present to the LORD I give to you and your sons and daughters as your regular share. It is an everlasting covenant of salt before the LORD for both you and your offspring."
NUM|18|20|The LORD said to Aaron, "You will have no inheritance in their land, nor will you have any share among them; I am your share and your inheritance among the Israelites.
NUM|18|21|"I give to the Levites all the tithes in Israel as their inheritance in return for the work they do while serving at the Tent of Meeting.
NUM|18|22|From now on the Israelites must not go near the Tent of Meeting, or they will bear the consequences of their sin and will die.
NUM|18|23|It is the Levites who are to do the work at the Tent of Meeting and bear the responsibility for offenses against it. This is a lasting ordinance for the generations to come. They will receive no inheritance among the Israelites.
NUM|18|24|Instead, I give to the Levites as their inheritance the tithes that the Israelites present as an offering to the LORD. That is why I said concerning them: 'They will have no inheritance among the Israelites.'"
NUM|18|25|The LORD said to Moses,
NUM|18|26|"Speak to the Levites and say to them: 'When you receive from the Israelites the tithe I give you as your inheritance, you must present a tenth of that tithe as the LORD's offering.
NUM|18|27|Your offering will be reckoned to you as grain from the threshing floor or juice from the winepress.
NUM|18|28|In this way you also will present an offering to the LORD from all the tithes you receive from the Israelites. From these tithes you must give the LORD's portion to Aaron the priest.
NUM|18|29|You must present as the LORD's portion the best and holiest part of everything given to you.'
NUM|18|30|"Say to the Levites: 'When you present the best part, it will be reckoned to you as the product of the threshing floor or the winepress.
NUM|18|31|You and your households may eat the rest of it anywhere, for it is your wages for your work at the Tent of Meeting.
NUM|18|32|By presenting the best part of it you will not be guilty in this matter; then you will not defile the holy offerings of the Israelites, and you will not die.'"
NUM|19|1|The LORD said to Moses and Aaron:
NUM|19|2|"This is a requirement of the law that the LORD has commanded: Tell the Israelites to bring you a red heifer without defect or blemish and that has never been under a yoke.
NUM|19|3|Give it to Eleazar the priest; it is to be taken outside the camp and slaughtered in his presence.
NUM|19|4|Then Eleazar the priest is to take some of its blood on his finger and sprinkle it seven times toward the front of the Tent of Meeting.
NUM|19|5|While he watches, the heifer is to be burned-its hide, flesh, blood and offal.
NUM|19|6|The priest is to take some cedar wood, hyssop and scarlet wool and throw them onto the burning heifer.
NUM|19|7|After that, the priest must wash his clothes and bathe himself with water. He may then come into the camp, but he will be ceremonially unclean till evening.
NUM|19|8|The man who burns it must also wash his clothes and bathe with water, and he too will be unclean till evening.
NUM|19|9|"A man who is clean shall gather up the ashes of the heifer and put them in a ceremonially clean place outside the camp. They shall be kept by the Israelite community for use in the water of cleansing; it is for purification from sin.
NUM|19|10|The man who gathers up the ashes of the heifer must also wash his clothes, and he too will be unclean till evening. This will be a lasting ordinance both for the Israelites and for the aliens living among them.
NUM|19|11|"Whoever touches the dead body of anyone will be unclean for seven days.
NUM|19|12|He must purify himself with the water on the third day and on the seventh day; then he will be clean. But if he does not purify himself on the third and seventh days, he will not be clean.
NUM|19|13|Whoever touches the dead body of anyone and fails to purify himself defiles the LORD's tabernacle. That person must be cut off from Israel. Because the water of cleansing has not been sprinkled on him, he is unclean; his uncleanness remains on him.
NUM|19|14|"This is the law that applies when a person dies in a tent: Anyone who enters the tent and anyone who is in it will be unclean for seven days,
NUM|19|15|and every open container without a lid fastened on it will be unclean.
NUM|19|16|"Anyone out in the open who touches someone who has been killed with a sword or someone who has died a natural death, or anyone who touches a human bone or a grave, will be unclean for seven days.
NUM|19|17|"For the unclean person, put some ashes from the burned purification offering into a jar and pour fresh water over them.
NUM|19|18|Then a man who is ceremonially clean is to take some hyssop, dip it in the water and sprinkle the tent and all the furnishings and the people who were there. He must also sprinkle anyone who has touched a human bone or a grave or someone who has been killed or someone who has died a natural death.
NUM|19|19|The man who is clean is to sprinkle the unclean person on the third and seventh days, and on the seventh day he is to purify him. The person being cleansed must wash his clothes and bathe with water, and that evening he will be clean.
NUM|19|20|But if a person who is unclean does not purify himself, he must be cut off from the community, because he has defiled the sanctuary of the LORD. The water of cleansing has not been sprinkled on him, and he is unclean.
NUM|19|21|This is a lasting ordinance for them. "The man who sprinkles the water of cleansing must also wash his clothes, and anyone who touches the water of cleansing will be unclean till evening.
NUM|19|22|Anything that an unclean person touches becomes unclean, and anyone who touches it becomes unclean till evening."
NUM|20|1|In the first month the whole Israelite community arrived at the Desert of Zin, and they stayed at Kadesh. There Miriam died and was buried.
NUM|20|2|Now there was no water for the community, and the people gathered in opposition to Moses and Aaron.
NUM|20|3|They quarreled with Moses and said, "If only we had died when our brothers fell dead before the LORD!
NUM|20|4|Why did you bring the LORD's community into this desert, that we and our livestock should die here?
NUM|20|5|Why did you bring us up out of Egypt to this terrible place? It has no grain or figs, grapevines or pomegranates. And there is no water to drink!"
NUM|20|6|Moses and Aaron went from the assembly to the entrance to the Tent of Meeting and fell facedown, and the glory of the LORD appeared to them.
NUM|20|7|The LORD said to Moses,
NUM|20|8|"Take the staff, and you and your brother Aaron gather the assembly together. Speak to that rock before their eyes and it will pour out its water. You will bring water out of the rock for the community so they and their livestock can drink."
NUM|20|9|So Moses took the staff from the LORD's presence, just as he commanded him.
NUM|20|10|He and Aaron gathered the assembly together in front of the rock and Moses said to them, "Listen, you rebels, must we bring you water out of this rock?"
NUM|20|11|Then Moses raised his arm and struck the rock twice with his staff. Water gushed out, and the community and their livestock drank.
NUM|20|12|But the LORD said to Moses and Aaron, "Because you did not trust in me enough to honor me as holy in the sight of the Israelites, you will not bring this community into the land I give them."
NUM|20|13|These were the waters of Meribah, where the Israelites quarreled with the LORD and where he showed himself holy among them.
NUM|20|14|Moses sent messengers from Kadesh to the king of Edom, saying: "This is what your brother Israel says: You know about all the hardships that have come upon us.
NUM|20|15|Our forefathers went down into Egypt, and we lived there many years. The Egyptians mistreated us and our fathers,
NUM|20|16|but when we cried out to the LORD, he heard our cry and sent an angel and brought us out of Egypt. "Now we are here at Kadesh, a town on the edge of your territory.
NUM|20|17|Please let us pass through your country. We will not go through any field or vineyard, or drink water from any well. We will travel along the king's highway and not turn to the right or to the left until we have passed through your territory."
NUM|20|18|But Edom answered: "You may not pass through here; if you try, we will march out and attack you with the sword."
NUM|20|19|The Israelites replied: "We will go along the main road, and if we or our livestock drink any of your water, we will pay for it. We only want to pass through on foot-nothing else."
NUM|20|20|Again they answered: "You may not pass through." Then Edom came out against them with a large and powerful army.
NUM|20|21|Since Edom refused to let them go through their territory, Israel turned away from them.
NUM|20|22|The whole Israelite community set out from Kadesh and came to Mount Hor.
NUM|20|23|At Mount Hor, near the border of Edom, the LORD said to Moses and Aaron,
NUM|20|24|"Aaron will be gathered to his people. He will not enter the land I give the Israelites, because both of you rebelled against my command at the waters of Meribah.
NUM|20|25|Get Aaron and his son Eleazar and take them up Mount Hor.
NUM|20|26|Remove Aaron's garments and put them on his son Eleazar, for Aaron will be gathered to his people; he will die there."
NUM|20|27|Moses did as the LORD commanded: They went up Mount Hor in the sight of the whole community.
NUM|20|28|Moses removed Aaron's garments and put them on his son Eleazar. And Aaron died there on top of the mountain. Then Moses and Eleazar came down from the mountain,
NUM|20|29|and when the whole community learned that Aaron had died, the entire house of Israel mourned for him thirty days.
NUM|21|1|When the Canaanite king of Arad, who lived in the Negev, heard that Israel was coming along the road to Atharim, he attacked the Israelites and captured some of them.
NUM|21|2|Then Israel made this vow to the LORD: "If you will deliver these people into our hands, we will totally destroy their cities."
NUM|21|3|The LORD listened to Israel's plea and gave the Canaanites over to them. They completely destroyed them and their towns; so the place was named Hormah.
NUM|21|4|They traveled from Mount Hor along the route to the Red Sea, to go around Edom. But the people grew impatient on the way;
NUM|21|5|they spoke against God and against Moses, and said, "Why have you brought us up out of Egypt to die in the desert? There is no bread! There is no water! And we detest this miserable food!"
NUM|21|6|Then the LORD sent venomous snakes among them; they bit the people and many Israelites died.
NUM|21|7|The people came to Moses and said, "We sinned when we spoke against the LORD and against you. Pray that the LORD will take the snakes away from us." So Moses prayed for the people.
NUM|21|8|The LORD said to Moses, "Make a snake and put it up on a pole; anyone who is bitten can look at it and live."
NUM|21|9|So Moses made a bronze snake and put it up on a pole. Then when anyone was bitten by a snake and looked at the bronze snake, he lived.
NUM|21|10|The Israelites moved on and camped at Oboth.
NUM|21|11|Then they set out from Oboth and camped in Iye Abarim, in the desert that faces Moab toward the sunrise.
NUM|21|12|From there they moved on and camped in the Zered Valley.
NUM|21|13|They set out from there and camped alongside the Arnon, which is in the desert extending into Amorite territory. The Arnon is the border of Moab, between Moab and the Amorites.
NUM|21|14|That is why the Book of the Wars of the LORD says: "...Waheb in Suphah and the ravines, the Arnon
NUM|21|15|and the slopes of the ravines that lead to the site of Ar and lie along the border of Moab."
NUM|21|16|From there they continued on to Beer, the well where the LORD said to Moses, "Gather the people together and I will give them water."
NUM|21|17|Then Israel sang this song: "Spring up, O well! Sing about it,
NUM|21|18|about the well that the princes dug, that the nobles of the people sank- the nobles with scepters and staffs." Then they went from the desert to Mattanah,
NUM|21|19|from Mattanah to Nahaliel, from Nahaliel to Bamoth,
NUM|21|20|and from Bamoth to the valley in Moab where the top of Pisgah overlooks the wasteland.
NUM|21|21|Israel sent messengers to say to Sihon king of the Amorites:
NUM|21|22|"Let us pass through your country. We will not turn aside into any field or vineyard, or drink water from any well. We will travel along the king's highway until we have passed through your territory."
NUM|21|23|But Sihon would not let Israel pass through his territory. He mustered his entire army and marched out into the desert against Israel. When he reached Jahaz, he fought with Israel.
NUM|21|24|Israel, however, put him to the sword and took over his land from the Arnon to the Jabbok, but only as far as the Ammonites, because their border was fortified.
NUM|21|25|Israel captured all the cities of the Amorites and occupied them, including Heshbon and all its surrounding settlements.
NUM|21|26|Heshbon was the city of Sihon king of the Amorites, who had fought against the former king of Moab and had taken from him all his land as far as the Arnon.
NUM|21|27|That is why the poets say: "Come to Heshbon and let it be rebuilt; let Sihon's city be restored.
NUM|21|28|"Fire went out from Heshbon, a blaze from the city of Sihon. It consumed Ar of Moab, the citizens of Arnon's heights.
NUM|21|29|Woe to you, O Moab! You are destroyed, O people of Chemosh! He has given up his sons as fugitives and his daughters as captives to Sihon king of the Amorites.
NUM|21|30|"But we have overthrown them; Heshbon is destroyed all the way to Dibon. We have demolished them as far as Nophah, which extends to Medeba."
NUM|21|31|So Israel settled in the land of the Amorites.
NUM|21|32|After Moses had sent spies to Jazer, the Israelites captured its surrounding settlements and drove out the Amorites who were there.
NUM|21|33|Then they turned and went up along the road toward Bashan, and Og king of Bashan and his whole army marched out to meet them in battle at Edrei.
NUM|21|34|The LORD said to Moses, "Do not be afraid of him, for I have handed him over to you, with his whole army and his land. Do to him what you did to Sihon king of the Amorites, who reigned in Heshbon."
NUM|21|35|So they struck him down, together with his sons and his whole army, leaving them no survivors. And they took possession of his land.
NUM|22|1|Then the Israelites traveled to the plains of Moab and camped along the Jordan across from Jericho.
NUM|22|2|Now Balak son of Zippor saw all that Israel had done to the Amorites,
NUM|22|3|and Moab was terrified because there were so many people. Indeed, Moab was filled with dread because of the Israelites.
NUM|22|4|The Moabites said to the elders of Midian, "This horde is going to lick up everything around us, as an ox licks up the grass of the field." So Balak son of Zippor, who was king of Moab at that time,
NUM|22|5|sent messengers to summon Balaam son of Beor, who was at Pethor, near the River, in his native land. Balak said: "A people has come out of Egypt; they cover the face of the land and have settled next to me.
NUM|22|6|Now come and put a curse on these people, because they are too powerful for me. Perhaps then I will be able to defeat them and drive them out of the country. For I know that those you bless are blessed, and those you curse are cursed."
NUM|22|7|The elders of Moab and Midian left, taking with them the fee for divination. When they came to Balaam, they told him what Balak had said.
NUM|22|8|"Spend the night here," Balaam said to them, "and I will bring you back the answer the LORD gives me." So the Moabite princes stayed with him.
NUM|22|9|God came to Balaam and asked, "Who are these men with you?"
NUM|22|10|Balaam said to God, "Balak son of Zippor, king of Moab, sent me this message:
NUM|22|11|'A people that has come out of Egypt covers the face of the land. Now come and put a curse on them for me. Perhaps then I will be able to fight them and drive them away.'"
NUM|22|12|But God said to Balaam, "Do not go with them. You must not put a curse on those people, because they are blessed."
NUM|22|13|The next morning Balaam got up and said to Balak's princes, "Go back to your own country, for the LORD has refused to let me go with you."
NUM|22|14|So the Moabite princes returned to Balak and said, "Balaam refused to come with us."
NUM|22|15|Then Balak sent other princes, more numerous and more distinguished than the first.
NUM|22|16|They came to Balaam and said: "This is what Balak son of Zippor says: Do not let anything keep you from coming to me,
NUM|22|17|because I will reward you handsomely and do whatever you say. Come and put a curse on these people for me."
NUM|22|18|But Balaam answered them, "Even if Balak gave me his palace filled with silver and gold, I could not do anything great or small to go beyond the command of the LORD my God.
NUM|22|19|Now stay here tonight as the others did, and I will find out what else the LORD will tell me."
NUM|22|20|That night God came to Balaam and said, "Since these men have come to summon you, go with them, but do only what I tell you."
NUM|22|21|Balaam got up in the morning, saddled his donkey and went with the princes of Moab.
NUM|22|22|But God was very angry when he went, and the angel of the LORD stood in the road to oppose him. Balaam was riding on his donkey, and his two servants were with him.
NUM|22|23|When the donkey saw the angel of the LORD standing in the road with a drawn sword in his hand, she turned off the road into a field. Balaam beat her to get her back on the road.
NUM|22|24|Then the angel of the LORD stood in a narrow path between two vineyards, with walls on both sides.
NUM|22|25|When the donkey saw the angel of the LORD, she pressed close to the wall, crushing Balaam's foot against it. So he beat her again.
NUM|22|26|Then the angel of the LORD moved on ahead and stood in a narrow place where there was no room to turn, either to the right or to the left.
NUM|22|27|When the donkey saw the angel of the LORD, she lay down under Balaam, and he was angry and beat her with his staff.
NUM|22|28|Then the LORD opened the donkey's mouth, and she said to Balaam, "What have I done to you to make you beat me these three times?"
NUM|22|29|Balaam answered the donkey, "You have made a fool of me! If I had a sword in my hand, I would kill you right now."
NUM|22|30|The donkey said to Balaam, "Am I not your own donkey, which you have always ridden, to this day? Have I been in the habit of doing this to you?No," he said.
NUM|22|31|Then the LORD opened Balaam's eyes, and he saw the angel of the LORD standing in the road with his sword drawn. So he bowed low and fell facedown.
NUM|22|32|The angel of the LORD asked him, "Why have you beaten your donkey these three times? I have come here to oppose you because your path is a reckless one before me.
NUM|22|33|The donkey saw me and turned away from me these three times. If she had not turned away, I would certainly have killed you by now, but I would have spared her."
NUM|22|34|Balaam said to the angel of the LORD, "I have sinned. I did not realize you were standing in the road to oppose me. Now if you are displeased, I will go back."
NUM|22|35|The angel of the LORD said to Balaam, "Go with the men, but speak only what I tell you." So Balaam went with the princes of Balak.
NUM|22|36|When Balak heard that Balaam was coming, he went out to meet him at the Moabite town on the Arnon border, at the edge of his territory.
NUM|22|37|Balak said to Balaam, "Did I not send you an urgent summons? Why didn't you come to me? Am I really not able to reward you?"
NUM|22|38|"Well, I have come to you now," Balaam replied. "But can I say just anything? I must speak only what God puts in my mouth."
NUM|22|39|Then Balaam went with Balak to Kiriath Huzoth.
NUM|22|40|Balak sacrificed cattle and sheep, and gave some to Balaam and the princes who were with him.
NUM|22|41|The next morning Balak took Balaam up to Bamoth Baal, and from there he saw part of the people.
NUM|23|1|Balaam said, "Build me seven altars here, and prepare seven bulls and seven rams for me."
NUM|23|2|Balak did as Balaam said, and the two of them offered a bull and a ram on each altar.
NUM|23|3|Then Balaam said to Balak, "Stay here beside your offering while I go aside. Perhaps the LORD will come to meet with me. Whatever he reveals to me I will tell you." Then he went off to a barren height.
NUM|23|4|God met with him, and Balaam said, "I have prepared seven altars, and on each altar I have offered a bull and a ram."
NUM|23|5|The LORD put a message in Balaam's mouth and said, "Go back to Balak and give him this message."
NUM|23|6|So he went back to him and found him standing beside his offering, with all the princes of Moab.
NUM|23|7|Then Balaam uttered his oracle: "Balak brought me from Aram, the king of Moab from the eastern mountains. 'Come,' he said, 'curse Jacob for me; come, denounce Israel.'
NUM|23|8|How can I curse those whom God has not cursed? How can I denounce those whom the LORD has not denounced?
NUM|23|9|From the rocky peaks I see them, from the heights I view them. I see a people who live apart and do not consider themselves one of the nations.
NUM|23|10|Who can count the dust of Jacob or number the fourth part of Israel? Let me die the death of the righteous, and may my end be like theirs!"
NUM|23|11|Balak said to Balaam, "What have you done to me? I brought you to curse my enemies, but you have done nothing but bless them!"
NUM|23|12|He answered, "Must I not speak what the LORD puts in my mouth?"
NUM|23|13|Then Balak said to him, "Come with me to another place where you can see them; you will see only a part but not all of them. And from there, curse them for me."
NUM|23|14|So he took him to the field of Zophim on the top of Pisgah, and there he built seven altars and offered a bull and a ram on each altar.
NUM|23|15|Balaam said to Balak, "Stay here beside your offering while I meet with him over there."
NUM|23|16|The LORD met with Balaam and put a message in his mouth and said, "Go back to Balak and give him this message."
NUM|23|17|So he went to him and found him standing beside his offering, with the princes of Moab. Balak asked him, "What did the LORD say?"
NUM|23|18|Then he uttered his oracle: "Arise, Balak, and listen; hear me, son of Zippor.
NUM|23|19|God is not a man, that he should lie, nor a son of man, that he should change his mind. Does he speak and then not act? Does he promise and not fulfill?
NUM|23|20|I have received a command to bless; he has blessed, and I cannot change it.
NUM|23|21|"No misfortune is seen in Jacob, no misery observed in Israel. The LORD their God is with them; the shout of the King is among them.
NUM|23|22|God brought them out of Egypt; they have the strength of a wild ox.
NUM|23|23|There is no sorcery against Jacob, no divination against Israel. It will now be said of Jacob and of Israel, 'See what God has done!'
NUM|23|24|The people rise like a lioness; they rouse themselves like a lion that does not rest till he devours his prey and drinks the blood of his victims."
NUM|23|25|Then Balak said to Balaam, "Neither curse them at all nor bless them at all!"
NUM|23|26|Balaam answered, "Did I not tell you I must do whatever the LORD says?"
NUM|23|27|Then Balak said to Balaam, "Come, let me take you to another place. Perhaps it will please God to let you curse them for me from there."
NUM|23|28|And Balak took Balaam to the top of Peor, overlooking the wasteland.
NUM|23|29|Balaam said, "Build me seven altars here, and prepare seven bulls and seven rams for me."
NUM|23|30|Balak did as Balaam had said, and offered a bull and a ram on each altar.
NUM|24|1|Now when Balaam saw that it pleased the LORD to bless Israel, he did not resort to sorcery as at other times, but turned his face toward the desert.
NUM|24|2|When Balaam looked out and saw Israel encamped tribe by tribe, the Spirit of God came upon him
NUM|24|3|and he uttered his oracle: "The oracle of Balaam son of Beor, the oracle of one whose eye sees clearly,
NUM|24|4|the oracle of one who hears the words of God, who sees a vision from the Almighty, who falls prostrate, and whose eyes are opened:
NUM|24|5|"How beautiful are your tents, O Jacob, your dwelling places, O Israel!
NUM|24|6|"Like valleys they spread out, like gardens beside a river, like aloes planted by the LORD, like cedars beside the waters.
NUM|24|7|Water will flow from their buckets; their seed will have abundant water. "Their king will be greater than Agag; their kingdom will be exalted.
NUM|24|8|"God brought them out of Egypt; they have the strength of a wild ox. They devour hostile nations and break their bones in pieces; with their arrows they pierce them.
NUM|24|9|Like a lion they crouch and lie down, like a lioness-who dares to rouse them? "May those who bless you be blessed and those who curse you be cursed!"
NUM|24|10|Then Balak's anger burned against Balaam. He struck his hands together and said to him, "I summoned you to curse my enemies, but you have blessed them these three times.
NUM|24|11|Now leave at once and go home! I said I would reward you handsomely, but the LORD has kept you from being rewarded."
NUM|24|12|Balaam answered Balak, "Did I not tell the messengers you sent me,
NUM|24|13|'Even if Balak gave me his palace filled with silver and gold, I could not do anything of my own accord, good or bad, to go beyond the command of the LORD -and I must say only what the LORD says'?
NUM|24|14|Now I am going back to my people, but come, let me warn you of what this people will do to your people in days to come."
NUM|24|15|Then he uttered his oracle: "The oracle of Balaam son of Beor, the oracle of one whose eye sees clearly,
NUM|24|16|the oracle of one who hears the words of God, who has knowledge from the Most High, who sees a vision from the Almighty, who falls prostrate, and whose eyes are opened:
NUM|24|17|"I see him, but not now; I behold him, but not near. A star will come out of Jacob; a scepter will rise out of Israel. He will crush the foreheads of Moab, the skulls of all the sons of Sheth.
NUM|24|18|Edom will be conquered; Seir, his enemy, will be conquered, but Israel will grow strong.
NUM|24|19|A ruler will come out of Jacob and destroy the survivors of the city."
NUM|24|20|Then Balaam saw Amalek and uttered his oracle: "Amalek was first among the nations, but he will come to ruin at last."
NUM|24|21|Then he saw the Kenites and uttered his oracle: "Your dwelling place is secure, your nest is set in a rock;
NUM|24|22|yet you Kenites will be destroyed when Asshur takes you captive."
NUM|24|23|Then he uttered his oracle: "Ah, who can live when God does this?
NUM|24|24|Ships will come from the shores of Kittim; they will subdue Asshur and Eber, but they too will come to ruin."
NUM|24|25|Then Balaam got up and returned home and Balak went his own way.
NUM|25|1|While Israel was staying in Shittim, the men began to indulge in sexual immorality with Moabite women,
NUM|25|2|who invited them to the sacrifices to their gods. The people ate and bowed down before these gods.
NUM|25|3|So Israel joined in worshiping the Baal of Peor. And the LORD's anger burned against them.
NUM|25|4|The LORD said to Moses, "Take all the leaders of these people, kill them and expose them in broad daylight before the LORD, so that the LORD's fierce anger may turn away from Israel."
NUM|25|5|So Moses said to Israel's judges, "Each of you must put to death those of your men who have joined in worshiping the Baal of Peor."
NUM|25|6|Then an Israelite man brought to his family a Midianite woman right before the eyes of Moses and the whole assembly of Israel while they were weeping at the entrance to the Tent of Meeting.
NUM|25|7|When Phinehas son of Eleazar, the son of Aaron, the priest, saw this, he left the assembly, took a spear in his hand
NUM|25|8|and followed the Israelite into the tent. He drove the spear through both of them-through the Israelite and into the woman's body. Then the plague against the Israelites was stopped;
NUM|25|9|but those who died in the plague numbered 24,000.
NUM|25|10|The LORD said to Moses,
NUM|25|11|"Phinehas son of Eleazar, the son of Aaron, the priest, has turned my anger away from the Israelites; for he was as zealous as I am for my honor among them, so that in my zeal I did not put an end to them.
NUM|25|12|Therefore tell him I am making my covenant of peace with him.
NUM|25|13|He and his descendants will have a covenant of a lasting priesthood, because he was zealous for the honor of his God and made atonement for the Israelites."
NUM|25|14|The name of the Israelite who was killed with the Midianite woman was Zimri son of Salu, the leader of a Simeonite family.
NUM|25|15|And the name of the Midianite woman who was put to death was Cozbi daughter of Zur, a tribal chief of a Midianite family.
NUM|25|16|The LORD said to Moses,
NUM|25|17|"Treat the Midianites as enemies and kill them,
NUM|25|18|because they treated you as enemies when they deceived you in the affair of Peor and their sister Cozbi, the daughter of a Midianite leader, the woman who was killed when the plague came as a result of Peor."
NUM|26|1|After the plague the LORD said to Moses and Eleazar son of Aaron, the priest,
NUM|26|2|"Take a census of the whole Israelite community by families-all those twenty years old or more who are able to serve in the army of Israel."
NUM|26|3|So on the plains of Moab by the Jordan across from Jericho, Moses and Eleazar the priest spoke with them and said,
NUM|26|4|"Take a census of the men twenty years old or more, as the LORD commanded Moses." These were the Israelites who came out of Egypt:
NUM|26|5|The descendants of Reuben, the firstborn son of Israel, were: through Hanoch, the Hanochite clan; through Pallu, the Palluite clan;
NUM|26|6|through Hezron, the Hezronite clan; through Carmi, the Carmite clan.
NUM|26|7|These were the clans of Reuben; those numbered were 43,730.
NUM|26|8|The son of Pallu was Eliab,
NUM|26|9|and the sons of Eliab were Nemuel, Dathan and Abiram. The same Dathan and Abiram were the community officials who rebelled against Moses and Aaron and were among Korah's followers when they rebelled against the LORD.
NUM|26|10|The earth opened its mouth and swallowed them along with Korah, whose followers died when the fire devoured the 250 men. And they served as a warning sign.
NUM|26|11|The line of Korah, however, did not die out.
NUM|26|12|The descendants of Simeon by their clans were: through Nemuel, the Nemuelite clan; through Jamin, the Jaminite clan; through Jakin, the Jakinite clan;
NUM|26|13|through Zerah, the Zerahite clan; through Shaul, the Shaulite clan.
NUM|26|14|These were the clans of Simeon; there were 22,200 men.
NUM|26|15|The descendants of Gad by their clans were: through Zephon, the Zephonite clan; through Haggi, the Haggite clan; through Shuni, the Shunite clan;
NUM|26|16|through Ozni, the Oznite clan; through Eri, the Erite clan;
NUM|26|17|through Arodi, the Arodite clan; through Areli, the Arelite clan.
NUM|26|18|These were the clans of Gad; those numbered were 40,500.
NUM|26|19|Er and Onan were sons of Judah, but they died in Canaan.
NUM|26|20|The descendants of Judah by their clans were: through Shelah, the Shelanite clan; through Perez, the Perezite clan; through Zerah, the Zerahite clan.
NUM|26|21|The descendants of Perez were: through Hezron, the Hezronite clan; through Hamul, the Hamulite clan.
NUM|26|22|These were the clans of Judah; those numbered were 76,500.
NUM|26|23|The descendants of Issachar by their clans were: through Tola, the Tolaite clan; through Puah, the Puite clan;
NUM|26|24|through Jashub, the Jashubite clan; through Shimron, the Shimronite clan.
NUM|26|25|These were the clans of Issachar; those numbered were 64,300.
NUM|26|26|The descendants of Zebulun by their clans were: through Sered, the Seredite clan; through Elon, the Elonite clan; through Jahleel, the Jahleelite clan.
NUM|26|27|These were the clans of Zebulun; those numbered were 60,500.
NUM|26|28|The descendants of Joseph by their clans through Manasseh and Ephraim were:
NUM|26|29|The descendants of Manasseh: through Makir, the Makirite clan (Makir was the father of Gilead); through Gilead, the Gileadite clan.
NUM|26|30|These were the descendants of Gilead: through Iezer, the Iezerite clan; through Helek, the Helekite clan;
NUM|26|31|through Asriel, the Asrielite clan; through Shechem, the Shechemite clan;
NUM|26|32|through Shemida, the Shemidaite clan; through Hepher, the Hepherite clan.
NUM|26|33|(Zelophehad son of Hepher had no sons; he had only daughters, whose names were Mahlah, Noah, Hoglah, Milcah and Tirzah.)
NUM|26|34|These were the clans of Manasseh; those numbered were 52,700.
NUM|26|35|These were the descendants of Ephraim by their clans: through Shuthelah, the Shuthelahite clan; through Beker, the Bekerite clan; through Tahan, the Tahanite clan.
NUM|26|36|These were the descendants of Shuthelah: through Eran, the Eranite clan.
NUM|26|37|These were the clans of Ephraim; those numbered were 32,500. These were the descendants of Joseph by their clans.
NUM|26|38|The descendants of Benjamin by their clans were: through Bela, the Belaite clan; through Ashbel, the Ashbelite clan; through Ahiram, the Ahiramite clan;
NUM|26|39|through Shupham, the Shuphamite clan; through Hupham, the Huphamite clan.
NUM|26|40|The descendants of Bela through Ard and Naaman were: through Ard, the Ardite clan; through Naaman, the Naamite clan.
NUM|26|41|These were the clans of Benjamin; those numbered were 45,600.
NUM|26|42|These were the descendants of Dan by their clans: through Shuham, the Shuhamite clan. These were the clans of Dan:
NUM|26|43|All of them were Shuhamite clans; and those numbered were 64,400.
NUM|26|44|The descendants of Asher by their clans were: through Imnah, the Imnite clan; through Ishvi, the Ishvite clan; through Beriah, the Beriite clan;
NUM|26|45|and through the descendants of Beriah: through Heber, the Heberite clan; through Malkiel, the Malkielite clan.
NUM|26|46|(Asher had a daughter named Serah.)
NUM|26|47|These were the clans of Asher; those numbered were 53,400.
NUM|26|48|The descendants of Naphtali by their clans were: through Jahzeel, the Jahzeelite clan; through Guni, the Gunite clan;
NUM|26|49|through Jezer, the Jezerite clan; through Shillem, the Shillemite clan.
NUM|26|50|These were the clans of Naphtali; those numbered were 45,400.
NUM|26|51|The total number of the men of Israel was 601,730.
NUM|26|52|The LORD said to Moses,
NUM|26|53|"The land is to be allotted to them as an inheritance based on the number of names.
NUM|26|54|To a larger group give a larger inheritance, and to a smaller group a smaller one; each is to receive its inheritance according to the number of those listed.
NUM|26|55|Be sure that the land is distributed by lot. What each group inherits will be according to the names for its ancestral tribe.
NUM|26|56|Each inheritance is to be distributed by lot among the larger and smaller groups."
NUM|26|57|These were the Levites who were counted by their clans: through Gershon, the Gershonite clan; through Kohath, the Kohathite clan; through Merari, the Merarite clan.
NUM|26|58|These also were Levite clans: the Libnite clan, the Hebronite clan, the Mahlite clan, the Mushite clan, the Korahite clan. (Kohath was the forefather of Amram;
NUM|26|59|the name of Amram's wife was Jochebed, a descendant of Levi, who was born to the Levites in Egypt. To Amram she bore Aaron, Moses and their sister Miriam.
NUM|26|60|Aaron was the father of Nadab and Abihu, Eleazar and Ithamar.
NUM|26|61|But Nadab and Abihu died when they made an offering before the LORD with unauthorized fire.)
NUM|26|62|All the male Levites a month old or more numbered 23,000. They were not counted along with the other Israelites because they received no inheritance among them.
NUM|26|63|These are the ones counted by Moses and Eleazar the priest when they counted the Israelites on the plains of Moab by the Jordan across from Jericho.
NUM|26|64|Not one of them was among those counted by Moses and Aaron the priest when they counted the Israelites in the Desert of Sinai.
NUM|26|65|For the LORD had told those Israelites they would surely die in the desert, and not one of them was left except Caleb son of Jephunneh and Joshua son of Nun.
NUM|27|1|The daughters of Zelophehad son of Hepher, the son of Gilead, the son of Makir, the son of Manasseh, belonged to the clans of Manasseh son of Joseph. The names of the daughters were Mahlah, Noah, Hoglah, Milcah and Tirzah. They approached
NUM|27|2|the entrance to the Tent of Meeting and stood before Moses, Eleazar the priest, the leaders and the whole assembly, and said,
NUM|27|3|"Our father died in the desert. He was not among Korah's followers, who banded together against the LORD, but he died for his own sin and left no sons.
NUM|27|4|Why should our father's name disappear from his clan because he had no son? Give us property among our father's relatives."
NUM|27|5|So Moses brought their case before the LORD
NUM|27|6|and the LORD said to him,
NUM|27|7|"What Zelophehad's daughters are saying is right. You must certainly give them property as an inheritance among their father's relatives and turn their father's inheritance over to them.
NUM|27|8|"Say to the Israelites, 'If a man dies and leaves no son, turn his inheritance over to his daughter.
NUM|27|9|If he has no daughter, give his inheritance to his brothers.
NUM|27|10|If he has no brothers, give his inheritance to his father's brothers.
NUM|27|11|If his father had no brothers, give his inheritance to the nearest relative in his clan, that he may possess it. This is to be a legal requirement for the Israelites, as the LORD commanded Moses.'"
NUM|27|12|Then the LORD said to Moses, "Go up this mountain in the Abarim range and see the land I have given the Israelites.
NUM|27|13|After you have seen it, you too will be gathered to your people, as your brother Aaron was,
NUM|27|14|for when the community rebelled at the waters in the Desert of Zin, both of you disobeyed my command to honor me as holy before their eyes." (These were the waters of Meribah Kadesh, in the Desert of Zin.)
NUM|27|15|Moses said to the LORD,
NUM|27|16|"May the LORD, the God of the spirits of all mankind, appoint a man over this community
NUM|27|17|to go out and come in before them, one who will lead them out and bring them in, so the LORD's people will not be like sheep without a shepherd."
NUM|27|18|So the LORD said to Moses, "Take Joshua son of Nun, a man in whom is the spirit, and lay your hand on him.
NUM|27|19|Have him stand before Eleazar the priest and the entire assembly and commission him in their presence.
NUM|27|20|Give him some of your authority so the whole Israelite community will obey him.
NUM|27|21|He is to stand before Eleazar the priest, who will obtain decisions for him by inquiring of the Urim before the LORD. At his command he and the entire community of the Israelites will go out, and at his command they will come in."
NUM|27|22|Moses did as the LORD commanded him. He took Joshua and had him stand before Eleazar the priest and the whole assembly.
NUM|27|23|Then he laid his hands on him and commissioned him, as the LORD instructed through Moses.
NUM|28|1|The LORD said to Moses,
NUM|28|2|"Give this command to the Israelites and say to them: 'See that you present to me at the appointed time the food for my offerings made by fire, as an aroma pleasing to me.'
NUM|28|3|Say to them: 'This is the offering made by fire that you are to present to the LORD: two lambs a year old without defect, as a regular burnt offering each day.
NUM|28|4|Prepare one lamb in the morning and the other at twilight,
NUM|28|5|together with a grain offering of a tenth of an ephah of fine flour mixed with a quarter of a hin of oil from pressed olives.
NUM|28|6|This is the regular burnt offering instituted at Mount Sinai as a pleasing aroma, an offering made to the LORD by fire.
NUM|28|7|The accompanying drink offering is to be a quarter of a hin of fermented drink with each lamb. Pour out the drink offering to the LORD at the sanctuary.
NUM|28|8|Prepare the second lamb at twilight, along with the same kind of grain offering and drink offering that you prepare in the morning. This is an offering made by fire, an aroma pleasing to the LORD.
NUM|28|9|"'On the Sabbath day, make an offering of two lambs a year old without defect, together with its drink offering and a grain offering of two-tenths of an ephah of fine flour mixed with oil.
NUM|28|10|This is the burnt offering for every Sabbath, in addition to the regular burnt offering and its drink offering.
NUM|28|11|"'On the first of every month, present to the LORD a burnt offering of two young bulls, one ram and seven male lambs a year old, all without defect.
NUM|28|12|With each bull there is to be a grain offering of three-tenths of an ephah of fine flour mixed with oil; with the ram, a grain offering of two-tenths of an ephah of fine flour mixed with oil;
NUM|28|13|and with each lamb, a grain offering of a tenth of an ephah of fine flour mixed with oil. This is for a burnt offering, a pleasing aroma, an offering made to the LORD by fire.
NUM|28|14|With each bull there is to be a drink offering of half a hin of wine; with the ram, a third of a hin; and with each lamb, a quarter of a hin. This is the monthly burnt offering to be made at each new moon during the year.
NUM|28|15|Besides the regular burnt offering with its drink offering, one male goat is to be presented to the LORD as a sin offering.
NUM|28|16|"'On the fourteenth day of the first month the LORD's Passover is to be held.
NUM|28|17|On the fifteenth day of this month there is to be a festival; for seven days eat bread made without yeast.
NUM|28|18|On the first day hold a sacred assembly and do no regular work.
NUM|28|19|Present to the LORD an offering made by fire, a burnt offering of two young bulls, one ram and seven male lambs a year old, all without defect.
NUM|28|20|With each bull prepare a grain offering of three-tenths of an ephah of fine flour mixed with oil; with the ram, two-tenths;
NUM|28|21|and with each of the seven lambs, one-tenth.
NUM|28|22|Include one male goat as a sin offering to make atonement for you.
NUM|28|23|Prepare these in addition to the regular morning burnt offering.
NUM|28|24|In this way prepare the food for the offering made by fire every day for seven days as an aroma pleasing to the LORD; it is to be prepared in addition to the regular burnt offering and its drink offering.
NUM|28|25|On the seventh day hold a sacred assembly and do no regular work.
NUM|28|26|"'On the day of firstfruits, when you present to the LORD an offering of new grain during the Feast of Weeks, hold a sacred assembly and do no regular work.
NUM|28|27|Present a burnt offering of two young bulls, one ram and seven male lambs a year old as an aroma pleasing to the LORD.
NUM|28|28|With each bull there is to be a grain offering of three-tenths of an ephah of fine flour mixed with oil; with the ram, two-tenths;
NUM|28|29|and with each of the seven lambs, one-tenth.
NUM|28|30|Include one male goat to make atonement for you.
NUM|28|31|Prepare these together with their drink offerings, in addition to the regular burnt offering and its grain offering. Be sure the animals are without defect.
NUM|29|1|"'On the first day of the seventh month hold a sacred assembly and do no regular work. It is a day for you to sound the trumpets.
NUM|29|2|As an aroma pleasing to the LORD, prepare a burnt offering of one young bull, one ram and seven male lambs a year old, all without defect.
NUM|29|3|With the bull prepare a grain offering of three-tenths of an ephah of fine flour mixed with oil; with the ram, two-tenths;
NUM|29|4|and with each of the seven lambs, one-tenth.
NUM|29|5|Include one male goat as a sin offering to make atonement for you.
NUM|29|6|These are in addition to the monthly and daily burnt offerings with their grain offerings and drink offerings as specified. They are offerings made to the LORD by fire-a pleasing aroma.
NUM|29|7|"'On the tenth day of this seventh month hold a sacred assembly. You must deny yourselves and do no work.
NUM|29|8|Present as an aroma pleasing to the LORD a burnt offering of one young bull, one ram and seven male lambs a year old, all without defect.
NUM|29|9|With the bull prepare a grain offering of three-tenths of an ephah of fine flour mixed with oil; with the ram, two-tenths;
NUM|29|10|and with each of the seven lambs, one-tenth.
NUM|29|11|Include one male goat as a sin offering, in addition to the sin offering for atonement and the regular burnt offering with its grain offering, and their drink offerings.
NUM|29|12|"'On the fifteenth day of the seventh month, hold a sacred assembly and do no regular work. Celebrate a festival to the LORD for seven days.
NUM|29|13|Present an offering made by fire as an aroma pleasing to the LORD, a burnt offering of thirteen young bulls, two rams and fourteen male lambs a year old, all without defect.
NUM|29|14|With each of the thirteen bulls prepare a grain offering of three-tenths of an ephah of fine flour mixed with oil; with each of the two rams, two-tenths;
NUM|29|15|and with each of the fourteen lambs, one-tenth.
NUM|29|16|Include one male goat as a sin offering, in addition to the regular burnt offering with its grain offering and drink offering.
NUM|29|17|"'On the second day prepare twelve young bulls, two rams and fourteen male lambs a year old, all without defect.
NUM|29|18|With the bulls, rams and lambs, prepare their grain offerings and drink offerings according to the number specified.
NUM|29|19|Include one male goat as a sin offering, in addition to the regular burnt offering with its grain offering, and their drink offerings.
NUM|29|20|"'On the third day prepare eleven bulls, two rams and fourteen male lambs a year old, all without defect.
NUM|29|21|With the bulls, rams and lambs, prepare their grain offerings and drink offerings according to the number specified.
NUM|29|22|Include one male goat as a sin offering, in addition to the regular burnt offering with its grain offering and drink offering.
NUM|29|23|"'On the fourth day prepare ten bulls, two rams and fourteen male lambs a year old, all without defect.
NUM|29|24|With the bulls, rams and lambs, prepare their grain offerings and drink offerings according to the number specified.
NUM|29|25|Include one male goat as a sin offering, in addition to the regular burnt offering with its grain offering and drink offering.
NUM|29|26|"'On the fifth day prepare nine bulls, two rams and fourteen male lambs a year old, all without defect.
NUM|29|27|With the bulls, rams and lambs, prepare their grain offerings and drink offerings according to the number specified.
NUM|29|28|Include one male goat as a sin offering, in addition to the regular burnt offering with its grain offering and drink offering.
NUM|29|29|"'On the sixth day prepare eight bulls, two rams and fourteen male lambs a year old, all without defect.
NUM|29|30|With the bulls, rams and lambs, prepare their grain offerings and drink offerings according to the number specified.
NUM|29|31|Include one male goat as a sin offering, in addition to the regular burnt offering with its grain offering and drink offering.
NUM|29|32|"'On the seventh day prepare seven bulls, two rams and fourteen male lambs a year old, all without defect.
NUM|29|33|With the bulls, rams and lambs, prepare their grain offerings and drink offerings according to the number specified.
NUM|29|34|Include one male goat as a sin offering, in addition to the regular burnt offering with its grain offering and drink offering.
NUM|29|35|"'On the eighth day hold an assembly and do no regular work.
NUM|29|36|Present an offering made by fire as an aroma pleasing to the LORD, a burnt offering of one bull, one ram and seven male lambs a year old, all without defect.
NUM|29|37|With the bull, the ram and the lambs, prepare their grain offerings and drink offerings according to the number specified.
NUM|29|38|Include one male goat as a sin offering, in addition to the regular burnt offering with its grain offering and drink offering.
NUM|29|39|"'In addition to what you vow and your freewill offerings, prepare these for the LORD at your appointed feasts: your burnt offerings, grain offerings, drink offerings and fellowship offerings. '"
NUM|29|40|Moses told the Israelites all that the LORD commanded him.
NUM|30|1|Moses said to the heads of the tribes of Israel: "This is what the LORD commands:
NUM|30|2|When a man makes a vow to the LORD or takes an oath to obligate himself by a pledge, he must not break his word but must do everything he said.
NUM|30|3|"When a young woman still living in her father's house makes a vow to the LORD or obligates herself by a pledge
NUM|30|4|and her father hears about her vow or pledge but says nothing to her, then all her vows and every pledge by which she obligated herself will stand.
NUM|30|5|But if her father forbids her when he hears about it, none of her vows or the pledges by which she obligated herself will stand; the LORD will release her because her father has forbidden her.
NUM|30|6|"If she marries after she makes a vow or after her lips utter a rash promise by which she obligates herself
NUM|30|7|and her husband hears about it but says nothing to her, then her vows or the pledges by which she obligated herself will stand.
NUM|30|8|But if her husband forbids her when he hears about it, he nullifies the vow that obligates her or the rash promise by which she obligates herself, and the LORD will release her.
NUM|30|9|"Any vow or obligation taken by a widow or divorced woman will be binding on her.
NUM|30|10|"If a woman living with her husband makes a vow or obligates herself by a pledge under oath
NUM|30|11|and her husband hears about it but says nothing to her and does not forbid her, then all her vows or the pledges by which she obligated herself will stand.
NUM|30|12|But if her husband nullifies them when he hears about them, then none of the vows or pledges that came from her lips will stand. Her husband has nullified them, and the LORD will release her.
NUM|30|13|Her husband may confirm or nullify any vow she makes or any sworn pledge to deny herself.
NUM|30|14|But if her husband says nothing to her about it from day to day, then he confirms all her vows or the pledges binding on her. He confirms them by saying nothing to her when he hears about them.
NUM|30|15|If, however, he nullifies them some time after he hears about them, then he is responsible for her guilt."
NUM|30|16|These are the regulations the LORD gave Moses concerning relationships between a man and his wife, and between a father and his young daughter still living in his house.
NUM|31|1|The LORD said to Moses,
NUM|31|2|"Take vengeance on the Midianites for the Israelites. After that, you will be gathered to your people."
NUM|31|3|So Moses said to the people, "Arm some of your men to go to war against the Midianites and to carry out the LORD's vengeance on them.
NUM|31|4|Send into battle a thousand men from each of the tribes of Israel."
NUM|31|5|So twelve thousand men armed for battle, a thousand from each tribe, were supplied from the clans of Israel.
NUM|31|6|Moses sent them into battle, a thousand from each tribe, along with Phinehas son of Eleazar, the priest, who took with him articles from the sanctuary and the trumpets for signaling.
NUM|31|7|They fought against Midian, as the LORD commanded Moses, and killed every man.
NUM|31|8|Among their victims were Evi, Rekem, Zur, Hur and Reba-the five kings of Midian. They also killed Balaam son of Beor with the sword.
NUM|31|9|The Israelites captured the Midianite women and children and took all the Midianite herds, flocks and goods as plunder.
NUM|31|10|They burned all the towns where the Midianites had settled, as well as all their camps.
NUM|31|11|They took all the plunder and spoils, including the people and animals,
NUM|31|12|and brought the captives, spoils and plunder to Moses and Eleazar the priest and the Israelite assembly at their camp on the plains of Moab, by the Jordan across from Jericho.
NUM|31|13|Moses, Eleazar the priest and all the leaders of the community went to meet them outside the camp.
NUM|31|14|Moses was angry with the officers of the army-the commanders of thousands and commanders of hundreds-who returned from the battle.
NUM|31|15|"Have you allowed all the women to live?" he asked them.
NUM|31|16|"They were the ones who followed Balaam's advice and were the means of turning the Israelites away from the LORD in what happened at Peor, so that a plague struck the LORD's people.
NUM|31|17|Now kill all the boys. And kill every woman who has slept with a man,
NUM|31|18|but save for yourselves every girl who has never slept with a man.
NUM|31|19|"All of you who have killed anyone or touched anyone who was killed must stay outside the camp seven days. On the third and seventh days you must purify yourselves and your captives.
NUM|31|20|Purify every garment as well as everything made of leather, goat hair or wood."
NUM|31|21|Then Eleazar the priest said to the soldiers who had gone into battle, "This is the requirement of the law that the LORD gave Moses:
NUM|31|22|Gold, silver, bronze, iron, tin, lead
NUM|31|23|and anything else that can withstand fire must be put through the fire, and then it will be clean. But it must also be purified with the water of cleansing. And whatever cannot withstand fire must be put through that water.
NUM|31|24|On the seventh day wash your clothes and you will be clean. Then you may come into the camp."
NUM|31|25|The LORD said to Moses,
NUM|31|26|"You and Eleazar the priest and the family heads of the community are to count all the people and animals that were captured.
NUM|31|27|Divide the spoils between the soldiers who took part in the battle and the rest of the community.
NUM|31|28|From the soldiers who fought in the battle, set apart as tribute for the LORD one out of every five hundred, whether persons, cattle, donkeys, sheep or goats.
NUM|31|29|Take this tribute from their half share and give it to Eleazar the priest as the LORD's part.
NUM|31|30|From the Israelites' half, select one out of every fifty, whether persons, cattle, donkeys, sheep, goats or other animals. Give them to the Levites, who are responsible for the care of the LORD's tabernacle."
NUM|31|31|So Moses and Eleazar the priest did as the LORD commanded Moses.
NUM|31|32|The plunder remaining from the spoils that the soldiers took was 675,000 sheep,
NUM|31|33|72,000 cattle,
NUM|31|34|61,000 donkeys
NUM|31|35|and 32,000 women who had never slept with a man.
NUM|31|36|The half share of those who fought in the battle was: 337,500 sheep,
NUM|31|37|of which the tribute for the LORD was 675;
NUM|31|38|36,000 cattle, of which the tribute for the LORD was 72;
NUM|31|39|30,500 donkeys, of which the tribute for the LORD was 61;
NUM|31|40|16,000 people, of which the tribute for the LORD was 32.
NUM|31|41|Moses gave the tribute to Eleazar the priest as the LORD's part, as the LORD commanded Moses.
NUM|31|42|The half belonging to the Israelites, which Moses set apart from that of the fighting men-
NUM|31|43|the community's half-was 337,500 sheep,
NUM|31|44|36,000 cattle,
NUM|31|45|30,500 donkeys
NUM|31|46|and 16,000 people.
NUM|31|47|From the Israelites' half, Moses selected one out of every fifty persons and animals, as the LORD commanded him, and gave them to the Levites, who were responsible for the care of the LORD's tabernacle.
NUM|31|48|Then the officers who were over the units of the army-the commanders of thousands and commanders of hundreds-went to Moses
NUM|31|49|and said to him, "Your servants have counted the soldiers under our command, and not one is missing.
NUM|31|50|So we have brought as an offering to the LORD the gold articles each of us acquired-armlets, bracelets, signet rings, earrings and necklaces-to make atonement for ourselves before the LORD."
NUM|31|51|Moses and Eleazar the priest accepted from them the gold-all the crafted articles.
NUM|31|52|All the gold from the commanders of thousands and commanders of hundreds that Moses and Eleazar presented as a gift to the LORD weighed 16,750 shekels.
NUM|31|53|Each soldier had taken plunder for himself.
NUM|31|54|Moses and Eleazar the priest accepted the gold from the commanders of thousands and commanders of hundreds and brought it into the Tent of Meeting as a memorial for the Israelites before the LORD.
NUM|32|1|The Reubenites and Gadites, who had very large herds and flocks, saw that the lands of Jazer and Gilead were suitable for livestock.
NUM|32|2|So they came to Moses and Eleazar the priest and to the leaders of the community, and said,
NUM|32|3|"Ataroth, Dibon, Jazer, Nimrah, Heshbon, Elealeh, Sebam, Nebo and Beon-
NUM|32|4|the land the LORD subdued before the people of Israel-are suitable for livestock, and your servants have livestock.
NUM|32|5|If we have found favor in your eyes," they said, "let this land be given to your servants as our possession. Do not make us cross the Jordan."
NUM|32|6|Moses said to the Gadites and Reubenites, "Shall your countrymen go to war while you sit here?
NUM|32|7|Why do you discourage the Israelites from going over into the land the LORD has given them?
NUM|32|8|This is what your fathers did when I sent them from Kadesh Barnea to look over the land.
NUM|32|9|After they went up to the Valley of Eshcol and viewed the land, they discouraged the Israelites from entering the land the LORD had given them.
NUM|32|10|The LORD's anger was aroused that day and he swore this oath:
NUM|32|11|'Because they have not followed me wholeheartedly, not one of the men twenty years old or more who came up out of Egypt will see the land I promised on oath to Abraham, Isaac and Jacob-
NUM|32|12|not one except Caleb son of Jephunneh the Kenizzite and Joshua son of Nun, for they followed the LORD wholeheartedly.'
NUM|32|13|The LORD's anger burned against Israel and he made them wander in the desert forty years, until the whole generation of those who had done evil in his sight was gone.
NUM|32|14|"And here you are, a brood of sinners, standing in the place of your fathers and making the LORD even more angry with Israel.
NUM|32|15|If you turn away from following him, he will again leave all this people in the desert, and you will be the cause of their destruction."
NUM|32|16|Then they came up to him and said, "We would like to build pens here for our livestock and cities for our women and children.
NUM|32|17|But we are ready to arm ourselves and go ahead of the Israelites until we have brought them to their place. Meanwhile our women and children will live in fortified cities, for protection from the inhabitants of the land.
NUM|32|18|We will not return to our homes until every Israelite has received his inheritance.
NUM|32|19|We will not receive any inheritance with them on the other side of the Jordan, because our inheritance has come to us on the east side of the Jordan."
NUM|32|20|Then Moses said to them, "If you will do this-if you will arm yourselves before the LORD for battle,
NUM|32|21|and if all of you will go armed over the Jordan before the LORD until he has driven his enemies out before him-
NUM|32|22|then when the land is subdued before the LORD, you may return and be free from your obligation to the LORD and to Israel. And this land will be your possession before the LORD.
NUM|32|23|"But if you fail to do this, you will be sinning against the LORD; and you may be sure that your sin will find you out.
NUM|32|24|Build cities for your women and children, and pens for your flocks, but do what you have promised."
NUM|32|25|The Gadites and Reubenites said to Moses, "We your servants will do as our lord commands.
NUM|32|26|Our children and wives, our flocks and herds will remain here in the cities of Gilead.
NUM|32|27|But your servants, every man armed for battle, will cross over to fight before the LORD, just as our lord says."
NUM|32|28|Then Moses gave orders about them to Eleazar the priest and Joshua son of Nun and to the family heads of the Israelite tribes.
NUM|32|29|He said to them, "If the Gadites and Reubenites, every man armed for battle, cross over the Jordan with you before the LORD, then when the land is subdued before you, give them the land of Gilead as their possession.
NUM|32|30|But if they do not cross over with you armed, they must accept their possession with you in Canaan."
NUM|32|31|The Gadites and Reubenites answered, "Your servants will do what the LORD has said.
NUM|32|32|We will cross over before the LORD into Canaan armed, but the property we inherit will be on this side of the Jordan."
NUM|32|33|Then Moses gave to the Gadites, the Reubenites and the half-tribe of Manasseh son of Joseph the kingdom of Sihon king of the Amorites and the kingdom of Og king of Bashan-the whole land with its cities and the territory around them.
NUM|32|34|The Gadites built up Dibon, Ataroth, Aroer,
NUM|32|35|Atroth Shophan, Jazer, Jogbehah,
NUM|32|36|Beth Nimrah and Beth Haran as fortified cities, and built pens for their flocks.
NUM|32|37|And the Reubenites rebuilt Heshbon, Elealeh and Kiriathaim,
NUM|32|38|as well as Nebo and Baal Meon (these names were changed) and Sibmah. They gave names to the cities they rebuilt.
NUM|32|39|The descendants of Makir son of Manasseh went to Gilead, captured it and drove out the Amorites who were there.
NUM|32|40|So Moses gave Gilead to the Makirites, the descendants of Manasseh, and they settled there.
NUM|32|41|Jair, a descendant of Manasseh, captured their settlements and called them Havvoth Jair.
NUM|32|42|And Nobah captured Kenath and its surrounding settlements and called it Nobah after himself.
NUM|33|1|Here are the stages in the journey of the Israelites when they came out of Egypt by divisions under the leadership of Moses and Aaron.
NUM|33|2|At the LORD's command Moses recorded the stages in their journey. This is their journey by stages:
NUM|33|3|The Israelites set out from Rameses on the fifteenth day of the first month, the day after the Passover. They marched out boldly in full view of all the Egyptians,
NUM|33|4|who were burying all their firstborn, whom the LORD had struck down among them; for the LORD had brought judgment on their gods.
NUM|33|5|The Israelites left Rameses and camped at Succoth.
NUM|33|6|They left Succoth and camped at Etham, on the edge of the desert.
NUM|33|7|They left Etham, turned back to Pi Hahiroth, to the east of Baal Zephon, and camped near Migdol.
NUM|33|8|They left Pi Hahiroth and passed through the sea into the desert, and when they had traveled for three days in the Desert of Etham, they camped at Marah.
NUM|33|9|They left Marah and went to Elim, where there were twelve springs and seventy palm trees, and they camped there.
NUM|33|10|They left Elim and camped by the Red Sea.
NUM|33|11|They left the Red Sea and camped in the Desert of Sin.
NUM|33|12|They left the Desert of Sin and camped at Dophkah.
NUM|33|13|They left Dophkah and camped at Alush.
NUM|33|14|They left Alush and camped at Rephidim, where there was no water for the people to drink.
NUM|33|15|They left Rephidim and camped in the Desert of Sinai.
NUM|33|16|They left the Desert of Sinai and camped at Kibroth Hattaavah.
NUM|33|17|They left Kibroth Hattaavah and camped at Hazeroth.
NUM|33|18|They left Hazeroth and camped at Rithmah.
NUM|33|19|They left Rithmah and camped at Rimmon Perez.
NUM|33|20|They left Rimmon Perez and camped at Libnah.
NUM|33|21|They left Libnah and camped at Rissah.
NUM|33|22|They left Rissah and camped at Kehelathah.
NUM|33|23|They left Kehelathah and camped at Mount Shepher.
NUM|33|24|They left Mount Shepher and camped at Haradah.
NUM|33|25|They left Haradah and camped at Makheloth.
NUM|33|26|They left Makheloth and camped at Tahath.
NUM|33|27|They left Tahath and camped at Terah.
NUM|33|28|They left Terah and camped at Mithcah.
NUM|33|29|They left Mithcah and camped at Hashmonah.
NUM|33|30|They left Hashmonah and camped at Moseroth.
NUM|33|31|They left Moseroth and camped at Bene Jaakan.
NUM|33|32|They left Bene Jaakan and camped at Hor Haggidgad.
NUM|33|33|They left Hor Haggidgad and camped at Jotbathah.
NUM|33|34|They left Jotbathah and camped at Abronah.
NUM|33|35|They left Abronah and camped at Ezion Geber.
NUM|33|36|They left Ezion Geber and camped at Kadesh, in the Desert of Zin.
NUM|33|37|They left Kadesh and camped at Mount Hor, on the border of Edom.
NUM|33|38|At the LORD's command Aaron the priest went up Mount Hor, where he died on the first day of the fifth month of the fortieth year after the Israelites came out of Egypt.
NUM|33|39|Aaron was a hundred and twenty-three years old when he died on Mount Hor.
NUM|33|40|The Canaanite king of Arad, who lived in the Negev of Canaan, heard that the Israelites were coming.
NUM|33|41|They left Mount Hor and camped at Zalmonah.
NUM|33|42|They left Zalmonah and camped at Punon.
NUM|33|43|They left Punon and camped at Oboth.
NUM|33|44|They left Oboth and camped at Iye Abarim, on the border of Moab.
NUM|33|45|They left Iyim and camped at Dibon Gad.
NUM|33|46|They left Dibon Gad and camped at Almon Diblathaim.
NUM|33|47|They left Almon Diblathaim and camped in the mountains of Abarim, near Nebo.
NUM|33|48|They left the mountains of Abarim and camped on the plains of Moab by the Jordan across from Jericho.
NUM|33|49|There on the plains of Moab they camped along the Jordan from Beth Jeshimoth to Abel Shittim.
NUM|33|50|On the plains of Moab by the Jordan across from Jericho the LORD said to Moses,
NUM|33|51|"Speak to the Israelites and say to them: 'When you cross the Jordan into Canaan,
NUM|33|52|drive out all the inhabitants of the land before you. Destroy all their carved images and their cast idols, and demolish all their high places.
NUM|33|53|Take possession of the land and settle in it, for I have given you the land to possess.
NUM|33|54|Distribute the land by lot, according to your clans. To a larger group give a larger inheritance, and to a smaller group a smaller one. Whatever falls to them by lot will be theirs. Distribute it according to your ancestral tribes.
NUM|33|55|"'But if you do not drive out the inhabitants of the land, those you allow to remain will become barbs in your eyes and thorns in your sides. They will give you trouble in the land where you will live.
NUM|33|56|And then I will do to you what I plan to do to them.'"
NUM|34|1|The LORD said to Moses,
NUM|34|2|"Command the Israelites and say to them: 'When you enter Canaan, the land that will be allotted to you as an inheritance will have these boundaries:
NUM|34|3|"'Your southern side will include some of the Desert of Zin along the border of Edom. On the east, your southern boundary will start from the end of the Salt Sea,
NUM|34|4|cross south of Scorpion Pass, continue on to Zin and go south of Kadesh Barnea. Then it will go to Hazar Addar and over to Azmon,
NUM|34|5|where it will turn, join the Wadi of Egypt and end at the Sea.
NUM|34|6|"'Your western boundary will be the coast of the Great Sea. This will be your boundary on the west.
NUM|34|7|"'For your northern boundary, run a line from the Great Sea to Mount Hor
NUM|34|8|and from Mount Hor to Lebo Hamath. Then the boundary will go to Zedad,
NUM|34|9|continue to Ziphron and end at Hazar Enan. This will be your boundary on the north.
NUM|34|10|"'For your eastern boundary, run a line from Hazar Enan to Shepham.
NUM|34|11|The boundary will go down from Shepham to Riblah on the east side of Ain and continue along the slopes east of the Sea of Kinnereth.
NUM|34|12|Then the boundary will go down along the Jordan and end at the Salt Sea. "'This will be your land, with its boundaries on every side.'"
NUM|34|13|Moses commanded the Israelites: "Assign this land by lot as an inheritance. The LORD has ordered that it be given to the nine and a half tribes,
NUM|34|14|because the families of the tribe of Reuben, the tribe of Gad and the half-tribe of Manasseh have received their inheritance.
NUM|34|15|These two and a half tribes have received their inheritance on the east side of the Jordan of Jericho, toward the sunrise."
NUM|34|16|The LORD said to Moses,
NUM|34|17|"These are the names of the men who are to assign the land for you as an inheritance: Eleazar the priest and Joshua son of Nun.
NUM|34|18|And appoint one leader from each tribe to help assign the land.
NUM|34|19|These are their names: Caleb son of Jephunneh, from the tribe of Judah;
NUM|34|20|Shemuel son of Ammihud, from the tribe of Simeon;
NUM|34|21|Elidad son of Kislon, from the tribe of Benjamin;
NUM|34|22|Bukki son of Jogli, the leader from the tribe of Dan;
NUM|34|23|Hanniel son of Ephod, the leader from the tribe of Manasseh son of Joseph;
NUM|34|24|Kemuel son of Shiphtan, the leader from the tribe of Ephraim son of Joseph;
NUM|34|25|Elizaphan son of Parnach, the leader from the tribe of Zebulun;
NUM|34|26|Paltiel son of Azzan, the leader from the tribe of Issachar;
NUM|34|27|Ahihud son of Shelomi, the leader from the tribe of Asher;
NUM|34|28|Pedahel son of Ammihud, the leader from the tribe of Naphtali."
NUM|34|29|These are the men the LORD commanded to assign the inheritance to the Israelites in the land of Canaan.
NUM|35|1|On the plains of Moab by the Jordan across from Jericho, the LORD said to Moses,
NUM|35|2|"Command the Israelites to give the Levites towns to live in from the inheritance the Israelites will possess. And give them pasturelands around the towns.
NUM|35|3|Then they will have towns to live in and pasturelands for their cattle, flocks and all their other livestock.
NUM|35|4|"The pasturelands around the towns that you give the Levites will extend out fifteen hundred feet from the town wall.
NUM|35|5|Outside the town, measure three thousand feet on the east side, three thousand on the south side, three thousand on the west and three thousand on the north, with the town in the center. They will have this area as pastureland for the towns.
NUM|35|6|"Six of the towns you give the Levites will be cities of refuge, to which a person who has killed someone may flee. In addition, give them forty-two other towns.
NUM|35|7|In all you must give the Levites forty-eight towns, together with their pasturelands.
NUM|35|8|The towns you give the Levites from the land the Israelites possess are to be given in proportion to the inheritance of each tribe: Take many towns from a tribe that has many, but few from one that has few."
NUM|35|9|Then the LORD said to Moses:
NUM|35|10|"Speak to the Israelites and say to them: 'When you cross the Jordan into Canaan,
NUM|35|11|select some towns to be your cities of refuge, to which a person who has killed someone accidentally may flee.
NUM|35|12|They will be places of refuge from the avenger, so that a person accused of murder may not die before he stands trial before the assembly.
NUM|35|13|These six towns you give will be your cities of refuge.
NUM|35|14|Give three on this side of the Jordan and three in Canaan as cities of refuge.
NUM|35|15|These six towns will be a place of refuge for Israelites, aliens and any other people living among them, so that anyone who has killed another accidentally can flee there.
NUM|35|16|"'If a man strikes someone with an iron object so that he dies, he is a murderer; the murderer shall be put to death.
NUM|35|17|Or if anyone has a stone in his hand that could kill, and he strikes someone so that he dies, he is a murderer; the murderer shall be put to death.
NUM|35|18|Or if anyone has a wooden object in his hand that could kill, and he hits someone so that he dies, he is a murderer; the murderer shall be put to death.
NUM|35|19|The avenger of blood shall put the murderer to death; when he meets him, he shall put him to death.
NUM|35|20|If anyone with malice aforethought shoves another or throws something at him intentionally so that he dies
NUM|35|21|or if in hostility he hits him with his fist so that he dies, that person shall be put to death; he is a murderer. The avenger of blood shall put the murderer to death when he meets him.
NUM|35|22|"'But if without hostility someone suddenly shoves another or throws something at him unintentionally
NUM|35|23|or, without seeing him, drops a stone on him that could kill him, and he dies, then since he was not his enemy and he did not intend to harm him,
NUM|35|24|the assembly must judge between him and the avenger of blood according to these regulations.
NUM|35|25|The assembly must protect the one accused of murder from the avenger of blood and send him back to the city of refuge to which he fled. He must stay there until the death of the high priest, who was anointed with the holy oil.
NUM|35|26|"'But if the accused ever goes outside the limits of the city of refuge to which he has fled
NUM|35|27|and the avenger of blood finds him outside the city, the avenger of blood may kill the accused without being guilty of murder.
NUM|35|28|The accused must stay in his city of refuge until the death of the high priest; only after the death of the high priest may he return to his own property.
NUM|35|29|"'These are to be legal requirements for you throughout the generations to come, wherever you live.
NUM|35|30|"'Anyone who kills a person is to be put to death as a murderer only on the testimony of witnesses. But no one is to be put to death on the testimony of only one witness.
NUM|35|31|"'Do not accept a ransom for the life of a murderer, who deserves to die. He must surely be put to death.
NUM|35|32|"'Do not accept a ransom for anyone who has fled to a city of refuge and so allow him to go back and live on his own land before the death of the high priest.
NUM|35|33|"'Do not pollute the land where you are. Bloodshed pollutes the land, and atonement cannot be made for the land on which blood has been shed, except by the blood of the one who shed it.
NUM|35|34|Do not defile the land where you live and where I dwell, for I, the LORD, dwell among the Israelites.'"
NUM|36|1|The family heads of the clan of Gilead son of Makir, the son of Manasseh, who were from the clans of the descendants of Joseph, came and spoke before Moses and the leaders, the heads of the Israelite families.
NUM|36|2|They said, "When the LORD commanded my lord to give the land as an inheritance to the Israelites by lot, he ordered you to give the inheritance of our brother Zelophehad to his daughters.
NUM|36|3|Now suppose they marry men from other Israelite tribes; then their inheritance will be taken from our ancestral inheritance and added to that of the tribe they marry into. And so part of the inheritance allotted to us will be taken away.
NUM|36|4|When the Year of Jubilee for the Israelites comes, their inheritance will be added to that of the tribe into which they marry, and their property will be taken from the tribal inheritance of our forefathers."
NUM|36|5|Then at the LORD's command Moses gave this order to the Israelites: "What the tribe of the descendants of Joseph is saying is right.
NUM|36|6|This is what the LORD commands for Zelophehad's daughters: They may marry anyone they please as long as they marry within the tribal clan of their father.
NUM|36|7|No inheritance in Israel is to pass from tribe to tribe, for every Israelite shall keep the tribal land inherited from his forefathers.
NUM|36|8|Every daughter who inherits land in any Israelite tribe must marry someone in her father's tribal clan, so that every Israelite will possess the inheritance of his fathers.
NUM|36|9|No inheritance may pass from tribe to tribe, for each Israelite tribe is to keep the land it inherits."
NUM|36|10|So Zelophehad's daughters did as the LORD commanded Moses.
NUM|36|11|Zelophehad's daughters-Mahlah, Tirzah, Hoglah, Milcah and Noah-married their cousins on their father's side.
NUM|36|12|They married within the clans of the descendants of Manasseh son of Joseph, and their inheritance remained in their father's clan and tribe.
NUM|36|13|These are the commands and regulations the LORD gave through Moses to the Israelites on the plains of Moab by the Jordan across from Jericho.
