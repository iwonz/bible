MARK|1|1|上帝的兒子 ，耶穌基督福音的起頭。
MARK|1|2|正如 以賽亞 先知書上記著： 「看哪，我要差遣我的使者在你面前， 他要為你預備道路。
MARK|1|3|在曠野有聲音呼喊著： 預備主的道， 修直他的路。」
MARK|1|4|照這話，施洗 約翰 來到曠野 ，宣講悔改的洗禮，使罪得赦。
MARK|1|5|猶太 全地和全 耶路撒冷 的人都出去，到 約翰 那裏，承認他們的罪，在 約旦河 裏受他的洗。
MARK|1|6|約翰 穿駱駝毛的衣服，腰束皮帶，吃的是蝗蟲和野蜜。
MARK|1|7|他宣講，說：「有一位在我以後來的，能力比我更大，我就是彎腰給他解鞋帶也不配。
MARK|1|8|我用水給你們施洗，他卻要用聖靈給你們施洗。」
MARK|1|9|那時，耶穌從 加利利 的 拿撒勒 來，在 約旦河 裏受了 約翰 的洗。
MARK|1|10|他從水裏一上來，就看見天裂開了，聖靈彷彿鴿子降在他身上。
MARK|1|11|又有聲音從天上來，說：「你是我的愛子，我喜愛你。」
MARK|1|12|聖靈立刻把耶穌催促到曠野裏去。
MARK|1|13|他在曠野四十天，受撒但的試探，並與野獸同在一起，且有天使來伺候他。
MARK|1|14|約翰 下監以後，耶穌來到 加利利 ，宣講上帝的福音，
MARK|1|15|說：「日期滿了，上帝的國近了。你們要悔改，信福音！」
MARK|1|16|耶穌沿著 加利利 的海邊走，看見 西門 和 西門 的弟弟 安得烈 在海上撒網；他們本是打魚的。
MARK|1|17|耶穌對他們說：「來跟從我，我要叫你們得人如得魚一樣。」
MARK|1|18|他們立刻捨了網，跟從他。
MARK|1|19|耶穌稍往前走，又見 西庇太 的兒子 雅各 和他弟弟 約翰 在船上補網。
MARK|1|20|耶穌隨即呼召他們，他們就把父親 西庇太 和雇工留在船上，跟從了耶穌。
MARK|1|21|他們到了 迦百農 ，耶穌就在安息日進了會堂教導人。
MARK|1|22|他們對他的教導感到很驚奇，因為他教導他們正像有權柄的人，不像文士。
MARK|1|23|當時，會堂裏有一個污靈附身的人，他在喊叫，
MARK|1|24|說：「 拿撒勒 人耶穌，你為甚麼干擾我們？你來消滅我們嗎？我知道你是誰，你是上帝的聖者。」
MARK|1|25|耶穌斥責他說：「不要作聲，從這人身上出來吧！」
MARK|1|26|污靈使那人抽了一陣風，大聲喊叫，就出來了。
MARK|1|27|眾人都驚訝，以致彼此對問：「這是甚麼事？是個新的教導啊！他用權柄命令污靈，連污靈也聽從了他。」
MARK|1|28|於是耶穌的名聲立刻傳遍了全 加利利 周圍地區。
MARK|1|29|他們一出會堂，就同 雅各 和 約翰 進了 西門 和 安得烈 的家。
MARK|1|30|西門 的岳母正發燒躺著，就有人告訴耶穌。
MARK|1|31|耶穌進前拉著她的手，扶她起來，燒就退了，於是她服事他們。
MARK|1|32|傍晚日落的時候，有人帶著一切害病的和被鬼附的，來到耶穌跟前。
MARK|1|33|全城的人都聚集在門前。
MARK|1|34|耶穌治好了許多害各樣病的人，又趕出許多鬼，不許鬼說話，因為鬼認識他。
MARK|1|35|次日早晨，天未亮的時候，耶穌起來，到曠野地方去，在那裏禱告。
MARK|1|36|西門 和同伴出去找他，
MARK|1|37|找到了就對他說：「眾人都在找你！」
MARK|1|38|耶穌對他們說：「讓我們往別處去，到鄰近的鄉村，我也好在那裏傳道，因為我是為這事出來的。」
MARK|1|39|於是他走遍全 加利利 ，在他們的會堂傳道，並且趕鬼。
MARK|1|40|有一個痲瘋病人來求耶穌，向他跪下 ，說：「你若肯，你能使我潔淨。」
MARK|1|41|耶穌動了慈心，就伸手摸他，說：「我肯，你潔淨了吧！」
MARK|1|42|痲瘋病立刻離開他，他就潔淨了。
MARK|1|43|耶穌嚴嚴地叮囑他，立刻打發他走，
MARK|1|44|對他說：「你要注意，千萬不可告訴任何人，只要去，讓祭司為你檢查，又因為你已經潔淨，獻上 摩西 所吩咐的祭物，作為證據給眾人看。」
MARK|1|45|那人出去，倒說許多的話，把這件事傳揚開了，使耶穌不能再公開進城，只好留在外邊曠野地方，人從各處都到他跟前來。
MARK|2|1|過了些日子，耶穌又進了 迦百農 。人聽說他在屋裏，
MARK|2|2|於是許多人聚集，甚至連門前都沒有空地；耶穌就對他們講道。
MARK|2|3|有人帶著一個癱子來見耶穌，是由四個人抬來的；
MARK|2|4|因為人多，無法抬到耶穌跟前，就把他所在那房子的屋頂拆了，既拆通了，就把癱子連所躺臥的褥子都縋下去。
MARK|2|5|耶穌見他們的信心，就對癱子說：「孩子，你的罪赦了。」
MARK|2|6|有幾個文士坐在那裏，心裏議論，說：
MARK|2|7|「這個人為甚麼這樣說呢？他說褻瀆的話了。除了上帝一位之外，誰能赦罪呢？」
MARK|2|8|耶穌心中立刻知道他們心裏這樣議論，就說：「你們心裏為甚麼這樣議論呢？
MARK|2|9|對癱子說『你的罪赦了』，或說『起來！拿你的褥子行走』，哪一樣容易呢？
MARK|2|10|但要讓你們知道，人子在地上有赦罪的權柄。」就對癱子說：
MARK|2|11|「我吩咐你，起來！拿你的褥子回家去吧。」
MARK|2|12|那人就起來，立刻拿著褥子，當著眾人面前出去了，以致眾人都驚奇，歸榮耀給上帝，說：「我們從來沒有見過這樣的事！」
MARK|2|13|耶穌又到海邊去，眾人都到他跟前來，他就教導他們。
MARK|2|14|耶穌往前走，看見 亞勒腓 的兒子 利未 在稅關坐著，就對他說：「來跟從我！」他就起來跟從耶穌。
MARK|2|15|耶穌在 利未 家裏坐席的時候，有好些稅吏和罪人與耶穌和他的門徒一同坐席，因為有很多人也跟隨耶穌。
MARK|2|16|法利賽人中的文士 看見耶穌與罪人和稅吏一同吃飯，就對他的門徒說：「他與稅吏和罪人一同吃飯嗎？」
MARK|2|17|耶穌聽見，就對他們說：「健康的人用不著醫生，有病的人才用得著。我不是來召義人，而是召罪人。」
MARK|2|18|那時， 約翰 的門徒和法利賽人都禁食。他們來問耶穌說：「 約翰 的門徒和法利賽人的門徒禁食，你的門徒卻不禁食，這是為甚麼呢？」
MARK|2|19|耶穌對他們說：「新郎和賓客在一起的時候，賓客怎麼能禁食呢？只要新郎和他們在一起，他們不能禁食。
MARK|2|20|但日子將到，新郎要被帶走，那日他們就要禁食了。
MARK|2|21|「沒有人把新布縫在舊衣服上，若是這樣，所補上的新布會撕破舊衣服，裂口就更大了。
MARK|2|22|也沒有人把新酒裝在舊皮袋裏，若是這樣，酒會脹破皮袋，酒和皮袋都糟蹋了 。相反地，新酒要裝在新皮袋裏 。」
MARK|2|23|有一個安息日，耶穌從麥田經過。他的門徒走路的時候，摘起麥穗來。
MARK|2|24|法利賽人對耶穌說：「看哪！他們為甚麼做安息日不合法的事呢？」
MARK|2|25|耶穌對他們說：「 大衛 和跟從他的人飢餓需要食物時所做的事，你們沒有念過嗎？
MARK|2|26|他在 亞比亞他 作大祭司的時候，怎麼進了上帝的居所，吃了供餅，又給跟從他的人吃呢？這餅除了祭司以外，人都不可以吃。」
MARK|2|27|他又對他們說：「安息日是為人設立的，人不是為安息日設立的。
MARK|2|28|所以，人子也是安息日的主。」
MARK|3|1|耶穌又進了會堂，在那裏有一個人，他的一隻手萎縮了。
MARK|3|2|眾人為了要控告耶穌，就窺探他會不會在安息日醫治那人。
MARK|3|3|耶穌對那手萎縮了的人說：「起來站在當中！」
MARK|3|4|他又問眾人：「在安息日行善行惡，救命害命，哪樣是合法的呢？」他們都不作聲。
MARK|3|5|耶穌怒目環視他們，因他們的心剛硬而憂傷，就對那人說：「伸出手來！」他把手一伸，手就復原了。
MARK|3|6|法利賽人出去，立刻同 希律 一黨的人商議怎樣除掉耶穌。
MARK|3|7|耶穌和門徒退到海邊去，有許多人從 加利利 跟隨他。還有許多人聽見他所做的事，就從 猶太 、 耶路撒冷 、 以土買 、 約旦河 的東邊，以及 推羅 和 西頓 的附近地方來到他那裏。
MARK|3|8|
MARK|3|9|因為人多，他吩咐門徒為他預備一隻小船，免得眾人擁擠他。
MARK|3|10|他治好了許多人，所以凡有疾病的，都擠著要摸他。
MARK|3|11|每當污靈看見他，就俯伏在他面前，喊著說：「你是上帝的兒子。」
MARK|3|12|耶穌再三囑咐他們不要把他宣揚出去。
MARK|3|13|耶穌上了山，把自己所要的人召來，他們就來到他那裏。
MARK|3|14|於是他設立十二個人，又稱他們為使徒 ，要他們常和自己同在，也要差他們去傳道，
MARK|3|15|並給他們權柄趕鬼。
MARK|3|16|他設立的十二個人 有 西門 －耶穌又給他起名叫 彼得 ，
MARK|3|17|還有 西庇太 的兒子 雅各 和 雅各 的弟弟 約翰 —耶穌又給他們起名叫 半尼其 ，就是雷的兒子—
MARK|3|18|又有 安得烈 、 腓力 、 巴多羅買 、 馬太 、 多馬 、 亞勒腓 的兒子 雅各 、 達太 和激進黨的 西門 ，
MARK|3|19|還有出賣耶穌的 加略 人 猶大 。
MARK|3|20|耶穌進了屋子，眾人又聚集，甚至他連飯也顧不得吃。
MARK|3|21|耶穌的家人聽見，就出來要拉住他，因為他們說他癲狂了。
MARK|3|22|從 耶路撒冷 下來的文士說：「他是被 別西卜 附身的」，又說：「他是靠著鬼王趕鬼的。」
MARK|3|23|耶穌叫他們來，用比喻對他們說：「撒但怎能趕出撒但呢？
MARK|3|24|一國若自相紛爭，那國就立不住；
MARK|3|25|一家若自相紛爭，那家就立不住。
MARK|3|26|撒但若自相攻打紛爭，他就立不住，必定滅亡。
MARK|3|27|沒有人能進壯士家裏，搶奪他的東西；除非先綁住那壯士，否則無法搶奪他的家。
MARK|3|28|我實在告訴你們，世人一切的罪和一切褻瀆的話都可以得到赦免；
MARK|3|29|凡褻瀆聖靈的，卻永不得赦免，而要擔當永遠的罪。」
MARK|3|30|因為他們說：「他是被污靈附身的。」
MARK|3|31|那時，耶穌的母親和他兄弟來，站在外邊，打發人去叫他。
MARK|3|32|有許多人在耶穌周圍坐著，他們就告訴他說：「看哪！你母親、你兄弟和你姊妹 在外邊找你。」
MARK|3|33|耶穌回答他們：「誰是我的母親？誰是我的兄弟？」
MARK|3|34|就環視那周圍坐著的人，說：「看哪，我的母親，我的兄弟！
MARK|3|35|凡遵行上帝旨意的人就是我的兄弟姊妹和母親。」
MARK|4|1|耶穌又在海邊教導人。有一大群人到他那裏聚集，他只好上船坐下。船在海裏，眾人都靠近海，站在岸上。
MARK|4|2|耶穌就用許多比喻教導他們。在教導的時候，他對他們說：
MARK|4|3|「你們聽啊，有一個撒種的出去撒種。
MARK|4|4|他撒的時候，有的落在路旁，飛鳥來把它吃掉了。
MARK|4|5|有的落在土淺的石頭地上，因為土不深，很快就長出苗來，
MARK|4|6|太陽出來一曬，因為沒有根就枯乾了。
MARK|4|7|有的落在荊棘裏，荊棘長起來，把它擠住了，就結不出果實。
MARK|4|8|又有的落在好土裏，就發芽長大，結出果實，有三十倍的，有六十倍的，有一百倍的。」
MARK|4|9|耶穌又說：「有耳可聽的，就應當聽！」
MARK|4|10|耶穌獨自一人的時候，跟隨他的人和十二使徒問他這些比喻的意思。
MARK|4|11|耶穌對他們說：「上帝國的奧祕只讓你們知道，若是對外人講，凡事就用比喻，
MARK|4|12|要 他們看了又看，卻看不清， 聽了又聽，卻不明白， 免得他們回轉過來，獲得赦免。」
MARK|4|13|耶穌又對他們說：「你們不明白這比喻嗎？這樣怎能明白一切的比喻呢？
MARK|4|14|撒種的人所撒的就是道。
MARK|4|15|那撒在路旁的種子，就是人聽了道，撒但立刻來，把撒在他們心裏的道奪了去。
MARK|4|16|那撒在石頭地上的，就是人聽了道，立刻歡喜領受，
MARK|4|17|因心裏沒有根，不過是暫時的，一旦為道遭受患難或迫害，立刻就跌倒。
MARK|4|18|還有那撒在荊棘裏的，就是人聽了道，
MARK|4|19|後來有世上的憂慮、錢財的迷惑，和別樣的私慾進來，把道擠住了，結不出果實。
MARK|4|20|那撒在好土裏的，就是人聽了道，領受了，並且結了果實，有三十倍的，有六十倍的，有一百倍的。」
MARK|4|21|耶穌又對他們說：「人拿燈來，難道是要放在斗底下，床底下，而不放在燈臺上嗎？
MARK|4|22|因為掩藏的事沒有不顯出來的，隱瞞的事也沒有不露出來的。
MARK|4|23|有耳可聽的，就應當聽！」
MARK|4|24|他又說：「你們要留心所聽的。你們用甚麼量器來量，也將要用甚麼來量給你們，並且要多給你們。
MARK|4|25|因為有的，還要給他；沒有的，連他所有的也要奪去。」
MARK|4|26|耶穌又說：「上帝的國如同人把種子撒在地上，
MARK|4|27|黑夜睡覺，白日起來，這種子就發芽生長，那人卻不知道如何會這樣。
MARK|4|28|土地自然而然地出產五穀，先發苗，後長穗，然後穗上結成飽滿的穀子。
MARK|4|29|五穀熟了，就用鐮刀去割，因為收成的時候到了。」
MARK|4|30|耶穌又說：「我們可用甚麼來比擬上帝的國呢？可用甚麼比喻來說明呢？
MARK|4|31|它像一粒芥菜種，種在地裏的時候，雖比地上所有的種子都小，
MARK|4|32|但種下去以後，它長起來，比各樣的菜都大，又長出大枝，以致天上的飛鳥可以在它的蔭下築巢。」
MARK|4|33|耶穌用許多這樣的比喻，照他們所能聽的，對他們講道；
MARK|4|34|若不用比喻，他就不對他們講，但私下沒有人的時候，就把一切的道講給門徒聽。
MARK|4|35|那天晚上，耶穌對門徒說：「我們渡到對岸去吧。」
MARK|4|36|門徒離開眾人，耶穌已在船上，他們就請他一同去；也有別的船和他同行。
MARK|4|37|忽然狂風大作，波浪打入船內，以致船灌滿了水。
MARK|4|38|耶穌在船尾上，枕著枕頭睡覺。門徒叫醒他，說：「老師！我們快沒命了，你不管嗎？」
MARK|4|39|耶穌醒了，斥責那風，向海說：「住了吧！靜了吧！」風就止住，大大平靜了。
MARK|4|40|耶穌對他們說：「為甚麼膽怯？你們還沒有信心嗎？」
MARK|4|41|他們就非常懼怕，彼此說：「這到底是誰？連風和海都聽從他。」
MARK|5|1|他們渡到海的對岸，到 格拉森 人 的地區。
MARK|5|2|耶穌一下船，就有一個污靈附身的人從墳墓迎著他走來。
MARK|5|3|那人常住在墳墓裏，沒有人能捆住他，就是用鐵鏈也不能；
MARK|5|4|因為人屢次用腳鐐和鐵鏈捆鎖他，鐵鏈被他掙斷，腳鐐也被他弄碎了，總沒有人能制伏他。
MARK|5|5|他晝夜常在墳墓裏和山中喊叫，又用石頭打自己。
MARK|5|6|他遠遠看見耶穌，就跑過來拜他，
MARK|5|7|大聲呼叫說：「至高上帝的兒子耶穌，你為甚麼干擾我？我指著上帝懇求你，不要叫我受苦！」
MARK|5|8|這是因耶穌曾吩咐他說：「污靈啊，從這人身上出來！」
MARK|5|9|耶穌問他：「你叫甚麼名字？」他說：「我名叫 群 ，因為我們數目眾多。」
MARK|5|10|他就再三求耶穌不要叫他們離開那地方。
MARK|5|11|在山坡那裏，有一大群豬正在吃食；
MARK|5|12|污靈就央求耶穌，說：「求你打發我們進入豬群，好附著牠們。」
MARK|5|13|耶穌准了他們，污靈就出來，進入豬裏，那群豬就闖下山崖，投進海裏，淹死了。豬的數目約有二千。
MARK|5|14|放豬的逃跑了，去告訴城裏和鄉下的人。眾人就來，要看發生了甚麼事。
MARK|5|15|他們來到耶穌那裏，看見那被鬼附的人，就是曾被群鬼所附的，坐著，穿著衣服，神智清醒，他們就害怕。
MARK|5|16|看見這事的人把被鬼附的人所遇見的，和那群豬的事，都告訴了眾人，
MARK|5|17|眾人就央求耶穌離開他們的地區。
MARK|5|18|耶穌上船的時候，那曾被鬼附的人懇求要和耶穌在一起。
MARK|5|19|耶穌不許，卻對他說：「你回家去，到你的親友那裏，將主為你所做多麼大的事和他怎樣憐憫你，都告訴他們。」
MARK|5|20|那人就走了，開始在 低加坡里 傳揚耶穌為他做了多麼大的事，眾人就都驚訝。
MARK|5|21|耶穌又坐船 渡到對岸，有一大群人聚集到他身邊；他正在海邊。
MARK|5|22|有一個會堂主管，名叫 葉魯 ，也來了，一見到耶穌，就俯伏在他腳前，
MARK|5|23|再三求他，說：「我的小女兒快要死了，求你去為她按手，使她痊癒，可以活下去。」
MARK|5|24|耶穌就和他同去。 有一大群人跟隨他，擁擠著他。
MARK|5|25|有一個女人，患了經血不止的病有十二年，
MARK|5|26|在好多醫生手裏受了許多苦，又花盡了她所有的，一點也不見好，反而更重了。
MARK|5|27|她聽見耶穌的事，就夾在眾人中間，從後面來摸耶穌的衣裳，
MARK|5|28|因她想：「我只摸到他的衣裳，就會痊癒。」
MARK|5|29|於是她的流血立刻止住，她覺得身上的疾病好了。
MARK|5|30|耶穌頓時心裏覺得有能力從自己身上出去，就在眾人中間轉過來，說：「誰摸我的衣裳？」
MARK|5|31|門徒對他說：「你看眾人擁擠著你，還說『誰摸我』呢？」
MARK|5|32|耶穌周圍觀看，要見做這事的女人。
MARK|5|33|那女人知道在自己身上所成的事，就恐懼戰兢，來俯伏在耶穌跟前，將實情全告訴他。
MARK|5|34|耶穌對她說：「女兒，你的信救了你，平安地回去吧！你的疾病痊癒了。」
MARK|5|35|耶穌還在說話的時候，有人從會堂主管的家裏來，說：「你的女兒死了，何必還勞駕老師呢？」
MARK|5|36|耶穌不理會他們所說的話，就對會堂主管說：「不要怕，只要信！」
MARK|5|37|於是他帶著 彼得 、 雅各 和 雅各 的弟弟 約翰 同去，不許別人跟著他。
MARK|5|38|他們來到會堂主管的家裏，耶穌看到一片吵鬧，並有人大聲哭泣哀號，
MARK|5|39|就進到裏面，對他們說：「為甚麼大吵大哭呢？孩子不是死了，是睡著了。」
MARK|5|40|他們就嘲笑耶穌。耶穌把他們都趕出去，帶著孩子的父母和跟隨的人進了孩子所在的地方，
MARK|5|41|就拉著孩子的手，對她說：「大利大，古米！」翻出來就是說：「女孩，我吩咐你，起來！」
MARK|5|42|那女孩子立刻起來走動—她已經十二歲了；他們就非常驚奇。
MARK|5|43|耶穌切切地囑咐他們，不要讓人知道這事，又吩咐給她東西吃。
MARK|6|1|耶穌離開那裏，來到自己的家鄉；門徒也跟從他。
MARK|6|2|到了安息日，他在會堂裏教導人。眾人聽見，就很驚奇，說：「這人哪來這本事呢？所賜給他的是甚麼智慧？他手所做的是何等的異能呢？
MARK|6|3|這不是那木匠嗎？不是 馬利亞 的兒子 雅各 、 約西 、 猶大 、 西門 的長兄嗎？他姊妹們不也是在我們這裏嗎？」他們就厭棄他。
MARK|6|4|耶穌對他們說：「先知除了在本鄉、本族和自己的家之外，沒有不被尊敬的。」
MARK|6|5|耶穌在那裏不能行甚麼異能，不過為幾個病人按手，治好他們。
MARK|6|6|他也詫異他們不信。 耶穌走遍周圍鄉村教導人。
MARK|6|7|他叫了十二個使徒來，差遣他們兩個兩個地出去，也賜給他們權柄制伏污靈，
MARK|6|8|並且吩咐他們：途中不要帶食物和行囊，腰袋裏也不要帶錢，除了手杖以外，甚麼都不要帶；
MARK|6|9|只要穿鞋子，也不要穿兩件內衣。
MARK|6|10|他又對他們說：「你們無論到何處，進哪家，就住在哪裏，直到離開那地方。
MARK|6|11|若有甚麼地方的人不接待你們，不聽你們，你們離開那裏的時候，要跺掉你們腳上的塵土，證明他們的不是。」
MARK|6|12|使徒就出去傳道，叫人悔改，
MARK|6|13|又趕出許多鬼，用油抹了許多病人，治好他們。
MARK|6|14|耶穌的名聲傳開了， 希律 王也聽見。有人說：「施洗的 約翰 從死人中復活了，因此才有這些異能在他裏面運行。」
MARK|6|15|但別人說：「他是 以利亞 。」又有人說：「是先知，正如先知中的一位。」
MARK|6|16|希律 聽見卻說：「是我所斬的 約翰 ，他復活了。」
MARK|6|17|原來， 希律 為他兄弟 腓力 的妻子 希羅底 的緣故，派人去抓了 約翰 ，把他綁了在監獄裏，因為 希律 已經娶了那婦人。
MARK|6|18|約翰 曾對 希律 說：「你佔有你兄弟的妻子是不合法的。」
MARK|6|19|於是 希羅底 懷恨他，想要殺他，只是不能。
MARK|6|20|因為 希律 怕 約翰 ，知道他是義人，是聖人，所以就保護他，雖然聽了他的講論十分困惑 ，仍然樂意聽他。
MARK|6|21|有一天，恰巧是 希律 的生日， 希律 擺設宴席，請了大臣、千夫長和 加利利 的領袖。
MARK|6|22|他的女兒 希羅底 進來跳舞，使 希律 和同席的人都很高興。王就對女孩說：「無論你要甚麼，向我求，我都會給你」；
MARK|6|23|又對她多次 起誓說：「無論你向我求甚麼，就是我國家的一半，我也會給你。」
MARK|6|24|她就出去對她母親說：「我該求甚麼呢？」她母親說：「施洗 約翰 的頭。」
MARK|6|25|她就急忙進去見王，求他說：「我願王立刻把施洗 約翰 的頭放在盤子裏給我。」
MARK|6|26|王就很憂愁，然而因他所發的誓，又因同席的人，不願食言，
MARK|6|27|就立刻派一個衛兵，吩咐拿 約翰 的頭來。衛兵就去，在監獄裏斬了 約翰 ，
MARK|6|28|把頭放在盤子裏，拿來給那女孩，她就給她母親。
MARK|6|29|約翰 的門徒聽到了，就來把他的屍體領去，放在墳墓裏。
MARK|6|30|使徒們聚集到耶穌那裏，把一切所做的事、所傳的道全告訴他。
MARK|6|31|他就說：「你們來，同我私下到荒野的地方去歇一歇。」這是因為來往的人多，他們連吃飯的時間也沒有。
MARK|6|32|他們就坐船，私下往荒野的地方去。
MARK|6|33|眾人看見他們走了，有許多認識他們的，就從各城步行，一同跑到那裏，比他們先趕到了。
MARK|6|34|耶穌出來，見有一大群的人，就憐憫他們，因為他們如同羊沒有牧人一般，於是開始教導他們許多事。
MARK|6|35|天已經很晚，門徒進前來，說：「這地方偏僻，而且天已經很晚了，
MARK|6|36|請叫眾人散去，他們好往四面的鄉鎮村莊去，自己買些東西吃。」
MARK|6|37|耶穌回答他們說：「你們給他們吃吧！」門徒對他說：「我們要拿兩百個銀幣去買餅給他們吃嗎？」
MARK|6|38|耶穌說：「你們有多少餅？去看看。」他們知道後就說：「有五個，還有兩條魚。」
MARK|6|39|耶穌吩咐他們，叫眾人一組一組地坐在青草地上。
MARK|6|40|眾人就一群一群地坐下，有一百的，有五十的。
MARK|6|41|耶穌拿著這五個餅和兩條魚，望著天祝福，擘開餅，遞給門徒，擺在眾人面前，也把那兩條魚分給眾人。
MARK|6|42|他們都吃，並且吃飽了。
MARK|6|43|門徒把餅和魚的碎屑收拾起來，裝滿了十二個籃子。
MARK|6|44|吃餅的男人共有五千。
MARK|6|45|耶穌隨即催門徒上船，先渡到對岸，到 伯賽大 去，等他叫眾人散去。
MARK|6|46|他辭別了他們，就往山上去禱告。
MARK|6|47|到了晚上，船在海中，耶穌獨自在岸上。
MARK|6|48|他看見門徒因風不順，搖櫓很苦。天快亮的時候，他在海面上走，往他們那裏去，想要超過他們。
MARK|6|49|但門徒看見他在海面上走，以為是鬼怪，就喊叫起來；
MARK|6|50|因為他們都看見了他，甚為驚慌。耶穌連忙對他們說：「放心！是我，不要怕！」
MARK|6|51|於是他到他們那裏，一上船，風就停了；他們心裏十分驚奇。
MARK|6|52|這是因為他們不明白那分餅的事，心裏還是愚頑。
MARK|6|53|他們渡過了海，在 革尼撒勒 靠岸，泊了船，
MARK|6|54|他們一下來，眾人立刻認出是耶穌，
MARK|6|55|就跑遍那整個地區，聽到他在哪裏，就把有病的人用褥子抬到哪裏。
MARK|6|56|耶穌所到的地方，或村中、或城裏、或鄉間，他們都把病人放在街市上，求耶穌讓他們摸一摸他的衣裳繸子，摸著的人就都好了。
MARK|7|1|有法利賽人和幾個從 耶路撒冷 來的文士聚集到耶穌那裏。
MARK|7|2|他們曾看見他的門徒中有人用不潔淨的手，就是沒有洗的手吃飯。
MARK|7|3|法利賽人和所有的 猶太 人都拘守古人的傳統，若不按規矩洗手就不吃飯；
MARK|7|4|從市場來，若不洗淨也不吃飯；他們還拘守好些別的規矩，如洗杯、罐、銅器、床鋪 等。
MARK|7|5|法利賽人和文士問他說：「你的門徒為甚麼不照古人的傳統，竟然用不潔淨的手吃飯呢？」
MARK|7|6|耶穌對他們說：「 以賽亞 指著你們假冒為善的人所預言的說得好。如經上所記： 『這百姓用嘴唇尊敬我， 他們的心卻遠離我。
MARK|7|7|他們把人的規條當作教義教導人； 他們拜我也是枉然。』
MARK|7|8|你們是離棄上帝的誡命，拘守人的傳統。」
MARK|7|9|耶穌又說：「你們誠然是廢棄上帝的誡命，為要守自己的傳統。
MARK|7|10|摩西 說：『當孝敬父母』；又說：『咒罵父母的，必須處死。』
MARK|7|11|你們倒說：『人若對父母說：我所當供奉你的已經作了各耳板』（各耳板就是奉獻的意思），
MARK|7|12|你們就容許他不必再奉養父母。
MARK|7|13|這就是你們藉著繼承傳統，廢了上帝的話。你們還做許多這樣的事。」
MARK|7|14|耶穌又叫眾人來，對他們說：「你們都要聽我的話，也要明白。
MARK|7|15|從外面進去的不能玷污人，惟有從裏面出來的才玷污人。 」
MARK|7|16|
MARK|7|17|耶穌離開眾人，進了屋子，門徒就問他這比喻的意思。
MARK|7|18|耶穌對他們說：「你們也是這樣不明白嗎？難道你們不了解，凡從外面進去的不能玷污人嗎？
MARK|7|19|因為不是進入他的心，而是進入他的肚子，又排入廁所。」（這是說，各樣的食物都是潔淨的。）
MARK|7|20|耶穌又說：「從人裏面出來的，那才玷污人；
MARK|7|21|因為從人心裏發出種種惡念，如淫亂、偷盜、兇殺、
MARK|7|22|姦淫、貪婪、邪惡、詭詐、淫蕩、嫉妒、毀謗、驕傲、狂妄。
MARK|7|23|這一切的惡都是從裏面出來，且能玷污人。」
MARK|7|24|耶穌從那裏起身，往 推羅 境內去，進了一家，他不願意人知道，卻隱藏不住。
MARK|7|25|立刻有一個婦人，她的小女兒被污靈附著，一聽見耶穌的事，就來俯伏在他腳前。
MARK|7|26|這婦人是 希臘 人，屬 敘利亞 的 腓尼基 族。她求耶穌從她女兒身上趕出那鬼。
MARK|7|27|耶穌對她說：「讓孩子們先吃飽，拿孩子的餅丟給小狗吃是不妥的。」
MARK|7|28|婦人回答：「主啊，桌子底下的小狗也吃小孩子的碎屑呀！」
MARK|7|29|耶穌對她說：「憑著這句話，你回去吧，鬼已經離開你的女兒了。」
MARK|7|30|她就回家去，見小孩子躺在床上，鬼已經出去了。
MARK|7|31|耶穌又離開了 推羅 地區，經過 西頓 ，就從 低加坡里 境內來到 加利利海 。
MARK|7|32|有人帶著一個耳聾舌結的人來見耶穌，求他為他按手。
MARK|7|33|耶穌領他離開眾人，到一邊去，就用指頭探他的耳朵，吐唾沫抹他的舌頭，
MARK|7|34|望天嘆息，對他說：「以法大！」就是說「開了吧！」
MARK|7|35|他的耳朵立刻 開了，舌結也解了，他說話也清楚了。
MARK|7|36|耶穌囑咐他們不要告訴人；但他越囑咐，他們越發傳揚。
MARK|7|37|眾人分外驚奇，說：「他所做的事樣樣都好，他甚至使聾子聽見，啞巴說話。」
MARK|8|1|那時，又有一大群人聚集，沒有甚麼吃的。耶穌叫門徒來，說：
MARK|8|2|「我憐憫這群人，因為他們同我在這裏已經三天，沒有吃的東西了。
MARK|8|3|我若叫他們餓著回家，他們會在路上餓昏，因為其中有從遠處來的。」
MARK|8|4|門徒回答：「在這野地，從哪裏能得餅使這些人吃飽呢？」
MARK|8|5|耶穌問他們：「你們有多少餅？」他們說：「七個。」
MARK|8|6|他吩咐眾人坐在地上，就拿著這七個餅祝謝了，擘開，遞給門徒，叫他們擺開，門徒就擺在眾人面前。
MARK|8|7|他們還有幾條小魚；耶穌祝謝了，就吩咐也擺在眾人面前。
MARK|8|8|他們都吃，並且吃飽了，收拾剩下的碎屑，有七筐子。
MARK|8|9|人數約有四千。耶穌打發他們走了，
MARK|8|10|隨即同門徒上船，來到 大瑪努他 境內。
MARK|8|11|法利賽人出來盤問耶穌，要求他從天上顯個神蹟給他們看，想要試探他。
MARK|8|12|耶穌心裏深深嘆息，說：「這世代為甚麼求神蹟呢？我實在告訴你們，沒有神蹟給這世代看。」
MARK|8|13|他就離開他們，又上船往海的對岸去了。
MARK|8|14|門徒忘了帶餅，在船上除了一個餅，沒有別的食物。
MARK|8|15|耶穌囑咐他們說：「你們要謹慎，要防備法利賽人的酵和 希律 的酵。」
MARK|8|16|他們彼此議論說：「這是因為我們沒有餅吧。」
MARK|8|17|耶穌知道了，就說：「你們為甚麼因為沒有餅就議論呢？你們還不領悟，還不明白嗎？你們的心還是愚頑嗎？
MARK|8|18|你們有眼睛，看不見嗎？有耳朵，聽不到嗎？也不記得嗎？
MARK|8|19|我擘開那五個餅分給五千人，你們收拾的碎屑裝滿了多少個籃子呢？」他們說：「十二個。」
MARK|8|20|「又擘開那七個餅分給四千人，你們收拾的碎屑裝滿了多少個筐子呢？」他們說：「七個。」
MARK|8|21|耶穌說：「你們還不明白嗎？」
MARK|8|22|他們來到 伯賽大 ，有人帶一個盲人來，求耶穌摸他。
MARK|8|23|耶穌拉著盲人的手，領他到村外，就吐唾沫在他眼睛上，為他按手，問他：「你看見甚麼？」
MARK|8|24|他抬頭一看，說：「我看見人，他們好像樹木，並且行走。」
MARK|8|25|隨後耶穌又按手在他眼睛上，他定睛一看，就復原了，樣樣都看得清楚了。
MARK|8|26|耶穌打發他回家，說：「連這村子你也不要進去。」
MARK|8|27|耶穌和門徒出去，往 凱撒利亞．腓立比 附近的村莊去。在路上，他問門徒：「人們說我是誰？」
MARK|8|28|他們對他說：「是施洗的 約翰 ；有人說是 以利亞 ；又有人說是先知中的一位。」
MARK|8|29|他又問他們：「你們說我是誰？」 彼得 回答他：「你是基督。」
MARK|8|30|於是耶穌切切地囑咐他們不可對任何人說起他。
MARK|8|31|從此，他教導他們說：「人子必須受許多的苦，被長老、祭司長和文士棄絕，並且被殺，三天後復活。」
MARK|8|32|耶穌明白地說了這話， 彼得 就拉著他，責備他。
MARK|8|33|耶穌轉過來看著門徒，斥責 彼得 說：「撒但，退到我後邊去！因為你不體會上帝的心意，而是體會人的意思。」
MARK|8|34|於是他叫眾人和門徒來，對他們說：「若有人要跟從我，就當捨己，背起自己的十字架來跟從我。
MARK|8|35|因為凡要救自己生命的，必喪失生命；凡為我和福音喪失生命的，必救自己的生命。
MARK|8|36|人就是賺得全世界，賠上自己的生命，有甚麼益處呢？
MARK|8|37|人還能拿甚麼換生命呢？
MARK|8|38|凡在這淫亂罪惡的世代，把我和我的道當作可恥的，人子在他父的榮耀裏與聖天使一同來臨的時候，也要把那人當作可恥的。」
MARK|9|1|耶穌又對他們說：「我實在告訴你們，站在這裏的，有人在沒經歷死亡以前，必定看見上帝的國帶著能力臨到。」
MARK|9|2|過了六天，耶穌帶著 彼得 、 雅各 、 約翰 ，領他們悄悄地上了高山。他在他們面前變了形像，
MARK|9|3|衣服放光，極其潔白，地上漂布的人沒有一個能漂得那樣白。
MARK|9|4|有 以利亞 和 摩西 向他們顯現，並且與耶穌說話。
MARK|9|5|彼得 對耶穌說：「拉比 ，我們在這裏真好！我們來搭三座棚，一座為你，一座為 摩西 ，一座為 以利亞 。」
MARK|9|6|彼得 不知道說甚麼才好，因為他們很害怕。
MARK|9|7|有一朵雲彩來遮蓋他們，又有聲音從雲彩裏出來，說：「這是我的愛子，你們要聽從他！」
MARK|9|8|門徒連忙向周圍觀看，不再看見任何人，只見耶穌同他們在一起。
MARK|9|9|下山的時候，耶穌囑咐他們說：「人子還沒有從死人中復活，你們不要把所看到的告訴人。」
MARK|9|10|門徒將這話存記在心，彼此議論「從死人中復活」是甚麼意思。
MARK|9|11|他們就問耶穌：「文士為甚麼說 以利亞 必須先來？」
MARK|9|12|耶穌說：「 以利亞 的確先來復興萬事。經上不是指著人子說，他要受許多的苦和被人輕慢嗎？
MARK|9|13|我告訴你們， 以利亞 已經來了，他們任意待他，正如經上指著他說的。」
MARK|9|14|他們到了門徒那裏，看見有一大群人圍著他們，又有文士和他們辯論。
MARK|9|15|眾人一見耶穌，都很驚奇，就跑上去向他問安。
MARK|9|16|耶穌問他們：「你們和他們辯論甚麼？」
MARK|9|17|眾人中的一個回答：「老師，我帶了我的兒子到你這裏來，他被啞巴的靈附著。
MARK|9|18|無論在哪裏，那靈拿住他，把他摔倒，他就口吐白沫，牙關緊鎖，身體僵硬。我請過你的門徒把那靈趕出去，他們卻不能。」
MARK|9|19|耶穌回答：「唉！這不信的世代啊，我和你們在一起要到幾時呢？我忍耐你們要到幾時呢？把他帶到我這裏！」
MARK|9|20|他們就帶了他來。那靈一見耶穌，就使他重重地抽風，倒在地上，翻來覆去，口吐白沫。
MARK|9|21|耶穌問他父親：「他得這病有多久了呢？」父親說：「從小的時候。
MARK|9|22|那靈屢次把他扔在火裏、水裏，要治死他。你若能做甚麼，求你憐憫我們，幫助我們。」
MARK|9|23|耶穌對他說：「『你若能』，在信的人，凡事都能。」
MARK|9|24|孩子的父親立刻喊著說：「我信；求你幫助我的不信！」
MARK|9|25|耶穌看見眾人都跑上來，就斥責那污靈說：「你這聾啞的靈，我命令你從他裏頭出來，再不要進去！」
MARK|9|26|那靈大喊一聲，使孩子猛烈地抽了一陣風，就出來了。孩子好像死了一般，以致眾人多半說：「他死了。」
MARK|9|27|但耶穌拉著他的手，扶他起來，他就站起來了。
MARK|9|28|耶穌進了屋子，門徒就私下問他：「我們為甚麼不能趕出那靈呢？」
MARK|9|29|耶穌對他們說：「非用禱告 ，這一類的邪靈總趕不出來。」
MARK|9|30|他們離開那地方，經過 加利利 ；耶穌不願意人知道，
MARK|9|31|因為他正教導門徒說：「人子將要被交在人手裏，他們要殺害他；被殺以後，三天後他要復活。」
MARK|9|32|門徒卻不明白這話，又不敢問他。
MARK|9|33|他們來到 迦百農 。耶穌在屋裏問門徒說：「你們在路上議論的是甚麼？」
MARK|9|34|門徒不作聲，因為他們在路上彼此爭論誰最大。
MARK|9|35|耶穌坐下，叫十二個使徒來，說：「若有人願意為首，他要作眾人之後，作眾人的用人。」
MARK|9|36|於是耶穌領一個小孩過來，讓他站在門徒當中，又抱起他來，對他們說：
MARK|9|37|「凡為我的名接納一個像這小孩子的，就是接納我；凡接納我的，不是接納我，而是接納那差我來的。」
MARK|9|38|約翰 對耶穌說：「老師，我們看見一個人奉你的名趕鬼，我們就阻止他，因為他不跟從我們。」
MARK|9|39|耶穌說：「不要阻止他，因為沒有人奉我的名行異能，反倒輕易毀謗我。
MARK|9|40|不抵擋我們的，就是幫助我們的。
MARK|9|41|凡因你們是屬基督，給你們一杯水喝的，我實在告訴你們，他一定會得到賞賜。」
MARK|9|42|「凡使這些信我的小子 中的一個跌倒的，倒不如把大磨石拴在這人的頸項上，扔在海裏。
MARK|9|43|如果你一隻手使你跌倒，就把它砍下來；你缺一隻手進入永生，比有兩隻手落到地獄，入那不滅的火裏去還好。
MARK|9|44|
MARK|9|45|如果你一隻腳使你跌倒，就把它砍下來；你瘸腿進入永生，比有兩隻腳被扔進地獄裏還好。
MARK|9|46|
MARK|9|47|如果你一隻眼使你跌倒，就去掉它；你只有一隻眼進入上帝的國，比有兩隻眼被扔進地獄裏還好。
MARK|9|48|在那裏，蟲是不死的，火是不滅的。
MARK|9|49|因為每個人必被火像鹽一般醃起來。
MARK|9|50|鹽本是好的，若失了鹹味，你們怎能用它調味呢？你們中間要有鹽，彼此和睦。」
MARK|10|1|耶穌從那裏起身，來到 猶太 的境內， 約旦河 的東邊。眾人又聚集到他那裏，他又照常教導他們。
MARK|10|2|有法利賽人來問他說：「男人休妻合不合法？」意思是要試探他。
MARK|10|3|耶穌回答他們說：「 摩西 吩咐你們的是甚麼？」
MARK|10|4|他們說：「 摩西 准許寫了休書就可以休妻。」
MARK|10|5|耶穌對他們說：「 摩西 因為你們的心硬，所以寫這誡命給你們。
MARK|10|6|但從起初創造的時候，上帝造人是造男造女。
MARK|10|7|因此，人要離開他的父母，與妻子結合 ，
MARK|10|8|二人成為一體。既然如此，夫妻不再是兩個人，而是一體的了。
MARK|10|9|所以，上帝配合的，人不可分開。」
MARK|10|10|他們到了屋裏，門徒又問他這事。
MARK|10|11|耶穌對他們說：「凡休妻另娶的，就是犯姦淫，辜負他的妻子；
MARK|10|12|妻子若離棄丈夫另嫁，也是犯姦淫了。」
MARK|10|13|有人帶著小孩子來見耶穌，要他摸他們，門徒就責備那些人。
MARK|10|14|耶穌看見就很生氣，對門徒說：「讓小孩到我這裏來，不要阻止他們，因為在上帝國的正是這樣的人。
MARK|10|15|我實在告訴你們，凡要接受上帝國的，若不像小孩子，絕不能進去。」
MARK|10|16|於是他抱著小孩子，給他們按手，為他們祝福。
MARK|10|17|耶穌剛上路的時候，有一個人跑來，跪在他面前，問他：「善良的老師，我該做甚麼事才能承受永生？」
MARK|10|18|耶穌對他說：「你為甚麼稱我是善良的？除了上帝一位之外，再沒有善良的。
MARK|10|19|誡命你是知道的：『不可殺人；不可姦淫；不可偷盜；不可作假見證；不可虧負人；當孝敬父母。』」
MARK|10|20|他對耶穌說：「老師，這一切我從小都遵守了。」
MARK|10|21|耶穌看著他，就愛他，對他說：「你還缺少一件：去變賣你所有的，分給窮人，就必有財寶在天上；然後來跟從我。」
MARK|10|22|他聽見這話，臉就變了色，憂憂愁愁地走了，因為他的產業很多。
MARK|10|23|耶穌看了看周圍，對門徒說：「有錢財的人進上帝的國是何等的難哪！」
MARK|10|24|門徒對他的話非常驚奇。耶穌又對他們說：「孩子們， 要進上帝的國是何等的難哪！
MARK|10|25|駱駝穿過針眼比財主進上帝的國還容易呢！」
MARK|10|26|門徒就更為驚訝，彼此對問：「這樣，誰能得救呢？」
MARK|10|27|耶穌看著他們，說：「在人不能，在上帝卻不然，因為在上帝凡事都能。」
MARK|10|28|彼得 就對他說：「看哪，我們已經撇下一切跟從你了。」
MARK|10|29|耶穌說：「我實在告訴你們，凡為我和福音撇下房屋，或是兄弟、姊妹、父親、母親、兒女、田地，
MARK|10|30|沒有不在今世得百倍的，就是房屋、兄弟、姊妹、母親、兒女、田地，並且要受迫害，在來世得永生。
MARK|10|31|然而，有許多在前的，將要在後；在後的，將要在前。」
MARK|10|32|他們行路上 耶路撒冷 去。耶穌在前頭走，他們很驚訝，跟從的人也害怕。耶穌又叫十二使徒來，把自己將要遭遇的事告訴他們，
MARK|10|33|說：「看哪，我們上 耶路撒冷 去，人子將被交給祭司長和文士；他們要定他死罪，又交給外邦人。
MARK|10|34|他們要戲弄他，向他吐唾沫，鞭打他，殺害他；三天後，他要復活。」
MARK|10|35|西庇太 的兒子 雅各 和 約翰 進前來，對耶穌說：「老師，我們無論求你甚麼，願你為我們做。」
MARK|10|36|耶穌對他們說：「要我為你們做甚麼？」
MARK|10|37|他們對他說：「在你的榮耀裏，請賜我們一個坐在你右邊，一個坐在你左邊。」
MARK|10|38|耶穌對他們說：「你們不知道所求的是甚麼。我所喝的杯，你們能喝嗎？我所受的洗，你們能受嗎？」
MARK|10|39|他們對他說：「我們能。」耶穌對他們說：「我所喝的杯，你們要喝；我所受的洗，你們也要受。
MARK|10|40|可是坐在我的左右，不是我可以賜的，而是為誰預備就賜給誰。」
MARK|10|41|其餘十個門徒聽見，就對 雅各 和 約翰 很生氣。
MARK|10|42|耶穌叫了他們來，對他們說：「你們知道，外邦人有君王作主治理他們，有大臣操權管轄他們。
MARK|10|43|但是在你們中間，不可這樣。你們中間誰願為大，就要作你們的用人；
MARK|10|44|在你們中間誰願為首，就要作眾人的僕人。
MARK|10|45|因為人子來，並不是要受人的服事，乃是要服事人，並且要捨命作多人的贖價。」
MARK|10|46|他們到了 耶利哥 。耶穌同門徒並許多人離開 耶利哥 的時候，有一個討飯的盲人，是 底買 的兒子 巴底買 ，坐在路旁。
MARK|10|47|他聽見是 拿撒勒 的耶穌，就喊了起來，說：「 大衛 之子耶穌啊，可憐我吧！」
MARK|10|48|有許多人責備他，不許他作聲，他卻越發喊著：「 大衛 之子啊，可憐我吧！」
MARK|10|49|耶穌就站住，說：「叫他過來。」他們就叫那盲人，對他說：「放心，起來！他在叫你啦。」
MARK|10|50|盲人就丟下衣服，跳起來，走到耶穌那裏。
MARK|10|51|耶穌回答他說：「你要我為你做甚麼？」盲人對他說：「拉波尼 ，我要能看見。」
MARK|10|52|耶穌對他說：「你去吧！你的信救了你。」盲人立刻看得見，就在路上跟隨耶穌。
MARK|11|1|耶穌和門徒快到 耶路撒冷 ，來到 伯法其 和 伯大尼 ，在 橄欖山 那裏。耶穌打發兩個門徒，
MARK|11|2|對他們說：「你們往對面村子裏去，一進去的時候會看見一匹驢駒拴在那裏，是從來沒有人騎過的，把牠解開，牽來。
MARK|11|3|若有人對你們說：『為甚麼做這事？』你們就說：『主要用牠，但會立刻把牠牽回到這裏來。』」
MARK|11|4|他們去了，看見一匹驢駒拴在門外街道上，就把牠解開。
MARK|11|5|在那裏站著的人，有幾個說：「你們解開驢駒做甚麼？」
MARK|11|6|門徒照著耶穌的話說，那些人就任憑他們牽去了。
MARK|11|7|他們把驢駒牽到耶穌那裏，把自己的衣服搭在上面，耶穌就騎上。
MARK|11|8|有許多人把衣服鋪在路上，還有人把田間的樹枝砍下來鋪上。
MARK|11|9|前呼後擁的人都喊著說： 「和散那 ！ 奉主名來的是應當稱頌的！
MARK|11|10|那將要來的我祖 大衛 之國是應當稱頌的！ 至高無上的，和散那！」
MARK|11|11|耶穌到了 耶路撒冷 ，進入聖殿，看了周圍的一切。天色已晚，他就和十二使徒出城，往 伯大尼 去。
MARK|11|12|第二天，他們從 伯大尼 出來，耶穌餓了。
MARK|11|13|他遠遠地看見一棵無花果樹，樹上有葉子，就過去，看是不是在樹上可以找到甚麼。他到了樹下，竟找不到甚麼，只有葉子，因為不是無花果的季節。
MARK|11|14|耶穌就對樹說：「從今以後，永沒有人吃你的果子。」他的門徒都聽到了。
MARK|11|15|他們來到 耶路撒冷 。耶穌一進聖殿，就趕出在聖殿裏做買賣的人，推倒兌換銀錢之人的桌子和賣鴿子之人的凳子；
MARK|11|16|也不許人拿著器具從聖殿裏經過。
MARK|11|17|他教導他們說：「經上不是記著： 『我的殿要稱為萬國禱告的殿嗎？ 你們倒使它成為賊窩了。』」
MARK|11|18|祭司長和文士聽見這話，就想法子要除掉耶穌，卻又怕他，因為眾人都對他的教導感到驚奇。
MARK|11|19|每天晚上，他們 都到城外去。
MARK|11|20|早晨，他們從那裏經過，看見無花果樹連根都枯乾了。
MARK|11|21|彼得 想起耶穌的話來，就對他說：「拉比，你看！你所詛咒的無花果樹已經枯乾了。」
MARK|11|22|耶穌回答：「你們對上帝要有信心。
MARK|11|23|我實在告訴你們，無論何人對這座山說：『離開此地，投在海裏！』他心裏若不疑惑，只信所說的必成，就為他實現。
MARK|11|24|所以我告訴你們，凡你們禱告祈求的，無論是甚麼，只要信你們已經得著了，就為你們實現。
MARK|11|25|你們站著禱告的時候，若想起有人得罪你們，就該饒恕他，好讓你們在天上的父也饒恕你們的過犯。 」
MARK|11|26|
MARK|11|27|他們又來到 耶路撒冷 。耶穌在聖殿裏行走的時候，祭司長、文士和長老進前來，
MARK|11|28|問他說：「你仗著甚麼權柄做這些事？給你權柄做這些事的是誰呢？」
MARK|11|29|耶穌對他們說：「我要問你們一句話，你們回答我，我就告訴你們我仗著甚麼權柄做這些事。
MARK|11|30|約翰 的洗禮是從天上來的，還是從人間來的呢？你們回答我吧。」
MARK|11|31|他們彼此商議說：「我們若說『從天上來的』，他會說：『這樣，你們為甚麼不信他呢？』
MARK|11|32|但若說『從人間來的』，卻又怕眾人，因為大家認為 約翰 確是先知。」
MARK|11|33|於是他們回答耶穌：「我們不知道。」耶穌說：「我也不告訴你們，我仗著甚麼權柄做這些事。」
MARK|12|1|耶穌就用比喻對他們說：「有人開墾了一個葡萄園，四周圍上籬笆，挖了一個榨酒池，蓋了一座守望樓，租給園戶，就出外遠行去了。
MARK|12|2|到了時候，他打發一個僕人到園戶那裏，要向他們收葡萄園的果子。
MARK|12|3|他們拿住他，打了他，叫他空手回去。
MARK|12|4|園主再打發一個僕人到他們那裏。他們打傷他的頭，並且侮辱他。
MARK|12|5|園主又打發一個僕人去，他們就殺了他。以後又打發好些僕人去，有的被他們打了，有的被他們殺了。
MARK|12|6|園主還有一位，是他的愛子，最後又打發他去，說：『他們會尊敬我的兒子。』
MARK|12|7|那些園戶卻彼此說：『這是承受產業的。來，我們殺了他，產業就歸我們了！』
MARK|12|8|於是他們拿住他，殺了他，把他扔出葡萄園。
MARK|12|9|這樣，葡萄園主要怎麼做呢？他要來除滅那些園戶，將葡萄園轉給別人。
MARK|12|10|『匠人所丟棄的石頭 已作了房角的頭塊石頭。 這是主所做的， 在我們眼中看為奇妙。』 這經文你們沒有念過嗎？」
MARK|12|11|
MARK|12|12|他們看出這比喻是指著他們說的，就想要捉拿他，但是懼怕眾人，於是離開他走了。
MARK|12|13|後來，他們打發幾個法利賽人和 希律 黨人到耶穌那裏，要用他自己的話陷害他。
MARK|12|14|他們來了，就對他說：「老師，我們知道你是誠實的，無論誰你都一視同仁；因為你不看人的面子，而是誠誠實實傳上帝的道。納稅給凱撒合不合法？
MARK|12|15|我們該不該納？」耶穌知道他們的虛偽，就對他們說：「你們為甚麼試探我？拿一個銀幣來給我看。」
MARK|12|16|他們就拿了來。耶穌問他們：「這像和這名號是誰的？」他們對他說：「是凱撒的。」
MARK|12|17|耶穌對他們說：「凱撒的歸凱撒；上帝的歸上帝。」他們對他非常驚訝。
MARK|12|18|撒都該人來見耶穌。他們說沒有復活這回事，於是問耶穌：
MARK|12|19|「老師， 摩西 為我們寫下這話：『某人的哥哥若死了，撇下妻子，沒有孩子，他該娶哥哥的妻子，為哥哥生子立後。』
MARK|12|20|那麼，有兄弟七人，第一個娶了妻，死了，沒有留下孩子。
MARK|12|21|第二個娶了她，也死了，沒有留下孩子。第三個也是這樣。
MARK|12|22|那七個人都沒有留下孩子。最後，那婦人也死了。
MARK|12|23|在復活的時候， 她是哪一個的妻子呢？因為他們七個人都娶過她。」
MARK|12|24|耶穌說：「你們錯了，不正是因為不明白聖經，也不知道上帝的大能嗎？
MARK|12|25|當人從死人中復活後，也不娶也不嫁，而是像天上的天使一樣。
MARK|12|26|論到死人復活，你們沒有念過 摩西 書中《荊棘篇》上所記載的嗎？上帝對 摩西 說：『我是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。』
MARK|12|27|上帝不是死人的上帝，而是活人的上帝。你們是大錯了。」
MARK|12|28|有一個文士來，聽見他們的辯論，知道耶穌回答得好，就問他說：「誡命中哪一條是第一呢？」
MARK|12|29|耶穌回答：「第一是：『 以色列 啊，你要聽，主—我們的上帝是獨一的主。
MARK|12|30|你要盡心、盡性、盡意、盡力愛主—你的上帝。』
MARK|12|31|第二是：『要愛鄰 如己。』再沒有比這兩條誡命更大的了。」
MARK|12|32|那文士對耶穌說：「好，老師，你說得對，上帝是一位，除了他以外，再沒有別的了；
MARK|12|33|並且盡心、盡智、盡力愛他，又愛鄰如己，要比一切燔祭和祭祀好得多。」
MARK|12|34|耶穌見他回答得有智慧，就對他說：「你離上帝的國不遠了。」從此以後，沒有人敢再問他甚麼。
MARK|12|35|耶穌在聖殿裏教導人，問他們說：「文士怎麼說基督是 大衛 的後裔呢？
MARK|12|36|大衛 被聖靈感動，說： 『主對我主說： 你坐在我的右邊， 等我把你的仇敵放在你腳下 。』
MARK|12|37|大衛 親自稱他為主，他怎麼又是 大衛 的後裔呢？」一大群的人都喜歡聽他。
MARK|12|38|他在教導的時候，說：「你們要防備文士。他們好穿長袍走來走去，喜歡人們在街市上向他們問安，
MARK|12|39|又喜愛會堂裏的高位，宴席上的首座。
MARK|12|40|他們侵吞寡婦的家產，假意作很長的禱告。這些人要受更重的懲罰！」
MARK|12|41|耶穌面向聖殿銀庫坐著，看眾人怎樣把錢投入銀庫。有好些財主投了許多錢。
MARK|12|42|有一個窮寡婦來，投了兩個小文錢 ，就是一個大文錢 。
MARK|12|43|耶穌叫門徒來，對他們說：「我實在告訴你們，這窮寡婦投入銀庫裏的比眾人所投的更多。
MARK|12|44|因為，眾人都是拿有餘的捐獻，但這寡婦，雖然自己不足，卻把她一生所有的全都投進去了。」
MARK|13|1|耶穌從聖殿裏出來的時候，有一個門徒對他說：「老師，請看，這是多麼了不起的石頭！多麼了不起的建築！」
MARK|13|2|耶穌對他說：「你看見這些宏偉的建築嗎？這裏將沒有一塊石頭會留在另一塊石頭上而不被拆毀的。」
MARK|13|3|耶穌在 橄欖山 上，面向聖殿坐著； 彼得 、 雅各 、 約翰 和 安得烈 私下問他說：
MARK|13|4|「請告訴我們，甚麼時候有這些事呢？這一切事將成的時候有甚麼預兆呢？」
MARK|13|5|耶穌說：「你們要謹慎，免得有人迷惑你們。
MARK|13|6|將有好些人冒我的名來，說『我是基督』，並且要迷惑許多人。
MARK|13|7|當你們聽見打仗和打仗的風聲，不要驚慌；這些事必須發生，但這還不是終結。
MARK|13|8|民要攻打民，國要攻打國，多處必有地震、饑荒。這都是災難 的起頭。
MARK|13|9|但你們自己要謹慎；因為有人要把你們交給議會，並且你們在會堂裏要受鞭打，又為我的緣故站在統治者和君王面前，對他們作見證。
MARK|13|10|然而，福音必須先傳給萬民。
MARK|13|11|有人把你們解送去受審的時候，不要事先擔心說甚麼；到那時候，賜給你們甚麼話，你們就說甚麼；因為說話的不是你們，而是聖靈。
MARK|13|12|兄弟要把兄弟、父親要把兒女置於死地；兒女要起來與父母為敵，害死他們；
MARK|13|13|而且你們要為我的名被眾人憎恨。但堅忍到底的終必得救。」
MARK|13|14|「當你們看見那『施行毀滅的褻瀆者』站在不當站的地方（讀這經的人要會意），那時，在 猶太 的，應當逃到山上；
MARK|13|15|在屋頂上的，不要下來，也不要進家裏去拿東西；
MARK|13|16|在田裏的，不要回去取衣裳。
MARK|13|17|在那些日子，懷孕的和奶孩子的就苦了。
MARK|13|18|你們要祈求，叫這事不在冬天發生。
MARK|13|19|因為，在那些日子必有災難，自從上帝創造萬物直到如今，從沒有這樣的災難，將來也不會有。
MARK|13|20|若不是主減少那些日子，凡血肉之軀的，就沒有一個能得救；但是為了他所揀選的選民，他將那些日子減少了。
MARK|13|21|那時，若有人對你們說：『看哪，基督在這裏！看哪，在那裏！』你們不要信。
MARK|13|22|因為假基督和假先知將要起來，顯神蹟奇事，如果可能，連選民也迷惑了。
MARK|13|23|你們要謹慎！凡事我都預先告訴你們了。」
MARK|13|24|「在那些日子、那災難以後， 太陽要變黑，月亮也不放光，
MARK|13|25|眾星要從天上墜落， 天上的萬象都要震動。
MARK|13|26|那時，他們要看見人子帶著大能力和榮耀駕雲來臨。
MARK|13|27|他要差遣天使，從四方，從地極直到天邊，召集他的選民。」
MARK|13|28|「你們要從無花果樹學習功課：當樹枝發芽長葉的時候，你們就知道夏天近了。
MARK|13|29|同樣，當你們看見這些事發生，就知道那時候近了，就在門口了。
MARK|13|30|我實在告訴你們，這世代還沒有過去，這一切都要發生。
MARK|13|31|天地要廢去，我的話卻絕不廢去。」
MARK|13|32|「但那日子，那時辰，沒有人知道，連天上的天使也不知道，子也不知道，惟有父知道。
MARK|13|33|你們要謹慎，要警醒 ，因為你們不知道那時刻幾時來到。
MARK|13|34|這事正如一個人離家遠行，授權給僕人們，分派各人的工作，又吩咐看門的警醒。
MARK|13|35|所以，你們要警醒，因為你們不知道這家的主人甚麼時候來，是晚上，或半夜，或雞叫時，或早晨，
MARK|13|36|免得他忽然來到，看見你們睡著了。
MARK|13|37|我對你們所說的話，也是對眾人說的：要警醒！」
MARK|14|1|過兩天是逾越節，又是除酵節，祭司長和文士在想法子怎樣設計捉拿耶穌，把他殺掉。
MARK|14|2|他們說：「不可在過節的日子，恐怕百姓生亂。」
MARK|14|3|耶穌在 伯大尼 痲瘋病人 西門 家裏坐席的時候，有一個女人拿著一玉瓶極貴的純哪噠 香膏來，打破玉瓶，把膏澆在耶穌的頭上。
MARK|14|4|有幾個人心中很不高興，說：「何必這樣浪費香膏呢？
MARK|14|5|這香膏可以賣三百多個銀幣賙濟窮人。」他們就對那女人生氣。
MARK|14|6|耶穌說：「由她吧！為甚麼難為她呢？她在我身上做的是一件美事。
MARK|14|7|因為常有窮人和你們在一起，要向他們行善，隨時都可以，但是你們不常有我。
MARK|14|8|她所做的是盡她所能的；她是為了我的安葬，把香膏預先澆在我身上。
MARK|14|9|我實在告訴你們，普天之下，無論在甚麼地方傳這福音，都要述說這女人所做的，來記念她。」
MARK|14|10|十二使徒中有一個 加略 人 猶大 ，去見祭司長，要把耶穌交給他們。
MARK|14|11|他們聽見就很高興，又應許給他銀子；他就想怎樣找機會把耶穌交給他們。
MARK|14|12|除酵節的第一天，就是宰逾越節羔羊的那一天，門徒對耶穌說：「你要我們到哪裏去預備你吃逾越節的宴席呢？」
MARK|14|13|耶穌就打發兩個門徒，對他們說：「你們進城去，會有人拿著一罐水迎面而來，你們就跟著他。
MARK|14|14|無論他進哪一家，你們就對那家的主人說：『老師問：我的客房在哪裏？我和我的門徒要在那裏吃逾越節的宴席。』
MARK|14|15|他會帶你們看一間擺設齊全、準備妥當的樓上大廳，你們就在那裏為我們預備。」
MARK|14|16|門徒出去，進了城，所看到的正如耶穌所說的。他們就預備了逾越節的宴席。
MARK|14|17|到了晚上，耶穌和十二使徒都來了。
MARK|14|18|他們坐席，正吃的時候，耶穌說：「我實在告訴你們，你們中間有一個與我同吃的人要出賣我了。」
MARK|14|19|他們就憂愁起來，一個個地問他：「不是我吧？」
MARK|14|20|耶穌對他們說：「是十二人中的一個，就是同我蘸餅在盤子裏的那個人。
MARK|14|21|人子要去了，正如經上所寫有關他的；但出賣人子的人有禍了！那人沒有出生倒好。」
MARK|14|22|他們吃的時候，耶穌拿起餅來，祝福了，就擘開，遞給他們，說：「你們拿去，這是我的身體。」
MARK|14|23|他又拿起杯來，祝謝了，遞給他們；他們都喝了。
MARK|14|24|耶穌對他們說：「這是我立約的血，為許多人流出來的。
MARK|14|25|我實在告訴你們，我不再喝這葡萄汁，直到我在上帝的國裏喝新的那日子。」
MARK|14|26|他們唱了詩，就出來往 橄欖山 去。
MARK|14|27|耶穌對他們說：「你們都要跌倒，因為經上記著： 『我要擊打牧人， 羊就分散了。』，　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　
MARK|14|28|但我復活以後，要在你們之前往 加利利 去。」
MARK|14|29|彼得 說：「雖然眾人跌倒，但我不會。」
MARK|14|30|耶穌對他說：「我實在告訴你，今天夜裏，雞叫兩遍 以前，你要三次不認我。」
MARK|14|31|彼得 卻極力地說：「我就是必須和你同死，也絕不會不認你。」所有的門徒 都是這樣說。
MARK|14|32|他們來到一個地方，名叫 客西馬尼 。耶穌對門徒說：「你們坐在這裏，我去禱告。」
MARK|14|33|於是他帶著 彼得 、 雅各 和 約翰 同去。他驚恐起來，極其難過，
MARK|14|34|對他們說：「我心裏非常憂傷，幾乎要死；你們留在這裏，要警醒。」
MARK|14|35|他就稍往前走，俯伏在地，禱告說，如果可能，就叫那時候離開他。
MARK|14|36|他說：「阿爸，父啊！在你凡事都能；求你將這杯撤去。然而，不是照我所願的，而是照你所願的。」
MARK|14|37|耶穌回來，見他們睡著了，就對 彼得 說：「 西門 ，你睡著了嗎？不能警醒一小時嗎？
MARK|14|38|總要警醒禱告，免得陷入試探。你們心靈固然願意，肉體卻軟弱了。」
MARK|14|39|耶穌又去禱告，說的話跟先前一樣。
MARK|14|40|他又來，見他們睡著了，因為他們的眼睛很困倦；他們也不知道怎麼回答他。
MARK|14|41|他第三次來對他們說：「現在你們仍在睡覺安歇嗎？夠了，時候到了。看哪，人子被出賣在罪人手裏了。
MARK|14|42|起來，我們走吧！看哪，那出賣我的人快來了。」
MARK|14|43|耶穌還在說話的時候，忽然十二使徒之一的 猶大 來了，還有一群人帶著刀棒，從祭司長、文士和長老那裏跟他同來。
MARK|14|44|那出賣耶穌的人曾給他們一個暗號，說：「我親誰，誰就是。你們把他抓住，穩妥地帶走。」
MARK|14|45|猶大 來了，隨即到耶穌跟前，說：「拉比」，就跟他親吻。
MARK|14|46|他們就下手抓住他。
MARK|14|47|旁邊站著的人，有一個拔出刀來，把大祭司的僕人砍了一刀，削掉了他一隻耳朵。
MARK|14|48|耶穌回應他們說：「你們帶著刀棒出來拿我，如同拿強盜嗎？
MARK|14|49|我天天教導人，同你們在殿裏，你們並沒有抓我。但這是要應驗經上的話。」
MARK|14|50|門徒都離開他，逃走了。
MARK|14|51|有一個青年光著身子，只披一塊麻布，跟隨耶穌，眾人就抓住他。
MARK|14|52|他卻丟下麻布，赤身逃走了。
MARK|14|53|他們把耶穌帶到大祭司那裏，又有眾祭司長、長老和文士都來一同聚集。
MARK|14|54|彼得 遠遠地跟著耶穌，直到進了大祭司的院子，和警衛一同坐在火邊取暖。
MARK|14|55|祭司長和全議會尋找見證控告耶穌，要處死他，卻找不到實據。
MARK|14|56|因為有好些人作假見證告他，他們的見證又各不相符。
MARK|14|57|又有幾個人站起來，作假見證告他說：
MARK|14|58|「我們聽見他說：『我要拆毀這人手所造的殿，三日內另造一座不是人手所造的。』」
MARK|14|59|就是這樣，他們的見證還是不相符。
MARK|14|60|大祭司起來站在中間，問耶穌說：「這些人作證告你的事，你甚麼都不回答嗎？」
MARK|14|61|耶穌卻不言語，一句也不回答。大祭司又問他：「你是不是基督，那當稱頌者的兒子？」
MARK|14|62|耶穌說：「我是。 你們要看見人子 坐在那權能者的右邊， 駕著天上的雲來臨。」
MARK|14|63|大祭司就撕裂衣服，說：「我們何必再要證人呢？
MARK|14|64|你們已經聽見他這褻瀆的話了。你們的決定如何？」他們都判定他該處死。
MARK|14|65|於是有人開始向他吐唾沫，又蒙著他的臉，用拳頭打他，對他說：「你說預言吧！」警衛把他拉過來，打他耳光。
MARK|14|66|彼得 在下邊院子裏，大祭司的一個使女來了，
MARK|14|67|見 彼得 取暖，就看著他，說：「你素來也是同 拿撒勒 人耶穌一起的。」
MARK|14|68|彼得 卻不承認，說：「我不知道，也不明白你說的是甚麼！」於是他出來，到了前院，雞就叫了 。
MARK|14|69|那使女看見他，又對旁邊站著的人說：「這個人也是他們一夥的。」
MARK|14|70|彼得 又不承認。過了不久，旁邊站著的人又對 彼得 說：「你真是他們一夥的，因為你也是 加利利 人。」
MARK|14|71|彼得 就賭咒發誓說：「我不認得你們說的這個人。」
MARK|14|72|立刻，雞叫了第二遍。 彼得 想起耶穌對他所說的話：「雞叫兩遍以前，你要三次不認我。」他就忍不住哭了。
MARK|15|1|一到早晨，眾祭司長、長老、文士，和全議會的人大家商議，就把耶穌綁著，解去，交給 彼拉多 。
MARK|15|2|彼拉多 問他：「你是 猶太 人的王嗎？」耶穌回答：「是你說的。」
MARK|15|3|祭司長們告他許多的事。
MARK|15|4|彼拉多 又問他：「你看，他們告你這麼多的事，你甚麼都不回答嗎？」
MARK|15|5|耶穌仍不回答，以致 彼拉多 覺得驚訝。
MARK|15|6|每逢這節期， 彼拉多 照眾人所求的，釋放一個囚犯給他們。
MARK|15|7|有一個人名叫 巴拉巴 ，和作亂的人監禁在一起。他們作亂的時候曾殺過人。
MARK|15|8|眾人上去求 彼拉多 照常例給他們辦理。
MARK|15|9|彼拉多 說：「你們要我釋放 猶太 人的王給你們嗎？」
MARK|15|10|他原知道祭司長們是因嫉妒才把耶穌解了來。
MARK|15|11|但是祭司長們煽動眾人，寧可要他釋放 巴拉巴 給他們。
MARK|15|12|彼拉多 又說：「那麼，你們稱為 猶太 人的王的 ，要 我怎麼辦他呢？」
MARK|15|13|他們又再喊著：「把他釘十字架！」
MARK|15|14|彼拉多 說：「為甚麼？他做了甚麼惡事呢？」他們更加喊著：「把他釘十字架！」
MARK|15|15|彼拉多 要討好眾人，就釋放 巴拉巴 給他們，把耶穌鞭打後交給人釘十字架。
MARK|15|16|士兵把耶穌帶進總督府的庭院裏，叫齊了全營的兵。
MARK|15|17|他們給他穿上紫袍，又用荊棘編了冠冕給他戴上，
MARK|15|18|然後向他致敬，說：「萬歲， 猶太 人的王！」
MARK|15|19|他們又拿一根蘆葦稈打他的頭，向他吐唾沫，屈膝拜他。
MARK|15|20|他們戲弄完了，就給他脫了紫袍，又穿上他自己的衣服，帶他出去，要把他釘十字架。
MARK|15|21|有一個 古利奈 人 西門 ，就是 亞歷山大 和 魯孚 的父親，從鄉下來，經過那地方，他們就強迫他同去，好背耶穌的十字架。
MARK|15|22|他們帶耶穌到了一個地方叫 各各他 （翻出來就是「髑髏地」），
MARK|15|23|拿沒藥調和的酒給耶穌，他卻不受。
MARK|15|24|於是他們把他釘在十字架上，抽籤分他的衣服，看誰得甚麼。
MARK|15|25|他們把他釘十字架的時候是上午九點鐘。
MARK|15|26|罪狀牌上寫的是：「 猶太 人的王。」
MARK|15|27|他們又把兩個強盜和他同釘十字架，一個在右邊，一個在左邊。
MARK|15|28|
MARK|15|29|從那裏經過的人譏笑他，搖著頭，說：「哼！你這拆毀殿、三日又建造起來的，
MARK|15|30|救救你自己，從十字架上下來呀！」
MARK|15|31|眾祭司長和文士也這樣嘲笑他，彼此說：「他救了別人，不能救自己。
MARK|15|32|以色列 的王基督，現在從十字架上下來，好讓我們看見就信了呀！」那和他同釘的人也譏諷他。
MARK|15|33|到了正午，全地都黑暗了，直到下午三點鐘。
MARK|15|34|下午三點鐘的時候，耶穌大聲呼喊：「以羅伊！以羅伊！拉馬撒巴各大尼？」（翻出來就是：我的上帝！我的上帝！為甚麼離棄我？）
MARK|15|35|旁邊站著的人，有的聽見就說：「看哪，他叫 以利亞 呢！」
MARK|15|36|有一個人跑去，把海綿蘸滿了醋，綁在蘆葦稈上，送給他喝，說：「且等著，看 以利亞 會不會來把他放下來。」
MARK|15|37|耶穌大喊一聲，氣就斷了。
MARK|15|38|殿的幔子從上到下裂為兩半。
MARK|15|39|對面站著的百夫長看見耶穌這樣斷氣 ，就說：「這人真是上帝的兒子！」
MARK|15|40|還有些婦女遠遠地觀看，其中有 抹大拉 的 馬利亞 ，又有小 雅各 和 約西 的母親 馬利亞 ，並有 撒羅米 ，
MARK|15|41|就是耶穌在 加利利 的時候，跟隨他、服事他的那些人，還有同耶穌上 耶路撒冷 的好些婦女。
MARK|15|42|到了晚上，因為這是預備日，就是安息日的前一日，
MARK|15|43|有 亞利馬太 的 約瑟 前來，他是尊貴的議員，也是盼望著上帝國的，他放膽進去見 彼拉多 ，請求要耶穌的身體。
MARK|15|44|彼拉多 詫異耶穌已經死了，就叫百夫長來，問他耶穌是不是死了很久；
MARK|15|45|既從百夫長得知實情，就把耶穌的身體賜給 約瑟 。
MARK|15|46|約瑟 買了細麻布，把耶穌取下來，用細麻布裹好，安放在巖石中鑿出來的墓穴裏，又滾來一塊石頭擋住墓門。
MARK|15|47|抹大拉 的 馬利亞 和 約西 的母親 馬利亞 都看見安放他的地方。
MARK|16|1|過了安息日， 抹大拉 的 馬利亞 、 雅各 的母親 馬利亞 ，和 撒羅米 ，買了香料，要去膏耶穌的身體。
MARK|16|2|七日的第一日清早，太陽出來後，她們來到墳墓那裏，
MARK|16|3|彼此說：「誰要替我們把石頭從墓門滾開呢？」
MARK|16|4|她們抬頭一看，看見石頭已經滾開了，原來那石頭很大。
MARK|16|5|她們進了墳墓，看見一個年輕人坐在右邊，穿著白袍，就很驚奇。
MARK|16|6|那年輕人對她們說：「不要驚慌！你們尋找那釘十字架的 拿撒勒 人耶穌，他已經復活了，不在這裏。來看安放他的地方。
MARK|16|7|你們去，對他的門徒和 彼得 說：『他要比你們先到 加利利 去，在那裏你們會看見他，正如他從前所告訴你們的。』」
MARK|16|8|於是她們出來，從墳墓那裏逃走，又發抖又驚訝，甚麼也沒有告訴人，因為她們害怕。 〔
MARK|16|9|凡耶穌所吩咐的，她們簡潔地告訴 彼得 和他周圍的人。這些事以後，耶穌親自藉著他的門徒，從東到西，把那神聖、不朽、永遠拯救的福音傳出去。阿們！〕 〔 在七日的第一日清早，耶穌復活了，先向 抹大拉 的 馬利亞 顯現；耶穌曾從她身上趕出七個鬼。
MARK|16|10|她去告訴那向來跟隨耶穌的人；那時他們正哀慟哭泣。
MARK|16|11|他們聽見耶穌活了，被 馬利亞 看見，可是不信。〕 〔
MARK|16|12|這些事以後，門徒中有兩個人往鄉下去；正走著的時候，耶穌以另一種形像向他們顯現。
MARK|16|13|他們去告訴其餘的門徒，那些門徒還是不信。〕 〔
MARK|16|14|後來十一使徒坐席的時候，耶穌向他們顯現，責備他們不信，心裏剛硬，因為他們不信那些在他復活以後看見他的人。
MARK|16|15|他又對他們說：「你們往普天下去，傳福音給萬民 聽。
MARK|16|16|信而受洗的必然得救，不信的必被定罪。
MARK|16|17|信的人將有神蹟隨著他們：就是奉我的名趕鬼；說新方言；
MARK|16|18|手 能拿蛇；若喝了甚麼毒物，也不會受害；手按病人，病人就好了。」〕 〔
MARK|16|19|主耶穌 和他們說完了話以後，被接到天上，坐在上帝的右邊。
MARK|16|20|門徒出去，到處傳福音。主和他們同工，藉著伴隨的神蹟證實所傳的道。 〕
