2SAM|1|1|After the death of Saul, David returned from defeating the Amalekites and stayed in Ziklag two days.
2SAM|1|2|On the third day a man arrived from Saul's camp, with his clothes torn and with dust on his head. When he came to David, he fell to the ground to pay him honor.
2SAM|1|3|"Where have you come from?" David asked him. He answered, "I have escaped from the Israelite camp."
2SAM|1|4|"What happened?" David asked. "Tell me." He said, "The men fled from the battle. Many of them fell and died. And Saul and his son Jonathan are dead."
2SAM|1|5|Then David said to the young man who brought him the report, "How do you know that Saul and his son Jonathan are dead?"
2SAM|1|6|"I happened to be on Mount Gilboa," the young man said, "and there was Saul, leaning on his spear, with the chariots and riders almost upon him.
2SAM|1|7|When he turned around and saw me, he called out to me, and I said, 'What can I do?'
2SAM|1|8|"He asked me, 'Who are you?'"'An Amalekite,' I answered.
2SAM|1|9|"Then he said to me, 'Stand over me and kill me! I am in the throes of death, but I'm still alive.'
2SAM|1|10|"So I stood over him and killed him, because I knew that after he had fallen he could not survive. And I took the crown that was on his head and the band on his arm and have brought them here to my lord."
2SAM|1|11|Then David and all the men with him took hold of their clothes and tore them.
2SAM|1|12|They mourned and wept and fasted till evening for Saul and his son Jonathan, and for the army of the LORD and the house of Israel, because they had fallen by the sword.
2SAM|1|13|David said to the young man who brought him the report, "Where are you from?I am the son of an alien, an Amalekite," he answered.
2SAM|1|14|David asked him, "Why were you not afraid to lift your hand to destroy the LORD's anointed?"
2SAM|1|15|Then David called one of his men and said, "Go, strike him down!" So he struck him down, and he died.
2SAM|1|16|For David had said to him, "Your blood be on your own head. Your own mouth testified against you when you said, 'I killed the LORD's anointed.'"
2SAM|1|17|David took up this lament concerning Saul and his son Jonathan,
2SAM|1|18|and ordered that the men of Judah be taught this lament of the bow (it is written in the Book of Jashar):
2SAM|1|19|"Your glory, O Israel, lies slain on your heights. How the mighty have fallen!
2SAM|1|20|"Tell it not in Gath, proclaim it not in the streets of Ashkelon, lest the daughters of the Philistines be glad, lest the daughters of the uncircumcised rejoice.
2SAM|1|21|"O mountains of Gilboa, may you have neither dew nor rain, nor fields that yield offerings of grain. For there the shield of the mighty was defiled, the shield of Saul-no longer rubbed with oil.
2SAM|1|22|From the blood of the slain, from the flesh of the mighty, the bow of Jonathan did not turn back, the sword of Saul did not return unsatisfied.
2SAM|1|23|"Saul and Jonathan- in life they were loved and gracious, and in death they were not parted. They were swifter than eagles, they were stronger than lions.
2SAM|1|24|"O daughters of Israel, weep for Saul, who clothed you in scarlet and finery, who adorned your garments with ornaments of gold.
2SAM|1|25|"How the mighty have fallen in battle! Jonathan lies slain on your heights.
2SAM|1|26|I grieve for you, Jonathan my brother; you were very dear to me. Your love for me was wonderful, more wonderful than that of women.
2SAM|1|27|"How the mighty have fallen! The weapons of war have perished!"
2SAM|2|1|In the course of time, David inquired of the LORD. "Shall I go up to one of the towns of Judah?" he asked. The LORD said, "Go up." David asked, "Where shall I go?To Hebron," the LORD answered.
2SAM|2|2|So David went up there with his two wives, Ahinoam of Jezreel and Abigail, the widow of Nabal of Carmel.
2SAM|2|3|David also took the men who were with him, each with his family, and they settled in Hebron and its towns.
2SAM|2|4|Then the men of Judah came to Hebron and there they anointed David king over the house of Judah. When David was told that it was the men of Jabesh Gilead who had buried Saul,
2SAM|2|5|he sent messengers to the men of Jabesh Gilead to say to them, "The LORD bless you for showing this kindness to Saul your master by burying him.
2SAM|2|6|May the LORD now show you kindness and faithfulness, and I too will show you the same favor because you have done this.
2SAM|2|7|Now then, be strong and brave, for Saul your master is dead, and the house of Judah has anointed me king over them."
2SAM|2|8|Meanwhile, Abner son of Ner, the commander of Saul's army, had taken Ish-Bosheth son of Saul and brought him over to Mahanaim.
2SAM|2|9|He made him king over Gilead, Ashuri and Jezreel, and also over Ephraim, Benjamin and all Israel.
2SAM|2|10|Ish-Bosheth son of Saul was forty years old when he became king over Israel, and he reigned two years. The house of Judah, however, followed David.
2SAM|2|11|The length of time David was king in Hebron over the house of Judah was seven years and six months.
2SAM|2|12|Abner son of Ner, together with the men of Ish-Bosheth son of Saul, left Mahanaim and went to Gibeon.
2SAM|2|13|Joab son of Zeruiah and David's men went out and met them at the pool of Gibeon. One group sat down on one side of the pool and one group on the other side.
2SAM|2|14|Then Abner said to Joab, "Let's have some of the young men get up and fight hand to hand in front of us.All right, let them do it," Joab said.
2SAM|2|15|So they stood up and were counted off-twelve men for Benjamin and Ish-Bosheth son of Saul, and twelve for David.
2SAM|2|16|Then each man grabbed his opponent by the head and thrust his dagger into his opponent's side, and they fell down together. So that place in Gibeon was called Helkath Hazzurim.
2SAM|2|17|The battle that day was very fierce, and Abner and the men of Israel were defeated by David's men.
2SAM|2|18|The three sons of Zeruiah were there: Joab, Abishai and Asahel. Now Asahel was as fleet-footed as a wild gazelle.
2SAM|2|19|He chased Abner, turning neither to the right nor to the left as he pursued him.
2SAM|2|20|Abner looked behind him and asked, "Is that you, Asahel?It is," he answered.
2SAM|2|21|Then Abner said to him, "Turn aside to the right or to the left; take on one of the young men and strip him of his weapons." But Asahel would not stop chasing him.
2SAM|2|22|Again Abner warned Asahel, "Stop chasing me! Why should I strike you down? How could I look your brother Joab in the face?"
2SAM|2|23|But Asahel refused to give up the pursuit; so Abner thrust the butt of his spear into Asahel's stomach, and the spear came out through his back. He fell there and died on the spot. And every man stopped when he came to the place where Asahel had fallen and died.
2SAM|2|24|But Joab and Abishai pursued Abner, and as the sun was setting, they came to the hill of Ammah, near Giah on the way to the wasteland of Gibeon.
2SAM|2|25|Then the men of Benjamin rallied behind Abner. They formed themselves into a group and took their stand on top of a hill.
2SAM|2|26|Abner called out to Joab, "Must the sword devour forever? Don't you realize that this will end in bitterness? How long before you order your men to stop pursuing their brothers?"
2SAM|2|27|Joab answered, "As surely as God lives, if you had not spoken, the men would have continued the pursuit of their brothers until morning. "
2SAM|2|28|So Joab blew the trumpet, and all the men came to a halt; they no longer pursued Israel, nor did they fight anymore.
2SAM|2|29|All that night Abner and his men marched through the Arabah. They crossed the Jordan, continued through the whole Bithron and came to Mahanaim.
2SAM|2|30|Then Joab returned from pursuing Abner and assembled all his men. Besides Asahel, nineteen of David's men were found missing.
2SAM|2|31|But David's men had killed three hundred and sixty Benjamites who were with Abner.
2SAM|2|32|They took Asahel and buried him in his father's tomb at Bethlehem. Then Joab and his men marched all night and arrived at Hebron by daybreak.
2SAM|3|1|The war between the house of Saul and the house of David lasted a long time. David grew stronger and stronger, while the house of Saul grew weaker and weaker.
2SAM|3|2|Sons were born to David in Hebron: His firstborn was Amnon the son of Ahinoam of Jezreel;
2SAM|3|3|his second, Kileab the son of Abigail the widow of Nabal of Carmel; the third, Absalom the son of Maacah daughter of Talmai king of Geshur;
2SAM|3|4|the fourth, Adonijah the son of Haggith; the fifth, Shephatiah the son of Abital;
2SAM|3|5|and the sixth, Ithream the son of David's wife Eglah. These were born to David in Hebron.
2SAM|3|6|During the war between the house of Saul and the house of David, Abner had been strengthening his own position in the house of Saul.
2SAM|3|7|Now Saul had had a concubine named Rizpah daughter of Aiah. And Ish-Bosheth said to Abner, "Why did you sleep with my father's concubine?"
2SAM|3|8|Abner was very angry because of what Ish-Bosheth said and he answered, "Am I a dog's head-on Judah's side? This very day I am loyal to the house of your father Saul and to his family and friends. I haven't handed you over to David. Yet now you accuse me of an offense involving this woman!
2SAM|3|9|May God deal with Abner, be it ever so severely, if I do not do for David what the LORD promised him on oath
2SAM|3|10|and transfer the kingdom from the house of Saul and establish David's throne over Israel and Judah from Dan to Beersheba."
2SAM|3|11|Ish-Bosheth did not dare to say another word to Abner, because he was afraid of him.
2SAM|3|12|Then Abner sent messengers on his behalf to say to David, "Whose land is it? Make an agreement with me, and I will help you bring all Israel over to you."
2SAM|3|13|"Good," said David. "I will make an agreement with you. But I demand one thing of you: Do not come into my presence unless you bring Michal daughter of Saul when you come to see me."
2SAM|3|14|Then David sent messengers to Ish-Bosheth son of Saul, demanding, "Give me my wife Michal, whom I betrothed to myself for the price of a hundred Philistine foreskins."
2SAM|3|15|So Ish-Bosheth gave orders and had her taken away from her husband Paltiel son of Laish.
2SAM|3|16|Her husband, however, went with her, weeping behind her all the way to Bahurim. Then Abner said to him, "Go back home!" So he went back.
2SAM|3|17|Abner conferred with the elders of Israel and said, "For some time you have wanted to make David your king.
2SAM|3|18|Now do it! For the LORD promised David, 'By my servant David I will rescue my people Israel from the hand of the Philistines and from the hand of all their enemies.'"
2SAM|3|19|Abner also spoke to the Benjamites in person. Then he went to Hebron to tell David everything that Israel and the whole house of Benjamin wanted to do.
2SAM|3|20|When Abner, who had twenty men with him, came to David at Hebron, David prepared a feast for him and his men.
2SAM|3|21|Then Abner said to David, "Let me go at once and assemble all Israel for my lord the king, so that they may make a compact with you, and that you may rule over all that your heart desires." So David sent Abner away, and he went in peace.
2SAM|3|22|Just then David's men and Joab returned from a raid and brought with them a great deal of plunder. But Abner was no longer with David in Hebron, because David had sent him away, and he had gone in peace.
2SAM|3|23|When Joab and all the soldiers with him arrived, he was told that Abner son of Ner had come to the king and that the king had sent him away and that he had gone in peace.
2SAM|3|24|So Joab went to the king and said, "What have you done? Look, Abner came to you. Why did you let him go? Now he is gone!
2SAM|3|25|You know Abner son of Ner; he came to deceive you and observe your movements and find out everything you are doing."
2SAM|3|26|Joab then left David and sent messengers after Abner, and they brought him back from the well of Sirah. But David did not know it.
2SAM|3|27|Now when Abner returned to Hebron, Joab took him aside into the gateway, as though to speak with him privately. And there, to avenge the blood of his brother Asahel, Joab stabbed him in the stomach, and he died.
2SAM|3|28|Later, when David heard about this, he said, "I and my kingdom are forever innocent before the LORD concerning the blood of Abner son of Ner.
2SAM|3|29|May his blood fall upon the head of Joab and upon all his father's house! May Joab's house never be without someone who has a running sore or leprosy or who leans on a crutch or who falls by the sword or who lacks food."
2SAM|3|30|(Joab and his brother Abishai murdered Abner because he had killed their brother Asahel in the battle at Gibeon.)
2SAM|3|31|Then David said to Joab and all the people with him, "Tear your clothes and put on sackcloth and walk in mourning in front of Abner." King David himself walked behind the bier.
2SAM|3|32|They buried Abner in Hebron, and the king wept aloud at Abner's tomb. All the people wept also.
2SAM|3|33|The king sang this lament for Abner: "Should Abner have died as the lawless die?
2SAM|3|34|Your hands were not bound, your feet were not fettered. You fell as one falls before wicked men." And all the people wept over him again.
2SAM|3|35|Then they all came and urged David to eat something while it was still day; but David took an oath, saying, "May God deal with me, be it ever so severely, if I taste bread or anything else before the sun sets!"
2SAM|3|36|All the people took note and were pleased; indeed, everything the king did pleased them.
2SAM|3|37|So on that day all the people and all Israel knew that the king had no part in the murder of Abner son of Ner.
2SAM|3|38|Then the king said to his men, "Do you not realize that a prince and a great man has fallen in Israel this day?
2SAM|3|39|And today, though I am the anointed king, I am weak, and these sons of Zeruiah are too strong for me. May the LORD repay the evildoer according to his evil deeds!"
2SAM|4|1|When Ish-Bosheth son of Saul heard that Abner had died in Hebron, he lost courage, and all Israel became alarmed.
2SAM|4|2|Now Saul's son had two men who were leaders of raiding bands. One was named Baanah and the other Recab; they were sons of Rimmon the Beerothite from the tribe of Benjamin-Beeroth is considered part of Benjamin,
2SAM|4|3|because the people of Beeroth fled to Gittaim and have lived there as aliens to this day.
2SAM|4|4|(Jonathan son of Saul had a son who was lame in both feet. He was five years old when the news about Saul and Jonathan came from Jezreel. His nurse picked him up and fled, but as she hurried to leave, he fell and became crippled. His name was Mephibosheth.)
2SAM|4|5|Now Recab and Baanah, the sons of Rimmon the Beerothite, set out for the house of Ish-Bosheth, and they arrived there in the heat of the day while he was taking his noonday rest.
2SAM|4|6|They went into the inner part of the house as if to get some wheat, and they stabbed him in the stomach. Then Recab and his brother Baanah slipped away.
2SAM|4|7|They had gone into the house while he was lying on the bed in his bedroom. After they stabbed and killed him, they cut off his head. Taking it with them, they traveled all night by way of the Arabah.
2SAM|4|8|They brought the head of Ish-Bosheth to David at Hebron and said to the king, "Here is the head of Ish-Bosheth son of Saul, your enemy, who tried to take your life. This day the LORD has avenged my lord the king against Saul and his offspring."
2SAM|4|9|David answered Recab and his brother Baanah, the sons of Rimmon the Beerothite, "As surely as the LORD lives, who has delivered me out of all trouble,
2SAM|4|10|when a man told me, 'Saul is dead,' and thought he was bringing good news, I seized him and put him to death in Ziklag. That was the reward I gave him for his news!
2SAM|4|11|How much more-when wicked men have killed an innocent man in his own house and on his own bed-should I not now demand his blood from your hand and rid the earth of you!"
2SAM|4|12|So David gave an order to his men, and they killed them. They cut off their hands and feet and hung the bodies by the pool in Hebron. But they took the head of Ish-Bosheth and buried it in Abner's tomb at Hebron.
2SAM|5|1|All the tribes of Israel came to David at Hebron and said, "We are your own flesh and blood.
2SAM|5|2|In the past, while Saul was king over us, you were the one who led Israel on their military campaigns. And the LORD said to you, 'You will shepherd my people Israel, and you will become their ruler.'"
2SAM|5|3|When all the elders of Israel had come to King David at Hebron, the king made a compact with them at Hebron before the LORD, and they anointed David king over Israel.
2SAM|5|4|David was thirty years old when he became king, and he reigned forty years.
2SAM|5|5|In Hebron he reigned over Judah seven years and six months, and in Jerusalem he reigned over all Israel and Judah thirty-three years.
2SAM|5|6|The king and his men marched to Jerusalem to attack the Jebusites, who lived there. The Jebusites said to David, "You will not get in here; even the blind and the lame can ward you off." They thought, "David cannot get in here."
2SAM|5|7|Nevertheless, David captured the fortress of Zion, the City of David.
2SAM|5|8|On that day, David said, "Anyone who conquers the Jebusites will have to use the water shaft to reach those 'lame and blind' who are David's enemies. "That is why they say, "The 'blind and lame' will not enter the palace."
2SAM|5|9|David then took up residence in the fortress and called it the City of David. He built up the area around it, from the supporting terraces inward.
2SAM|5|10|And he became more and more powerful, because the LORD God Almighty was with him.
2SAM|5|11|Now Hiram king of Tyre sent messengers to David, along with cedar logs and carpenters and stonemasons, and they built a palace for David.
2SAM|5|12|And David knew that the LORD had established him as king over Israel and had exalted his kingdom for the sake of his people Israel.
2SAM|5|13|After he left Hebron, David took more concubines and wives in Jerusalem, and more sons and daughters were born to him.
2SAM|5|14|These are the names of the children born to him there: Shammua, Shobab, Nathan, Solomon,
2SAM|5|15|Ibhar, Elishua, Nepheg, Japhia,
2SAM|5|16|Elishama, Eliada and Eliphelet.
2SAM|5|17|When the Philistines heard that David had been anointed king over Israel, they went up in full force to search for him, but David heard about it and went down to the stronghold.
2SAM|5|18|Now the Philistines had come and spread out in the Valley of Rephaim;
2SAM|5|19|so David inquired of the LORD, "Shall I go and attack the Philistines? Will you hand them over to me?" The LORD answered him, "Go, for I will surely hand the Philistines over to you."
2SAM|5|20|So David went to Baal Perazim, and there he defeated them. He said, "As waters break out, the LORD has broken out against my enemies before me." So that place was called Baal Perazim.
2SAM|5|21|The Philistines abandoned their idols there, and David and his men carried them off.
2SAM|5|22|Once more the Philistines came up and spread out in the Valley of Rephaim;
2SAM|5|23|so David inquired of the LORD, and he answered, "Do not go straight up, but circle around behind them and attack them in front of the balsam trees.
2SAM|5|24|As soon as you hear the sound of marching in the tops of the balsam trees, move quickly, because that will mean the LORD has gone out in front of you to strike the Philistine army."
2SAM|5|25|So David did as the LORD commanded him, and he struck down the Philistines all the way from Gibeon to Gezer.
2SAM|6|1|David again brought together out of Israel chosen men, thirty thousand in all.
2SAM|6|2|He and all his men set out from Baalah of Judah to bring up from there the ark of God, which is called by the Name, the name of the LORD Almighty, who is enthroned between the cherubim that are on the ark.
2SAM|6|3|They set the ark of God on a new cart and brought it from the house of Abinadab, which was on the hill. Uzzah and Ahio, sons of Abinadab, were guiding the new cart
2SAM|6|4|with the ark of God on it, and Ahio was walking in front of it.
2SAM|6|5|David and the whole house of Israel were celebrating with all their might before the LORD, with songs and with harps, lyres, tambourines, sistrums and cymbals.
2SAM|6|6|When they came to the threshing floor of Nacon, Uzzah reached out and took hold of the ark of God, because the oxen stumbled.
2SAM|6|7|The LORD's anger burned against Uzzah because of his irreverent act; therefore God struck him down and he died there beside the ark of God.
2SAM|6|8|Then David was angry because the LORD's wrath had broken out against Uzzah, and to this day that place is called Perez Uzzah.
2SAM|6|9|David was afraid of the LORD that day and said, "How can the ark of the LORD ever come to me?"
2SAM|6|10|He was not willing to take the ark of the LORD to be with him in the City of David. Instead, he took it aside to the house of Obed-Edom the Gittite.
2SAM|6|11|The ark of the LORD remained in the house of Obed-Edom the Gittite for three months, and the LORD blessed him and his entire household.
2SAM|6|12|Now King David was told, "The LORD has blessed the household of Obed-Edom and everything he has, because of the ark of God." So David went down and brought up the ark of God from the house of Obed-Edom to the City of David with rejoicing.
2SAM|6|13|When those who were carrying the ark of the LORD had taken six steps, he sacrificed a bull and a fattened calf.
2SAM|6|14|David, wearing a linen ephod, danced before the LORD with all his might,
2SAM|6|15|while he and the entire house of Israel brought up the ark of the LORD with shouts and the sound of trumpets.
2SAM|6|16|As the ark of the LORD was entering the City of David, Michal daughter of Saul watched from a window. And when she saw King David leaping and dancing before the LORD, she despised him in her heart.
2SAM|6|17|They brought the ark of the LORD and set it in its place inside the tent that David had pitched for it, and David sacrificed burnt offerings and fellowship offerings before the LORD.
2SAM|6|18|After he had finished sacrificing the burnt offerings and fellowship offerings, he blessed the people in the name of the LORD Almighty.
2SAM|6|19|Then he gave a loaf of bread, a cake of dates and a cake of raisins to each person in the whole crowd of Israelites, both men and women. And all the people went to their homes.
2SAM|6|20|When David returned home to bless his household, Michal daughter of Saul came out to meet him and said, "How the king of Israel has distinguished himself today, disrobing in the sight of the slave girls of his servants as any vulgar fellow would!"
2SAM|6|21|David said to Michal, "It was before the LORD, who chose me rather than your father or anyone from his house when he appointed me ruler over the LORD's people Israel-I will celebrate before the LORD.
2SAM|6|22|I will become even more undignified than this, and I will be humiliated in my own eyes. But by these slave girls you spoke of, I will be held in honor."
2SAM|6|23|And Michal daughter of Saul had no children to the day of her death.
2SAM|7|1|After the king was settled in his palace and the LORD had given him rest from all his enemies around him,
2SAM|7|2|he said to Nathan the prophet, "Here I am, living in a palace of cedar, while the ark of God remains in a tent."
2SAM|7|3|Nathan replied to the king, "Whatever you have in mind, go ahead and do it, for the LORD is with you."
2SAM|7|4|That night the word of the LORD came to Nathan, saying:
2SAM|7|5|"Go and tell my servant David, 'This is what the LORD says: Are you the one to build me a house to dwell in?
2SAM|7|6|I have not dwelt in a house from the day I brought the Israelites up out of Egypt to this day. I have been moving from place to place with a tent as my dwelling.
2SAM|7|7|Wherever I have moved with all the Israelites, did I ever say to any of their rulers whom I commanded to shepherd my people Israel, "Why have you not built me a house of cedar?"'
2SAM|7|8|"Now then, tell my servant David, 'This is what the LORD Almighty says: I took you from the pasture and from following the flock to be ruler over my people Israel.
2SAM|7|9|I have been with you wherever you have gone, and I have cut off all your enemies from before you. Now I will make your name great, like the names of the greatest men of the earth.
2SAM|7|10|And I will provide a place for my people Israel and will plant them so that they can have a home of their own and no longer be disturbed. Wicked people will not oppress them anymore, as they did at the beginning
2SAM|7|11|and have done ever since the time I appointed leaders over my people Israel. I will also give you rest from all your enemies. "'The LORD declares to you that the LORD himself will establish a house for you:
2SAM|7|12|When your days are over and you rest with your fathers, I will raise up your offspring to succeed you, who will come from your own body, and I will establish his kingdom.
2SAM|7|13|He is the one who will build a house for my Name, and I will establish the throne of his kingdom forever.
2SAM|7|14|I will be his father, and he will be my son. When he does wrong, I will punish him with the rod of men, with floggings inflicted by men.
2SAM|7|15|But my love will never be taken away from him, as I took it away from Saul, whom I removed from before you.
2SAM|7|16|Your house and your kingdom will endure forever before me; your throne will be established forever.'"
2SAM|7|17|Nathan reported to David all the words of this entire revelation.
2SAM|7|18|Then King David went in and sat before the LORD, and he said: "Who am I, O Sovereign LORD, and what is my family, that you have brought me this far?
2SAM|7|19|And as if this were not enough in your sight, O Sovereign LORD, you have also spoken about the future of the house of your servant. Is this your usual way of dealing with man, O Sovereign LORD?
2SAM|7|20|"What more can David say to you? For you know your servant, O Sovereign LORD.
2SAM|7|21|For the sake of your word and according to your will, you have done this great thing and made it known to your servant.
2SAM|7|22|"How great you are, O Sovereign LORD! There is no one like you, and there is no God but you, as we have heard with our own ears.
2SAM|7|23|And who is like your people Israel-the one nation on earth that God went out to redeem as a people for himself, and to make a name for himself, and to perform great and awesome wonders by driving out nations and their gods from before your people, whom you redeemed from Egypt?
2SAM|7|24|You have established your people Israel as your very own forever, and you, O LORD, have become their God.
2SAM|7|25|"And now, LORD God, keep forever the promise you have made concerning your servant and his house. Do as you promised,
2SAM|7|26|so that your name will be great forever. Then men will say, 'The LORD Almighty is God over Israel!' And the house of your servant David will be established before you.
2SAM|7|27|"O LORD Almighty, God of Israel, you have revealed this to your servant, saying, 'I will build a house for you.' So your servant has found courage to offer you this prayer.
2SAM|7|28|O Sovereign LORD, you are God! Your words are trustworthy, and you have promised these good things to your servant.
2SAM|7|29|Now be pleased to bless the house of your servant, that it may continue forever in your sight; for you, O Sovereign LORD, have spoken, and with your blessing the house of your servant will be blessed forever."
2SAM|8|1|In the course of time, David defeated the Philistines and subdued them, and he took Metheg Ammah from the control of the Philistines.
2SAM|8|2|David also defeated the Moabites. He made them lie down on the ground and measured them off with a length of cord. Every two lengths of them were put to death, and the third length was allowed to live. So the Moabites became subject to David and brought tribute.
2SAM|8|3|Moreover, David fought Hadadezer son of Rehob, king of Zobah, when he went to restore his control along the Euphrates River.
2SAM|8|4|David captured a thousand of his chariots, seven thousand charioteers and twenty thousand foot soldiers. He hamstrung all but a hundred of the chariot horses.
2SAM|8|5|When the Arameans of Damascus came to help Hadadezer king of Zobah, David struck down twenty-two thousand of them.
2SAM|8|6|He put garrisons in the Aramean kingdom of Damascus, and the Arameans became subject to him and brought tribute. The LORD gave David victory wherever he went.
2SAM|8|7|David took the gold shields that belonged to the officers of Hadadezer and brought them to Jerusalem.
2SAM|8|8|From Tebah and Berothai, towns that belonged to Hadadezer, King David took a great quantity of bronze.
2SAM|8|9|When Tou king of Hamath heard that David had defeated the entire army of Hadadezer,
2SAM|8|10|he sent his son Joram to King David to greet him and congratulate him on his victory in battle over Hadadezer, who had been at war with Tou. Joram brought with him articles of silver and gold and bronze.
2SAM|8|11|King David dedicated these articles to the LORD, as he had done with the silver and gold from all the nations he had subdued:
2SAM|8|12|Edom and Moab, the Ammonites and the Philistines, and Amalek. He also dedicated the plunder taken from Hadadezer son of Rehob, king of Zobah.
2SAM|8|13|And David became famous after he returned from striking down eighteen thousand Edomites in the Valley of Salt.
2SAM|8|14|He put garrisons throughout Edom, and all the Edomites became subject to David. The LORD gave David victory wherever he went.
2SAM|8|15|David reigned over all Israel, doing what was just and right for all his people.
2SAM|8|16|Joab son of Zeruiah was over the army; Jehoshaphat son of Ahilud was recorder;
2SAM|8|17|Zadok son of Ahitub and Ahimelech son of Abiathar were priests; Seraiah was secretary;
2SAM|8|18|Benaiah son of Jehoiada was over the Kerethites and Pelethites; and David's sons were royal advisers.
2SAM|9|1|David asked, "Is there anyone still left of the house of Saul to whom I can show kindness for Jonathan's sake?"
2SAM|9|2|Now there was a servant of Saul's household named Ziba. They called him to appear before David, and the king said to him, "Are you Ziba?Your servant," he replied.
2SAM|9|3|The king asked, "Is there no one still left of the house of Saul to whom I can show God's kindness?" Ziba answered the king, "There is still a son of Jonathan; he is crippled in both feet."
2SAM|9|4|"Where is he?" the king asked. Ziba answered, "He is at the house of Makir son of Ammiel in Lo Debar."
2SAM|9|5|So King David had him brought from Lo Debar, from the house of Makir son of Ammiel.
2SAM|9|6|When Mephibosheth son of Jonathan, the son of Saul, came to David, he bowed down to pay him honor. David said, "Mephibosheth!Your servant," he replied.
2SAM|9|7|"Don't be afraid," David said to him, "for I will surely show you kindness for the sake of your father Jonathan. I will restore to you all the land that belonged to your grandfather Saul, and you will always eat at my table."
2SAM|9|8|Mephibosheth bowed down and said, "What is your servant, that you should notice a dead dog like me?"
2SAM|9|9|Then the king summoned Ziba, Saul's servant, and said to him, "I have given your master's grandson everything that belonged to Saul and his family.
2SAM|9|10|You and your sons and your servants are to farm the land for him and bring in the crops, so that your master's grandson may be provided for. And Mephibosheth, grandson of your master, will always eat at my table." (Now Ziba had fifteen sons and twenty servants.)
2SAM|9|11|Then Ziba said to the king, "Your servant will do whatever my lord the king commands his servant to do." So Mephibosheth ate at David's table like one of the king's sons.
2SAM|9|12|Mephibosheth had a young son named Mica, and all the members of Ziba's household were servants of Mephibosheth.
2SAM|9|13|And Mephibosheth lived in Jerusalem, because he always ate at the king's table, and he was crippled in both feet.
2SAM|10|1|In the course of time, the king of the Ammonites died, and his son Hanun succeeded him as king.
2SAM|10|2|David thought, "I will show kindness to Hanun son of Nahash, just as his father showed kindness to me." So David sent a delegation to express his sympathy to Hanun concerning his father. When David's men came to the land of the Ammonites,
2SAM|10|3|the Ammonite nobles said to Hanun their lord, "Do you think David is honoring your father by sending men to you to express sympathy? Hasn't David sent them to you to explore the city and spy it out and overthrow it?"
2SAM|10|4|So Hanun seized David's men, shaved off half of each man's beard, cut off their garments in the middle at the buttocks, and sent them away.
2SAM|10|5|When David was told about this, he sent messengers to meet the men, for they were greatly humiliated. The king said, "Stay at Jericho till your beards have grown, and then come back."
2SAM|10|6|When the Ammonites realized that they had become a stench in David's nostrils, they hired twenty thousand Aramean foot soldiers from Beth Rehob and Zobah, as well as the king of Maacah with a thousand men, and also twelve thousand men from Tob.
2SAM|10|7|On hearing this, David sent Joab out with the entire army of fighting men.
2SAM|10|8|The Ammonites came out and drew up in battle formation at the entrance to their city gate, while the Arameans of Zobah and Rehob and the men of Tob and Maacah were by themselves in the open country.
2SAM|10|9|Joab saw that there were battle lines in front of him and behind him; so he selected some of the best troops in Israel and deployed them against the Arameans.
2SAM|10|10|He put the rest of the men under the command of Abishai his brother and deployed them against the Ammonites.
2SAM|10|11|Joab said, "If the Arameans are too strong for me, then you are to come to my rescue; but if the Ammonites are too strong for you, then I will come to rescue you.
2SAM|10|12|Be strong and let us fight bravely for our people and the cities of our God. The LORD will do what is good in his sight."
2SAM|10|13|Then Joab and the troops with him advanced to fight the Arameans, and they fled before him.
2SAM|10|14|When the Ammonites saw that the Arameans were fleeing, they fled before Abishai and went inside the city. So Joab returned from fighting the Ammonites and came to Jerusalem.
2SAM|10|15|After the Arameans saw that they had been routed by Israel, they regrouped.
2SAM|10|16|Hadadezer had Arameans brought from beyond the River; they went to Helam, with Shobach the commander of Hadadezer's army leading them.
2SAM|10|17|When David was told of this, he gathered all Israel, crossed the Jordan and went to Helam. The Arameans formed their battle lines to meet David and fought against him.
2SAM|10|18|But they fled before Israel, and David killed seven hundred of their charioteers and forty thousand of their foot soldiers. He also struck down Shobach the commander of their army, and he died there.
2SAM|10|19|When all the kings who were vassals of Hadadezer saw that they had been defeated by Israel, they made peace with the Israelites and became subject to them. So the Arameans were afraid to help the Ammonites anymore.
2SAM|11|1|In the spring, at the time when kings go off to war, David sent Joab out with the king's men and the whole Israelite army. They destroyed the Ammonites and besieged Rabbah. But David remained in Jerusalem.
2SAM|11|2|One evening David got up from his bed and walked around on the roof of the palace. From the roof he saw a woman bathing. The woman was very beautiful,
2SAM|11|3|and David sent someone to find out about her. The man said, "Isn't this Bathsheba, the daughter of Eliam and the wife of Uriah the Hittite?"
2SAM|11|4|Then David sent messengers to get her. She came to him, and he slept with her. (She had purified herself from her uncleanness.) Then she went back home.
2SAM|11|5|The woman conceived and sent word to David, saying, "I am pregnant."
2SAM|11|6|So David sent this word to Joab: "Send me Uriah the Hittite." And Joab sent him to David.
2SAM|11|7|When Uriah came to him, David asked him how Joab was, how the soldiers were and how the war was going.
2SAM|11|8|Then David said to Uriah, "Go down to your house and wash your feet." So Uriah left the palace, and a gift from the king was sent after him.
2SAM|11|9|But Uriah slept at the entrance to the palace with all his master's servants and did not go down to his house.
2SAM|11|10|When David was told, "Uriah did not go home," he asked him, "Haven't you just come from a distance? Why didn't you go home?"
2SAM|11|11|Uriah said to David, "The ark and Israel and Judah are staying in tents, and my master Joab and my lord's men are camped in the open fields. How could I go to my house to eat and drink and lie with my wife? As surely as you live, I will not do such a thing!"
2SAM|11|12|Then David said to him, "Stay here one more day, and tomorrow I will send you back." So Uriah remained in Jerusalem that day and the next.
2SAM|11|13|At David's invitation, he ate and drank with him, and David made him drunk. But in the evening Uriah went out to sleep on his mat among his master's servants; he did not go home.
2SAM|11|14|In the morning David wrote a letter to Joab and sent it with Uriah.
2SAM|11|15|In it he wrote, "Put Uriah in the front line where the fighting is fiercest. Then withdraw from him so he will be struck down and die."
2SAM|11|16|So while Joab had the city under siege, he put Uriah at a place where he knew the strongest defenders were.
2SAM|11|17|When the men of the city came out and fought against Joab, some of the men in David's army fell; moreover, Uriah the Hittite died.
2SAM|11|18|Joab sent David a full account of the battle.
2SAM|11|19|He instructed the messenger: "When you have finished giving the king this account of the battle,
2SAM|11|20|the king's anger may flare up, and he may ask you, 'Why did you get so close to the city to fight? Didn't you know they would shoot arrows from the wall?
2SAM|11|21|Who killed Abimelech son of Jerub-Besheth? Didn't a woman throw an upper millstone on him from the wall, so that he died in Thebez? Why did you get so close to the wall?' If he asks you this, then say to him, 'Also, your servant Uriah the Hittite is dead.'"
2SAM|11|22|The messenger set out, and when he arrived he told David everything Joab had sent him to say.
2SAM|11|23|The messenger said to David, "The men overpowered us and came out against us in the open, but we drove them back to the entrance to the city gate.
2SAM|11|24|Then the archers shot arrows at your servants from the wall, and some of the king's men died. Moreover, your servant Uriah the Hittite is dead."
2SAM|11|25|David told the messenger, "Say this to Joab: 'Don't let this upset you; the sword devours one as well as another. Press the attack against the city and destroy it.' Say this to encourage Joab."
2SAM|11|26|When Uriah's wife heard that her husband was dead, she mourned for him.
2SAM|11|27|After the time of mourning was over, David had her brought to his house, and she became his wife and bore him a son. But the thing David had done displeased the LORD.
2SAM|12|1|The LORD sent Nathan to David. When he came to him, he said, "There were two men in a certain town, one rich and the other poor.
2SAM|12|2|The rich man had a very large number of sheep and cattle,
2SAM|12|3|but the poor man had nothing except one little ewe lamb he had bought. He raised it, and it grew up with him and his children. It shared his food, drank from his cup and even slept in his arms. It was like a daughter to him.
2SAM|12|4|"Now a traveler came to the rich man, but the rich man refrained from taking one of his own sheep or cattle to prepare a meal for the traveler who had come to him. Instead, he took the ewe lamb that belonged to the poor man and prepared it for the one who had come to him."
2SAM|12|5|David burned with anger against the man and said to Nathan, "As surely as the LORD lives, the man who did this deserves to die!
2SAM|12|6|He must pay for that lamb four times over, because he did such a thing and had no pity."
2SAM|12|7|Then Nathan said to David, "You are the man! This is what the LORD, the God of Israel, says: 'I anointed you king over Israel, and I delivered you from the hand of Saul.
2SAM|12|8|I gave your master's house to you, and your master's wives into your arms. I gave you the house of Israel and Judah. And if all this had been too little, I would have given you even more.
2SAM|12|9|Why did you despise the word of the LORD by doing what is evil in his eyes? You struck down Uriah the Hittite with the sword and took his wife to be your own. You killed him with the sword of the Ammonites.
2SAM|12|10|Now, therefore, the sword will never depart from your house, because you despised me and took the wife of Uriah the Hittite to be your own.'
2SAM|12|11|"This is what the LORD says: 'Out of your own household I am going to bring calamity upon you. Before your very eyes I will take your wives and give them to one who is close to you, and he will lie with your wives in broad daylight.
2SAM|12|12|You did it in secret, but I will do this thing in broad daylight before all Israel.'"
2SAM|12|13|Then David said to Nathan, "I have sinned against the LORD." Nathan replied, "The LORD has taken away your sin. You are not going to die.
2SAM|12|14|But because by doing this you have made the enemies of the LORD show utter contempt, the son born to you will die."
2SAM|12|15|After Nathan had gone home, the LORD struck the child that Uriah's wife had borne to David, and he became ill.
2SAM|12|16|David pleaded with God for the child. He fasted and went into his house and spent the nights lying on the ground.
2SAM|12|17|The elders of his household stood beside him to get him up from the ground, but he refused, and he would not eat any food with them.
2SAM|12|18|On the seventh day the child died. David's servants were afraid to tell him that the child was dead, for they thought, "While the child was still living, we spoke to David but he would not listen to us. How can we tell him the child is dead? He may do something desperate."
2SAM|12|19|David noticed that his servants were whispering among themselves and he realized the child was dead. "Is the child dead?" he asked. "Yes," they replied, "he is dead."
2SAM|12|20|Then David got up from the ground. After he had washed, put on lotions and changed his clothes, he went into the house of the LORD and worshiped. Then he went to his own house, and at his request they served him food, and he ate.
2SAM|12|21|His servants asked him, "Why are you acting this way? While the child was alive, you fasted and wept, but now that the child is dead, you get up and eat!"
2SAM|12|22|He answered, "While the child was still alive, I fasted and wept. I thought, 'Who knows? The LORD may be gracious to me and let the child live.'
2SAM|12|23|But now that he is dead, why should I fast? Can I bring him back again? I will go to him, but he will not return to me."
2SAM|12|24|Then David comforted his wife Bathsheba, and he went to her and lay with her. She gave birth to a son, and they named him Solomon. The LORD loved him;
2SAM|12|25|and because the LORD loved him, he sent word through Nathan the prophet to name him Jedidiah.
2SAM|12|26|Meanwhile Joab fought against Rabbah of the Ammonites and captured the royal citadel.
2SAM|12|27|Joab then sent messengers to David, saying, "I have fought against Rabbah and taken its water supply.
2SAM|12|28|Now muster the rest of the troops and besiege the city and capture it. Otherwise I will take the city, and it will be named after me."
2SAM|12|29|So David mustered the entire army and went to Rabbah, and attacked and captured it.
2SAM|12|30|He took the crown from the head of their king -its weight was a talent of gold, and it was set with precious stones-and it was placed on David's head. He took a great quantity of plunder from the city
2SAM|12|31|and brought out the people who were there, consigning them to labor with saws and with iron picks and axes, and he made them work at brickmaking. He did this to all the Ammonite towns. Then David and his entire army returned to Jerusalem.
2SAM|13|1|In the course of time, Amnon son of David fell in love with Tamar, the beautiful sister of Absalom son of David.
2SAM|13|2|Amnon became frustrated to the point of illness on account of his sister Tamar, for she was a virgin, and it seemed impossible for him to do anything to her.
2SAM|13|3|Now Amnon had a friend named Jonadab son of Shimeah, David's brother. Jonadab was a very shrewd man.
2SAM|13|4|He asked Amnon, "Why do you, the king's son, look so haggard morning after morning? Won't you tell me?" Amnon said to him, "I'm in love with Tamar, my brother Absalom's sister."
2SAM|13|5|"Go to bed and pretend to be ill," Jonadab said. "When your father comes to see you, say to him, 'I would like my sister Tamar to come and give me something to eat. Let her prepare the food in my sight so I may watch her and then eat it from her hand.'"
2SAM|13|6|So Amnon lay down and pretended to be ill. When the king came to see him, Amnon said to him, "I would like my sister Tamar to come and make some special bread in my sight, so I may eat from her hand."
2SAM|13|7|David sent word to Tamar at the palace: "Go to the house of your brother Amnon and prepare some food for him."
2SAM|13|8|So Tamar went to the house of her brother Amnon, who was lying down. She took some dough, kneaded it, made the bread in his sight and baked it.
2SAM|13|9|Then she took the pan and served him the bread, but he refused to eat. "Send everyone out of here," Amnon said. So everyone left him.
2SAM|13|10|Then Amnon said to Tamar, "Bring the food here into my bedroom so I may eat from your hand." And Tamar took the bread she had prepared and brought it to her brother Amnon in his bedroom.
2SAM|13|11|But when she took it to him to eat, he grabbed her and said, "Come to bed with me, my sister."
2SAM|13|12|"Don't, my brother!" she said to him. "Don't force me. Such a thing should not be done in Israel! Don't do this wicked thing.
2SAM|13|13|What about me? Where could I get rid of my disgrace? And what about you? You would be like one of the wicked fools in Israel. Please speak to the king; he will not keep me from being married to you."
2SAM|13|14|But he refused to listen to her, and since he was stronger than she, he raped her.
2SAM|13|15|Then Amnon hated her with intense hatred. In fact, he hated her more than he had loved her. Amnon said to her, "Get up and get out!"
2SAM|13|16|"No!" she said to him. "Sending me away would be a greater wrong than what you have already done to me." But he refused to listen to her.
2SAM|13|17|He called his personal servant and said, "Get this woman out of here and bolt the door after her."
2SAM|13|18|So his servant put her out and bolted the door after her. She was wearing a richly ornamented robe, for this was the kind of garment the virgin daughters of the king wore.
2SAM|13|19|Tamar put ashes on her head and tore the ornamented robe she was wearing. She put her hand on her head and went away, weeping aloud as she went.
2SAM|13|20|Her brother Absalom said to her, "Has that Amnon, your brother, been with you? Be quiet now, my sister; he is your brother. Don't take this thing to heart." And Tamar lived in her brother Absalom's house, a desolate woman.
2SAM|13|21|When King David heard all this, he was furious.
2SAM|13|22|Absalom never said a word to Amnon, either good or bad; he hated Amnon because he had disgraced his sister Tamar.
2SAM|13|23|Two years later, when Absalom's sheepshearers were at Baal Hazor near the border of Ephraim, he invited all the king's sons to come there.
2SAM|13|24|Absalom went to the king and said, "Your servant has had shearers come. Will the king and his officials please join me?"
2SAM|13|25|"No, my son," the king replied. "All of us should not go; we would only be a burden to you." Although Absalom urged him, he still refused to go, but gave him his blessing.
2SAM|13|26|Then Absalom said, "If not, please let my brother Amnon come with us." The king asked him, "Why should he go with you?"
2SAM|13|27|But Absalom urged him, so he sent with him Amnon and the rest of the king's sons.
2SAM|13|28|Absalom ordered his men, "Listen! When Amnon is in high spirits from drinking wine and I say to you, 'Strike Amnon down,' then kill him. Don't be afraid. Have not I given you this order? Be strong and brave."
2SAM|13|29|So Absalom's men did to Amnon what Absalom had ordered. Then all the king's sons got up, mounted their mules and fled.
2SAM|13|30|While they were on their way, the report came to David: "Absalom has struck down all the king's sons; not one of them is left."
2SAM|13|31|The king stood up, tore his clothes and lay down on the ground; and all his servants stood by with their clothes torn.
2SAM|13|32|But Jonadab son of Shimeah, David's brother, said, "My lord should not think that they killed all the princes; only Amnon is dead. This has been Absalom's expressed intention ever since the day Amnon raped his sister Tamar.
2SAM|13|33|My lord the king should not be concerned about the report that all the king's sons are dead. Only Amnon is dead."
2SAM|13|34|Meanwhile, Absalom had fled. Now the man standing watch looked up and saw many people on the road west of him, coming down the side of the hill. The watchman went and told the king, "I see men in the direction of Horonaim, on the side of the hill."
2SAM|13|35|Jonadab said to the king, "See, the king's sons are here; it has happened just as your servant said."
2SAM|13|36|As he finished speaking, the king's sons came in, wailing loudly. The king, too, and all his servants wept very bitterly.
2SAM|13|37|Absalom fled and went to Talmai son of Ammihud, the king of Geshur. But King David mourned for his son every day.
2SAM|13|38|After Absalom fled and went to Geshur, he stayed there three years.
2SAM|13|39|And the spirit of the king longed to go to Absalom, for he was consoled concerning Amnon's death.
2SAM|14|1|Joab son of Zeruiah knew that the king's heart longed for Absalom.
2SAM|14|2|So Joab sent someone to Tekoa and had a wise woman brought from there. He said to her, "Pretend you are in mourning. Dress in mourning clothes, and don't use any cosmetic lotions. Act like a woman who has spent many days grieving for the dead.
2SAM|14|3|Then go to the king and speak these words to him." And Joab put the words in her mouth.
2SAM|14|4|When the woman from Tekoa went to the king, she fell with her face to the ground to pay him honor, and she said, "Help me, O king!"
2SAM|14|5|The king asked her, "What is troubling you?" She said, "I am indeed a widow; my husband is dead.
2SAM|14|6|I your servant had two sons. They got into a fight with each other in the field, and no one was there to separate them. One struck the other and killed him.
2SAM|14|7|Now the whole clan has risen up against your servant; they say, 'Hand over the one who struck his brother down, so that we may put him to death for the life of his brother whom he killed; then we will get rid of the heir as well.' They would put out the only burning coal I have left, leaving my husband neither name nor descendant on the face of the earth."
2SAM|14|8|The king said to the woman, "Go home, and I will issue an order in your behalf."
2SAM|14|9|But the woman from Tekoa said to him, "My lord the king, let the blame rest on me and on my father's family, and let the king and his throne be without guilt."
2SAM|14|10|The king replied, "If anyone says anything to you, bring him to me, and he will not bother you again."
2SAM|14|11|She said, "Then let the king invoke the LORD his God to prevent the avenger of blood from adding to the destruction, so that my son will not be destroyed.As surely as the LORD lives," he said, "not one hair of your son's head will fall to the ground."
2SAM|14|12|Then the woman said, "Let your servant speak a word to my lord the king.Speak," he replied.
2SAM|14|13|The woman said, "Why then have you devised a thing like this against the people of God? When the king says this, does he not convict himself, for the king has not brought back his banished son?
2SAM|14|14|Like water spilled on the ground, which cannot be recovered, so we must die. But God does not take away life; instead, he devises ways so that a banished person may not remain estranged from him.
2SAM|14|15|"And now I have come to say this to my lord the king because the people have made me afraid. Your servant thought, 'I will speak to the king; perhaps he will do what his servant asks.
2SAM|14|16|Perhaps the king will agree to deliver his servant from the hand of the man who is trying to cut off both me and my son from the inheritance God gave us.'
2SAM|14|17|"And now your servant says, 'May the word of my lord the king bring me rest, for my lord the king is like an angel of God in discerning good and evil. May the LORD your God be with you.'"
2SAM|14|18|Then the king said to the woman, "Do not keep from me the answer to what I am going to ask you.Let my lord the king speak," the woman said.
2SAM|14|19|The king asked, "Isn't the hand of Joab with you in all this?" The woman answered, "As surely as you live, my lord the king, no one can turn to the right or to the left from anything my lord the king says. Yes, it was your servant Joab who instructed me to do this and who put all these words into the mouth of your servant.
2SAM|14|20|Your servant Joab did this to change the present situation. My lord has wisdom like that of an angel of God-he knows everything that happens in the land."
2SAM|14|21|The king said to Joab, "Very well, I will do it. Go, bring back the young man Absalom."
2SAM|14|22|Joab fell with his face to the ground to pay him honor, and he blessed the king. Joab said, "Today your servant knows that he has found favor in your eyes, my lord the king, because the king has granted his servant's request."
2SAM|14|23|Then Joab went to Geshur and brought Absalom back to Jerusalem.
2SAM|14|24|But the king said, "He must go to his own house; he must not see my face." So Absalom went to his own house and did not see the face of the king.
2SAM|14|25|In all Israel there was not a man so highly praised for his handsome appearance as Absalom. From the top of his head to the sole of his foot there was no blemish in him.
2SAM|14|26|Whenever he cut the hair of his head-he used to cut his hair from time to time when it became too heavy for him-he would weigh it, and its weight was two hundred shekels by the royal standard.
2SAM|14|27|Three sons and a daughter were born to Absalom. The daughter's name was Tamar, and she became a beautiful woman.
2SAM|14|28|Absalom lived two years in Jerusalem without seeing the king's face.
2SAM|14|29|Then Absalom sent for Joab in order to send him to the king, but Joab refused to come to him. So he sent a second time, but he refused to come.
2SAM|14|30|Then he said to his servants, "Look, Joab's field is next to mine, and he has barley there. Go and set it on fire." So Absalom's servants set the field on fire.
2SAM|14|31|Then Joab did go to Absalom's house and he said to him, "Why have your servants set my field on fire?"
2SAM|14|32|Absalom said to Joab, "Look, I sent word to you and said, 'Come here so I can send you to the king to ask, "Why have I come from Geshur? It would be better for me if I were still there!"' Now then, I want to see the king's face, and if I am guilty of anything, let him put me to death."
2SAM|14|33|So Joab went to the king and told him this. Then the king summoned Absalom, and he came in and bowed down with his face to the ground before the king. And the king kissed Absalom.
2SAM|15|1|In the course of time, Absalom provided himself with a chariot and horses and with fifty men to run ahead of him.
2SAM|15|2|He would get up early and stand by the side of the road leading to the city gate. Whenever anyone came with a complaint to be placed before the king for a decision, Absalom would call out to him, "What town are you from?" He would answer, "Your servant is from one of the tribes of Israel."
2SAM|15|3|Then Absalom would say to him, "Look, your claims are valid and proper, but there is no representative of the king to hear you."
2SAM|15|4|And Absalom would add, "If only I were appointed judge in the land! Then everyone who has a complaint or case could come to me and I would see that he gets justice."
2SAM|15|5|Also, whenever anyone approached him to bow down before him, Absalom would reach out his hand, take hold of him and kiss him.
2SAM|15|6|Absalom behaved in this way toward all the Israelites who came to the king asking for justice, and so he stole the hearts of the men of Israel.
2SAM|15|7|At the end of four years, Absalom said to the king, "Let me go to Hebron and fulfill a vow I made to the LORD.
2SAM|15|8|While your servant was living at Geshur in Aram, I made this vow: 'If the LORD takes me back to Jerusalem, I will worship the LORD in Hebron. '"
2SAM|15|9|The king said to him, "Go in peace." So he went to Hebron.
2SAM|15|10|Then Absalom sent secret messengers throughout the tribes of Israel to say, "As soon as you hear the sound of the trumpets, then say, 'Absalom is king in Hebron.'"
2SAM|15|11|Two hundred men from Jerusalem had accompanied Absalom. They had been invited as guests and went quite innocently, knowing nothing about the matter.
2SAM|15|12|While Absalom was offering sacrifices, he also sent for Ahithophel the Gilonite, David's counselor, to come from Giloh, his hometown. And so the conspiracy gained strength, and Absalom's following kept on increasing.
2SAM|15|13|A messenger came and told David, "The hearts of the men of Israel are with Absalom."
2SAM|15|14|Then David said to all his officials who were with him in Jerusalem, "Come! We must flee, or none of us will escape from Absalom. We must leave immediately, or he will move quickly to overtake us and bring ruin upon us and put the city to the sword."
2SAM|15|15|The king's officials answered him, "Your servants are ready to do whatever our lord the king chooses."
2SAM|15|16|The king set out, with his entire household following him; but he left ten concubines to take care of the palace.
2SAM|15|17|So the king set out, with all the people following him, and they halted at a place some distance away.
2SAM|15|18|All his men marched past him, along with all the Kerethites and Pelethites; and all the six hundred Gittites who had accompanied him from Gath marched before the king.
2SAM|15|19|The king said to Ittai the Gittite, "Why should you come along with us? Go back and stay with King Absalom. You are a foreigner, an exile from your homeland.
2SAM|15|20|You came only yesterday. And today shall I make you wander about with us, when I do not know where I am going? Go back, and take your countrymen. May kindness and faithfulness be with you."
2SAM|15|21|But Ittai replied to the king, "As surely as the LORD lives, and as my lord the king lives, wherever my lord the king may be, whether it means life or death, there will your servant be."
2SAM|15|22|David said to Ittai, "Go ahead, march on." So Ittai the Gittite marched on with all his men and the families that were with him.
2SAM|15|23|The whole countryside wept aloud as all the people passed by. The king also crossed the Kidron Valley, and all the people moved on toward the desert.
2SAM|15|24|Zadok was there, too, and all the Levites who were with him were carrying the ark of the covenant of God. They set down the ark of God, and Abiathar offered sacrifices until all the people had finished leaving the city.
2SAM|15|25|Then the king said to Zadok, "Take the ark of God back into the city. If I find favor in the LORD's eyes, he will bring me back and let me see it and his dwelling place again.
2SAM|15|26|But if he says, 'I am not pleased with you,' then I am ready; let him do to me whatever seems good to him."
2SAM|15|27|The king also said to Zadok the priest, "Aren't you a seer? Go back to the city in peace, with your son Ahimaaz and Jonathan son of Abiathar. You and Abiathar take your two sons with you.
2SAM|15|28|I will wait at the fords in the desert until word comes from you to inform me."
2SAM|15|29|So Zadok and Abiathar took the ark of God back to Jerusalem and stayed there.
2SAM|15|30|But David continued up the Mount of Olives, weeping as he went; his head was covered and he was barefoot. All the people with him covered their heads too and were weeping as they went up.
2SAM|15|31|Now David had been told, "Ahithophel is among the conspirators with Absalom." So David prayed, "O LORD, turn Ahithophel's counsel into foolishness."
2SAM|15|32|When David arrived at the summit, where people used to worship God, Hushai the Arkite was there to meet him, his robe torn and dust on his head.
2SAM|15|33|David said to him, "If you go with me, you will be a burden to me.
2SAM|15|34|But if you return to the city and say to Absalom, 'I will be your servant, O king; I was your father's servant in the past, but now I will be your servant,' then you can help me by frustrating Ahithophel's advice.
2SAM|15|35|Won't the priests Zadok and Abiathar be there with you? Tell them anything you hear in the king's palace.
2SAM|15|36|Their two sons, Ahimaaz son of Zadok and Jonathan son of Abiathar, are there with them. Send them to me with anything you hear."
2SAM|15|37|So David's friend Hushai arrived at Jerusalem as Absalom was entering the city.
2SAM|16|1|When David had gone a short distance beyond the summit, there was Ziba, the steward of Mephibosheth, waiting to meet him. He had a string of donkeys saddled and loaded with two hundred loaves of bread, a hundred cakes of raisins, a hundred cakes of figs and a skin of wine.
2SAM|16|2|The king asked Ziba, "Why have you brought these?" Ziba answered, "The donkeys are for the king's household to ride on, the bread and fruit are for the men to eat, and the wine is to refresh those who become exhausted in the desert."
2SAM|16|3|The king then asked, "Where is your master's grandson?" Ziba said to him, "He is staying in Jerusalem, because he thinks, 'Today the house of Israel will give me back my grandfather's kingdom.'"
2SAM|16|4|Then the king said to Ziba, "All that belonged to Mephibosheth is now yours.I humbly bow," Ziba said. "May I find favor in your eyes, my lord the king."
2SAM|16|5|As King David approached Bahurim, a man from the same clan as Saul's family came out from there. His name was Shimei son of Gera, and he cursed as he came out.
2SAM|16|6|He pelted David and all the king's officials with stones, though all the troops and the special guard were on David's right and left.
2SAM|16|7|As he cursed, Shimei said, "Get out, get out, you man of blood, you scoundrel!
2SAM|16|8|The LORD has repaid you for all the blood you shed in the household of Saul, in whose place you have reigned. The LORD has handed the kingdom over to your son Absalom. You have come to ruin because you are a man of blood!"
2SAM|16|9|Then Abishai son of Zeruiah said to the king, "Why should this dead dog curse my lord the king? Let me go over and cut off his head."
2SAM|16|10|But the king said, "What do you and I have in common, you sons of Zeruiah? If he is cursing because the LORD said to him, 'Curse David,' who can ask, 'Why do you do this?'"
2SAM|16|11|David then said to Abishai and all his officials, "My son, who is of my own flesh, is trying to take my life. How much more, then, this Benjamite! Leave him alone; let him curse, for the LORD has told him to.
2SAM|16|12|It may be that the LORD will see my distress and repay me with good for the cursing I am receiving today."
2SAM|16|13|So David and his men continued along the road while Shimei was going along the hillside opposite him, cursing as he went and throwing stones at him and showering him with dirt.
2SAM|16|14|The king and all the people with him arrived at their destination exhausted. And there he refreshed himself.
2SAM|16|15|Meanwhile, Absalom and all the men of Israel came to Jerusalem, and Ahithophel was with him.
2SAM|16|16|Then Hushai the Arkite, David's friend, went to Absalom and said to him, "Long live the king! Long live the king!"
2SAM|16|17|Absalom asked Hushai, "Is this the love you show your friend? Why didn't you go with your friend?"
2SAM|16|18|Hushai said to Absalom, "No, the one chosen by the LORD, by these people, and by all the men of Israel-his I will be, and I will remain with him.
2SAM|16|19|Furthermore, whom should I serve? Should I not serve the son? Just as I served your father, so I will serve you."
2SAM|16|20|Absalom said to Ahithophel, "Give us your advice. What should we do?"
2SAM|16|21|Ahithophel answered, "Lie with your father's concubines whom he left to take care of the palace. Then all Israel will hear that you have made yourself a stench in your father's nostrils, and the hands of everyone with you will be strengthened."
2SAM|16|22|So they pitched a tent for Absalom on the roof, and he lay with his father's concubines in the sight of all Israel.
2SAM|16|23|Now in those days the advice Ahithophel gave was like that of one who inquires of God. That was how both David and Absalom regarded all of Ahithophel's advice.
2SAM|17|1|Ahithophel said to Absalom, "I would choose twelve thousand men and set out tonight in pursuit of David.
2SAM|17|2|I would attack him while he is weary and weak. I would strike him with terror, and then all the people with him will flee. I would strike down only the king
2SAM|17|3|and bring all the people back to you. The death of the man you seek will mean the return of all; all the people will be unharmed."
2SAM|17|4|This plan seemed good to Absalom and to all the elders of Israel.
2SAM|17|5|But Absalom said, "Summon also Hushai the Arkite, so we can hear what he has to say."
2SAM|17|6|When Hushai came to him, Absalom said, "Ahithophel has given this advice. Should we do what he says? If not, give us your opinion."
2SAM|17|7|Hushai replied to Absalom, "The advice Ahithophel has given is not good this time.
2SAM|17|8|You know your father and his men; they are fighters, and as fierce as a wild bear robbed of her cubs. Besides, your father is an experienced fighter; he will not spend the night with the troops.
2SAM|17|9|Even now, he is hidden in a cave or some other place. If he should attack your troops first, whoever hears about it will say, 'There has been a slaughter among the troops who follow Absalom.'
2SAM|17|10|Then even the bravest soldier, whose heart is like the heart of a lion, will melt with fear, for all Israel knows that your father is a fighter and that those with him are brave.
2SAM|17|11|"So I advise you: Let all Israel, from Dan to Beersheba-as numerous as the sand on the seashore-be gathered to you, with you yourself leading them into battle.
2SAM|17|12|Then we will attack him wherever he may be found, and we will fall on him as dew settles on the ground. Neither he nor any of his men will be left alive.
2SAM|17|13|If he withdraws into a city, then all Israel will bring ropes to that city, and we will drag it down to the valley until not even a piece of it can be found."
2SAM|17|14|Absalom and all the men of Israel said, "The advice of Hushai the Arkite is better than that of Ahithophel." For the LORD had determined to frustrate the good advice of Ahithophel in order to bring disaster on Absalom.
2SAM|17|15|Hushai told Zadok and Abiathar, the priests, "Ahithophel has advised Absalom and the elders of Israel to do such and such, but I have advised them to do so and so.
2SAM|17|16|Now send a message immediately and tell David, 'Do not spend the night at the fords in the desert; cross over without fail, or the king and all the people with him will be swallowed up.'"
2SAM|17|17|Jonathan and Ahimaaz were staying at En Rogel. A servant girl was to go and inform them, and they were to go and tell King David, for they could not risk being seen entering the city.
2SAM|17|18|But a young man saw them and told Absalom. So the two of them left quickly and went to the house of a man in Bahurim. He had a well in his courtyard, and they climbed down into it.
2SAM|17|19|His wife took a covering and spread it out over the opening of the well and scattered grain over it. No one knew anything about it.
2SAM|17|20|When Absalom's men came to the woman at the house, they asked, "Where are Ahimaaz and Jonathan?" The woman answered them, "They crossed over the brook." The men searched but found no one, so they returned to Jerusalem.
2SAM|17|21|After the men had gone, the two climbed out of the well and went to inform King David. They said to him, "Set out and cross the river at once; Ahithophel has advised such and such against you."
2SAM|17|22|So David and all the people with him set out and crossed the Jordan. By daybreak, no one was left who had not crossed the Jordan.
2SAM|17|23|When Ahithophel saw that his advice had not been followed, he saddled his donkey and set out for his house in his hometown. He put his house in order and then hanged himself. So he died and was buried in his father's tomb.
2SAM|17|24|David went to Mahanaim, and Absalom crossed the Jordan with all the men of Israel.
2SAM|17|25|Absalom had appointed Amasa over the army in place of Joab. Amasa was the son of a man named Jether, an Israelite who had married Abigail, the daughter of Nahash and sister of Zeruiah the mother of Joab.
2SAM|17|26|The Israelites and Absalom camped in the land of Gilead.
2SAM|17|27|When David came to Mahanaim, Shobi son of Nahash from Rabbah of the Ammonites, and Makir son of Ammiel from Lo Debar, and Barzillai the Gileadite from Rogelim
2SAM|17|28|brought bedding and bowls and articles of pottery. They also brought wheat and barley, flour and roasted grain, beans and lentils,
2SAM|17|29|honey and curds, sheep, and cheese from cows' milk for David and his people to eat. For they said, "The people have become hungry and tired and thirsty in the desert."
2SAM|18|1|David mustered the men who were with him and appointed over them commanders of thousands and commanders of hundreds.
2SAM|18|2|David sent the troops out-a third under the command of Joab, a third under Joab's brother Abishai son of Zeruiah, and a third under Ittai the Gittite. The king told the troops, "I myself will surely march out with you."
2SAM|18|3|But the men said, "You must not go out; if we are forced to flee, they won't care about us. Even if half of us die, they won't care; but you are worth ten thousand of us. It would be better now for you to give us support from the city."
2SAM|18|4|The king answered, "I will do whatever seems best to you." So the king stood beside the gate while all the men marched out in units of hundreds and of thousands.
2SAM|18|5|The king commanded Joab, Abishai and Ittai, "Be gentle with the young man Absalom for my sake." And all the troops heard the king giving orders concerning Absalom to each of the commanders.
2SAM|18|6|The army marched into the field to fight Israel, and the battle took place in the forest of Ephraim.
2SAM|18|7|There the army of Israel was defeated by David's men, and the casualties that day were great-twenty thousand men.
2SAM|18|8|The battle spread out over the whole countryside, and the forest claimed more lives that day than the sword.
2SAM|18|9|Now Absalom happened to meet David's men. He was riding his mule, and as the mule went under the thick branches of a large oak, Absalom's head got caught in the tree. He was left hanging in midair, while the mule he was riding kept on going.
2SAM|18|10|When one of the men saw this, he told Joab, "I just saw Absalom hanging in an oak tree."
2SAM|18|11|Joab said to the man who had told him this, "What! You saw him? Why didn't you strike him to the ground right there? Then I would have had to give you ten shekels of silver and a warrior's belt."
2SAM|18|12|But the man replied, "Even if a thousand shekels were weighed out into my hands, I would not lift my hand against the king's son. In our hearing the king commanded you and Abishai and Ittai, 'Protect the young man Absalom for my sake. '
2SAM|18|13|And if I had put my life in jeopardy -and nothing is hidden from the king-you would have kept your distance from me."
2SAM|18|14|Joab said, "I'm not going to wait like this for you." So he took three javelins in his hand and plunged them into Absalom's heart while Absalom was still alive in the oak tree.
2SAM|18|15|And ten of Joab's armor-bearers surrounded Absalom, struck him and killed him.
2SAM|18|16|Then Joab sounded the trumpet, and the troops stopped pursuing Israel, for Joab halted them.
2SAM|18|17|They took Absalom, threw him into a big pit in the forest and piled up a large heap of rocks over him. Meanwhile, all the Israelites fled to their homes.
2SAM|18|18|During his lifetime Absalom had taken a pillar and erected it in the King's Valley as a monument to himself, for he thought, "I have no son to carry on the memory of my name." He named the pillar after himself, and it is called Absalom's Monument to this day.
2SAM|18|19|Now Ahimaaz son of Zadok said, "Let me run and take the news to the king that the LORD has delivered him from the hand of his enemies."
2SAM|18|20|"You are not the one to take the news today," Joab told him. "You may take the news another time, but you must not do so today, because the king's son is dead."
2SAM|18|21|Then Joab said to a Cushite, "Go, tell the king what you have seen." The Cushite bowed down before Joab and ran off.
2SAM|18|22|Ahimaaz son of Zadok again said to Joab, "Come what may, please let me run behind the Cushite." But Joab replied, "My son, why do you want to go? You don't have any news that will bring you a reward."
2SAM|18|23|He said, "Come what may, I want to run." So Joab said, "Run!" Then Ahimaaz ran by way of the plain and outran the Cushite.
2SAM|18|24|While David was sitting between the inner and outer gates, the watchman went up to the roof of the gateway by the wall. As he looked out, he saw a man running alone.
2SAM|18|25|The watchman called out to the king and reported it. The king said, "If he is alone, he must have good news." And the man came closer and closer.
2SAM|18|26|Then the watchman saw another man running, and he called down to the gatekeeper, "Look, another man running alone!" The king said, "He must be bringing good news, too."
2SAM|18|27|The watchman said, "It seems to me that the first one runs like Ahimaaz son of Zadok.He's a good man," the king said. "He comes with good news."
2SAM|18|28|Then Ahimaaz called out to the king, "All is well!" He bowed down before the king with his face to the ground and said, "Praise be to the LORD your God! He has delivered up the men who lifted their hands against my lord the king."
2SAM|18|29|The king asked, "Is the young man Absalom safe?" Ahimaaz answered, "I saw great confusion just as Joab was about to send the king's servant and me, your servant, but I don't know what it was."
2SAM|18|30|The king said, "Stand aside and wait here." So he stepped aside and stood there.
2SAM|18|31|Then the Cushite arrived and said, "My lord the king, hear the good news! The LORD has delivered you today from all who rose up against you."
2SAM|18|32|The king asked the Cushite, "Is the young man Absalom safe?" The Cushite replied, "May the enemies of my lord the king and all who rise up to harm you be like that young man."
2SAM|18|33|The king was shaken. He went up to the room over the gateway and wept. As he went, he said: "O my son Absalom! My son, my son Absalom! If only I had died instead of you-O Absalom, my son, my son!"
2SAM|19|1|Joab was told, "The king is weeping and mourning for Absalom."
2SAM|19|2|And for the whole army the victory that day was turned into mourning, because on that day the troops heard it said, "The king is grieving for his son."
2SAM|19|3|The men stole into the city that day as men steal in who are ashamed when they flee from battle.
2SAM|19|4|The king covered his face and cried aloud, "O my son Absalom! O Absalom, my son, my son!"
2SAM|19|5|Then Joab went into the house to the king and said, "Today you have humiliated all your men, who have just saved your life and the lives of your sons and daughters and the lives of your wives and concubines.
2SAM|19|6|You love those who hate you and hate those who love you. You have made it clear today that the commanders and their men mean nothing to you. I see that you would be pleased if Absalom were alive today and all of us were dead.
2SAM|19|7|Now go out and encourage your men. I swear by the LORD that if you don't go out, not a man will be left with you by nightfall. This will be worse for you than all the calamities that have come upon you from your youth till now."
2SAM|19|8|So the king got up and took his seat in the gateway. When the men were told, "The king is sitting in the gateway," they all came before him. Meanwhile, the Israelites had fled to their homes.
2SAM|19|9|Throughout the tribes of Israel, the people were all arguing with each other, saying, "The king delivered us from the hand of our enemies; he is the one who rescued us from the hand of the Philistines. But now he has fled the country because of Absalom;
2SAM|19|10|and Absalom, whom we anointed to rule over us, has died in battle. So why do you say nothing about bringing the king back?"
2SAM|19|11|King David sent this message to Zadok and Abiathar, the priests: "Ask the elders of Judah, 'Why should you be the last to bring the king back to his palace, since what is being said throughout Israel has reached the king at his quarters?
2SAM|19|12|You are my brothers, my own flesh and blood. So why should you be the last to bring back the king?'
2SAM|19|13|And say to Amasa, 'Are you not my own flesh and blood? May God deal with me, be it ever so severely, if from now on you are not the commander of my army in place of Joab.'"
2SAM|19|14|He won over the hearts of all the men of Judah as though they were one man. They sent word to the king, "Return, you and all your men."
2SAM|19|15|Then the king returned and went as far as the Jordan. Now the men of Judah had come to Gilgal to go out and meet the king and bring him across the Jordan.
2SAM|19|16|Shimei son of Gera, the Benjamite from Bahurim, hurried down with the men of Judah to meet King David.
2SAM|19|17|With him were a thousand Benjamites, along with Ziba, the steward of Saul's household, and his fifteen sons and twenty servants. They rushed to the Jordan, where the king was.
2SAM|19|18|They crossed at the ford to take the king's household over and to do whatever he wished. When Shimei son of Gera crossed the Jordan, he fell prostrate before the king
2SAM|19|19|and said to him, "May my lord not hold me guilty. Do not remember how your servant did wrong on the day my lord the king left Jerusalem. May the king put it out of his mind.
2SAM|19|20|For I your servant know that I have sinned, but today I have come here as the first of the whole house of Joseph to come down and meet my lord the king."
2SAM|19|21|Then Abishai son of Zeruiah said, "Shouldn't Shimei be put to death for this? He cursed the LORD's anointed."
2SAM|19|22|David replied, "What do you and I have in common, you sons of Zeruiah? This day you have become my adversaries! Should anyone be put to death in Israel today? Do I not know that today I am king over Israel?"
2SAM|19|23|So the king said to Shimei, "You shall not die." And the king promised him on oath.
2SAM|19|24|Mephibosheth, Saul's grandson, also went down to meet the king. He had not taken care of his feet or trimmed his mustache or washed his clothes from the day the king left until the day he returned safely.
2SAM|19|25|When he came from Jerusalem to meet the king, the king asked him, "Why didn't you go with me, Mephibosheth?"
2SAM|19|26|He said, "My lord the king, since I your servant am lame, I said, 'I will have my donkey saddled and will ride on it, so I can go with the king.' But Ziba my servant betrayed me.
2SAM|19|27|And he has slandered your servant to my lord the king. My lord the king is like an angel of God; so do whatever pleases you.
2SAM|19|28|All my grandfather's descendants deserved nothing but death from my lord the king, but you gave your servant a place among those who eat at your table. So what right do I have to make any more appeals to the king?"
2SAM|19|29|The king said to him, "Why say more? I order you and Ziba to divide the fields."
2SAM|19|30|Mephibosheth said to the king, "Let him take everything, now that my lord the king has arrived home safely."
2SAM|19|31|Barzillai the Gileadite also came down from Rogelim to cross the Jordan with the king and to send him on his way from there.
2SAM|19|32|Now Barzillai was a very old man, eighty years of age. He had provided for the king during his stay in Mahanaim, for he was a very wealthy man.
2SAM|19|33|The king said to Barzillai, "Cross over with me and stay with me in Jerusalem, and I will provide for you."
2SAM|19|34|But Barzillai answered the king, "How many more years will I live, that I should go up to Jerusalem with the king?
2SAM|19|35|I am now eighty years old. Can I tell the difference between what is good and what is not? Can your servant taste what he eats and drinks? Can I still hear the voices of men and women singers? Why should your servant be an added burden to my lord the king?
2SAM|19|36|Your servant will cross over the Jordan with the king for a short distance, but why should the king reward me in this way?
2SAM|19|37|Let your servant return, that I may die in my own town near the tomb of my father and mother. But here is your servant Kimham. Let him cross over with my lord the king. Do for him whatever pleases you."
2SAM|19|38|The king said, "Kimham shall cross over with me, and I will do for him whatever pleases you. And anything you desire from me I will do for you."
2SAM|19|39|So all the people crossed the Jordan, and then the king crossed over. The king kissed Barzillai and gave him his blessing, and Barzillai returned to his home.
2SAM|19|40|When the king crossed over to Gilgal, Kimham crossed with him. All the troops of Judah and half the troops of Israel had taken the king over.
2SAM|19|41|Soon all the men of Israel were coming to the king and saying to him, "Why did our brothers, the men of Judah, steal the king away and bring him and his household across the Jordan, together with all his men?"
2SAM|19|42|All the men of Judah answered the men of Israel, "We did this because the king is closely related to us. Why are you angry about it? Have we eaten any of the king's provisions? Have we taken anything for ourselves?"
2SAM|19|43|Then the men of Israel answered the men of Judah, "We have ten shares in the king; and besides, we have a greater claim on David than you have. So why do you treat us with contempt? Were we not the first to speak of bringing back our king?" But the men of Judah responded even more harshly than the men of Israel.
2SAM|20|1|Now a troublemaker named Sheba son of Bicri, a Benjamite, happened to be there. He sounded the trumpet and shouted, "We have no share in David, no part in Jesse's son! Every man to his tent, O Israel!"
2SAM|20|2|So all the men of Israel deserted David to follow Sheba son of Bicri. But the men of Judah stayed by their king all the way from the Jordan to Jerusalem.
2SAM|20|3|When David returned to his palace in Jerusalem, he took the ten concubines he had left to take care of the palace and put them in a house under guard. He provided for them, but did not lie with them. They were kept in confinement till the day of their death, living as widows.
2SAM|20|4|Then the king said to Amasa, "Summon the men of Judah to come to me within three days, and be here yourself."
2SAM|20|5|But when Amasa went to summon Judah, he took longer than the time the king had set for him.
2SAM|20|6|David said to Abishai, "Now Sheba son of Bicri will do us more harm than Absalom did. Take your master's men and pursue him, or he will find fortified cities and escape from us."
2SAM|20|7|So Joab's men and the Kerethites and Pelethites and all the mighty warriors went out under the command of Abishai. They marched out from Jerusalem to pursue Sheba son of Bicri.
2SAM|20|8|While they were at the great rock in Gibeon, Amasa came to meet them. Joab was wearing his military tunic, and strapped over it at his waist was a belt with a dagger in its sheath. As he stepped forward, it dropped out of its sheath.
2SAM|20|9|Joab said to Amasa, "How are you, my brother?" Then Joab took Amasa by the beard with his right hand to kiss him.
2SAM|20|10|Amasa was not on his guard against the dagger in Joab's hand, and Joab plunged it into his belly, and his intestines spilled out on the ground. Without being stabbed again, Amasa died. Then Joab and his brother Abishai pursued Sheba son of Bicri.
2SAM|20|11|One of Joab's men stood beside Amasa and said, "Whoever favors Joab, and whoever is for David, let him follow Joab!"
2SAM|20|12|Amasa lay wallowing in his blood in the middle of the road, and the man saw that all the troops came to a halt there. When he realized that everyone who came up to Amasa stopped, he dragged him from the road into a field and threw a garment over him.
2SAM|20|13|After Amasa had been removed from the road, all the men went on with Joab to pursue Sheba son of Bicri.
2SAM|20|14|Sheba passed through all the tribes of Israel to Abel Beth Maacah and through the entire region of the Berites, who gathered together and followed him.
2SAM|20|15|All the troops with Joab came and besieged Sheba in Abel Beth Maacah. They built a siege ramp up to the city, and it stood against the outer fortifications. While they were battering the wall to bring it down,
2SAM|20|16|a wise woman called from the city, "Listen! Listen! Tell Joab to come here so I can speak to him."
2SAM|20|17|He went toward her, and she asked, "Are you Joab?I am," he answered. She said, "Listen to what your servant has to say.I'm listening," he said.
2SAM|20|18|She continued, "Long ago they used to say, 'Get your answer at Abel,' and that settled it.
2SAM|20|19|We are the peaceful and faithful in Israel. You are trying to destroy a city that is a mother in Israel. Why do you want to swallow up the LORD's inheritance?"
2SAM|20|20|"Far be it from me!" Joab replied, "Far be it from me to swallow up or destroy!
2SAM|20|21|That is not the case. A man named Sheba son of Bicri, from the hill country of Ephraim, has lifted up his hand against the king, against David. Hand over this one man, and I'll withdraw from the city." The woman said to Joab, "His head will be thrown to you from the wall."
2SAM|20|22|Then the woman went to all the people with her wise advice, and they cut off the head of Sheba son of Bicri and threw it to Joab. So he sounded the trumpet, and his men dispersed from the city, each returning to his home. And Joab went back to the king in Jerusalem.
2SAM|20|23|Joab was over Israel's entire army; Benaiah son of Jehoiada was over the Kerethites and Pelethites;
2SAM|20|24|Adoniram was in charge of forced labor; Jehoshaphat son of Ahilud was recorder;
2SAM|20|25|Sheva was secretary; Zadok and Abiathar were priests;
2SAM|20|26|and Ira the Jairite was David's priest.
2SAM|21|1|During the reign of David, there was a famine for three successive years; so David sought the face of the LORD. The LORD said, "It is on account of Saul and his blood-stained house; it is because he put the Gibeonites to death."
2SAM|21|2|The king summoned the Gibeonites and spoke to them. (Now the Gibeonites were not a part of Israel but were survivors of the Amorites; the Israelites had sworn to spare them, but Saul in his zeal for Israel and Judah had tried to annihilate them.)
2SAM|21|3|David asked the Gibeonites, "What shall I do for you? How shall I make amends so that you will bless the LORD's inheritance?"
2SAM|21|4|The Gibeonites answered him, "We have no right to demand silver or gold from Saul or his family, nor do we have the right to put anyone in Israel to death.What do you want me to do for you?" David asked.
2SAM|21|5|They answered the king, "As for the man who destroyed us and plotted against us so that we have been decimated and have no place anywhere in Israel,
2SAM|21|6|let seven of his male descendants be given to us to be killed and exposed before the LORD at Gibeah of Saul-the Lord 's chosen one." So the king said, "I will give them to you."
2SAM|21|7|The king spared Mephibosheth son of Jonathan, the son of Saul, because of the oath before the LORD between David and Jonathan son of Saul.
2SAM|21|8|But the king took Armoni and Mephibosheth, the two sons of Aiah's daughter Rizpah, whom she had borne to Saul, together with the five sons of Saul's daughter Merab, whom she had borne to Adriel son of Barzillai the Meholathite.
2SAM|21|9|He handed them over to the Gibeonites, who killed and exposed them on a hill before the LORD. All seven of them fell together; they were put to death during the first days of the harvest, just as the barley harvest was beginning.
2SAM|21|10|Rizpah daughter of Aiah took sackcloth and spread it out for herself on a rock. From the beginning of the harvest till the rain poured down from the heavens on the bodies, she did not let the birds of the air touch them by day or the wild animals by night.
2SAM|21|11|When David was told what Aiah's daughter Rizpah, Saul's concubine, had done,
2SAM|21|12|he went and took the bones of Saul and his son Jonathan from the citizens of Jabesh Gilead. (They had taken them secretly from the public square at Beth Shan, where the Philistines had hung them after they struck Saul down on Gilboa.)
2SAM|21|13|David brought the bones of Saul and his son Jonathan from there, and the bones of those who had been killed and exposed were gathered up.
2SAM|21|14|They buried the bones of Saul and his son Jonathan in the tomb of Saul's father Kish, at Zela in Benjamin, and did everything the king commanded. After that, God answered prayer in behalf of the land.
2SAM|21|15|Once again there was a battle between the Philistines and Israel. David went down with his men to fight against the Philistines, and he became exhausted.
2SAM|21|16|And Ishbi-Benob, one of the descendants of Rapha, whose bronze spearhead weighed three hundred shekels and who was armed with a new sword, said he would kill David.
2SAM|21|17|But Abishai son of Zeruiah came to David's rescue; he struck the Philistine down and killed him. Then David's men swore to him, saying, "Never again will you go out with us to battle, so that the lamp of Israel will not be extinguished."
2SAM|21|18|In the course of time, there was another battle with the Philistines, at Gob. At that time Sibbecai the Hushathite killed Saph, one of the descendants of Rapha.
2SAM|21|19|In another battle with the Philistines at Gob, Elhanan son of Jaare-Oregim the Bethlehemite killed Goliath the Gittite, who had a spear with a shaft like a weaver's rod.
2SAM|21|20|In still another battle, which took place at Gath, there was a huge man with six fingers on each hand and six toes on each foot-twenty-four in all. He also was descended from Rapha.
2SAM|21|21|When he taunted Israel, Jonathan son of Shimeah, David's brother, killed him.
2SAM|21|22|These four were descendants of Rapha in Gath, and they fell at the hands of David and his men.
2SAM|22|1|David sang to the LORD the words of this song when the LORD delivered him from the hand of all his enemies and from the hand of Saul.
2SAM|22|2|He said: "The LORD is my rock, my fortress and my deliverer;
2SAM|22|3|my God is my rock, in whom I take refuge, my shield and the horn of my salvation. He is my stronghold, my refuge and my savior- from violent men you save me.
2SAM|22|4|I call to the LORD, who is worthy of praise, and I am saved from my enemies.
2SAM|22|5|"The waves of death swirled about me; the torrents of destruction overwhelmed me.
2SAM|22|6|The cords of the grave coiled around me; the snares of death confronted me.
2SAM|22|7|In my distress I called to the LORD; I called out to my God. From his temple he heard my voice; my cry came to his ears.
2SAM|22|8|"The earth trembled and quaked, the foundations of the heavens shook; they trembled because he was angry.
2SAM|22|9|Smoke rose from his nostrils; consuming fire came from his mouth, burning coals blazed out of it.
2SAM|22|10|He parted the heavens and came down; dark clouds were under his feet.
2SAM|22|11|He mounted the cherubim and flew; he soared on the wings of the wind.
2SAM|22|12|He made darkness his canopy around him- the dark rain clouds of the sky.
2SAM|22|13|Out of the brightness of his presence bolts of lightning blazed forth.
2SAM|22|14|The LORD thundered from heaven; the voice of the Most High resounded.
2SAM|22|15|He shot arrows and scattered the enemies, bolts of lightning and routed them.
2SAM|22|16|The valleys of the sea were exposed and the foundations of the earth laid bare at the rebuke of the LORD, at the blast of breath from his nostrils.
2SAM|22|17|"He reached down from on high and took hold of me; he drew me out of deep waters.
2SAM|22|18|He rescued me from my powerful enemy, from my foes, who were too strong for me.
2SAM|22|19|They confronted me in the day of my disaster, but the LORD was my support.
2SAM|22|20|He brought me out into a spacious place; he rescued me because he delighted in me.
2SAM|22|21|"The LORD has dealt with me according to my righteousness; according to the cleanness of my hands he has rewarded me.
2SAM|22|22|For I have kept the ways of the LORD; I have not done evil by turning from my God.
2SAM|22|23|All his laws are before me; I have not turned away from his decrees.
2SAM|22|24|I have been blameless before him and have kept myself from sin.
2SAM|22|25|The LORD has rewarded me according to my righteousness, according to my cleanness in his sight.
2SAM|22|26|"To the faithful you show yourself faithful, to the blameless you show yourself blameless,
2SAM|22|27|to the pure you show yourself pure, but to the crooked you show yourself shrewd.
2SAM|22|28|You save the humble, but your eyes are on the haughty to bring them low.
2SAM|22|29|You are my lamp, O LORD; the LORD turns my darkness into light.
2SAM|22|30|With your help I can advance against a troop; with my God I can scale a wall.
2SAM|22|31|"As for God, his way is perfect; the word of the LORD is flawless. He is a shield for all who take refuge in him.
2SAM|22|32|For who is God besides the LORD? And who is the Rock except our God?
2SAM|22|33|It is God who arms me with strength and makes my way perfect.
2SAM|22|34|He makes my feet like the feet of a deer; he enables me to stand on the heights.
2SAM|22|35|He trains my hands for battle; my arms can bend a bow of bronze.
2SAM|22|36|You give me your shield of victory; you stoop down to make me great.
2SAM|22|37|You broaden the path beneath me, so that my ankles do not turn.
2SAM|22|38|"I pursued my enemies and crushed them; I did not turn back till they were destroyed.
2SAM|22|39|I crushed them completely, and they could not rise; they fell beneath my feet.
2SAM|22|40|You armed me with strength for battle; you made my adversaries bow at my feet.
2SAM|22|41|You made my enemies turn their backs in flight, and I destroyed my foes.
2SAM|22|42|They cried for help, but there was no one to save them- to the LORD, but he did not answer.
2SAM|22|43|I beat them as fine as the dust of the earth; I pounded and trampled them like mud in the streets.
2SAM|22|44|"You have delivered me from the attacks of my people; you have preserved me as the head of nations. People I did not know are subject to me,
2SAM|22|45|and foreigners come cringing to me; as soon as they hear me, they obey me.
2SAM|22|46|They all lose heart; they come trembling from their strongholds.
2SAM|22|47|"The LORD lives! Praise be to my Rock! Exalted be God, the Rock, my Savior!
2SAM|22|48|He is the God who avenges me, who puts the nations under me,
2SAM|22|49|who sets me free from my enemies. You exalted me above my foes; from violent men you rescued me.
2SAM|22|50|Therefore I will praise you, O LORD, among the nations; I will sing praises to your name.
2SAM|22|51|He gives his king great victories; he shows unfailing kindness to his anointed, to David and his descendants forever."
2SAM|23|1|These are the last words of David: "The oracle of David son of Jesse, the oracle of the man exalted by the Most High, the man anointed by the God of Jacob, Israel's singer of songs:
2SAM|23|2|"The Spirit of the LORD spoke through me; his word was on my tongue.
2SAM|23|3|The God of Israel spoke, the Rock of Israel said to me: 'When one rules over men in righteousness, when he rules in the fear of God,
2SAM|23|4|he is like the light of morning at sunrise on a cloudless morning, like the brightness after rain that brings the grass from the earth.'
2SAM|23|5|"Is not my house right with God? Has he not made with me an everlasting covenant, arranged and secured in every part? Will he not bring to fruition my salvation and grant me my every desire?
2SAM|23|6|But evil men are all to be cast aside like thorns, which are not gathered with the hand.
2SAM|23|7|Whoever touches thorns uses a tool of iron or the shaft of a spear; they are burned up where they lie."
2SAM|23|8|These are the names of David's mighty men: Josheb-Basshebeth, a Tahkemonite, was chief of the Three; he raised his spear against eight hundred men, whom he killed in one encounter.
2SAM|23|9|Next to him was Eleazar son of Dodai the Ahohite. As one of the three mighty men, he was with David when they taunted the Philistines gathered at Pas Dammim for battle. Then the men of Israel retreated,
2SAM|23|10|but he stood his ground and struck down the Philistines till his hand grew tired and froze to the sword. The LORD brought about a great victory that day. The troops returned to Eleazar, but only to strip the dead.
2SAM|23|11|Next to him was Shammah son of Agee the Hararite. When the Philistines banded together at a place where there was a field full of lentils, Israel's troops fled from them.
2SAM|23|12|But Shammah took his stand in the middle of the field. He defended it and struck the Philistines down, and the LORD brought about a great victory.
2SAM|23|13|During harvest time, three of the thirty chief men came down to David at the cave of Adullam, while a band of Philistines was encamped in the Valley of Rephaim.
2SAM|23|14|At that time David was in the stronghold, and the Philistine garrison was at Bethlehem.
2SAM|23|15|David longed for water and said, "Oh, that someone would get me a drink of water from the well near the gate of Bethlehem!"
2SAM|23|16|So the three mighty men broke through the Philistine lines, drew water from the well near the gate of Bethlehem and carried it back to David. But he refused to drink it; instead, he poured it out before the LORD.
2SAM|23|17|"Far be it from me, O LORD, to do this!" he said. "Is it not the blood of men who went at the risk of their lives?" And David would not drink it. Such were the exploits of the three mighty men.
2SAM|23|18|Abishai the brother of Joab son of Zeruiah was chief of the Three. He raised his spear against three hundred men, whom he killed, and so he became as famous as the Three.
2SAM|23|19|Was he not held in greater honor than the Three? He became their commander, even though he was not included among them.
2SAM|23|20|Benaiah son of Jehoiada was a valiant fighter from Kabzeel, who performed great exploits. He struck down two of Moab's best men. He also went down into a pit on a snowy day and killed a lion.
2SAM|23|21|And he struck down a huge Egyptian. Although the Egyptian had a spear in his hand, Benaiah went against him with a club. He snatched the spear from the Egyptian's hand and killed him with his own spear.
2SAM|23|22|Such were the exploits of Benaiah son of Jehoiada; he too was as famous as the three mighty men.
2SAM|23|23|He was held in greater honor than any of the Thirty, but he was not included among the Three. And David put him in charge of his bodyguard.
2SAM|23|24|Among the Thirty were: Asahel the brother of Joab, Elhanan son of Dodo from Bethlehem,
2SAM|23|25|Shammah the Harodite, Elika the Harodite,
2SAM|23|26|Helez the Paltite, Ira son of Ikkesh from Tekoa,
2SAM|23|27|Abiezer from Anathoth, Mebunnai the Hushathite,
2SAM|23|28|Zalmon the Ahohite, Maharai the Netophathite,
2SAM|23|29|Heled son of Baanah the Netophathite, Ithai son of Ribai from Gibeah in Benjamin,
2SAM|23|30|Benaiah the Pirathonite, Hiddai from the ravines of Gaash,
2SAM|23|31|Abi-Albon the Arbathite, Azmaveth the Barhumite,
2SAM|23|32|Eliahba the Shaalbonite, the sons of Jashen, Jonathan
2SAM|23|33|son of Shammah the Hararite, Ahiam son of Sharar the Hararite,
2SAM|23|34|Eliphelet son of Ahasbai the Maacathite, Eliam son of Ahithophel the Gilonite,
2SAM|23|35|Hezro the Carmelite, Paarai the Arbite,
2SAM|23|36|Igal son of Nathan from Zobah, the son of Hagri,
2SAM|23|37|Zelek the Ammonite, Naharai the Beerothite, the armor-bearer of Joab son of Zeruiah,
2SAM|23|38|Ira the Ithrite, Gareb the Ithrite
2SAM|23|39|and Uriah the Hittite. There were thirty-seven in all.
2SAM|24|1|Again the anger of the LORD burned against Israel, and he incited David against them, saying, "Go and take a census of Israel and Judah."
2SAM|24|2|So the king said to Joab and the army commanders with him, "Go throughout the tribes of Israel from Dan to Beersheba and enroll the fighting men, so that I may know how many there are."
2SAM|24|3|But Joab replied to the king, "May the LORD your God multiply the troops a hundred times over, and may the eyes of my lord the king see it. But why does my lord the king want to do such a thing?"
2SAM|24|4|The king's word, however, overruled Joab and the army commanders; so they left the presence of the king to enroll the fighting men of Israel.
2SAM|24|5|After crossing the Jordan, they camped near Aroer, south of the town in the gorge, and then went through Gad and on to Jazer.
2SAM|24|6|They went to Gilead and the region of Tahtim Hodshi, and on to Dan Jaan and around toward Sidon.
2SAM|24|7|Then they went toward the fortress of Tyre and all the towns of the Hivites and Canaanites. Finally, they went on to Beersheba in the Negev of Judah.
2SAM|24|8|After they had gone through the entire land, they came back to Jerusalem at the end of nine months and twenty days.
2SAM|24|9|Joab reported the number of the fighting men to the king: In Israel there were eight hundred thousand able-bodied men who could handle a sword, and in Judah five hundred thousand.
2SAM|24|10|David was conscience-stricken after he had counted the fighting men, and he said to the LORD, "I have sinned greatly in what I have done. Now, O LORD, I beg you, take away the guilt of your servant. I have done a very foolish thing."
2SAM|24|11|Before David got up the next morning, the word of the LORD had come to Gad the prophet, David's seer:
2SAM|24|12|"Go and tell David, 'This is what the LORD says: I am giving you three options. Choose one of them for me to carry out against you.'"
2SAM|24|13|So Gad went to David and said to him, "Shall there come upon you three years of famine in your land? Or three months of fleeing from your enemies while they pursue you? Or three days of plague in your land? Now then, think it over and decide how I should answer the one who sent me."
2SAM|24|14|David said to Gad, "I am in deep distress. Let us fall into the hands of the LORD, for his mercy is great; but do not let me fall into the hands of men."
2SAM|24|15|So the LORD sent a plague on Israel from that morning until the end of the time designated, and seventy thousand of the people from Dan to Beersheba died.
2SAM|24|16|When the angel stretched out his hand to destroy Jerusalem, the LORD was grieved because of the calamity and said to the angel who was afflicting the people, "Enough! Withdraw your hand." The angel of the LORD was then at the threshing floor of Araunah the Jebusite.
2SAM|24|17|When David saw the angel who was striking down the people, he said to the LORD, "I am the one who has sinned and done wrong. These are but sheep. What have they done? Let your hand fall upon me and my family."
2SAM|24|18|On that day Gad went to David and said to him, "Go up and build an altar to the LORD on the threshing floor of Araunah the Jebusite."
2SAM|24|19|So David went up, as the LORD had commanded through Gad.
2SAM|24|20|When Araunah looked and saw the king and his men coming toward him, he went out and bowed down before the king with his face to the ground.
2SAM|24|21|Araunah said, "Why has my lord the king come to his servant?To buy your threshing floor," David answered, "so I can build an altar to the LORD, that the plague on the people may be stopped."
2SAM|24|22|Araunah said to David, "Let my lord the king take whatever pleases him and offer it up. Here are oxen for the burnt offering, and here are threshing sledges and ox yokes for the wood.
2SAM|24|23|O king, Araunah gives all this to the king." Araunah also said to him, "May the LORD your God accept you."
2SAM|24|24|But the king replied to Araunah, "No, I insist on paying you for it. I will not sacrifice to the LORD my God burnt offerings that cost me nothing." So David bought the threshing floor and the oxen and paid fifty shekels of silver for them.
2SAM|24|25|David built an altar to the LORD there and sacrificed burnt offerings and fellowship offerings. Then the LORD answered prayer in behalf of the land, and the plague on Israel was stopped.
