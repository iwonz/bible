ESTH|1|1|И было во дни Артаксеркса, – этот Артаксеркс царствовал над ста двадцатью семью областями от Индии и до Ефиопии, –
ESTH|1|2|в то время, как царь Артаксеркс сел на царский престол свой, что в Сузах, городе престольном,
ESTH|1|3|в третий год своего царствования он сделал пир для всех князей своих и для служащих при нем, для главных начальников войска Персидского и Мидийского и для правителей областей своих,
ESTH|1|4|показывая великое богатство царства своего и отличный блеск величия своего [в течение] многих дней, ста восьмидесяти дней.
ESTH|1|5|По окончании сих дней, сделал царь для народа своего, находившегося в престольном городе Сузах, от большого до малого, пир семидневный на садовом дворе дома царского.
ESTH|1|6|Белые, бумажные и яхонтового цвета шерстяные ткани, прикрепленные виссонными и пурпуровыми шнурами, [висели] на серебряных кольцах и мраморных столбах.
ESTH|1|7|Золотые и серебряные ложа [были] на помосте, устланном камнями зеленого цвета и мрамором, и перламутром, и камнями черного цвета.
ESTH|1|8|Напитки подаваемы [были] в золотых сосудах и сосудах разнообразных, ценою в тридцать тысяч талантов; и вина царского было множество, по богатству царя. Питье [шло] чинно, никто не принуждал, потому что царь дал такое приказание всем управляющим в доме его, чтобы делали по воле каждого.
ESTH|1|9|И царица Астинь сделала также пир для женщин в царском доме царя Артаксеркса.
ESTH|1|10|В седьмой день, когда развеселилось сердце царя от вина, он сказал Мегуману, Бизфе, Харбоне, Бигфе и Авагфе, Зефару и Каркасу – семи евнухам, служившим пред лицем царя Артаксеркса,
ESTH|1|11|чтобы они привели царицу Астинь пред лице царя в венце царском для того, чтобы показать народам и князьям красоту ее; потому что она была очень красива.
ESTH|1|12|Но царица Астинь не захотела прийти по приказанию царя, [объявленному] чрез евнухов.
ESTH|1|13|И разгневался царь сильно, и ярость его загорелась в нем. И сказал царь мудрецам, знающим [прежние] времена – ибо дела царя [делались] пред всеми знающими закон и права, –
ESTH|1|14|приближенными же к нему [тогда были]: Каршена, Шефар, Адмафа, Фарсис, Мерес, Марсена, Мемухан – семь князей Персидских и Мидийских, которые могли видеть лице царя [и] сидели первыми в царстве:
ESTH|1|15|как поступить по закону с царицею Астинь за то, что она не сделала по слову царя Артаксеркса, [объявленному] чрез евнухов?
ESTH|1|16|И сказал Мемухан пред лицем царя и князей: не пред царем одним виновна царица Астинь, а пред всеми князьями и пред всеми народами, которые по всем областям царя Артаксеркса;
ESTH|1|17|потому что поступок царицы дойдет до всех жен, и они будут пренебрегать мужьями своими и говорить: царь Артаксеркс велел привести царицу Астинь пред лице свое, а она не пошла.
ESTH|1|18|Теперь княгини Персидские и Мидийские, которые услышат о поступке царицы, будут [то же] говорить всем князьям царя; и пренебрежения и огорчения будет довольно.
ESTH|1|19|Если благоугодно царю, пусть выйдет от него царское постановление и впишется в законы Персидские и Мидийские и не отменяется, о том, что Астинь не будет входить пред лице царя Артаксеркса, а царское достоинство ее царь передаст другой, которая лучше ее.
ESTH|1|20|Когда услышат о сем постановлении царя, которое разойдется по всему царству его, как оно ни велико, тогда все жены будут почитать мужей своих, от большого до малого.
ESTH|1|21|И угодно было слово сие в глазах царя и князей; и сделал царь по слову Мемухана.
ESTH|1|22|И послал во все области царя письма, писанные в каждую область письменами ее и к каждому народу на языке его, чтобы всякий муж был господином в доме своем, и чтобы это было объявлено каждому на природном языке его.
ESTH|2|1|После сего, когда утих гнев царя Артаксеркса, он вспомнил об Астинь и о том, что она сделала, и что было определено о ней.
ESTH|2|2|И сказали отроки царя, служившие при нем: пусть бы поискали царю молодых красивых девиц,
ESTH|2|3|и пусть бы назначил царь наблюдателей во все области своего царства, которые собрали бы всех молодых девиц, красивых видом, в престольный город Сузы, в дом жен под надзор Гегая, царского евнуха, стража жен, и пусть бы выдавали им притиранья,
ESTH|2|4|и девица, которая понравится глазам царя, пусть будет царицею вместо Астинь. И угодно было слово это в глазах царя, и он так и сделал.
ESTH|2|5|Был в Сузах, городе престольном, один Иудеянин, имя его Мардохей, сын Иаира, сын Семея, сын Киса, из колена Вениаминова.
ESTH|2|6|Он был переселен из Иерусалима вместе с пленниками, выведенными с Иехониею, царем Иудейским, которых переселил Навуходоносор, царь Вавилонский.
ESTH|2|7|И был он воспитателем Гадассы, – она же Есфирь, – дочери дяди его, так как не было у нее ни отца, ни матери. Девица эта была красива станом и пригожа лицем. И по смерти отца ее и матери ее, Мардохей взял ее к себе вместо дочери.
ESTH|2|8|Когда объявлено было повеление царя и указ его, и когда собраны были многие девицы в престольный город Сузы под надзор Гегая, тогда взята была и Есфирь в царский дом под надзор Гегая, стража жен.
ESTH|2|9|И понравилась эта девица глазам его и приобрела у него благоволение, и он поспешил выдать ей притиранья и [все, назначенное на] часть ее, и приставить к ней семь девиц, достойных быть при ней, из дома царского, и переместил ее и девиц ее в лучшее отделение женского дома.
ESTH|2|10|Не сказывала Есфирь ни о народе своем, ни о родстве своем, потому что Мардохей дал ей приказание, чтобы она не сказывала.
ESTH|2|11|И всякий день Мардохей приходил ко двору женского дома, чтобы наведываться о здоровье Есфири и о том, что делается с нею.
ESTH|2|12|Когда наступало время каждой девице входить к царю Артаксерксу, после того, как в течение двенадцати месяцев выполнено было над нею все, определенное женщинам, – ибо столько времени продолжались дни притиранья их: шесть месяцев мирровым маслом и шесть месяцев ароматами и другими притираньями женскими, –
ESTH|2|13|тогда девица входила к царю. Чего бы она ни потребовала, ей давали все для выхода из женского дома в дом царя.
ESTH|2|14|Вечером она входила и утром возвращалась в другой дом женский под надзор Шаазгаза, царского евнуха, стража наложниц; и уже не входила к царю, разве только царь пожелал бы ее, и она призывалась бы по имени.
ESTH|2|15|Когда настало время Есфири, дочери Аминадава, дяди Мардохея, который взял ее к себе вместо дочери, – идти к царю, тогда она не просила ничего, кроме того, о чем сказал ей Гегай, евнух царский, страж жен. И приобрела Есфирь расположение [к себе] в глазах всех, видевших ее.
ESTH|2|16|И взята была Есфирь к царю Артаксерксу, в царский дом его, в десятом месяце, то есть в месяце Тебефе, в седьмой год его царствования.
ESTH|2|17|И полюбил царь Есфирь более всех жен, и она приобрела его благоволение и благорасположение более всех девиц; и он возложил царский венец на голову ее и сделал ее царицею на место Астинь.
ESTH|2|18|И сделал царь большой пир для всех князей своих и для служащих при нем, – пир ради Есфири, и сделал льготу областям и роздал дары с царственною щедростью.
ESTH|2|19|И когда во второй раз собраны были девицы, и Мардохей сидел у ворот царских,
ESTH|2|20|Есфирь все еще не сказывала о родстве своем и о народе своем, как приказал ей Мардохей; а слово Мардохея Есфирь выполняла [и теперь] так же, как тогда, когда была у него на воспитании.
ESTH|2|21|В это время, как Мардохей сидел у ворот царских, два царских евнуха, Гавафа и Фарра, оберегавшие порог, озлобились, и замышляли наложить руку на царя Артаксеркса.
ESTH|2|22|Узнав о том, Мардохей сообщил царице Есфири, а Есфирь сказала царю от имени Мардохея.
ESTH|2|23|Дело было исследовано и найдено [верным], и их обоих повесили на дереве. И было вписано о благодеянии Мардохея в книгу дневных записей у царя.
ESTH|3|1|После сего возвеличил царь Артаксеркс Амана, сына Амадафа, Вугеянина, и вознес его, и поставил седалище его выше всех князей, которые у него;
ESTH|3|2|и все служащие при царе, которые [были] у царских ворот, кланялись и падали ниц пред Аманом, ибо так приказал царь. А Мардохей не кланялся и не падал ниц.
ESTH|3|3|И говорили служащие при царе, которые у царских ворот, Мардохею: зачем ты преступаешь повеление царское?
ESTH|3|4|И как они говорили ему каждый день, а он не слушал их, то они донесли Аману, чтобы посмотреть, устоит ли в слове [своем] Мардохей, ибо он сообщил им, что он Иудеянин.
ESTH|3|5|И когда увидел Аман, что Мардохей не кланяется и не падает ниц пред ним, то исполнился гнева Аман.
ESTH|3|6|И показалось ему ничтожным наложить руку на одного Мардохея; но так как сказали ему, из какого народа Мардохей, то задумал Аман истребить всех Иудеев, которые [были] во всем царстве Артаксеркса, [как] народ Мардохеев.
ESTH|3|7|в первый месяц, который есть месяц Нисан, в двенадцатый год царя Артаксеркса, и бросали пур, то есть жребий, пред лицем Амана изо дня в день и из месяца в месяц, [и пал жребий] на двенадцатый [месяц], то есть на месяц Адар.
ESTH|3|8|И сказал Аман царю Артаксерксу: есть один народ, разбросанный и рассеянный между народами по всем областям царства твоего; и законы их отличны от [законов] всех народов, и законов царя они не выполняют; и царю не следует [так] оставлять их.
ESTH|3|9|Если царю благоугодно, то пусть будет предписано истребить их, и десять тысяч талантов серебра я отвешу в руки приставников, чтобы внести в казну царскую.
ESTH|3|10|Тогда снял царь перстень свой с руки своей и отдал его Аману, сыну Амадафа, Вугеянину, чтобы скрепить указ против Иудеев.
ESTH|3|11|И сказал царь Аману: отдаю тебе [это] серебро и народ; поступи с ним, как тебе угодно.
ESTH|3|12|И призваны были писцы царские в первый месяц, в тринадцатый день его, и написано было, как приказал Аман, к сатрапам царским и к начальствующим над каждою областью и к князьям у каждого народа, в каждую область письменами ее и к каждому народу на языке его: [все] было написано от имени царя Артаксеркса и скреплено царским перстнем.
ESTH|3|13|И посланы были письма через гонцов во все области царя, чтобы убить, погубить и истребить всех Иудеев, малого и старого, детей и женщин в один день, в тринадцатый день двенадцатого месяца, то есть месяца Адара, и имение их разграбить.
ESTH|3|14|Список с указа отдать в каждую область [как] закон, объявляемый для всех народов, чтобы они были готовы к тому дню.
ESTH|3|15|Гонцы отправились быстро с царским повелением. Объявлен был указ и в Сузах, престольном городе; и царь и Аман сидели и пили, а город Сузы [был] в смятении.
ESTH|4|1|Когда Мардохей узнал все, что делалось, разодрал одежды свои и возложил на себя вретище и пепел, и вышел на средину города и взывал с воплем великим и горьким.
ESTH|4|2|И дошел до царских ворот; так как нельзя было входить в царские ворота во вретище.
ESTH|4|3|Равно и во всякой области и месте, куда [только] доходило повеление царя и указ его, было большое сетование у Иудеев, и пост, и плач, и вопль; вретище и пепел служили постелью для многих.
ESTH|4|4|И пришли служанки Есфири и евнухи ее и рассказали ей, и сильно встревожилась царица. И послала одежды, чтобы Мардохей надел их и снял с себя вретище свое. Но он не принял.
ESTH|4|5|Тогда позвала Есфирь Гафаха, одного из евнухов царя, которого он приставил к ней, и послала его к Мардохею узнать: что это и отчего это?
ESTH|4|6|И пошел Гафах к Мардохею на городскую площадь, которая пред царскими воротами.
ESTH|4|7|И рассказал ему Мардохей обо всем, что с ним случилось, и об определенном числе серебра, которое обещал Аман отвесить в казну царскую за Иудеев, чтобы истребить их;
ESTH|4|8|и вручил ему список с указа, обнародованного в Сузах, об истреблении их, чтобы показать Есфири и дать ей знать [обо всем]; притом наказывал ей, чтобы она пошла к царю и молила его о помиловании и просила его за народ свой.
ESTH|4|9|И пришел Гафах и пересказал Есфири слова Мардохея.
ESTH|4|10|И сказала Есфирь Гафаху и послала его [сказать] Мардохею:
ESTH|4|11|все служащие при царе и народы в областях царских знают, что всякому, и мужчине и женщине, кто войдет к царю во внутренний двор, не быв позван, один суд – смерть; только тот, к кому прострет царь свой золотой скипетр, останется жив. А я не звана к царю вот уже тридцать дней.
ESTH|4|12|И пересказали Мардохею слова Есфири.
ESTH|4|13|И сказал Мардохей в ответ Есфири: не думай, что ты [одна] спасешься в доме царском из всех Иудеев.
ESTH|4|14|Если ты промолчишь в это время, то свобода и избавление придет для Иудеев из другого места, а ты и дом отца твоего погибнете. И кто знает, не для такого ли времени ты и достигла достоинства царского?
ESTH|4|15|И сказала Есфирь в ответ Мардохею:
ESTH|4|16|пойди, собери всех Иудеев, находящихся в Сузах, и поститесь ради меня, и не ешьте и не пейте три дня, ни днем, ни ночью, и я с служанками моими буду также поститься и потом пойду к царю, хотя это против закона, и если погибнуть – погибну.
ESTH|4|17|И пошел Мардохей и сделал, как приказала ему Есфирь.
ESTH|5|1|На третий день Есфирь оделась по–царски, и стала она на внутреннем дворе царского дома, перед домом царя; царь же сидел [тогда] на царском престоле своем, в царском доме, прямо против входа в дом, Когда царь увидел царицу Есфирь, стоящую на дворе, она нашла милость в глазах его.
ESTH|5|2|И простер царь к Есфири золотой скипетр, который был в руке его, и подошла Есфирь и коснулась конца скипетра,
ESTH|5|3|И сказал ей царь: что тебе, царица Есфирь, и какая просьба твоя? Даже до полуцарства будет дано тебе.
ESTH|5|4|И сказала Есфирь: если царю благоугодно, пусть придет царь с Аманом сегодня на пир, который я приготовила ему.
ESTH|5|5|И сказал царь: сходите скорее за Аманом, чтобы сделать по слову Есфири. И пришел царь с Аманом на пир, который приготовила Есфирь.
ESTH|5|6|И сказал царь Есфири при питье вина: какое желание твое? оно будет удовлетворено; и какая просьба твоя? [хотя бы] до полуцарства, она будет исполнена.
ESTH|5|7|И отвечала Есфирь, и сказала: [вот] мое желание и моя просьба:
ESTH|5|8|если я нашла благоволение в очах царя, и если царю благоугодно удовлетворить желание мое и исполнить просьбу мою, то пусть царь с Аманом придет на пир, который я приготовлю для них, и завтра я исполню слово царя.
ESTH|5|9|И вышел Аман в тот день веселый и благодушный. Но когда увидел Аман Мардохея у ворот царских, и тот не встал и с места не тронулся пред ним, тогда исполнился Аман гневом на Мардохея.
ESTH|5|10|Однако же скрепился Аман. А когда пришел в дом свой, то послал позвать друзей своих и Зерешь, жену свою.
ESTH|5|11|И рассказывал им Аман о великом богатстве своем и о множестве сыновей своих и обо всем том, как возвеличил его царь и как вознес его над князьями и слугами царскими.
ESTH|5|12|И сказал Аман: да и царица Есфирь никого не позвала с царем на пир, который она приготовила, кроме меня; так и на завтра я зван к ней с царем.
ESTH|5|13|Но всего этого не довольно для меня, доколе я вижу Мардохея Иудеянина сидящим у ворот царских.
ESTH|5|14|И сказала ему Зерешь, жена его, и все друзья его: пусть приготовят дерево вышиною в пятьдесят локтей, и утром скажи царю, чтобы повесили Мардохея на нем, и тогда весело иди на пир с царем. И понравилось это слово Аману, и он приготовил дерево.
ESTH|6|1|В ту ночь Господь отнял сон от царя, и он велел принести памятную книгу дневных записей; и читали их пред царем,
ESTH|6|2|и найдено записанным [там], как донес Мардохей на Гавафу Ифарру, двух евнухов царских, оберегавших порог, которые замышляли наложить руку на царя Артаксеркса.
ESTH|6|3|И сказал царь: какая дана почесть и отличие Мардохею за это? И сказали отроки царя, служившие при нем: ничего не сделано ему.
ESTH|6|4|И сказал царь: кто на дворе? Аман же пришел [тогда] на внешний двор царского дома поговорить с царем, чтобы повесили Мардохея на дереве, которое он приготовил для него.
ESTH|6|5|И сказали отроки царю: вот, Аман стоит на дворе. И сказал царь: пусть войдет.
ESTH|6|6|И вошел Аман. И сказал ему царь: что сделать бы тому человеку, которого царь хочет отличить почестью? Аман подумал в сердце своем: кому [другому] захочет царь оказать почесть, кроме меня?
ESTH|6|7|И сказал Аман царю: тому человеку, которого царь хочет отличить почестью,
ESTH|6|8|пусть принесут одеяние царское, в которое одевается царь, и [приведут] коня, на котором ездит царь, возложат царский венец на голову его,
ESTH|6|9|и пусть подадут одеяние и коня в руки одному из первых князей царских, – и облекут того человека, которого царь хочет отличить почестью, и выведут его на коне на городскую площадь, и провозгласят пред ним: так делается тому человеку, которого царь хочет отличить почестью!
ESTH|6|10|И сказал царь Аману: тотчас же возьми одеяние и коня, как ты сказал, и сделай это Мардохею Иудеянину, сидящему у царских ворот; ничего не опусти из всего, что ты говорил.
ESTH|6|11|И взял Аман одеяние и коня и облек Мардохея, и вывел его на коне на городскую площадь и провозгласил пред ним: так делается тому человеку, которого царь хочет отличить почестью!
ESTH|6|12|И возвратился Мардохей к царским воротам. Аман же поспешил в дом свой, печальный и закрыв голову.
ESTH|6|13|И пересказал Аман Зереши, жене своей, и всем друзьям своим все, что случилось с ним. И сказали ему мудрецы его и Зерешь, жена его: если из племени Иудеев Мардохей, из–за которого ты начал падать, то не пересилишь его, а наверно падешь пред ним.
ESTH|6|14|Они еще разговаривали с ним, [как] пришли евнухи царя и стали торопить Амана идти на пир, который приготовила Есфирь.
ESTH|7|1|И пришел царь с Аманом пировать у Есфири царицы.
ESTH|7|2|И сказал царь Есфири также и в [этот] второй день во время пира: какое желание твое, царица Есфирь? оно будет удовлетворено; и какая просьба твоя? [хотя бы] до полуцарства, она будет исполнена.
ESTH|7|3|И отвечала царица Есфирь и сказала: если я нашла благоволение в очах твоих, царь, и если царю благоугодно, то да будут дарованы мне жизнь моя, по желанию моему, и народ мой, по просьбе моей!
ESTH|7|4|Ибо проданы мы, я и народ мой, на истребление, убиение и погибель. Если бы мы проданы были в рабы и рабыни, я молчала бы, хотя враг не вознаградил бы ущерба царя.
ESTH|7|5|И отвечал царь Артаксеркс и сказал царице Есфири: кто это такой, и где тот, который отважился в сердце своем сделать так?
ESTH|7|6|И сказала Есфирь: враг и неприятель – этот злобный Аман! И Аман затрепетал пред царем и царицею.
ESTH|7|7|И царь встал во гневе своем с пира [и пошел] в сад при дворце; Аман же остался умолять о жизни своей царицу Есфирь, ибо видел, что определена ему злая участь от царя.
ESTH|7|8|Когда царь возвратился из сада при дворце в дом пира, Аман был припавшим к ложу, на котором находилась Есфирь. И сказал царь: даже и насиловать царицу [хочет] в доме у меня! Слово вышло из уст царя, – и накрыли лице Аману.
ESTH|7|9|И сказал Харбона, один из евнухов при царе: вот и дерево, которое приготовил Аман для Мардохея, говорившего доброе для царя, стоит у дома Амана, вышиною в пятьдесят локтей. И сказал царь: повесьте его на нем.
ESTH|7|10|И повесили Амана на дереве, которое он приготовил для Мардохея. И гнев царя утих.
ESTH|8|1|В тот день царь Артаксеркс отдал царице Есфири дом Амана, врага Иудеев; а Мардохей вошел пред лице царя, ибо Есфирь объявила, что он для нее.
ESTH|8|2|И снял царь перстень свой, который он отнял у Амана, и отдал его Мардохею; Есфирь же поставила Мардохея смотрителем над домом Амана.
ESTH|8|3|И продолжала Есфирь говорить пред царем и пала к ногам его, и плакала и умоляла его отвратить злобу Амана Вугеянина и замысел его, который он замыслил против Иудеев.
ESTH|8|4|И простер царь к Есфири золотой скипетр; и поднялась Есфирь, и стала пред лицем царя,
ESTH|8|5|и сказала: если царю благоугодно, и если я нашла благоволение пред лицем его, и справедливо дело сие пред лицем царя, и нравлюсь я очам его, то пусть было бы написано, чтобы возвращены были письма по замыслу Амана, сына Амадафа, Вугеянина, писанные им об истреблении Иудеев во всех областях царя;
ESTH|8|6|ибо, как я могу видеть бедствие, которое постигнет народ мой, и как я могу видеть погибель родных моих?
ESTH|8|7|И сказал царь Артаксеркс царице Есфири и Мардохею Иудеянину: вот, я дом Амана отдал Есфири, и его самого повесили на дереве за то, что он налагал руку свою на Иудеев;
ESTH|8|8|напишите и вы о Иудеях, что вам угодно, от имени царя и скрепите царским перстнем, ибо письма, написанного от имени царя и скрепленного перстнем царским, нельзя изменить.
ESTH|8|9|И позваны были тогда царские писцы в третий месяц, то есть в месяц Сиван, в двадцать третий день его, и написано было все так, как приказал Мардохей, к Иудеям, и к сатрапам, и областеначальникам, и правителям областей от Индии до Ефиопии, ста двадцати семи областей, в каждую область письменами ее и к каждому народу на языке его, и к Иудеям письменами их и на языке их.
ESTH|8|10|И написал он от имени царя Артаксеркса, и скрепил царским перстнем, и послал письма чрез гонцов на конях, на дромадерах и мулах царских,
ESTH|8|11|о том, что царь позволяет Иудеям, находящимся во всяком городе, собраться и стать на защиту жизни своей, истребить, убить и погубить всех сильных в народе и в области, которые во вражде с ними, детей и жен, и имение их разграбить,
ESTH|8|12|в один день по всем областям царя Артаксеркса, в тринадцатый день двенадцатого месяца, то есть месяца Адара.
ESTH|8|13|Список с сего указа отдать в каждую область, [как] закон, объявляемый для всех народов, чтоб Иудеи готовы были к тому дню мстить врагам своим.
ESTH|8|14|Гонцы, поехавшие верхом на быстрых конях царских, погнали скоро и поспешно, с царским повелением. Объявлен был указ и в Сузах, престольном городе.
ESTH|8|15|И Мардохей вышел от царя в царском одеянии яхонтового и белого цвета и в большом золотом венце, и в мантии виссонной и пурпуровой. И город Сузы возвеселился и возрадовался.
ESTH|8|16|А у Иудеев было [тогда] освещение и радость, и веселье, и торжество.
ESTH|8|17|И во всякой области и во всяком городе, во [всяком] месте, куда [только] доходило повеление царя и указ его, была радость у Иудеев и веселье, пиршество и праздничный день. И многие из народов страны сделались Иудеями, потому что напал на них страх пред Иудеями.
ESTH|9|1|В двенадцатый месяц, то есть в месяц Адар, в тринадцатый день его, в который пришло время исполниться повелению царя и указу его, в тот день, когда надеялись неприятели Иудеев взять власть над ними, а вышло наоборот, что сами Иудеи взяли власть над врагами своими, –
ESTH|9|2|собрались Иудеи в городах своих по всем областям царя Артаксеркса, чтобы наложить руку на зложелателей своих; и никто не мог устоять пред лицем их, потому что страх пред ними напал на все народы.
ESTH|9|3|И все князья в областях и сатрапы, и областеначальники, и исполнители дел царских поддерживали Иудеев, потому что напал на них страх пред Мардохеем.
ESTH|9|4|Ибо велик был Мардохей в доме у царя, и слава о нем ходила по всем областям, так как сей человек, Мардохей, поднимался выше и выше.
ESTH|9|5|И избивали Иудеи всех врагов своих, побивая мечом, умерщвляя и истребляя, и поступали с неприятелями своими по своей воле.
ESTH|9|6|В Сузах, городе престольном, умертвили Иудеи и погубили пятьсот человек;
ESTH|9|7|и Паршандафу и Далфона и Асфафу,
ESTH|9|8|и Порафу и Адалью и Аридафу,
ESTH|9|9|и Пармашфу и Арисая и Аридая и Ваиезафу, –
ESTH|9|10|десятерых сыновей Амана, сына Амадафа, врага Иудеев, умертвили они, а на грабеж не простерли руки своей.
ESTH|9|11|В тот же день донесли царю о числе умерщвленных в Сузах, престольном городе.
ESTH|9|12|И сказал царь царице Есфири: в Сузах, городе престольном, умертвили Иудеи и погубили пятьсот человек и десятерых сыновей Амана; что же сделали они в прочих областях царя? Какое желание твое? и оно будет удовлетворено. И какая еще просьба твоя? она будет исполнена.
ESTH|9|13|И сказала Есфирь: если царю благоугодно, то пусть бы позволено было Иудеям, которые в Сузах, делать то же и завтра, что сегодня, и десятерых сыновей Амановых пусть бы повесили на дереве.
ESTH|9|14|И приказал царь сделать так; и дан [на это] указ в Сузах, и десятерых сыновей Амановых повесили.
ESTH|9|15|И собрались Иудеи, которые в Сузах, также и в четырнадцатый день месяца Адара и умертвили в Сузах триста человек, а на грабеж не простерли руки своей.
ESTH|9|16|И прочие Иудеи, находившиеся в царских областях, собрались, чтобы стать на защиту жизни своей и быть покойными от врагов своих, и умертвили из неприятелей своих семьдесят пять тысяч, а на грабеж не простерли руки своей.
ESTH|9|17|[Это было] в тринадцатый день месяца Адара; а в четырнадцатый день сего же месяца они успокоились и сделали его днем пиршества и веселья.
ESTH|9|18|Иудеи же, которые в Сузах, собирались в тринадцатый день его и в четырнадцатый день его, а в пятнадцатый день его успокоились и сделали его днем пиршества и веселья.
ESTH|9|19|Поэтому Иудеи сельские, живущие в селениях открытых, проводят четырнадцатый день месяца Адара в веселье и пиршестве, как день праздничный, посылая подарки друг ко другу.
ESTH|9|20|И описал Мардохей эти происшествия и послал письма ко всем Иудеям, которые в областях царя Артаксеркса, к близким и к дальним,
ESTH|9|21|[о том], чтобы они установили каждогодно празднование у себя четырнадцатого дня месяца Адара и пятнадцатого дня его,
ESTH|9|22|как таких дней, в которые Иудеи сделались покойны от врагов своих, и [как] такого месяца, в который превратилась у них печаль в радость, и сетование – в день праздничный, – чтобы сделали их днями пиршества и веселья, посылая подарки друг другу и подаяния бедным.
ESTH|9|23|И приняли Иудеи то, что уже сами начали делать, и о чем Мардохей написал к ним,
ESTH|9|24|как Аман, сын Амадафа, Вугеянин, враг всех Иудеев, думал погубить Иудеев и бросал пур, [жребий], об истреблении и погублении их,
ESTH|9|25|и как Есфирь дошла до царя, и как царь приказал новым письмом, чтобы злой замысл Амана, который он задумал на Иудеев, обратился на голову его, и чтобы повесили его и сыновей его на дереве.
ESTH|9|26|Потому и назвали эти дни Пурим, от имени: пур. Поэтому, согласно со всеми словами сего письма и с тем, что сами видели и до чего доходило у них,
ESTH|9|27|постановили Иудеи и приняли на себя и на детей своих и на всех, присоединяющихся к ним, неотменно, чтобы праздновать эти два дня, по предписанному о них и в свое для них время, каждый год;
ESTH|9|28|и чтобы дни эти были памятны и празднуемы во все роды в каждом племени, в каждой области и в каждом городе; и чтобы дни эти Пурим не отменялись у Иудеев, и память о них не исчезла у детей их.
ESTH|9|29|Написала также царица Есфирь, дочь Абихаила, и Мардохей Иудеянин, со всею настойчивостью, чтобы исполняли это новое письмо о Пуриме;
ESTH|9|30|и послали письма ко всем Иудеям в сто двадцать семь областей царства Артаксерксова со словами мира и правды,
ESTH|9|31|чтобы они твердо наблюдали эти дни Пурим в свое время, какое уставил о них Мардохей Иудеянин и царица Есфирь, и как они сами назначали их для себя и для детей своих в дни пощения и воплей.
ESTH|9|32|Так повеление Есфири подтвердило это слово о Пуриме, и оно вписано в книгу.
ESTH|10|1|Потом наложил царь Артаксеркс подать на землю и на острова морские.
ESTH|10|2|Впрочем, все дела силы его и могущества его и обстоятельное показание о величии Мардохея, которым возвеличил его царь, записаны в книге дневных записей царей Мидийских и Персидских,
ESTH|10|3|[равно как и то], что Мардохей Иудеянин [был] вторым по царе Артаксерксе и великим у Иудеев и любимым у множества братьев своих, [ибо] искал добра народу своему и говорил во благо всего племени своего.
