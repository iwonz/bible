ESTH|1|1|Et fuit in diebus Asueri, qui regnavit ab India usque Aethiopiam super centum viginti septem provincias,
ESTH|1|2|quando sedit in solio regni sui in castris Susan,
ESTH|1|3|tertio igitur anno imperii sui, fecit grande convivium cunctis principibus et pueris suis, fortissimis Persarum et Medorum, inclitis et praefectis provinciarum coram se,
ESTH|1|4|ut ostenderet divitias gloriae regni sui ac splendorem atque iactantiam magnitudinis suae multo tempore, centum videlicet et octoginta diebus.
ESTH|1|5|Cumque implerentur dies convivii, invitavit omnem populum, qui inventus est in Susan, a maximo usque ad minimum; et septem diebus iussit convivium praeparari in vestibulo horti palatii regis.
ESTH|1|6|Et pendebant ex omni parte tentoria lintea et carbasina ac hyacinthina sustentata funibus byssinis atque purpureis, qui argenteis circulis inserti erant et columnis marmoreis fulciebantur; lectuli quoque aurei et argentei dispositi erant super pavimentum smaragdino et pario stratum lapide aliisque varii coloris.
ESTH|1|7|Bibebant autem, qui invitati erant, aureis poculis, aliis atque aliis; vinum quoque, ut magnificentia regia dignum erat, abundans et praecipuum ponebatur.
ESTH|1|8|Nec erat qui cogeret ad bibendum, quoniam sic rex statuerat omnibus praepositis domus suae, ut facerent secundum uniuscuiusque voluntatem.
ESTH|1|9|Vasthi quoque regina fecit convivium feminarum in palatio regio, ubi rex Asuerus manere consueverat.
ESTH|1|10|Itaque die septimo, cum rex esset hilarior potione meri, praecepit Mauman et Bazatha et Harbona et Bagatha et Abgatha et Zethar et Charchas, septem eunuchis, qui in conspectu eius ministrabant,
ESTH|1|11|ut introducerent reginam Vasthi coram rege, posito super caput eius diademate regni, ut ostenderet cunctis populis et principibus pulchritudinem illius; erat enim pulchra valde.
ESTH|1|12|Quae renuit et ad regis imperium, quod per eunuchos mandaverat, venire contempsit; unde iratus rex et nimio furore succensus
ESTH|1|13|interrogavit sapientes, qui tempora noverant, et illorum faciebat cuncta consilio scientium leges ac iura maiorum -
ESTH|1|14|erant autem ei proximi Charsena et Sethar et Admatha et Tharsis et Mares et Marsana et Mamuchan, septem duces Persarum atque Medorum, qui videbant faciem regis et primi sedebant in regno C:
ESTH|1|15|" Secundum legem quid oportet fieri Vasthi reginae, quae Asueri regis imperium, quod per eunuchos mandaverat, facere noluit? ".
ESTH|1|16|Responditque Mamuchan, audiente rege atque principibus: " Non solum regem laesit regina Vasthi, sed et omnes principes et populos, qui sunt in cunctis provinciis regis Asueri.
ESTH|1|17|Egredietur enim sermo reginae ad omnes mulieres, ut contemnant viros suos et dicant: "Rex Asuerus iussit, ut regina Vasthi intraret ad eum, et illa noluit".
ESTH|1|18|Atque hac ipsa die dicent omnes principum coniuges Persarum atque Medorum quem audierint sermonem reginae principibus regis; unde despectio et indignatio.
ESTH|1|19|Si tibi, rex, placet, egrediatur edictum a facie tua et scribatur inter leges Persarum atque Medorum, quas immutari illicitum est, ut nequaquam ultra Vasthi ingrediatur ad regem, sed regnum illius altera, quae melior illa est, accipiat.
ESTH|1|20|Et hoc in omne, quod latissimum est, provinciarum tuarum divulgetur imperium, et cunctae uxores, tam maiorum quam minorum, deferent maritis suis honorem ".
ESTH|1|21|Placuit consilium eius regi et principibus, fecitque rex iuxta consilium Mamuchan.
ESTH|1|22|Et misit epistulas ad universas provincias regni sui, ut quaeque gens audire et legere poterat, diversis linguis et litteris, esse viros principes ac maiores in domibus suis et subditas habere omnes mulieres, quae essent cum eis.
ESTH|2|1|His ita gestis, postquam regis Asueri deferbuerat indignatio, recordatus est Vasthi, et quae fecisset vel quae passa esset.
ESTH|2|2|Dixeruntque pueri regis ac ministri eius: " Quaerantur regi puellae virgines ac speciosae,
ESTH|2|3|et constituantur, qui considerent per universas provincias puellas speciosas et virgines et adducant eas ad civitatem Susan et tradant in domum feminarum sub manu Egei eunuchi, qui est praepositus et custos mulierum regiarum; et accipiant mundum muliebrem.
ESTH|2|4|Et, quaecumque inter omnes oculis regis placuerit, ipsa regnet pro Vasthi ". Placuit sermo regi; et ita, ut suggesserant, iussit fieri.
ESTH|2|5|Erat vir Iudaeus in Susan civitate vocabulo Mardochaeus filius Iair filii Semei filii Cis de tribu Beniamin,
ESTH|2|6|qui translatus fuerat de Ierusalem cum captivis, qui ducti fuerant cum Iechonia rege Iudae, quem Nabuchodonosor rex Babylonis transtulerat.
ESTH|2|7|Qui fuit nutricius filiae patrui sui Edissae, quae altero nomine Esther vocabatur et utrumque parentem amiserat: pulchra aspectu et decora facie. Mortuisque patre eius ac matre, Mardochaeus sibi eam adoptavit in filiam.
ESTH|2|8|Et factum est, cum percrebruisset regis imperium, et iuxta mandatum illius multae virgines pulchrae adducerentur Susan et Egeo traderentur, Esther quoque in domum regis in manus Egei custodis feminarum tradita est.
ESTH|2|9|Quae placuit ei et invenit gratiam in conspectu illius; et acceleravit mundum muliebrem et tradidit ei partes suas et septem puellas speciosissimas de domo regis, et tam ipsam quam pedisequas eius transtulit in optimam partem domus feminarum.
ESTH|2|10|Quae non indicaverat ei populum et cognationem suam; Mardochaeus enim praeceperat, ut de hac re omnino reticeret.
ESTH|2|11|Qui deambulabat cotidie ante vestibulum domus, in qua electae virgines servabantur, curam agens salutis Esther et scire volens quid ei accideret.
ESTH|2|12|Cum autem venisset tempus singularum per ordinem puellarum, ut intrarent ad regem, expletis omnibus, quae ad cultum muliebrem pertinebant, per menses duodecim; ita dumtaxat, ut sex mensibus oleo ungerentur myrrhino et aliis sex feminarum pigmentis et aromatibus uterentur,
ESTH|2|13|ingredientesque ad regem, quidquid postulassent, accipiebant, ut portarent secum de triclinio feminarum ad regis cubiculum.
ESTH|2|14|Et, quae intraverat vespere, mane iterum in domum feminarum deducebatur, sub manu Sasagazi eunuchi, qui concubinis praesidebat. Nec habebat potestatem ad regem ultra redeundi, nisi voluisset rex et eam venire iussisset ex nomine.
ESTH|2|15|Evoluto autem tempore per ordinem, instabat dies, quo Esther filia Abihail patrui Mardochaei, quam sibi adoptaverat in filiam, intrare deberet ad regem. Quae non quaesivit quidquam, nisi quae voluit Egeus eunuchus custos feminarum, et omnium oculis gratiosa et amabilis videbatur.
ESTH|2|16|Ducta est itaque ad cubiculum regis Asueri mense decimo, qui vocatur Tebeth, septimo anno regni eius.
ESTH|2|17|Et amavit eam rex plus quam omnes mulieres; habuitque gratiam et favorem coram eo super omnes virgines, et posuit diadema regni in capite eius fecitque eam regnare in loco Vasthi.
ESTH|2|18|Et iussit convivium praeparari magnificum cunctis principibus et servis suis, convivium Esther; et dedit remissionem tributi universis provinciis ac dona largitus est iuxta magnificentiam principalem.
ESTH|2|19|Mardochaeus autem manebat ad regis ianuam,
ESTH|2|20|necdum prodiderat Esther cognationem et populum suum iuxta mandatum eius; quidquid enim ille praecipiebat, observabat Esther, ut eo tempore solita erat, quo eam parvulam nutriebat.
ESTH|2|21|Eo igitur tempore, quo Mardochaeus ad regis ianuam morabatur, irati sunt Bagathan et Thares, duo eunuchi regis, qui ianitores erant volueruntque in regem mittere manus.
ESTH|2|22|Quod Mardochaeum non latuit; statimque nuntiavit reginae Esther, et illa regi ex nomine Mardochaei.
ESTH|2|23|Quaesitum est et inventum, et appensus uterque eorum in patibulo; mandatumque est libro annalium coram rege.
ESTH|3|1|Post haec rex Asuerus exaltavit Aman filium Amadathi, qui erat de stirpe Agag, et posuit solium eius super omnes principes, quos habebat.
ESTH|3|2|Cunctique servi regis, qui in foribus palatii versabantur, flectebant genua et adorabant Aman; sic enim praeceperat rex pro illo. Solus Mardochaeus non flectebat genu neque adorabat eum.
ESTH|3|3|Cui dixerunt pueri regis, qui ad fores palatii praesidebant: " Cur non observas mandatum regis? ".
ESTH|3|4|Cumque hoc crebrius dicerent, et ille nollet audire, nuntiaverunt Aman scire cupientes utrum perseveraret in sententia; dixerat enim eis se esse Iudaeum.
ESTH|3|5|Cumque Aman experimento probasset quod Mardochaeus non sibi flecteret genu nec se adoraret, iratus est valde
ESTH|3|6|et pro nihilo duxit in unum Mardochaeum mittere manus suas - audierat enim quod esset gentis Iudaeae - magisque voluit omnem Iudaeorum, qui erant in regno Asueri, perdere nationem.
ESTH|3|7|Mense primo, cuius vocabulum est Nisan, anno duodecimo regni Asueri, missa est in urnam sors, quae dicitur Phur, coram Aman, quo die et quo mense gens Iudaeorum deberet interfici; et exivit dies tertia decima mensis duodecimi, qui vocatur Adar.
ESTH|3|8|Dixitque Aman regi Asuero: " Est populus per omnes provincias regni tui dispersus, segregatus inter populos alienisque utens legibus, quas ceteri non cognoscunt, insuper et regis scita contemnens; non expedit regi, ut det illis requiem.
ESTH|3|9|Si tibi placet, scriptis decerne, ut pereat, et decem milia talentorum argenti appendam arcariis gazae tuae ".
ESTH|3|10|Tulit ergo rex anulum, quo utebatur, de manu sua et dedit eum Aman filio Amadathi de progenie Agag, hosti Iudaeorum.
ESTH|3|11|Dixitque ad eum: " Argentum, quod polliceris, tuum sit; de populo age, quod tibi placet ".
ESTH|3|12|Vocatique sunt scribae regis mense primo, tertia decima die eius, et scriptum est, ut iusserat Aman, ad omnes satrapas regis et duces provinciarum et principes diversarum gentium, ut quaeque gens legere poterat et audire pro varietate linguarum, ex nomine regis Asueri; et litterae ipsius signatae anulo.
ESTH|3|13|Missae sunt epistulae per cursores ad universas provincias regis, ut perderent, occiderent atque delerent omnes Iudaeos, a puero usque ad senem, parvulos et mulieres uno die, hoc est tertio decimo mensis duodecimi, qui vocatur Adar, et bona eorum diriperent.
ESTH|3|14|Exemplar autem epistularum ut lex in omnibus provinciis promulgandum erat, ut scirent omnes populi et pararent se ad praedictam diem.
ESTH|3|15|Festinabant cursores, qui missi erant, regis imperium explere; statimque in Susan pependit edictum, rege et Aman celebrante convivium, dum civitas ipsa esset conturbata.
ESTH|4|1|Cum comperisset Mardochaeus omnia, quae acciderant, scidit vestimenta sua et indutus est sacco spargens cinerem capiti. Et in platea mediae civitatis voce magna et amara clamabat
ESTH|4|2|usque ad fores palatii gradiens; non enim erat licitum indutum sacco aulam regis intrare.
ESTH|4|3|In omnibus quoque provinciis, quocumque edictum et dogma regis pervenerat, planctus ingens erat apud Iudaeos, ieiunium, ululatus et fletus, sacco et cinere multis pro strato utentibus.
ESTH|4|4|Ingressae sunt autem puellae Esther et eunuchi nuntiaveruntque ei. Quod audiens consternata est valde et misit vestem, ut, ablato sacco, induerent eum; quam accipere noluit.
ESTH|4|5|Accitoque Athach eunucho, quem rex ministrum ei dederat, praecepit ei, ut iret ad Mardochaeum et disceret ab eo cur hoc faceret.
ESTH|4|6|Egressusque Athach ivit ad Mardochaeum stantem in platea civitatis ante ostium palatii.
ESTH|4|7|Qui indicavit ei omnia, quae ei acciderant, quantum Aman promisisset, ut in thesauros regis pro Iudaeorum nece inferret argentum.
ESTH|4|8|Exemplar quoque edicti, quod pendebat in Susan ad perdendum eos, dedit ei, ut reginae ostenderet et moneret eam, ut intraret ad regem et deprecaretur eum et rogaret pro populo suo. 8a " Memor, inquit, dierum humilitatis tuae, quando nutrita sis in manu mea, quia Aman secundus a rege locutus est contra nos in mortem. Et tu, invoca Dominum et loquere regi pro nobis et libera nos de morte ".
ESTH|4|9|Regressus Athach nuntiavit Esther omnia, quae Mardochaeus dixerat.
ESTH|4|10|Quae respondit ei et iussit, ut diceret Mardochaeo:
ESTH|4|11|" Omnes servi regis et cunctae, quae sub dicione eius sunt, norunt provinciae, quod cuique sive viro sive mulieri, qui non vocatus interius atrium regis intraverit, una lex sit, ut statim interficiatur, nisi forte rex auream virgam ad eum tetenderit, ut possit vivere; ego autem triginta iam diebus non sum vocata ad regem ".
ESTH|4|12|Quod cum audisset Mardochaeus,
ESTH|4|13|rursum mandavit Esther dicens: " Ne putes quod animam tuam tantum liberes, quia in domo regis es, prae cunctis Iudaeis.
ESTH|4|14|Si enim nunc silueris, aliunde Iudaeis liberatio et salvatio exsurget, et tu et domus patris tui peribitis; et quis novit utrum idcirco ad regnum veneris, ut in tali tempore parareris? ".
ESTH|4|15|Rursumque Esther haec Mardochaeo verba mandavit:
ESTH|4|16|" Vade et congrega omnes Iudaeos, qui in Susan reperiuntur; et ieiunate pro me. Non comedatis et non bibatis tribus diebus et tribus noctibus, et ego cum ancillis meis similiter ieiunabo; et tunc ingrediar ad regem contra legem faciens; si pereo, pereo ".
ESTH|4|17|Ivit itaque Mardochaeus et fecit omnia, quae ei Esther mandaverat.
ESTH|5|1|Et factum est die tertio, induta Esther regalibus vestimentis ste tit in atrio domus regiae, quod erat interius contra basilicam regis. At ille sedebat super solium suum in consistorio palatii contra ostium domus.
ESTH|5|2|Et factum est, cum vidisset Esther reginam stantem, placuit oculis eius, et extendit contra eam virgam auream, quam tenebat manu; quae accedens tetigit summitatem virgae eius.
ESTH|5|3|Dixitque ad eam rex: " Quid vis, Esther regina? Quae est petitio tua? Etiamsi dimidiam partem regni petieris, dabitur tibi ".
ESTH|5|4|At illa respondit: " Si regi placet, obsecro, ut venias ad me hodie et Aman tecum ad convivium, quod paravi ".
ESTH|5|5|Statimque rex: " Vocate, inquit, cito Aman, ut fiat verbum Esther ".Venerunt itaque rex et Aman ad convivium, quod eis regina paraverat.
ESTH|5|6|Dixitque ei rex, postquam vinum biberat: " Quid petis, ut detur tibi, et pro qua re postulas? Etiamsi dimidiam partem regni mei petieris, impetrabis ".
ESTH|5|7|Cui respondit Esther: " Petitio mea et preces:
ESTH|5|8|Si inveni in conspectu regis gratiam, et si regi placet, ut det mihi, quod postulo, et meam impleat petitionem, veniat rex et Aman ad convivium, quod parabo eis, et cras faciam secundum verbum regis ".
ESTH|5|9|Egressus est itaque illo die Aman laetus et alacer corde. Cumque vidisset Mardochaeum sedentem in foribus palatii, et non solum non assurrexisse sibi, sed nec motum quidem de loco sessionis suae, indignatus est valde.
ESTH|5|10|Et, dissimulata ira, reversus in domum suam convocavit ad se amicos suos et Zares uxorem suam
ESTH|5|11|et exposuit illis magnitudinem divitiarum suarum filiorumque turbam, et quanta eum gloria super omnes principes et servos suos rex elevasset.
ESTH|5|12|Et post haec ait: " Regina quoque Esther nullum alium vocavit ad convivium cum rege praeter me; apud quam etiam cras cum rege pransurus sum.
ESTH|5|13|Et, cum omnia haec habeam, nihil me habere puto, quamdiu videro Mardochaeum Iudaeum sedentem in foribus regis ".
ESTH|5|14|Responderuntque ei Zares uxor eius et ceteri amici: " Iube parari excelsam trabem habentem altitudinis quinquaginta cubitos et dic mane regi, ut appendatur super eam Mardochaeus; et sic ibis cum rege laetus ad convivium ". Placuit ei consilium et iussit excelsam parari trabem.
ESTH|6|1|Noctem illam duxit rex insomnem iussitque afferri sibi librum memorialium, annales priorum temporum. Quae cum illo praesente legerentur,
ESTH|6|2|ventum est ad eum locum, ubi scriptum erat quomodo nuntiasset Mardochaeus insidias Bagathan et Thares duorum eunuchorum ianitorum, qui voluerant manus mittere in regem Asuerum.
ESTH|6|3|Quod cum audisset rex, ait: " Quid pro hac fide honoris ac praemii Mardochaeus consecutus est? ". Dixeruntque ei servi illius ac ministri: " Nihil omnino mercedis accepit ".
ESTH|6|4|Statimque rex: " Quis est, inquit, in atrio? ". Aman quippe exterius atrium domus regiae intraverat, ut suggereret regi, ut iuberet Mardochaeum suspendi in patibulo, quod ei fuerat praeparatum.
ESTH|6|5|Responderunt pueri: " Ecce Aman stat in atrio ". Dixitque rex: " Ingrediatur ".
ESTH|6|6|Cumque esset ingressus, ait illi: " Quid debet fieri viro, quem rex honorare desiderat? ". Cogitans autem in corde suo Aman et reputans quod nullum alium rex nisi se vellet honorare
ESTH|6|7|respondit: " Homo, quem rex honorare cupit,
ESTH|6|8|debet indui vestibus regiis, quibus rex indutus erat, et imponi super equum, qui de sella regis est, et acceperit regium diadema super caput suum;
ESTH|6|9|et primus de regiis principibus nobilissimis induat eum et teneat equum eius et per plateam civitatis incedens clamet et dicat: "Sic honorabitur quemcumque voluerit rex honorare" ".
ESTH|6|10|Dixitque ei rex: " Festina et, sumpta stola et equo, fac, ut locutus es, Mardochaeo Iudaeo, qui sedet in foribus palatii; cave, ne quidquam de his, quae locutus es, praetermittas ".
ESTH|6|11|Tulit itaque Aman stolam et equum; indutumque Mardochaeum et impositum equo praecedebat in platea civitatis atque clamabat: " Hoc honore condignus est quemcumque rex voluerit honorare ".
ESTH|6|12|Reversusque est Mardochaeus ad ianuam palatii; et Aman festinavit ire in domum suam lugens et operto capite.
ESTH|6|13|Narravitque Zares uxori suae et amicis omnia, quae evenissent sibi; cui responderunt sapientes, quos habebat in consilio, et uxor eius: " Si de semine Iudaeorum est Mardochaeus, ante quem cadere coepisti, non poteris praevalere contra eum, sed cades in conspectu eius ".
ESTH|6|14|Adhuc illis loquentibus, venerunt eunuchi regis et cito eum ad convivium, quod regina paraverat, pergere compulerunt.
ESTH|7|1|Intravit itaque rex et Aman, ut biberent cum regina.
ESTH|7|2|Dixitque ei rex etiam in secundo die, postquam vino incaluerat: " Quae est petitio tua, Esther, ut detur tibi, et quid vis fieri? Etiamsi dimidiam regni mei partem petieris, impetrabis ".
ESTH|7|3|Ad quem illa respondit: " Si inveni gratiam in oculis tuis, o rex, et si tibi placet, dona mihi animam meam, pro qua rogo, et populum meum, pro quo obsecro.
ESTH|7|4|Traditi enim sumus, ego et populus meus, ut conteramur, iugulemur et pereamus. Atque utinam in servos et famulas venderemur: tacuissem, quia tribulatio haec non esset digna conturbare regem ".
ESTH|7|5|Respondensque rex Asuerus ait: " Quis est iste et ubi est, ut haec audeat facere? ".
ESTH|7|6|Dixit Esther: " Hostis et inimicus noster pessimus iste est Aman ". Quod ille audiens ilico obstupuit coram rege ac regina.
ESTH|7|7|Rex autem surrexit iratus et de loco convivii intravit in hortum palatii. Aman quoque surrexit, ut rogaret Esther reginam pro anima sua; intellexit enim a rege sibi decretum esse malum.
ESTH|7|8|Qui cum reversus esset de horto et intrasset convivii locum, repperit Aman super lectulum corruisse, in quo iacebat Esther, et ait: " Etiam reginam vult opprimere, me praesente, in domo mea? ". Necdum verbum de ore regis exierat, et statim operuerunt faciem eius.
ESTH|7|9|Dixitque Harbona, unus de eunuchis, qui stabant in ministerio regis: " En etiam lignum, quod paraverat Mardochaeo, qui locutus est bonum pro rege, stat in domo Aman habens altitudinis quinquaginta cubitos ". Cui dixit rex: " Appendite eum in eo ".
ESTH|7|10|Suspensus est itaque Aman in patibulo, quod paraverat Mardochaeo; et regis ira quievit.
ESTH|8|1|Die illo dedit rex Asuerus Esther reginae domum Aman adversarii Iudaeorum, et Mardochaeus ingressus est ante faciem regis; confessa est enim ei Esther quid esset sibi.
ESTH|8|2|Tulitque rex anulum suum, quem ab Aman recipi iusserat, et tradidit Mardochaeo; Esther autem constituit Mardochaeum super domum Aman.
ESTH|8|3|Et adiecit Esther loqui coram rege et procidit ad pedes eius flevitque et locuta ad eum oravit, ut malitiam Aman Agagitae et machinationes eius pessimas, quas excogitaverat contra Iudaeos, iuberet irritas fieri.
ESTH|8|4|At ille ex more sceptrum aureum protendit manu; illaque consurgens stetit ante eum
ESTH|8|5|et ait: " Si placet regi, et si inveni gratiam coram eo, et deprecatio mea non ei videtur esse contraria, et accepta sum in oculis eius, obsecro, ut novis epistulis veteres litterae Aman filii Amadathi, Agagitae, insidiatoris et hostis Iudaeorum, quibus eos in cunctis regis provinciis perire praeceperat, corrigantur.
ESTH|8|6|Quomodo enim potero sustinere malum, quod passurus est populus meus, et interitum cognationis meae? ".
ESTH|8|7|Responditque rex Asuerus Esther reginae et Mardochaeo Iudaeo: " Domum Aman concessi Esther et ipsum iussi appendi in patibulo, quia ausus est manum in Iudaeos mittere.
ESTH|8|8|Scribite ergo Iudaeis sicut vobis placet, ex regis nomine, signantes litteras anulo meo, quia epistulae ex regis nomine scriptae et illius anulo signatae non possunt immutari ".
ESTH|8|9|Accitisque scribis regis - erat autem tempus tertii mensis, qui appellatur Sivan, vicesima et tertia illius die - scriptae sunt epistulae, ut Mardochaeus voluerat, ad Iudaeos et ad satrapas procuratoresque et principes, qui centum viginti septem provinciis ab India usque ad Aethiopiam praesidebant, provinciae atque provinciae, populo et populo, iuxta linguas et litteras suas, et Iudaeis iuxta linguam et litteras suas.
ESTH|8|10|Ipsaeque epistulae, quae ex regis nomine mittebantur, anulo ipsius obsignatae sunt et missae per veredarios electis equis regiis discurrentes.
ESTH|8|11|Quibus permisit rex Iudaeis in singulis civitatibus, ut in unum congregarentur et starent pro animabus suis et omnes inimicos suos cum coniugibus ac liberis interficerent atque delerent et spolia eorum diriperent;
ESTH|8|12|et constituta est per omnes provincias una ultionis dies, id est tertia decima mensis duodecimi, qui vocatur Adar.
ESTH|8|13|Exemplar epistulae in forma legis in omnibus provinciis promulgandum erat, ut omnibus populis notum fieret paratos esse Iudaeos in diem illam ad capiendam vindictam de hostibus suis.
ESTH|8|14|Egressique sunt veredarii celeres nuntios perferentes, et edictum regis pependit in Susan.
ESTH|8|15|Mardochaeus autem de palatio et de conspectu regis egrediens fulgebat vestibus regiis, hyacinthinis videlicet et albis, coronam magnam auream portans in capite et amictus pallio serico atque purpureo; omnisque civitas exsultavit atque laetata est.
ESTH|8|16|Iudaeis autem nova lux oriri visa est, gaudium, honor et tripudium.
ESTH|8|17|Apud omnes populos, urbes atque provincias, quocumque regis iussa veniebant, Iudaeis fuit exsultatio, epulae atque convivia et festus dies, in tantum ut plures alterius gentis et sectae eorum religioni et caeremoniis iungerentur; grandis enim cunctos Iudaici nominis terror invaserat.
ESTH|9|1|Igitur duodecimi mensis - id est Adar - tertia decima die, quando verbum et edictum regis explendum erat, et hostes Iudaeorum sperabant quod dominarentur ipsis, versa vice Iudaei superaverunt adversarios suos.
ESTH|9|2|Congregatique sunt per singulas civitates, ut extenderent manum contra inimicos et persecutores suos; nullusque ausus est resistere, eo quod omnes populos invaserat formido eorum.
ESTH|9|3|Nam et omnes provinciarum principes et satrapae et procuratores omnisque dignitas, quae singulis locis ac operibus praeerat, sustinebant Iudaeos timore Mardochaei,
ESTH|9|4|quem principem esse palatii et plurimum posse cognoverant; fama quoque nominis eius crescebat cotidie et per cunctorum ora volitabat.
ESTH|9|5|Itaque percusserunt Iudaei omnes inimicos suos plaga gladii et necis et interitus, reddentes eis, quod sibi paraverant facere.
ESTH|9|6|In Susan quingentos viros interfecerunt, extra decem filios Aman Agagitae hostis Iudaeorum, quorum ista sunt nomina:
ESTH|9|7|Pharsandatha et Delphon et Esphatha
ESTH|9|8|et Phoratha et Adalia et Aridatha
ESTH|9|9|et Phermesta et Arisai et Aridai et Iezatha.
ESTH|9|10|Quos cum occidissent, praedas de substantiis eorum tangere noluerunt.
ESTH|9|11|Statimque numerus eorum, qui occisi erant in Susan, ad regem relatus est.
ESTH|9|12|Qui dixit reginae: " In urbe Susan interfecerunt et deleverunt Iudaei quingentos viros et decem filios Aman. Quantam putas eos exercuisse caedem in universis provinciis? Quid ultra postulas et quid vis, ut fieri iubeam?.
ESTH|9|13|Cui illa respondit: " Si regi placet, detur potestas Iudaeis, qui in Susan sunt, ut sicut hodie fecerunt, sic et cras faciant, et decem filii Aman in patibulo suspendantur ".
ESTH|9|14|Praecepitque rex, ut ita fieret. Statimque in Susan pependit edictum, et decem filii Aman suspensi sunt.
ESTH|9|15|Congregatis igitur Iudaeis, qui in Susan erant, quarta decima die mensis Adar, interfecti sunt in Susan trecenti viri, nec eorum ab illis direpta substantia est.
ESTH|9|16|Reliqui autem Iudaei per omnes provincias, quae dicioni regis subiacebant, congregati pro animabus suis steterunt, ut requiescerent ab hostibus, ac interfecerunt de persecutoribus suis septuaginta quinque milia, sed nullus de substantiis eorum quidquam contigit.
ESTH|9|17|Dies autem tertius decimus mensis Adar, dies apud omnes interfectionis fuit, et quarta decima die requieverunt. Quem constituerunt esse diem epularum et laetitiae.
ESTH|9|18|At hi, qui in urbe Susan congregati sunt, tertio decimo et quarto decimo die eiusdem mensis in caede versati sunt, quinto decimo autem die requieverunt; et idcirco eundem diem constituerunt sollemnem epularum atque laetitiae.
ESTH|9|19|Hi vero Iudaei, qui in oppidis non muratis ac villis morabantur, quartum decimum diem mensis Adar conviviorum et gaudii decreverunt, ita ut exsultent in eo et mittant sibi mutuo partes epularum. Illi autem, qui in urbibus habitant, agunt etiam quintum decimum diem mensis Adar cum gaudio et convivio et ut diem festum, in quo mittunt sibi mutuo partes epularum.
ESTH|9|20|Scripsit itaque Mardochaeus omnia haec et litteris comprehensa misit ad omnes Iudaeos, qui in omnibus regis provinciis morabantur, tam in vicino positis quam procul,
ESTH|9|21|ut quartam decimam et quintam decimam diem mensis Adar pro festis susciperent et, revertente semper anno, sollemni honore celebrarent
ESTH|9|22|secundum dies, in quibus requieverunt Iudaei ab inimicis suis, et mensem, qui de luctu atque tristitia in hilaritatem gaudiumque ipsis conversus est, essentque istae dies epularum atque laetitiae, et mitterent sibi invicem ciborum partes et pauperibus munuscula largirentur.
ESTH|9|23|Susceperuntque Iudaei in sollemnem ritum cuncta, quae eo tempore facere coeperant, et quae Mardochaeus litteris facienda mandaverat.
ESTH|9|24|Aman enim filius Amadathi stirpis Agag, adversarius omnium Iudaeorum, cogitavit contra eos malum, ut deleret illos, et misit Phur, id est sortem, ut eos conturbaret atque deleret.
ESTH|9|25|Sed postquam ingressa est Esther ad regem, mandavit ille simul cum litteris, ut malum, quod iste contra Iudaeos cogitaverat, reverteretur in caput eius, et suspenderentur ipse et filii eius in patibulo.
ESTH|9|26|Atque ex illo tempore dies isti appellati sunt Phurim propter nomen Phur. Propter cuncta illa, quae in hac epistula continentur,
ESTH|9|27|et propter ea, quae de his viderant et quae eis acciderant, statuerunt et in sollemnem ritum numquam mutandum susceperunt Iudaei super se et semen suum et super cunctos, qui religioni eorum voluerint copulari, ut duos hos dies secundum praeceptum et tempus eorum singulis annis celebrarent.
ESTH|9|28|Isti dies memorarentur et celebrarentur per singulas generationes in singulis cognationibus, provinciis et civitatibus, nec esset ulla civitas, in qua dies Phurim non observarentur a Iudaeis et ab eorum progenie.
ESTH|9|29|Scripseruntque Esther regina filia Abihail et Mardochaeus Iudaeus omni studio ad confirmandam hanc secundam epistulam Phurim.
ESTH|9|30|Et miserunt ad omnes Iudaeos, qui in centum viginti septem provinciis regis Asueri versabantur, verba pacis et veritatis,
ESTH|9|31|statuentes dies Phurim pro temporibus suis, sicut constituerant Mardochaeus et Esther, et sicut illi statuerant pro seipsis et pro semine suo, praecepta ieiuniorum et clamorum.
ESTH|9|32|Et mandatum Esther confirmavit praecepta Phurim et scriptum est in libro.
ESTH|10|1|Rex vero Asuerus terrae et maris insulis imposuit tribu tum.
ESTH|10|2|Cuius fortitudo et imperium et dignitas atque sublimitas, qua exaltavit Mardochaeum, scripta sunt in libro annalium regum Medorum atque Persarum,
ESTH|10|3|et quomodo Mardochaeus Iudaici generis secundus a rege Asuero fuerit et magnus apud Iudaeos et acceptabilis plebi fratrum suorum, quaerens bona populo suo et loquens ea, quae ad pacem seminis sui pertinerent.
