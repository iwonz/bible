EZEK|1|1|І сталося тридцятого року, четвертого місяця, п'ятого дня місяця, коли я був серед полонених над річкою Кевар, відкрилося небо, і побачив я Божі видіння.
EZEK|1|2|П'ятого дня місяця, це п'ятий рік полону царя Єгоякима,
EZEK|1|3|сталося Господнє слово до Єзекіїля, сина Бузі, священика, у халдейському краї над річкою Кевар, і була там над ним Господня рука.
EZEK|1|4|І побачив я, аж ось бурхливий вітер насував із півночі, велика хмара та палючий огонь; а навколо неї сяйво, а з середини його ніби блискуча мідь, з-посеред огню.
EZEK|1|5|А з середини його подоба чотирьох живих істот, а оце їхній вид: вони мали подобу людини.
EZEK|1|6|І кожна мала чотири обличчі, і кожна з них мала чотири крилі.
EZEK|1|7|А їхня нога нога проста, а стопа їхньої ноги як стопа телячої ноги, і вони сяяли, як ніби блискуча мідь.
EZEK|1|8|А під їхніми крилами були людські руки на чотирьох сторонах їхніх, і вони четверо мали свої обличчя та свої крила.
EZEK|1|9|Їхні крила прилягали одне до одного, не оберталися в ході своїй, кожне ходило просто наперед себе.
EZEK|1|10|А подоба їхнього обличчя обличчя людини та обличчя лева мали вони четверо з правиці, а обличчя вола мали вони четверо з лівиці, і обличчя орла мали вони четверо.
EZEK|1|11|А їхні обличчя та їхні крила були розділені вгорі; у кожного двоє крил злучувалися одне з одним, і двоє закривали їхнє тіло.
EZEK|1|12|І кожна ходила просто перед себе. Туди, куди бажав дух ходити, вони йшли, не оберталися в ході своїй.
EZEK|1|13|А подоба тих істот була на вид вугілля з огню, вони палали на вигляд смолоскипів; той огонь проходжувався поміж істотами. І огонь мав сяйво, і з огню виходила блискавка.
EZEK|1|14|І ті живі істоти бігали й верталися, немов блискавка.
EZEK|1|15|І придивився я до тих істот, аж ось по одному колесі на землі при тих живих істотах, при чотирьох їхніх обличчях.
EZEK|1|16|Вид тих колес та їхній виріб як вигляд хризоліту, й одна подоба їм чотирьом, а їхній вид та їхній виріб ніби колесо в колесі.
EZEK|1|17|Вони ходили в ході своїй на чотири боки, не оберталися в ході своїй.
EZEK|1|18|А їхні обіддя були високі та страшні; і їхнє обіддя довкола в чотирьох їх було повне очей.
EZEK|1|19|І коли ходили ті живі істоти, ходили й ті колеса при них; а коли ті істоти підіймалися з-над землі, підіймалися й ті колеса.
EZEK|1|20|Куди бажав дух ходити, ішли, куди мав той дух іти; і ті колеса підіймалися з ними, бо в колесах був дух істот.
EZEK|1|21|Коли ті йшли, ходили й вони; а коли ті стояли стояли й вони; а коли ті підіймалися з-над землі, підіймалися з ними й ті колеса, бо був дух істот у тих колесах.
EZEK|1|22|А на головах тих живих істот була подоба небозводу, ніби грізний кришталь, розтягнений над їхніми головами згори.
EZEK|1|23|А під цим небозводом були їхні прості крила, звернені одне до одного. У кожної було по двоє крил, що закривали їм їхні тіла.
EZEK|1|24|А коли вони йшли, чув я шум їхніх крил, як шум великої води, як голос Всемогутнього, звук гамору, як табору. А коли вони ставали, опадали їхні крила.
EZEK|1|25|І розлягався голос з-над небозводу, що над їхньою головою. І коли вони ставали, опадали їхні крила.
EZEK|1|26|А згори небозводу, що над їхньою головою, була подоба трону на вигляд каменя сапфіру; а на подобі трону була подоба на вигляд людини, на ньому згори.
EZEK|1|27|І бачив я ніби блискучу мідь, на вид огню в середині його навколо, від виду стегон його й вище, а від виду стегон його й до долу бачив я ніби огонь та сяйво навколо нього.
EZEK|1|28|Як вигляд веселки, що буває в хмарі в дощовий день, такий був вигляд сяйва навколо. Це був вигляд подоби Господньої слави! І коли я це побачив, я впав на обличчя своє, і почув голос, що говорив.
EZEK|2|1|І сказав Він до мене: Сину людський, зведися на ноги свої, і Я буду говорити з тобою!
EZEK|2|2|І ввійшов в мене дух, коли Він говорив до мене, і звів мене на мої ноги, і я чув Того, Хто говорив до мене.
EZEK|2|3|І сказав Він до мене: Сину людський, Я посилаю тебе до Ізраїлевих синів, до людей бунтівників, що бунтуються проти Мене. Вони та їхні батьки відпали від Мене аж до цього дня!
EZEK|2|4|А ці сини, що Я посилаю тебе до них, зухвалого обличчя та твердого серця. І ти скажеш до них: Так говорить Господь Бог!
EZEK|2|5|А вони чи послухаються, чи занехають, бо вони дім ворохобний, то пізнають, що пророк був серед них.
EZEK|2|6|А ти, сину людський, не бійся їх, і не бійся їхніх слів, хоч вони для тебе будяччя та тернина, і ти сидиш між скорпіонами. Слів їхніх не бійся, а їхнього вигляду не лякайся, бо вони дім ворохобний.
EZEK|2|7|І будеш говорити до них Мої слова, чи вони послухаються, чи занехають, бо вони ворохобні.
EZEK|2|8|А ти, сину людський, послухай, що кажу Я тобі: Не будь ворохобний, як цей дім ворохобности, відкрий свої уста та з'їж, що Я тобі дам.
EZEK|2|9|І побачив я, аж ось до мене простягнена рука, а в ній звій книжковий.
EZEK|2|10|І Він розгорнув його перед моїм обличчям, а він пописаний спереду та ззаду. І було на ньому написано пісні плачу, стогін та горе...
EZEK|3|1|І сказав Він до мене: Сину людський, з'їж, що знайдеш! З'їж цього звоя, і йди, говори до Ізраїлевого дому!
EZEK|3|2|І відкрив я свої уста, і Він дав мені з'їсти цього звоя.
EZEK|3|3|І сказав Він до мене: Сину людський, нагодуй свого живота, і наповни своє нутро тим звоєм, що даю Я тобі! І я з'їв. І був він в устах моїх солодкий, як мед.
EZEK|3|4|І сказав Він до мені: Сину людський, іди, ввійди до Ізраїлевого дому, і говори до них Моїми словами.
EZEK|3|5|Бо ти посланий не до народу чужої мови та тяжкого язика, але до Ізраїлевого дому,
EZEK|3|6|не до численних народів чужої мови та тяжкого язика, що ти не розумієш їхніх слів. Та коли б і до них послав тебе, вони будуть слухати тебе!
EZEK|3|7|Але Ізраїлів дім не захоче слухатися тебе, бо вони не хочуть слухатися Мене, бо ввесь Ізраїлів дім твердолобі та жорстокосерді вони!
EZEK|3|8|Ось Я зробив твоє обличчя твердим проти їхнього обличчя, і чоло твоє твердим проти лоба їхнього.
EZEK|3|9|Як той діямант, твердішим від скелі, зробив Я чоло твоє, не бійся їх, і не лякайся перед ними, бо вони дім ворохобности!
EZEK|3|10|І сказав Він до мене: Сину людський, усі Мої слова, які говорю Я до тебе, візьми в своє серце та слухай вухами своїми.
EZEK|3|11|І йди, піди до вигнанців, до синів твого народу, і будеш говорити до них і скажеш їм: Так говорить Господь Бог, а вони чи послухаються, чи занехають.
EZEK|3|12|І підійняв мене Дух, і я почув за собою гуркіт громового голосу: Благословенна слава Господня! із свого місця,
EZEK|3|13|і шум крил живих істот, що дотикались одне об одне, і цокіт коліс рівночасно з ними, і гуркіт громового голосу!...
EZEK|3|14|І Дух підійняв мене, і взяв мене, і йшов я огірчений в лютості духа свого, а Господня рука була надо мною сильна!
EZEK|3|15|І прийшов я до вигнанців в Тел-Авіві, що сидять при річці Кевар, і там, де вони сидять, сидів і я там серед них сім день остовпілий.
EZEK|3|16|І сталося в кінці семи день, і було слово Господнє до мене таке:
EZEK|3|17|Сину людський, Я настановив тебе вартовим для Ізраїлевого дому, і як почуєш ти слово з уст Моїх, то остережи їх від Мене.
EZEK|3|18|Коли Я скажу безбожному: Конче помреш, а ти не остережеш його й не будеш говорити, щоб остерегти несправедливого від його несправедливої дороги, щоб він жив, то цей безбожний помре за свою провину, а його кров Я зажадаю з твоєї руки!
EZEK|3|19|Але ти, коли остережеш несправедливого, а він не вернеться від своєї несправедливости та від своєї несправедливої дороги, він помре за свою провину, а ти душу свою врятував.
EZEK|3|20|А коли праведний відвернеться від своєї справедливости та зробить кривду, то я покладу спотикання перед ним, і він помре, бо ти не остеріг його. Він за гріх свій помре, і не згадаються його праведні вчинки, які він робив, і кров його з твоєї руки Я буду жадати!
EZEK|3|21|А ти, коли остережеш справедливого, щоб справедливий не грішив, і він не згрішив, то жити буде він жити, бо був остережений, а ти душу свою врятував.
EZEK|3|22|І була там надо мною Господня рука, і сказав Він до мене: Устань, вийди до долини, і там Я буду говорити з тобою.
EZEK|3|23|І встав я, і вийшов до долини, аж ось там стояла слава Господня, як та слава, яку я бачив над річкою Кевар. І впав я на обличчя своє...
EZEK|3|24|Та ввійшов у мене Дух, і звів мене на ноги мої. І Він говорив зо мною й сказав мені: Увійди, замкнися в середині свого дому!
EZEK|3|25|А ти, сину людський, ось дадуть на тебе шнури, і зв'яжуть тебе ними, і ти не вийдеш з-поміж них!
EZEK|3|26|А язик твій приліплю до твого піднебіння, і ти занімієш, і не будеш їм більш докоряти, бо вони дім ворохобний.
EZEK|3|27|А коли Я говоритиму з тобою, то відкрию твої уста, і ти скажеш до них: Так говорить Господь Бог. Хто хоче слухати нехай слухає, а хто хоче занехати нехай занехає, бо вони дім ворохобний!
EZEK|4|1|А ти, сину людський, візьми собі цеглину, і поклади її перед собою, і накреслиш на ній місто Єрусалим.
EZEK|4|2|І постав проти нього облогу, і збудуй проти нього башту, і висип вала навколо нього, і постав проти нього табори війська, і постав проти нього муроломи.
EZEK|4|3|І візьми собі залізну сковороду, і постав її ніби залізною стіною поміж собою та між тим містом, і зверни своє обличчя до нього, і буде воно в облозі, і ти обляжеш його. Це ознака для Ізраїлевого дому!
EZEK|4|4|А ти лягай на лівий свій бік, і поклади на нього провину Ізраїлевого дому. За числом днів, що будеш лежати на ньому, ти будеш носити їхню провину.
EZEK|4|5|І Я призначив тобі роки їхньої провини за числом днів, три сотні й дев'ятдесят днів, і ти будеш носити провину Ізраїлевого дому.
EZEK|4|6|А коли ти це скінчиш, то ляжеш удруге, на правий свій бік, і будеш носити провину Юдиного дому сорок день, один день за один рік Я тобі призначив.
EZEK|4|7|І на облогу Єрусалиму зверни своє обличчя та відкрите рамено своє, і будеш пророкувати на нього.
EZEK|4|8|І ось Я накладу на тебе шнури, і ти не повернешся з боку одного на інший бік, аж поки ти не закінчиш днів своєї облоги.
EZEK|4|9|А ти візьми собі пшениці та ячменю, і бобів та сочевиці, і проса та вики, і даси їх до одного посуду, і зробиш із них собі хліб, за кількістю днів, що лежатимеш на боці своєму, три сотні й дев'ятдесят день будеш те їсти.
EZEK|4|10|А їжа твоя, яку будеш ти їсти, буде вагою двадцять шеклів на день, час від часу будеш це їсти.
EZEK|4|11|І воду будеш пити мірою, шоста частина гіна, час від часу будеш пити.
EZEK|4|12|І їстимеш це, як ячмінного калача, і будеш пекти це на кавалках людського калу, перед їхніми очима...
EZEK|4|13|І сказав Господь: Так будуть їсти Ізраїлеві сини свій нечистий хліб серед тих народів, куди Я їх вижену...
EZEK|4|14|А я відказав: О Господи, Боже, ось душа моя не занечищена, і падла та розшматованого звірями я не їв від молодости своєї й аж дотепер, і м'ясо нечисте не входило в мої уста.
EZEK|4|15|І сказав Він до мене: Дивися, Я дав тобі товарячий гній замість людського калу, і ти зроби на ньому свій хліб!
EZEK|4|16|І сказав Він до мене: Сину людський, ось Я поламаю підпору хліба в Єрусалимі, і будуть їсти хліб за вагою та в страху, а воду будуть пити за мірою та зо смутком,
EZEK|4|17|щоб відчули вони брак хліба та води, і жахнулися один з одним, і вони знидіють за свій гріх!
EZEK|5|1|А ти, сину людський, візьми собі гострого меча, як бритву стрижіїв; візьми його собі, і проведи ним по голові своїй та по бороді своїй. І візьми собі вагові шальки, і поділи те волосся.
EZEK|5|2|Третину спали в огні посеред міста, коли виповняться дні облоги; і візьми другу третину, і посічи мечем навколо нього, а третину розпороши на вітер, і Я витягну меча за ними.
EZEK|5|3|І візьми звідти мале число волосся, і зав'яжи його в своїх полах.
EZEK|5|4|І візьми із нього ще, і кинь його до середини огню, і спали його в огні, з нього вийде огонь на ввесь Ізраїлів дім...
EZEK|5|5|Так говорить Господь Бог: Цей Єрусалим Я поставив його в середині народів, а довкілля його країни.
EZEK|5|6|Та він став проти постанов Моїх більше від поганів, а проти устав Моїх більше від тих країн, що навколо нього, бо права Мої вони відкинули, а устави Мої не ходили вони ними.
EZEK|5|7|Тому так говорить Господь Бог: За те, що ви ворохобилися більше від тих поган, що навколо вас, й уставами Моїми не ходили, і постанов Моїх не виконували, а робили за постановами тих поган, що навколо вас,
EZEK|5|8|тому так говорить Господь Бог: Ось Я проти тебе, Сам Я, і зроблю серед тебе суди перед очима тих поган!
EZEK|5|9|І зроблю на тобі те, чого Я не робив, і нічого подібного вже не зроблю, за гидоти твої.
EZEK|5|10|Тому серед тебе батьки будуть їсти синів, а сини будуть їсти батьків своїх, і виконаю над тобою присуди, і розпорошу ввесь останок твій на всі вітри!...
EZEK|5|11|Тому, як живий Я, говорить Господь Бог, за те, що ти занечистив святиню Мою всіма гидотами своїми та всіма обридженнями своїми, то теж Я відкину тебе, й око Моє не матиме милосердя, і Сам Я не змилосерджуся!
EZEK|5|12|Третина твоя помре від моровиці й загине від голоду серед тебе, а третина попадає від меча в твоїх околицях, а третину розпорошу на всі вітри, і витягну за ними меча!
EZEK|5|13|І докінчиться гнів Мій, і Я заспокою Свою лють проти них, і задовольнюся. І пізнають вони, що Я, Господь, говорив у горливості Своїй, коли доконаю Свою лютість на них!
EZEK|5|14|І зроблю тебе руїною та ганьбою серед людів, що навколо тебе, перед очима кожного, хто буде проходити...
EZEK|5|15|І станеш ганьбою та посміховиськом, осторогою та остовпінням для народів, що навколо тебе, коли буду виконувати на тобі присуди гнівом та люттю, та лютими картаннями. Я, Господь, оце говорив!
EZEK|5|16|Коли Я пошлю на них злі стріли голоду, що будуть нищівними, що пошлю їх понищити вас та примножу голод на вас, то Я зламаю вам підпору хліба,
EZEK|5|17|і пошлю на вас голод та злу звірину, і позбавлю тебе дітей, і моровиця та кров перейде серед тебе, і спроваджу на тебе меча. Я, Господь, оце говорив!
EZEK|6|1|І було мені слово Господнє таке:
EZEK|6|2|Сину людський, зверни своє обличчя до Ізраїлевих гір, і пророкуй на них,
EZEK|6|3|та й скажеш: Гори Ізраїлеві, послухайте слова Господа Бога! Так говорить Господь Бог горам та підгіркам, і річищам та долинам: Ось Я спроваджу на вас меча, і вигублю ваші пагірки,
EZEK|6|4|і будуть опустошені ваші жертівники, і будуть розбиті ваші фіґури сонця, і кину Я ваших побитих перед вашими божками!
EZEK|6|5|І дам трупи Ізраїлевих синів перед їхніми божками, і розпорошу ваші кості навколо ваших жертівників...
EZEK|6|6|По всіх місцях вашого перебування міста будуть поруйновані, а пагірки попустошені, щоб ваші жертівники були поруйновані та побезчещені, і щоб були розтрощені й перестали існувати ваші божки, і були розбиті ваші фіґури сонця, і були стерті ваші діла...
EZEK|6|7|І впаде забитий між вами, і ви пізнаєте, що Я Господь!
EZEK|6|8|А Я позоставлю з вас решту, бо будете мати врятованих від меча серед народів, коли ви будете розпорошені серед країн.
EZEK|6|9|І ваші врятовані згадають про Мене серед народів, куди будуть забрані до полону, коли Я зламаю їхнє блудне серце, що відпало від Мене, та їхні очі, що перелюб чинили з своїми божками, і вони самі будуть бридитися тих злих речей, що робили, щодо всіх їхніх гидот.
EZEK|6|10|І пізнають вони, що Я Господь, і що Я не надармо говорив, що вчиню їм оцю злу річ!
EZEK|6|11|Так говорить Господь Бог: Удар своєю долонею й тупни ногою своєю, і скажи: Горе за всі злі вчинки Ізраїлевого дому, за які вони попадають від меча, голоду та моровиці!
EZEK|6|12|Той, хто далекий, помре від моровиці, а хто близький впаде від меча, а хто позостане та буде врятований помре від голоду. І так Я викінчу Свою лютість на них!
EZEK|6|13|І пізнаєте ви, що Я Господь, коли їхні забиті будуть лежати серед їхніх божків навколо їхніх жертівників на всякім високім підгір'ї, на всіх щитах гір, і під усяким зеленим деревом, і під усяким густим дубом, на місці, де вони приносили приємні пахощі для всіх своїх божків.
EZEK|6|14|І Я витягну руку Свою на них, і зроблю цей Край спустошенням та пусткою, від пустині аж до Рівли, по всіх місцях їхнього сидіння... І пізнають вони, що Я Господь!
EZEK|7|1|І було мені слово Господнє таке:
EZEK|7|2|А ти, сину людський, послухай: Отак Господь Бог промовляє до Краю Ізраїлевого: Кінець, надійшов той кінець на чотири окрайки землі!
EZEK|7|3|На тебе тепер цей кінець, і пошлю Я на тебе Свій гнів, і тебе розсуджу за твоїми дорогами, і на тебе складу всі гидоти твої.
EZEK|7|4|І око Моє над тобою не змилується, і милосердя не буду Я мати, бо дороги твої Я на тебе складу, а гидоти твої серед тебе зостануть, і пізнаєте ви, що Я то Господь!
EZEK|7|5|Отак Господь Бог промовляє: Ось приходить біда на біду!
EZEK|7|6|Приходить кінець, приходить кінець, він збудився на тебе, приходить ось він!
EZEK|7|7|Надійшла твоя доля для тебе, о мешканче Краю, приходить цей час, близький той день заколоту, нема на горах крику радости...
EZEK|7|8|Тепер лютість Свою незабаром Я виллю на тебе, і Свій гнів докінчу проти тебе, і тебе осуджу за твоїми дорогами, і на тебе складу всі гидоти твої!
EZEK|7|9|І око Моє над тобою не змилується, і милосердя не буду Я мати, бо дороги твої Я на тебе складу, а гидоти твої серед тебе залишаться, і пізнаєте ви, що Я Господь, що карає!
EZEK|7|10|Ось той день, ось приходить, доля виходить, виростає кий, розцвітає пиха,
EZEK|7|11|розвилося насильство для кия безбожности! Нічого із них не залишиться: ані з численности їхньої, ані з їхнього заворушення, ані з їхньої пишноти...
EZEK|7|12|Надходить той час, наближається день... Хто купує, нехай не радіє, а хто продає, хай не буде в жалобі, бо сунеться лютість на все многолюддя його!
EZEK|7|13|Бо до проданого не повернеться вже продавець, хоча б залишився при житті між живими, бо пророцтво про все многолюддя їхнє не відміниться, і ніхто беззаконням своїм не зміцнить свого життя...
EZEK|7|14|Засурмлять у сурму та все приготують, та не піде ніхто на війну, бо на все многолюддя його Моя лютість!
EZEK|7|15|На вулиці меч, моровиця ж та голод у домі, хто на полі помре від меча, з хто в місті зжере того голод та мор...
EZEK|7|16|І врятовані з них повтікають, і будуть на горах, немов голуби із долин, всі будуть стогнати, кожен за гріх свій...
EZEK|7|17|Усі руки ослабнуть, затремтять, як вода, всі коліна,
EZEK|7|18|і веретами попідперізуються, і покриє їх страх, і на кожнім лиці буде сором, а на всіх головах їхніх жалобна та лисина...
EZEK|7|19|Вони повикидають на вулицю срібло своє, і за ніщо їхнє золото стане, їхнє срібло та золото їхнє не буде могти врятувати їх у день гніву Господнього, ним не наситять своєї душі й свого нутра вони не наповнять, бо їхня провина була перешкодою!
EZEK|7|20|А гордість вчинили за славну оздобу свою, у ній наробили бовванів гидоти своєї й обриджень своїх, тому їм оберну Я її на нечистість,
EZEK|7|21|і віддам її в руку чужих на грабунок, а нечестивим землі на здобич...
EZEK|7|22|І обличчя Своє відверну Я від них, і вони побезчестять Мій скарб, і ввійдуть до нього насильники та й побезчестять його...
EZEK|7|23|Зроби ланцюга, бо земля переповнилась правом кривавим, а місто насильством наповнилось...
EZEK|7|24|І наведу Я найзліших із народів, і посядуть вони доми їхні, і гордість вельможних спиню, і святощі їхні побезчещені будуть!
EZEK|7|25|Загибіль іде, й вони будуть шукати спокою та не буде його...
EZEK|7|26|Прийде біда до біди, й буде звістка до звістки, і будуть шукати пророцтва в пророка, та згине Закон у священиків і рада у старших...
EZEK|7|27|Цар буде в жалобі, і страхом зодягнеться князь, а руки народу землі затремтять... За дорогами їхніми їм учиню, і судитиму їх їхніми судами, і пізнають, що Я то Господь!
EZEK|8|1|І сталося за шостого року, шостого місяця, п'ятого дня місяця сидів я в своєму домі, а Юдині старші сиділи передо мною, то впала там на мене рука Господа Бога.
EZEK|8|2|І побачив я, аж ось подоба, на вигляд чоловіка: від виду стегон його й додолу огонь, а від стегон його й догори на вигляд сяйва, ніби палаюча мідь.
EZEK|8|3|І витягнув Він подобу руки, і взяв мене за волосся моєї голови, а Дух підійняв мене між землею та між небом, і впровадив мене до Єрусалиму в Божих видіннях, до входу внутрішньої брами, зверненої на північ, де місце перебування ідола, що викликує заздрість.
EZEK|8|4|І ось була там слава Ізраїлевого Бога, як той вид, що я бачив у долині!
EZEK|8|5|І сказав Він до мене: Сину людський, зведи очі свої в напрямі на північ! І звів я очі свої в напрямі на північ, аж ось з півночі, від брами жертівника, був той ідол заздрости при вході.
EZEK|8|6|І сказав Він до мене: Сину людський, чи ти бачиш, що вони роблять! Це великі гидоти, що Ізраїлів дім робить тут, щоб віддалитися від Моєї святині! Та ти знову побачиш іще більші гидоти.
EZEK|8|7|І привів мене до входу подвір'я, і побачив я, аж ось дірка в стіні!
EZEK|8|8|І сказав Він мені: Сину людський, прокопай дірку в стіні! І прокопав я в стіні, аж ось вхід!
EZEK|8|9|І сказав Він до мене: Увійди, і побач ті злі гидоти, які вони роблять отут!
EZEK|8|10|І ввійшов я й побачив, аж ось усякий вид плазуна та огидливої звірини, і всякі божки Ізраїлевого дому, накреслені на стіні навколо кругом...
EZEK|8|11|А сімдесят чоловіка зо старших Ізраїлевого дому та Яазанія, Шафанів син, що стояв посеред них, стояли перед ними, і кожен мав у своїй руці свою кадильницю, і підіймалися пахощі з хмари кадила.
EZEK|8|12|І сказав Він до мене: Чи бачив ти, сину людський, що роблять Ізраїлеві старші в темноті, кожен у кімнатах своїх ідолів? Бо говорять вони: Господь нас не бачить, Господь покинув цей Край...
EZEK|8|13|І сказав Він до мене: Ти знову побачиш ще більші гидоти, які вони роблять.
EZEK|8|14|І Він запровадив мене до входу до брами Господнього дому що на півночі, аж ось там сидять жінки, що оплакували Таммуза.
EZEK|8|15|І сказав Він до мене: Чи ти бачив, сину людський? Ти знову побачиш гидоти ще більші від цих!
EZEK|8|16|І Він запровадив мене до внутрішнього подвір'я Господнього дому. Аж ось при вході до Господнього храму, між притвором та між жертівником, було біля двадцяти й п'яти чоловіка: спини їхні до Господнього храму, а їхні обличчя на схід, і вони кланялися до сходу, до сонця.
EZEK|8|17|І сказав Він до мене: Чи ти бачив, сину людський? Чи легко Юдиному дому, щоб не робити тих гидот, які вони роблять отут? Бо вони наповнили Край насильством, і знову гнівають Мене, й ось вони держать зелені галузки при носі своїм.
EZEK|8|18|Тому то й Я зроблю з лютістю: око Моє не змилується, і милосердя не буду Я мати. І вони будуть кликати сильним голосом в вуха Мої, та Я їх не почую!...
EZEK|9|1|І кликнув Він в уші мої сильним голосом, кажучи: Наблизьте карателів міста, і кожен нехай має в своїй руці свої нищівні знаряддя.
EZEK|9|2|І ось прийшли шість чоловіка з дороги горішньої брами, що звернена на північ, і кожен мав у своїй руці свої знаряддя розбивання, а серед них один чоловік був одягнений в льняне, а писарський каламар був при стегнах його. І вони прийшли, і стали при мідяному жертівнику.
EZEK|9|3|А слава Ізраїлевого Бога піднялася з-над Херувима, що була над ним, до порога дому. І закликав Він чоловіка, одягненого в льняне, що писарський каламар був при стегнах його.
EZEK|9|4|І сказав Господь до нього: Перейди серединою міста, серединою Єрусалиму, і зроби знака на чолах людей, що зідхають та стогнуть над усіма тими гидотами, що робляться в його середині.
EZEK|9|5|А до інших Він сказав при мені: Ходіть за ним у місті, і вбивайте; нехай ваше око не має милосердя, і ви не змилуйтеся!
EZEK|9|6|Старого, юнака, і дівчину, і дітей та жінок позабивайте дощенту, а до кожної людини, що на ній цей знак, не підійдете; а зачнете від Моєї святині... І зачали вони від тих старих людей, що були перед домом.
EZEK|9|7|І сказав Він до них: Занечистіть цей дім, і наповніть подвір'я трупами, і вийдіть! І вони повиходили, і вбивали в місті.
EZEK|9|8|І сталося, коли вони вбивали, то я позостався, і впав на своє обличчя, і кликав та казав: О Господи, Боже, чи Ти вигубиш увесь останок Ізраїлів, виливаючи гнів Свій на Єрусалим?
EZEK|9|9|І сказав Він до мене: Провина дому Ізраїля й Юди дуже-дуже велика, і земля наповнена душогубствами, а місто повне кривди. Бо вони кажуть: Господь покинув цей Край, і Господь не бачить...
EZEK|9|10|І також Я, не змилосердиться око Моє, і не змилуюсь Я, їхню дорогу Я дам на їхню голову!
EZEK|9|11|І ось чоловік, одягнений в льняне, що каламар був при стегнах його, приніс відповідь, кажучи: Я зробив, як мені наказав Ти!
EZEK|10|1|І побачив я, аж ось на небозводі, що на голові Херувимів, було щось, як камінь сапфір, на вигляд подоби трону бачилося на них.
EZEK|10|2|І Він промовив до того чоловіка, одягненого в льняне, та й сказав: Увійди поміж колеса під Херувимом, і наповни свої жмені вуглинами огню з-поміж Херувимів, і кинь на місто! І він увійшов перед моїми очима.
EZEK|10|3|А Херувими стояли з правого боку дому, коли входив чоловік, і хмара наповнила внутрішнє подвір'я.
EZEK|10|4|І піднялася слава Господня з-над Херувима на поріг дому, і наповнився дім хмарою, а подвір'я наповнилося сяйвом Господньої слави.
EZEK|10|5|А шум крил Херувимів був чутий аж до зовнішнього подвір'я, як голос Бога Всемогутнього, коли Він говорить.
EZEK|10|6|І сталося, коли Він наказав чоловікові, одягненому в льняне, кажучи: Візьми огонь поміж колесами з-під Херувимів, то той прийшов і став при колесі.
EZEK|10|7|І Херувим простягнув свою руку з-поміж Херувимів до огню, що поміж Херувимами, і взяв, і дав до жмені одягненого в льняне, а той узяв і вийшов.
EZEK|10|8|І показалася в Херувимів подоба людської руки під їхніми крилами.
EZEK|10|9|І я побачив, аж ось чотири колесі при Херувимах, по одному колесі при кожному Херувимі, а вид тих колес, ніби вигляд каменя хризоліта.
EZEK|10|10|А їхній вигляд подоба одна чотирьом їм, як коли б колесо було в колесі.
EZEK|10|11|В ході своїй вони йшли на чотири свої боки, не оберталися в ході своїй, бо до того місця, куди обернеться голова, за нею йшли вони, не оберталися в ході своїй.
EZEK|10|12|А все їхнє тіло, і їхня спина, і їхні руки, і їхні крила, і ті колеса були повні очей навколо, всі чотири мали колеса.
EZEK|10|13|А ці колеса були кликані при мені Ґалґал.
EZEK|10|14|А в кожного чотири обличчі: обличчя одного обличчя Херувима, обличчя другого обличчя людини, а третій обличчя лева, а четвертий обличчя орла.
EZEK|10|15|І піднялися ті Херувими. Це та жива істота, яку я бачив на річці Кевар.
EZEK|10|16|А коли йшли ті Херувими, то йшли й ті колеса при них, а коли ті Херувими підіймають свої крила, щоб знятись із землі, не відвертаються також ті колеса від них.
EZEK|10|17|Коли ті ставали, ставали й вони, а коли ті підіймалися, підіймалися й вони, бо в них був дух живої істоти.
EZEK|10|18|І вийшла слава Господня з-над порога дому, і стала над Херувимами.
EZEK|10|19|І підняли Херувими свої крила, і знялися з землі на моїх очах, коли вони йшли, а ті колеса побіч них, і стали при вході до східньої брами Господнього дому, а слава Ізраїлевого Бога зверху над ними.
EZEK|10|20|Це та жива істота, яку я бачив під Богом Ізраїлевим над річкою Кевар. І я пізнав, що це Херувими.
EZEK|10|21|У кожного було по чотири обличчі, у кожного чотири крилі, а під їхніми крилами подоба людських рук.
EZEK|10|22|А подоба їхнього обличчя це ті обличчя, які я бачив над річкою Кевар, їхній вигляд та вони самі. Кожен ішов просто вперед.
EZEK|11|1|І підійняв мене Дух, і привів мене до східньої брами Господнього дому, що обернена на схід. І ось при вході до брам двадцять і п'ять чоловіка, а серед них бачив я Яазанію, сина Аззурового, та Пелатію, сина Бенаїного, князів народу.
EZEK|11|2|І сказав Він до мене: Сину людський, оце ті люди, що задумують кривду, і радять злу раду в цьому місті,
EZEK|11|3|що говорять: Не скоро будувати доми. Воно казан, а ми м'ясо.
EZEK|11|4|Тому пророкуй на них, пророкуй, сину людський!
EZEK|11|5|І зійшов на мене Дух Господній, та й до мене сказав: Скажи: Так говорить Господь: Отак кажете, доме Ізраїлів, і заміри вашого духа Я знаю їх.
EZEK|11|6|Ви намножили своїх забитих у цьому місті, і наповнили його вулиці трупами.
EZEK|11|7|Тому так говорить Господь Бог: Ваші забиті, що ви їх поклали серед нього, вони те м'ясо, а воно той казан. Та Я випроваджу вас із нього!
EZEK|11|8|Ви боїтеся меча і меча наведу Я на вас, говорить Господь Бог.
EZEK|11|9|І випроваджу вас із нього, і дам вас у руку чужих, і зроблю між вами присуди!
EZEK|11|10|Від меча ви попадаєте; на границі Ізраїля розсуджу вас, і ви пізнаєте, що Я то Господь!
EZEK|11|11|Воно не буде вам казаном, і ви не станете в ньому м'ясом. При границі Ізраїля розсуджу вас!
EZEK|11|12|І пізнаєте ви, що Я Господь, бо за уставами Його ви не ходили, а постанов Моїх не виконували, але виконували за постановами тих народів, що навколо вас.
EZEK|11|13|І сталося, коли я пророкував, то Пелатія, син Бенаніїн, помер. І впав я на своє обличчя, і закричав сильним голосом та й сказав: О Господи Боже, Ти робиш кінець з Ізраїлевим останком!...
EZEK|11|14|І було мені слово Господнє таке:
EZEK|11|15|Сину людський, брати твої, брати твої мужі рідні тобі, а ввесь Ізраїлів дім увесь той, що до них говорили мешканці Єрусалиму: Віддаліться від Господа, нам даний цей Край на володіння,
EZEK|11|16|тому скажи: Так говорить Господь Бог: Хоч Я віддалив їх поміж народи, і хоч розпорошив їх по краях, проте буду для них хоч малою святинею в тих краях, куди вони ввійшли.
EZEK|11|17|Тому скажи: Так говорить Господь Бог: І позбираю Я вас із народів, зберу з тих країв, серед яких ви розпорошені, і дам вам Ізраїлеву землю.
EZEK|11|18|І вони ввійдуть туди, і викинуть з неї усі мерзоти її та всі гидоти її.
EZEK|11|19|І дам їм одне серце, і нового духа дам у вас, і вийму з їхнього тіла серце камінне, і дам їм серце із м'яса,
EZEK|11|20|щоб вони ходили за уставами Моїми, і додержували Мої постанови та виконували їх. І вони стануть Мені народом, а Я буду їм Богом!
EZEK|11|21|А щодо тих, що їхнє серце ходить за гидотами своїми та мерзотами своїми, то поверну їхню дорогу на їхню голову, говорить Господь Бог...
EZEK|11|22|І попідіймали Херувими крила свої, а колеса при них, і слава Ізраїлевого Бога зверху над ними.
EZEK|11|23|І піднялася слава Господня з-над середини міста, і стала на горі, що зо сходу міста.
EZEK|11|24|І дух підніс мене, і ввів мене в Халдею до полонян у видінні, Духом Божим. І підійнялося від мене те видіння, яке я бачив.
EZEK|11|25|І я говорив до полонян усі Господні слова, які Він наказав був мені.
EZEK|12|1|І було мені слово Господнє таке:
EZEK|12|2|Сину людський, ти живеш серед дому ворохобного, вони мають очі, щоб бачити, та не бачать, мають вуха, щоб слухати, та не чують, бо вони дім ворохобний.
EZEK|12|3|А ти, сину людський, пороби собі речі для мандрівки, і йди на вигнання вдень на їхніх очах, і підеш на вигнання з свого місця до іншого місця на їхніх очах, може побачать вони, що вони дім ворохобности.
EZEK|12|4|І повиносиш свої речі, як речі для мандрівки, удень на їхніх очах, а ти вийдеш увечорі на їхніх очах, як виходять вигнанці.
EZEK|12|5|На їхніх очах пробий собі дірку в стіні, і повиносиш нею.
EZEK|12|6|На їхніх очах на рамені повиносиш, винесеш потемки, закриєш обличчя своє, і не побачиш землі, бо Я поставив тебе знаком для Ізраїлевого дому.
EZEK|12|7|І зробив я так, як наказано мені: речі свої я повиносив удень, а ввечорі пробив собі рукою дірку в стіні, потемки повиносив, на рамені носив на їхніх очах.
EZEK|12|8|А ранком було мені слово Господнє таке:
EZEK|12|9|Сину людський, чи ж не сказав до тебе дім Ізраїлів, дім ворохобности: Що ти робиш?
EZEK|12|10|Скажи до них: Так сказав Господь Бог: Це пророцтво про начальника Єрусалиму та ввесь Ізраїлів дім, що в ньому вони.
EZEK|12|11|Скажи: Я ваш знак. Як зробив Я, так буде зроблено їм, підуть на вигнання в полон!
EZEK|12|12|А той начальник, що серед них, на рамені буде нести потемки й вийде; у стіні проб'ють дірку, щоб вивести його; обличчя своє він закриє, щоб не бачити землі очима.
EZEK|12|13|І розтягну на нього сітку Свою, і він буде схоплений в пастку Мою, і відведу його до Вавилону, до халдейського краю, та його він не побачить, і там помре.
EZEK|12|14|А все, що навколо нього, його помічники та всі війська його, розпорошу на всі вітри, і витягну за ними меча...
EZEK|12|15|І пізнають вони, що Я Господь, коли розвію їх поміж народами та розпорошу їх по країнах!
EZEK|12|16|А нечисленних з них людей збережу від меча, від голоду та від зарази, щоб вони оповідали про свої гидоти серед народів, куди поприходять. І вони пізнають, що Я Господь!
EZEK|12|17|І було мені слово Господнє таке:
EZEK|12|18|Сину людський, їж свій хліб у дрижанні, а воду свою пий у тремтінні та в журбі.
EZEK|12|19|І скажеш до народу цього Краю: Так говорить Господь Бог на мешканців Єрусалиму, на Ізраїлеву землю: Вони хліб свій в журбі будуть їсти, а воду свою будуть пити в остовпінні, бо спустошів їхній Край від своєї повні за насилля всіх, що мешкають у ньому.
EZEK|12|20|І поруйнуються населені міста, а Край стане спустошенням, і пізнаєте ви, що Я Господь!
EZEK|12|21|І було мені слово Господнє таке:
EZEK|12|22|Сину людський, що це в вас за приповістка така в Ізраїлевій землі: Продовжаться дні, і зникне всіляке видіння?
EZEK|12|23|Тому скажи їм: Так говорить Господь Бог: Припиню Я цю приповістку, і більше не будуть її приповісткувати в Ізраїлі, але говори їм: Наблизилися оті дні й слово всякого видіння.
EZEK|12|24|Бо не буде вже жодного марного видіння та підлесливого чарування в Ізраїлевім домі.
EZEK|12|25|Бо Я, Господь, буду говорити, а яке слово говоритиму, то буде воно здійснене, не відтягнеться вже, бо за ваших днів, доме ворохобности, буду говорити слово, і його виконаю, говорить Господь Бог.
EZEK|12|26|І було мені слово Господнє таке:
EZEK|12|27|Сину людський, ось говорить Ізраїлів дім: Те видіння, яке він бачить, воно про далекі дні, і про далекі часи він пророкує.
EZEK|12|28|Тому їм скажи: Так говорить Господь Бог: Не відтягнуться вже всі слова Мої, яке слово говоритиму, те буде виконане, говорить Господь Бог!
EZEK|13|1|І було мені слово Господнє таке:
EZEK|13|2|Сину людський, пророкуй на Ізраїлевих пророків, що пророкують, і скажи пророкам, що провіщають із власного серця: Послухайте Господнього слова!
EZEK|13|3|Так говорить Господь Бог: Горе на пророків безумних, що ходять за своїм духом та за тим, чого не бачили!
EZEK|13|4|Твої пророки, Ізраїлю, як ті лисиці в руїнах!
EZEK|13|5|Не ввійшли ви в проломи, і не загородили загороди над Ізраїлевим домом, щоб стати на бій Господнього дня.
EZEK|13|6|Вони бачать марноту та фальшиве чарування, говорячи: Говорить Господь, а Господь не посилав їх, та вони мають надію, що сповниться слово.
EZEK|13|7|Хіба ж не марне видіння ви бачили, і не фальшиве чарування ви говорили? А ви кажете: Говорить Господь, а Я не говорив!
EZEK|13|8|Тому так говорить Господь Бог: За те, що ви говорите марноту, і бачите лжу, тому ось Я проти вас, говорить Господь Бог.
EZEK|13|9|І буде рука Моя проти пророків, що бачать марноту й чарують ілжею. Вони не будуть на раді народу Мого, і в перепису Ізраїлевого дому не будуть записані, і до землі Ізраїлевої не ввійдуть. І пізнаєте ви, що Я Господь Бог!
EZEK|13|10|Саме за те, що вони впровадили народ Мій у помилку, говорячи мир, а миру нема. І він будує мура, а вони тинкують його будьяким тинком.
EZEK|13|11|Скажи до тих, що тинкують будьяким тинком, що мур упаде. Буде дощ заливний, і ви, каміння великого граду, впадете, і вітер бурхливий розвалить мура.
EZEK|13|12|І ось стіна впаде. Чи ж не скажуть вам: Де той тинк, яким ви тинкували?
EZEK|13|13|Тому так говорить Господь Бог: Я вчиню, що бурхливий вітер валитиме в лютості Моїй, і буде дощ заливний в Моїм гніві, і каміння великого граду в лютості на вигублення.
EZEK|13|14|І розіб'ю Я ту стіну, яку ви обтинкували будьяким тинком, і повалю її до землі, й оголиться підвалина її, і впаде, і ви загинете в середині його, Єрусалима, і пізнаєте, що Я Господь!
EZEK|13|15|І докінчу Я лютість Свою на стіні та на тих, що тинкують її якимбудь тинком, і скажу вам: Немає стіни та її тинкувальників,
EZEK|13|16|Ізраїлевих пророків, що пророкували на Єрусалим і бачили для нього видіння миру, та немає миру, говорить Господь!
EZEK|13|17|А ти, сину людський, зверни своє обличчя до дочок свого народу, що пророкують з власного серця, і пророкуй на них,
EZEK|13|18|та й скажи: Так говорить Господь Бог: Горе тим, що шиють чародійні обв'язки на суглоби рук, і роблять хустки на голову всякого зросту, щоб ловити душі. Невже, ловлячи душі Мого народу, ви свої душі спасете?
EZEK|13|19|І ви безчестите Мене в Мого народу за жмені ячменю та за кришки хліба, забиваючи душі, що не повинні б умирати, та лишаючи при житті душі, що не повинні б жити, своїми обманами Моєму народові, що слухають лжу.
EZEK|13|20|Тому так говорить Господь Бог: Ось Я проти ваших чародійних обв'язок, ув які ви ловите душі. І позриваю їх із ваших рамен, і повипускаю ті душі, ті душі, що ви ловите, щоб були вільні, як птахи.
EZEK|13|21|І позриваю ваші хустки, і врятую народ Свій з вашої руки, і не будуть вони вже в вашій руці за здобич, і пізнаєте ви, що Я Господь.
EZEK|13|22|За те, що ви лжею заподіяли біль серцю праведного, хоч Я не зробив йому болю, і за те, що ви зміцнюєте руки безбожного, щоб він не відвернувся від своєї злої дороги, щоб спасти його при житті,
EZEK|13|23|тому більш не будете бачити марноти та не будете віщувати, і Я врятую народ Свій з вашої руки, і ви пізнаєте, що Я Господь!
EZEK|14|1|І прийшли до мене мужі з Ізраїлевих старших, і посідали передо мною.
EZEK|14|2|І було мені слово Господнє таке:
EZEK|14|3|Сину людський, ці мужі допустили своїх божків у своє серце, а спотикання провини своєї поклали перед обличчям своїм. Чи ж можуть вони запитувати Мене?
EZEK|14|4|Тому говори з ними, та й скажеш до них: Так говорить Господь Бог: Кожен чоловік з Ізраїлевого дому, що допустить своїх божків у своє серце, а спотикання провини своєї покладе перед обличчям своїм, і прийде до пророка, тому Я, Господь, відповім, згідно з цим, згідно з многотою його божків,
EZEK|14|5|щоб схопити тих з Ізраїлевого дому за їхнє серце, бо всі вони віддалилися від Мене через своїх божків!
EZEK|14|6|Тому скажи до Ізраїлевого дому: Так говорить Господь Бог: Наверніться, і відступіть від ваших божків, і від усіх ваших гидот відверніть свої обличчя!
EZEK|14|7|Бо кожен чоловік із Ізраїлевого дому або з чужинців, що мешкають серед Ізраїля, коли відступить від Мене, і допустить своїх божків у своє серце, і покладе спотикання своєї провини перед обличчям своїм, і прийде до пророка, щоб запитати Мене, тому Я, Господь, відповім від Себе.
EZEK|14|8|І зверну Я лице Своє проти цього чоловіка, і вчиню його за знака та за приповістку, і вигублю його з-посеред Свого народу, і пізнаєте ви, що Я Господь!
EZEK|14|9|А пророк, коли б був зведений, і говорив би слово, Я, Господь, зведу цього пророка, і простягну руку Свою на нього, і вигублю його з-посеред Свого народу Ізраїлевого!
EZEK|14|10|І понесуть вони свою провину, яка провина того, хто питається, така буде провина пророка,
EZEK|14|11|щоб не блудив уже Ізраїлів дім від Мене, і не занечищувався вже всіма своїми гріхами. І будуть вони Мені народом, а Я буду їм Богом, говорить Господь Бог!
EZEK|14|12|І було мені слово Господнє таке:
EZEK|14|13|Сину людський, коли згрішить проти Мене земля, спроневірюючи, то Я простягну Свою руку на неї, і зламаю їй хлібну підпору, і пошлю на неї голод, і вигублю з неї людину й скотину.
EZEK|14|14|А коли б серед неї були три мужі: Ной, Даниїл та Йов, вони в своїй справедливості врятували б лише свою власну душу, говорить Господь Бог.
EZEK|14|15|Коли б Я перепровадив по землі люту звірину, й обезлюдніла б вона, і стала б вона спустошенням, так що ніхто не проходив би нею через ту звірину,
EZEK|14|16|той й ці три мужі серед неї, як живий Я, говорить Господь Бог, не врятують вони ні синів, ні дочок! Самі вони будуть врятовані, а Край стане спустошенням...
EZEK|14|17|Або коли б Я спровадив на цю землю меча, та й мечеві сказав: Пройди по Краю, і вигуби з нього людину й скотину,
EZEK|14|18|то ці три мужі серед нього, як живий Я! говорить Господь Бог, не врятують синів, ні дочок, бо врятуються самі тільки вони!
EZEK|14|19|Або коли б Я моровицю послав до цієї землі, і вилив би на неї свою лютість у крові, щоб вигубити з неї людину й скотину,
EZEK|14|20|а Ной, Даниїл та Йов були б серед неї, як живий Я! говорить Господь Бог, ані сина, ані дочки не врятували б вони! Вони в своїй справедливості врятують тільки свою власну душу.
EZEK|14|21|Бо так говорить Господь Бог: Хоч послав би Я на Єрусалим чотири Свої лихі присуди: меча, і голод, і люту звірину та моровицю, щоб вигубити з нього людину та скотину,
EZEK|14|22|то все таки залишаться в ньому рештки, що будуть випроваджені, сини та дочки. Ось вони вийдуть до вас, і ви побачите їхню дорогу та їхні вчинки, і будете потішені за те лихо, що Я навів на Єрусалим, за все, що Я навів був на нього.
EZEK|14|23|І потішать вони вас, коли ви побачите їхню дорогу та їхні вчинки, і пізнаєте, що не надармо зробив Я все, що зробив серед нього, говорить Господь Бог.
EZEK|15|1|І було мені слово Господнє таке:
EZEK|15|2|Сину людський, чим краще виноградове дерево від усякого дерева, та виноградна галузка, що була серед дерев лісових?
EZEK|15|3|Чи візьметься з нього кусок дерева, щоб зробити яку роботу? Чи візьмуть із нього кілка, щоб повісити на ньому всяку річ?
EZEK|15|4|Ось воно дане огневі на пожертя... Обидва кінці його пожер огонь, а середина його надгоріла, чи надається воно до роботи?
EZEK|15|5|Як було воно непорушним воно не надавалося на роботу, що ж тепер, коли огонь пожер його, і воно надгоріло, то ще буде надаватися на роботу?
EZEK|15|6|Тому так говорить Господь Бог: Як виноградове дерево між лісними деревами, що Я дав його огневі на пожертя, так дам Я мешканців Єрусалиму!
EZEK|15|7|І оберну Я лице Своє проти них, з одного огню вони вийшли, та пожере їх другий огонь. І пізнаєте, ви, що Я Господь, коли зверну Своє лице проти них!
EZEK|15|8|І віддам цей Край на спустошення, за те, що вони спроневірилися, говорить Господь Бог.
EZEK|16|1|І було мені слово Господнє таке:
EZEK|16|2|Сину людський, повідом Єрусалим про його гидоти,
EZEK|16|3|та й скажи: Так говорить Господь Бог до дочки Єрусалиму: Походження твоє й народження твоє з краю ханаанського, твій батько амореєць, а мати твоя хіттеянка.
EZEK|16|4|При твоєму народженні, того дня, як ти народилася, не був обрізаний пупок твій, і водою не була ти обмита на очищення, ані не була ти посолена, ані не була ти сповита.
EZEK|16|5|Не змилувалося над тобою жодне око, щоб зробити тобі одну з цих речей з милосердя над тобою, але була ти викинена на відкрите поле, так мало ціновано душу твою в день твойого народження!
EZEK|16|6|І проходив Я повз тебе, і бачив тебе, як ти валялася в своїй крові, і сказав Я до тебе: Живи в своїй крові! Так, Я сказав тобі: Живи в своїй крові!
EZEK|16|7|Рости ж, зробив Я тебе, як польову ростину, і ти зросла та стала велика, і дійшла ти до найвродливішої вроди: перса випростались, волос твій виріс, а ти була зовсім нага!
EZEK|16|8|І проходив Я повз тебе, і побачив тебе, аж ось час твій наспів, час кохання. І простягнув Я полу Свою над тобою, і закрив твою наготу, і присягнув тобі, і ввійшов з тобою в заповіт, говорить Господь Бог, і стала ти Моєю.
EZEK|16|9|І обмив Я тебе водою, і сполоскав Я кров твою з тебе, і натер тебе оливою.
EZEK|16|10|І зодягнув тебе різнокольоровим, взув тебе в тахаш, і сповив тебе в віссон, і покрив тебе шовком.
EZEK|16|11|І приоздобив тебе оздобою, і дав нараменники на руки твої, а ланцюга на шию твою.
EZEK|16|12|І дав Я носову сережку до носа твого, і сережки на вуха твої, а пишну корону на твою голову.
EZEK|16|13|І приоздобилась ти золотом та сріблом, а одіж твоя віссон та шовк, і різнокольорове; булку й мед та оливу ти їла, і стала ти гарна-прегарна, і вдалося тобі досягти царської гідности!
EZEK|16|14|І розійшлося ім'я твоє поміж народами за твою красу, бо досконала вона, через пишноту Мою, яку Я на тебе поклав, говорить Господь Бог!
EZEK|16|15|І покладалася ти на красу свою, і стала розпусною через славу свою, і виливала ти розпусту свою на кожного перехожого, його ти була.
EZEK|16|16|І брала ти з шат своїх, і робила собі різнокольорові пагірки, і чинила розпусту на них, як не бувало й не буде.
EZEK|16|17|І брала ти речі з пишноти своєї, з Мого золота та зо срібла Мого, що дав тобі Я, і наробила собі подоб чоловічої статі, і чинила розпусту із ними.
EZEK|16|18|І брала ти свою різнокольорову одіж, і покривала їх, а оливу Мою та Моє кадило клала перед ними.
EZEK|16|19|А Мій хліб, що давав Я тобі, булку й оливу та мед, що ними годував Я тебе, то віддавала ти те перед їхнє обличчя на любі пахощі. І сталося це, говорить Господь Бог.
EZEK|16|20|І брала ти синів своїх та дочок своїх, що породила Мені, і приносила їх на їжу їм. Чи мало було розпусти твоєї,
EZEK|16|21|що ти різала дітей Моїх і давала їм, перепроваджуючи через огонь для них?
EZEK|16|22|І при всіх гидотах твоїх та розпустах твоїх ти не пам'ятала про дні своєї молодости, коли була нагою-пренагою, коли валялася в крові своїй...
EZEK|16|23|І сталося по всьому тому твоєму злі, горе, горе тобі! говорить Господь Бог,
EZEK|16|24|і побудувала ти собі місця розпусти, і поробила собі підвищення на кожному майдані.
EZEK|16|25|На кожному роздоріжжі побудувала ти свої підвищення, і знеславила красу свою, і розхиляла ноги свої для кожного перехожого, і побільшувала свою розпусту...
EZEK|16|26|І чинила ти розпусту з синами Єгипту, з своїми сусідами великотелесими, і побільшувала свою розпусту, щоб гнівити Мене.
EZEK|16|27|І ось простягнув Я Свою руку на тебе, і відняв належну частину твою, і дав тебе на волю твоїх ненависниць, филистимських дочок, засоромлених твоєю нечистою дорогою.
EZEK|16|28|Бо чинила ти розпусту з синами Ашшуровими, і не могла насититись, і блудила з ними, і теж не наситилась.
EZEK|16|29|І побільшила ти свою розпусту до купецького краю халдеїв, та теж цим не наситилася.
EZEK|16|30|Як змучилося серце твоє, говорить Господь Бог, коли ти робила всі оці вчинки свавільної розпусної жінки!
EZEK|16|31|Коли ти будувала місця своєї розпусти на кожному роздоріжжі, а підвищення своє робила на кожному майдані, то не була ти, як блудниця, щоб збирати заплату за розпусту,
EZEK|16|32|але як перелюбна жінка, що замість свого чоловіка бере собі чужих.
EZEK|16|33|Усім блудницям дають дарунка, а ти сама давала дарунки свої всім коханцям своїм, і підкуповувала їх, щоб приходили до тебе звідусіль на розпусту з тобою.
EZEK|16|34|І було тобі при твоїй розпусті навпаки від інших жінок, бо не волочились за тобою, а через те, що ти давала заплату за розпусту, і заплата за розпусту не давалась тобі, то сталось тобі навпаки.
EZEK|16|35|Тому то, розпуснице, послухай Господнього слова:
EZEK|16|36|Так говорить Господь Бог: За те, що виливалась твоя розпуста, і відкривалась твоя нагота в блудодійстві твоїм з твоїми коханцями та зо всіма божками гидоти твоєї, і за кров синів твоїх, яких ти давала їм,
EZEK|16|37|тому ось Я позбираю всіх коханців твоїх, яким була ти приємна, і всіх, кого ти кохала, разом з тими, кого ти зненавиділа, і зберу їх коло тебе знавкола, і відкрию їм наготу твою, і вони побачать увесь твій сором!
EZEK|16|38|І засуджу тебе присудом на перелюбниць та тих, що кров проливають, і дам тебе на кров лютости та заздрости...
EZEK|16|39|І віддам тебе в їхню руку, і вони зруйнують твоє місце розпусти, і порозвалюють підвищення твої, і постягають з тебе шати твої, і позабирають пишні вбрання твої, і покладуть тебе зовсім нагою...
EZEK|16|40|І зберуть проти тебе збори, і закидають тебе камінням, і порубають тебе своїми мечами...
EZEK|16|41|І попалять доми твої огнем, і зроблять на тебе присуди на очах багатьох жінок. І зроблю Я кінець, щоб не була ти розпусницею, і ти вже не будеш давати дарунка за розпусту!
EZEK|16|42|І заспокоїться Моя лютість на тебе, і відійде від тебе Моя заздрість, і я заспокоюся, і не буду вже гніватися.
EZEK|16|43|За те, що ти не пам'ятала про дні своєї молодости, і гнівила Мене всім тим, то й Я ось поверну дорогу твою на твою голову, говорить Господь Бог, щоб не чинила ти розпусти після всіх гидот своїх!...
EZEK|16|44|Ось кожен приповістник говоритиме про тебе приповістку, кажучи: Яка мати така її донька!
EZEK|16|45|Ти дочка своєї матері, що покинула свого чоловіка та своїх синів, і ти сестра своїх сестер, що покидали своїх чоловіків та своїх синів. Мати ваша хіттейка, а ваш батько амореєць!
EZEK|16|46|А старша сестра твоя Самарія та дочки її, що сидять по лівиці твоїй, а сестра твоя, менша від тебе, що сидить по правиці твоїй це Содома та дочки її.
EZEK|16|47|А ти хіба не ходила їхніми дорогами й не робила за їхніми гидотами? Мало бракувало, і зіпсулася б ти більше від них на всіх своїх дорогах!
EZEK|16|48|Як живий Я, говорить Господь Бог, не зробила Содома, сестра твоя, вона та дочки її, як зробила ти та твої дочки!
EZEK|16|49|Ось оце була провина твоєї сестри Содоми: пиха, ситість їжі та преспокійний спокій були в неї та в її дочок, а руки вбогого та бідного вона не зміцняла.
EZEK|16|50|І запишались вони, і робили гидоти перед Моїм обличчям. І Я їх відкинув, як побачив оце.
EZEK|16|51|А Самарія не нагрішила й половини гріхів твоїх, та ти побільшила гидоти свої більш від них, і оправдала сестер своїх усіма своїми гидотами, які ти зробила.
EZEK|16|52|Тож носи свою ганьбу ти, що чинила її для своїх сестер, через твої гріхи, якими гидоти чинила ти більше за них, вони будуть справедливіші за тебе! І також посоромся, і носи свій сором за твоє всправедливлення своїх сестер!
EZEK|16|53|І поверну Я їхню долю, долю Содоми та дочок її, і Самарію та дочок її, і поверну долю твою серед них,
EZEK|16|54|щоб носила ти свій сором, і соромилася всього того, що ти наробила, потішаючи їх.
EZEK|16|55|А твої сестри, Содома та дочки її, вернуться до свого попереднього стану, і Самарія та дочки її вернуться до свого попереднього стану, і ти та дочки твої вернетесь до свого попереднього стану.
EZEK|16|56|І не була сестра твоя Содома згадувана в устах твоїх за днів твоїх гордощів,
EZEK|16|57|поки не відкрилося зло твоє, коли ганьбили тебе дочки Сирії та всіх околиць його, і дочки филистимські погорджували тебе звідусіль.
EZEK|16|58|Свою розпусту та гидоти свої, ти їх понесеш, говорить Господь.
EZEK|16|59|Бо так говорить Господь Бог: І зроблю Я з тобою, як робила ти, що погордила присягою, щоб зламати заповіта.
EZEK|16|60|І згадаю Я Свого заповіта з тобою за днів твоєї молодости, і поставлю тобі заповіта вічного.
EZEK|16|61|І ти згадаєш про свої дороги й засоромишся, коли ти візьмеш сестер своїх, старших від тебе, разом з меншими від тебе і дам їх тобі за дочок, але не з твого заповіту.
EZEK|16|62|І відновлю Я Свого заповіта з тобою, і ти пізнаєш, що Я Господь,
EZEK|16|63|щоб згадала ти й засоромилася, і не могла більше відкривати уста перед ганьбою своєю, коли прощу тобі все, що ти наробила, говорить Господь Бог.
EZEK|17|1|І було мені слово Господнє таке:
EZEK|17|2|Сину людський, загадай загадку, і склади притчу Ізраїлевому домові,
EZEK|17|3|та й скажи: Так говорить Господь Бог: великий орел великокрилий, з широко розгорненими крилами, повний різнокольорового пір'я, прилетів до Ливану, і взяв верховіття кедру.
EZEK|17|4|Чубка галузок його обірвав, і приніс його до купецького краю, у місті гандлярів поклав його.
EZEK|17|5|І взяв він з насіння тієї землі, і посіяв його до насінневого поля, узяв і засадив його над великими водами, немов ту вербу.
EZEK|17|6|І воно виросло, і стало гіллястим виноградом, низькорослим, що обертав свої галузки до нього, а його коріння були під ним. І стало воно виноградом, і вигнало віття, і пустило галузки.
EZEK|17|7|Та був ще один великий орел, великокрилий та густоперий. І ось той виноград витянув пожадливо своє коріння на нього, і свої галузки пустив до нього, щоб він напоїв його з грядок свого засадження.
EZEK|17|8|Він був посаджений на доброму полі при великих водах, щоб пустив галузки та приніс плід, щоб став пишним виноградом.
EZEK|17|9|Скажи: Так говорить Господь Бог: Чи поведеться йому? Чи не вирвуть коріння його, і не позривають плоду його, так що він засохне? Усе зелене галуззя його посохне, і не треба великого рамена та численного народу, щоб вирвати його з його коріння.
EZEK|17|10|І ось хоч він засаджений, чи поведеться йому? Чи всихаючи, не всохне він, як тільки доторкнеться його східній вітер? Він усохне на грядках, де посаджений...
EZEK|17|11|І було мені слово Господнє таке:
EZEK|17|12|Скажи ж домові ворохобному: чи ви не пізнали, що це? Скажи: Ось прийшов вавилонський цар до Єрусалиму, і взяв його царя та його князів, і відвів їх до себе до Вавилону.
EZEK|17|13|І взяв із царського насіння, і склав з ним умову, і ввів його в присягу, і забрав потужних землі,
EZEK|17|14|щоб це було царство низьке, щоб воно не підіймалося, щоб дотримувало його умову, і було їй вірним.
EZEK|17|15|Але той збунтувався проти нього, послав своїх послів до Єгипту, щоб дали йому коней та багато народу. Чи йому поведеться? Чи втече той, хто робить таке? А коли зламає умову, то чи врятується він?
EZEK|17|16|Як живий Я, говорить Господь Бог, у місці царя, який поставив його царем, той, що погордив його присягою та зламав свою умову з ним, помре в нього в Вавилоні!
EZEK|17|17|І фараон не поможе йому на війні великим військом та численним народом, коли насиплють вала та збудують башту, щоб вигубити багато душ.
EZEK|17|18|І погордив він присягою, щоб зламати умову, хоч дав був свою руку, і все те зробив, тому він не врятується.
EZEK|17|19|Тому так говорить Господь Бог: Як живий Я, присягу Мою, якою він погордив, та умову Мою, яку він зламав, дам це на його голову!
EZEK|17|20|І розтягну над ним Свою сітку, і буде він схоплений в пастку Мою, і спроваджу його до Вавилону, і розсуджуся з ним там за його спроневірення, яке він спроневірив проти Мене.
EZEK|17|21|І всі втікачі його з усіх його полків попадають від меча, а позосталі будуть розпорошені на всі вітри. І пізнаєте ви, що Я, Господь, говорив!
EZEK|17|22|Так говорить Господь Бог: І візьму Я з верховіття високого кедру, і дам до землі. З чубка галузок його вирву тендітну, і Сам посаджу на високій та стрімкій горі.
EZEK|17|23|На високій горі Ізраїлевій посаджу її, і вона випустить галузку й принесе плід, і стане сильною кедриною. І буде пробувати під ними усяке птаство, усяке крилате буде перебувати в тіні його галузок.
EZEK|17|24|І пізнають усі польові дерева, що Я, Господь, понизив високе дерево, повищив дерево низьке, висушив дерево зелене, і дав розцвістися дереву сухому. Я, Господь, говорив і вчинив!
EZEK|18|1|І було мені слово Господнє таке:
EZEK|18|2|Що це вам, що ви складаєте приповістку на Ізраїлеву землю, говорячи: Батьки їли неспіле, а оскома в синів на зубах!
EZEK|18|3|Як живий Я, говорить Господь Бог, не будете вже складати тієї приповістки в Ізраїлі!
EZEK|18|4|Тож усі душі Мої: як душа батькова, так і душа синова Мої вони! Душа, що грішить, вона помре.
EZEK|18|5|А чоловік, коли він справедливий, і робить право та справедливість,
EZEK|18|6|на горах жертвенного не їсть, і очей своїх не зводить до божків Ізраїлевого дому, і жінки свого ближнього не занечищує, а до жінки в часі її нечистоти не наближується,
EZEK|18|7|і нікого не тисне, боржникові заставу його конче звертає, грабунку не чинить, хліб свій дає голодному, а голого покриває одежею,
EZEK|18|8|на лихву не дає, а відсотків не бере, від кривди відвертає руку свою, чинить правдивий суд поміж чоловіком та чоловіком,
EZEK|18|9|уставами Моїми ходить, а прав Моїх дотримує, щоб чинити правду, справедливий такий конче буде жити, говорить Господь Бог!
EZEK|18|10|А як породить він сина насильника, що кров проливає, і робить хоч тільки одне з того,
EZEK|18|11|чого він усього того не робив, а також на горах жертвенне їв, і жінку свого ближнього занечищував,
EZEK|18|12|убогого й бідаря утискав, грабунки чинив, застави боржникові не звертав, і до божків зводив свої очі, гидоту робив,
EZEK|18|13|на лихву давав, і відсоток брав, то чи буде він жити? Не буде він жити! Він усі ті гидоти чинив, він мусить конче померти, кров його буде на ньому!
EZEK|18|14|А ось породив він сина, і той побачив усі гріхи свого батька, які той робив, і хоч бачив, та не робив, як той:
EZEK|18|15|на горах жертвенного не їв, і очей своїх до божків Ізраїлевого дому не зводив, жінки свого ближнього не занечищував,
EZEK|18|16|і нікого не утискав, застави у застав не брав, і грабунку не чинив, хліб свій голодному давав, а голого одежею покривав,
EZEK|18|17|від кривди свою руку відвертав, лихви та відсотків не брав, права Мої чинив, уставами Моїми ходив, такий не помре за провину свого батька, він конче буде жити!
EZEK|18|18|Батько ж його, за те, що утиском тиснув, грабунком грабував брата, і що недобре чинив серед народу свого, то ось він помре за провину свою!
EZEK|18|19|А скажете ви: Чому той син не поніс провину за батька? Але ж син той чинив право та справедливість, дотримував усі устави Мої й виконував їх, він конче буде жити!
EZEK|18|20|Та душа, що грішить, вона помре. Син не понесе кари за батькову провину, а батько не понесе за провину синову, справедливість справедливого буде на ньому, а несправедливість несправедливого на тому буде.
EZEK|18|21|А коли б несправедливий відвернувся від усіх гріхів своїх, яких наробив, і виконував усі устави Мої, і робив право та справедливість, буде конче він жити, не помре!
EZEK|18|22|Усі його гріхи, які наробив він, не згадаються йому, він буде жити в своїй справедливості, яку чинив!
EZEK|18|23|Чи Я маю вподобання в смерті несправедливого? говорить Господь Бог, чи ж не в тому, щоб він повернувся з доріг своїх та й жив?
EZEK|18|24|А коли б справедливий відвернувся від своєї справедливости й став робити кривду, усі ті гидоти, які робить несправедливий, то чи такий буде жити? Усі справедливості його, які він робив, не згадаються, за своє спроневірення, що він спроневірив, і за гріх свій що згрішив, за них він помре!
EZEK|18|25|А ви кажете: Неправа Господня дорога! Послухайте но, доме Ізраїлів, чи ж дорога Моя неправа? Чи не ваші дороги неправі?
EZEK|18|26|Коли б справедливий відвернувся від своєї справедливости й чинив кривду, і за те помер, то він помре за кривду свою, яку він чинив.
EZEK|18|27|А коли б несправедливий відвернувся від своєї несправедливости, яку він чинив, і чинив би право та справедливість, він душу свою при житті збереже.
EZEK|18|28|І коли б він побачив, і відвернувся від усіх своїх гріхів, які він чинив, то конче буде він жити, не помре!
EZEK|18|29|А Ізраїлів дім каже: Неправа Господня дорога! Чи ж Мої дороги неправі, доме Ізраїлів? Чи ж то не ваші дороги неправі?
EZEK|18|30|Тому буду судити вас, доме Ізраїлів, кожного за дорогами його, говорить Господь Бог. Покайтеся, і відверніться від усіх ваших гріхів, і не буде вам провина на спотикання!
EZEK|18|31|Поскидайте з себе всі ваші гріхи, якими ви грішили, і створіть собі нове серце та нового духа! І нащо маєте померти, Ізраїлів доме?
EZEK|18|32|Бо не жадаю Я смерти помираючого, говорить Господь Бог, але покайтеся та й живіть!
EZEK|19|1|А ти пісню жалобну здійми про князів Ізраїлевих,
EZEK|19|2|та й скажи: Яка твоя мати левиця: Лягла поміж левів, серед левчуків вона викохала левенят!
EZEK|19|3|І одне із своїх левенят вона вигодувала, левчуком воно стало, і здобич ловити навчився, людину він жер!
EZEK|19|4|І похід розголосили народи на нього, в їхню яму він схоплений був, і його в ланцюгах до краю єгипетського відвели...
EZEK|19|5|Як левиця побачила, що надаремно чекає, що пропала надія її, то взяла вона знову одне із своїх левенят, і вчинила його левчуком.
EZEK|19|6|І ходив він між левами й став левчуком, і здобич ловити навчився, людину він жер!
EZEK|19|7|І він розбивав їхні палати, і руйнував їхні міста, і від голосу рику його остовпіла земля й що на ній!
EZEK|19|8|Та пастку на нього поставили люди знавкола з округ, і свою сітку на нього розкинули, і він схоплений був в їхню яму!
EZEK|19|9|І кинули в клітку його в ланцюгах, і його відвели до царя вавилонського, і в твердиню його запроторили, щоб голос його вже не чувся на горах Ізраїлевих...
EZEK|19|10|Твоя мати, як той виноград у винограднику, посадженому над водою, плодюча й гілляста була через води великі.
EZEK|19|11|І виросли пруття міцні, й надавались на берла володарів, і височів між гущавинами його зріст, і він показався в своїй висоті, у численних галузках своїх!
EZEK|19|12|Та була вона вирвана в лютості, об землю кинена, і вітер зо сходу зсушив її плід, поламалися й повисихали вони, а її міцний прут огонь його зжер...
EZEK|19|13|А тепер посадили її на пустині, у краї сухому й безвідному,
EZEK|19|14|і вийшов огонь із прута її вітки та й пожер її плід, і немає у неї міцного прута, берла на панування... Це пісня жалобна, і буде за пісню жалоби вона.
EZEK|20|1|І сталося за сьомого року, в п'ятому місяці, у десятому дні місяця, поприходили люди з Ізраїлевих старших, щоб запитатися в Господа, і посідали передо мною.
EZEK|20|2|І було мені слово Господнє таке:
EZEK|20|3|Сину людський, говори з Ізраїлевими старшими та й скажеш до них: Так говорить Господь Бог: Чи ви прийшли, щоб запитатися в Мене? Як живий Я, не відповім вам, говорить Господь Бог!
EZEK|20|4|Чи ти розсудиш їх, чи ти їх розсудиш, сину людський? Завідом їх про гидоти їхніх батьків,
EZEK|20|5|та й скажеш до них: Так говорить Господь Бог: Того дня, коли Я був вибрав Ізраїля, і підніс Свою руку до насіння Якового дому, і відкрився їм в єгипетському краї, і підніс Свою руку до них, говорячи: Я Господь, Бог ваш,
EZEK|20|6|того дня Я підніс Свою руку до них, щоб вивести їх з єгипетського краю до Краю, що Я вислідив для них, що тече молоком та медом, що він окраса для всіх країв.
EZEK|20|7|І сказав Я до них: Відкидайте кожен гидоти від очей своїх, і не занечищуйтеся божками Єгипту. Я Господь, Бог ваш!
EZEK|20|8|Та були вони ворохобні проти Мене, і не хотіли слухатися Мене, не відкидали кожен гидот від очей своїх, і не покинули єгипетських божків. І подумав Я, що виллю на них Свою лютість, що докінчу на них Свій гнів посеред єгипетського краю.
EZEK|20|9|І зробив Я ради Свого Ймення, щоб воно не безчестилося на очах тих народів, що вони серед них, що Я відкрився їм на їхніх очах, щоб вивести їх з єгипетського краю.
EZEK|20|10|І вивів Я їх з єгипетського краю, і спровадив їх до пустині.
EZEK|20|11|І дав їм постанови Свої, і познайомив їх з постановами Моїми, які коли чинитиме людина, то житиме ними.
EZEK|20|12|І також дав Я їм Свої суботи, щоб були вони знаком поміж Мною та між ними, щоб пізнати, що Я Господь, що освячує їх.
EZEK|20|13|Та став ворохобним проти мене Ізраїлів дім на пустині, уставами Моїми не ходили вони, і повідкидали Мої постанови, які коли чинить людина, то житиме ними, а суботи Мої дуже зневажали. Тому Я сказав був, що виллю лютість Свою на них на пустині, щоб вигубити їх.
EZEK|20|14|Та зробив Я ради Ймення Свого, щоб воно не зневажалося на очах тих народів, що на їхніх очах Я вивів їх.
EZEK|20|15|Але й Я, прирікаючи, підніс їм Свою руку на пустині, що не впроваджу їх до Краю, якого Я дав, що тече молоком та медом, що окраса він для всіх країв,
EZEK|20|16|за те, що постанови Мої вони відкинули, а устави Мої не ходили вони ними, і суботи Мої зневажали, бо за своїми божками ходило їхнє серце...
EZEK|20|17|І змилувалось Моє око над ними, щоб не нищити їх, і не зробив Я з ними кінця на пустині.
EZEK|20|18|І сказав Я їхнім синам на пустині: Уставами ваших батьків не ходіть, і постанов їхніх не перестерігайте, і божками їхніми не занечищуйтесь!
EZEK|20|19|Я Господь, Бог ваш, уставами Моїми ходіть, і постанови Мої перестерігайте й виконуйте їх.
EZEK|20|20|І святіть суботи Мої, і вони стануть знаком поміж Мною та між вами, щоб пізнати, що Я Господь, Бог ваш!
EZEK|20|21|Та стали ворохобні ті сини проти Мене, уставами Моїми не ходили, а постанов Моїх не перестерігали, щоб виконувати їх, які коли робить людина, то житиме ними, і суботи Мої зневажали. І подумав Я був, що виллю лютість Свою на них, щоб заспокоїти гнів Мій на них на пустині.
EZEK|20|22|І відвернув Я Свою руку, і зробив ради Ймення Свого, щоб не зневажати його на очах тих народів, що на їхніх очах Я їх вивів.
EZEK|20|23|Та й Я, прирікаючи, підніс їм Свою руку на пустині, щоб розпорошити їх серед народів і порозсипати їх по краях,
EZEK|20|24|за те, що постанов Моїх не чинили, і устави Мої відкинули, а суботи Мої зневажали, і до божків своїх батьків були їхні очі.
EZEK|20|25|І тому Я дав їм мати устави недобрі, і постанови, що не будуть вони жити ними.
EZEK|20|26|І занечистив Я їх їхніми дарунками, перепровадженням через огонь кожного, хто відкриває утробу, щоб спустошити їх, щоб пізнали вони, що Я Господь!
EZEK|20|27|Тому говори до Ізраїлевого дому, сину людський, і скажи до них: Так говорить Господь Бог: Ще оцим зневажали Мене батьки ваші, коли спроневірилися проти Мене:
EZEK|20|28|коли Я ввів їх до Краю, що про нього, прирікаючи, підносив Я Свою руку дати його їм, то коли вони бачили всякий високий пагірок і всяке густе дерево, то приносили там свої жертви, і давали там свої дари, що гнівили Мене, і складали там свої любі пахощі, і приносили там свої литі жертви.
EZEK|20|29|І сказав Я до них: Що це за висота, що ви ходите туди? І зветься вона Бама аж до цього дня.
EZEK|20|30|Тому скажи до Ізраїлевого дому: Так говорить Господь Бог: Чи ви будете занечищуватися дорогою своїх батьків і будете ходити в розпусті за гидотами їхніми?
EZEK|20|31|А приношенням ваших дарів, перепровадженням ваших синів через огонь ви занечищуєтеся при всіх ваших божках аж до сьогодні. А ви хочете питати Мене, Ізраїлів доме? Як живий Я, говорить Господь Бог, не дам Я вам відповіді!
EZEK|20|32|А що входить вам на серце, зовсім не станеться те, що ви говорите: Будемо, як інші народи, як племена Краю, служити дереву та каменю.
EZEK|20|33|Як живий Я, говорить Господь Бог, рукою потужною й витягненим раменом та виливаною лютістю буду царювати над вами!
EZEK|20|34|І виведу вас із тих народів, і позбираю вас із тих країв, де ви розпорошені рукою потужною й витягненим раменом та виливаною лютістю.
EZEK|20|35|І заведу вас до пустині народів, і буду там судитися з вами лицем до лиця,
EZEK|20|36|як судився Я з вашими батьками на пустині єгипетського краю, так буду судитися з вами, говорить Господь Бог!
EZEK|20|37|І проведу вас під палицею, і введу вас у зв'язок заповіту.
EZEK|20|38|І повибираю з вас бунтівників та тих, що грішать проти Мене, повипроваджую їх з краю їхнього пробування, і до Ізраїлевої землі вже не ввійдуть вони! І пізнаєте ви, що Я Господь!
EZEK|20|39|А ви, Ізраїлів доме, так говорить Господь Бог: Кожен ідіть, служіть своїм божкам! Але потім ви напевно будете слухатися Мене, і святого Ймення Мого ви вже не зневажите своїми дарунками та своїми божками...
EZEK|20|40|Бо на Моїй святій горі, на високій Ізраїлевій горі, говорить Господь Бог, там буде служити Мені ввесь Ізраїлів дім, увесь він, що в Краю, там Я їх уподобаю Собі, і там зажадаю ваших приношень і первоплодів ваших приношень у всіх ваших святощах!
EZEK|20|41|Любими пахощами вподобаю Собі вас, коли вас виведу з народів, і зберу вас із тих країв, де ви розпорошені, і буду Я святитися між вами на очах усіх поган.
EZEK|20|42|І пізнаєте ви, що Я Господь, коли впроваджу вас до Ізраїлевої землі, до того Краю, що про нього, прирікаючи, підніс Я Свою руку дати його вашим батькам.
EZEK|20|43|І згадаєте там свої дороги, і всі свої вчинки, якими ви занечистилися, і почуєте огидження перед самими собою за всі ваші лиха, які наробили...
EZEK|20|44|І пізнаєте, що я Господь, коли Я чинитиму з вами ради Ймення Свого, а не за вашими злими дорогами та за вашими зіпсутими вчинками, доме Ізраїлів, говорить Господь Бог.
EZEK|20|45|(21-1) І було мені слово Господнє таке:
EZEK|20|46|(21-2) Сину людський, зверни обличчя своє в напрямі на південь, і крапай словами на полудень, і пророкуй на ліс південного поля.
EZEK|20|47|(21-3) І скажи до південного лісу: Послухай Господнього слова: Так говорить Господь Бог: Ось у тобі запалю Я огонь, і поїсть він у тебе кожне дерево зелене, і кожне дерево сухе; полум'яний огонь не погасне, і будуть попалені ним всі простори від півдня до півночі.
EZEK|20|48|(21-4) І побачить кожне тіло, що Я, Господь, розпалив його, і він не погасне!
EZEK|20|49|(21-5) І сказав я: О Господи, Боже, вони мені кажуть: Чи він не говорить самі тільки притчі?
EZEK|21|1|(21-6) І було мені слово Господнє таке:
EZEK|21|2|(21-7) Сину людський, зверни ти обличчя своє до Єрусалиму, і крапай словами на святині, і пророкуй на землю Ізраїлеву.
EZEK|21|3|(21-8) І скажи Ізраїлевій землі: Так говорить Господь: Ото Я проти тебе, і меча Свого витягну з піхви його, і витну з тебе справедливого й несправедливого.
EZEK|21|4|(21-9) Через те, що Я витну з тебе справедливого й несправедливого, тому вийде Мій меч проти кожного тіла від півдня на північ.
EZEK|21|5|(21-10) І кожне тіло пізнає, що Я Господь, витяг меча Свого з піхви його, уже не вернеться він!
EZEK|21|6|(21-11) А ти, сину людський, стогни, ніби мав би ти зламані стегна, і гірко стогни на їхніх очах!
EZEK|21|7|(21-12) І буде, коли тобі скажуть: Чого то ти стогнеш? то скажеш: На звістку, що йде, і кожне серце розтане, і всякі руки ослабнуть, і погасне всякий дух, і всі коліна зайдуться водою! Оце прийде та станеться, каже Господь Бог.
EZEK|21|8|(21-13) І було мені слово Господнє таке:
EZEK|21|9|(21-14) Сину людський, пророкуй і кажи: Так говорить Господь: Скажи: Меч, меч, нагострений він та блискучий!
EZEK|21|10|(21-15) Щоб приносити жертву нагострений він, щоб блищати він був полірований. Хіба будемо радіти? Хіба жезло сина Мого легковажить усякеє дерево?
EZEK|21|11|(21-16) І дали його виполірувати, щоб узяти в долоню. Це нагострений меч, і він полірований, щоб дати його в руку вбивця...
EZEK|21|12|(21-17) Кричи та реви, сину людський, бо він проти народу Мого, він проти всіх князів Ізраїлевих, їх віддано мечеві з народом Моїм, тому вдарся по стегнах!
EZEK|21|13|(21-18) Та він уже випробуваний. Та що ж тепер, коли йому жезло обридло? Він не встоїть, каже Господь Бог.
EZEK|21|14|(21-19) А ти, сину людський, пророкуй, і вдар долонею об долоню, і нехай меч подвоїться та потроїться! Це меч побитих, великий меч забитого, що кружляє довкола них.
EZEK|21|15|(21-20) Щоб стопилося серце й полягло якнайбільше при всіх їхніх брамах, Я дам різанину меча. О горе, він справді зроблений блискучим, виполіруваним на різанину!
EZEK|21|16|(21-21) Об'єднайся, праворуч іди, зверни ліворуч, іди, куди тільки звернене буде вістря твоє...
EZEK|21|17|(21-22) І Я вдарю долоню Свою об долоню Свою, і Свою лють заспокою. Я, Господь, це прорік!
EZEK|21|18|(21-23) І було мені слово Господнє таке:
EZEK|21|19|(21-24) А ти, сину людський, признач собі дві дорозі, якими прибуде меч вавилонського царя. Вони вийдуть обидві із краю одного, а ти вистругай дороговказну руку, на початку дороги до міста її вистругай.
EZEK|21|20|(21-25) Признач дорогу, якою прибуде меч до Рабби Аммонових синів та до Юди в укріплений Єрусалим.
EZEK|21|21|(21-26) Бо цар вавилонський став на роздоріжжі, на початку двох доріг. Щоб ворожити чарами, трясе він стрілами, питає домашніх божків, розглядає печінку.
EZEK|21|22|(21-27) У правиці його був чар на Єрусалим, щоб поставити муроломи, щоб відкрити уста на крик, щоб підняти голос окриком, щоб поставити муроломи на брами, щоб насипати вала, щоб збудувати башту.
EZEK|21|23|(21-28) Але буде це їм в їхніх очах, як чарування марнотне, буде для них заприсяження присягами, та він згадає провину, щоб були вони схоплені.
EZEK|21|24|(21-29) Тому так говорить Господь Бог: За те, що ви згадуєте свої провини, що відкриваєте ваші гріхи, щоб бачені були ваші гріхи ваших учинків, за те, що ви пригадуєте, у ворожі руки схоплені будете!
EZEK|21|25|(21-30) А ти, недостойний, несправедливий князю Ізраїлів, що надійшов його день у час провини кінцевої,
EZEK|21|26|(21-31) так говорить Господь Бог: Зняти завоя й скинути корону! Це не зостанеться так, піднесеться низьке, а високе понизиться!
EZEK|21|27|(21-32) Руїною, руїною, руїною покладу його! Та цього не станеться, аж поки не прийде Той, Хто має право, і Я Йому дам!
EZEK|21|28|(21-33) А ти, сину людський, пророкуй та й скажеш: Так говорить Господь Бог на Аммонових синів та про їхню ганьбу: І скажеш: Меч, меч відкритий на різанину, блискучий, щоб блищав, як та блискавка,
EZEK|21|29|(21-34) для тебе бачили обманні видіння, пророкували для тебе неправду, щоб посадити його на шию недостойних злочинців, яких день прийде в час кари кінцевої.
EZEK|21|30|(21-35) Верни ж меча до піхви його! У місці, де створений ти, у краю походження твого осуджу Я тебе!
EZEK|21|31|(21-36) І виллю на тебе Свій гнів, в огні пересердя Свого на тебе дмухну, і дам тебе в руку людей зухвалих, які знищення замишляють!
EZEK|21|32|(21-37) Ти станеш огневі на їжу, твоя кров буде серед землі, не згадають про тебе, бо Я, Господь, говорив це!
EZEK|22|1|І було мені слово Господнє таке:
EZEK|22|2|А ти, сину людський, чи будеш судити, чи судитимеш ти місто крови? І завідом його про всі гидоти його,
EZEK|22|3|та й скажеш: Так говорить Господь Бог: Місто проливає кров у своїй середині, щоб прийшов його час, і робить божків собі, щоб занечищуватися!
EZEK|22|4|Кров'ю, що ти проливала, о дочко Єрусалиму, грішила ти, а божками, яких ти робила, занечистилася, і наблизила свої дні, і прийшла аж до своїх років. Тому дам тебе народам на ганьбу, і на посміховисько для всіх країв!
EZEK|22|5|Близькі та далекі від тебе насміхаються з тебе, нечистойменна, багатозаколотна!
EZEK|22|6|Ось Ізраїлеві князі, кожен за раменом своїм, були в тебе, щоб кров проливати.
EZEK|22|7|Батька та матір у тебе легковажать, чужинцеві роблять утиск серед тебе, сироту та вдову пригнічуть у тебе.
EZEK|22|8|Моїми святощами ти погорджуєш, а суботи Мої зневажаєш.
EZEK|22|9|У тебе є наклепники, щоб кров проливати, і на пагірках їдять у тебе, розпусту чинять серед тебе.
EZEK|22|10|Наготу батька в тебе відкривають, жінку, у часі її місячної нечистоти, безчестять у тебе.
EZEK|22|11|І один робить гидоту з жінкою свого ближнього, а той занечищує розпустою невістку свою, а той безчестить у тебе сестру свою, дочку батька свого...
EZEK|22|12|Підкуп беруть у тебе, щоб кров проливати, лихву та відсотка береш ти й ошукуєш утиском ближніх своїх. А Мене ти забуваєш, говорить Господь Бог...
EZEK|22|13|І ось сплеснув Я руками Своїми за твою кривду, яку ти робила, та за кровопролиття твої, що були в тебе.
EZEK|22|14|Чи встоїть твоє серце, чи будуть міцні твої руки на ті дні, що Я буду з тобою чинити? Я, Господь, говорив це й зробив!
EZEK|22|15|І розпорошу тебе серед народів, і розсиплю тебе по краях, і викину твою нечистість із тебе.
EZEK|22|16|І станеш ти збезчещеною через себе на очах народів, і пізнаєш, що Я Господь!...
EZEK|22|17|І було мені слово Господнє таке:
EZEK|22|18|Сину людський, дім Ізраїлів став мені за жужелицю; усі вони мідь, і цина, і залізо, і оливо в середині горна, жужелицею срібла сталися.
EZEK|22|19|Тому так говорить Господь Бог: За те, що всі ви стали жужелицею, тому ось Я позбираю вас до середині Єрусалиму.
EZEK|22|20|Як збирають срібло, і мідь, і залізо, і оливо, і цину до середини горна, щоб дмухати на нього огнем, щоб розтопити, так зберу у Своїм гніві та в люті Своїй, і покладу, і розтоплю вас!
EZEK|22|21|І позбираю вас, і дмухну на вас огнем Свого гніву, і ви будете розтоплені в середині його...
EZEK|22|22|Як розтоплюється срібло в середині горна, так будете розтоплені ви в середині його, і пізнаєте, що Я, Господь, вилив гнів Свій на вас!...
EZEK|22|23|І було мені слово Господнє таке:
EZEK|22|24|Сину людський, скажи до неї: Ти земля неочищена, у дні гніву дощем не политая!
EZEK|22|25|Змова її пророків серед нього, як ревучий лев, що здобич шматує: жеруть душу, маєток та багатство забирають, прибільшують удів її в середині її.
EZEK|22|26|Священики її ламають Закона Мого, і зневажають Мої святощі, не розрізняють між святим та несвятим, і не оголошують різниці між нечистим та чистим, від субіт Моїх закривають свої очі. І був Я зневажений серед них.
EZEK|22|27|Князі її в середині її, немов ті вовки, що здобич шматують, щоб розливати кров, щоб губити душі ради користи.
EZEK|22|28|А пророки її все замазують болотом, бачать марноту, і чарують собі неправдою, вони кажуть: Так говорить Господь Бог, а Господь не говорив...
EZEK|22|29|Народи Краю тиснуть утиском та грабують грабунком, а вбогого та бідака гноблять, а чужинця тиснуть у безправ'ї...
EZEK|22|30|І шукав Я між ними чоловіка, що поставив би загороду, і став би в виломі перед Моїм обличчям за цей Край, щоб Я не знищив його, та Я не знайшов!
EZEK|22|31|І Я вилив на них Свій гнів, огнем пересердя Свого повигублював їх, їхню дорогу Я дав на їхню голову, каже Господь Бог...
EZEK|23|1|І було мені слово Господнє таке:
EZEK|23|2|Сину людський, були собі дві жінки, дочки однієї матері.
EZEK|23|3|І чинили вони в Єгипті розпусту, у своїй молодості чинили розпусту, там почавлені їхні груди, там замацані їхні перса дівочі.
EZEK|23|4|А їхні імена: Огола старша та Оголива сестра її. І стали вони Мої, і породили синів та дочок. А їхні імена: Самарія Огола, а Єрусалим Оголива.
EZEK|23|5|І стала розпусною Огола, бувши Моєю, і кохалася з своїми коханцями, з асиріянами, хто був їй близький,
EZEK|23|6|що їхнє убрання блакить, намісники та заступники вони, усі вони юнаки вродливі, вершники, що гарцюють на конях.
EZEK|23|7|І дала вона свою розпусту їм, що всі вони добірні Ашшурові сини, і всіма, яких кохала, і всіма своїми божками була вона занечищена.
EZEK|23|8|Та не відкидала вона своєї розпусти й від єгиптян, бо вони лежали з нею в її молодості, і вони стискали дівочі її перса, і виливали свою розпусту на неї...
EZEK|23|9|Тому й дав Я її в руку її коханків, у руку Ашшурових синів, що з ними кохалась вона.
EZEK|23|10|Вони відкрили її наготу, позабирали синів її та дочок її, а її забили мечем... І стала вона неславним ім'ям для жінок, і присуди зробили на ній.
EZEK|23|11|А сестра її Оголива бачила це, але вчинила любов свою гіршою від неї, а розпусту свою більшою від розпусти своєї сестри.
EZEK|23|12|Вона кохалася з синами Ашшуровими, з близькими їй намісниками та заступниками, досконало зодягненими, з верхівцями, що гарцюють на конях, усі вони юнаки вродливі.
EZEK|23|13|І побачив Я, що вона обезчещена, що дорога одна їм обом.
EZEK|23|14|Та вона ще додала до розпусти своєї, бо коли побачила мужів, вирізьблених на стіні, зображення халдеїв, креслених і запущених червонилом,
EZEK|23|15|підперезаних поясом по стегнах своїх, вони з опадаючим завоєм на голові їхній, усі вони на вигляд військові старшини, подоба синів вавилонських, Халдея край народження їхнього,
EZEK|23|16|то пожадала вона їх через сам погляд очей своїх, і послала посланців по них, до Халдеї.
EZEK|23|17|І прийшли до неї сини Вавилону на ложе любовне, і занечистили її своєю розпустою, і вона занечистилася ними, і відвернулася душа її від них...
EZEK|23|18|І відкрила вона розпусту свою, і відкрила свою наготу, тому відвернулася душа Моя від неї, як відвернулася душа Моя від її сестри.
EZEK|23|19|І побільшила вона розпусту свою на згадку днів своєї молодости, коли чинила розпусту в єгипетському краї.
EZEK|23|20|І жадала вона собі на коханців тих, що їхня плоть плоть ослина, а їхня похіть похіть жеребця.
EZEK|23|21|І згадала ти розпусту своєї молодости, коли єгиптяни стискали груди твої ради перс твоєї молодости.
EZEK|23|22|Тому, Оголиво, так говорить Господь Бог: Ось Я збуджу коханців твоїх на тебе, що від них відвернулася душа твоя, і спроваджу їх на тебе з довкілля,
EZEK|23|23|синів Вавилону, і всіх халдеїв, Пекод, і Шоа, і Коа, і всіх синів Ашшурових з ними, уродливі то юнаки, усі вони начальники та заступники, військові старшини та славні, усі вони гарцюють на конях.
EZEK|23|24|І прийдуть на тебе з півночі, з колесницями та з колесами, та зо збором народів; щита великого й щита малого та шоломи покладуть проти тебе навколо. І дам їм право, і вони засудять тебе за своїми правами.
EZEK|23|25|І зверну Я лютість Свою на тебе, і вони зроблять з тобою в гніві: пообтинають носа твого та вуха твої, а що полишиться в тебе, від меча упаде. Вони позабирають синів твоїх та дочок твоїх, а що залишиться в тебе, буде пожерте огнем...
EZEK|23|26|І постягають із тебе шати твої, і позабирають речі пишноти твоєї.
EZEK|23|27|І спиню Я розпусту твою в тебе, і розпусту твою з єгипетського краю, і ти не зведеш очей своїх на них, а про Єгипта вже не згадаєш.
EZEK|23|28|Бо так говорить Господь Бог: Ось Я даю тебе в руку того, кого ти зненавиділа, у руку тих, що від них відвернулася душа твоя.
EZEK|23|29|І зроблять з тобою в ненависті, і візьмуть здобуток твій, і поставлять тебе нагою та голою, і буде відкрита нагота перелюбу твого, і розпуста твоя та твій блуд...
EZEK|23|30|Будуть робити це тобі за твоє ходіння в розпусті з народами, за те, що ти збезчестилась їхніми божками.
EZEK|23|31|Дорогою своєї сестри ти ходила, тому дам її келіха в твою руку.
EZEK|23|32|Так говорить Господь Бог: Келіха своєї сестри ти вип'єш, глибокого та широкого; станеш за жарт та за посміховисько, це багатомісткий келіх.
EZEK|23|33|П'янством та смутком будеш наповнена, буде це келіх спустошення й розруху, келіх твоєї сестри Самарії.
EZEK|23|34|І ти вип'єш його, і витягнеш усе, а череп'я його порозбиваєш, і перса свої порозриваєш, бо це Я говорив, каже Господь Бог.
EZEK|23|35|Тому так говорить Господь Бог: Через те, що ти забула Мене, і кинула мене за спину свою, то й ти носи розпусту свою та свій блуд!
EZEK|23|36|І сказав Господь до мене: Сину людський, чи будеш судити Оголу та Оголиву? То викажи їм їхні гидоти!
EZEK|23|37|Бо вони перелюб чинили, і кров на їхніх руках, і з божками своїми перелюб чинили, і також синів своїх, яких породили Мені, перепроваджували через огонь для них на їжу...
EZEK|23|38|Ще оце чинили Мені: Занечистили святиню Мою того дня, і суботи Мої зневажили.
EZEK|23|39|А коли вони різали синів своїх для своїх божків, то приходили до Моєї святині того дня, щоб збезчестити її, і оце так робили вони в середині Мого дому...
EZEK|23|40|А що більше, посилали до мужів, що здалека приходять, що до них був посланий посланець, і ось поприходили ті, що для них ти вмилася, нафарбувала блакитом очі свої й оздобою приоздобилася.
EZEK|23|41|І сіла ти на дорогоцінному ліжку, а перед ним накритий стіл, і поклала на ньому кадило Моє та оливу Мою.
EZEK|23|42|І голос заспокоєної товпи лунав при ньому, і до мужів тієї товпи спроваджували ще п'яних з пустині, і давали нараменники на їхні руки та пишні корони на їхні голови.
EZEK|23|43|І сказав Я до тієї, що в'янула від перелюбу: Буде тепер вона ще далі чинити розпусту?
EZEK|23|44|І прийшли до неї, як приходять до блудниці, так приходили до Оголи та Оголиви, розпусних жінок.
EZEK|23|45|А люди справедливі вони розсудять їх правом про тих, що чинять перелюб, та правом про тих, що кров проливають, бо вони чинять перелюб, і кров на їхніх руках.
EZEK|23|46|Бо так говорить Господь Бог: Скликати б на них збори, і дати їх на страх та на здобич!
EZEK|23|47|І збори закидають їх камінням, і порозсікають їх своїми мечами, синів їхніх та їхніх дочок повбивають, а їхні доми попалять огнем...
EZEK|23|48|І спиню Я розпусту в Краю, і буде наука всім жінкам, і вони не будуть робити такого, як ваша розпуста!
EZEK|23|49|І покладуть вони вашу розпусту на вас, і ви будете носити гріхи ваших божків. І ви пізнаєте, що Я Господь Бог!
EZEK|24|1|А за дев'ятого року, десятого місяця, десятого дня місяця було мені слово Господнє таке:
EZEK|24|2|Сину людський, напиши собі ім'я цього дня, цього самого дня, бо вавилонський цар саме цього дня наступив на Єрусалим.
EZEK|24|3|І розкажи притчу на дім ворохобности, та й скажеш їм: Так говорить Господь Бог: Пристав ти котла, пристав та й налий води в нього.
EZEK|24|4|Повкладай його кусні до нього, усякий добрий кусок, стегно та лопатку, наповни кістками добірними.
EZEK|24|5|Візьми добірніше з отари, розклади під ним дрова, звари його кусні, і щоб у ньому зварилися кості його.
EZEK|24|6|Тому так Господь Бог промовляє: Горе місту цьому душогубному, котлові, що іржа його в ньому, і що його іржа не сходить із нього! Кусок за куском повитягуй це з нього; на нього нехай не впаде жеребок!
EZEK|24|7|Кров бо його серед нього, він на голу скелю її помістив, не вилив на землю її, щоб порохом вкрити її.
EZEK|24|8|Щоб лютість підійняти, щоб помститися, Я дам його кров на голу скелю, щоб вона непокрита була.
EZEK|24|9|Тому так Господь Бог промовляє: Горе місту цьому душогубному, збільшу огнище й Я!
EZEK|24|10|Підклади дров, розпали цей огонь, довари м'ясо, і вилий росіл, а кості хай спалені будуть.
EZEK|24|11|І постав його порожнім на вугілля його, щоб він розігрівся, і щоб мідь його розпалилась, і щоб розтопилась у ньому нечистість його, щоб іржа його зникла.
EZEK|24|12|Увесь труд надармо пішов, і не зійшла з нього його велика іржа, в огонь його з його іржею!
EZEK|24|13|У твоїй нечистоті є розпуста. За те, що Я чистив тебе, але чистим не став ти, ти з своєї нечистости вже не відчистишся, аж поки Я не заспокою Свою лютість на тобі.
EZEK|24|14|Я, Господь, це казав, і надійде воно! І зроблю, не звільню, і не змилуюся, за твоїми дорогами та за твоїми ділами засудять тебе, це Господь Бог промовляє!
EZEK|24|15|І було мені слово Господнє таке:
EZEK|24|16|Сину людський, ось Я візьму від тебе несподіваним ударом утіху очей твоїх, а ти не голоси й не плач, і нехай не виступить сльоза твоя.
EZEK|24|17|Стогни собі тихо, жалоби по померлих не роби, прикрасу голови своєї обвий на себе, а взуття своє взуй на ноги свої, і не закривай вусів, і не їж жалобного хліба.
EZEK|24|18|І говорив я до народу рано, а ввечері померла мені жінка... І зробив я рано, як наказано мені.
EZEK|24|19|І сказав мені той народ: Чи не розповіси нам, що це нам таке, що ти робиш?
EZEK|24|20|І я їм сказав: Було мені слово Господнє таке:
EZEK|24|21|Скажи Ізраїлевому дому: Так говорить Господь Бог: Ось Я збезчещу святиню Мою, опору вашої сили, утіху ваших очей та любе вашій душі. А ваші сини та ваші дочки, що ви покинули їх, попадають від меча...
EZEK|24|22|І ви зробите, як зробив я: вусів не закриєте, і хліба жалобного не будете їсти...
EZEK|24|23|А прикраси ваші будуть на ваших головах, і взуття ваше на ваших ногах, не будете голосити, і не будете плакати, а будете сохнути через свої гріхи, і будете стогнати один до одного...
EZEK|24|24|І стане Єзекіїль вам за знака: усе, що робив він, будете робити і ви. І коли те прийде, то пізнаєте ви, що Я Господь Бог.
EZEK|24|25|А ти, сину людський, того дня, коли візьму від них їхню силу, радість пишноти їхньої, утіху очей їхніх, прагнення їхньої душі, їхніх синів та дочок їхніх,
EZEK|24|26|того дня прийде до тебе врятований, щоб сповістити про це в твої вуха.
EZEK|24|27|Цього дня відкриються твої уста разом з цим урятованим, і будеш говорити, і не будеш уже німий, і станеш для них знаком. І пізнають, що Я Господь!
EZEK|25|1|І було мені слово Господнє таке:
EZEK|25|2|Сину людський, зверни своє обличчя до Аммонових синів, і пророкуй на них.
EZEK|25|3|І скажеш Аммоновим синам: Послухайте слова Господа Бога: Так говорить Господь Бог: За те, що ти говориш Ага! про Мою святиню, бо вона збезчещена, і про Ізраїлеву землю, бо спустошена, і про Юдин дім, бо пішов у полон,
EZEK|25|4|тому ось Я дам тебе синам сходу на спадок, і поставлять вони в тебе шатра свої, і зроблять у тебе місця свого пробування. Вони будуть їсти твій плід, і вони будуть пити твоє молоко.
EZEK|25|5|І дам я Раббу на стайню для верблюдів, а Аммонових синів на лігво отари, і ви пізнаєте, що Я Господь!
EZEK|25|6|Бо так Господь Бог промовляє: За твоє плескання рукою, і твоє тупотіння ногою, і що в душі тішишся ти всією своєю погордою до Ізраїлевої землі,
EZEK|25|7|тому ось Я витягну Свою руку на тебе, і дам тебе на здобич для народів, і витну тебе з народів, і вигублю тебе з країв, знищу тебе, і пізнаєш, що Я Господь!
EZEK|25|8|Так сказав Господь Бог: За те, що Моав та Сеїр говорять: Ось Юдин дім як усі народи,
EZEK|25|9|тому ось Я відкрию Моавове збіччя від міст, від його міст, від його кінця, пишноту землі: Бен-Гаєшімот, Баал-Меон аж до Кір'ятаїму.
EZEK|25|10|Я дам його на спадок для синів сходу разом з синами Аммоновими, щоб не згадувались Аммонові сини серед народів.
EZEK|25|11|А над Моавом зроблю присуди, і пізнають вони, що Я Господь!
EZEK|25|12|Так говорить Господь Бог: За те, що Едом мстився мстою над Юдиним домом, і тяжко грішили, через те, що мстилися над ними,
EZEK|25|13|тому так говорить Господь Бог: І витягну Я руку Свою на Едома, і витну з нього людину й скотину, і вчиню його руїною, від Теману й аж до Дедану вони попадають від меча!
EZEK|25|14|І дам Я Свою помсту над Едомом у руку Мого народу Ізраїля, і вчиню в Едомі за гнівом Своїм, за лютістю Своєю, і зазнають вони Моєї помсти, говорить Господь Бог!
EZEK|25|15|Так говорить Господь Бог: За те, що филистимляни чинили в помсті, і мстилися мстою через погорду в душі, щоб нищити в вічній ненависті,
EZEK|25|16|тому так говорить Господь Бог: Ось Я витягну Свою руку на филистимлян, і витну керетян, і вигублю останок морського берега,
EZEK|25|17|і вчиню над ними жорстокі помсти лютими карами. І пізнають вони, що Я Господь, коли Я вчиню Свою помсту серед них!
EZEK|26|1|І сталося одинадцятого року, першого дня місяця, було слово Господнє до мене таке:
EZEK|26|2|Сину людський, за те, що Тир говорить на Єрусалим: Ага! зламалися це двері народів, він звертається до мене, і я насичуся, бо він знищений,
EZEK|26|3|тому так говорить Господь Бог: Ось Я на тебе, Тире, і підійму на тебе багато народів, як море підіймає свої хвилі...
EZEK|26|4|І понищать вони мури Тиру, і повалять башти його, і вимету з нього порох його, і оберну його на голу скелю...
EZEK|26|5|Він буде серед моря місцем розтягнення неводу, бо Я сказав це, говорить Господь Бог, і стане він за здобич для народів,
EZEK|26|6|а його дочки, що на полі, будуть побиті мечем, і пізнають вони, що Я Господь!
EZEK|26|7|Бо так говорить Господь Бог: Ось Я спроваджу до Тиру Навуходоносора, вавилонського царя, з півночі, царя над царями, з конем і колесницею та з верхівцями, і з ними натовп, і численний народ.
EZEK|26|8|Він позабиває на полі дочок твоїх мечем, і зробить на тебе башту, і насипле на тебе вала, і поставить проти тебе щита...
EZEK|26|9|І дасть муролома на мури твої, і порозбиває мечами своїми він башти твої!
EZEK|26|10|Від надміру коней його закриє тебе їхня курява, від цокоту вершника, колеса та колесниці затремтять твої мури, як буде він входити в брами твої, як входять до міста з розламаним муром...
EZEK|26|11|Копитами коней своїх він потопче усі твої вулиці, позабиває мечем твій народ, і на землю попадають пам'ятники твоєї могутности...
EZEK|26|12|І вони розграбують багатство твоє, і пограбують товари твої, і порозвалюють мури твої, і порозбивають доми твої пишні, а каміння твоє, і дерева твої, і навіть твій порох вони поскидають у воду!...
EZEK|26|13|І Я припиню розлягання пісень твоїх, і бренькіт гусел твоїх більше чутий не буде...
EZEK|26|14|І зроблю тебе голою скелею, станеш місцем розтягнення сітки, і більше не будеш збудований, бо я, Господь, це сказав, Господь Бог промовляє!
EZEK|26|15|Отак Господь Бог промовляє до Тиру: Чи ж від шуму падіння твого, коли будуть стогнати ранені, коли забиватимуть посеред тебе, не затремтять острови?
EZEK|26|16|І всі князі моря посходять із тронів своїх, і поздіймають вони свої мантії, і постягають свої кольорові одежі, і зодягнуться страхом, посідають на землю, і будуть тремтіти щохвилі, і стовпом постають над тобою...
EZEK|26|17|І пісню жалобну про тебе вони заспівають, і скажуть тобі: Як загинуло ти, як одірване ти від морів, славне місто, що сильним на морі було, воно й його мешканці, що наводили страх свій на всіх його мешканців!
EZEK|26|18|Тепер затремтять острови в дні упадку твого, і жахнуться всі ті острови, що на морі, твоєю загубою...
EZEK|26|19|Бо так Господь Бог промовляє: Коли Я тебе оберну на спустошене місто, немов ті міста, що вони не замешкані, коли підійму Я безодню на тебе, і велика вода тебе вкриє,
EZEK|26|20|то знижу тебе разом з тими, що сходять в могилу, до предавнього люду, і в підземній землі осаджу я тебе, як руїни відвічні, із тими, що сходять в могилу, щоб ізнову ти не заселився, і в країні живих більш не жив!...
EZEK|26|21|За пострах тебе учиню, і не буде тебе, і будуть шукати тебе, та вже більше не знайдуть навіки, говорить оце Господь Бог!
EZEK|27|1|І було мені слово Господнє таке:
EZEK|27|2|А ти, сину людський, здійми пісню жалобну про Тир!
EZEK|27|3|І скажеш до Тиру: Ти, що при входах морських пробуваєш, що торгуєш з народами на численних островах: Так говорить Господь Бог: Тире, ти сказав: я то корона краси!
EZEK|27|4|У серці морів границі твої; будівничі твої довершили твою красу!
EZEK|27|5|З кипарису з Сеніру вони збудували для тебе всі дошки подвійні, взяли кедра з Ливану, щоб щоглу зробити на тобі.
EZEK|27|6|З башанських дубів твої весла зробили, твій поклад зробили із кости слонової, із смереки з островів тих Кіттійських.
EZEK|27|7|Сорокатий з Єгипту віссон був вітрилом твоїм, щоб за прапора бути тобі; блакить та пурпура з островів Еліші стали твоїм покриттям.
EZEK|27|8|Мешканці Сидону й Арваду були веслярами тобі, мудреці твої, Тире, у тебе були, вони мореплавці твої.
EZEK|27|9|Старші із Ґевалу й його мудреці були в тебе за тих, що латали проломи твої. Всі морські кораблі й мореплавці їхні в тебе були, щоб міняти крам твій.
EZEK|27|10|Перс, і Луд, і Пут були в війську твоїм вояками твоїми, вішали в тебе щита та шолома, вони то давали тобі пишноту.
EZEK|27|11|Синове Арваду та військо твоє навколо на мурах твоїх, а Ґаммадеї на баштах твоїх пробували, щити свої вішали навколо на мурах твоїх, вони довершили окрасу твою.
EZEK|27|12|Таршіш був для тебе купцем через многоту багатства усякого; сріблом, залізом, циною й оливом платили вони за крам твій.
EZEK|27|13|Яван, Тувал та Мешех це купці твої, людську душу та мідяні речі давали вони за замінний крам твій.
EZEK|27|14|З дому Тоґарми давали коні, і верхівців, і мулів за крам твій.
EZEK|27|15|Синове Дедану твої покупці; численні острови торгували з тобою, рогами слонової кости й гебановим деревом звертали данину твою.
EZEK|27|16|Арам твій купець через многість виробів твоїх; рубин, пурпуру, і квітчасту тканину, і віссон, і коралі та дорогоцінний камінь давали тобі за крам твій.
EZEK|27|17|Юда й Ізраїлів Край це купці твої; пшеницю з Мінніту, солодощі, і мед, і оливу й бальзам давали вони за замінний крам твій.
EZEK|27|18|Дамаск твій купець через многість виробів твоїх, через многість багатства усякого, вином із Хелбону та білою вовною.
EZEK|27|19|Ведан та Яван із Уззалу давали тобі за крам залізо оброблене, бальзам та очерет, було це замінним крамом твоїм.
EZEK|27|20|Дедан твій купець килимками до сідел при їждженні.
EZEK|27|21|Арабія та всі кедарські князі покупці це твоєї руки; ягнятами, і баранами, і козлами, ними торгівля твоя.
EZEK|27|22|Купці Шеви й Рами покупці це твої, коштовним бальзамом, і дорогим усіляким камінням та злотом давали вони за товар твій.
EZEK|27|23|Харан, і Ханне, і Еден, купці Шеви, Ашшур та Кілмад це твої покупці.
EZEK|27|24|Це твої покупці коштовним убранням: покривалами блакитними, і квітчастими, і багатокольоровими тканими виробами, міцними шнурами пов'язаними за крам твій.
EZEK|27|25|Кораблі із Таршішу твої каравани, для краму твого замінного, і став ти багатим, і став дуже славним у серці морів.
EZEK|27|26|На воду велику тебе завели твої веслярі, і в серці морів східній вітер розіб'є тебе.
EZEK|27|27|Багатство твоє та крам твій, і вироби твої замінні, мореплавці твої і твої щоглярі, ті, що латають пробої твої, і ті, що міняють замінний крам твій, і всі твої вояки, які в тебе, і всі збори твої, що серед тебе, попадають в серці морів в дні упадку твого!
EZEK|27|28|На лемент твоїх щоглярів затремтять вали морські,
EZEK|27|29|і посходять з своїх кораблів усі веслярі, мореплавці, всі морські щоглярі, на землі постають.
EZEK|27|30|І заголосять за тебе вони тужним голосом, і кричатимуть гірко, і свої голови порохом пообсипають, у попелі будуть качатись!
EZEK|27|31|І зроблять собі ради тебе жалобную лисину, і себе опережуть веретами, і плакатимуть за тобою в гіркоті душі гірким голосінням....
EZEK|27|32|І пісню жалоби сини їхні здіймуть про тебе, і над тобою співатимуть жалібно: Хто інший, як Тир, посередині моря зруйнований?
EZEK|27|33|Коли припливали вироби твої із морів, насищав ти численні народи; многотою багатства твого та виробів замінних твоїх ти збагачував земських царів!
EZEK|27|34|Тепер же, коли ти розбитий на морі, у водних глибинах, то замінний виріб твій і всі збори твої серед тебе попадали...
EZEK|27|35|Над тобою стовпіють усі остров'яни, а їхні царі затремтіли від жаху, засльозилися їхні обличчя!
EZEK|27|36|Купці серед народів глузливо свистять над тобою, ти пострахом став, і не буде навіки тебе!...
EZEK|28|1|І було мені слово Господнє таке:
EZEK|28|2|Сину людський, скажи князеві Тиру: Так говорить Господь Бог: за те, що повищилось серце твоє й ти сказав: Я Бог, сиджу на Божому престолі в серці морів, а ти тільки людина, а не Бог, хоч ставив своє серце нарівні з серцем Божим...
EZEK|28|3|Ось ти мудріший від Даниїла, кожен мудрець не прилучиться до тебе.
EZEK|28|4|Своєю мудрістю та своїм розумом набув ти собі багатство, і назгромадив золота та срібла в скарбницях своїх.
EZEK|28|5|Великою своєю мудрістю та торгівлею свою помножив ти багатство своє, і повищилось твоє серце багатством своїм!
EZEK|28|6|Тому так говорить Господь Бог: За те, що ти ставиш своє серце нарівні з серцем Божим,
EZEK|28|7|тому ось Я спроваджу на тебе чужих, насильників поміж народами, і вони повитягають мечі свої на красу твоєї мудрости, і зневажать красу твою.
EZEK|28|8|Вони скинуть тебе в могилу, і помреш ти смертю пробитого в серці морів.
EZEK|28|9|Чи справді ти скажеш: Я бог! перед убивником своїм, а ти ж тільки людина, а не Бог, у руці тих, що зневажають тебе?
EZEK|28|10|Ти помреш смертю необрізанців, від руки чужих, бо Я це сказав, говорить Господь Бог!
EZEK|28|11|І було мені слово Господнє таке:
EZEK|28|12|Сину людський, здійми жалобну пісню на тирського царя, та й скажеш йому: Так говорить Господь Бог: Ти печать досконалости, повен мудрости, і корона краси.
EZEK|28|13|Ти пробував ув Едені, садку Божому: усякий дорогий камінь на одежі твоїй: карнеоль, топаз і яспіс, хризоліт, согам, і онікс, сапфір, рубін і смарагд, і золото; знаряддя бубнів твоїх та сопілок твоїх були в тебе що дня, коли був ти створений, були вони наготовлені.
EZEK|28|14|Ти помазаний Херувим хоронитель, і Я дав тебе на святу гору Божу, ти ходив посеред огнистого каміння.
EZEK|28|15|Ти був бездоганний у своїх дорогах від дня твого створення, аж поки не знайшлася на тобі несправедливість.
EZEK|28|16|Через велику торгівлю твою твоє нутро переповнилось насиллям, і ти прогрішив. Тому Я зневажив тебе, щоб не був ти на Божій горі, і погубив тебе, хоронителю Херувиме, з середини огнистого каміння.
EZEK|28|17|Стало високим твоє серце через красу твою, ти занапастив свою мудрість через свою красу. Кинув Я тебе на землю, дав тебе перед царями, щоб дивились на тебе.
EZEK|28|18|Многотою провин своїх, через кривду торгівлі своєї зневажив ти святині свої. І вивів Я огонь з твоєї середини, і він пожер тебе, і Я зробив тебе попелом на землі на очах усіх, хто бачить тебе.
EZEK|28|19|Усі, хто знає тебе серед народів, остовпіють над тобою; ти пострахом станеш, і не буде тебе аж навіки!...
EZEK|28|20|І було мені слово Господнє таке:
EZEK|28|21|Сину людський, зверни своє обличчя до Сидону, і пророкуй на нього,
EZEK|28|22|та й скажеш: так говорить Господь Бог: Ось Я на тебе, Сидоне, і буду шанований серед тебе, і пізнають, що Я Господь, коли робитиму на нього присуди, і коли покажу Свою святість серед нього.
EZEK|28|23|І пошлю на нього моровицю та кров на його вулиці, і впаде серед нього пробитий, що прийде на нього знавкола, і пізнають, що Я Господь.
EZEK|28|24|І не буде вже для Ізраїлевого дому колючої тернини та будяччя, що приносить біль зо всіх їхніх околиць, що погорджують ними, і пізнають вони, що Я Господь Бог.
EZEK|28|25|Так говорить Господь Бог: Коли Я позбираю Ізраїлів дім із народів, між якими вони розпорошені, то Я покажу на ньому Свою святість на очах народів, і вони осядуть на землі своїй, яку Я дав Своєму рабові Якову.
EZEK|28|26|І осядуть вони на ній безпечно, і будуватимуть доми та садитимуть виноградники, і будуть сидіти безпечно, коли Я чинитиму присуди на всіх тих, що погорджують ними з їхнього довкілля. І пізнають вони, що Я Господь, їхній Бог!
EZEK|29|1|За десятого року, десятого місяця, дванадцятого дня місяця, було мені слово Господнє таке:
EZEK|29|2|Сину людський, зверни своє обличчя до фараона, єгипетського царя, і пророкуй на нього та на ввесь Єгипет.
EZEK|29|3|Говори та й скажеш: Так говорить Господь Бог: Ось Я на тебе, фараоне, царю єгипетський, крокодиле великий, що лежиш серед своїх рік, що говориш: Моя річка моя, і я утворив її для себе!
EZEK|29|4|І вкладу гачки в щелепи твої, і поприліплюю рибу твоїх річок до твоєї луски, і підійму тебе з середини твоїх річок, і всі риби твоїх річок поприліплюються до твоєї луски!
EZEK|29|5|І вирву тебе й кину в пустиню, тебе та всі риби річок твоїх; ти впадеш на поверхні поля, не будеш згромаджений і не будеш позбираний, для земної звірини та для птаства небесного дам Я на їжу тебе...
EZEK|29|6|І пізнають усі мешканці Єгипту, що Я Господь, бо вони були для Ізраїлевого дому очеретяною палицею.
EZEK|29|7|Коли вони хапались за тебе долонею, ти ламався й роздирав їм усе рамено; а коли вони опиралися на тебе, ти ламався й чинив, що їм тряслися всі стегна.
EZEK|29|8|Тому так говорить Господь Бог: Ось Я наведу на тебе меча, і витну з-між тебе людину й скотину.
EZEK|29|9|І стане єгипетський край спустошенням та руїною, і пізнають вони, що Я Господь, за те, що він говорив: Річка моя, і то я її утворив!
EZEK|29|10|Тому ось Я проти тебе та проти річок твоїх, і оберну єгипетський край на поруйновані руїни, на спустошення від Міґдолу аж до Севене, і аж до границі Етіопії,
EZEK|29|11|не перейде по ньому нога людська, і нога звірини не перейде по ньому, і не буде він замешканий сорок років...
EZEK|29|12|І оберну Я єгипетський край на спустошення серед спустошених країв, а його міста серед поруйнованих міст будуть спустошенням сорок років, і розпорошу Єгипет серед народів, і порозсипаю їх по краях...
EZEK|29|13|Бо так говорить Господь Бог: Наприкінці сорока років позбираю Єгипет з-між народів, де вони були розпорошені.
EZEK|29|14|І верну долю Єгипту, і верну їх до краю Патрос, до краю їхнього походження, і вони будуть там царством слабим.
EZEK|29|15|З-поміж царств воно буде найнижче, і не підійметься вже понад народами, і поменшу їх, щоб не панували над народами.
EZEK|29|16|І не буде вже воно для Ізраїлевого дому надією, яка пригадувала б беззаконня, коли вони, зверталися до нього. І пізнають вони що Я Господь Бог!
EZEK|29|17|І сталося за двадцятого й сьомого року, першого місяця, першого дня місяця, було мені слово Господнє таке:
EZEK|29|18|Сину людський, Навуходоносор, цар вавилонський, змусив своє військо робити велику працю проти Тиру. Кожна голова вилисіла, і всяке рамено витерте, та нема нагороди ані йому, ані війську його від Тиру за ту працю, яку він робив проти нього.
EZEK|29|19|Тому так говорить Господь Бог: Ось Я дам Навуходоносорові, цареві вавилонському, єгипетську землю, і він забере багатство її, і ограбує грабунком її, і забере її здобиччю, і вона стане нагородою для війська його.
EZEK|29|20|За працю його, яку він робив у ній, Я даю йому єгипетську землю, бо вони це зробили Мені, говорить Господь Бог.
EZEK|29|21|Того дня вирощу рога Ізраїлевому домові, а тобі відкрию уста серед них. І вони пізнають, що Я Господь.
EZEK|30|1|І було мені слово Господнє таке:
EZEK|30|2|Сину людський, пророкуй, і скажеш: Так говорить Господь Бог: Голосіть Ой! цього дня!
EZEK|30|3|Бо близький день, і близький день Господній, день хмарний, настає час народів!
EZEK|30|4|І прийде меч на Єгипет, і буде тремтіння в Етіопії, коли будуть падати забиті в Єгипті, і заберуть багатство його, і будуть розбиті основи його.
EZEK|30|5|Куш, і Пут, і Луд, і ввесь помішаний народ, і Кув, і сини землі заповіту попадають з ними від меча.
EZEK|30|6|Так говорить Господь: І попадають підпори Єгипту, і так упаде гординя сили його, від Міґдолу аж до Севене, від меча попадають у ньому, говорить Господь Бог.
EZEK|30|7|І буде він спустошений серед попустошених країв, а міста його будуть серед міст поруйнованих.
EZEK|30|8|І пізнають вони, що Я Господь, коли Я дам огонь на Єгипет, і будуть поторощені всі, хто йому помагає.
EZEK|30|9|Того дня повиходять посланці з-перед Мого лиця на кораблях, щоб налякати безпечну Етіопію, і буде через них жах, як у день Єгипту, бо це ось надходить!
EZEK|30|10|Так говорить Господь Бог: І Я зроблю кінець єгипетському многолюдству рукою Навуходоносора, вавилонського царя.
EZEK|30|11|Він та народ його з ним, насильники людів, будуть спроваджені знищити землю, і вони повитягують мечі свої на Єгипет, і наповнять край побитими!
EZEK|30|12|І оберну Я річки на суходіл, і передам землю в руку злочинців, і спустошу край та все, що в ньому, рукою чужих. Я, Господь, це сказав!
EZEK|30|13|Так говорить Господь Бог: І повигублюю божків, і зроблю кінець бовванам з Нофу, і не буде вже князів в єгипетському краї, і дам пострах на єгипетську землю.
EZEK|30|14|І Патрос спустошу, і дам огонь у Цоан, і буду виконувати присуди в Но.
EZEK|30|15|І виллю Я гнів Свій на Сіна, твердиню єгипетську, і витну многолюдство Но.
EZEK|30|16|І пошлю Я огонь на Єгипет, сильно буде корчитись Сін, а Но буде проламаний, а на Ноф нападуть вороги вдень.
EZEK|30|17|Юнаки Авену та Пі-Весету попадають від меча, а інші підуть у полон.
EZEK|30|18|А в Тахпанхесі потемніє день, коли Я ламатиму там єгипетські ярма, і скінчиться в ньому пиха сили його. Самого його хмара закриє, а його дочки підуть у полон...
EZEK|30|19|І буду виконувати присуди над Єгиптом, і вони пізнають, що Я Господь!
EZEK|30|20|І сталося, за одинадцятого року, першого місяця, сьомого дня місяця, було мені слово Господнє таке:
EZEK|30|21|Сину людський, Я зламав рамено фараона, єгипетського царя, і ось воно не буде перев'язане, щоб дати ліки, щоб покласти пов'язку, щоб обвинути його, і щоб зміцнити його вхопитися за меча.
EZEK|30|22|Тому так говорить Господь Бог: Ось Я на фараона, єгипетського царя, і поламаю рамена його, те дуже та те зламане, і викину меча з його руки.
EZEK|30|23|І розпорошу Єгипет серед народів, і порозсипаю їх по краях.
EZEK|30|24|І зміцню рамена вавилонського царя, і дам меча Свого в його руку, і зламаю Я фараонові рамена, і він буде стогнати стогоном проколеного перед ним.
EZEK|30|25|І зміцню Я рамена вавилонського царя, а фараонові рамена опадуть. І пізнають вони, що Я Господь, коли Я дам Свого меча в руку вавилонського царя, і простягну його на єгипетську землю.
EZEK|30|26|І розпорошу Єгипет серед народів, і порозсипаю їх по краях. І пізнають вони, що Я Господь!
EZEK|31|1|І сталося за одинадцятого року, третього місяця, першого дня місяця, було мені слово Господнє таке:
EZEK|31|2|Сину людський, скажи фараонові, цареві єгипетському, та до його многолюдства: До кого ти вподоблюєшся в своїй величі?
EZEK|31|3|Ось Ашшур, кедр на Ливані, з прекрасними галузками, з тінистою гущавиною, і високорослий, і аж між хмарами буде верховіття його.
EZEK|31|4|Води його виховали, безодня його викохала, він річки свої попровадив навколо свого насадження, а канали свої посилав до всіх дерев польових.
EZEK|31|5|Тому його зріст став вищий від усіх польових дерев, і помножилися галузки його, і від великої води його віття повидовжувалось, коли вигнався він.
EZEK|31|6|В його віттях кублилося все птаство небесне, а під його галузками родилася всяка польова звірина, а в його тіні сиділи всі численні народи.
EZEK|31|7|І був він уродливий висотою свого зросту, довготою галузок своїх, бо його корінь був при великих водах.
EZEK|31|8|Кедри в Божому садку не були рівні йому, кипариси не були подібні до галузок його, а платани не були, як його віття. Жодне дерево в Божому садку не було подібне до нього красою своєю!
EZEK|31|9|Я оздобив його ряснотою галузок його, і йому заздрили всі еденські дерева, що в Божому садку.
EZEK|31|10|Тому так сказав Господь Бог: За те, що ти повищився зростом, і дав верховіття своє аж між хмари, і повищилося серце його, коли він став високим,
EZEK|31|11|то дай його в руку сильного з народів, він конче зробить йому за його беззаконня, за це Я вигнав його!
EZEK|31|12|І витяли його чужі, насильники народів, і повідкидали його. На гори й на всі долини попадали галузки його, і було поламане віття його по всіх потоках землі, а всі народи землі повиходили з тіні його й покинули його.
EZEK|31|13|Над його руїнами пробувало все небесне птаство, а при галуззях його була всяка польова звірина,
EZEK|31|14|щоб не повищувалися своїм зростом усі дерева при воді, і не давали свого верховіття поміж хмари, і не ставали у своїй величі сильні між ними, що п'ють воду, бо всі вони віддані смерті до підземного краю серед людських синів, до тих, хто сходить до могили.
EZEK|31|15|Так говорить Господь Бог: Того дня, коли він зійшов до шеолу, учинив Я жалобу, закрив над ними безодню, затримав його річки, і була стримана велика вода, і затемнив над ним Лівана, а всі польові дерева помліли над ним.
EZEK|31|16|Від гуку упадку його Я вчинив тремтячими народи, коли Я знизив його до шеолу з тими, що сходять до гробу. І потішилися в підземному краї всі еденські дерева, добірне та добре Ливанське, всі, що п'ють воду.
EZEK|31|17|Також вони зійшли з ними до шеолу, до побитих мечем, що сиділи, як його помічники, в його тіні серед народів.
EZEK|31|18|До кого став ти так подібний у славі та в великості серед еденських дерев? І будеш ти знижений з еденськими деревами до підземного краю, посеред необрізанців будеш лежати з пробитими мечем. Це фараон та все многолюдство його, говорить Господь Бог.
EZEK|32|1|І сталося за дванадцятого року, дванадцятого місяця, третього дня місяця, було мені слово Господнє таке:
EZEK|32|2|Сину людський, здійми пісню жалобную на фараона, єгипетського царя, та й скажеш йому: Левчукові з народів подібний ти був, а тепер ти мов морська потвора, виприскуєш воду по ріках своїх, і скаламучуєш воду ногами своїми, болотиш ти їхні річки!
EZEK|32|3|Отак Господь Бог промовляє: Але сітку Свою розтягну Я на тебе через збори численних народів, і тебе Своїм неводом витягну!
EZEK|32|4|І викину зразу на землю тебе, і кину тебе Я на поле широке, і над тобою спочине всяке птаство небесне, і тобою насичу звірину всієї землі...
EZEK|32|5|І дам твоє м'ясо на гори, а трупом твоїм Я долини наповню...
EZEK|32|6|І землю, де пливаєш ти, аж до гір напою її кров'ю твоєю, тобою наповняться річища...
EZEK|32|7|А коли Я тебе погашу, то небо закрию, а зорі його позатемнюю, сонце хмарою вкрию його, а місяць не буде світити свого світла...
EZEK|32|8|Всі світила, що світять на небі, позатемнюю їх над тобою, і дам темноту понад краєм твоїм, говорить Господь Бог!
EZEK|32|9|І занепокою Я серце численних народів, коли вість рознесу про руїну твою між народами аж до країв, яких ти не знав.
EZEK|32|10|І остовпіють численні народи з-за тебе, а їхні царі затремтять через тебе в страху, як буду махати мечем Своїм Я перед їхнім обличчям, і тремтітиме кожен щохвилі за душу свою в дні упадку твого...
EZEK|32|11|Бо так Господь Бог промовляє: Меч царя вавилонського прийде на тебе!
EZEK|32|12|Мечами хоробрих Я порозкидаю твоє многолюдство. Усі вони насильники народів, і гордість Єгипту понищать вони, і все многолюдство його буде вигублене...
EZEK|32|13|І вигублю ввесь його скот при водах великих, і не буде вже їх каламутити людська нога, і копито скотини не буде вже їх каламутити.
EZEK|32|14|Тоді їхні води очищу, а їхні річки попроваджу, неначе оливу, говорить Господь Бог.
EZEK|32|15|Коли оберну Я єгипетський край на спустошення, і край опустошений буде від усього, що в нім, коли Я поб'ю всіх тих, що замешкують в ньому, то пізнають вони, що Я то Господь!...
EZEK|32|16|Оце пісня жалобна, і будуть жалобно співати її, дочки народів будуть співати жалобно її, про Єгипет та про все многолюдство його будуть жалобно співати її, говорить Господь Бог.
EZEK|32|17|І сталося за дванадцятого року, п'ятнадцятого дня місяця, було мені слово Господнє таке:
EZEK|32|18|Сину людський, жалобно заголоси про многолюдство Єгипту, і скинь його, його та дочок потужних народів до підземного краю із тими, хто сходить в могилу!
EZEK|32|19|Від кого ти став приємніший? Зійди й покладись з необрізанцями!
EZEK|32|20|Попадають серед пробитих мечем, меч даний на те, із ним ляжуть його всі народи...
EZEK|32|21|Будуть йому говорити сильніші з хоробрих з-посеред шеолу із помічниками: Посходили, полягали ці необрізанці, побиті мечем:
EZEK|32|22|Там Ашшур і всі збори його, навколо нього гроби його, всі побиті вони, від меча всі попадали,
EZEK|32|23|що були його гроби найглибше в могилі, і був його полк біля гробу його, всі побиті вони, від меча всі попадали, що ширили жах по краю живих...
EZEK|32|24|Там Елам та ввесь натовп його коло гробу його, всі побиті вони, від меча всі попадали, що зійшли необрізанцями до підземного краю, що ширили жах свій по краю живих, і понесли ганьбу свою з тими, хто сходить в могилу...
EZEK|32|25|Дали йому ложе посеред побитих зо всім многолюдством його, гроби його коло нього, всі вони необрізанці, побиті мечем, бо ширили жах свій по краю живих і понесли ганьбу свою з тими, хто сходить в могилу, посеред побитих покладений він...
EZEK|32|26|Там Мешех, Тувал та все многолюдство його, гроби його коло нього, всі вони необрізанці, побиті мечем, бо ширили жах свій по краю живих...
EZEK|32|27|І не будуть лежати із лицарями, що попадали із необрізанців, що зійшли до шеолу з військовим знаряддям своїм, і поклали свої мечі під свої голови, і їхня провина на їхніх костях, бо жах перед лицарями був у краї живих,
EZEK|32|28|а ти розпорошений між необрізанцями, і поляжеш із тими, хто побитий мечем...
EZEK|32|29|Там Едом, і царі його, і князі всі його, що при всій своїй силі були зложені з побитими мечами, вони ляжуть з необрізанцями та з тими, хто сходить в могилу...
EZEK|32|30|Там північні князі, всі вони й всі сидоняни, що посходили разом з побитими, хоч був жах від їхньої міці, були посоромлені, і полягали вони, необрізанці, з побитими мечем, і свою ганьбу понесли із тими, хто сходить в могилу...
EZEK|32|31|Фараон їх побачить, і потішиться всім многолюдством своїм, мечем побитий фараон та все його військо, говорить Господь Бог!...
EZEK|32|32|Бо поширю Я жах Свій на землю живих, і буде покладений серед необрізанців з побитими мечем фараон та усе многолюдство його, говорить Господь Бог!
EZEK|33|1|І було мені слово Господнє таке:
EZEK|33|2|Сину людський, говори синам свого народу, та й скажеш до них: Коли б Я спровадив на який край меча, і взяв би народ цього краю одного чоловіка з-поміж себе, і поставив би його собі вартовим,
EZEK|33|3|і коли б він побачив меча, що йде на цей край, і засурмив би в сурму, й остеріг народ,
EZEK|33|4|і почув би хто голос сурми, та не був би обережний, і прийшов би меч та й захопив би його, то кров його на голові його буде!
EZEK|33|5|Голос сурми він чув, та не був обережний, кров його буде на ньому, а він, коли б був обережний, урятував би свою душу.
EZEK|33|6|А той вартовий, коли б побачив меча, що йде, і не засурмив би в сурму, а народ не був би обережний, і прийшов би меч, і захопив би одного з них, то він був би узятий за гріх свій, а його кров Я зажадаю з руки вартового.
EZEK|33|7|А ти, сину людський, Я дав тебе вартовим для Ізраїлевого дому, і ти почуєш з уст Моїх слово, й остережеш їх від Мене.
EZEK|33|8|Коли б Я сказав до безбожного: Безбожнику, ти конче помреш!, а ти не говорив би, щоб остерегти безбожного від дороги його, то він, несправедливий, помре за свій гріх, а його кров Я вимагатиму з твоєї руки.
EZEK|33|9|А ти, коли остережеш несправедливого від дороги його, щоб вернувся з неї, і він не вернеться з своєї дороги, він помре за гріх свій, а ти душу свою врятував.
EZEK|33|10|А ти, сину людський, скажи до Ізраїлевого дому: Ви кажете так, говорячи: Коли наші провини та наші гріхи на нас, і через них ми гинемо, то як будемо жити?
EZEK|33|11|Скажи їм Як живий Я, говорить Господь Бог, не прагну смерти несправедливого, а тільки щоб вернути несправедливого з дороги його, і буде він жити! Наверніться, наверніться з ваших злих доріг, і нащо вам умирати, доме Ізраїлів?
EZEK|33|12|А ти, сину людський, скажи до синів свого народу: Справедливість справедливого не врятує його в дні гріха його, а несправедливість несправедливого не спіткнеться він об неї в дні навернення від своєї несправедливости, а справедливий не зможе жити в ній в дні свого гріха.
EZEK|33|13|Коли Я скажу справедливому: Буде конче він жити, а він надіявся б на свою справедливість, та робив би кривду, то вся його справедливість не буде згадана, і за кривду свою, що зробив, він помре!
EZEK|33|14|А коли Я скажу до несправедливого: Конче помреш ти, а він навернеться від свого гріха, і робитиме право та справедливість:
EZEK|33|15|заставу поверне несправедливий, грабунок відшкодує, ходитиме уставами життя, щоб не чинити кривди, то конче буде він жити, не помре!
EZEK|33|16|Усі гріхи його, які він нагрішив, не будуть йому згадані, право та справедливість робив він, конче буде він жити!
EZEK|33|17|І кажуть сини твого народу: Несправедлива Господня дорога! тоді як несправедлива їхня власна дорога.
EZEK|33|18|Коли справедливий відвернеться від своєї справедливости, і робитиме кривду, то помре він за те!
EZEK|33|19|А коли несправедливий відвернеться від своєї несправедливости, і чинитиме право та справедливість, то на них він буде жити!
EZEK|33|20|А ви кажете: Несправедлива Господня дорога! Кожного з вас Я буду судити, Ізраїлів доме, за його дорогами!
EZEK|33|21|І сталося за дванадцятого року, десятого місяця, п'ятого дня місяця від нашого вигнання, прийшов був до мене втікач з Єрусалиму, говорячи: Побите це місто!...
EZEK|33|22|А Господня рука була прийшла до мене ввечорі перед приходом цього втікача, і Він відкрив мої уста, поки прийшов той до мене вранці. І були відкриті мої уста, і не був уже я більше німий!
EZEK|33|23|І було мені слово Господнє таке:
EZEK|33|24|Сину людський, мешканці цих руїн на Ізраїлевій землі говорять так: Авраам був один, та проте посів цей Край, а нас багато, нам даний цей Край на спадщину!
EZEK|33|25|Тому скажи їм: Так сказав Господь Бог: Ви на крові їсте, а свої очі зводите до бовванів своїх, і кров проливаєте, і цей Край посядете ви?
EZEK|33|26|Ви спираєтесь на свого меча, робите гидоту, і кожен безчестить жінку свого ближнього, і цей Край посядете ви?
EZEK|33|27|Так скажеш до них: Так говорить Господь Бог: Як живий Я, ті, хто в руїнах, попадають від меча, а той, хто на широкім полі, того віддам звірині, щоб пожерла його, а ті, хто в твердинях та в печерах, помруть від моровиці!
EZEK|33|28|І оберну Я цей Край на спустошення та на сплюндрування, і скінчиться пиха сили його, і опустошіють Ізраїлеві гори, так що не буде й перехожого...
EZEK|33|29|І пізнають вони, що Я Господь, коли Я оберну цей Край на спустошення та на сплюндрування за всі їхні гидоти, що зробили вони.
EZEK|33|30|А ти, сину людський, сини твого народу умовляються про тебе при стінах і в дверях домів, і говорять один з одним, кожен зо своїм братом, кажучи: Увійдіть та послухайте, що це за слово, що виходить від Господа?
EZEK|33|31|І прийдуть до тебе, як приходить народ, і сядуть перед тобою як Мій народ, і послухають твоїх слів, але їх не виконають, бо що приємне в устах їхніх, те вони зроблять, а серце їхнє ходить за захланністю їхньою.
EZEK|33|32|І ось ти для них, як пісня кохання, красноголосий і добрий грач, і вони слухають слова твої, але їх не виконують!
EZEK|33|33|А коли оце прийде, ось воно вже приходить! то пізнають вони, що серед них був пророк.
EZEK|34|1|І було мені слово Господнє таке:
EZEK|34|2|Сину людський, пророкуй на Ізраїлевих пастирів, пророкуй та й скажеш до них, до тих пастирів: Так говорить Господь Бог: Горе Ізраїлевим пастирям, які пасуть самих себе! Хіба ж не отару повинні пасти пастирі?
EZEK|34|3|Жир ви їсте, та вовну вдягаєте, ситу вівцю ріжете, але отари не пасете!
EZEK|34|4|Слабих не зміцняєте, а хворої не лікуєте, і пораненої не перев'язуєте, сполошеної не вертаєте, і загинулої не шукаєте, але пануєте над ними силою та жорстокістю!
EZEK|34|5|І порозпорошувалися вони з браку пастиря, і стали за їжу для всякої польової звірини, і порозбігалися...
EZEK|34|6|Блукає отара Моя по всіх горах та по всіх високих згір'ях, і по всій широкій землі розпорошена отара Моя, і немає нікого, хто турбувався б про них, і немає нікого, хто б їх шукав!...
EZEK|34|7|Тому, пастирі, послухайте слова Господнього:
EZEK|34|8|Як живий Я, говорить Господь Бог, за те, що отара Моя полишена на здобич, і стала отара Моя за їжу для всякої польової звірини через брак пастиря, і пастирі Мої не шукають Моєї отари, а себе самих пасуть пастирі Мої, а отари Моєї не пасуть,
EZEK|34|9|тому, пастирі, послухайте слова Господнього:
EZEK|34|10|Так говорить Господь Бог: Ось Я на тих пастирів, і зажадаю з їхньої руки отари Моєї, і відірву їх від пасіння отари, і ті пастирі не будуть уже пасти самих себе, й Я врятую Свою отару з їхніх уст, і вони не будуть їм за їжу.
EZEK|34|11|Бо так Господь Бог промовляє: Ось Я Сам, і зажадаю отару Мою, і перегляну їх.
EZEK|34|12|Як пастух переглядає своє стадо того дня, коли він серед своєї розпорошеної отари, так Я перегляну отару Свою, і вирятую їх зо всіх тих місць, куди вони були розпорошені за хмарного та імлистого дня.
EZEK|34|13|І випроваджу їх від народів, і позбираю їх із країв, і приведу їх до їхньої землі, і буду їх пасти на Ізраїлевих горах, при річищах та по всіх оселях Краю.
EZEK|34|14|На пасовищі доброму пастиму їх, і на високих Ізраїлевих горах буде їхній випас, там вони будуть лежати на випасі доброму, і випасатимуть сите пасовище на Ізраїлевих горах!
EZEK|34|15|Я буду пасти отару Свою, і Я їх покладу на спочинок, говорить Господь Бог.
EZEK|34|16|Загинулу вівцю відшукаю, а сполошену поверну, а поранену перев'яжу, а хвору зміцню, а ситу та сильну погублю, буду пасти її правосуддям!
EZEK|34|17|А ви, отаро Моя, так говорить Господь Бог: Ось Я буду судити між вівцею й вівцею, між бараном і козлами.
EZEK|34|18|Чи мало вам того, що ви спасуєте хороше пасовище, а решту ваших пасовищ ви топчете своїми ногами? І воду чисту ви п'єте, а позосталу ногами своїми каламутите?
EZEK|34|19|І отара Моя мусить випасати потоптане вашими ногами, і пити скаламучене вашими ногами!
EZEK|34|20|Тому так Господь Бог промовляє до них: Ось Я Сам і розсуджу між вівцею ситою й між вівцею худою.
EZEK|34|21|За те, що ви боком і раменом попихаєте, і рогами вашими колете всіх слабих, аж поки не порозпорошуєте їх геть,
EZEK|34|22|то Я спасу отару Свою, і вона не буде вже за здобич, і Я розсуджу між вівцею та вівцею!
EZEK|34|23|І поставлю над ними одного пастиря, і він буде їх пасти, раба Мого Давида, він їх буде пасти, і він їм буде за пастиря!
EZEK|34|24|А Я, Господь, буду їм Богом, а раб Мій Давид князем серед них. Я, Господь, це сказав!
EZEK|34|25|І складу Я з ними заповіта миру, і прикінчу на землі злу звірину, і вони пробуватимуть в пустині безпечно, і будуть спати по лісах.
EZEK|34|26|І вчиню їх та довкілля Мого взгір'я благословенням, і спущу дощ в його часі, будуть це дощі благословенні.
EZEK|34|27|І польове дерево видасть свій плід, а земля видасть свій урожай, і будуть вони безпечні на своїй землі, і пізнають, що Я Господь, коли зламаю занози їхнього ярма, і врятую їх від руки тих, хто їх поневолив.
EZEK|34|28|І не будуть уже вони за здобич для народів, і звірина земна не жертиме їх, і будуть вони сидіти безпечно, і не буде нікого, хто б їх настрашив.
EZEK|34|29|І викохаю їм саджанця на славу, і не будуть вони вже забрані голодом із землі, і не понесуть уже ганьби народів.
EZEK|34|30|І пізнають вони, що Я Господь, Бог їхній, з ними, а вони народ Мій, дім Ізраїлів, говорить Господь Бог.
EZEK|34|31|А ви отара Моя, отара Мого випасу, ви люди, а Я Бог ваш, говорить Господь Бог.
EZEK|35|1|І було мені слово Господнє таке:
EZEK|35|2|Сину людський, зверни своє обличчя до гори Сеїр, і пророкуй на неї
EZEK|35|3|та й скажеш їй: Так говорить Господь Бог: Ось Я на тебе, горо Сеїре, і витягну руку Свою на тебе, й оберну тебе на спустошення та на сплюндрування.
EZEK|35|4|Міста твої оберну на руїну, а ти будеш спустошенням, і пізнаєте ви, що Я Господь!
EZEK|35|5|За те, що ти маєш вічну ворожнечу, і валила Ізраїлевих синів через меча в часі їхнього нещастя, в часі загибелі кінцевої,
EZEK|35|6|тому як живий Я, говорить Господь Бог, на кров оберну тебе, і кров буде гнати тебе. Отож кров ти зненавиділа, то кров буде гнати тебе!
EZEK|35|7|Оберну Я гору Сеїр на спустошення та на сплюндрування, і витну з неї того, хто йде та вертається.
EZEK|35|8|І наповню його гори трупами його! Згір'я твої й долини твої та всі твої річища, побиті мечем попадають у них!
EZEK|35|9|На вічні руїни оберну Я тебе, а міста твої не заселяться, і пізнаєте ви, що Я Господь!
EZEK|35|10|За те, що ти кажеш: Два ці народи, і два ці краї будуть мої, і ми посядемо те, де Господь був,
EZEK|35|11|тому, як живий Я, говорить Господь Бог, зроблю Я за гнівом твоїм та за заздрістю твоєю, які ти робив із своєї ненависти до них, і вони пізнають Мене, коли буду судити тебе.
EZEK|35|12|І пізнаєш ти, що Я Господь, чув усі образи твої, які ти казав на Ізраїлеві гори, говорячи: Вони опустошілі, дані нам на їжу!
EZEK|35|13|І ви величалися проти Мене своїми устами, і збільшували проти Мене слова свої, Я це чув!
EZEK|35|14|Так говорить Господь Бог: Коли буде радіти вся земля, тоді вчиню її тобі спустошенням!
EZEK|35|15|Як радієш ти зо спадку Ізраїлевого дому через те, що опустошіло воно, так зроблю Я й тобі. Спустошенням станеш, горо Сеїре, та ввесь Едом, увесь він, і пізнають вони, що Я Господь!
EZEK|36|1|А ти, сину людський, пророкуй на Ізраїлеві гори, та й скажеш: Ізраїлеві гори, послухайте слова Господнього!
EZEK|36|2|Так говорить Господь Бог: За те, що ворог говорить на вас Ага! і вічні пагірки стали вам за спадщину,
EZEK|36|3|тому пророкуй та й скажеш: Так говорить Господь Бог: За те, що пустошено й топтано вас знавкола, щоб були ви спадком для останку народів, і були ви взяті на кінчик язика й на балаканину народу,
EZEK|36|4|тому, Ізраїлеві гори, послухайте слова Господа Бога: Так говорить Господь Бог до гір та до згір'їв, до річищ та до долин, і до спустошілих руїн, і до опущених міст, що стали за здобич та за посміховисько для решти тих народів, що навколо.
EZEK|36|5|Так говорить Господь Бог: Поправді кажу, що огнем Своєї ревности говорив Я на решту тих народів та на ввесь Едом, що взяли собі Мій Край за спадок у радості всього серця, у погорді душі, щоб вигнати його на здобич.
EZEK|36|6|Тому пророкуй на Ізраїлеву землю, та й скажеш до гір, до згір'їв, до річищ та до долин: Так говорить Господь Бог: Ось Я говорив у ревності Своїй та в гніві Своїм за те, що ви носили ганьбу народів.
EZEK|36|7|Тому так говорить Господь Бог: Прирікаючи, Я підняв Свою руку, що ті люди, які навколо вас, вони понесуть свою ганьбу!
EZEK|36|8|А ви, Ізраїлеві гори, розпустіть ваше віття, і будете приносити плід свій для Мого народу Ізраїля, бо вони зблизилися, щоб прийти.
EZEK|36|9|Бо ось Я прийду до вас, і звернуся до вас, і ви будете оброблені та обсіяні.
EZEK|36|10|І розмножу на вас людину, увесь Ізраїлів дім, усього його, і будуть заселені ці міста, а руїни будуть забудовані.
EZEK|36|11|І розмножу на вас людину та скотину, і вони помножаться та розплодяться, і позаселюю вас, як за вашої давнини, і буду чинити вам краще, як за ваших початків, і ви пізнаєте, що Я Господь!
EZEK|36|12|І попроваджу на вас людину, мій народ Ізраїлів, і вони посядуть тебе, і станеш ти їм на спадок, і не будеш уже більше позбавляти їх дітей.
EZEK|36|13|Так говорить Господь Бог: За те, що говорять про вас: Ти їси людину, і позбавляєш народ свій дітей,
EZEK|36|14|тому ти не будеш уже їсти людини, і більше не позбавиш свій народ дітей, говорить Господь Бог!
EZEK|36|15|І не почуєш уже ти більше ганьби від поган, і наруги народів не будеш більше носити, і не вчиниш більше, щоб народ твій спотикався, говорить Господь Бог!
EZEK|36|16|І було мені слово Господнє таке:
EZEK|36|17|Сину людський, Ізраїлів дім вони жили на землі своїй, та й занечистили її своєю дорогою та своїми вчинками, як нечистість жінки в час нечистоти її стала їхня дорога перед Моїм лицем!
EZEK|36|18|І вилив Я гнів Свій на них за ту кров, яку вилили вони на землю, та бовванами своїми занечистили її.
EZEK|36|19|І розсіяв Я їх серед народів, і вони були розпорошені по країнах. За їхньою дорогою та за їхніми вчинками розсудив Я їх.
EZEK|36|20|І коли прийшли вони до тих народів, куди поприходили, то зневажили святе Моє Ймення, коли стали до них говорити: Вони народ Господа, та з землі Його повиходили!
EZEK|36|21|І змилувався Я над Своїм святим Ім'ям, що його зневажив Ізраїлів дім серед народів, куди вони поприходили.
EZEK|36|22|Тому скажи до Ізраїлевого дому: Так говорить Господь Бог: Не для вас Я роблю це, Ізраїлів доме, а тільки для святого Свого Ймення, яке ви зневажили серед народів, куди ви поприходили.
EZEK|36|23|І освячу Я велике Ім'я Своє, зневажене серед народів, що ви зневажили серед них, і пізнають ті люди, що Я Господь, говорить Господь Бог, коли Я покажу Свою святість серед вас на їхніх очах.
EZEK|36|24|І візьму вас із тих народів, і позбираю вас зо всіх країв, і приведу вас до вашої землі.
EZEK|36|25|І покроплю вас чистою водою, і станете чисті; зо всіх ваших нечистот і зо всіх ваших бовванів очищу вас.
EZEK|36|26|І дам вам нове серце, і нового духа дам у ваше нутро, і викину камінне серце з вашого тіла, і дам вам серце із плоті.
EZEK|36|27|І духа Свого дам Я до вашого нутра, і зроблю Я те, що уставами Моїми будете ходити, а постанови Мої будете стерегти та виконувати.
EZEK|36|28|І ви будете сидіти в Краю, якого Я дав вашим батькам, і будете Мені народом, а Я буду вам Богом!
EZEK|36|29|І спасу вас від усіх ваших нечистот, і покличу збіжжя, і помножу його, і не дам на вас голоду.
EZEK|36|30|І намножу плід дерева та врожай поля, щоб ви більше не набиралися сорому через голод між народами.
EZEK|36|31|І згадаєте ви про ваші дороги лихі та про ваші вчинки, що не добрі, і будете бридитися самих себе за свої провини та за гидоти свої.
EZEK|36|32|Не для вас Я це робитиму, говорить Господь Бог, нехай буде це вам відоме! Зашарійтеся та посоромтеся ваших доріг, Ізраїлів доме!
EZEK|36|33|Так говорить Господь Бог: Того дня, коли Я очищу вас зо всіх ваших провин, то позаселюю ці міста, і будуть забудовані руїни.
EZEK|36|34|А спустошена земля буде оброблювана за те, що була спустошенням на очах кожного перехожого.
EZEK|36|35|І скажуть: Цей опустошілий Край став як той еденський садок, а ці міста, повалені й попустошені та поруйновані, тепер укріплені та замешкані!
EZEK|36|36|І пізнають народи, які зостануться навколо вас, що Я, Господь, забудував поруйноване, засадив спустошіле. Я, Господь, говорив це і зробив!
EZEK|36|37|Так говорить Господь Бог: Ще на це прихилюся до Ізраїлевого дому, щоб зробити їм: помножу їх, як людську отару!
EZEK|36|38|Як освячена отара, як отара Єрусалиму в його свята, такі будуть ці поруйновані міста, повні отари людської, і пізнають вони, що Я Господь!
EZEK|37|1|Була надо мною Господня рука, і Дух Господній випровадив мене, і спинив мене серед долини, а вона повна кісток!
EZEK|37|2|І Він обвів мене біля них навколо, аж ось їх дуже багато на поверхні долини, і ось вони стали дуже сухі!
EZEK|37|3|І сказав Він мені: Сину людський, чи оживуть оці кості? А я відказав: Господи Боже, Ти знаєш!
EZEK|37|4|І сказав Він мені: Пророкуй про ці кості, та й скажеш до них: Сухі кості, послухайте слова Господнього!
EZEK|37|5|Так говорить Господь Бог до цих кісток: Ось Я введу у вас духа і ви оживете!
EZEK|37|6|І дам на вас жили, і виросте на вас тіло, і простягну на вас шкіру, і дам у вас духа, і ви оживете. І пізнаєте ви, що Я Господь!
EZEK|37|7|І пророкував я, як наказано. І знявся шум, коли я пророкував, і ось гуркіт, а кості зближалися, кістка до кістки своєї.
EZEK|37|8|І побачив я, аж ось на них жили, і виросло тіло, і була натягнена на них шкіра зверху, та духа не було в них.
EZEK|37|9|І сказав Він мені: Пророкуй до духа, пророкуй, сину людський, та й скажеш до духа: Так говорить Господь Бог: Прилинь, духу, з чотирьох вітрів, і дихни на цих забитих, і нехай оживуть!
EZEK|37|10|І я пророкував, як Він наказав був мені, і ввійшов у них дух, і вони ожили, і поставали на ноги свої, військо дуже-дуже велике!...
EZEK|37|11|І сказав Він мені: Сину людський, ці кості вони ввесь Ізраїлів дім. Ось вони кажуть: Повисихали наші кості, і загинула наша надія, нам кінець!
EZEK|37|12|Тому пророкуй та й скажеш до них: Так говорить Господь Бог: Ось Я повідчиняю ваші гроби, і позводжу вас із ваших гробів, мій народе, і введу вас до Ізраїлевої землі!
EZEK|37|13|І пізнаєте ви, що Я Господь, коли Я повідчиняю ваші гроби, і коли позводжу вас із ваших гробів, Мій народе!
EZEK|37|14|І дам Я в вас Свого Духа, і ви оживете, і вміщу вас на вашій землі, і пізнаєте ви, що Я, Господь, сказав це й зробив, говорить Господь!
EZEK|37|15|І було мені слово Господнє таке:
EZEK|37|16|А ти, сину людський, візьми собі один кусок дерева, і напиши на ньому: Юді та синам Ізраїля, його друзям. І візьми ще один кусок дерева, і напиши на ньому: Йосипові дерево Єфрема та всьому домові Ізраїля, друзям його.
EZEK|37|17|І зблизь їх собі одне до одного на один кусок дерева, і вони стануть за одне в твоїй руці!
EZEK|37|18|І як скажуть до тебе сини твого народу, говорячи: Чи не оголосиш нам, що це в тебе таке?
EZEK|37|19|то скажи їм: Так говорить Господь Бог: Ось Я візьму дерево Йосипа, що в Єфремовій руці, та племена Ізраїлеві, його друзів, і дам на нього дерево Юди, і вчиню їх за одне дерево, і стануть вони одним у Моїй руці!
EZEK|37|20|І будуть ці дерева, що напишеш на них, у руці твоїй на їхніх очах.
EZEK|37|21|І скажи до них: Так говорить Господь Бог: Ось Я візьму Ізраїлевих синів з-посеред народів, куди вони пішли, і позбираю їх знавкола, і введу їх до їхньої землі.
EZEK|37|22|І зроблю їх за один народ у Краї на Ізраїлевих горах, і буде для всіх них один цар за царя, і не будуть уже двома народами, і не будуть уже більш поділені на двоє царств.
EZEK|37|23|І більш не будуть вони занечищуватися своїми бовванами й гидотами своїми та всіма своїми переступами, спасу їх зо всіх їхніх осель, де вони грішили, й очищу їх. І будуть вони мені народом, а Я буду їм Богом!
EZEK|37|24|А раб Мій Давид буде царем над ними, і один пастир буде для всіх них, і постановами Моїми вони будуть ходити, а устави Мої будуть стерегти й виконувати їх.
EZEK|37|25|І осядуть вони на тій землі, яку Я дав був Моєму рабові Яковові, що сиділи на ній їхні батьки, і осядуть на ній вони та їхні сини, та сини синів їхніх аж навіки, а Мій раб Давид буде їм князем навіки!
EZEK|37|26|І складу з ними заповіта миру, це буде вічний заповіт із ними. І зміцню їх, і намножу їх, і дам Свою святиню серед них на віки!
EZEK|37|27|І буде місце Мого пробування над ними, і Я буду їм Богом, а вони Мені будуть народом.
EZEK|37|28|І пізнають ці народи, що Я Господь, що освятив Ізраїля, коли буде Моя святиня серед них навіки!
EZEK|38|1|І було мені слово Господнє таке:
EZEK|38|2|Сину людський, зверни своє обличчя до Ґоґа, краю Маґоґа, князя Рошу, Мешеху та Тувалу, і пророкуй на нього
EZEK|38|3|та й скажеш: Так сказав Господь: Ось Я проти тебе, Ґоґу, княже Рошу, Мешеху та Тувалу!
EZEK|38|4|І заверну тебе, і вкладу гачки в щелепи твої, і виведу тебе та все військо твоє, коней та верхівців, усі вони досконало озброєні, велике зборище, зо щитами та щитками, усі озброєні мечами.
EZEK|38|5|Парас, Куш і Пут із ними, усі вони зо щитом та з шоломом.
EZEK|38|6|Ґомер і всі орди його, дім Тоґарми, кінці північні та всі відділи його, численні народи з тобою.
EZEK|38|7|Приготуйся, і приготуй собі ти та все зборище твоє, зібрані при тобі, і будеш для них сторожею.
EZEK|38|8|По багатьох днях ти будеш потрібний, у кінці років прийдеш до Краю, що повернений від меча, що зібраний від численних народів, на Ізраїлеві гори, що завжди були руїною, а він був виведений від народів, і всі вони сидять безпечно.
EZEK|38|9|І вийдеш, прийдеш як буря, будеш як хмара, щоб покрити землю, ти та всі відділи твої, та численні народи з тобою.
EZEK|38|10|Так говорить Господь Бог: І станеться того дня, увійдуть слова на твоє серце, і ти будеш думати злу думку,
EZEK|38|11|та й скажеш: Піду на неукріплений край, знайду спокійних, що безпечно сидять, усі вони сидять в осадах без муру, і нема в них засува та воріт,
EZEK|38|12|щоб набрати здобичі, і чинити грабунок, щоб повернути свою руку на заселені руїни, і на народ, зібраний з народів, що набувають добуток та маєток, що сидять посеред землі.
EZEK|38|13|Шева та Дедан, і купці Таршішу, і всі левчуки його скажуть тобі: Чи ти прийшов набрати здобичі, чи ти зібрав своє зборище, щоб чинити грабунок, щоб винести срібло та золото, щоб набрати добутку та маєтку, щоб набрати великої здобичі?
EZEK|38|14|Тому пророкуй, сину людський, та й скажеш до Ґоґа: Так говорить Господь Бог: Чи того дня, коли народ Мій сидітиме безпечно, ти не довідаєшся про це?
EZEK|38|15|І прийдеш із свого місця, із північних кінців, ти та численні народи з тобою, всі вони гарцюють на конях, зборище велике й військо численне!
EZEK|38|16|І здіймешся на народ Мій Ізраїлів, як хмара, щоб покрити землю. Буде це на кінці днів, і виведу тебе на Мій Край, щоб народи пізнали Мене, коли Я покажу Свою святість тобі, Ґоґу, на їхніх очах.
EZEK|38|17|Так говорить Господь Бог: Чи ти той, що про нього говорив Я за давніх днів через Моїх рабів, Ізраїлевих пророків, що пророкували за тих днів про роки, щоб привести тебе на них?
EZEK|38|18|І станеться того дня, у дні приходу Ґоґа на Ізраїлеву землю, говорить Господь Бог, увійде ревність Моя в ніздрі Мої.
EZEK|38|19|І в ревності своїй, в огні Свого гніву Я сказав: цього дня буде великий трус на Ізраїлевій землі.
EZEK|38|20|І затремтять перед Моїм лицем морські риби та птаство небесне, і польова звірина, всяке гаддя, що плазує по землі, і всяка людина, що на поверхні землі, і будуть поруйновані гори, і поваляться урвища, і всякий мур на землю впаде.
EZEK|38|21|І покличу проти нього меча на всіх горах Моїх, говорить Господь Бог, меч кожного буде на брата його!
EZEK|38|22|І буду судитися з ними моровицею та кров'ю, і пущу заливний дощ та камінний град, огонь та сірку на нього та на відділи його, та на численні народи, що з ним.
EZEK|38|23|І звеличуся, і покажу Свою святість, і буду пізнаний на очах численних народів, і вони пізнають, що Я Господь!
EZEK|39|1|А ти, сину людський, пророкуй на Ґоґа та й скажеш: Так говорить Господь Бог: Ото Я на тебе, княже Рошу, Мешеху та Тувалу!
EZEK|39|2|І верну тебе, і попроваджу тебе, і підійму тебе з північних кінців, і впроваджу тебе на Ізраїлеві гори.
EZEK|39|3|І виб'ю лука твого з твоєї лівиці, а твої стріли кину з твоєї правиці.
EZEK|39|4|Упадеш на Ізраїлевих горах ти й усі відділи твої та народи, що з тобою; віддам тебе на з'їдження хижому птаству, усякому крилатому та польовій звірині.
EZEK|39|5|На відкритому полі впадеш ти, бо це Я говорив, говорить Господь Бог!
EZEK|39|6|І пошлю Я огонь на Маґоґа та на тих, що безпечно замешкують острови, і пізнають вони, що Я Господь!
EZEK|39|7|А Своє святе Ім'я розголошу посеред Мого народу Ізраїля, і більше не дам зневажити святе Моє Ймення, і народи пізнають, що Я Господь, Святий Ізраїлів!
EZEK|39|8|Ось прийде і станеться, говорить Господь Бог, це той день, що Я говорив.
EZEK|39|9|І повиходять мешканці Ізраїлевих міст, і накладуть огонь, і палитимуть зброю та щитка й щита, лука та стріли, і ручноно кия та ратище, і будуть ними палити огонь сім років.
EZEK|39|10|І не будуть носити дров з поля, і не будуть рубати з лісів, бо зброєю будуть палити огонь, і візьмуть здобич із тих, хто брав здобич із них, і пограбують тих, хто їх грабував, говорить Господь Бог.
EZEK|39|11|І станеться того дня, дам Я там Ґоґові місце гробу в Ізраїлі, Долину Перехожих, на схід від моря, і що замикає дорогу перехожим. І поховають там Ґоґа й усе його многолюдство, та й назвуть: Долина Многолюдства Ґоґа.
EZEK|39|12|І буде ховати їх Ізраїлів дім, щоб очистити землю, сім місяців.
EZEK|39|13|І буде ховати ввесь народ краю, і він стане для них за пам'ятку, того дня, коли Я прославлю Себе, говорить Господь Бог.
EZEK|39|14|І відділять людей, які без перерви ходитимуть по краю й ховатимуть з перехожими позосталих ще на поверхні землі, щоб її очистити. По семи місяцях вони ще будуть вишукувати.
EZEK|39|15|І перейдуть ті обхідники по краю, і коли хто побачить людську кістку, то поставить при ній знака, аж поки не поховають її похоронники в Долині Многолюдства Ґоґа.
EZEK|39|16|А ім'я міста Гамона. І очистять землю.
EZEK|39|17|А ти, сину людський, так говорить Господь Бог: Скажи птахові, усякому крилатому, та всій польовій звірині: Згромадьтеся й прийдіть, зберіться навколо над жертвою, що Я принесу для вас, велика жертва на Ізраїлевих горах, і ви будете їсти м'ясо, і будете пити кров.
EZEK|39|18|Ви будете їсти тіло лицарів, а кров князів землі будете пити, барани, і вівці, і козли, бики, ситі башанські бики всі вони.
EZEK|39|19|І будете їсти лій аж до ситости, і будете пити кров аж до впоєння з Моєї жертви, яку Я приніс для вас,
EZEK|39|20|і насититеся при Моєму столі кіньми та верхівцями, лицарями та всякими вояками, говорить Господь Бог!
EZEK|39|21|І дам Свою славу між народами, і побачать усі народи Мій суд, що зроблю Я, та Мою руку, що на них покладу.
EZEK|39|22|І пізнає Ізраїлів дім, що Я Господь, їхній Бог, від цього дня й далі.
EZEK|39|23|І пізнають народи, що Ізраїлів дім пішов на вигнання за провини свої, за те, що спроневірилися Мені, а Я сховав був від них лице Своє, і віддав їх у руку їхніх неприятелів, і всі вони попадали від меча.
EZEK|39|24|За їхньою нечистістю та за їхнє беззаконня зробив Я це з ними, і сховав від них лице Своє.
EZEK|39|25|Тому так говорить Господь Бог: Тепер поверну долю Якова, і змилуюся над усім Ізраїлевим домом, і буду ревний за Своє святе Ймення.
EZEK|39|26|І відчують вони свою ганьбу та все своє спроневірення, яким спроневірилися Мені, коли сядуть безпечно на своїй землі, і не буде вже нікого, хто б їх страшив,
EZEK|39|27|коли поверну їх з народів, і позбираю їх із країв їхніх ворогів, і покажу Свою святість у них на очах численних народів.
EZEK|39|28|І пізнають вони, що Я Господь, Бог їхній, коли вижену їх у полон до народів, а потому позбираю їх на їхню землю, і більш не позоставлю там нікого з них.
EZEK|39|29|І не сховаю вже від них Свого лиця, бо виллю Духа Свого на Ізраїлів дім, говорить Господь Бог!
EZEK|40|1|Двадцятого й п'ятого року нашого вигнання, на початку року, десятого дня місяця, чотирнадцятого року по тому, як було зруйноване місто, того самого дня була на мені Господня рука, і Він упровадив мене туди.
EZEK|40|2|У Божих видіннях упровадив Він мене до Ізраїлевого Краю, і дав спочити мені на дуже високій горі, а на ній була ніби будова міста, з полудня.
EZEK|40|3|І привів мене туди, і ось чоловік, що його вид, ніби вид блискучої міді, а в його руці льняна нитка та мірнича палиця, і він стояв у брамі.
EZEK|40|4|І сказав мені цей чоловік: Сину людський, дивися своїми очима й слухай своїми вухами, і зверни своє серце на все, що я покажу тобі, бо ти приведений сюди, щоб показати тобі. Усе, що ти побачиш, об'яви Ізраїлевому домові.
EZEK|40|5|І ось мур назовні храму навколо, а в руці того чоловіка мірнича палиця на шість ліктів, на міру ліктем та долонею. І зміряв він ширину тієї будівлі одна палиця, і заввишки одна палиця.
EZEK|40|6|І прийшов він до брами, що її перед у напрямі до сходу, і ввійшов її сходами, і зміряв порога тієї брами одна палиця завширшки, і другий поріг одна палиця завширшки.
EZEK|40|7|А вартівня одна палиця завдовжки й одна палиця завширшки, а поміж вартівнями п'ять ліктів; а поріг брами з боку сінечок тієї брами, зсередини одна палиця.
EZEK|40|8|І зміряв він сіни тієї брами зсередини одна палиця.
EZEK|40|9|І зміряв сіни брами вісім ліктів, а стовпи її два лікті, а сіни брами зсередини.
EZEK|40|10|А брамні вартівні в напрямі на схід три звідси й три звідти, і міра одна їм трьом, і міра одна стовпам звідси та звідти.
EZEK|40|11|І зміряв він ширину входу до брами десять ліктів, довжина брами тринадцять ліктів.
EZEK|40|12|А розмежування перед вартівнями один лікоть, і один лікоть звідти, а вартівня шість ліктів звідси й шість ліктів звідти.
EZEK|40|13|І зміряв браму з даху вартівні до даху її, завширшки двадцять і п'ять ліктів, двері навпроти дверей.
EZEK|40|14|І поробив стовпи, шістдесят ліктів, і до стовпів підходить подвір'я, навколо брами.
EZEK|40|15|А від переду брамного входу аж до переду сіней внутрішньої брами п'ятдесят ліктів.
EZEK|40|16|І були вікна, широкі знадвору й вузькі в середині, до вартівень та до їхніх стовпів у середині брами навколо, і так до сіней, і вікна навколо до середини, а на стовпах вирізьблені пальми.
EZEK|40|17|І він впровадив мене до зовнішнього подвір'я. І ось комори та підлога, викладена з каміння, зроблена для подвір'я навколо, тридцять комір на підлозі.
EZEK|40|18|А ця підлога була позад брам, по довжині брам, долішня підлога.
EZEK|40|19|І зміряв він ширину від переду долішньої брами до переду внутрішнього подвір'я назовні, сто ліктів, на схід та на північ.
EZEK|40|20|А та брама, що перед її в напрямі на північ до зовнішнього подвір'я, він зміряв довжину її та ширину її.
EZEK|40|21|І вартівні її три звідси й три звідти, і стовпи її, і сіни її були за мірою першої брами, п'ятдесят ліктів довжина її, а ширина двадцять і п'ять на міру ліктем.
EZEK|40|22|А вікна її, і сіни її та вирізьблені пальми її за мірою брами, що перед її в напрямі на схід, а сімома східцями входять у неї, а її сіни перед ними.
EZEK|40|23|І брама внутрішнього подвір'я навпроти брами на північ та на схід. І зміряв він від брами до брами сто ліктів.
EZEK|40|24|І він попровадив мене в напрямі на південь, аж ось брама в напрямі на південь. І він зміряв стовпи її та сіни її за тими мірами.
EZEK|40|25|А в неї вікна та сіни її навколо, які ті вікна, п'ятдесят ліктів завдовжки, а завширшки двадцять і п'ять ліктів.
EZEK|40|26|А семеро східців вхід до неї, і сіни її перед ними, а вирізьблені пальми її одна звідси, а одна звідти при стовпах її.
EZEK|40|27|А брама внутрішнього подвір'я у напрямі на південь, і він зміряв від брами до брами в напрямі на південь сто ліктів.
EZEK|40|28|І впровадив мене до внутрішнього подвір'я південною брамою, і зміряв південну браму за тими мірами.
EZEK|40|29|І вартівні її, і стовпи її, і сіни її за тими мірами, і вікна її, і в сінях її навколо п'ятдесят ліктів завдовжки, а завширшки двадцять і п'ять ліктів.
EZEK|40|30|А сіни її навколо завдовжки двадцять і п'ять ліктів, а завширшки п'ять ліктів.
EZEK|40|31|І сіни її при зовнішньому подвір'ї, і пальми при стовпах її, а вісім сходів її вхід.
EZEK|40|32|І він упровадив мене до внутрішнього подвір'я в напрямі на схід, і зміряв брами за тими мірами.
EZEK|40|33|І вартівні її, і стовпи її, і сіни її за тими мірами, а в неї вікна та в її сінях навколо, завдовжки п'ятдесят ліктів, а завширшки двадцять і п'ять ліктів.
EZEK|40|34|А її сіни були до зовнішнього подвір'я, а пальми її при її стовпах звідси й звідти, а вісім східців її вхід.
EZEK|40|35|І впровадив мене до північної брами, і зміряв тими мірами.
EZEK|40|36|Вартівні її, стовпи її, і її сіни та вікна в неї навколо, завдовжки п'ятдесят ліктів, а завширшки двадцять і п'ять ліктів.
EZEK|40|37|А стовпи її до зовнішнього подвір'я, а пальми при стовпах її з цього й з того боку, а вісім сходів її вхід.
EZEK|40|38|І комора, і її вхід у стовпах брам, там полощуть цілопалення.
EZEK|40|39|А в сінях брами два столи звідси й два столи звідти, щоб різати на них цілопалення й жертви за гріх та жертви за провину.
EZEK|40|40|А при зовнішньому боці, що підіймається до входу північної брами, два столи, і при боці іншому, що при сінях брами, два столи.
EZEK|40|41|Чотири столи звідси й чотири столи звідти при боці брами, вісім столів, що на них ріжуть.
EZEK|40|42|І чотири столи на цілопалення, каміння тесане, завдовжки лікоть один і і пів, а заввишки один лікоть; на них кладуть знаряддя, що ними ріжуть цілопалення та жертву.
EZEK|40|43|І гаки, на одну долоню, були приготовлені в домі навколо, а на столах жертовне м'ясо.
EZEK|40|44|А назовні внутрішньої брами були дві кімнаті у внутрішньому подвір'ї, що при північному боці брами, а їхній перед у напрямі на південь, одна при боці східньої брами, перед її у напрямі на північ.
EZEK|40|45|І сказав він до мене: Ця кімната, що перед її в напрямі на південь, для священиків, що стережуть сторожу храму.
EZEK|40|46|А та кімната, що перед її в напрямі на північ, для священиків, що виконують сторожу жертівника. Це Садокові сини, що з Левієвих синів наближуються до Господа, щоб служити Йому.
EZEK|40|47|І зміряв подвір'я завдовжки сто ліктів, і завширшки сто ліктів, чотирикутнє, а жертівник був перед храмом.
EZEK|40|48|І впровадив мене до сіней храму, і зміряв стовпа сіней, п'ять ліктів звідси, і п'ять ліктів звідти, а ширина брами три лікті звідси й три лікті звідти.
EZEK|40|49|Довжина сіней двадцять ліктів, а завширшки одинадцять ліктів, а десятьма сходами ходять до нього; а стовпи при стовпах, один звідси, а один звідти.
EZEK|41|1|І впровадив мене до храму, і він зміряв стовпи, шість ліктів завширшки звідси, і шість ліктів завширшки звідти, ширина скинії.
EZEK|41|2|А ширина входу десять ліктів, а боки входу п'ять ліктів звідси й п'ять ліктів звідти; і зміряв довжину його сорок ліктів, а завширшки двадцять ліктів.
EZEK|41|3|І ввійшов він до середини, і зміряв входового стовпа два лікті, а вхід шість ліктів, а ширина входу сім ліктів.
EZEK|41|4|І зміряв довжину його двадцять ліктів, а завширшки двадцять ліктів на переді храму. І сказав він мені: Це Святеє Святих!
EZEK|41|5|І зміряв він стіну храму шість ліктів, а ширина бічної кімнати чотири лікті кругом навколо храму.
EZEK|41|6|А кімнати бічні, кімната при кімнаті, тридцять в трьох поверхах, і входили в стіну, що храм мав для бічних кімнат навколо кругом, щоб держалися, і не держалися в стіні того храму.
EZEK|41|7|І він ставав ширший, і обертався все більше вгору до бічних кімнат, бо той храм був обернений більше вгору, кругом навколо храму, тому храм був ширший вгору, і так долішній поверх входить на горішній через середній.
EZEK|41|8|І бачив я вишину храму навколо, підвалини бічних кімнат повна палиця, шість ліктів.
EZEK|41|9|Ширина стіни, що в бічній кімнаті назовні, п'ять ліктів, а вільне місце між бічними кімнатами, що належить до храму.
EZEK|41|10|І поміж коморами завширшки двадцять ліктів кругом навколо храму.
EZEK|41|11|А вхід з бічної кімнати до вільного місця вхід один у напрямі на північ, і вхід один на південь, а ширина вільного місця п'ять ліктів кругом навколо.
EZEK|41|12|А будівля, що перед відгородженим майданом у напрямі на захід, завширшки сімдесят ліктів, а стіна будівлі п'ять ліктів, ширина кругом навколо, а довжина її дев'ятдесят ліктів.
EZEK|41|13|І він зміряв той храм, завдовжки сто ліктів, а відгороджений майдан і будівля та стіни її, завдовжки сто ліктів.
EZEK|41|14|А ширина передньої частини храму та відгородженого майдану на схід сто ліктів.
EZEK|41|15|І зміряв він довжину будівлі до переду відгородженого майдану, що позад неї, ґалерія звідси й звідти, сто ліктів, і так внутрішній храм і сінечки подвір'я.
EZEK|41|16|Пороги та вікна, широкі знадвору, і вузькі всередині, ґалерія навколо них трьох, навпроти порогу дерев'яний обклад навколо й земля до вікон, а вікна зачинені.
EZEK|41|17|Усе понад входом і аж до внутрішнього храму, і назовні при кожній стіні кругом навколо, у внутрішньому й у зовнішньому, вирізьблене,
EZEK|41|18|і було зроблене херувимами та пальмами, і пальма була між херувимом та херувимом, два обличчя в херувима.
EZEK|41|19|І людське обличчя мали пальми звідси, а обличчя левчука мали пальми звідти, пороблені при всьому домі навколо.
EZEK|41|20|Від землі аж понад вхід пороблені херувими та пальми на стіні храму.
EZEK|41|21|Храм мав чотирикутні одвірки, а перед святині мав такий самий вигляд.
EZEK|41|22|Жертівник був із дерева, три лікті високий, а довжина його два лікті, а в нього його кути й підніжжя його та стіни його дерево. І сказав він мені: Це той стіл, що перед Господнім лицем!
EZEK|41|23|А в храмі та в святині було двоє дверей.
EZEK|41|24|І в тих дверях було по дві дошці, обидві дошки оберталися, дві в одних дверях, і дві в інших дверях.
EZEK|41|25|І були зроблені на них, на дверях храму, херувими та пальми, як пороблені були в стінах, а дерев'яний ґанок при переді сіней назовні.
EZEK|41|26|І вікна, широкі знадвору й вузькі всередині, і пальми звідси та звідти при боках сіней, і такі бічні кімнати храму та стріхи.
EZEK|42|1|І він вивів мене до зовнішнього подвір'я дорогою в напрямі на північ, і ввів мене до кімнат, що навпроти відгородженої площі, і що навпроти будівлі на північ.
EZEK|42|2|Навпроти завдовжки сто ліктів, вхід північний, а завширшки п'ятдесят ліктів.
EZEK|42|3|Навпроти двадцять ліктів, що у внутрішньому подвір'ї, і навпроти викладеної підлоги, що в зовнішньому подвір'ї, ґалерія до переду ґалерії на три поверхи.
EZEK|42|4|А перед кімнатами був хід на десять ліктів ширини до внутрішнього подвір'я, дорогою ста ліктів, а виходи їхні на північ.
EZEK|42|5|А горішні кімнати були коротші, бо ґалерії забирали від них більше місця, ніж з долішніх та з середніх тієї будівлі.
EZEK|42|6|Бо вони були триповерхові, і не було в них стовпів, як стовпи подвір'я, тому вони були вужчі від долішніх та від середніх на землі.
EZEK|42|7|А мур, що назовні навпроти кімнат, у напрямі зовнішнього подвір'я, до переду кімнат довжина його п'ятдесят ліктів.
EZEK|42|8|Бо довжина тих кімнат, що в зовнішнього подвір'я, п'ятдесят ліктів, і ось на переді храму сто ліктів.
EZEK|42|9|А під тими кімнатами хід від сходу, коли входити до них з зовнішнього подвір'я.
EZEK|42|10|По ширині муру подвір'я в напрямі на схід до переду вільного місця й до переду будівлі кімнати.
EZEK|42|11|А дорога перед ними як вид кімнат, що в напрямі на північ; яка довжина, така ширина їхня, а всі виходи були за їхніми способами та за їхніми виходами.
EZEK|42|12|І як входи кімнат, що в напрямі півдня, такий був вхід на початку дороги, дороги перед відповідним муром у напрямі на схід, коли йти до них.
EZEK|42|13|І сказав він мені: Кімнати північні і кімнати південні, що на переді вільного місця, це кімнати священні, де їдять священики, що наближуються до Господа, найсвятіше, там складають найсвятіше, і жертву хлібну, і жертву за гріх, і жертву за провину, бо це місце святе.
EZEK|42|14|Коли священики ввійдуть, то не сміють виходити зо святині до зовнішнього подвір'я, і мають там складати свої шати, в яких служать, бо вони святощі. І зодягнуть вони інші шати, і тоді тільки можуть зближатися до того, що належить народові.
EZEK|42|15|І скінчив він вимірювання внутрішнього храму, і випровадив мене в напрямі брами, що перед її в напрямі на схід, і зміряв те кругом навколо.
EZEK|42|16|Він зміряв мірничою палицею східній бік, п'ять сотень палиць мірничою палицею навколо.
EZEK|42|17|Зміряв північний бік, п'ять сотень палиць мірничною палицею навколо.
EZEK|42|18|Зміряв південний бік, п'ять сотень палиць мірничою палицею.
EZEK|42|19|Обернувся до західнього боку, наміряв п'ять сотень палиць мірничою палицею.
EZEK|42|20|На чотири сторони відміряв те. Мало воно мур кругом навколо, завдовжки п'ять сотень, і завширшки п'ять сотень, щоб відділити між святим та звичайним.
EZEK|43|1|І попровадив мене до брами, до брами, що звернена в напрямі сходу.
EZEK|43|2|І ось слава Ізраїлевого Бога йшла в напрямі від сходу, а голос Його був, як шум великої води, а земля засвітилася від слави Його!
EZEK|43|3|І вид був такий же, як я бачив: як те видиво, що я бачив, коли я приходив руйнувати місто, і види були, як той вид, що я бачив при річці Кевар. І впав я на обличчя своє!
EZEK|43|4|І слава Господня ввійшла в храм у напрямі брами, що перед її в напрямі сходу!
EZEK|43|5|І підняв мене Дух, і впровадив мене до внутрішнього подвір'я, і ось слава Господня наповнила храм!
EZEK|43|6|І почув я Промовляючого до мене з храму, а той муж стояв при мені.
EZEK|43|7|І сказав Він мені: Сину людський, це місце престолу Мого, і місце стіп Моїх ніг, де Я буду перебувати навіки посеред Ізраїлевих синів, не занечистить уже Ізраїлів дім святе Ім'я Моє, вони та їхні царі розпустою своєю та трупами їхніх царів при їхньому вмиранні!
EZEK|43|8|Вони ставили свого порога при Моєму порозі, і свої одвірки при одвірках Моїх, так що тільки стіна була між Мною та між ними, і вони занечистили святе Ім'я Моє своїми гидотами, яких наробили, і Я вигубив їх у Своїм гніві...
EZEK|43|9|Тепер нехай вони віддалять від Мене розпусту свою та трупи своїх царів, і Я буду пробувати між ними навіки.
EZEK|43|10|Ти, сину людський, об'яви Ізраїлевому домові про цей храм, і вони посоромляться від своїх провин, і зміряють міру.
EZEK|43|11|А якщо вони засоромляться від усього, чого наробили, то виясни їм вигляд храму, і план його, і виходи його та його входи, і всі устави його, і всі начерки його, і всі закони його, і напиши це на очах їх, і нехай вони стережуть усякий начерк його, і всі устави його, і нехай вони роблять їх!
EZEK|43|12|Оце закон храму: на вершині гори вся границя його кругом навколо має бути Святеє Святих. Ось це закон храму.
EZEK|43|13|А оце міри жертівника ліктями, лікоть це лікоть та долоня. І основа жертівника лікоть, і лікоть завширшки, а його границя до його краю навколо одна п'ядь, і це задня сторона жертівника.
EZEK|43|14|А від основи на землі аж до долішнього обкладу жертівника два лікті, а завширшки один лікоть, а від малого відступу жертівника аж до великого чотири лікті, а завширшки лікоть.
EZEK|43|15|А жертівник чотири лікті високий, а від жертівника й вище чотири роги.
EZEK|43|16|А огнище дванадцять ліктів завдовжки на дванадцять завширшки, чотирикутнє при чотирьох своїх боках.
EZEK|43|17|А долішній обклад чотирнадцять ліктів завдовжки на чотирнадцять завширшки при чотирьох боках її, а границя навколо нього півліктя, а основа його лікоть навколо, а сходи його звернені на схід.
EZEK|43|18|І сказав Він мені: Сину людський, так говорить Господь Бог: Оце устави жертівника на день, коли він буде зроблений, щоб приносити на ньому цілопалення, і кропити на нього кров.
EZEK|43|19|І даси священикам-Левитам, що вони з Садокового насіння, що наближуються до Мене, говорить Господь Бог, щоб служили Мені, молодого бика з великої худоби на жертву за гріх.
EZEK|43|20|І візьмеш з його крови, і покропи на чотири його роги й до чотирьох кутів оправи та до границі навколо, і очисти його та освяти його.
EZEK|43|21|І візьмеш бика тієї жертви за гріх, і спалять його на означеному місці храму назовні святині.
EZEK|43|22|А другого дня принесеш у жертву козла безвадного на жертву за гріх, і очистять жертівника, як очистили биком.
EZEK|43|23|А коли покінчиш очищати, принесеш у жертву молодого бика з великої худоби, безвадного, і безвадного барана з отари.
EZEK|43|24|І приведи їх перед Господнє лице, і кинуть священики на них сіль, і принесуть їх цілопаленням для Господа.
EZEK|43|25|Сім день будеш приготовляти козла жертви за гріх на кожен день, і молодого бика з великої худоби, і барана з отари, безвадних приготовлять.
EZEK|43|26|Сім день будуть очищати того жертівника, і очистять його, і освятять його.
EZEK|43|27|І скінчаться ті дні, і станеться, восьмого дня й далі приготовлять священики на жертівнику ваші цілопалення та ваші жертви мирні, і вподобаю Собі вас, говорить Господь Бог!
EZEK|44|1|І вернув мене в напрямі брами зовнішньої святині, що обернена на схід, а вона замкнена.
EZEK|44|2|І сказав мені Господь: Брама ця буде замкнена, не буде відчинена, і ніхто не ввійде в неї, бо в неї ввійшов Господь, Бог Ізраїлів, і вона буде замкнена.
EZEK|44|3|Князь, сам князь буде сидіти в ній, щоб їсти хліб перед Господнім лицем; сіньми брами він увійде, і сіньми вийде.
EZEK|44|4|І випровадив мене в напрямі північної брами до переду храму, і побачив я, аж ось слава Господня наповнила Господній дім! І впав я на обличчя своє...
EZEK|44|5|І сказав мені Господь: Сину людський, зверни своє серце, і побач своїми очима, а своїми вухами послухай усе, що Я говоритиму з тобою щодо всіх постанов Господнього дому, і щодо всяких законів його, і звернеш своє серце до входу того храму в усіх виходах святині.
EZEK|44|6|І скажеш до ворохобників, до Ізраїлевого дому: Так говорить Господь Бог: Досить вам усіх ваших гидот, Ізраїлів доме,
EZEK|44|7|що ви вводили чужинців, необрізаносердих та необрізанотілих, щоб були в Моїй святині, щоб зневажити його, Мій храм, коли приносили Мій хліб, лій та кров, і, крім усіх ваших гидот, зламали Мого заповіта.
EZEK|44|8|І ви не несли сторожі святощів Моїх, але поставили їх собі за сторожів Моєї варти в Моїй святині.
EZEK|44|9|Так говорить Господь Бог: Кожен чужинець, необрізаносердий та необрізанотілий не ввійде до Моєї святині; це і про всякого чужинця, що живе серед Ізраїлевих синів.
EZEK|44|10|І навіть Левити, що були віддалилися від Мене, коли блукав Ізраїль, що були зблудили від Мене за своїми божками, і вони понесуть кару за свою вину,
EZEK|44|11|і будуть вони в святині Моїй служити сторожами при брамах храму, і обслуговувати храм, вони будуть приносити цілопалення й жертву народові, і вони будуть ставати перед ними, щоб служити їм.
EZEK|44|12|За те, що вони служили їм перед їхніми бовванами, і стали для Ізраїлевого дому за спотикання на провину, тому підняв Я Свою руку на них, говорить Господь Бог, і вони понесуть провину свою!
EZEK|44|13|І вони не підійдуть до Мене, щоб бути священиками Мені, і щоб підходити до всіх святощів Моїх, до Святого Святих, і будуть носити ганьбу свою та гидоти свої, які наробили...
EZEK|44|14|І дам Я їх сторожами варти храму щодо всієї його праці, і щодо всього, що робиться в ньому.
EZEK|44|15|А священики-Левити, Садокові сини, що несли сторожу Моєї святині, коли Ізраїлеві сини зблудили були від Мене, вони наблизяться до Мене на службу Мені, і будуть стояти перед Моїм лицем, щоб приносити Мені лій та кров, говорить Господь Бог.
EZEK|44|16|Вони ввійдуть до Моєї святині, і вони наблизяться до Мого столу на службу Мені, і будуть нести Мої сторожі.
EZEK|44|17|І станеться, коли вони входитимуть до брами внутрішнього подвір'я, то зодягатимуть льняну одіж, і не ввійде на них вовна, коли вони служитимуть у брамах внутрішнього подвір'я та назовні.
EZEK|44|18|Льняні завої будуть на їхній голові, а льняна спідня одежа буде на їхніх стегнах; не будуть оперізуватися тим, що викликає піт.
EZEK|44|19|А коли вони будуть виходити до зовнішнього подвір'я, до народу, здійматимуть шати свої, в яких служили, і поскладають їх у священних кімнатах, і зодягнуть іншу одежу, щоб своїми священними шатами не торкатися народу.
EZEK|44|20|А голови своєї вони не будуть голити, і волосся не запустять, конче будуть стригти волосся своє.
EZEK|44|21|І вина не будуть пити кожен із священиків, коли мають входити до внутрішнього подвір'я.
EZEK|44|22|А вдів та розвідок не братимуть собі за жінок, а братимуть тільки дівчат із насіння Ізраїлевого дому, та вдову, що буде вдовою по священикові.
EZEK|44|23|А народ Мій будуть вони навчати розрізняти між святим та звичайним, і зроблять їх знаючими різницю між нечистим та чистим.
EZEK|44|24|А в суперечці вони стануть, щоб судити, правосуддям Моїм розсудять її, і будуть стерегти Закони Мої, і устави Мої при всіх святах Моїх, і суботи Мої будуть святити!
EZEK|44|25|І до мертвої людини не підійдуть, щоб не занечистити себе, а тільки ради батька й матері, і ради сина, і дочки, і ради брата й сестри, що не належала чоловікові, занечистяться.
EZEK|44|26|А по його очищенні прирахують йому ще сім день.
EZEK|44|27|А того дня, коли він входить до святині, до внутрішнього подвір'я, щоб служити в святині, він принесе свою жертву за гріх, говорить Господь Бог.
EZEK|44|28|І оце буде їм за спадщину: Я їхня спадщина, а володіння не дасте їм в Ізраїлі, Я їхнє володіння!
EZEK|44|29|Жертву хлібну, і жертву за гріх, і жертву за провину, оце будуть вони їсти, і все закляте в Ізраїлі буде їхнє.
EZEK|44|30|І перше з усяких первонароджених зо всього, і всякі приношення всього зо всіх ваших приношень буде священикам, і початок ваших діж дасте священикові, щоб він поклав благословення на вашому домі.
EZEK|44|31|Усякого падла та пошматованого з птаства та скотини священики не будуть їсти.
EZEK|45|1|А коли ви будете кидати жеребка про землю в спадщину, то дасте приношення Господеві, святе із землі, двадцять і п'ять тисяч ліктів завдовжки, а десять тисяч завширшки йому. Це буде святе в усій його границі навколо.
EZEK|45|2|З того буде для святині чотирикутнє місце довкола, п'ять сотень на п'ять сотень, і п'ятдесят ліктів вигін йому навколо.
EZEK|45|3|А з цієї міри відміряєш двадцять і п'ять тисяч ліктів завдовж та десять тисяч завшир, і в цьому буде святиня, Святеє Святих.
EZEK|45|4|Це святість із землі; вона буде для священиків, що служать святині, для тих, що наближуються, щоб служити Господеві, і буде їм місцем для домів і святим місцем.
EZEK|45|5|А двадцять і п'ять тисяч ліктів завдовж і десять тисяч завшир буде для Левитів, що служать храмові, їм на володіння, міста на сидіння.
EZEK|45|6|А на володіння місту дасте п'ять тисяч завшир і двадцять і п'ять тисяч завдовж, навпроти святого приношення; воно буде для всього Ізраїлевого дому.
EZEK|45|7|А для князя буде з того й з того боку святого приношення й володіння міста, навпроти святого приношення й на переді володіння міста від західнього краю на захід, і від східнього краю на схід, а завдовж відповідно одній частині племена від західньої границі до границі східньої
EZEK|45|8|землі; це буде йому за володіння в Ізраїлі, і Мої князі не будуть уже тиснути народу Мого, а Край дадуть Ізраїлевому домові, їхнім племенам.
EZEK|45|9|Так говорить Господь Бог: Досить вам, Ізраїлеві князі! Насильство та утиски відсуньте, а робіть правосуддя та правду, перестаньте випихати народ Мій з його землі, говорить Господь Бог!
EZEK|45|10|Майте справедливу вагу, і справедливу ефу та справедливого бата.
EZEK|45|11|Ефа й бат буде однакова міра, щоб бат виносив десяту частину хомеру, а десята частина хомеру ефа; згідно з хомером буде міра його.
EZEK|45|12|А шекель двадцять ґерів; двадцять шеклів, двадцять і п'ять шеклів, та п'ятнадцять шеклів буде вам міна.
EZEK|45|13|Оце те приношення, що ви принесете: шоста частина ефи з хомеру пшениці й шоста частина ефи з хомеру ячменю.
EZEK|45|14|А постанова про оливу з бата оливи: десята частина бата з кору, десять батів хомер, бо десять батів хомер.
EZEK|45|15|І одна штука з отари з двохсот штук з доброго пасовиська Ізраїлевого на жертву хлібну, і на цілопалення, і на жертви мирні, щоб очистити їх, говорить Господь Бог.
EZEK|45|16|Увесь народ цього Краю повинен давати приношення для князя в Ізраїлі.
EZEK|45|17|А на обов'язку князя буде: цілопалення, і жертва хлібна та жертва лита в свята, і в новомісяччя та в суботи, в усі свята Ізраїлевого дому, він приготує жертву за гріх, і жертву хлібну, і цілопалення, і жертви мирні на очищення за Ізраїлів дім.
EZEK|45|18|Так говорить Господь Бог: У першому місяці, першого дня місяця візьмеш молодого бика з великої худоби, безвадного, й очистиш святиню.
EZEK|45|19|І візьме священик з крови жертви за гріх, і покропить на одвірок храму та на чотири кути відступу жертівника, і на одвірок брами внутрішнього подвір'я.
EZEK|45|20|І так зробиш сьомого дня першого місяця за кожного, хто прогрішиться через помилку або з глупоти, і очистите храма.
EZEK|45|21|У першому місяці, чотирнадцятого дня місяця буде вам Пасха, свято семиденне; будете їсти опрісноки.
EZEK|45|22|І приготує того дня князь за себе та за ввесь народ Краю бика на жертву за гріх.
EZEK|45|23|І сім день свята буде він приготовлювати цілопалення для Господа, сім биків і сім баранів безвадних на день, сім день, і жертву за гріх, козла на день.
EZEK|45|24|І приготовить жертву хлібну, ефу на бика й ефу на барана, а оливи гін на ефу.
EZEK|45|25|Сьомого місяця, п'ятнадцятого дня місяця в свято буде він приготовлювати те саме, сім день, як жертву за гріх, як цілопалення, так і жертву хлібну, так і оливу.
EZEK|46|1|Так говорить Господь Бог: Брама внутрішнього подвір'я, що звернена на схід, буде замкнена шість день праці, а суботнього дня буде відчинена, і в день новомісяччя буде відчинена.
EZEK|46|2|І ввійде князь ходом сіней брами ззовні, і стане при одвірку брами, а священики приготують його цілопалення та його мирну жертву, і він поклониться на порозі брами. А брама не буде замкнена аж до вечора.
EZEK|46|3|І буде вклонятися народ Краю при вході цієї брами в суботи та в новомісяччя перед Господнім лицем.
EZEK|46|4|А те цілопалення, що князь принесе Господеві суботнього дня, це шість безвадних овець та безвадний баран.
EZEK|46|5|А жертва мучна ефа на барана, а на овець жертва хлібна, скільки дасть рука його, а оливи гін на ефу.
EZEK|46|6|А в день новомісяччя молодий бик з великої худоби, безвадний, і шестеро овець та баран будуть безвадні.
EZEK|46|7|І ефу на бика, і ефу на барана приготує він хлібну жертву, а на овець як сягне рука його, а оливи гін на ефу.
EZEK|46|8|А коли приходитиме князь, то він увійде ходом сіней брами, і тим же ходом своїм вийде.
EZEK|46|9|А коли народ Краю буде приходити перед Господнє лице в свята, то хто входить ходом північної брама, щоб поклонитися, вийде ходом брами південної, а хто входить ходом брами південної, вийде ходом брами північної, не вернеться ходом тієї брами, яким увійшов, але вийде протилеглою йому.
EZEK|46|10|А князь буде серед них: при вході їх ввійде, і при виході їх вийде.
EZEK|46|11|А в свята та в урочисті дні буде хлібна жертва, ефа на бика й ефа на барана, а на вівці скільки дасть рука його, а оливи гін на ефу.
EZEK|46|12|А коли князь приготує добровільного дара, цілопалення або мирні жертви, дар для Господа, то відчинять йому браму, що звернена на схід, і приготує своє цілопалення та свої мирні жертви, як готує за суботи, і вийде, і замкнуть браму по його виході.
EZEK|46|13|А вівцю однорічну, безвадну, приготовиш на цілопалення кожен день для Господа, щоранку приготовиш його.
EZEK|46|14|А жертву хлібну приготовиш до нього щоранку, шосту частину ефи, а оливи третину гіна, щоб покропити пшеничну муку, це хлібна жертва для Господа, постанови вічні назавжди.
EZEK|46|15|І приготують вівцю й жертву хлібну та оливу щоранку на стале цілопалення.
EZEK|46|16|Так говорить Господь Бог: Коли князь дасть кому зо своїх синів дара зо спадку свого, це буде належати його синам, як їхнє володіння в спадщині.
EZEK|46|17|А коли він дасть дара з свого спадку одному з своїх рабів, то це буде належати йому аж до року волі його, та й вернеться князеві, бо це його спадок, тільки синам його він належатиме.
EZEK|46|18|А князь не візьме зо спадку народу, витискаючи їх з їхнього володіння, із свого володіння дасть своїм синам спадок, щоб ніхто з народу Мого не розпорошився зо свого володіння.
EZEK|46|19|І впровадив мене входом, що при боці брами, до священних кімнат для священиків, що звернені на північ; і ось там є місце на їхньому задньому боці на захід.
EZEK|46|20|І сказав він мені: Оце місце, де священики будуть варити жертву за провину та жертву за гріх, де будуть пекти жертву хлібну, щоб не виносити до зовнішнього подвір'я, і не посвятити народа.
EZEK|46|21|І він вивів мене до зовнішнього подвір'я, і провів мене по чотирьох рогах подвір'я, і ось ще подвір'я на кожному розі подвір'я.
EZEK|46|22|На чотирьох рогах подвір'я були малі подвір'я, сорок ліктів завдовж і тридцять завшир, міра одна для них чотирьох, простокутні.
EZEK|46|23|І був ряд каміння навколо них, навколо них чотирьох, і пороблені кухні під горожею навколо.
EZEK|46|24|І сказав він мені: Оце дім кухарів, що там варять слуги храму жертву народові.
EZEK|47|1|І він вернув мене до дверей храму, аж ось виходить вода з-під порога храму на схід, бо перед того храму на схід. А вода сходила здолу, з правого боку храму, з півдня від жертівника.
EZEK|47|2|І він випровадив мене в напрямі брами на північ, і провів мене навколо зовнішньою дорогою до зовнішньої брами, дорогою, зверненою на схід; і ось вода виприскувала з правого боку.
EZEK|47|3|І вийшов цей чоловік на схід, а шнур був у його руці, і він відміряв тисячу ліктів, і перепровадив мене водою, водою по кістки.
EZEK|47|4|І відміряв ще тисячу, і перепровадив мене водою, водою по коліна; і відміряв ще тисячу, і перепровадив мене водою по стегна.
EZEK|47|5|І відміряв він ще тисячу, і був потік, якого я не міг перейти, бо стала великою та вода на пливання, потік, що був неперехідний.
EZEK|47|6|І сказав він мені: Чи ти бачив це, сину людський? І повів мене, і вернув мене на берег цього потоку.
EZEK|47|7|А коли я вернувся, то ось на березі потоку дуже багато дерев з цього й з того боку.
EZEK|47|8|І сказав він до мене: Ця вода виходить до східньої округи, і сходить на степ, і сходить до моря, до води солоної, і вздоровиться вода.
EZEK|47|9|І станеться, всяка жива душа, що роїться скрізь, куди приходить той потік, буде жити, і буде дуже багато риби, бо ввійшла туди та вода, і буде вздоровлена, і буде жити все, куди пройде той потік.
EZEK|47|10|І станеться, стануть при ньому рибаки від Ен-Ґеді й аж до Ен-Еґлаїму; вода буде місцем розтягнення неводу, їхня риба буде за родом своїм, як риба Великого моря, дуже численна.
EZEK|47|11|Його ж багна та калюжі його не будуть уздоровлені, на сіль вони дані.
EZEK|47|12|А над потоком виросте на його березі з цього й з того боку всяке дерево їстивне; не опаде його листя, і не перестане плід його, кожного місяця буде давати первоплоди, бо вода його вона зо святині виходить, і буде плід його на їжу, а його листя на лік.
EZEK|47|13|Так говорить Господь Бог: Оце границя, що ви посядете собі цю землю для дванадцяти Ізраїлевих племен; Йосип матиме два уділи.
EZEK|47|14|І посядете її як один, так і другий, бо, прирікаючи, підняв Я був руку Свою дати її вашим батькам, і припаде цей Край вам у спадщину.
EZEK|47|15|А оце границя Краю: на північному кінці від Великого моря напрямець до Хетлону, як іти до Цедаду,
EZEK|47|16|Хамат, Берота, Сівраїм, що між границею Дамаску та між границею Хамату, середущий Хацар, що при границі Хаврану.
EZEK|47|17|І буде границя від моря: Хацар-Енон, границя Дамаску на північ, і границя Хамату. Це північний кінець.
EZEK|47|18|А східній кінець, з-між Хаврану та з-між Дамаску, і з-між Ґілеаду та з-між Ізраїлевого краю Йордан; від границі аж до східнього моря відміряєте. Це східній кінець.
EZEK|47|19|А південний кінець, на південь: від Тамару аж до води Мерівот-Кадешу, потоку, до Великого моря. Це південний кінець, на південь.
EZEK|47|20|А західній кінець Велике море, від границі аж навпроти того, де йти на Хамат. Це західній кінець.
EZEK|47|21|І поділите цю землю собі, Ізраїлевим племенам.
EZEK|47|22|І станеться, поділите її жеребком на спадок собі та чужинцям, що мешкають серед вас, що породили синів серед вас, і стануть вам, як тубільці між синами Ізраїлевими; з вами вони кинуть жеребка про спадок серед Ізраїлевих племен.
EZEK|47|23|І станеться, у тому племені, де мешкатиме з ним той чужинець, там дасте його спадок, говорить Господь Бог.
EZEK|48|1|А оце імена племен: Від північного кінця по боці дороги до Хетлону, де йти до Хамату, Хацар-Енан, на границі Дамаску на північ, по боці Хамату, і будуть вони йому від східнього кінця аж до моря, один уділ Данові.
EZEK|48|2|А при границі Дана від східнього кінця й аж до кінця західнього, один уділ Ассирові.
EZEK|48|3|А при границі Ассира від східнього кінця аж до кінця західнього, один уділ Нефталимові.
EZEK|48|4|А при границі Нефталима від східнього кінця аж до кінця західнього, один уділ Манасії.
EZEK|48|5|А при границі Манасії від східнього кінця аж до кінця західнього, один уділ Єфремові.
EZEK|48|6|А при границі Єфрема від східнього кінця й аж до кінця західнього, один уділ Рувимові.
EZEK|48|7|А при границі Рувима від східнього кінця аж до кінця західнього, один уділ Юді.
EZEK|48|8|А при границі Юди від східнього кінця аж до кінця західнього буде те приношення, що ви принесете, ділянка на двадцять і п'ять тисяч завшир, а завдовж як одна з частин племен зо східнього кінця аж до кінця західнього, і буде в ній святиня.
EZEK|48|9|Те приношення, що принесете Господеві, ділянка буде завдовж двадцять і п'ять тисяч, а завшир двадцять тисяч.
EZEK|48|10|А святе приношення буде для оцих: ділянка священикам на північ двадцять і п'ять тисяч, а на захід завшир десять тисяч, а на схід завшир десять тисяч, а на південь завдовж двадцять і п'ять тисяч, і Господня святиня буде серед того.
EZEK|48|11|Священиками, посвяченим із синів Садока, що виконували Мою сторожу, що не блукали блуканиною Ізраїлевих синів, як блукали Левити,
EZEK|48|12|то буде їм приношення з приношення цієї землі, найсвятіша святість, при границі Левитів.
EZEK|48|13|А Левити відповідно границі священиків, ділянка їм на двадцять і п'ять тисяч завдовж, а завшир десять тисяч, уся довжина двадцять і п'ять тисяч, а ширина десять тисяч.
EZEK|48|14|І вони не продадуть із цього, і не виміняють, і первоплід землі ні до кого не перейде, бо це святість для Господа.
EZEK|48|15|А ділянка на п'ять тисяч завширшки й на двадцять і п'ять тисяч завдовжки призначається на оселення й на пасовиська, а саме те місто буде всередині.
EZEK|48|16|А оце розміри його: північний край чотири тисячі й п'ять сотень, і південний край чотири тисячі й п'ять сотень, і від східнього краю чотири тисячі й п'ять сотень, а західній край чотири тисячі й п'ять сотень.
EZEK|48|17|І буде пасовисько для міста, на північ двісті й п'ятдесят, і на південь двісті й п'ятдесят, і на схід двісті й п'ятдесят, і на захід двісті й п'ятдесят.
EZEK|48|18|А позостале на довжину навпроти святого приношення десять тисяч на схід і десять тисяч на захід, і буде воно навпроти святого приношення, і буде плід його на хліб робітникам міста.
EZEK|48|19|А робітники міста будуть оброблювати його зо всіх Ізраїлевих племен.
EZEK|48|20|Усе приношення ділянка на двадцять і п'ять тисяч завдовж і на двадцять і п'ять тисяч завшир, чотирикутнє, і піднесене святе приношення понад володіння міста.
EZEK|48|21|А позостале для князя, з цього й з того боку святого приношення та володіння міста перед тими двадцятьма й п'ятьма тисячами приношення аж до границі на схід та на захід, навпроти тих двадцяти й п'яти тисяч аж до границі на захід, навпроти частин племен, це князеві, і буде святе приношення, а святиня дому серед них.
EZEK|48|22|А з володіння Левитів і з володіння міста серед того, що буде князеві, між границею Юди й між границею Веніямина, буде це князеві.
EZEK|48|23|А решта племен від східнього кінця аж до кінця західнього, один уділ Веніяминові.
EZEK|48|24|А при границі Веніямина від східнього кінця аж до кінця західнього, один уділ Симеонові.
EZEK|48|25|А при границі Симеона від східнього кінця аж до кінця західнього, один уділ Іссахарові.
EZEK|48|26|А при границі Іссахара від східнього кінця аж до кінця західнього, один уділ Завулонові.
EZEK|48|27|А при границі Завулона від східнього кінця аж до кінця західнього, один уділ Ґадові.
EZEK|48|28|А при границі Ґада до границі південної, на півдні, то буде границя від Тамару до води Меріват-Кадешу, потоку, до Великого моря.
EZEK|48|29|Оце Край, що поділите жеребком у спадок Ізраїлевим племенам, і це їхні уділи, говорить Господь Бог.
EZEK|48|30|А оце виходи міста: з північного кінця чотири тисячі й п'ять сотень міри.
EZEK|48|31|А міські брами на імена Ізраїлевих племен, три брамі на північ: одна брама Рувимова, одна брама Юдина, одна брама Левієва.
EZEK|48|32|А при східньому кінці чотири тисячі й п'ять сотень, а брам троє: одна брама Йосипова, одна брама Веніяминова, одна брама Данова.
EZEK|48|33|І південний край чотири тисячі й п'ять сотень міри, а брам троє: одна брама Симеонова, одна брама Іссахарова, одна брама Завулонова.
EZEK|48|34|Західній кінець чотири тисячі й п'ятьсот, три їхні брамі: одна брама Ґадова, одна брама Ассирова, одна брама Нефталимова.
EZEK|48|35|Навколо вісімнадцять тисяч. А ім'я міста з того дня: Тут Господь.
