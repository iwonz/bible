ZEPH|1|1|當 亞們 的兒子 猶大 王 約西亞 在位的時候，耶和華的話臨到 希西家 的玄孫， 亞瑪利雅 的曾孫， 基大利 的孫子， 古示 的兒子 西番雅 。
ZEPH|1|2|耶和華說： 「我必從地面上徹底除滅萬物。
ZEPH|1|3|我必除滅人與牲畜， 除滅空中的鳥、海裏的魚、 絆腳石和惡人； 我必把人從地面上剪除， 這是耶和華說的。
ZEPH|1|4|我必伸手攻擊 猶大 和 耶路撒冷 所有的居民； 從這地方剪除剩下的 巴力 、 事奉偶像之祭司的名字與祭司；
ZEPH|1|5|還有那些在屋頂拜天上萬象的， 那些敬拜耶和華指著他起誓， 卻又指著 米勒公 起誓的；
ZEPH|1|6|並那些轉去不跟從耶和華， 不尋求耶和華，也不求問他的。」
ZEPH|1|7|在主耶和華面前要靜默無聲， 因為耶和華的日子快到了。 耶和華已經預備祭物， 將召來的人分別為聖。
ZEPH|1|8|「到了獻祭給耶和華的日子， 我要懲罰領袖和王子， 及所有穿外邦衣服的人。
ZEPH|1|9|到那日，我必懲罰所有跳過門檻， 以殘暴和詭詐塞滿主人房屋的人。
ZEPH|1|10|「當那日，從 魚門 必發出悲哀的聲音， 從第二城區發出哀號的聲音， 從山間發出破裂的大響聲。 這是耶和華說的。
ZEPH|1|11|瑪革提施 的居民哪，你們要哀號， 因為所有的商人 都滅亡了， 滿載銀子的人都被剪除。
ZEPH|1|12|那時，我必用燈巡查 耶路撒冷 ， 懲罰那些沉湎在酒渣上的人； 他們心裏說： 『耶和華必不降福，也不降禍。』
ZEPH|1|13|他們的財寶成為掠物， 房屋變為廢墟。 他們建造房屋，卻不得住在其內； 栽葡萄園，卻不得喝其中所出的酒。」
ZEPH|1|14|耶和華的大日臨近， 臨近而且甚快； 那是耶和華日子的風聲， 勇士必在那裏痛痛地哭號。
ZEPH|1|15|那日是憤怒的日子， 急難困苦的日子， 荒廢淒涼的日子， 黑暗幽冥的日子， 烏雲密佈的日子，
ZEPH|1|16|是吹角吶喊的日子， 要攻擊堅固的城， 攻擊高大的城樓。
ZEPH|1|17|我必使災禍臨到人身上， 使他們行走如同盲人， 因為他們得罪了耶和華； 他們的血必倒出如灰塵， 肉身拋棄如糞土。
ZEPH|1|18|當耶和華發怒的日子， 他們的金銀不能救自己； 耶和華妒忌的火必燒滅全地， 要向地上所有的居民施行可怕的毀滅。
ZEPH|2|1|不知羞恥的國民哪， 趁命令尚未發出， 日子流逝如糠秕， 耶和華的烈怒尚未臨到你們， 他發怒的日子未到以先， 你們應當聚集，聚集起來。
ZEPH|2|2|
ZEPH|2|3|世上遵守耶和華典章的謙卑人哪， 你們都當尋求耶和華， 尋求公義，尋求謙卑； 或許在耶和華發怒的日子得以隱藏。
ZEPH|2|4|迦薩 必遭遺棄 ， 亞實基倫 必然荒涼； 亞實突 人必在正午被趕出， 以革倫 也要連根拔除 。
ZEPH|2|5|禍哉，住沿海之地的 基利提 人！ 迦南 、 非利士 人之地啊，耶和華的話攻擊你們： 我必毀滅你，以致無人居住。
ZEPH|2|6|沿海之地要變為草場， 牧人的住處 和羊群的圈。
ZEPH|2|7|這地必為 猶大 家的餘民所得； 他們要在那裏放牧， 晚上躺臥在 亞實基倫 的房屋中； 因為耶和華－他們的上帝必眷顧他們， 使被擄的人歸回。
ZEPH|2|8|我聽見 摩押 毀謗， 亞捫 人辱罵； 他們辱罵我的百姓， 自誇自大，侵犯他們的疆土。」
ZEPH|2|9|萬軍之耶和華－ 以色列 的上帝說： 因此，我指著我的永生起誓： 摩押 必如 所多瑪 ， 亞捫 人必像 蛾摩拉 ， 都變為刺草、鹽坑、永遠荒廢之地。 我百姓中剩餘的必擄掠他們， 我國中的倖存者必得他們的地。
ZEPH|2|10|這事臨到他們是因他們的驕傲， 他們自誇自大， 辱罵萬軍之耶和華的百姓。
ZEPH|2|11|耶和華必向他們顯為可畏， 因他使地上的眾神衰微； 列國的海島各在自己的地方敬拜他。
ZEPH|2|12|你們 古實 人， 也是被我的刀所殺的。
ZEPH|2|13|耶和華要伸手攻擊北方， 毀滅 亞述 ， 使 尼尼微 荒涼， 乾旱如同曠野。
ZEPH|2|14|群畜，就是各類 的走獸必臥在其中， 鵜鶘和豪豬要宿在柱頂； 窗戶有鳴叫的聲音， 門檻毀壞 ， 他要毀壞香柏木板 。
ZEPH|2|15|這素來歡樂、安然居住的城， 心裏說：「惟有我，除我以外再沒有別的」， 現在竟然荒涼，成為野獸躺臥之處！ 凡經過的人都必搖著手嗤笑它。
ZEPH|3|1|禍哉，這欺壓的城！ 悖逆，污穢，
ZEPH|3|2|不聽從命令， 不領受訓誨， 不倚靠耶和華， 不親近它的上帝。
ZEPH|3|3|其中的領袖是咆哮的獅子， 審判官是晚上 的野狼， 不留一點到早晨。
ZEPH|3|4|它的先知是虛浮詭詐的人， 祭司褻瀆聖所，強解律法。
ZEPH|3|5|耶和華在它中間行公義， 斷不做非義的事， 每早晨顯明他的公義，無日不然； 只是不義的人不知羞恥。
ZEPH|3|6|「我已經除滅列國， 使他們的城樓荒廢。 我使他們街道荒涼， 無人經過； 他們的城鎮毀壞， 沒有人，沒有居民。
ZEPH|3|7|我說：『只要你敬畏我， 領受訓誨； 其住處就不會照我原先所定的被剪除 。』 然而，他們從早起來就在各樣事上敗壞自己。
ZEPH|3|8|「你們要等候我， 直到我興起擄掠 的日子； 因為我已定意招聚列邦，聚集列國， 將我的惱怒，我一切的烈怒，都傾倒在它們身上。 我妒忌的火必燒滅全地。 這是耶和華說的。
ZEPH|3|9|「那時，我要改變萬民， 使他們有清潔的嘴唇， 好求告耶和華的名， 同心合意事奉我。
ZEPH|3|10|那些向我祈求的， 我所分散的子民 ， 必從 古實河 的那一邊， 獻供物給我。
ZEPH|3|11|「當那日，你必不再因一切得罪我的事蒙羞， 因為那時我必從你中間除掉狂喜高傲的人， 在我的聖山上你也不再狂傲。
ZEPH|3|12|我卻要在你中間留下困苦貧寒的百姓， 他們必投靠耶和華的名。
ZEPH|3|13|以色列 的餘民必不行惡， 不說謊，口中沒有詭詐的舌頭； 他們吃喝躺臥， 無人使他們驚嚇。」
ZEPH|3|14|錫安 哪，應當歌唱！ 以色列 啊，應當歡呼！ 耶路撒冷 啊，應當滿心歡喜快樂！
ZEPH|3|15|耶和華已經免去對你的審判， 趕出你的仇敵。 以色列 的王－耶和華在你中間； 你必不再懼怕災禍。
ZEPH|3|16|當那日，必有話對 耶路撒冷 說： 「不要懼怕！ 錫安 哪，不要手軟！
ZEPH|3|17|耶和華－你的上帝在你中間 大有能力，施行拯救。 他必因你歡欣喜樂， 他在愛中靜默， 且因你而喜樂歡呼。
ZEPH|3|18|我要聚集那些因無節期而愁煩的人， 他們曾遠離你， 是你的重擔和羞辱 。
ZEPH|3|19|那時，看哪，我必對付所有苦待你的人， 拯救瘸腿的，召集被趕出的； 那些在全地受羞辱的， 我必使他們得稱讚，享名聲。
ZEPH|3|20|那時，我必領你們回來，召集你們； 我使你們被擄之人歸回的時候， 我必使你們在地上的萬民中享名聲，得稱讚； 這是耶和華說的。」
