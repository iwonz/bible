2KGS|1|1|亞哈 死後， 摩押 背叛 以色列 。
2KGS|1|2|亞哈謝 在 撒瑪利亞 ，一日從樓上的欄杆跌下來，就病了。於是他派使者，對他們說：「你們去問 以革倫 的神明 巴力‧西卜 ，我這病是否能痊癒。」
2KGS|1|3|但耶和華的使者對 提斯比 人 以利亞 說：「你起來，上去迎見 撒瑪利亞 王的使者，對他們說：『你們去問 以革倫 的神明 巴力‧西卜 ，是因為 以色列 中沒有上帝嗎？』
2KGS|1|4|所以耶和華如此說：『你必不能下你所上的床，因為你一定會死！』」 以利亞 就去了。
2KGS|1|5|使者回到王那裏，王對他們說：「你們為甚麼回來了呢？」
2KGS|1|6|他們對王說：「有一個人上來迎見我們，對我們說：『去，回到差你們來的王那裏，對他說：耶和華如此說，你派人去問 以革倫 的神明 巴力‧西卜 ，是因為 以色列 中沒有上帝嗎？所以你必不能下所上的床，你一定會死。』」
2KGS|1|7|王對他們說：「上來迎見你們，告訴你們這些話的人是甚麼樣子呢？」
2KGS|1|8|他們對王說：「這人身穿毛衣 ，腰束皮帶。」王說：「他一定是 提斯比 人 以利亞 。」
2KGS|1|9|於是，王派了一個五十夫長，帶領五十人到 以利亞 那裏。他上來，看哪， 以利亞 正坐在山頂上。五十夫長對他說：「神人哪，王吩咐你下來！」
2KGS|1|10|以利亞 回答五十夫長說：「我若是神人，願火從天上降下來，吞滅你和你的五十個人！」於是有火從天上降下來，吞滅五十夫長和他的五十個人。
2KGS|1|11|王又派另一個五十夫長，帶領五十人到 以利亞 那裏。五十夫長對他說：「神人哪，王這樣吩咐，快快下來！」
2KGS|1|12|以利亞 回答他們說：「我若是神人，願火從天上降下來，吞滅你和你的五十個人！」於是上帝的火 從天上降下來，吞滅五十夫長和他的五十個人。
2KGS|1|13|王第三次又派一個五十夫長，帶領五十人去。第三個五十夫長上去，雙膝跪在 以利亞 面前，哀求他說：「神人哪，願我的性命和你這五十個僕人的性命在你眼中看為寶貴！
2KGS|1|14|看哪，已經有火從天上降下來，吞滅前兩次來的五十夫長和他們的五十個人，現在願我的性命在你眼中看為寶貴！」
2KGS|1|15|耶和華的使者對 以利亞 說：「你跟他下去，不要怕他！」 以利亞 就起來，跟他下到王那裏去。
2KGS|1|16|他對王說：「耶和華如此說：『你派人去問 以革倫 的神明 巴力‧西卜 ，是因為 以色列 中沒有上帝可以讓你求問他的話嗎？所以你必不能下所上的床，你一定會死！』」
2KGS|1|17|亞哈謝 死了，正如耶和華藉 以利亞 所說的話。 猶大 王 約沙法 的兒子 約蘭 第二年， 亞哈謝 的兄弟 約蘭 接續他作王，因 亞哈謝 沒有兒子。
2KGS|1|18|亞哈謝 其餘所做的事，不都寫在《以色列諸王記》上嗎？
2KGS|2|1|耶和華要用旋風接 以利亞 升天的時候， 以利亞 與 以利沙 從 吉甲 往前行。
2KGS|2|2|以利亞 對 以利沙 說：「耶和華差遣我往 伯特利 去，你可以留在這裏。」 以利沙 說：「我指著永生的耶和華，又指著你的性命起誓，我必不離開你。」於是二人下到 伯特利 。
2KGS|2|3|在 伯特利 的先知的門徒出來，到 以利沙 那裏，對他說：「耶和華今日要接你的師父離開你 ，你知不知道？」他說：「我知道，你們不要作聲。」
2KGS|2|4|以利亞 對 以利沙 說：「耶和華差遣我往 耶利哥 去，你可以留在這裏。」 以利沙 說：「我指著永生的耶和華，又指著你的性命起誓，我必不離開你。」於是二人到了 耶利哥 。
2KGS|2|5|在 耶利哥 的先知的門徒來靠近 以利沙 ，對他說：「耶和華今日要接你的師父離開你，你知不知道？」他說：「我知道，你們不要作聲。」
2KGS|2|6|以利亞 對 以利沙 說：「耶和華差遣我往 約旦河 去，你可以留在這裏。」 以利沙 說：「我指著永生的耶和華，又指著你的性命起誓，我必不離開你。」於是二人一同往前行。
2KGS|2|7|有五十個先知的門徒同去，遠遠地站在他們對面；他們二人在 約旦河 邊站住。
2KGS|2|8|以利亞 捲起自己的外衣，用來打水，水就左右分開，二人走乾地過去。
2KGS|2|9|過去之後， 以利亞 對 以利沙 說：「我未被接去離開你以前，你要我為你做甚麼，只管求。」 以利沙 說：「願感動你的靈雙倍感動我。」
2KGS|2|10|以利亞 說：「你求的是一件難事。我被接去離開你的時候，你若看見我，就必得著；若不然，就得不著了。」
2KGS|2|11|他們邊走邊說話的時候，看哪，有火馬和火焰車出現，把二人隔開， 以利亞 就乘旋風升天去了。
2KGS|2|12|以利沙 看見，就呼叫說：「我父啊！我父啊！ 以色列 的戰車騎兵啊！」 以利沙 不再看見他的時候，就把自己的衣服撕為兩片。
2KGS|2|13|他拾起 以利亞 身上掉下來的外衣，回去站在 約旦河 邊。
2KGS|2|14|他用 以利亞 身上掉下來的外衣打水，說：「耶和華－ 以利亞 的上帝在哪裏呢？」打水之後，水也左右分開， 以利沙 就過去了。
2KGS|2|15|在 耶利哥 的先知的門徒從對面看見他，說：「感動 以利亞 的靈臨到 以利沙 身上了。」他們就來迎接他，俯伏於地，向他下拜，
2KGS|2|16|對他說：「看哪，僕人這裏有五十個壯士，請你讓他們去尋找你師父，或者耶和華的靈將他提起來，投在某山某谷。」 以利沙 說：「你們不必派人去。」
2KGS|2|17|他們再三催促，直到他不好意思，就說：「你們派人去吧！」他們就派了五十個人去，尋找了三天，也沒有找著他。
2KGS|2|18|以利沙 仍然留在 耶利哥 ，他們回到他那裏，他對他們說：「我不是告訴你們不必去嗎？」
2KGS|2|19|耶利哥城 的人對 以利沙 說：「看哪，這城的地勢美好，正如我主所看見的，只是水質惡劣，地也沒有生產。」
2KGS|2|20|以利沙 說：「你們拿一個新的瓶子來，裏面裝鹽。」他們就拿給他。
2KGS|2|21|他出去到了水源，把鹽倒在那裏，說：「耶和華如此說：『我治好了這水，從那裏不會再有死亡和不生產的事了。』」
2KGS|2|22|於是那水治好了，直到今日，正如 以利沙 所說的話。
2KGS|2|23|以利沙 從那裏上 伯特利 去。正上路的時候，有些孩童從城裏出來，譏笑他，對他說：「禿頭的，上去吧！禿頭的，上去吧！」
2KGS|2|24|他轉過身來瞪著他們，奉耶和華的名詛咒他們。於是有兩隻母熊從林中出來，撕裂他們當中的四十二個孩童。
2KGS|2|25|以利沙 從 伯特利 上 迦密山 ，又從那裏回到 撒瑪利亞 。
2KGS|3|1|猶大 王 約沙法 第十八年， 亞哈 的兒子 約蘭 在 撒瑪利亞 登基，作 以色列 王十二年。
2KGS|3|2|他行耶和華眼中看為惡的事，但不致像他父母所行的，因為他除掉他父所造 巴力 的柱像。
2KGS|3|3|然而，他依戀 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪，總不離開。
2KGS|3|4|摩押 王 米沙 牧養許多羊，曾向 以色列 王進貢十萬羔羊和十萬公綿羊的毛。
2KGS|3|5|亞哈 死後， 摩押 王背叛 以色列 王。
2KGS|3|6|那時 約蘭 王出 撒瑪利亞 ，數點 以色列 眾人。
2KGS|3|7|他向前行，派人到 猶大 王 約沙法 那裏，說：「 摩押 王背叛我，你肯同我去攻打 摩押 嗎？」 約沙法 說：「我肯上去，你我不分彼此，我的軍隊就是你的軍隊，我的馬就是你的馬。」
2KGS|3|8|然後 約沙法 說：「我們從哪條路上去呢？」 約蘭 說：「從 以東 曠野的路上去。」
2KGS|3|9|於是， 以色列 王和 猶大 王，以及 以東 王，都一同去。他們繞行了七日的路程，軍隊和所帶的牲畜都沒有水喝。
2KGS|3|10|以色列 王說：「哀哉！耶和華召集我們這三王，是要交在 摩押 人的手裏。」
2KGS|3|11|約沙法 說：「這裏不是有耶和華的先知嗎？我們可以託他求問耶和華。」 以色列 王的一個大臣回答說：「這裏有 沙法 的兒子 以利沙 ，就是從前服事 以利亞 的 。」
2KGS|3|12|約沙法 說：「他必有耶和華的話。」於是 以色列 王、 約沙法 和 以東 王都下去見他。
2KGS|3|13|以利沙 對 以色列 王說：「我跟你有甚麼關係呢？去問你父親的先知和你母親的先知吧！」 以色列 王對他說：「不，因為耶和華召集我們這三王，是要交在 摩押 人的手裏。」
2KGS|3|14|以利沙 說：「我指著所事奉永生的萬軍之耶和華起誓，我若不看 猶大 王 約沙法 的情面，必不理你，不睬你。
2KGS|3|15|現在你們給我找一個彈琴的人來。」彈琴的人彈奏的時候，耶和華的手就按在 以利沙 身上。
2KGS|3|16|他就說：「耶和華如此說：『你們要在這谷中到處挖溝。』
2KGS|3|17|因為耶和華如此說：『你們雖不見風，也不見雨，這谷卻必滿了水，使你們和你們的牛羊牲畜都有水喝。』
2KGS|3|18|在耶和華眼中這還算是小事，他也必將 摩押 人交在你們手中。
2KGS|3|19|你們必攻破一切堡壘和美好的城鎮，砍伐各種好樹，塞住一切水泉，用石頭毀壞一切良田。」
2KGS|3|20|到了早晨，約在獻祭的時候，看哪，有水從 以東 而來，遍地就滿了水。
2KGS|3|21|摩押 眾人聽見這三王上來要與他們打仗，凡能束上腰帶的，無論老少，都被召集站在邊界上。
2KGS|3|22|摩押 人清早起來，日光照在水上，他們看見對面水紅如血，
2KGS|3|23|就說：「這是血啊！必是三王互相擊殺，全都滅亡了。 摩押 人哪，我們現在去搶奪財物吧！」
2KGS|3|24|摩押 人到了 以色列 營， 以色列 人起來攻打他們，他們就在 以色列 人面前逃跑。 以色列 人追殺 摩押 人，直殺入 摩押 境內 。
2KGS|3|25|他們拆毀 摩押 的城鎮，各人拋石頭填滿一切良田，塞住一切水泉，砍伐各種好樹，只剩下 吉珥‧哈列設 的石牆，但甩石的兵仍然包圍攻打那城。
2KGS|3|26|摩押 王見戰事激烈，對他不利，就率領七百個拿刀的兵，想突圍逃到 以東 王那裏，卻沒有成功。
2KGS|3|27|於是他在城牆上，把那應當接續他作王的長子獻為燔祭。 有極大的憤怒臨到 以色列 ，於是三王離開 摩押 王，各自回本地去了。
2KGS|4|1|有個先知門徒的妻子哀求 以利沙 說：「你的僕人，我丈夫死了，他敬畏耶和華是你所知道的。現在有債主來，要帶走我的兩個孩子給他作奴隸。」
2KGS|4|2|以利沙 對她說：「我可以為你做甚麼呢？告訴我，你家裏有甚麼？」她說：「婢女家中除了一瓶油之外，甚麼也沒有。」
2KGS|4|3|以利沙 說：「你到外面去向所有的鄰舍借器皿，要空的器皿，不要少借。
2KGS|4|4|然後你回家，關上門，你和你兒子在裏面把油倒在所有的器皿裏，倒滿了就放在一邊。」
2KGS|4|5|於是婦人離開 以利沙 去了。她關上門，把自己和兒子關在家裏。他們把器皿拿給她，她就倒油。
2KGS|4|6|器皿都滿了，她對兒子說：「再給我拿器皿來。」兒子對她說：「沒有器皿了。」油就止住了。
2KGS|4|7|婦人去告訴神人，神人說：「你去賣了油還債，你和你兩個兒子可以靠著所剩的過活。」
2KGS|4|8|一日， 以利沙 經過 書念 ，在那裏有一個富有的婦人強留他吃飯。此後， 以利沙 每次經過就轉到那裏去吃飯。
2KGS|4|9|婦人對丈夫說：「看哪，我知道那常從我們這裏經過的是神聖的神人。
2KGS|4|10|我們可以為他蓋一間有牆的小閣樓，裏面安放床榻、桌子、椅子、燈臺。每當他來到我們這裏，就可以住在那裏。」
2KGS|4|11|一日， 以利沙 來到那裏，轉進那閣樓，躺臥在那裏。
2KGS|4|12|以利沙 吩咐僕人 基哈西 說：「你叫這 書念 婦人來。」他把婦人叫了來，婦人就站在 以利沙 面前。
2KGS|4|13|以利沙 吩咐僕人說：「你對她說：『看哪，你為我們費了許多心思，我可以為你做甚麼呢？我可以為你向王或元帥求甚麼呢？』」她說：「我已住在自己百姓之中。」
2KGS|4|14|以利沙 說：「究竟可以為她做甚麼呢？」 基哈西 說：「她真的沒有兒子，她丈夫也老了。」
2KGS|4|15|以利沙 說：「叫她回來。」於是他叫了她來，她就站在門口。
2KGS|4|16|以利沙 說：「明年這時候 ，你必抱一個兒子。」她說：「神人，我主啊，不要這樣欺哄婢女。」
2KGS|4|17|婦人果然懷孕，到了明年那時候，生了一個兒子，正如 以利沙 向她所說的。
2KGS|4|18|孩子長大，一日出去到他父親和收割的人那裏。
2KGS|4|19|他對父親說：「我的頭啊，我的頭啊！」他父親對僕人說：「把他抱到他母親那裏。」
2KGS|4|20|僕人抱去，交給他母親。孩子坐在母親的膝上，到中午就死了。
2KGS|4|21|他母親上去，把他放在神人的床上，關了門出來，
2KGS|4|22|呼叫她丈夫說：「你叫一個僕人給我牽一匹驢來，我要趕去見神人，然後回來。」
2KGS|4|23|丈夫說：「今日不是初一，也不是安息日，你為何要到他那裏去呢？」婦人說：「平安無事。」
2KGS|4|24|於是她備上驢，對僕人說：「走，趕緊走，除非我吩咐你，不要為了我而慢下來。」
2KGS|4|25|婦人往 迦密山 去，到了神人那裏。 神人遠遠看見她，對僕人 基哈西 說：「看哪， 書念 的婦人來了！
2KGS|4|26|現在你跑去迎接她，對她說，你平安嗎？你丈夫平安嗎？孩子平安嗎？」她說：「平安。」
2KGS|4|27|婦人上了山，到神人那裏，就抱住神人的腳。 基哈西 前來要推開她，神人說：「由她吧！因為她心裏愁苦。但耶和華向我隱瞞這事，沒有告訴我。」
2KGS|4|28|婦人說：「我何嘗向我主求過兒子呢？我豈不是說過，不要欺哄我嗎？」
2KGS|4|29|以利沙 吩咐 基哈西 說：「你束上腰，手拿我的杖前去。若遇見人，不要向他問安，人若向你問安，也不要回答。要把我的杖放在孩子臉上。」
2KGS|4|30|孩子的母親說：「我指著永生的耶和華，又指著你的性命起誓，我必不離開你。」於是 以利沙 起身，隨著她去了。
2KGS|4|31|基哈西 在他們以先去了，把杖放在孩子臉上，卻沒有聲音，也沒有動靜。 基哈西 回去，迎見 以利沙 ，告訴他說：「孩子還沒有醒過來。」
2KGS|4|32|以利沙 進了屋子，看哪，孩子死了，放在自己的床上。
2KGS|4|33|他進去，關上門，只有他們兩個人，他就向耶和華祈禱。
2KGS|4|34|他上去伏在孩子身上，口對口，眼對眼，手對手。他伏在孩子身上，孩子的身體就漸漸暖和了。
2KGS|4|35|然後他下來，在屋裏來回走了一趟，又上去伏在孩子身上。孩子打了七個噴嚏，眼睛就睜開了。
2KGS|4|36|以利沙 叫 基哈西 說：「你叫這 書念 婦人來。」於是他叫了她來。婦人來到 以利沙 那裏， 以利沙 說：「把你兒子抱起來。」
2KGS|4|37|婦人就進來，在 以利沙 腳前俯伏於地，向他下拜，然後抱起她兒子出去了。
2KGS|4|38|以利沙 回到 吉甲 ，那地正有饑荒。先知的門徒坐在他面前，他吩咐僕人說：「你把大鍋放在火上，給先知的門徒熬湯。」
2KGS|4|39|有一個人去到田野摘菜，發現一棵野瓜藤，就摘了滿滿一兜的野瓜回來，切了放進熬湯的鍋中，並不知道那是甚麼。
2KGS|4|40|他們把湯倒出來給大家吃。他們吃湯裏東西的時候，喊叫說：「神人哪，鍋子裏的東西會死人！」所以他們不能吃了。
2KGS|4|41|以利沙 說：「拿點麵來。」他把麵撒在鍋中，說：「倒出來，給大家吃吧！」鍋中就沒有毒了。
2KGS|4|42|有一個人從 巴力‧沙利沙 來，帶著初熟果子的食物、二十個大麥做的餅和新麥穗，裝在袋子裏送給神人。神人說：「把這些給大家吃。」
2KGS|4|43|僕人說：「這些豈可擺在一百人面前呢？」 以利沙 說：「你只管給大家吃吧！因為耶和華如此說，他們必吃了，還有剩下的。」
2KGS|4|44|僕人就擺在他們面前，他們吃了，還有剩下，正如耶和華所說的。
2KGS|5|1|亞蘭 王的元帥 乃縵 在他主人面前是一個偉大的人，得王的喜悅，因為耶和華曾藉他使 亞蘭 人得勝。他雖然是大能的勇士，卻染上了痲瘋 。
2KGS|5|2|亞蘭 人成群出征的時候，從 以色列 地擄了一個小女孩，她就服事 乃縵 的妻子。
2KGS|5|3|她對女主人說：「我希望主人去見 撒瑪利亞 的先知，他必能治好主人的痲瘋。」
2KGS|5|4|乃縵 去告訴他主人說，從 以色列 地來的女孩如此如此說。
2KGS|5|5|亞蘭 王說：「你可以去，我也會送信給 以色列 王。」於是 乃縵 手裏帶十他連得銀子、六千舍客勒金子和十套衣裳去了。
2KGS|5|6|他帶著這信給 以色列 王，說：「現在你接到這信，看哪，我派臣僕 乃縵 到你這裏來，你要治好他的痲瘋。」
2KGS|5|7|以色列 王讀了信就撕裂衣服，說：「我豈是上帝，能使人死使人活呢？這人竟派人來，叫我治好一個人的痲瘋。你們要知道，看，這人是找機會來跟我吵架的。」
2KGS|5|8|神人 以利沙 聽見 以色列 王撕裂衣服，就派人到王那裏，說：「你為甚麼撕裂衣服呢？讓那人到我這裏來，他會知道 以色列 中有先知。」
2KGS|5|9|於是 乃縵 帶著車馬到了 以利沙 的家，站在門前。
2KGS|5|10|以利沙 派一個使者，對 乃縵 說：「去，在 約旦河 中沐浴七次，你的肉就必復原，你會得潔淨。」
2KGS|5|11|乃縵 卻發怒走了。他說：「看哪，我以為他必定會出來，到我這裏，站著求告耶和華－他上帝的名，在患處上搖手，治好這痲瘋。
2KGS|5|12|大馬士革 的 亞瑪拿河 和 法珥法河 豈不比 以色列 的一切水更好嗎？我難道不可以在那裏沐浴而得潔淨嗎？」於是他生氣，轉身走了。
2KGS|5|13|他的僕人近前來，對他說：「我父啊，先知若吩咐你做一件大事，你豈不做嗎？何況是吩咐你去沐浴，得潔淨呢？」
2KGS|5|14|於是 乃縵 下去，照著神人的話，在 約旦河 裏浸了七次。他的肉復原，好像小孩的肉，他就潔淨了。
2KGS|5|15|乃縵 帶著所有跟隨他的人，回到神人那裏，站在他面前，說：「看哪，我知道，除了 以色列 ，全地沒有上帝。現在請你收下僕人的禮物。」
2KGS|5|16|以利沙 說：「我指著所事奉永生的耶和華起誓，我必不接受。」 乃縵 再三請他收下，他卻不肯。
2KGS|5|17|乃縵 說：「你若不肯，請把兩匹騾子能馱的土賜給僕人，僕人必不再把燔祭或祭物獻給別神，只獻給耶和華。
2KGS|5|18|惟有一件事，願耶和華饒恕你僕人：我主人進 臨門 廟在那裏叩拜的時候，他總是扶著我的手，所以我也在 臨門 廟叩拜。我在 臨門 廟叩拜的這事，願耶和華饒恕你僕人。」
2KGS|5|19|以利沙 對他說：「你平安地回去吧！」 乃縵 離開他去了。走了一小段路，
2KGS|5|20|神人 以利沙 的僕人 基哈西 說：「看哪，我主人不願從這 亞蘭 人 乃縵 手裏接受他帶來的禮物，我指著永生的耶和華起誓，我必跑去追上他，向他拿些東西。」
2KGS|5|21|於是 基哈西 去追 乃縵 。 乃縵 看見有人追來，就下車迎著他，說：「都平安嗎？」
2KGS|5|22|他說：「都平安！我主人派我來說：『看哪，現在有兩個年輕人，是先知的門徒，從 以法蓮 山區來到我這裏，請你給他們一他連得銀子，兩套衣裳。』」
2KGS|5|23|乃縵 說：「好啊，請收下二他連得。」他再三請求，就把二他連得銀子裝在兩個袋子裏，連同兩套衣裳交給兩個僕人；他們就在 基哈西 前頭抬著走。
2KGS|5|24|到了山岡， 基哈西 從他們手中接過來，放在屋裏，打發這些人走了。
2KGS|5|25|基哈西 進去，站在主人面前。 以利沙 對他說：「 基哈西 ，你從哪裏來？」他說：「僕人哪裏也沒去。」
2KGS|5|26|以利沙 對他說：「那人下車轉過來迎著你的時候，我的心豈沒有去呢？這豈是接受銀子，接受衣裳、橄欖園、葡萄園、牛羊、僕婢的時候呢？
2KGS|5|27|因此， 乃縵 的痲瘋必緊隨你和你的後裔，直到永遠。」 基哈西 從 以利沙 面前出去，就長了痲瘋，像雪一樣。
2KGS|6|1|先知的門徒對 以利沙 說：「看哪，我們在你面前居住的地方，那裏對我們太窄小了。
2KGS|6|2|讓我們往 約旦河 去，各人從那裏取一根木料，在那裏為自己建造居住的地方。」他說：「你們去吧！」
2KGS|6|3|有一人說：「請你與僕人同去。」他說：「我可以去。」
2KGS|6|4|於是 以利沙 與他們同去。到了 約旦河 ，他們砍伐樹木。
2KGS|6|5|有一人砍樹的時候，斧子的頭掉在水裏，他就喊著說：「不好了！我主啊，斧子是借來的。」
2KGS|6|6|神人說：「掉在哪裏了？」他把那地方指給 以利沙 看。 以利沙 砍了一塊木頭，拋在水裏，就使斧子的頭浮上來了。
2KGS|6|7|以利沙 說：「拿起來吧！」那人就伸手拿起來了。
2KGS|6|8|亞蘭 王與 以色列 作戰，他和臣僕商議說：「我要在某處某處安營 。」
2KGS|6|9|神人派人到 以色列 王那裏，說：「你要小心，不要從某處經過，因為 亞蘭 人下到那裏去了。」
2KGS|6|10|以色列 王派人到神人告訴他的地方去。神人警告他，他就在那裏有所防備，不止一兩次。
2KGS|6|11|亞蘭 王因這事心裏氣憤，召了臣僕來，對他們說：「我們當中有誰幫助 以色列 王，你們不告訴我嗎？」
2KGS|6|12|有一個臣僕說：「不，我主，我王！只有 以色列 中的先知 以利沙 ，把王在臥房所說的話告訴 以色列 王。」
2KGS|6|13|王說：「你們去查看他在哪裏，我好派人去捉拿他。」有人告訴王說：「看哪，他在 多坍 。」
2KGS|6|14|王就派遣車馬和大軍往那裏去，夜間他們到了，圍困那城。
2KGS|6|15|神人的僕人清早起來出去，看哪，車馬軍兵圍困了城。僕人對神人說：「不好了！我主啊，我們該怎麼辦呢？」
2KGS|6|16|神人說：「不要懼怕！因與我們同在的比與他們同在的更多。」
2KGS|6|17|以利沙 禱告說：「耶和華啊，求你開他的眼目，使他能看見。」耶和華開了這年輕人的眼目，他就看見了，看哪，滿山有火馬和火焰車圍繞 以利沙 。
2KGS|6|18|亞蘭 人下到 以利沙 那裏， 以利沙 向耶和華禱告說：「求你擊打這國，使他們眼目失明。」耶和華就照 以利沙 的話，擊打他們，使他們眼目失明。
2KGS|6|19|以利沙 對他們說：「這不是那條路，也不是那座城。你們跟我走，我必領你們到你們要尋找的人那裏。」於是他領他們到了 撒瑪利亞 。
2KGS|6|20|他們進了 撒瑪利亞 ， 以利沙 說：「耶和華啊，求你開這些人的眼目，使他們能看見。」耶和華開了他們的眼目，他們就看見了，看哪，是在 撒瑪利亞城 中。
2KGS|6|21|以色列 王看見他們，就對 以利沙 說：「我父啊，我真的可以擊殺他們嗎？」
2KGS|6|22|他說：「不可擊殺！這些人豈是你用刀用弓擄來給你擊殺的呢？當在他們面前擺設飲食給他們吃喝，讓他們回到他們主人那裏。」
2KGS|6|23|王為他們預備了盛大的宴席。他們吃喝完了，王就送他們回到他們主人那裏。此後， 亞蘭 的軍隊不再侵犯 以色列 地了。
2KGS|6|24|此後， 亞蘭 王 便‧哈達 召集他的全軍，上來圍困 撒瑪利亞 。
2KGS|6|25|看哪，被圍困的時候， 撒瑪利亞 有大饑荒，甚至一個驢頭值八十舍客勒，四分之一卡布 的鴿子糞值五舍客勒。
2KGS|6|26|一日， 以色列 王在城牆上經過，有一個婦人向他呼叫說：「我主，我王啊！求你幫助。」
2KGS|6|27|王說：「耶和華不幫助你，我從哪裏幫助你呢？是從禾場，或從壓酒池嗎？」
2KGS|6|28|王對婦人說：「你有甚麼事？」她說：「這婦人對我說：『把你的兒子交出來，我們今日可以吃他，明日可以吃我的兒子。』
2KGS|6|29|我們就煮了我的兒子吃了。次日我對她說：『要把你的兒子交出來，我們可以吃。』她卻把她的兒子藏起來。」
2KGS|6|30|王聽見婦人的話，就撕裂衣服；那時，王在城牆上經過，百姓看見了，看哪，王貼身穿著麻布。
2KGS|6|31|王說：「我今日若容許 沙法 的兒子 以利沙 的頭還留在他身上，願上帝重重懲罰我！」
2KGS|6|32|那時， 以利沙 正坐在家中，有長老與他同坐。王派一個人先去，使者還沒有到， 以利沙 對長老說：「你們看，這兇手之子派人來斬我的頭。你們注意，當使者來到，你們就關上門，把他關在門外。在他後頭不就是他主人的腳步聲嗎？」
2KGS|6|33|正與他們說話的時候，看哪，使者 下到他那裏，說：「看哪，這災禍是從耶和華來的，我何必再仰望耶和華呢？」
2KGS|7|1|以利沙 說：「你們要聽耶和華的話，耶和華如此說：明日約這時候，在 撒瑪利亞 城門口，一細亞細麵只賣一舍客勒，二細亞大麥也賣一舍客勒。」
2KGS|7|2|有一個攙扶王的軍官回答神人說：「看哪，即使耶和華打開天上的窗戶，也不可能有這事。」 以利沙 說：「看哪，你必親眼看見，在那裏卻吃不到甚麼。」
2KGS|7|3|在城門口有四個長痲瘋的人，他們彼此說：「我們為何坐在這裏等死呢？
2KGS|7|4|我們若說要進城去，城裏有饑荒，我們必死在那裏。若我們在這裏坐著不動，也必死。現在，來吧，我們去向 亞蘭 人的軍隊投降。若他們饒我們的命，我們就活著；若殺我們，我們就死吧！」
2KGS|7|5|黃昏的時候，他們起來往 亞蘭 人的軍營去；到了營邊，看哪，沒有一人在那裏。
2KGS|7|6|因為主使 亞蘭 人的軍隊聽見戰車戰馬的聲音，大軍的聲音，他們就彼此說：「看哪，這必是 以色列 王雇用 赫 人諸王和 埃及 諸王來攻擊我們。」
2KGS|7|7|所以，在黃昏的時候他們起來逃跑，撇下帳棚、馬、驢，把軍營留在原處，只顧逃命。
2KGS|7|8|那些長痲瘋的人到了營邊，進了一座帳棚，吃了喝了，從當中拿走金銀和衣服，收藏起來。他們又回來，進了另一座帳棚，從當中拿走財物去收藏。
2KGS|7|9|那時，他們彼此說：「我們所做的不對了！這一天是有好消息的日子，我們竟不作聲！若等到天亮，我們就有罪了。現在，來，我們去向王室報信吧！」
2KGS|7|10|他們就去叫守城門的人，告訴他們說：「我們到了 亞蘭 人的軍營，看哪，沒有一人在那裏，也無人聲，只有拴著的馬和驢，帳棚都留在原處。」
2KGS|7|11|守城門的人就呼叫，他們向城內的王室報信。
2KGS|7|12|王夜間起來，對臣僕說：「我告訴你們 亞蘭 人向我們做的事。他們知道我們飢餓，所以離營，埋伏在田野，說：『 以色列 人出城的時候，我們活捉他們，我們就可以進到城裏去。』」
2KGS|7|13|王的一個臣僕回答說：「不如叫人從城裏剩下的馬中取五匹，看哪，這些馬像 以色列 大眾一樣 ，快要滅亡了；我們派人去窺探吧！」
2KGS|7|14|於是他們取了兩輛車和馬，王派人去跟蹤 亞蘭 人的軍隊，說：「你們去窺探吧。」
2KGS|7|15|他們去跟蹤 亞蘭 人，直到 約旦河 。看哪，整條路上都是 亞蘭 人匆忙逃跑時所丟棄的衣服和器具，使者就回來向王報告。
2KGS|7|16|百姓就出去，擄掠 亞蘭 人的軍營。於是一細亞細麵只賣一舍客勒，二細亞大麥也賣一舍客勒，正如耶和華所說的。
2KGS|7|17|王派攙扶他的那軍官在城門指揮，百姓在城門把他踩死了，正如神人在王下到他那裏的時候所說的。
2KGS|7|18|神人曾對王說：「明日約這時候，在 撒瑪利亞 城門口，二細亞大麥只賣一舍客勒，一細亞細麵也賣一舍客勒。」
2KGS|7|19|那軍官回答神人說：「看哪，即使耶和華打開天上的窗戶，也不可能有這事。」神人說：「看哪，你必親眼看見，在那裏卻吃不到甚麼。」
2KGS|7|20|這話果然應驗在他身上，因為百姓在城門把他踩死了。
2KGS|8|1|以利沙 曾對他救活的孩子的母親說：「你和你的全家要起身，往你可住的地方去住，因為耶和華已令饑荒降在這地七年。」
2KGS|8|2|婦人就起身，照神人的話去做，帶著全家往 非利士 人的地去，寄居了七年。
2KGS|8|3|過了七年，那婦人從 非利士 人的地回來，就出去為自己的房屋田地哀求王。
2KGS|8|4|那時王正與神人的僕人 基哈西 談話，說：「你把 以利沙 所做的一切大事告訴我。」
2KGS|8|5|基哈西 告訴王 以利沙 如何使死人復活，看哪， 以利沙 所救活的孩子的母親正為自己的房屋田地來哀求王。 基哈西 說：「我主我王，這就是那婦人，這是她的兒子，就是 以利沙 所救活的。」
2KGS|8|6|王問那婦人，她就把事情告訴王。於是王為她派一個官員，說：「凡屬這婦人的都還給她，自從她離開本地直到今日，她田地的出產也都還給她。」
2KGS|8|7|以利沙 來到 大馬士革 ， 亞蘭 王 便‧哈達 正患病。有人告訴王說：「神人來到這裏了。」
2KGS|8|8|王就吩咐 哈薛 說：「你帶著禮物去見神人，託他求問耶和華，我這病能不能好？」
2KGS|8|9|於是 哈薛 用四十匹駱駝，馱著 大馬士革 的各樣美物為禮物，去迎見 以利沙 。 哈薛 到了那裏，站在他面前，說：「你兒子 亞蘭 王 便‧哈達 派我到你這裏，問說：『我這病會不會好？』」
2KGS|8|10|以利沙 對 哈薛 說：「你回去告訴他說：『你一定會好。』但耶和華指示我，他必定會死。」
2KGS|8|11|神人定睛看著 哈薛 ，直到他感到羞愧。神人就哭了。
2KGS|8|12|哈薛 說：「我主為甚麼哭？」他說：「因為我知道你必虐待 以色列 人，用火焚燒他們的堡壘，用刀殺死他們的壯丁，摔死他們的嬰孩，剖開他們的孕婦。」
2KGS|8|13|哈薛 說：「僕人算甚麼，不過是一條狗，怎麼能行這大事呢？」 以利沙 說：「耶和華指示我，你必作 亞蘭 王。」
2KGS|8|14|哈薛 離開 以利沙 ，回到他主人那裏。主人對他說：「 以利沙 對你說了甚麼？」他說：「他告訴我你必能好。」
2KGS|8|15|次日， 哈薛 拿被子浸在水中，蒙住王的臉，王就死了。於是 哈薛 篡了他的位。
2KGS|8|16|亞哈 的兒子 以色列 王 約蘭 第五年－ 約沙法 曾作 猶大 王 － 猶大 王 約沙法 的兒子 約蘭 登基作了 猶大 王。
2KGS|8|17|約蘭 登基的時候年三十二歲，在 耶路撒冷 作王八年。
2KGS|8|18|他行 以色列 諸王的道，正如 亞哈 家所行的，因他娶了 亞哈 的女兒為妻，行耶和華眼中看為惡的事。
2KGS|8|19|耶和華卻因他僕人 大衛 的緣故，不肯滅絕 猶大 ，要照他所應許的，永遠賜燈光給 大衛 和他的子孫。
2KGS|8|20|約蘭 在位期間， 以東 背叛，自己立王治理他們，脫離 猶大 的權勢。
2KGS|8|21|約蘭 率領他所有的戰車過到 撒益 去。他夜間起來，攻打圍困他的 以東 人和戰車長； 猶大 軍兵逃跑，各回自己的帳棚去了；
2KGS|8|22|這樣， 以東 背叛，脫離 猶大 的管轄，直到今日。那時 立拿 也背叛了。
2KGS|8|23|約蘭 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|8|24|約蘭 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 亞哈謝 接續他作王。
2KGS|8|25|亞哈 的兒子 以色列 王 約蘭 第十二年， 猶大 王 約蘭 的兒子 亞哈謝 登基。
2KGS|8|26|他登基的時候年二十二歲，在 耶路撒冷 作王一年。他母親名叫 亞她利雅 ，是 以色列 王 暗利 的孫女。
2KGS|8|27|亞哈謝 行 亞哈 家的道，行耶和華眼中看為惡的事，與 亞哈 家一樣，因為他是 亞哈 家的女婿。
2KGS|8|28|他與 亞哈 的兒子 約蘭 同往 基列 的 拉末 去，與 亞蘭 王 哈薛 交戰。 亞蘭 人打傷了 約蘭 ，
2KGS|8|29|約蘭 王回到 耶斯列 ，醫治在 拉末 與 亞蘭 王 哈薛 打仗時，被 亞蘭 人擊打所受的傷。 約蘭 的兒子 猶大 王 亞哈謝 因為 亞哈 的兒子 約蘭 病了，就下到 耶斯列 看望他。
2KGS|9|1|以利沙 先知叫了一個先知的門徒來，吩咐他：「你束上腰，手拿這瓶膏油往 基列 的 拉末 去。
2KGS|9|2|你到了那裏，要在那裏尋找 寧示 的孫子， 約沙法 的兒子 耶戶 。你去，使他從弟兄中起來，帶他進最裏面的內室，
2KGS|9|3|把瓶裏的膏油倒在他頭上，說：『耶和華如此說：我膏你作 以色列 王。』然後你就開門逃跑，不要等候。」
2KGS|9|4|於是那青年，那年輕的先知往 基列 的 拉末 去了。
2KGS|9|5|他到了那裏，看哪，眾軍官都坐著，就說：「長官，我有話對你說。」 耶戶 說：「你要對我們哪一個說呢？」他說：「長官，我要對你說。」
2KGS|9|6|耶戶 就起來，進了內室，那青年把膏油倒在他頭上，對他說：「耶和華－ 以色列 的上帝如此說：『我膏你作耶和華百姓 以色列 的王。
2KGS|9|7|你要擊殺你主人 亞哈 的全家，我好在 耶洗別 身上，為我僕人眾先知和耶和華所有僕人的血伸冤。
2KGS|9|8|亞哈 全家都必滅亡，凡屬 亞哈 的男丁，無論是奴役的、自由的，我必從 以色列 中剪除。
2KGS|9|9|我必使 亞哈 的家像 尼八 兒子 耶羅波安 的家，又像 亞希雅 兒子 巴沙 的家。
2KGS|9|10|至於 耶洗別 ，狗必在 耶斯列 田裏吃她，無人埋葬。』」於是那青年就開門逃跑了。
2KGS|9|11|耶戶 出來，回到他主人的臣僕那裏，有一人問他說：「平安嗎？這瘋狂的人為甚麼到你這裏來呢？」他對他們說：「你們認得那人，也知道他在胡說。」
2KGS|9|12|他們說：「說謊！告訴我們吧。」他說：「他如此如此對我說：『耶和華如此說：我膏你作 以色列 的王。』」
2KGS|9|13|他們各人就急忙把自己的衣服鋪在臺階的上層，在 耶戶 的下面；他們吹角，說：「 耶戶 作王了！」
2KGS|9|14|這樣， 寧示 的孫子， 約沙法 的兒子 耶戶 背叛了 約蘭 。先前 約蘭 和 以色列 眾人因為 亞蘭 王 哈薛 的緣故，把守 基列 的 拉末 。
2KGS|9|15|後來 約蘭 王回到 耶斯列 ，醫治他與 亞蘭 王 哈薛 打仗時，被 亞蘭 人擊打所受的傷。 耶戶 說：「若你們有這樣的意思，就不要讓人溜出城，到 耶斯列 去報信。」
2KGS|9|16|於是 耶戶 駕戰車往 耶斯列 去，因為 約蘭 臥病在那裏。 猶大 王 亞哈謝 已經下去看望他。
2KGS|9|17|有一個守望的人站在 耶斯列 的城樓上，看見 耶戶 帶著一隊人來，就說：「我看見一隊人。」 約蘭 說：「派一個騎兵去迎接他們，問說：『平安嗎？』」
2KGS|9|18|騎兵就去迎接 耶戶 ，說：「王如此說：『平安嗎？』」耶戶說：「平安不平安跟你有甚麼關係呢？轉身跟在我後面吧！」守望的人說：「使者到了他們那裏，卻不回來。」
2KGS|9|19|王又派第二個騎兵去。這人到了他們那裏，說：「王如此說：『平安嗎？』」 耶戶 說：「平安不平安跟你有甚麼關係呢？轉身跟在我後面吧！」
2KGS|9|20|守望的人又說：「他到了他們那裏，也不回來。車駕得很兇猛，好像 寧示 的孫子 耶戶 在駕車。」
2KGS|9|21|約蘭 吩咐說：「套車！」人就給他套車。 以色列 王 約蘭 和 猶大 王 亞哈謝 各坐自己的車出去迎接 耶戶 ，在 耶斯列 人 拿伯 的田那裏遇見他。
2KGS|9|22|約蘭 見 耶戶 就說：「 耶戶 ，平安嗎？」 耶戶 說：「你母親 耶洗別 的淫行邪術這樣多，怎麼能平安呢？」
2KGS|9|23|約蘭 用手轉過車來逃跑，對 亞哈謝 說：「 亞哈謝 啊，反了！」
2KGS|9|24|耶戶 全力拉弓，射中 約蘭 兩臂中間，箭從心窩穿出， 約蘭 就仆倒在車上。
2KGS|9|25|耶戶 對他的軍官 畢甲 說：「把他拋在 耶斯列 人 拿伯 的田裏。你當記得，你我一同駕車跟隨他父親 亞哈 的時候，耶和華對 亞哈 說了預言，
2KGS|9|26|耶和華說：『我昨日看見 拿伯 的血和他眾子的血，我發誓我必在這塊田上報應你。』這是耶和華說的。現在你要照著耶和華的話，把他拋在這田裏。」
2KGS|9|27|猶大 王 亞哈謝 看見了，就沿著 伯．哈干 的路逃跑。 耶戶 追趕他，說：「把這人也擊殺在車上，在靠近 以伯蓮 的 姑珥 坡上 。」他逃到 米吉多 ，就死在那裏。
2KGS|9|28|他的臣僕用車把他的屍體運回 耶路撒冷 ，與他祖先同葬在 大衛城 ，他自己的墳墓裏。
2KGS|9|29|亞哈 的兒子 約蘭 第十一年， 亞哈謝 登基作了 猶大 王。
2KGS|9|30|耶戶 到了 耶斯列 。 耶洗別 聽見了，就畫眼影、梳頭，從窗戶往外觀看。
2KGS|9|31|耶戶 進了城門， 耶洗別 說：「殺主人的 心利 啊，平安嗎？」
2KGS|9|32|耶戶 向窗戶抬頭，說：「有誰順從我？誰？」有兩三個太監向外看他。
2KGS|9|33|耶戶 說：「把她拋下來！」他們就把她拋下來。她的血濺在牆上和馬上， 耶戶 踐踏在她身上。
2KGS|9|34|耶戶 進去，吃了喝了，說：「你們去處理這被詛咒的婦人，埋了她，因為她是王的女兒。」
2KGS|9|35|他們去了，要埋葬她，卻只找到她的頭骨和腳，以及手掌。
2KGS|9|36|他們回來報告 耶戶 ， 耶戶 說：「這正應驗耶和華藉他僕人 提斯比 人 以利亞 所說的話，說：『在 耶斯列 田裏，狗必吃 耶洗別 的肉，
2KGS|9|37|耶洗別 的屍體必在 耶斯列 田裏的地面上如同糞土，甚至沒有人可說：這是 耶洗別 。』」
2KGS|10|1|亞哈 有七十個兒子在 撒瑪利亞 。 耶戶 寫信送到 撒瑪利亞 ，給 耶斯列 的領袖和長老 ，以及教養 亞哈 眾兒子的人，說：
2KGS|10|2|「你們主人的眾兒子既然在你們那裏，你們又有戰車、馬匹、兵器、堅固城，現在你們接了這信，
2KGS|10|3|可以在你們主人的眾兒子中選一個賢能正直的，使他坐他父親的王位，你們也可以為你們主人的家作戰。」
2KGS|10|4|他們卻非常懼怕，說：「看哪，兩個王在他面前尚且站立不住，我們怎能站立得住呢？」
2KGS|10|5|王宮總管、市長和長老，並教養眾兒子的人，派人到 耶戶 那裏，說：「我們是你的僕人，凡你所吩咐的，我們都必遵行。我們不立誰作王，你看怎樣好就怎樣做吧。」
2KGS|10|6|耶戶 寫第二封信給他們，說：「你們若歸順我，聽從我的話，明日這時候，要帶著你們主人眾兒子的首級，來到 耶斯列 我這裏。」那時王的兒子七十人都住在城中教養他們的那些尊貴人家裏。
2KGS|10|7|信一到他們那裏，他們就把王的七十個兒子殺了，將首級裝在筐裏，送到 耶斯列 ， 耶戶 那裏。
2KGS|10|8|有使者來告訴 耶戶 說：「他們把王眾兒子的首級送來了。」 耶戶 說：「把首級分成兩堆，放在城門口，直到早晨。」
2KGS|10|9|次日早晨， 耶戶 出來，站著對眾百姓說：「你們都是公義的！看哪，我背叛了我的主人，把他殺了，但這所有的人又是誰殺的呢？
2KGS|10|10|由此可知，耶和華指著 亞哈 家所說的話一句也沒有落空，因為耶和華實現了他藉他僕人 以利亞 所說的話。」
2KGS|10|11|凡 亞哈 家在 耶斯列 所剩下的，他的大臣、密友、祭司， 耶戶 全都殺了，沒有留下一個倖存者。
2KGS|10|12|耶戶 起身往 撒瑪利亞 去。路途中，在牧人聚集的 伯．艾克特 ，
2KGS|10|13|耶戶 遇見 猶大 王 亞哈謝 的兄弟，說：「你們是誰？」他們說：「我們是 亞哈謝 的兄弟，現在下去要向王和太后的眾兒子問安。」
2KGS|10|14|耶戶 說：「活捉他們！」人就活捉了他們，把他們殺在 伯．艾克特 的坑邊，共四十二人，一個也沒有留下。
2KGS|10|15|耶戶 從那裏往前行，遇見 利甲 的兒子 約拿達 來迎接他， 耶戶 向他問安，對他說：「你的心 ，像我的心待你的心那樣正直嗎？」 約拿達 說：「是。」 耶戶 說：「若是這樣，請你伸出手來。」他伸出手， 耶戶 就拉他上車。
2KGS|10|16|耶戶 說：「你和我同去，看我為耶和華怎樣熱心。」於是他們請他坐在車上。
2KGS|10|17|到了 撒瑪利亞 ， 耶戶 把 亞哈 家在 撒瑪利亞 剩下的人全都殺了，直到滅盡，正如耶和華對 以利亞 所說的話。
2KGS|10|18|耶戶 召集眾百姓，對他們說：「 亞哈 事奉 巴力 還不夠熱心， 耶戶 更要熱心。
2KGS|10|19|現在你們召集 巴力 的眾先知和所有拜 巴力 的人，以及 巴力 的眾祭司，都到我這裏來，一個也不可缺少，因為我要給 巴力 獻大祭；凡不來的必不得活。」 耶戶 行詭詐，為要消滅拜 巴力 的人。
2KGS|10|20|耶戶 說：「要為 巴力 召集嚴肅會！」於是他們宣告了。
2KGS|10|21|耶戶 派人走遍 以色列 ；凡拜 巴力 的人都來齊了，沒有留下一個不來的。他們進了 巴力 廟， 巴力 廟中前後都擠滿了人。
2KGS|10|22|耶戶 對掌管服裝的人說：「拿出袍子來，給所有拜 巴力 的人穿。」他就拿出禮服來給了他們。
2KGS|10|23|耶戶 和 利甲 的兒子 約拿達 進了 巴力 廟，對拜 巴力 的人說：「你們要搜查察看，不可以有耶和華的僕人在你們這裏，只可以有拜 巴力 的人。」
2KGS|10|24|他們進去，獻上祭物和燔祭． 耶戶 先安排八十人在廟外，說：「我把這些人交在你們手中，誰放走其中一人，誰就要以命償命！」
2KGS|10|25|耶戶 獻完了燔祭，就對護衛兵和眾軍官說：「進去殺他們，不要讓一人逃脫！」護衛兵和軍官用刀殺了他們，將屍體拋出去，然後進入 巴力 廟的堡壘，
2KGS|10|26|將 巴力 廟中的柱像都 拿出來焚燒。
2KGS|10|27|他們毀壞 巴力 的柱像，拆毀了 巴力 廟當廁所，直到今日。
2KGS|10|28|這樣， 耶戶 在 以色列 中消滅了 巴力 。
2KGS|10|29|只是 耶戶 不離開 尼八 的兒子 耶羅波安 使 以色列 人陷入罪裏的那罪，就是拜 伯特利 和 但 的金牛犢。
2KGS|10|30|耶和華對 耶戶 說：「因你辦好我眼中看為正的事，照我的心意待 亞哈 家，你的子孫必接續你坐 以色列 的王位，直到第四代。」
2KGS|10|31|只是 耶戶 不盡心遵守耶和華－ 以色列 上帝的律法，不離開 耶羅波安 使 以色列 人陷入罪裏的那罪。
2KGS|10|32|在那些日子，耶和華開始削弱 以色列 。 哈薛 在 以色列 各邊界攻擊他們，
2KGS|10|33|就是 約旦河 東 基列 全地，從靠近 亞嫩谷 邊的 亞羅珥 起，包括 基列 和 巴珊 ，就是 迦得 人、 呂便 人、 瑪拿西 人的地。
2KGS|10|34|耶戶 其餘的事，凡他所做的和他英勇的事蹟，不都寫在《以色列諸王記》上嗎？
2KGS|10|35|耶戶 與他祖先同睡，葬在 撒瑪利亞 ，他兒子 約哈斯 接續他作王。
2KGS|10|36|耶戶 在 撒瑪利亞 作 以色列 王二十八年。
2KGS|11|1|亞哈謝 的母親 亞她利雅 見她兒子死了，就起來剿滅王室所有的後裔。
2KGS|11|2|但 約蘭 王的女兒， 亞哈謝 的妹妹 約示巴 ，將 亞哈謝 的兒子 約阿施 從被殺的王子中偷出來，把他和他的奶媽藏在臥房裏，躲避了 亞她利雅 ，沒有被殺。
2KGS|11|3|亞她利雅 治理這地的時候， 約阿施 和他的奶媽在耶和華的殿裏藏了六年。
2KGS|11|4|第七年， 耶何耶大 派人叫 迦利 人和護衛兵的眾百夫長來，領他們進耶和華的殿，與他們立約，使他們在耶和華殿裏起誓，又把王的兒子指給他們看，
2KGS|11|5|吩咐他們說：「你們要這樣做：你們當中在安息日值班的，三分之一要把守王宮，
2KGS|11|6|三分之一要在 蘇珥門 ，三分之一要在護衛兵院的後門；你們要這樣輪流把守王宮。
2KGS|11|7|你們安息日所有不值班的兩隊人員要在耶和華的殿裏護衛王；
2KGS|11|8|各人手拿兵器，四圍保護王。凡擅自闖入你們行列的，要被處死。王出入的時候，你們當跟隨他。」
2KGS|11|9|眾百夫長就照著 耶何耶大 祭司一切所吩咐的去做，各帶自己的人，無論安息日值班或不值班的，都到 耶何耶大 祭司那裏。
2KGS|11|10|祭司就把耶和華殿裏所藏 大衛 王的槍和盾牌交給百夫長。
2KGS|11|11|護衛兵手中各拿兵器，在祭壇和殿那裏，從殿南到殿北，站在王的四圍。
2KGS|11|12|耶何耶大 領 約阿施 出來，給他戴上冠冕，把律法書交給他，膏他作王；眾人都鼓掌說：「願王萬歲！」
2KGS|11|13|亞她利雅 聽見護衛兵和百姓的聲音，就進耶和華的殿，到百姓那裏。
2KGS|11|14|她觀看，看哪，王照儀式站在柱旁，百夫長和號手在王旁邊，國中的眾百姓歡樂吹號。 亞她利雅 就撕裂衣服，喊著說：「反了！反了！」
2KGS|11|15|耶何耶大 祭司吩咐管軍兵的百夫長，對他們說：「把她從行列之間趕出去，凡跟隨她的必用刀殺死！」因為祭司說：「不可在耶和華殿裏殺她。」
2KGS|11|16|他們就下手拿住她；她進入通往王宮的 馬門 ，就在那裏被殺。
2KGS|11|17|耶何耶大 使王和百姓與耶和華立約，作耶和華的子民，又使王與百姓立約。
2KGS|11|18|於是國中的眾百姓都到 巴力 廟去，拆毀了廟，徹底打碎祭壇和偶像，又在壇前把 巴力 的祭司 瑪坦 殺了。 耶何耶大 祭司派官員看守耶和華的殿，
2KGS|11|19|又率領百夫長， 迦利 人和護衛兵，以及國中的眾百姓，請王從耶和華的殿下來，由護衛兵的門進入王宮，他就坐上王位。
2KGS|11|20|國中的眾百姓都歡樂，合城也都平靜。他們已將 亞她利雅 在王宮那裏用刀殺了。
2KGS|11|21|約阿施 登基的時候年方七歲。
2KGS|12|1|耶戶 第七年， 約阿施 登基，在 耶路撒冷 作王四十年。他母親名叫 西比亞 ，是 別是巴 人。
2KGS|12|2|約阿施 在 耶何耶大 祭司教導他的一切日子，行耶和華眼中看為正的事。
2KGS|12|3|只是丘壇還沒有廢去，百姓仍在丘壇獻祭燒香。
2KGS|12|4|約阿施 對眾祭司說：「凡獻到耶和華殿分別為聖的銀子，無論是人的贖價，各人生命的贖價， 或自願獻給耶和華殿的銀子，
2KGS|12|5|祭司可以各自從認識的人收取，用來修理殿的破壞之處，就是在那裏發現的一切破壞之處。」
2KGS|12|6|然而，到了 約阿施 王第二十三年，祭司仍未修理殿的破壞之處。
2KGS|12|7|所以 約阿施 王召了 耶何耶大 祭司和眾祭司來，對他們說：「你們怎麼不修理殿的破壞之處呢？現在，不要再從認識的人收銀子了，但要為了殿的破壞之處，把銀子交出來。」
2KGS|12|8|眾祭司答應不再收百姓的銀子，也不再修理殿的破壞之處。
2KGS|12|9|耶何耶大 祭司取了一個櫃子，在櫃蓋上鑽了一個洞，放在祭壇旁，在進耶和華殿的右邊；守門的祭司將獻到耶和華殿的一切銀子投在櫃裏。
2KGS|12|10|他們見櫃裏的銀子多了，就叫王的書記和大祭司上來，將耶和華殿裏所得的銀子數點了，包起來。
2KGS|12|11|他們把秤好了的銀子交在管理耶和華殿督工的手裏，督工就支付給木匠和建造耶和華殿的工人，
2KGS|12|12|瓦匠和石匠，又買木料和鑿成的石頭，用來修理耶和華殿的破壞之處，以及其他修理殿的各項費用。
2KGS|12|13|但這些獻到耶和華殿的銀子，並沒有用來造耶和華殿裏的銀杯、鉗子、盤子、號筒和其他的金銀器皿。
2KGS|12|14|他們把這銀子交給工人，用來整修耶和華的殿。
2KGS|12|15|他們不用跟這些經手接受銀子去支付工人的人算賬，因為這些人辦事誠實。
2KGS|12|16|贖愆祭和贖罪祭的銀子沒有獻到耶和華的殿裏，都歸給祭司。
2KGS|12|17|那時， 亞蘭 王 哈薛 上來攻打 迦特 ，攻取了它。 哈薛 就定意上來攻打 耶路撒冷 。
2KGS|12|18|猶大 王 約阿施 將他祖先 猶大 王 約沙法 、 約蘭 、 亞哈謝 所分別為聖的物和自己所分別為聖的物，以及耶和華殿與王宮府庫裏所有的金子都送給 亞蘭 王 哈薛 ； 哈薛 就不上 耶路撒冷 來了。
2KGS|12|19|約阿施 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|12|20|約阿施 的臣僕起來背叛，在下到 悉拉 路上的 米羅 宮那裏把他殺了。
2KGS|12|21|殺他的臣僕就是 示米押 的兒子 約撒拔 和 朔默 的兒子 約薩拔 。他與祖先同葬在 大衛城 ，他兒子 亞瑪謝 接續他作王。
2KGS|13|1|亞哈謝 的兒子 猶大 王 約阿施 第二十三年， 耶戶 的兒子 約哈斯 在 撒瑪利亞 登基作 以色列 王十七年。
2KGS|13|2|約哈斯 行耶和華眼中看為惡的事，效法 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪，總不離開。
2KGS|13|3|於是，耶和華的怒氣向 以色列 發作，將他們屢次交在 亞蘭 王 哈薛 和他兒子 便‧哈達 的手裏。
2KGS|13|4|約哈斯 懇求耶和華，耶和華就應允他，因為耶和華看見 以色列 所受的欺壓，因 亞蘭 王欺壓他們。
2KGS|13|5|耶和華賜給 以色列 一位拯救者，使他們脫離 亞蘭 人的手，於是 以色列 人仍舊安居在自己的帳棚裏。
2KGS|13|6|然而他們不離開 耶羅波安 家使 以色列 陷入罪裏的那罪，仍行在罪中，並且在 撒瑪利亞 留下 亞舍拉 。
2KGS|13|7|亞蘭 王滅絕 約哈斯 的軍隊，踐踏他們如禾場上的塵沙，只給 約哈斯 留下五十騎兵，十輛戰車，一萬步兵。
2KGS|13|8|約哈斯 其餘的事，凡他所做的和他英勇的事蹟，不都寫在《以色列諸王記》上嗎？
2KGS|13|9|約哈斯 與他祖先同睡，葬在 撒瑪利亞 ，他兒子 約阿施 接續他作王。
2KGS|13|10|猶大 王 約阿施 第三十七年， 約哈斯 的兒子 約阿施 在 撒瑪利亞 登基作 以色列 王十六年。
2KGS|13|11|他行耶和華眼中看為惡的事，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的一切罪，仍行在罪中。
2KGS|13|12|約阿施 其餘的事，凡他所做的和他與 猶大 王 亞瑪謝 交戰的英勇事蹟，不都寫在《以色列諸王記》上嗎？
2KGS|13|13|約阿施 與他祖先同睡， 耶羅波安 坐上他的王位。 約阿施 與 以色列 諸王一同葬在 撒瑪利亞 。
2KGS|13|14|以利沙 得了致命的病， 以色列 王 約阿施 下來看他，伏在他臉上哭泣，說：「我父啊！我父啊！ 以色列 的戰車和騎兵啊！」
2KGS|13|15|以利沙 對他說：「把弓箭拿來。」王就拿了弓箭來。
2KGS|13|16|以利沙 對 以色列 王說：「你用手開弓。」王就用手開弓。 以利沙 按手在王的手上，
2KGS|13|17|說：「打開朝東的窗戶。」他就打開。 以利沙 說：「射箭！」他就射箭。 以利沙 說：「這是耶和華得勝的箭，是戰勝 亞蘭 人的箭，因為你必在 亞弗 攻打 亞蘭 人，直到滅盡他們。」
2KGS|13|18|以利沙 又說：「拿幾枝箭來。」他就拿了來。 以利沙 對 以色列 王說：「打地吧！」他打了三次，就停止了。
2KGS|13|19|神人向他發怒，說：「你應當擊打五六次，就能攻打 亞蘭 人直到滅盡；現在你只能打敗 亞蘭 人三次。」
2KGS|13|20|以利沙 死了，人把他埋葬了。新的一年， 摩押 人成群結隊入侵境內。
2KGS|13|21|有人正在埋葬死人，看哪，他們看見一群人來，就把死人拋在 以利沙 的墳墓裏，逃跑了。死人一碰到 以利沙 的骸骨，就活過來，用腳站了起來。
2KGS|13|22|約哈斯 在位年間， 亞蘭 王 哈薛 屢次欺壓 以色列 。
2KGS|13|23|耶和華卻因與 亞伯拉罕 、 以撒 、 雅各 所立的約，仍施恩給 以色列 人，憐憫他們，眷顧他們，不肯滅盡他們，直到現在 仍不趕逐他們離開自己面前。
2KGS|13|24|亞蘭 王 哈薛 死了，他兒子 便‧哈達 接續他作王。
2KGS|13|25|從前 哈薛 和 約阿施 的父親 約哈斯 交戰，攻取了些城鎮，現在 約哈斯 的兒子 約阿施 三次打敗 哈薛 的兒子 便‧哈達 ，從他手中收回了 以色列 的城鎮。
2KGS|14|1|約哈斯 的兒子 以色列 王 約阿施 第二年， 猶大 王 約阿施 的兒子 亞瑪謝 登基。
2KGS|14|2|他登基的時候年二十五歲，在 耶路撒冷 作王二十九年。他母親名叫 約耶但 ，是 耶路撒冷 人。
2KGS|14|3|亞瑪謝 行耶和華眼中看為正的事，但不如他祖先 大衛 。他效法他父親 約阿施 一切所行的。
2KGS|14|4|只是丘壇還沒有廢去，百姓仍在丘壇獻祭燒香。
2KGS|14|5|王國在他手裏鞏固的時候，他就把殺他父王的臣僕殺了，
2KGS|14|6|卻沒有處死殺王兇手的兒子，正如 摩西 律法書上耶和華所吩咐的說：「不可因子殺父，也不可因父殺子，各人要為自己的罪而死。」
2KGS|14|7|亞瑪謝 在 鹽谷 殺了一萬 以東 人，又在戰役中攻取了 西拉 ，稱它為 約帖 ，直到今日。
2KGS|14|8|那時， 亞瑪謝 派使者到 耶戶 的孫子， 約哈斯 的兒子 以色列 王 約阿施 那裏，說：「來，讓我們面對面較量吧！」
2KGS|14|9|以色列 王 約阿施 派人去見 猶大 王 亞瑪謝 ，說：「 黎巴嫩 的蒺藜派人去見 黎巴嫩 的香柏樹，說：『將你的女兒嫁給我的兒子。』但有一隻野獸經過 黎巴嫩 ，把蒺藜踐踏了。
2KGS|14|10|你果然打敗了 以東 ，就心高氣傲。你以此為榮，就待在自己家裏算了吧，為何要惹禍，使自己和 猶大 一同敗亡呢？」
2KGS|14|11|亞瑪謝 卻不肯聽從。於是 以色列 王 約阿施 上來，在 猶大 的 伯‧示麥 與 猶大 王 亞瑪謝 面對面較量。
2KGS|14|12|猶大 敗在 以色列 面前，他們逃跑，各人逃回自己的帳棚去了。
2KGS|14|13|以色列 王 約阿施 在 伯‧示麥 擒住 亞哈謝 的孫子， 約阿施 的兒子 猶大 王 亞瑪謝 ，就來到 耶路撒冷 ，拆毀 耶路撒冷 的城牆，從 以法蓮門 直到 角門 共四百肘。
2KGS|14|14|他又拿了耶和華殿裏與王宮府庫裏所有的金銀和器皿，並帶著人質，回 撒瑪利亞 去了。
2KGS|14|15|約阿施 其餘所做的事和他英勇的事蹟，以及他與 猶大 王 亞瑪謝 交戰的事，不都寫在《以色列諸王記》上嗎？
2KGS|14|16|約阿施 與他祖先同睡，與 以色列 諸王一同葬在 撒瑪利亞 ，他兒子 耶羅波安 接續他作王。
2KGS|14|17|約哈斯 的兒子 以色列 王 約阿施 死後， 猶大 王 約阿施 的兒子 亞瑪謝 又活了十五年。
2KGS|14|18|亞瑪謝 其餘的事，不都寫在《猶大列王記》上嗎？
2KGS|14|19|耶路撒冷 有人背叛 亞瑪謝 ， 亞瑪謝 逃往 拉吉 ；他們卻派人追到 拉吉 ，在那裏殺了他。
2KGS|14|20|有人用馬將他馱回，葬在 耶路撒冷 ，與他祖先一同葬在 大衛城 。
2KGS|14|21|猶大 眾百姓立 亞撒利雅 接續他父親 亞瑪謝 作王，那時他年十六歲。
2KGS|14|22|亞瑪謝 王與他祖先同睡之後， 亞撒利雅 收復 以拉他 回歸 猶大 ，又重新整修。
2KGS|14|23|約阿施 的兒子 猶大 王 亞瑪謝 第十五年， 以色列 王 約阿施 的兒子 耶羅波安 在 撒瑪利亞 登基，作王四十一年。
2KGS|14|24|他行耶和華眼中看為惡的事，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的一切罪。
2KGS|14|25|他收回 以色列 邊界之地，從 哈馬口 直到 亞拉巴海 ，正如耶和華－ 以色列 的上帝藉他僕人 迦特．希弗 人 亞米太 的兒子 約拿 先知所說的。
2KGS|14|26|因耶和華看見 以色列 非常艱苦的困境；沒有奴役的，沒有自由的，也沒有人來幫助 以色列 。
2KGS|14|27|耶和華並沒有說要將 以色列 的名從天下塗抹，卻要藉 約阿施 的兒子 耶羅波安 拯救他們。
2KGS|14|28|耶羅波安 其餘的事，凡他所做的和他英勇的事蹟，他怎樣作戰，怎樣收復 大馬士革 和先前屬 猶大 的 哈馬 回歸 以色列 ，不都寫在《以色列諸王記》上嗎？
2KGS|14|29|耶羅波安 與他祖先 以色列 諸王同睡，他兒子 撒迦利雅 接續他作王。
2KGS|15|1|以色列 王 耶羅波安 第二十七年， 猶大 王 亞瑪謝 的兒子 亞撒利雅 登基。
2KGS|15|2|他登基的時候年十六歲，在 耶路撒冷 作王五十二年。他母親名叫 耶可利雅 ，是 耶路撒冷 人。
2KGS|15|3|亞撒利雅 行耶和華眼中看為正的事，效法他父親 亞瑪謝 一切所行的。
2KGS|15|4|只是丘壇還沒有廢去，百姓仍在丘壇獻祭燒香。
2KGS|15|5|耶和華降災於王，使他長了痲瘋，直到死的那日。他住在隔離的行宮裏，他兒子 約坦 管理王的家，治理這地的百姓。
2KGS|15|6|亞撒利雅 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|15|7|亞撒利雅 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 約坦 接續他作王。
2KGS|15|8|猶大 王 亞撒利雅 第三十八年， 耶羅波安 的兒子 撒迦利雅 登基，在 撒瑪利亞 作 以色列 王六個月。
2KGS|15|9|他行耶和華眼中看為惡的事，效法他祖先所行的，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪。
2KGS|15|10|雅比 的兒子 沙龍 背叛他，在百姓面前 擊殺他，篡了他的位。
2KGS|15|11|撒迦利雅 其餘的事，看哪，都寫在《以色列諸王記》上。
2KGS|15|12|這就是耶和華應許 耶戶 的話：「你的子孫必坐 以色列 的王位，直到第四代。」這事果然發生了。
2KGS|15|13|猶大 王 烏西雅 第三十九年， 雅比 的兒子 沙龍 登基，在 撒瑪利亞 作王一個月。
2KGS|15|14|迦底 的兒子 米拿現 從 得撒 上 撒瑪利亞 ，殺了 雅比 的兒子 沙龍 ，篡了他的位。
2KGS|15|15|沙龍 其餘的事和他陰謀背叛的事，看哪，都寫在《以色列諸王記》上。
2KGS|15|16|那時， 米拿現 從 得撒 起擊殺 提斐薩 和城中所有的人，以及它周圍的地區，因為他們沒有給他開城門。他擊殺他們，剖開其中所有的孕婦。
2KGS|15|17|猶大 王 亞撒利雅 第三十九年， 迦底 的兒子 米拿現 登基，在 撒瑪利亞 作 以色列 王十年。
2KGS|15|18|他行耶和華眼中看為惡的事，終生不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪。
2KGS|15|19|亞述 王 普勒 來攻擊這地， 米拿現 給他一千他連得銀子，為了請 普勒 幫助他鞏固他所掌握的國度。
2KGS|15|20|米拿現 向 以色列 所有的富豪索取銀子，要他們各出五十舍客勒，交給 亞述 王。於是 亞述 王回去了，不在境內停留。
2KGS|15|21|米拿現 其餘的事，凡他所做的，不都寫在《以色列諸王記》上嗎？
2KGS|15|22|米拿現 與他祖先同睡，他兒子 比加轄 接續他作王。
2KGS|15|23|猶大 王 亞撒利雅 第五十年， 米拿現 的兒子 比加轄 登基，在 撒瑪利亞 作 以色列 王二年。
2KGS|15|24|他行耶和華眼中看為惡的事，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪。
2KGS|15|25|比加轄 的將軍， 利瑪利 的兒子 比加 背叛他，在 撒瑪利亞 王宮的堡壘殺了他。 亞珥歌伯 和 亞利耶 並 基列 的五十人幫助 比加 ； 比加 擊殺他，篡了他的位。
2KGS|15|26|比加轄 其餘的事，凡他所做的，看哪，都寫在《以色列諸王記》上。
2KGS|15|27|猶大 王 亞撒利雅 第五十二年， 利瑪利 的兒子 比加 登基，在 撒瑪利亞 作 以色列 王二十年。
2KGS|15|28|他行耶和華眼中看為惡的事，不離開 尼八 的兒子 耶羅波安 使 以色列 陷入罪裏的那罪。
2KGS|15|29|在 以色列 王 比加 的日子， 亞述 王 提革拉‧毗列色 來奪取 以雲 、 亞伯‧伯‧瑪迦 、 亞挪 、 基低斯 、 夏瑣 、 基列 、 加利利 和 拿弗他利 全地，把這些地方的居民都擄到 亞述 去了。
2KGS|15|30|烏西雅 的兒子 約坦 第二十年， 以拉 的兒子 何細亞 背叛 利瑪利 的兒子 比加 ，擊殺他，篡了他的位。
2KGS|15|31|比加 其餘的事，凡他所做的，看哪，都寫在《以色列諸王記》上。
2KGS|15|32|利瑪利 的兒子 以色列 王 比加 第二年， 猶大 王 烏西雅 的兒子 約坦 登基。
2KGS|15|33|他登基的時候年二十五歲，在 耶路撒冷 作王十六年。他母親名叫 耶路沙 ，是 撒督 的女兒。
2KGS|15|34|約坦 行耶和華眼中看為正的事，效法他父親 烏西雅 一切所行的。
2KGS|15|35|只是丘壇還沒有廢去，百姓仍在丘壇獻祭燒香。 約坦 建了耶和華殿的 上門 。
2KGS|15|36|約坦 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|15|37|在那些日子，耶和華開始差 亞蘭 王 利汛 和 利瑪利 的兒子 比加 去攻擊 猶大 。
2KGS|15|38|約坦 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 亞哈斯 接續他作王。
2KGS|16|1|利瑪利 的兒子 比加 第十七年， 猶大 王 約坦 的兒子 亞哈斯 登基。
2KGS|16|2|他登基的時候年二十歲，在 耶路撒冷 作王十六年。他不像他祖先 大衛 行耶和華－他上帝眼中看為正的事，
2KGS|16|3|卻行 以色列 諸王的道，又照著耶和華從 以色列 人面前趕出的外邦人所行可憎的事，使他的兒子經火，
2KGS|16|4|並在丘壇上、山岡上、各青翠樹下獻祭燒香。
2KGS|16|5|那時， 亞蘭 王 利汛 和 利瑪利 的兒子 以色列 王 比加 上來攻打 耶路撒冷 ，圍困 亞哈斯 ，卻不能打勝。
2KGS|16|6|當時 亞蘭 王 利汛 收復 以拉他 回歸 亞蘭 ，把 猶大 人從 以拉他 趕出去。 以東 人來到 以拉他 ，住在那裏，直到今日。
2KGS|16|7|亞哈斯 派使者到 亞述 王 提革拉‧毗列色 那裏，說：「我是你的僕人，你的兒子。現在 亞蘭 王和 以色列 王攻擊我，求你上來，救我脫離他們的手。」
2KGS|16|8|亞哈斯 將耶和華殿裏和王宮府庫裏所有的金銀都送給 亞述 王為禮物。
2KGS|16|9|亞述 王答應了他，上去攻打 大馬士革 ，攻下了城，殺了 利汛 ，把居民擄到 吉珥 。
2KGS|16|10|亞哈斯 王到 大馬士革 迎接 亞述 王 提革拉‧毗列色 ，在 大馬士革 看見一座壇。 亞哈斯 王把壇的規模和樣式，以及作法的細節，送到 烏利亞 祭司那裏。
2KGS|16|11|烏利亞 祭司照著 亞哈斯 王從 大馬士革 所送來的一切，在 亞哈斯 王還未從 大馬士革 回來之前，築了一座壇。
2KGS|16|12|王從 大馬士革 回來，看見壇，走近壇前，在壇上獻祭。
2KGS|16|13|他燒燔祭和素祭，獻澆酒祭，將平安祭牲的血灑在壇上。
2KGS|16|14|他移動耶和華面前的銅壇，從殿的前面，新壇和耶和華殿的中間，搬到新壇的北邊。
2KGS|16|15|亞哈斯 王吩咐 烏利亞 祭司說：「早晨的燔祭、晚上的素祭，王的燔祭、素祭，國內眾百姓的燔祭、素祭、澆酒祭都要燒在大壇上。燔祭牲和其他祭牲的血全都要灑在這壇上。至於銅壇，我要作求問之用。」
2KGS|16|16|烏利亞 祭司就照著 亞哈斯 王所吩咐的一切做了。
2KGS|16|17|亞哈斯 王把盆座四面的嵌邊拆下來，把盆從座上挪下來，又將銅海從馱銅海的銅牛上搬下來，放在石板鋪的地上。
2KGS|16|18|他為了 亞述 王的緣故，在耶和華的殿裏移動 殿裏為安息日所蓋的遮棚 和王從外面進來的入口。
2KGS|16|19|亞哈斯 其餘所做的事，不都寫在《猶大列王記》上嗎？
2KGS|16|20|亞哈斯 與他祖先同睡， 與他祖先同葬在 大衛城 ，他兒子 希西家 接續他作王。
2KGS|17|1|猶大 王 亞哈斯 第十二年， 以拉 的兒子 何細亞 在 撒瑪利亞 登基作 以色列 王九年。
2KGS|17|2|他行耶和華眼中看為惡的事，只是不像在他以前的 以色列 諸王。
2KGS|17|3|亞述 王 撒縵以色 上來攻擊 何細亞 ， 何細亞 就服事他，向他進貢。
2KGS|17|4|何細亞 背叛，派使者到 埃及 王 梭 那裏 ，不照往年所行的向 亞述 王進貢。 亞述 王知道了，就逮捕他，把他囚在監裏。
2KGS|17|5|亞述 王上來攻擊 以色列 全地，上到 撒瑪利亞 ，圍困這城三年。
2KGS|17|6|何細亞 第九年， 亞述 王攻取了 撒瑪利亞 ，把 以色列 人擄到 亞述 ，安置在 哈臘 與 歌散 的 哈博河 邊，以及 瑪代 人的城鎮。
2KGS|17|7|這是因為 以色列 人得罪了那領他們出 埃及 地、脫離 埃及 王法老之手的耶和華－他們的上帝，去敬畏別神，
2KGS|17|8|隨從耶和華在 以色列 人面前所趕出外邦人的風俗和 以色列 諸王所立的規條。
2KGS|17|9|以色列 人暗中行不正的事，違背耶和華－他們的上帝，在他們所有的城鎮，從瞭望樓直到堅固城，建築丘壇；
2KGS|17|10|在各高岡上、各青翠樹下立柱像和 亞舍拉 ；
2KGS|17|11|在各丘壇上燒香，效法耶和華在他們面前趕出的外邦人所行的，又行惡事，惹耶和華發怒。
2KGS|17|12|他們事奉偶像，耶和華對他們說：「你們不可做這事。」
2KGS|17|13|耶和華藉眾先知、先見勸戒 以色列 和 猶大 說：「當離開你們的惡行，謹守我的誡命律例，遵行我吩咐你們祖先、藉我僕人眾先知所傳給你們的一切律法。」
2KGS|17|14|他們卻不聽從，竟硬著頸項，像他們祖先一樣，不信服耶和華－他們的上帝。
2KGS|17|15|他們厭棄他的律例，和他與他們列祖所立的約，以及他勸戒他們的話，去隨從虛無的神明 ，自己成為虛妄，效法周圍的列國，就是耶和華囑咐他們不可效法的。
2KGS|17|16|他們離棄耶和華－他們上帝的一切誡命，為自己鑄造了兩個牛犢的像，立了 亞舍拉 ，敬拜天上的萬象，事奉 巴力 ，
2KGS|17|17|使他們的兒女經火，占卜，行法術，出賣自己，行耶和華眼中看為惡的事，惹他發怒。
2KGS|17|18|所以耶和華向 以色列 大大發怒，從自己面前趕出他們，只剩下 猶大 一個支派。
2KGS|17|19|但是， 猶大 也不遵守耶和華－他們上帝的誡命，效法 以色列 所立的規條。
2KGS|17|20|耶和華就厭棄 以色列 所有的後裔，使他們受苦，把他們交在搶奪他們的人手中，直到他把他們從自己面前趕出去。
2KGS|17|21|當他使 以色列 從 大衛 家分離出來的時候，他們立 尼八 的兒子 耶羅波安 作王。 耶羅波安 引誘 以色列 不隨從耶和華，陷入大罪中。
2KGS|17|22|以色列 人行 耶羅波安 所犯的一切罪，總不離開，
2KGS|17|23|以致耶和華把他們從自己面前趕出去，正如他藉他僕人眾先知所說的。這樣， 以色列 人從自己的土地被擄到 亞述 ，直到今日。
2KGS|17|24|亞述 王從 巴比倫 、 古他 、 亞瓦 、 哈馬 和 西法瓦音 遷移人來，安置在 撒瑪利亞 的城鎮，代替 以色列 人；他們就佔據了 撒瑪利亞 ，住在城中。
2KGS|17|25|他們開始住在那裏的時候，不敬畏耶和華，所以耶和華叫獅子進入他們中間，咬死了一些人。
2KGS|17|26|有人對 亞述 王說：「你所遷移安置在 撒瑪利亞 城鎮的各國的人，他們不知道那地之上帝的規矩，所以他叫獅子進入他們中間。看哪，獅子咬死了他們，因為他們不知道那地之上帝的規矩。」
2KGS|17|27|亞述 王吩咐說：「當派一個從那裏擄來的祭司回去，叫他住在那裏，將那地之上帝的規矩指導他們。」
2KGS|17|28|於是有一個從 撒瑪利亞 擄去的祭司回來，住在 伯特利 ，教導他們怎樣敬畏耶和華。
2KGS|17|29|然而，各國的人在所住的城裏為自己製造神像，安置在 撒瑪利亞 人所建有丘壇的廟中。
2KGS|17|30|巴比倫 人造 疏割‧比訥 像； 古他 人造 匿甲 像； 哈馬 人造 亞示瑪 像；
2KGS|17|31|亞瓦 人造 匿哈 和 他珥他 像； 西法瓦音 人用火焚燒兒女，獻給 西法瓦音 的神明 亞得米勒 和 亞拿米勒 。
2KGS|17|32|他們懼怕耶和華，卻從他們中間立丘壇的祭司，在丘壇的廟中為他們獻祭。
2KGS|17|33|他們懼怕耶和華，但又事奉自己的神明，從何邦遷來，就隨從那裏的風俗，
2KGS|17|34|直到如今仍照先前的風俗去行。 他們不敬畏耶和華，不遵守耶和華吩咐 雅各 後裔的律例、典章、律法、誡命； 雅各 就是從前耶和華起名叫 以色列 的。
2KGS|17|35|耶和華曾與他們立約，吩咐他們說：「不可敬畏別神，不可跪拜事奉它們，也不可向它們獻祭。
2KGS|17|36|惟有那用大能和伸出來的膀臂領你們出 埃及 地的耶和華，你們當敬畏他，向他跪拜，向他獻祭。
2KGS|17|37|他給你們寫的律例、典章、律法、誡命，你們應當永遠謹守遵行。你們不可敬畏別神。
2KGS|17|38|你們不可忘記我與你們所立的約，也不可敬畏別神。
2KGS|17|39|只要敬畏耶和華－你們的上帝，他必救你們脫離一切仇敵的手。」
2KGS|17|40|他們卻不聽從，仍照先前的風俗去行。
2KGS|17|41|這樣，這些國家又懼怕耶和華，又事奉他們的偶像。他們子子孫孫也都照樣行，效法他們的祖宗，直到今日。
2KGS|18|1|以拉 的兒子 以色列 王 何細亞 第三年， 猶大 王 亞哈斯 的兒子 希西家 登基。
2KGS|18|2|他登基的時候年二十五歲，在 耶路撒冷 作王二十九年。他母親名叫 亞比 ，是 撒迦利雅 的女兒。
2KGS|18|3|希西家 行耶和華眼中看為正的事，效法他祖先 大衛 一切所行的。
2KGS|18|4|他廢去丘壇，毀壞柱像，砍下 亞舍拉 ，打碎 摩西 所造的銅蛇，因為到那時 以色列 人仍向銅蛇燒香。人叫銅蛇為 尼忽士但 。
2KGS|18|5|希西家 倚靠耶和華－ 以色列 的上帝，在他之前和在他之後的 猶大 列王中沒有一個像他一樣的。
2KGS|18|6|因為他緊緊跟隨耶和華，謹守耶和華所吩咐 摩西 的誡命，總不離開。
2KGS|18|7|耶和華與他同在，他無論往何處去盡都亨通。他背叛 亞述 王，不服事他。
2KGS|18|8|希西家 攻擊 非利士 人，直到 迦薩 ，以及所屬的領土，從瞭望樓到堅固城。
2KGS|18|9|希西家 王第四年，也就是 以拉 的兒子 以色列 王 何細亞 第七年， 亞述 王 撒縵以色 上來圍困 撒瑪利亞 。
2KGS|18|10|過了三年，他們攻取了城。 希西家 第六年， 以色列 王 何細亞 第九年， 撒瑪利亞 被攻取了。
2KGS|18|11|亞述 王把 以色列 人擄到 亞述 ，安置在 哈臘 與 歌散 的 哈博河 邊，以及 瑪代 人的城鎮。
2KGS|18|12|這是因為他們不聽從耶和華－他們的上帝的話，違背了他的約；他們既不聽從，也不遵行耶和華僕人 摩西 一切所吩咐的。
2KGS|18|13|希西家 王十四年， 亞述 王 西拿基立 上來攻擊 猶大 的一切堅固的城，將城攻取。
2KGS|18|14|猶大 王 希西家 派人到 拉吉 ， 亞述 王那裏，說：「我錯了，求你撤退離開我；凡你罰我的，我必承當。」於是 亞述 王罰 猶大 王 希西家 三百他連得銀子，三十他連得金子。
2KGS|18|15|希西家 把耶和華殿裏和王宮府庫裏所有的銀子都給了他。
2KGS|18|16|那時， 猶大 王 希西家 將耶和華殿門上的金子和他自己包在柱子上的金子都刮下來，給了 亞述 王。
2KGS|18|17|亞述 王從 拉吉 差遣元帥 、太監長 和將軍 率領大軍前往 耶路撒冷 ，到 希西家 王那裏去。他們上來，到 耶路撒冷 。他們上來之後，站在 上池 的水溝旁，在往漂布地的大路上。
2KGS|18|18|他們呼叫王， 希勒家 的兒子 以利亞敬 宮廷總管， 舍伯那 書記和 亞薩 的兒子 約亞 史官就出來見他們。
2KGS|18|19|將軍對他們說：「你們去告訴 希西家 ，大王 亞述 王如此說：『你倚靠甚麼，讓你如此自信滿滿？
2KGS|18|20|你說，你有打仗的計謀和能力，我看不過是空話。你到底倚靠誰，竟敢背叛我呢？
2KGS|18|21|現在，看哪，你自己所倚靠的 埃及 是那斷裂的葦杖，人若倚靠這杖，它就刺進他的手，穿透它。 埃及 王法老向所有倚靠他的人都是這樣。
2KGS|18|22|你們若對我說：我們倚靠耶和華－我們的上帝， 希西家 豈不是將上帝的丘壇和祭壇廢去，並且吩咐 猶大 和 耶路撒冷 的人說：你們當在 耶路撒冷 這壇前敬拜嗎？
2KGS|18|23|現在你與我主 亞述 王打賭，我給你兩千匹馬，看你能否派得出騎士來騎牠們。
2KGS|18|24|若不然，怎能使我主臣僕中最小的一個軍官轉臉而逃呢？你難道要倚靠 埃及 的戰車和騎兵嗎？
2KGS|18|25|現在我上來攻擊毀滅這地方，豈不是出於耶和華嗎？耶和華吩咐我說，你上去攻擊這地，毀滅它吧！』」
2KGS|18|26|希勒家 的兒子 以利亞敬 ， 舍伯那 和 約亞 對將軍說：「求你用 亞蘭 話對僕人說，因為我們聽得懂；不要用 猶大 話對我們說，免得傳到城牆上百姓的耳中。」
2KGS|18|27|將軍對他們說：「我主差遣我來，豈是單對你和你的主人說這些話嗎？不也是對這些坐在城牆上、要與你們一同吃自己糞、喝自己尿的人說的嗎？」
2KGS|18|28|於是 亞述 將軍站著，用 猶大 話大聲喊著說：「你們當聽大王 亞述 王的話，
2KGS|18|29|王如此說：『你們不要被 希西家 欺哄了，因他不能救你們脫離我的手。
2KGS|18|30|不要聽憑 希西家 說服你們倚靠耶和華，他說，耶和華必要拯救我們，這城必不交在 亞述 王的手中。』
2KGS|18|31|你們不要聽 希西家 的話！因 亞述 王如此說：『你們要與我講和，出來投降我，各人就可以吃自己葡萄樹和無花果樹的果子，喝自己井裏的水，
2KGS|18|32|等我來領你們到一個地方，與你們本地一樣，就是有五穀和新酒之地，有糧食和葡萄園之地，有橄欖樹和蜂蜜之地，好使你們存活，不至於死。不要聽 希西家 的話，因為他誤導你們說：耶和華必拯救我們。
2KGS|18|33|列國的神明有哪一個曾救它本國脫離 亞述 王的手呢？
2KGS|18|34|哈馬 、 亞珥拔 的神明在哪裏呢？ 西法瓦音 、 希拿 、 以瓦 的神明在哪裏呢？ 它們曾救 撒瑪利亞 脫離我的手嗎？
2KGS|18|35|這些國的神明有誰曾救自己的國脫離我的手呢？難道耶和華能救 耶路撒冷 脫離我的手嗎？』」
2KGS|18|36|百姓靜默不言，一句不答，因為 希西家 王曾吩咐說：「不要回答他。」
2KGS|18|37|當下， 希勒家 的兒子 以利亞敬 宮廷總管、 舍伯那 書記和 亞薩 的兒子 約亞 史官，都撕裂衣服，來到 希西家 那裏，將 亞述 將軍的話告訴他。
2KGS|19|1|希西家 王聽見了，就撕裂衣服，披上麻布，進了耶和華的殿。
2KGS|19|2|他差遣 以利亞敬 宮廷總管和 舍伯那 書記，並祭司中年長的，都披上麻布，到 亞摩斯 的兒子 以賽亞 先知那裏去。
2KGS|19|3|他們對他說：「 希西家 如此說：『今日是急難、懲罰、凌辱的日子，就如嬰孩快要出生，卻沒有力氣生產。
2KGS|19|4|或許耶和華－你的上帝聽見 亞述 將軍一切的話，就是他主人 亞述 王差他來辱罵永生上帝的話，耶和華－你的上帝就斥責所聽見的這些話。求你為倖存的餘民揚聲禱告。』」
2KGS|19|5|希西家 王的臣僕來到 以賽亞 那裏的時候，
2KGS|19|6|以賽亞 對他們說：「要對你們的主人這樣說，耶和華如此說：『你聽見 亞述 王的僕人褻瀆我的話，不要懼怕。
2KGS|19|7|看哪，我必驚動他的心 ，他要聽見風聲就歸回本地，在那裏我必使他倒在刀下。』」
2KGS|19|8|亞述 將軍聽見 亞述 王已拔營離開 拉吉 ，就啟程返回，正遇見 亞述 王去攻打 立拿 。
2KGS|19|9|亞述 王聽見有人談論 古實 王 特哈加 說：「看哪，他出來要與你爭戰。」於是 亞述 王又差使者去見 希西家 ，說：
2KGS|19|10|「你們要對 猶大 王 希西家 如此說：『不要聽你所倚靠的上帝欺哄你說： 耶路撒冷 必不交在 亞述 王的手中。
2KGS|19|11|看哪，你總聽說 亞述 諸王向列國所行的是盡行滅絕，難道你能倖免嗎？
2KGS|19|12|我祖先所毀滅的，就是 歌散 、 哈蘭 、 利色 和 提‧拉撒 的 伊甸 人；這些國的神明何曾拯救他們呢？
2KGS|19|13|哈馬 的王， 亞珥拔 的王， 西法瓦音城 的王， 希拿 和 以瓦 的王，都在哪裏呢？』」
2KGS|19|14|希西家 從使者手裏接過書信，讀完了，就上耶和華的殿，在耶和華面前展開書信。
2KGS|19|15|希西家 向耶和華禱告說：「坐在基路伯之上耶和華－ 以色列 的上帝啊，你，惟有你是地上萬國的上帝，你創造了天和地。
2KGS|19|16|耶和華啊，求你側耳而聽；耶和華啊，求你睜眼而看，聽 西拿基立 差遣使者辱罵永生上帝的話。
2KGS|19|17|耶和華啊， 亞述 諸王果然使列國和列國之地變為荒蕪，
2KGS|19|18|將列國的神像扔在火裏，因為它們不是上帝，是人手所造的，是木頭、石頭，所以被滅絕了。
2KGS|19|19|耶和華－我們的上帝啊，現在求你救我們脫離 亞述 王的手，使地上萬國都知道惟獨你－耶和華是上帝！」
2KGS|19|20|亞摩斯 的兒子 以賽亞 差人去見 希西家 ，說：「耶和華－ 以色列 的上帝如此說：你因 亞述 王 西拿基立 的事向我祈求，我已聽見了。
2KGS|19|21|耶和華論他這樣說： 『少女 錫安 藐視你，嘲笑你； 耶路撒冷 向你搖頭。
2KGS|19|22|『你辱罵誰，褻瀆誰， 揚起聲來，高舉眼目攻擊誰呢？ 你攻擊的是 以色列 的聖者。
2KGS|19|23|你藉你的使者辱罵主說： 我率領許多戰車登上高山， 到 黎巴嫩 的頂端； 我要砍伐其中高大的香柏樹 和上好的松樹； 我必進到極遙遠的住所， 進入最茂盛的森林裏。
2KGS|19|24|我已經在外邦挖井喝水； 我必用腳掌踏乾 埃及 一切的河流。
2KGS|19|25|『你豈沒有聽見 我早先所定、古時所立、現今實現的事嗎？ 就是讓你去毀壞堅固的城鎮，使它們變為廢墟；
2KGS|19|26|城裏的居民力量微小， 他們驚惶羞愧； 像野草，像青菜， 如房頂上的草， 又如未長成而枯乾的禾稼。
2KGS|19|27|『你坐下，你出去，你進來， 你向我發烈怒，我都知道。
2KGS|19|28|因你向我發烈怒， 你的狂傲上達我耳中， 我要用鉤子鉤住你的鼻子， 將嚼環放在你口裏， 使你從原路轉回去。』
2KGS|19|29|「這是給你的預兆：你們今年要吃野生的，明年也要吃自長的；後年，你們就要耕種收割，栽葡萄園，吃其中的果子。
2KGS|19|30|猶大 家所逃脫剩餘的，仍要往下扎根，向上結果。
2KGS|19|31|必有剩餘的民從 耶路撒冷 而出，有逃脫的人從 錫安山 而來。萬軍之耶和華的熱心必成就這事。
2KGS|19|32|「所以耶和華論 亞述 王如此說：他必不得來到這城，也不在這裏射箭，不得拿盾牌到城前，也不建土堆攻城。
2KGS|19|33|他從哪條路來，必從那條路回去，必不得來到這城。這是耶和華說的。
2KGS|19|34|因我為自己的緣故，又為我僕人 大衛 的緣故，必保護拯救這城。」
2KGS|19|35|當夜，耶和華的使者出去，在 亞述 營中殺了十八萬五千人。清早有人起來，看哪，都是死屍。
2KGS|19|36|亞述 王 西拿基立 就拔營回去，住在 尼尼微 。
2KGS|19|37|一日，他在他的神明 尼斯洛 廟裏叩拜，他兒子 亞得米勒 和 沙利色 用刀殺了他，然後逃到 亞拉臘 地；他兒子 以撒．哈頓 接續他作王。
2KGS|20|1|那些日子， 希西家 病得要死， 亞摩斯 的兒子 以賽亞 先知來見他，對他說：「耶和華如此說：『你當留遺囑給你的家，因為你必死，不能活了。』」
2KGS|20|2|希西家 轉臉朝牆，向耶和華禱告說：
2KGS|20|3|「耶和華啊，求你記念我在你面前怎樣存完全的心，按誠實行事，又做你眼中看為善的事。」 希西家 就痛哭。
2KGS|20|4|以賽亞 出來，還沒有離開中院，耶和華的話就臨到他，說：
2KGS|20|5|「你回去告訴我百姓的君王 希西家 說：耶和華－你祖先 大衛 的上帝如此說：『我聽見了你的禱告，看見了你的眼淚。看哪，我必醫治你；到第三日，你必上到耶和華的殿。
2KGS|20|6|我必加添你十五年的壽數，並且我要救你和這城脫離 亞述 王的手。我為自己和我僕人 大衛 的緣故，必保護這城。』」
2KGS|20|7|以賽亞 說：「取一塊無花果餅來。」人就取了來，貼在瘡上，王就痊癒了。
2KGS|20|8|希西家 對 以賽亞 說：「耶和華必醫治我，到第三日我能上耶和華的殿，有甚麼預兆呢？」
2KGS|20|9|以賽亞 說：「耶和華必成就他所說的這話。這是耶和華給你的預兆：你要日影向前進十度呢？或是要往後退十度呢？」
2KGS|20|10|希西家 說：「日影向前進十度容易；不，讓日影往後退十度吧。」
2KGS|20|11|以賽亞 先知求告耶和華，耶和華就使 亞哈斯 日晷上照下來的日影，往後退了十度。
2KGS|20|12|那時， 巴拉但 的兒子， 巴比倫 王 米羅達‧巴拉但 聽見 希西家 生病了，就送書信和禮物給他。
2KGS|20|13|希西家 聽使者的話 ，就將自己一切寶庫裏的金子、銀子、香料、貴重的膏油和他軍械庫裏的兵器，以及他所有的財寶，都給他們看；在他家中和全國之內， 希西家 沒有一樣東西不給他們看的。
2KGS|20|14|於是 以賽亞 先知到 希西家 王那裏去，對他說：「這些人說了些甚麼？他們從哪裏來見你？」 希西家 說：「他們從遠方的 巴比倫 來。」
2KGS|20|15|以賽亞 說：「他們在你家裏看見了甚麼？」 希西家 說：「凡我家中所有的，他們都看見了；我財寶中沒有一樣東西不給他們看的。」
2KGS|20|16|以賽亞 對 希西家 說：「你要聽耶和華的話：
2KGS|20|17|耶和華說：『看哪，日子將到，凡你家裏所有的，並你祖先積蓄到如今的一切，都要被擄到 巴比倫 去，不留下一樣；
2KGS|20|18|從你本身所生的孩子，其中必有被擄到 巴比倫 王宮當太監的。』」
2KGS|20|19|希西家 對 以賽亞 說：「你所說耶和華的話甚好。」因為他想：「在我有生之年豈不是有太平和安穩嗎？」
2KGS|20|20|希西家 其餘的事和他一切英勇的事蹟，他怎樣造池、挖溝、引水入城，不都寫在《猶大列王記》上嗎？
2KGS|20|21|希西家 與他祖先同睡，他兒子 瑪拿西 接續他作王。
2KGS|21|1|瑪拿西 登基的時候年十二歲，在 耶路撒冷 作王五十五年。他母親名叫 協西巴 。
2KGS|21|2|瑪拿西 行耶和華眼中看為惡的事，效法耶和華在 以色列 人面前趕出的列國那些可憎的事。
2KGS|21|3|他重新建築他父親 希西家 所毀壞的丘壇，又為 巴力 築壇，造 亞舍拉 ，效法 以色列 王 亞哈 所行的，敬拜天上的萬象，事奉它們。
2KGS|21|4|他在耶和華殿中築壇，耶和華曾指著這殿說：「我必立我的名在 耶路撒冷 。」
2KGS|21|5|他在耶和華殿的兩個院子為天上的萬象築壇，
2KGS|21|6|並使他的兒子經火，又觀星象，行法術，求問招魂的和行巫術的，多行耶和華眼中看為惡的事，惹他發怒。
2KGS|21|7|他又把自己所造的 亞舍拉 雕像立在殿內，耶和華曾對 大衛 和他兒子 所羅門 說：「我在 以色列 眾支派中所選擇的 耶路撒冷 和這殿，必立我的名，直到永遠。
2KGS|21|8|只要 以色列 人謹守遵行我一切所吩咐的和我僕人 摩西 所吩咐的一切律法，我就不再使他們的腳挪移，離開我所賜給他們列祖之土地。」
2KGS|21|9|他們卻不聽從，並且 瑪拿西 引誘他們行惡，比耶和華在 以色列 人面前所滅的列國更嚴重。
2KGS|21|10|耶和華藉他僕人眾先知說：
2KGS|21|11|「因 猶大 王 瑪拿西 行這些可憎的惡事，比先前 亞摩利 人所行的一切更壞，使 猶大 人拜偶像，陷入罪裏，
2KGS|21|12|所以耶和華－ 以色列 的上帝如此說：看哪，我必降禍於 耶路撒冷 和 猶大 ，凡聽見的人都必雙耳齊鳴。
2KGS|21|13|我必用量 撒瑪利亞 的準繩和 亞哈 家的鉛垂線拉在 耶路撒冷 之上；我必擦拭 耶路撒冷 ，如人擦盤子，把盤子翻過來。
2KGS|21|14|我必撇棄我產業中的餘民，把他們交在仇敵手中，使他們成為所有仇敵的擄物和掠物，
2KGS|21|15|因為自從他們的祖先出 埃及 的那日直到今日，他們常行我眼中看為惡的事，惹我發怒。」
2KGS|21|16|瑪拿西 行耶和華眼中看為惡的事，使 猶大 陷入罪裏，又流許多無辜人的血，直到這血充滿了 耶路撒冷 ，從這邊到那邊。
2KGS|21|17|瑪拿西 其餘的事，凡他所做的和他所犯的罪，不都寫在《猶大列王記》上嗎？
2KGS|21|18|瑪拿西 與他祖先同睡，葬在自己王宮的園子， 烏撒 園裏，他兒子 亞們 接續他作王。
2KGS|21|19|亞們 登基的時候年二十二歲，在 耶路撒冷 作王二年。他母親名叫 米舒利密 ，是 約提巴 人 哈魯斯 的女兒。
2KGS|21|20|亞們 行耶和華眼中看為惡的事，效法他父親 瑪拿西 所行的。
2KGS|21|21|他行他父親一切所行的道，事奉他父親所事奉的偶像，敬拜它們，
2KGS|21|22|離棄耶和華－他列祖的上帝，不遵行耶和華的道。
2KGS|21|23|亞們 的臣僕背叛他，在宮裏殺了王。
2KGS|21|24|但這地的百姓殺了所有背叛 亞們 王的人；這地的百姓立他兒子 約西亞 接續他作王。
2KGS|21|25|亞們 其餘所做的事，不都寫在《猶大列王記》上嗎？
2KGS|21|26|亞們 葬在 烏撒 園內自己的墳墓裏，他兒子 約西亞 接續他作王。
2KGS|22|1|約西亞 登基的時候年八歲，在 耶路撒冷 作王三十一年。他母親名叫 耶底大 ，是 波斯加 人 亞大雅 的女兒。
2KGS|22|2|約西亞 行耶和華眼中看為正的事，行他祖先 大衛 一切所行的道，不偏左右。
2KGS|22|3|約西亞 王十八年，王派 米書蘭 的孫子， 亞薩利雅 的兒子 沙番 書記上耶和華殿去，說：
2KGS|22|4|「你上到 希勒家 大祭司那裏，請他把奉獻到耶和華殿的銀子，就是門口的守衛從百姓中收來的銀子，結算清楚，
2KGS|22|5|交在管理耶和華殿督工的手裏，由他們支付給在耶和華殿裏做工的人，好修理殿的破壞之處，
2KGS|22|6|就是木匠、工人和瓦匠，又買木料和鑿成的石頭，來整修殿宇。
2KGS|22|7|但他們不用跟這些經手接受銀子的人算帳，因為這些人辦事誠實。」
2KGS|22|8|希勒家 大祭司對 沙番 書記說：「我在耶和華殿裏發現了律法書。」 希勒家 把書遞給 沙番 ， 沙番 就讀了。
2KGS|22|9|沙番 書記到王那裏，把這事回覆王說：「你的僕人已把殿裏所發現的銀子倒出來，交在管理耶和華殿督工的手裏了。」
2KGS|22|10|沙番 書記又向王報告說：「 希勒家 祭司遞給我一卷書。」 沙番 就在王面前朗讀那書。
2KGS|22|11|王聽見律法書上的話，就撕裂衣服。
2KGS|22|12|王吩咐 希勒家 祭司與 沙番 的兒子 亞希甘 、 米該亞 的兒子 亞革波 、 沙番 書記和王的臣僕 亞撒雅 ，說：
2KGS|22|13|「你們去，以所發現這書上的話，為我、為百姓、為全 猶大 求問耶和華；因為我們祖先沒有聽從這書上的話，沒有遵照一切所寫有關我們的 去行，耶和華就向我們大發烈怒。」
2KGS|22|14|於是， 希勒家 祭司和 亞希甘 、 亞革波 、 沙番 、 亞撒雅 都去見 戶勒大 女先知，她是掌管禮服的 沙龍 的妻子； 沙龍 是 哈珥哈斯 的孫子， 特瓦 的兒子。 戶勒大 住在 耶路撒冷 第二區。他們向她請教。
2KGS|22|15|她對他們說：「耶和華－ 以色列 的上帝如此說：『你們可以回覆那派你們來見我的人說，
2KGS|22|16|耶和華如此說：看哪，我必照著 猶大 王所讀那書上的一切話，降禍於這地方和其上的居民。
2KGS|22|17|因為他們離棄我，向別神燒香，用他們手所做的一切惹我發怒，所以我的憤怒必向這地方發作，總不止息。』
2KGS|22|18|然而，派你們來求問耶和華的 猶大 王，你們要這樣回覆他：『耶和華－ 以色列 的上帝如此說：至於你所聽見的話，
2KGS|22|19|就是聽見我指著這地方和其上的居民說，要使這地方變為荒蕪、百姓受詛咒的話，你的心就軟化，在耶和華面前謙卑下來，撕裂衣服，向我哭泣，因此我應允你。這是耶和華說的。
2KGS|22|20|因此，看哪，我必使你歸到你祖先那裏，平安地進入墳墓；我要降於這地方的一切災禍，你不會親眼看見。』」他們就去把這話回覆王。
2KGS|23|1|王派人召集 猶大 和 耶路撒冷 的眾長老來。
2KGS|23|2|王和 猶大 眾人、 耶路撒冷 的居民、祭司、先知，以及所有的百姓，無論大小，都一同上到耶和華的殿去；王把耶和華殿裏所發現的約書上一切的話讀給他們聽。
2KGS|23|3|王站在柱子旁邊，在耶和華面前立約，要盡心盡性跟從耶和華，遵守他的誡命、法度、律例，實行這書上所寫這約的話。全體百姓都願遵守所立的約。
2KGS|23|4|王吩咐 希勒家 大祭司和副祭司，以及把守殿門的，把那些為 巴力 和 亞舍拉 ，以及天上萬象所造的器皿，都從耶和華殿裏搬出來，在 耶路撒冷 外 汲淪 的田間燒了，把灰拿到 伯特利 去。
2KGS|23|5|從前 猶大 列王所立拜偶像的祭司，在 猶大 城鎮的丘壇和 耶路撒冷 周圍燒香，現在王都廢去，他們是向 巴力 和日、月、行星，以及天上萬象燒香的人。
2KGS|23|6|他把 亞舍拉 從耶和華殿裏搬到 耶路撒冷 外的 汲淪溪 ，在 汲淪溪 邊焚燒，打碎成灰，把灰撒在平民的墳上。
2KGS|23|7|他又拆毀耶和華殿裏男的廟妓的屋子，就是婦女在那裏為 亞舍拉 編織衣服的屋子。
2KGS|23|8|他從 猶大 的城鎮將眾祭司帶來，從 迦巴 直到 別是巴 ，玷污祭司燒香的丘壇。他又拆毀城門旁的丘壇，這丘壇是在 約書亞 市長的城門前，在人進城門的左邊。
2KGS|23|9|只是丘壇的祭司不登 耶路撒冷 耶和華的壇，僅在他們弟兄中間吃無酵餅。
2KGS|23|10|他又玷污 欣嫩子谷 的 陀斐特 ，不許人在那裏使兒女經火獻給 摩洛 。
2KGS|23|11|他把在耶和華殿門旁、靠近 拿單‧米勒 官員走廊的屋子， 猶大 列王獻給太陽的馬廢去，且用火焚燒獻給太陽的戰車。
2KGS|23|12|猶大 列王在 亞哈斯 樓房頂上所築的壇和 瑪拿西 在耶和華殿兩院中所築的壇，王都拆毀，從那裏移走 ，把灰倒在 汲淪溪 中。
2KGS|23|13|從前 以色列 王 所羅門 在 耶路撒冷 東邊、 邪僻山 南邊為 西頓 人可憎的 亞斯她錄 、 摩押 人可憎的 基抹 、 亞捫 人可憎的 米勒公 所築的丘壇，王都玷污了，
2KGS|23|14|又打碎柱像，砍下 亞舍拉 ，用人的骨頭填滿那地方。
2KGS|23|15|此外，在 伯特利 丘壇的壇，就是 尼八 的兒子 耶羅波安 所築、使 以色列 人陷入罪裏的，他也把這壇和丘壇都拆毀了，又焚燒丘壇 ，打碎成灰，並焚燒了 亞舍拉 。
2KGS|23|16|約西亞 轉頭，看見山上的墳墓，就派人取出墳墓裏的骸骨，燒在壇上，玷污了壇，正如從前 耶羅波安 在節期中站在壇旁時，耶和華藉神人所宣告的話。 約西亞 轉頭看見了宣告這些話的神人的墳墓。
2KGS|23|17|他說：「我看見的這碑是甚麼呢？」那城裏的人對他說：「這是神人的墳墓，他從 猶大 來，宣告了王向 伯特利 的壇所做的這些事。」
2KGS|23|18|約西亞 說：「讓他安息吧！不要挪移他的骸骨。」他們就保存了他的骸骨和從 撒瑪利亞 來的那先知的骸骨。
2KGS|23|19|從前 以色列 諸王在 撒瑪利亞 的城鎮所建一切惹動怒氣的丘壇的廟， 約西亞 也都廢去了，正如他在 伯特利 所做的。
2KGS|23|20|他又把在那裏所有丘壇的祭司都殺在壇上，並在壇上燒人的骨頭。於是他回 耶路撒冷 去了。
2KGS|23|21|王吩咐眾百姓說：「你們當照這約書上所寫的，向耶和華－你們的上帝守逾越節。」
2KGS|23|22|自從士師治理 以色列 ，到 以色列 諸王、 猶大 列王在位的一切日子，從來沒有守過這樣的逾越節，
2KGS|23|23|只有在 約西亞 王十八年，才在 耶路撒冷 向耶和華守這逾越節。
2KGS|23|24|此外，在 猶大 地和 耶路撒冷 所見那些招魂的、行巫術的，家中的神像和偶像，以及一切可憎之物， 約西亞 盡都除掉，實行了 希勒家 祭司在耶和華殿裏所發現的律法書上所寫的話。
2KGS|23|25|在 約西亞 以前，沒有王像他盡心、盡性、盡力地歸向耶和華，遵行 摩西 的一切律法；在他以後，也沒有興起一個王像他。
2KGS|23|26|然而，耶和華向 猶大 所發猛烈的怒氣仍不止息，因為 瑪拿西 種種的惡事激怒了他。
2KGS|23|27|耶和華說：「我也必將 猶大 從我面前趕出，如同趕出 以色列 一樣。我必撇棄我從前所選擇的這城 耶路撒冷 和我所說我的名必留在那裏的殿。」
2KGS|23|28|約西亞 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|23|29|約西亞 的日子， 埃及 王法老 尼哥 上到 幼發拉底河 ，到 亞述 王那裏； 約西亞 王去迎擊他。 埃及 王在 米吉多 看見 約西亞 ，就殺了他。
2KGS|23|30|他的臣僕用車把他的屍體從 米吉多 送到 耶路撒冷 ，葬在他自己的墳墓裏。這地的百姓選 約西亞 的兒子 約哈斯 ，膏立他，接續他父親作王。
2KGS|23|31|約哈斯 登基的時候年二十三歲，在 耶路撒冷 作王三個月。他母親名叫 哈慕她 ，是 立拿 人 耶利米 的女兒。
2KGS|23|32|約哈斯 行耶和華眼中看為惡的事，效法他祖先一切所行的。
2KGS|23|33|法老 尼哥 把 約哈斯 監禁在 哈馬 地的 利比拉 ，不許他在 耶路撒冷 作王 ，又罰這地一百他連得銀子，一他連得金子。
2KGS|23|34|法老 尼哥 立 約西亞 的兒子 以利亞敬 接續他父親 約西亞 作王，給他改名叫 約雅敬 ，卻把 約哈斯 帶到 埃及 ，他就死在那裏。
2KGS|23|35|約雅敬 進貢金銀給法老，照著法老的指示在這地徵收銀子，向這地的百姓按各人的能力索取金銀，要送給法老 尼哥 。
2KGS|23|36|約雅敬 登基的時候年二十五歲，在 耶路撒冷 作王十一年。他母親名叫 西布大 ，是 魯瑪 人 毗大雅 的女兒。
2KGS|23|37|約雅敬 行耶和華眼中看為惡的事，效法他祖先一切所行的。
2KGS|24|1|約雅敬 的日子， 巴比倫 王 尼布甲尼撒 上來； 約雅敬 服事他三年，以後又背叛他。
2KGS|24|2|耶和華派 迦勒底 、 亞蘭 、 摩押 和 亞捫 人的軍隊來攻擊 約雅敬 ；耶和華派他們來攻擊 猶大 ，要毀滅它，正如耶和華藉他僕人眾先知所說的話。
2KGS|24|3|這事臨到 猶大 ，誠然是出於耶和華的命令 ，要把 猶大 從自己面前趕出去，是因 瑪拿西 所犯的一切罪，
2KGS|24|4|又因他流無辜人的血，使無辜人的血充滿 耶路撒冷 ；耶和華不願赦免。
2KGS|24|5|約雅敬 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
2KGS|24|6|約雅敬 與他祖先同睡，他兒子 約雅斤 接續他作王。
2KGS|24|7|埃及 王不再從他的國出征，因為 巴比倫 王把 埃及 王所管之地，從 埃及 溪谷直到 幼發拉底河 都奪去了。
2KGS|24|8|約雅斤 登基的時候年十八歲，在 耶路撒冷 作王三個月。他母親名叫 尼護施她 ，是 耶路撒冷 人 以利拿單 的女兒。
2KGS|24|9|約雅斤 行耶和華眼中看為惡的事，效法他父親一切所行的。
2KGS|24|10|那時， 巴比倫 王 尼布甲尼撒 的軍兵上到 耶路撒冷 ，城被圍困。
2KGS|24|11|當他的軍兵圍困城的時候， 巴比倫 王 尼布甲尼撒 親自來到 耶路撒冷 。
2KGS|24|12|猶大 王 約雅斤 和他母親、臣僕、王子、官員一同出來，向 巴比倫 王投降。 巴比倫 王俘擄了他，那時是 巴比倫 王第八年。
2KGS|24|13|巴比倫 王把耶和華殿裏和王宮裏一切的寶物從那裏拿走，又把 以色列 王 所羅門 所造耶和華殿裏一切的金器都毀壞了，正如耶和華所說的。
2KGS|24|14|他把全 耶路撒冷 眾領袖和所有大能的勇士，共一萬人，連同所有的木匠和鐵匠都擄了去，只留下這地最貧窮的百姓。
2KGS|24|15|他把 約雅斤 和他的母親、后妃、官員，以及這地的貴族，都從 耶路撒冷 擄到 巴比倫 去了，
2KGS|24|16|又把所有的勇士七千人，木匠和鐵匠一千人，全是能上陣的勇士，都擄到 巴比倫 去了。
2KGS|24|17|巴比倫 王立 約雅斤 的叔父 瑪探雅 取代他作王，給 瑪探雅 改名叫 西底家 。
2KGS|24|18|西底家 登基的時候年二十一歲，在 耶路撒冷 作王十一年。他母親名叫 哈慕她 ，是 立拿 人 耶利米 的女兒。
2KGS|24|19|西底家 行耶和華眼中看為惡的事，正如 約雅敬 一切所行的。
2KGS|24|20|因此，耶和華向 耶路撒冷 和 猶大 發怒，以致把他們從自己面前趕出去。 西底家 背叛 巴比倫 王。
2KGS|25|1|西底家 作王第九年十月初十， 巴比倫 王 尼布甲尼撒 率領全軍前來攻擊 耶路撒冷 ，對城安營，四圍築堡壘攻城。
2KGS|25|2|城被圍困，直到 西底家 王十一年。
2KGS|25|3|四月初九，城裏的饑荒非常嚴重，當地的百姓都沒有糧食。
2KGS|25|4|城被攻破，士兵全都在夜間從靠近王的花園、兩城牆中間的門逃跑。 迦勒底 人正在四圍攻城，王就往 亞拉巴 逃去。
2KGS|25|5|迦勒底 的軍隊追趕王，在 耶利哥 的平原追上他；他的全軍都離開他潰散了。
2KGS|25|6|迦勒底 人就拿住王，帶他到 利比拉 的 巴比倫 王那裏；他們就判他的罪。
2KGS|25|7|他們在 西底家 眼前殺了他的兒女，挖了 西底家 的眼睛，用銅鏈鎖著他，帶到 巴比倫 去。
2KGS|25|8|巴比倫 王 尼布甲尼撒 十九年五月初七， 巴比倫 王的臣僕 尼布撒拉旦 護衛長進入 耶路撒冷 ，
2KGS|25|9|他焚燒了耶和華的殿、王宮和 耶路撒冷 一切的房屋；用火焚燒所有大戶人家的房屋。
2KGS|25|10|跟從護衛長的 迦勒底 全軍拆毀了 耶路撒冷 四圍的城牆。
2KGS|25|11|那時 尼布撒拉旦 護衛長將城裏剩下的百姓和那些投降 巴比倫 王的人，以及其餘的眾人，都擄去了。
2KGS|25|12|但護衛長留下一些當地最窮的人，叫他們修整葡萄園，耕種田地。
2KGS|25|13|耶和華殿的銅柱並殿內的盆座和銅海， 迦勒底 人都打碎了，把那些銅運到 巴比倫 去。
2KGS|25|14|他們又帶走鍋、鏟子、鉗子、勺子和供奉用的一切銅器；
2KGS|25|15|火盆和碗，無論金的銀的，護衛長都帶走了；
2KGS|25|16|還有 所羅門 為耶和華殿所造的兩根柱子、一個銅海和盆座，這一切器皿的銅多得無法可秤。
2KGS|25|17|這一根柱子高十八肘，柱上有銅頂，銅頂高三肘；銅頂的周圍有網子和石榴，也都是銅的。第二根柱子與此相同，也有網子。
2KGS|25|18|護衛長拿住 西萊雅 大祭司、 西番亞 副祭司和門口的三個守衛，
2KGS|25|19|又從城中拿住一個管理士兵的官 ，並在城裏所找到王面前的五個親信，和召募當地百姓之將軍的書記官，以及在城中找到的六十個當地百姓。
2KGS|25|20|尼布撒拉旦 護衛長把這些人帶到 利比拉 的 巴比倫 王那裏。
2KGS|25|21|巴比倫 王擊殺他們，在 哈馬 地的 利比拉 把他們處死。這樣， 猶大 人就被擄去離開本地。
2KGS|25|22|至於 猶大 地剩下的百姓，就是 巴比倫 王 尼布甲尼撒 所留下的， 巴比倫 王立了 沙番 的孫子， 亞希甘 的兒子 基大利 作他們的省長。
2KGS|25|23|所有的軍官和屬他們的人聽見 巴比倫 王立了 基大利 作省長， 尼探雅 的兒子 以實瑪利 、 加利亞 的兒子 約哈難 、 尼陀法 人 單戶蔑 的兒子 西萊雅 、 瑪迦 人的兒子 雅撒尼亞 ，和屬他們的人，都來到 米斯巴 的 基大利 那裏。
2KGS|25|24|基大利 向他們和屬他們的人起誓說：「你們不必懼怕 迦勒底 臣僕，只管住在這地，服事 巴比倫 王，就可以得福。」
2KGS|25|25|七月中，王室後裔 以利沙瑪 的孫子， 尼探雅 的兒子 以實瑪利 帶著十個人來，擊殺了 基大利 和同他在 米斯巴 的 猶大 人與 迦勒底 人，把他們殺死。
2KGS|25|26|於是眾人，無論大小，連同軍官，因為懼怕 迦勒底 人，都起身逃到 埃及 去了。
2KGS|25|27|巴比倫 王 以未‧米羅達 作王的元年，就是 猶大 王 約雅斤 被擄後三十七年，十二月二十七日，他使 猶大 王 約雅斤 抬起頭來，提他出監，
2KGS|25|28|對他說好話，使他的位高過與他一同被擄在 巴比倫 眾王的位；
2KGS|25|29|又給他脫了囚服，使他終身常在 巴比倫 王面前吃飯。
2KGS|25|30|王賜給他日常需用的食物，每日一份，終身都是這樣。
