JUDG|1|1|約書亞 死後， 以色列 人求問耶和華說：「我們中間誰當首先上去攻打 迦南 人，與他們爭戰呢？」
JUDG|1|2|耶和華說：「 猶大 要先上去。看哪，我已將那地交在他手中。」
JUDG|1|3|猶大 對他哥哥 西緬 說：「請你同我上到我抽籤所得之地，與 迦南 人爭戰；我也同你去你抽籤所得之地。」於是 西緬 與他同去。
JUDG|1|4|猶大 就上去，耶和華把 迦南 人和 比利洗 人交在他們手中。他們在 比色 擊殺了一萬人。
JUDG|1|5|他們在 比色 遇見 亞多尼‧比色 ，與他爭戰，擊敗了 迦南 人和 比利洗 人。
JUDG|1|6|亞多尼‧比色 逃跑，他們追趕他，捉住他，砍斷他大拇指和大腳趾。
JUDG|1|7|亞多尼‧比色 說：「從前有七十個王，大拇指和大腳趾都被我砍斷，在我桌子底下拾取零碎食物。現在上帝照著我所做的報應我了。」他們把 亞多尼‧比色 帶到 耶路撒冷 ，他就死在那裏。
JUDG|1|8|猶大 人攻打 耶路撒冷 ，奪取了它，用刀殺城內的人，並且放火燒城。
JUDG|1|9|後來 猶大 人下去，與住山區、 尼革夫 和低地的 迦南 人爭戰。
JUDG|1|10|猶大 去攻打住 希伯崙 的 迦南 人，殺了 示篩 、 亞希幔 、 撻買 。 希伯崙 從前名叫 基列‧亞巴 。
JUDG|1|11|猶大 從那裏去攻擊 底壁 的居民。 底壁 從前名叫 基列‧西弗 。
JUDG|1|12|迦勒 說：「誰能攻打 基列‧西弗 ，奪取那城，我就把我女兒 押撒 嫁給他。」
JUDG|1|13|迦勒 的弟弟 基納斯 的兒子 俄陀聶 奪取了那城， 迦勒 就把女兒 押撒 嫁給他。
JUDG|1|14|押撒 來的時候，催促丈夫 向她父親要一塊田。 押撒 一下驢， 迦勒 就對她說：「你要甚麼？」
JUDG|1|15|她對 迦勒 說：「求你賜我福分；你既然把 尼革夫 給了我，求你也給我水泉。」 迦勒 就把上泉和下泉都賜給她。
JUDG|1|16|摩西 的岳父是 基尼 人，他的子孫與 猶大 人一起上到棕樹城，往 亞拉得 以南的 猶大 曠野 去，住在百姓當中 。
JUDG|1|17|猶大 和他哥哥 西緬 同去，擊殺了住 洗法 的 迦南 人，將城徹底毀滅。因此，那城名叫 何珥瑪 。
JUDG|1|18|猶大 攻取了 迦薩 和所屬的領土， 亞實基倫 和所屬的領土， 以革倫 和所屬的領土。
JUDG|1|19|耶和華與 猶大 同在， 猶大 取得了山區，卻不能趕出平原的居民，因為他們有鐵的戰車。
JUDG|1|20|以色列 人照 摩西 所說的，把 希伯崙 給了 迦勒 。 迦勒 從那裏趕出 亞衲 的三支後裔。
JUDG|1|21|至於住 耶路撒冷 的 耶布斯 人， 便雅憫 人沒有把他們趕出。於是， 耶布斯 人與 便雅憫 人同住在 耶路撒冷 ，直到今日。
JUDG|1|22|約瑟 家也上到 伯特利 去，耶和華與他們同在。
JUDG|1|23|約瑟 家去窺探 伯特利 ，那城起先名叫 路斯 。
JUDG|1|24|探子看見一個人從城裏出來，就對他說：「請你把進城的路指示我們，我們會厚待你。」
JUDG|1|25|那人把進城的路指示他們。他們就用刀擊殺了城中的居民，卻放走那人和他的全家。
JUDG|1|26|那人往 赫 人之地去，建造了一座城，起名叫 路斯 。那城到如今還叫這名。
JUDG|1|27|瑪拿西 沒有趕出 伯˙善 和所屬鄉鎮 的居民， 他納 和所屬鄉鎮的居民， 多珥 和所屬鄉鎮的居民， 以伯蓮 和所屬鄉鎮的居民， 米吉多 和所屬鄉鎮的居民； 迦南 人仍堅持住在這地。
JUDG|1|28|以色列 強盛的時候，就叫 迦南 人做苦工，沒有把他們全然趕走。
JUDG|1|29|以法蓮 沒有趕出住 基色 的 迦南 人。於是 迦南 人仍住在 基色 ，在 以法蓮 中間。
JUDG|1|30|西布倫 沒有趕出 基倫 的居民和 拿哈拉 的居民。於是 迦南 人仍住在 西布倫 中間，成了服勞役的人。
JUDG|1|31|亞設 沒有趕出 亞柯 的居民和 西頓 的居民，以及 亞黑拉 、 亞革悉 、 黑巴 、 亞弗革 和 利合 的居民。
JUDG|1|32|亞設 人因為沒有趕出那地的居民 迦南 人，就住在他們中間。
JUDG|1|33|拿弗他利 沒有趕出 伯˙示麥 和 伯˙亞納 的居民。於是 拿弗他利 就住在那地的居民 迦南 人中，而 伯˙示麥 和 伯˙亞納 的居民卻成了為他們服勞役的人。
JUDG|1|34|亞摩利 人強逼 但 人住在山區，不准他們下到平原。
JUDG|1|35|亞摩利 人仍堅持住在 希烈山 、 亞雅崙 和 沙賓 ；然而 約瑟 家權勢強盛的時候，他們成為服勞役的人。
JUDG|1|36|亞摩利 人 的地界是從 亞克拉濱 斜坡，從 西拉 延伸而上。
JUDG|2|1|耶和華的使者從 吉甲 上到 波金 ，說：「我領你們從 埃及 上來，帶你們到我向你們列祖起誓應許之地。我曾說：『我永不廢棄我與你們的約。
JUDG|2|2|你們不可與這地的居民立約，要拆毀他們的祭壇。』你們竟沒有聽從我的話。你們為何這樣做呢！
JUDG|2|3|因此我說：『我必不將他們從你們面前趕出。他們必作你們肋下的荊棘 ，他們的神明必成為你們的圈套。』」
JUDG|2|4|耶和華的使者向 以色列 眾人說這些話的時候，百姓放聲大哭。
JUDG|2|5|於是他們給那地方起名叫 波金 ，並在那裏向耶和華獻祭。
JUDG|2|6|約書亞 解散百姓， 以色列 人回到自己的地業，佔各自的地。
JUDG|2|7|約書亞 在世的日子和他死了以後，那些見過耶和華為 以色列 所做一切大事的長老還在世的時候，百姓都事奉耶和華。
JUDG|2|8|耶和華的僕人， 嫩 的兒子 約書亞 死了，那時他一百一十歲。
JUDG|2|9|以色列 人把他葬在他自己地業的境內， 以法蓮 山區的 亭拿‧希烈 ，在 迦實山 的北邊。
JUDG|2|10|那世代的人也都歸到自己的列祖。後來興起的另一世代不認識耶和華，也不知道他為 以色列 所做的事。
JUDG|2|11|以色列 人行耶和華眼中看為惡的事，去事奉諸 巴力 。
JUDG|2|12|他們離棄領他們出 埃及 地的耶和華－他們列祖的上帝，去隨從別神，就是四圍列國的神明，向它們叩拜，惹耶和華發怒。
JUDG|2|13|他們離棄了耶和華，去事奉 巴力 和 亞斯她錄 。
JUDG|2|14|耶和華的怒氣向 以色列 發作，把他們交在搶奪他們的人手中，又把他們交給四圍仇敵的手中 ，以致他們在仇敵面前再也不能站立得住。
JUDG|2|15|他們無論往何處去，耶和華的手都以災禍攻擊他們，正如耶和華所說的，又如耶和華向他們所起的誓；他們就極其困苦。
JUDG|2|16|耶和華興起士師，士師就拯救他們脫離搶奪他們之人的手。
JUDG|2|17|然而，他們卻不聽從士師，竟隨從別神而行淫，向它們叩拜。他們列祖所行的道，所聽從耶和華的命令，他們都速速偏離了，並不照樣遵行。
JUDG|2|18|耶和華為他們興起士師，耶和華與士師同在。士師在世的一切日子，耶和華拯救他們脫離仇敵的手。耶和華因他們受欺壓迫害所發出的哀聲，就憐憫他們。
JUDG|2|19|但士師一死，他們又轉去行惡，比他們祖宗更壞，去隨從別神，事奉叩拜它們，總不放棄他們的惡習和頑梗的行為。
JUDG|2|20|於是耶和華的怒氣向 以色列 發作，說：「因為這國違背我吩咐他們列祖當守的約，不聽從我的話，
JUDG|2|21|約書亞 死的時候所剩下的各國，我必不再從他們面前趕出任何一個，
JUDG|2|22|為要藉此考驗 以色列 是否肯謹守遵行耶和華的道，像他們列祖一樣地謹守。」
JUDG|2|23|耶和華留下那些國家，不將他們速速趕出，也不把他們交在 約書亞 的手中。
JUDG|3|1|耶和華留下這些國家，為要考驗所有未曾經歷 迦南 任何戰役的 以色列 人，
JUDG|3|2|只是為了要 以色列 人的後代認識戰爭，教導他們，尤其那些未曾認識這些事的人。
JUDG|3|3|留下的有 非利士 的五個領袖，所有的 迦南 人， 西頓 人，以及從 巴力‧黑門山 到 哈馬口 ，住 黎巴嫩山 的 希未 人。
JUDG|3|4|他們是為了要考驗 以色列 ，好知道他們是否肯聽從耶和華藉 摩西 吩咐他們列祖的命令。
JUDG|3|5|以色列 人住在 迦南 人、 赫 人、 亞摩利 人、 比利洗 人、 希未 人、 耶布斯 人中間，
JUDG|3|6|娶他們的女兒，將自己的女兒嫁給他們的兒子，並事奉他們的神明。
JUDG|3|7|以色列 人行耶和華眼中看為惡的事，忘記耶和華－他們的上帝，去事奉諸 巴力 和 亞舍拉 ，
JUDG|3|8|所以耶和華的怒氣向 以色列 發作，把他們交給 美索不達米亞 王 古珊‧利薩田 的手中。 以色列 人服事 古珊‧利薩田 八年。
JUDG|3|9|以色列 人呼求耶和華，耶和華就為 以色列 人興起一位拯救者來救他們，就是 迦勒 的弟弟 基納斯 的兒子 俄陀聶 。
JUDG|3|10|耶和華的靈降在他身上，他就作了 以色列 的士師。他出去爭戰，耶和華將 亞蘭 王 古珊‧利薩田 交在他手中，他的手戰勝了 古珊‧利薩田 。
JUDG|3|11|於是這地太平四十年。 基納斯 的兒子 俄陀聶 死了。
JUDG|3|12|以色列 人又行耶和華眼中看為惡的事。耶和華使 摩押 王 伊磯倫 強大，攻擊 以色列 ，因為他們行耶和華眼中看為惡的事。
JUDG|3|13|伊磯倫 召集 亞捫 人和 亞瑪力 人到他那裏，他就去攻打 以色列 ，佔據了棕樹城。
JUDG|3|14|於是 以色列 人服事 摩押 王 伊磯倫 十八年。
JUDG|3|15|以色列 人呼求耶和華，耶和華就為他們興起一位拯救者， 便雅憫 人 基拉 的兒子 以笏 ，他是個慣用左手的人 。 以色列 人託他送禮物給 摩押 王 伊磯倫 。
JUDG|3|16|以笏 打造了一把兩刃的劍，長一短肘 ，綁在右腿上衣服裏面。
JUDG|3|17|他把禮物獻給 摩押 王 伊磯倫 。 伊磯倫 是個很肥胖的人。
JUDG|3|18|以笏 獻完禮物的時候，就把抬禮物的人送走。
JUDG|3|19|但他自己卻從靠近 吉甲 的雕像那裏轉回來，說：「王啊，我有一件機密的事要奏告你。」王說：「迴避吧！」於是所有侍立在他左右的人都退去了。
JUDG|3|20|以笏 來到王那裏，那時他獨自一人坐在陰涼的頂樓。 以笏 說：「我有上帝的話向你報告。」王就從座位上站起來。
JUDG|3|21|以笏 伸出左手，從右腿上拔出劍來，刺入王的肚腹。
JUDG|3|22|劍柄連同劍刃都刺進去了，肥肉夾住了劍刃。他沒有把劍從王的肚腹拔出來，糞便就流出來了 。
JUDG|3|23|以笏 出到門廊，把王關在樓門裏面，就上了鎖。
JUDG|3|24|以笏 出來之後，王的僕人就來了。他們觀看，看哪，樓門鎖住，就說：「他必是在陰涼的房間裏大解。」
JUDG|3|25|他們等得不耐煩，看哪，樓門仍然不開，就拿鑰匙打開樓門，看哪，他們的主人已經倒在地上死了。
JUDG|3|26|他們耽延的時候， 以笏 就逃跑了。他經過雕像那裏，逃到 西伊拉 。
JUDG|3|27|他到了那裏，就在 以法蓮 山區吹角。 以色列 人跟隨他從山區下來，他在他們前面引路，
JUDG|3|28|對他們說：「緊跟著我！因為耶和華已經把你們的仇敵 摩押 交在你們手中。」於是他們跟著他下去，佔據了 摩押 對面 約旦河 的渡口，不准一人過去。
JUDG|3|29|那時，他們擊殺了約一萬 摩押 人，都是強壯的勇士，連一個也沒有逃脫。
JUDG|3|30|那日， 摩押 在 以色列 手下制伏了。於是這地太平八十年。
JUDG|3|31|以笏 之後，有 亞拿 的兒子 珊迦 ，他用趕牛的棍子打死六百 非利士 人。他也拯救了 以色列 。
JUDG|4|1|以笏 死後， 以色列 人又行耶和華眼中看為惡的事。
JUDG|4|2|耶和華把他們交給在 夏瑣 作王的 迦南 王 耶賓 手中；他的將軍是 西西拉 ，住在 夏羅設‧哈歌印 。
JUDG|4|3|以色列 人呼求耶和華，因為 耶賓 王有鐵的戰車九百輛，並且殘酷欺壓 以色列 人二十年。
JUDG|4|4|有一位女先知 底波拉 ，是 拉比多 的妻子，當時作 以色列 的士師。
JUDG|4|5|她住在 以法蓮 山區 拉瑪 和 伯特利 的中間，在 底波拉 的棕樹下。 以色列 人都上到她那裏去聽審判。
JUDG|4|6|她派人從 拿弗他利 的 基低斯 把 亞比挪菴 的兒子 巴拉 召來，對他說：「耶和華－ 以色列 的上帝吩咐你：『你要率領一萬 拿弗他利 人和 西布倫 人上 他泊山 去。
JUDG|4|7|我必使 耶賓 的將軍 西西拉 率領他的戰車和全軍往 基順河 ，到你那裏去，我必把他交在你手中。』」
JUDG|4|8|巴拉 對她說：「你若同我去，我就去；你若不同我去，我就不去。」
JUDG|4|9|底波拉 說：「我一定會與你同去，然而你在所行的路上必得不著榮耀，因為耶和華要把 西西拉 交給一個婦人的手裏。」於是 底波拉 起來，與 巴拉 一同往 基低斯 去了。
JUDG|4|10|巴拉 召集 西布倫 人和 拿弗他利 人到 基低斯 ，跟他上去的有一萬人。 底波拉 也同他上去。
JUDG|4|11|摩西 岳父 何巴 的後裔， 基尼 人 希百 離開了 基尼 族，到靠近 基低斯 的 撒拿音 橡樹旁支搭帳棚。
JUDG|4|12|有人告訴 西西拉 ：「 亞比挪菴 的兒子 巴拉 已經上了 他泊山 。」
JUDG|4|13|西西拉 就召集所有的鐵戰車九百輛和隨從的全軍，從 夏羅設‧哈歌印 出來，到了 基順河 。
JUDG|4|14|底波拉 對 巴拉 說：「起來，今日就是耶和華把 西西拉 交在你手中的日子。耶和華豈不在你前面行嗎?」於是 巴拉 下了 他泊山 ，跟隨他的有一萬人。
JUDG|4|15|耶和華使 西西拉 和他一切的戰車，以及全軍潰亂，在 巴拉 面前倒在刀下。 西西拉 下了車，徒步逃跑。
JUDG|4|16|巴拉 追趕戰車、軍隊，直到 夏羅設‧哈歌印 。 西西拉 的全軍都倒在刀下，一個也沒有留下。
JUDG|4|17|只有 西西拉 徒步逃跑到 基尼 人 希百 之妻 雅億 的帳棚，因為 夏瑣 王 耶賓 與 基尼 人的 希百 家和平共處。
JUDG|4|18|雅億 出來迎接 西西拉 ，對他說：「請我主進來，進到我這裏來，不要怕。」 西西拉 就進了她的帳棚， 雅億 用被子將他蓋住。
JUDG|4|19|西西拉 對 雅億 說：「我渴了，求你給我一點水喝。」 雅億 就打開裝奶的皮袋，給他喝，再把他蓋住。
JUDG|4|20|西西拉 對 雅億 說：「請你站在帳棚門口，若有人來問你說：『有人在這裏嗎？』你就說：『沒有。』」
JUDG|4|21|西西拉 疲乏沉睡了。 希百 的妻 雅億 取了帳棚的橛子，手拿著錘子，靜悄悄地到他那裏，將橛子從他的太陽穴釘進去，直釘到地裏。 西西拉 就死了。
JUDG|4|22|看哪， 巴拉 追趕 西西拉 ， 雅億 出來迎接他，對他說：「來，我給你看你要找的人。」他就進入帳棚，看哪， 西西拉 已經倒在地上死了，橛子還在他的太陽穴中。
JUDG|4|23|那日，上帝在 以色列 人面前制伏了 迦南 王 耶賓 。
JUDG|4|24|從此， 以色列 人的手對 迦南 王 耶賓 越來越強硬，直到將 迦南 王 耶賓 剪除。
JUDG|5|1|那日， 底波拉 和 亞比挪菴 的兒子 巴拉 唱歌，說：
JUDG|5|2|「 以色列 有領袖率領 ， 百姓甘心犧牲自己， 你們當稱頌耶和華！
JUDG|5|3|「君王啊，要聽！王子啊，要側耳！ 我要，我要向耶和華歌唱； 我要歌頌耶和華－ 以色列 的上帝。
JUDG|5|4|「耶和華啊，你從 西珥 出來， 從 以東 田野向前行， 地震動 天滴下， 雲也滴下雨水。
JUDG|5|5|眾山在耶和華面前搖動， 西奈山 在耶和華－ 以色列 上帝面前也搖動。
JUDG|5|6|「在 亞拿 之子 珊迦 的時候， 在 雅億 的日子， 大道無人行走， 過路人繞道而行。
JUDG|5|7|以色列 農村荒蕪， 空無一人， 直到我 底波拉 興起， 興起作 以色列 之母！
JUDG|5|8|以色列 人選擇新的諸神， 戰爭就臨到城門。 以色列 四萬人中， 看得見盾牌槍矛嗎？
JUDG|5|9|我心嚮往 以色列 的領袖， 他們在民中甘心犧牲自己。 你們應當稱頌耶和華！
JUDG|5|10|「騎淺色母驢的、 坐繡花毯子的、 行走在路上的， 你們都當思想！
JUDG|5|11|打水的聲音勝過弓箭的響聲， 那裏，人要述說耶和華公義的作為， 他對 以色列 鄉民公義的作為。 「那時，耶和華的子民下到城門。
JUDG|5|12|「 底波拉 啊，興起！興起！ 當興起，興起，唱歌！ 巴拉 啊，你當興起！ 亞比挪菴 的兒子啊，當俘擄你的俘虜！
JUDG|5|13|那時，貴族中的倖存者前進， 耶和華的百姓為我前進攻擊勇士。
JUDG|5|14|源自 亞瑪力 的人從 以法蓮 下來 ， 跟著你，你的族人 便雅憫 ； 有領袖從 瑪吉 下來， 手握官員權杖的從 西布倫 下來。
JUDG|5|15|以薩迦 的領袖與 底波拉 一起； 巴拉 怎樣， 以薩迦 也怎樣； 他跟隨 巴拉 衝下平原。 呂便 支派 有胸懷大志的人。
JUDG|5|16|你為何坐在羊圈內， 聽羊群中吹笛的聲音呢？ 呂便 支派具心有大謀的人。
JUDG|5|17|基列 安居在 約旦河 東。 但 為何住在船上呢？ 亞設 在海邊居住， 它在港口安居。
JUDG|5|18|西布倫 是拚命敢死的百姓， 拿弗他利 在田野的高處也是如此。 　
JUDG|5|19|「君王都來爭戰； 那時 迦南 諸王在 米吉多 水旁的 他納 爭戰， 卻得不到擄掠的銀錢。
JUDG|5|20|星宿從天上爭戰， 從它們的軌道攻擊 西西拉 。
JUDG|5|21|基順 的急流沖走他們， 古老的急流， 基順 的急流。 我的靈啊，努力前進！
JUDG|5|22|「那時馬蹄踢踏， 壯馬奔馳飛騰。
JUDG|5|23|「耶和華的使者說：『要詛咒 米羅斯 ， 重重詛咒其中的居民， 因為他們不來幫助耶和華， 不來幫助耶和華攻擊壯士。』
JUDG|5|24|「願 基尼 人 希百 的妻子 雅億 比眾婦人多得福氣， 比帳棚中的婦人更蒙福祉。
JUDG|5|25|西西拉 求水， 雅億 給他奶， 用貴重的碗裝乳酪給他。
JUDG|5|26|雅億 左手拿著帳棚的橛子， 右手拿著工匠的錘子， 擊打 西西拉 ，打碎他的頭， 打破穿透他的太陽穴。
JUDG|5|27|西西拉 在她腳下曲身，仆倒，躺臥， 在她腳下曲身，仆倒； 他在哪裏曲身，就在哪裏仆倒，死亡。
JUDG|5|28|「 西西拉 的母親從窗戶裏往外觀看， 她在窗格子中哀號： 『他的戰車為何遲遲未歸？ 他的車輪為何走得那麼慢呢？』
JUDG|5|29|她聰明的宮女回答她， 她也自言自語說：
JUDG|5|30|『或許他們得了戰利品而分， 每個壯士得了一兩個女子？ 西西拉 得了彩衣為擄物， 得了繡花的彩衣為掠物， 這兩面繡花的彩衣， 披在頸項上作為戰利品。』
JUDG|5|31|「耶和華啊，願你的仇敵都這樣滅亡！ 願愛你的人如太陽上升，大發光輝！」 於是這地太平四十年。
JUDG|6|1|以色列 人又行耶和華眼中看為惡的事，耶和華就把他們交在 米甸 手裏七年。
JUDG|6|2|米甸 的手戰勝 以色列 ； 以色列 人躲避 米甸 人，就在山中挖洞穴，挖洞建營寨。
JUDG|6|3|每當 以色列 人撒種之後， 米甸 、 亞瑪力 和東邊的人都上來攻打他們，
JUDG|6|4|對著他們安營，毀壞那地的農作物，直到 迦薩 ，沒有給 以色列 留下食物，牛、羊、驢也沒有留下。
JUDG|6|5|因為那些人帶著他們的牲畜和帳棚上來，像蝗蟲那樣多；人和駱駝無數，都進入境內，毀壞全地。
JUDG|6|6|以色列 因 米甸 的緣故極其窮乏， 以色列 人就呼求耶和華。
JUDG|6|7|以色列 人因 米甸 的緣故呼求耶和華的時候，
JUDG|6|8|耶和華就差遣先知到 以色列 人那裏，對他們說：「耶和華－ 以色列 的上帝如此說：『我曾領你們從 埃及 上來，從為奴之家出來，
JUDG|6|9|救你們脫離 埃及 人的手，脫離一切欺壓你們之人的手。我從你們面前趕出他們，把他們的地賜給你們。
JUDG|6|10|我對你們說，我是耶和華－你們的上帝。你們住在 亞摩利 人的地，不可敬畏他們的神明，但你們卻不聽從我的話。』」
JUDG|6|11|耶和華的使者到了 俄弗拉 ，坐在 亞比以謝 族 約阿施 的橡樹下。 約阿施 的兒子 基甸 正在醡酒池那裏打麥子，為了躲避 米甸 人。
JUDG|6|12|耶和華的使者向 基甸 顯現，對他說：「大能的勇士啊，耶和華與你同在！」
JUDG|6|13|基甸 對他說：「主啊，請容許我說，耶和華若與我們同在，我們怎麼會遭遇這一切事呢？我們的列祖告訴我們：『耶和華領我們從 埃及 上來』，他那奇妙的作為在哪裏呢？現在耶和華卻丟棄了我們，把我們交在 米甸 人的手掌中。」
JUDG|6|14|耶和華轉向 基甸 ，說：「去，靠著你這能力拯救 以色列 脫離 米甸 人的手掌。我豈不是已經差遣了你嗎？」
JUDG|6|15|基甸 對他說：「主啊，請容許我說，我怎能拯救 以色列 呢？看哪，我這一支在 瑪拿西 支派中是最貧寒的，我在我父家又是最微小的。」
JUDG|6|16|耶和華對他說：「我與你同在，你就必擊敗 米甸 ，如擊打一個人。」
JUDG|6|17|基甸 對他說：「我若在你眼前蒙恩，求你給我一個證據，證明是你在跟我說話。
JUDG|6|18|求你不要離開這裏，等我回來，將供物帶來，供在你面前。」他說：「我必等你回來。」
JUDG|6|19|基甸 去預備一隻小山羊，用一伊法細麵做了無酵餅，將肉放在籃子裏，將湯盛在壺中，帶到他那裏，在橡樹下獻上。
JUDG|6|20|上帝的使者對 基甸 說：「將肉和無酵餅放在這磐石上，把湯倒出來。」他就照樣做了。
JUDG|6|21|耶和華的使者伸出手裏的杖，杖頭一碰到肉和無酵餅，就有火從磐石中出來，吞滅了肉和無酵餅。耶和華的使者就從他眼前消失了。
JUDG|6|22|基甸 見他是耶和華的使者，就說：「哎呀！主耶和華啊！因為我真的面對面看見了耶和華的使者。」
JUDG|6|23|耶和華對他說：「安心吧，不要怕，你不會死。」
JUDG|6|24|於是 基甸 在那裏為耶和華築了一座壇，起名叫「耶和華沙龍」 。這壇至今還在 亞比以謝 族的 俄弗拉 。
JUDG|6|25|那夜，耶和華對 基甸 說：「你要把你父親的公牛，就是 那七歲的第二頭公牛取來，並拆毀你父親為 巴力 築的壇，砍下壇旁的 亞舍拉 ，
JUDG|6|26|在這堡壘頂上整整齊齊地為耶和華－你的上帝築一座壇，將第二頭公牛獻為燔祭，用你所砍下的 亞舍拉 當柴。」
JUDG|6|27|基甸 就從他僕人中選了十個人，照耶和華吩咐他的做了。他因怕父家和本城的人，不敢在白天做這事，就在夜間做。
JUDG|6|28|城裏的人清早起來，看哪， 巴力 的壇被拆毀，壇旁的 亞舍拉 被砍下，第二頭公牛獻在築好的壇上，
JUDG|6|29|就彼此問：「這是誰做的事呢？」他們尋找查訪之後，就說：「這是 約阿施 的兒子 基甸 做的事。」
JUDG|6|30|城裏的人對 約阿施 說：「把你的兒子交出來，我們要處死他，因為他拆毀了 巴力 的壇，砍下了壇旁的 亞舍拉 。」
JUDG|6|31|約阿施 對站著敵對他的眾人說：「你們是為 巴力 辯護嗎？你們要救它嗎？誰為它辯護，就在早晨把誰處死吧！ 巴力 如果是上帝，有人拆毀了它的壇，就讓它為自己辯護吧！」
JUDG|6|32|所以那日人稱 基甸 為 耶路巴力 ，意思是：「他拆毀了 巴力 的壇，讓 巴力 與他爭辯吧。」
JUDG|6|33|那時，所有的 米甸 人、 亞瑪力 人和東邊的人都聚集在一起，過了河，在 耶斯列 平原安營。
JUDG|6|34|耶和華的靈降在 基甸 身上；他吹角， 亞比以謝 族都聚集跟隨他。
JUDG|6|35|他派使者走遍 瑪拿西 ， 瑪拿西 人也聚集跟隨他。他又派使者到 亞設 、 西布倫 、 拿弗他利 ，他們也都上來會合。
JUDG|6|36|基甸 對上帝說：「你如果真的照你所說的，藉我的手拯救 以色列 ，
JUDG|6|37|看哪，我把一團羊毛放在禾場上，若單是羊毛上有露水，遍地都是乾的，我就知道你必照你所說的，藉我的手拯救 以色列 。」
JUDG|6|38|一切果然發生了。次日早晨 基甸 起來，把羊毛擰一擰，從羊毛中擠出露水來，裝滿一碗的水。
JUDG|6|39|基甸 又對上帝說：「求你不要向我發怒，我再說一次，讓我用羊毛再試一次，但願羊毛是乾的，遍地都有露水。」
JUDG|6|40|這夜，上帝也照樣做，遍地都有露水，只有羊毛是乾的。
JUDG|7|1|耶路巴力 ，就是 基甸 ，和所有跟隨他的人早晨起來，在 哈律泉 旁安營。 米甸 營在他北邊，靠近 摩利岡 的平原。
JUDG|7|2|耶和華對 基甸 說：「跟隨你的人太多，我不能把 米甸 交在他們手中，免得 以色列 向我自誇，說：『是我自己的手救了我。』
JUDG|7|3|現在你要向這百姓宣告說：『凡懼怕戰兢的，可以離開 基列山 回去。』」於是有二萬二千人回去，只剩下一萬人。
JUDG|7|4|耶和華對 基甸 說：「人還是太多。你要帶他們下到水旁，我好在那裏為你試試他們。我指著誰對你說：『這人可以跟你去』，他就可以跟你去；我指著誰對你說：『這人不可跟你去』，他就不可跟你去。」
JUDG|7|5|基甸 就帶百姓下到水旁。耶和華對 基甸 說：「凡用舌頭舔水像狗一樣舔的，要使他單獨站在一處；那些用雙膝跪下喝水的，也要使他單獨站在一處。」
JUDG|7|6|用手捧到嘴邊舔水的數目有三百人，其餘的百姓都用雙膝跪下喝水。
JUDG|7|7|耶和華對 基甸 說：「我要用這舔水的三百人拯救你們，把 米甸 交在你手中；其餘的百姓都可以各回自己的地方去。」
JUDG|7|8|百姓手裏拿著食物和角；其餘的 以色列 人， 基甸 都打發他們各自回到自己的帳棚，只留下這三百人。 米甸 營在他下邊的平原上。
JUDG|7|9|那夜，耶和華對 基甸 說：「起來，下去攻營，因我已把它交在你手中。
JUDG|7|10|倘若你害怕下去，可以帶你的僕人 普拉 下到那營裏去，
JUDG|7|11|你必聽見他們所說的，這樣你的手就有力量下去攻營。」於是 基甸 帶著僕人 普拉 下到軍營裏帶著兵器的人邊上。
JUDG|7|12|米甸 人、 亞瑪力 人和所有東邊的人都散佈在平原，如同蝗蟲那樣多。他們的駱駝無數，多如海邊的沙。
JUDG|7|13|基甸 到了那裏，看哪，有一人把夢告訴同伴說：「看哪，我做了一個夢。看哪，一個大麥餅滾入 米甸 營中，來到帳幕，把帳幕撞倒，帳幕就翻轉倒塌了。」
JUDG|7|14|同伴回答說：「這不是別的，而是 以色列 人 約阿施 的兒子 基甸 的刀。上帝已把 米甸 和全軍都交在他手中了。」
JUDG|7|15|基甸 聽見這夢的敘述和夢的解釋，就敬拜上帝。他回到 以色列 營中，說：「起來吧！耶和華已把 米甸 軍隊交在你們手中了。」
JUDG|7|16|於是 基甸 將三百人分成三隊，把角和空瓶交在每個人手中，瓶內有火把。
JUDG|7|17|他對他們說：「看著我，你們要照樣做。看哪，我來到營邊，我怎樣做，你們也要照樣做。
JUDG|7|18|我和所有跟隨我的人吹角的時候，你們也要在營的四圍吹角，喊叫：『為耶和華！為 基甸 ！』」
JUDG|7|19|基甸 和跟隨他的一百人，在半夜之初換崗哨的時候來到營旁。他們就吹角，打破手中的瓶；
JUDG|7|20|三隊的人都吹角，打破瓶子。他們左手拿著火把，右手拿著吹的角，喊叫：「耶和華和 基甸 的刀！」
JUDG|7|21|他們圍著軍營，各人站在自己的地方；全營的人都逃竄，一面喊，一面逃跑。
JUDG|7|22|三百人就吹角，耶和華使全營的人用刀自相擊殺。全營的人逃往 西利拉 的 伯‧哈示他 ，一直逃到靠近 他巴 的 亞伯‧米何拉 。
JUDG|7|23|從 拿弗他利 、 亞設 和 瑪拿西 全地來的 以色列 人被召來，追趕 米甸 人。
JUDG|7|24|基甸 也派人走遍 以法蓮 山區，說：「你們下來迎擊 米甸 人，在他們的前面沿著 約旦河 把守渡口，直到 伯‧巴拉 。」於是 以法蓮 眾人聚集，沿著 約旦河 把守渡口，直到 伯‧巴拉 。
JUDG|7|25|他們捉住了 米甸 的兩個領袖， 俄立 和 西伊伯 。他們在 俄立 磐石上殺了 俄立 ，在 西伊伯 酒池那裏殺了 西伊伯 。他們追趕 米甸 人，把 俄立 和 西伊伯 的首級帶到 約旦河 對岸，到 基甸 那裏。
JUDG|8|1|以法蓮 人對 基甸 說：「你去與 米甸 爭戰，沒有召我們同去，你為甚麼這樣待我們呢？」他們就和 基甸 激烈地爭吵。
JUDG|8|2|基甸 對他們說：「我現在所做的怎麼與你們所做的相比呢？ 以法蓮 拾取剩下的葡萄不強過 亞比以謝 族所摘的葡萄嗎？
JUDG|8|3|上帝已把 米甸 的兩個領袖 俄立 和 西伊伯 交在你們手中；我所做的怎能與你們所做的相比呢？」 基甸 說了這話，他們對他的怒氣就消了。
JUDG|8|4|基甸 和跟隨他的三百人來到 約旦河 ，渡了過去；他們雖然疲乏，還是追趕。
JUDG|8|5|基甸 對 疏割 人說：「請你們拿幾塊餅來給跟隨我的百姓，因為他們疲乏了。我正在追擊 米甸 王 西巴 和 撒慕拿 。」
JUDG|8|6|疏割 人的領袖回答說：「 西巴 和 撒慕拿 的手掌現在已經在你手裏，因此我們該將餅送給你的軍隊嗎？」
JUDG|8|7|基甸 說：「好吧！耶和華將 西巴 和 撒慕拿 交在我手之後，我必用曠野的荊棘和枳條鞭打你們。」
JUDG|8|8|基甸 從那裏上到 毗努伊勒 ，對那裏的人也提出同樣的請求； 毗努伊勒 人給他的答覆跟 疏割 人的答覆一樣。
JUDG|8|9|他也對 毗努伊勒 人說：「我平平安安回來的時候，必拆毀這城樓。」
JUDG|8|10|那時 西巴 和 撒慕拿 ，以及跟隨他們的軍隊都在 加各 ，約有一萬五千人，是東邊的人全軍所剩下的，因為拿刀戰死的約有十二萬人。
JUDG|8|11|基甸 從 挪巴 和 約比哈 的東邊，從住帳棚人 的路上去，趁 米甸 的軍兵以為安全的時候攻擊他們。
JUDG|8|12|西巴 和 撒慕拿 逃跑； 基甸 追趕他們，捉住 米甸 的兩個王 西巴 和 撒慕拿 ，使他們全軍潰散。
JUDG|8|13|約阿施 的兒子 基甸 從戰場，沿著 希列斯 斜坡回來，
JUDG|8|14|捉住 疏割 人的一個少年，查問他。他就為 基甸 寫下 疏割 的領袖和長老的名字，共七十七人。
JUDG|8|15|基甸 到了 疏割 人那裏，說：「你們從前譏笑我說：『 西巴 和 撒慕拿 的手掌現在已經在你手裏，因此我們該將餅送給跟隨你的疲乏的人嗎？』看哪， 西巴 和 撒慕拿 在這裏。」
JUDG|8|16|於是他拿住城內的長老，用曠野的荊棘和枳條責打 疏割 人。
JUDG|8|17|他又拆了 毗努伊勒 的城樓，殺了城裏的人。
JUDG|8|18|基甸 對 西巴 和 撒慕拿 說：「你們在 他泊山 所殺的人是甚麼樣子的？」他們說：「他們很像你，個個都有王子的樣子。」
JUDG|8|19|基甸 說：「他們都是我的兄弟，我母親的兒子。我指著永生的耶和華起誓，你們若存留他們的性命，我就不殺你們了。」
JUDG|8|20|他對他的長子 益帖 說：「你起來殺他們！」但是這少年害怕，不敢拔刀，因為他還是個少年。
JUDG|8|21|西巴 和 撒慕拿 說：「你自己起來殺我們吧！因為人如何，力量也如何。」 基甸 就起來，殺了 西巴 和 撒慕拿 ，取了他們駱駝頸項上的月牙圈。
JUDG|8|22|以色列 人對 基甸 說：「你既然救我們脫離 米甸 的手，願你治理我們，你的兒子孫子也治理我們。」
JUDG|8|23|基甸 對他們說：「我不治理你們，我的兒子也不治理你們，耶和華會治理你們。」
JUDG|8|24|基甸 又對他們說：「我有一件事求你們，請你們各人把所奪的耳環給我。」因敵人都戴金耳環，他們是 以實瑪利 人。
JUDG|8|25|以色列 人說：「我們情願送給你！」他們就鋪開一件外衣，各人將所奪的耳環丟在上面。
JUDG|8|26|基甸 所要求的金耳環，重一千七百舍客勒金子。此外還有 米甸 王所戴的月牙圈、耳環，和所穿的紫色衣服，以及駱駝頸項上的鏈子。
JUDG|8|27|基甸 以此造了一個以弗得，設立在他的本城 俄弗拉 。全 以色列 就在那裏拜這以弗得行淫，這就成了 基甸 和他全家的圈套。
JUDG|8|28|這樣， 米甸 就被 以色列 人制伏了，再也不能抬頭。 基甸 還在的日子，這地太平四十年。
JUDG|8|29|約阿施 的兒子 耶路巴力 回去，住在自己家裏。
JUDG|8|30|基甸 有七十個親生的兒子，因為他有許多妻子。
JUDG|8|31|他在 示劍 的妾也為他生了一個兒子， 基甸 給他起名叫 亞比米勒 。
JUDG|8|32|約阿施 的兒子 基甸 年紀老邁而死，葬在 亞比以謝 族的 俄弗拉 ，他父親 約阿施 的墳墓裏。
JUDG|8|33|基甸 死後， 以色列 人又去隨從諸 巴力 而行淫，以 巴力‧比利土 為他們的神明。
JUDG|8|34|以色列 人不記得耶和華－他們的上帝，就是那位拯救他們脫離四圍仇敵之手的，
JUDG|8|35|也不照著 耶路巴力 ，就是 基甸 向 以色列 所施的恩惠善待他的家。
JUDG|9|1|耶路巴力 的兒子 亞比米勒 到 示劍 他的母舅那裏，對他們和他外祖父全家的人說：
JUDG|9|2|「請你們問 示劍 所有的居民：『是 耶路巴力 的眾兒子七十人都治理你們好，還是一人治理你們好呢？』你們要記得，我是你們的骨肉。」
JUDG|9|3|他的母舅們為他把這一切話說給 示劍 所有的居民聽，他們的心就傾向 亞比米勒 ，因為他們說：「他是我們的弟兄。」
JUDG|9|4|他們從 巴力‧比利土 的廟中取了七十銀子給 亞比米勒 ， 亞比米勒 用這些錢雇了一些無賴匪徒跟隨他。
JUDG|9|5|他來到 俄弗拉 他父親的家，在一塊磐石上把他的兄弟，就是 耶路巴力 的七十個兒子都殺了，只剩下 耶路巴力 的小兒子 約坦 ，因為他躲了起來。
JUDG|9|6|示劍 所有的居民和全 伯‧米羅 都聚集在一起，到 示劍 橡樹旁的柱子那裏，立 亞比米勒 為王。
JUDG|9|7|有人將這事告訴 約坦 ，他就去站在 基利心山 頂上，高聲喊叫，對他們說：「 示劍 的居民哪，你們要聽我，上帝也就會聽你們。
JUDG|9|8|有一次，樹木要膏一王治理他們，就去對橄欖樹說：『請你來作王治理我們！』
JUDG|9|9|橄欖樹對它們說：『我豈可停止生產使神明和人得尊榮的油，而行走飄搖在眾樹之上呢？』
JUDG|9|10|樹木對無花果樹說：『請你來作王治理我們！』
JUDG|9|11|無花果樹對它們說：『我豈可停止結甜美的果子，而行走飄搖在眾樹之上呢？』
JUDG|9|12|樹木對葡萄樹說：『請你來作王治理我們！』
JUDG|9|13|葡萄樹對它們說：『我豈可停止出產使神明和人歡樂的新酒，而行走飄搖在眾樹之上呢。』
JUDG|9|14|眾樹對荊棘說：『請你來作王治理我們！』
JUDG|9|15|荊棘對眾樹說：『你們若真的要膏我作王治理你們，就要來到我的蔭下尋求庇護；不然，願火從荊棘裏出來，吞滅 黎巴嫩 的香柏樹。』
JUDG|9|16|「現在你們若以誠實正直立 亞比米勒 為王，若善待 耶路巴力 和他的家，若照他手所做的回報他─
JUDG|9|17|從前我父為你們爭戰，冒生命的危險救你們脫離 米甸 的手，
JUDG|9|18|但是你們如今起來攻擊我的父家，在一塊磐石上把他的七十個兒子全殺了，又立他使女所生的兒子 亞比米勒 為 示劍 居民的王，因為他是你們的弟兄─
JUDG|9|19|你們如今若以誠實正直對待 耶路巴力 和他的家，就可以因 亞比米勒 歡樂，他也可以因你們歡樂；
JUDG|9|20|不然，願火從 亞比米勒 發出，吞滅 示劍 居民和 伯‧米羅 ，又願火從 示劍 居民和 伯‧米羅 發出，吞滅 亞比米勒 。」
JUDG|9|21|約坦 因躲避他的兄弟 亞比米勒 就逃跑，去到 比珥 ，住在那裏。
JUDG|9|22|亞比米勒 治理 以色列 三年。
JUDG|9|23|上帝派邪靈到 亞比米勒 和 示劍 居民中間， 示劍 居民就以詭詐待 亞比米勒 。
JUDG|9|24|這是要使 耶路巴力 七十個兒子受害所流的血，歸於他們的兄弟 亞比米勒 ，因他殺害他們，也歸於那些出手幫助他殺害兄弟的 示劍 居民。
JUDG|9|25|示劍 居民在山頂上設下埋伏，等候 亞比米勒 。凡沿著那條路，從他們那裏經過的人，他們就搶劫。有人把這事告訴 亞比米勒 。
JUDG|9|26|以別 的兒子 迦勒 和他的弟兄經過，來到 示劍 ， 示劍 居民都信任他。
JUDG|9|27|他們出到田間，摘下葡萄，踹酒，作樂。他們進入他們神明的廟中吃喝，詛咒 亞比米勒 。
JUDG|9|28|以別 的兒子 迦勒 說：「 亞比米勒 是誰，我們 示劍 人是誰，叫我們服事他呢？他不是 耶路巴力 的兒子嗎？他的助手不是 西布勒 嗎？你們應當服事 示劍 的父親 哈抹 的後裔！我們為何要服事 亞比米勒 呢？
JUDG|9|29|惟願這民歸到我的手下，我就除掉 亞比米勒 。」他就對 亞比米勒 說：「增加你的軍兵，出來吧！」
JUDG|9|30|西布勒 市長聽見 以別 的兒子 迦勒 的話，就怒氣大發。
JUDG|9|31|他悄悄地派一些使者到 亞比米勒 那裏，說：「看哪， 以別 的兒子 迦勒 和他的弟兄到了 示劍 。看哪，他們煽動那城攻擊你。
JUDG|9|32|現在，你和跟隨你的百姓要夜間起來，在田間埋伏。
JUDG|9|33|早晨太陽一出，你就趁早攻城。看哪， 迦勒 和跟隨他的百姓出來攻擊你的時候，你就全力對付他們。」
JUDG|9|34|於是， 亞比米勒 和跟隨他的眾百姓夜間起來，兵分四隊，埋伏攻擊 示劍 。
JUDG|9|35|以別 的兒子 迦勒 出去，站在城門口。 亞比米勒 和跟隨他的百姓從埋伏之處起來。
JUDG|9|36|迦勒 看見百姓，就對 西布勒 說：「看哪，有百姓從山頂上下來。」 西布勒 對他說：「你把山的影子看作是人了。」
JUDG|9|37|迦勒 又繼續講，他說：「看哪，有百姓從地的高處下來，又有一隊從 米惡尼尼 橡樹 的路前來。」
JUDG|9|38|西布勒 對他說：「你所誇口的在哪裏呢？你曾說：『 亞比米勒 是誰，叫我們服事他呢？』這不是你所藐視的百姓嗎？你現在出去，與他們交戰吧！」
JUDG|9|39|於是 迦勒 率領 示劍 居民出去，與 亞比米勒 交戰。
JUDG|9|40|亞比米勒 追趕 迦勒 ， 迦勒 在他面前逃跑。有許多人被刺傷仆倒，直到城門口。
JUDG|9|41|亞比米勒 住在 亞魯瑪 。 西布勒 趕出 迦勒 和他的弟兄，不准他們住在 示劍 。
JUDG|9|42|次日，百姓出到田間，有人告訴 亞比米勒 ，
JUDG|9|43|他就帶領百姓，把他們分成三隊，埋伏在田間窺探。看哪， 示劍 居民從城裏出來，他就起來擊殺他們。
JUDG|9|44|亞比米勒 和跟隨他的一隊向前衝，站在城門口；另外兩隊直衝向田間，擊殺了眾人。
JUDG|9|45|亞比米勒 攻城一整天，將城奪取，殺了其中的百姓，把城拆毀，撒上了鹽。
JUDG|9|46|示劍 城樓裏所有的居民聽見了，就進入 伊勒‧比利土 廟的地窖裏。
JUDG|9|47|有人告訴 亞比米勒 ， 示劍 城樓裏所有的居民都聚在一起。
JUDG|9|48|亞比米勒 和所有跟隨他的百姓都上 撒們山 去。 亞比米勒 手拿斧子，砍下一根樹枝，舉起來，扛在肩上，對跟隨他的百姓說：「你們看我做甚麼，就趕快照樣做。」
JUDG|9|49|眾百姓也都各砍一根樹枝，跟 亞比米勒 走，把樹枝堆在地窖上，放火燒地窖。這樣， 示劍 城樓裏所有的人都死了，男女約有一千。
JUDG|9|50|亞比米勒 到 提備斯 ，對著 提備斯 安營，攻取了那城。
JUDG|9|51|城中有一座堅固的樓；城裏所有的居民，無論男女，都逃到那裏，關上門，上了樓頂。
JUDG|9|52|亞比米勒 到了樓前，攻打它。他挨近樓門，要放火焚燒。
JUDG|9|53|有一個婦人把一塊上磨石拋在 亞比米勒 的頭上，打破了他的頭蓋骨。
JUDG|9|54|他就急忙叫拿他兵器的青年來，對他說：「拔出你的刀來，殺了我吧！免得有人提到我說：『他被一個婦人殺了。』」於是那青年把他刺透，他就死了。
JUDG|9|55|以色列 人見 亞比米勒 死了，就各回自己的地方去了。
JUDG|9|56|這樣，上帝報應了 亞比米勒 向他父親所做的惡事，就是殺了自己七十個兄弟。
JUDG|9|57|示劍 人的一切惡事，上帝也都報應在他們頭上； 耶路巴力 的兒子 約坦 的詛咒都臨到他們身上了。
JUDG|10|1|亞比米勒 以後， 陀拉 興起，拯救 以色列 ，他是 朵多 的孫子， 普瓦 的兒子， 以薩迦 人，住在 以法蓮 山區的 沙密 。
JUDG|10|2|陀拉 作 以色列 的士師二十三年。他死了，葬在 沙密 。
JUDG|10|3|陀拉 以後有 基列 人 睚珥 興起，作 以色列 的士師二十二年。
JUDG|10|4|他有三十個兒子，騎著三十匹驢駒。他們有三十座城，叫作 哈倭特‧睚珥 ，直到如今，都在 基列 地。
JUDG|10|5|睚珥 死了，葬在 加們 。
JUDG|10|6|以色列 人又行耶和華眼中看為惡的事，去事奉諸 巴力 和 亞斯她錄 ，以及 亞蘭 的神明、 西頓 的神明、 摩押 的神明、 亞捫 人的神明、 非利士 人的神明。他們離棄耶和華，不事奉他。
JUDG|10|7|耶和華的怒氣向 以色列 發作，把他們交給 非利士 人和 亞捫 人的手中。
JUDG|10|8|從那年起，他們欺壓迫害 以色列 人，在 約旦河 東， 亞摩利 人境內， 基列 一帶所有的 以色列 人，長達十八年。
JUDG|10|9|亞捫 人渡過 約旦河 去攻打 猶大 和 便雅憫 ，以及 以法蓮 家族。 以色列 的處境非常困苦。
JUDG|10|10|以色列 人哀求耶和華說：「我們得罪了你，因為我們離棄了我們的上帝，去事奉諸 巴力 。」
JUDG|10|11|耶和華對 以色列 人說：「我豈沒有救你們脫離 埃及 人、 亞摩利 人、 亞捫 人和 非利士 人嗎？
JUDG|10|12|西頓 人、 亞瑪力 人和 馬雲 人 欺壓你們，你們哀求我，我也拯救你們脫離他們的手。
JUDG|10|13|你們竟離棄我去事奉別神！所以我不再救你們了。
JUDG|10|14|你們去哀求你們所選擇的神明；你們遭遇急難的時候，讓它們救你們吧！」
JUDG|10|15|以色列 人對耶和華說：「我們犯罪了，照你看為好的待我們，只求你今日拯救我們吧！」
JUDG|10|16|以色列 人就除掉他們中間的外邦神明，事奉耶和華。耶和華因 以色列 所受的苦難而心裏焦急。
JUDG|10|17|亞捫 人被召來，在 基列 安營； 以色列 人也聚集，在 米斯巴 安營。
JUDG|10|18|基列 百姓中的領袖彼此說：「誰領先出去攻打 亞捫 人，誰就作 基列 所有居民的領袖。」
JUDG|11|1|基列 人 耶弗他 是個大能的勇士，是妓女的兒子。 基列 生了 耶弗他 。
JUDG|11|2|基列 的妻子也給他生了幾個兒子。他妻子生的兒子長大後，就把 耶弗他 趕出去，說：「你不可在我們父家繼承產業，因為你是別的女人生的兒子。」
JUDG|11|3|耶弗他 就逃離他的兄弟，住在 陀伯 地。有些無賴的人聚集在他那裏，與他一同出入。
JUDG|11|4|過了些日子， 亞捫 人攻打 以色列 。
JUDG|11|5|亞捫 人攻打 以色列 的時候， 基列 的長老去請 耶弗他 從 陀伯 地回來。
JUDG|11|6|他們對 耶弗他 說：「請你來作我們的指揮官，好讓我們跟 亞捫 人打仗。」
JUDG|11|7|耶弗他 對 基列 的長老說：「你們不是恨我，把我趕出父家嗎？現在你們遭遇急難，為何到我這裏來呢？」
JUDG|11|8|基列 的長老對 耶弗他 說：「現在我們回到你這裏，是要請你同我們去跟 亞捫 人打仗，作 基列 所有居民的領袖。」
JUDG|11|9|耶弗他 對 基列 的長老說：「若你們請我回去跟 亞捫 人打仗，耶和華把他們交給我，我就作你們的領袖。」
JUDG|11|10|基列 的長老對 耶弗他 說：「有耶和華在你我之間作證，我們必定照你的話做。」
JUDG|11|11|於是 耶弗他 與 基列 的長老同去，百姓就立 耶弗他 作他們的領袖和指揮官。 耶弗他 在 米斯巴 將他一切的事陳述在耶和華面前。
JUDG|11|12|耶弗他 派使者到 亞捫 人的王那裏，說：「你與我有甚麼相干，竟來到我這裏攻打我的地呢？」
JUDG|11|13|亞捫 人的王對 耶弗他 的使者說：「因為 以色列 從 埃及 上來的時候佔據我的地，從 亞嫩河 到 雅博河 ，直到 約旦河 。現在你要和平歸還這些地方！」
JUDG|11|14|耶弗他 又派使者到 亞捫 人的王那裏，
JUDG|11|15|對他說：「 耶弗他 如此說： 以色列 並沒有佔據 摩押 地和 亞捫 人的地。
JUDG|11|16|以色列 人從 埃及 上來，是經過曠野到 紅海 ，來到 加低斯 。
JUDG|11|17|那時， 以色列 派使者去 以東 王那裏，說：『求你讓我穿越你的地。』 以東 王卻不聽。 以色列 又照樣派使者去 摩押 王那裏，他也不肯。於是 以色列 人就住在 加低斯 。
JUDG|11|18|他們又經過曠野，繞過 以東 地和 摩押 地，到 摩押 地的東邊 ，在 亞嫩河 邊安營，並沒有進入 摩押 的境內，因為 亞嫩河 是 摩押 的邊界。
JUDG|11|19|以色列 派使者去 亞摩利 王，就是 希實本 王 西宏 那裏； 以色列 對他說：『求你讓我們穿越你的地，到我自己的地方去。』
JUDG|11|20|西宏 卻不信任 以色列 ，不讓他們穿越他的疆界。他召集了他的眾百姓在 雅雜 安營，與 以色列 爭戰。
JUDG|11|21|耶和華－ 以色列 的上帝將 西宏 和他的眾百姓都交在 以色列 手中， 以色列 人就擊殺他們，佔領了那地居民 亞摩利 人的全地。
JUDG|11|22|他們佔領了 亞摩利 人所有的疆土，從 亞嫩河 到 雅博河 ，從曠野直到 約旦河 。
JUDG|11|23|耶和華－ 以色列 的上帝如今從他百姓 以色列 面前趕出 亞摩利 人，你竟要佔領它嗎？
JUDG|11|24|你不是已經得了你的神明 基抹 賜給你的地為業嗎？耶和華－我們的上帝在我們面前所趕出的，我們也要得它為業。
JUDG|11|25|現在你比 西撥 的兒子 摩押 王 巴勒 還強嗎？他真的曾與 以色列 爭執，或是真的與他們爭戰了嗎？
JUDG|11|26|以色列 人住 希實本 和所屬的鄉鎮， 亞羅珥 和所屬的鄉鎮，以及沿著 亞嫩河 的一切城鎮，已經有三百年了。在這期間，你們為甚麼不取回呢？
JUDG|11|27|我並沒有得罪你，你卻要攻打我，加害於我。願審判人的耶和華今日在 以色列 人和 亞捫 人之間判斷是非。」
JUDG|11|28|但 亞捫 人的王不聽 耶弗他 傳達給他的話。
JUDG|11|29|耶和華的靈降在 耶弗他 身上，他就經過 基列 和 瑪拿西 ，經過 基列 的 米斯巴 ，又從 基列 的 米斯巴 過到 亞捫 人那裏。
JUDG|11|30|耶弗他 向耶和華許願，說：「你若真的將 亞捫 人交在我手中，
JUDG|11|31|我從 亞捫 人那裏平平安安回來的時候，無論誰先從我家門出來迎接我，就要歸給耶和華，我必將他獻上作為燔祭。」
JUDG|11|32|於是 耶弗他 往 亞捫 人那裏去，與他們爭戰。耶和華將他們交在他手中，
JUDG|11|33|他就徹底擊敗他們，從 亞羅珥 到 米匿 ，直到 亞備勒‧基拉明 ，攻取了二十座城。這樣， 亞捫 人就在 以色列 人面前被制伏了。
JUDG|11|34|耶弗他 回 米斯巴 去，到了自己的家，看哪，他女兒拿著手鼓跳舞出來迎接他。她是 耶弗他 的獨生女，除她以外，沒有別的兒女。
JUDG|11|35|耶弗他一看見她，就撕裂衣服，說：「哀哉！我的女兒啊，你使我非常悲痛，叫我十分為難了。因為我已經向耶和華開了口，不能收回。」
JUDG|11|36|他女兒對他說：「我的父親啊，你既向耶和華開了口，就當照你口中所說的向我行，因為耶和華已經在你的仇敵 亞捫 人身上為你報了仇。」
JUDG|11|37|她又對父親說：「我只求你這一件事，給我兩個月，讓我和同伴下到山裏，好為我的童貞哀哭。」
JUDG|11|38|耶弗他 說：「你去吧！」他就讓她離開兩個月。她和同伴去了，在山裏為她的童貞哀哭。
JUDG|11|39|過了兩個月，她回到父親那裏，父親就照所許的願向她行了。她從來沒有親近男人。於是 以色列 中有個風俗，
JUDG|11|40|每年按著日期 以色列 的女子要去為 基列 人 耶弗他 的女兒哀哭四天。
JUDG|12|1|以法蓮 人被召來，渡河來到 撒分 。他們對 耶弗他 說：「你去與 亞捫 人爭戰，為甚麼沒有召我們同去呢？我們必用火將你和你的家燒了。」
JUDG|12|2|耶弗他 對他們說：「我和我的百姓與 亞捫 人有極大的衝突；我曾召你們來，你們卻沒有來救我脫離他們的手。
JUDG|12|3|我見你們不來救我，就拚了命前去攻打 亞捫 人，耶和華就將他們交在我手中。你們今日為甚麼上我這裏來攻打我呢？」
JUDG|12|4|於是 耶弗他 召集 基列 所有的人，要與 以法蓮 人爭戰。 基列 人擊殺 以法蓮 人，因 以法蓮 人曾說：「你們 基列 人在 以法蓮 和 瑪拿西 中，不過是 以法蓮 逃亡的人而已。」
JUDG|12|5|基列 人把守 約旦河 的渡口，不許 以法蓮 人過去。逃跑的 以法蓮 人若說：「讓我過河。」 基列 人就問他說：「你是不是 以法蓮 人？」他若說：「不是」，
JUDG|12|6|基列 人就對他說：「你說『示播列』。」 以法蓮 人因為發音不準，就會說成「西播列」。 基列 人就捉住他，在 約旦河 的渡口把他殺了。那時， 以法蓮 人被殺的有四萬二千人。
JUDG|12|7|耶弗他 作 以色列 的士師六年。 基列 人 耶弗他 死了，葬在 基列 的城裏 。
JUDG|12|8|耶弗他 以後，有 伯利恆 人 以比讚 作 以色列 的士師。
JUDG|12|9|他有三十個兒子。他把三十個女兒都嫁出去了，也為他的兒子從外面娶了三十個媳婦。他作 以色列 的士師七年。
JUDG|12|10|以比讚 死了，葬在 伯利恆 。
JUDG|12|11|以比讚 以後，有 西布倫 人 以倫 作 以色列 的士師，他作 以色列 的士師十年。
JUDG|12|12|西布倫 人 以倫 死了，葬在 西布倫 地的 亞雅崙 。
JUDG|12|13|以倫 以後，有 比拉頓 人 希列 的兒子 押頓 作 以色列 的士師。
JUDG|12|14|他有四十個兒子，三十個孫子，騎著七十匹驢駒。 押頓 作 以色列 的士師八年。
JUDG|12|15|比拉頓 人 希列 的兒子 押頓 死了，葬在 以法蓮 地的 比拉頓 ，就在 亞瑪力 人的山區。
JUDG|13|1|以色列 人又行耶和華眼中看為惡的事，耶和華將他們交在 非利士 人手中四十年。
JUDG|13|2|那時，有一個 但 支派的 瑣拉 人，名叫 瑪挪亞 。他的妻子不懷孕，不生育。
JUDG|13|3|耶和華的使者向那婦人顯現，對她說：「看哪，以前你不懷孕，不生育，如今你必懷孕生一個兒子。
JUDG|13|4|現在你要謹慎，清酒烈酒都不可喝，任何不潔之物都不可吃，
JUDG|13|5|看哪，你必懷孕，生一個兒子。不可用剃刀剃他的頭，因為這孩子一出母胎就歸給上帝作拿細耳人。他必開始拯救 以色列 脫離 非利士 人的手。」
JUDG|13|6|那婦人來對丈夫說：「有一個神人到我這裏來，他的容貌如上帝使者的容貌，非常可畏。我沒有問他從哪裏來，他也沒有把他的名字告訴我。
JUDG|13|7|他對我說：『看哪，你要懷孕，生一個兒子 。現在，清酒烈酒都不可喝，任何不潔之物都不可吃，因為這孩子從出母胎一直到死的那一天，要歸給上帝作拿細耳人。』」
JUDG|13|8|瑪挪亞 祈求耶和華說：「主啊，求你再差遣那神人到我們這裏來，指示我們對這將要生的孩子該怎樣作。」
JUDG|13|9|上帝垂聽了 瑪挪亞 的聲音。那婦人坐在田間的時候，上帝的使者又到她那裏，但是她的丈夫 瑪挪亞 沒有同她在一起。
JUDG|13|10|婦人急忙跑去告訴丈夫，對他說：「看哪，那日到我這裏來的人又向我顯現了。」
JUDG|13|11|瑪挪亞 起來，跟隨他的妻子來到那人那裏，對他說：「你就是跟這婦人說話的那個人嗎？」他說：「是我。」
JUDG|13|12|瑪挪亞 說：「現在，願你的話應驗！這孩子該如何管教呢？他當做甚麼呢？」
JUDG|13|13|耶和華的使者對 瑪挪亞 說：「我告訴這婦人的一切事，她都要遵守。
JUDG|13|14|葡萄樹所結的不可吃，清酒烈酒都不可喝，任何不潔之物也不可吃。凡我所吩咐的，她都當遵守。」
JUDG|13|15|瑪挪亞 對耶和華的使者說：「請容許我們留你下來，好為你預備一隻小山羊。」
JUDG|13|16|耶和華的使者對 瑪挪亞 說：「你雖然留我，我卻不吃你的食物。你若預備燔祭，就當獻給耶和華。」因 瑪挪亞 不知道他是耶和華的使者。
JUDG|13|17|瑪挪亞 對耶和華的使者說：「請問大名？好讓我們在你的話應驗的時候尊敬你。」
JUDG|13|18|耶和華的使者對他說：「你何必問我的名字呢？我的名字是奇妙的。」
JUDG|13|19|瑪挪亞 取一隻小山羊和素祭，在磐石上獻給耶和華。他行奇妙的事， 瑪挪亞 和他的妻子觀看，
JUDG|13|20|火焰從壇上往上升，耶和華的使者也在壇上的火焰中升上去了。 瑪挪亞 和他的妻子看見，就臉伏於地。
JUDG|13|21|耶和華的使者不再向 瑪挪亞 和他的妻子顯現了。那時， 瑪挪亞 才知道他是耶和華的使者。
JUDG|13|22|瑪挪亞 對他的妻子說：「我們一定會死，因為我們看見了上帝。」
JUDG|13|23|他的妻子卻對他說：「耶和華若有意要我們死，就不會從我們手中接受燔祭和素祭，不會將這一切事指示我們，這時也不會讓我們聽到這話。」
JUDG|13|24|後來婦人生了一個兒子，給他起名叫 參孫 。孩子漸漸長大，耶和華賜福給他。
JUDG|13|25|在 瑣拉 和 以實陶 之間的 瑪哈尼‧但 ，耶和華的靈開始感動 參孫 。
JUDG|14|1|參孫 下到 亭拿 ，在 亭拿 看見一個女子，是 非利士 人的女兒。
JUDG|14|2|他上來告訴他父母說：「我在 亭拿 看見一個女子，是 非利士 人的女兒，現在請你們給我娶她為妻。」
JUDG|14|3|他父母對他說：「在你弟兄的女兒中，或在本族所有的人中，難道沒有女子嗎？你何必在未受割禮的 非利士 人中去娶妻呢？」 參孫 對他父親說：「請你給我娶那女子，因為我喜歡她。」
JUDG|14|4|他的父母並不知道這事是出於耶和華，因為他在找機會攻擊 非利士 人。那時， 非利士 人轄制 以色列 人。
JUDG|14|5|參孫 跟他父母下 亭拿 去，他們到了 亭拿 的葡萄園。看哪，有一隻少壯獅子對著他吼叫。
JUDG|14|6|耶和華的靈大大感動 參孫 ，他就手無寸鐵撕裂獅子，如撕裂小山羊一樣。他做這事，並沒有告訴他的父母親。
JUDG|14|7|參孫 下去跟那女子說話，看著就喜歡她。
JUDG|14|8|過了些日子，他回來要娶那女子，繞道去看獅子的殘骸，看哪，有一群蜜蜂在獅子的屍體內，也有蜜在裏面。
JUDG|14|9|他就取了蜜，放在手掌上，邊走邊吃。他到了父母那裏，給他們蜜，他們也吃了。但他沒有告訴他們，這蜜是從獅子的屍體內取來的。
JUDG|14|10|他父親下到女子那裏去。 參孫 在那裏擺設宴席， 因為這是當時年輕人的習俗。
JUDG|14|11|他們看見 參孫 ，就請了三十個人陪伴他。
JUDG|14|12|參孫 對他們說：「我給你們出個謎語，你們若能在七日宴席之內，猜出謎底告訴我，我就給你們三十件細麻內衣和三十套更換的衣服。
JUDG|14|13|但你們若不能告訴我，你們就給我三十件細麻內衣和三十套更換的衣服。」他們對他說：「請把謎語說給我們聽。」
JUDG|14|14|參孫 對他們說： 「吃的從吃者出來； 甜的從強者出來」。 三日之久，他們都猜不出謎語來。
JUDG|14|15|第七日 ，他們對 參孫 的妻子說：「你哄騙你的丈夫，為我們探出謎底來，否則我們就用火燒你和你的父家。你們請我們來，是不是要奪走我們所有的呢？」
JUDG|14|16|參孫 的妻子在丈夫面前哭哭啼啼說：「你只是恨我，並不愛我。你給我本族的人出謎語，卻不把謎底告訴我。」 參孫 對她說：「看哪，連我的父母我都沒有說，我怎麼可以告訴你呢？」
JUDG|14|17|在七日宴席中，她一直在丈夫面前哭哭啼啼。第七日， 參孫 因妻子的催逼就把謎底告訴了她。她把謎底告訴了她本族的人。
JUDG|14|18|第七日日落以前，那城裏的人對 參孫 說： 「有甚麼比蜜還甜呢？ 有甚麼比獅子更強呢？」 參孫 對他們說： 「你們若不用我的母牛犢耕地， 就無法猜出我的謎底來。」
JUDG|14|19|耶和華的靈大大感動 參孫 ，他就下到 亞實基倫 ，擊殺了三十個人，奪了他們身上的衣服，把衣服給了猜出謎語的人。 參孫 怒氣大發，就上他父親的家去了。
JUDG|14|20|參孫 的妻子就歸了 參孫 的一個同伴，就是作過他伴郎的。
JUDG|15|1|過了些日子，在割麥子的時候， 參孫 帶著一隻小山羊去探望他的妻子，說：「我要進內室到我妻子那裏。」他岳父不許他進去。
JUDG|15|2|他岳父說：「我以為你極其恨她，因此我把她給了你的同伴。她妹妹不是比她更美麗嗎？你可以娶來代替她！」
JUDG|15|3|參孫 對他們說：「這一次我若加害 非利士 人，就不算是我的錯了。」
JUDG|15|4|於是 參孫 去捉了三百隻狐狸，把牠們的尾巴一對一對地綁住，再將火把綁在兩條尾巴中間。
JUDG|15|5|他點著火把，把狐狸放進 非利士 人直立的莊稼，把堆積的禾捆和直立的莊稼，葡萄園、橄欖園全都燒了。
JUDG|15|6|非利士 人說：「這事是誰做的呢？」有人說：「是 亭拿 人的女婿 參孫 做的，因為他岳父把他的妻子給了他的同伴。」於是 非利士 人上去，用火燒了女子和她的父親。
JUDG|15|7|參孫 對他們說：「你們既然這麼做，我必向你們報仇才肯罷休。」
JUDG|15|8|參孫 狠狠擊殺他們，把他們連腿帶腰都砍了。過後，他就下去，住在 以坦巖 的石洞裏。
JUDG|15|9|非利士 人上去，安營在 猶大 ，侵犯 利希 。
JUDG|15|10|猶大 人說：「你們為何上來攻擊我們呢？」他們說：「我們上來是要捆綁 參孫 ，照他向我們所做的對待他。」
JUDG|15|11|於是，三千 猶大 人下到 以坦巖 的石洞裏，對 參孫 說：「 非利士 人轄制我們，你不知道嗎？你向我們做的是甚麼事呢？」他說：「他們向我怎樣做，我也要向他們怎樣做。」
JUDG|15|12|猶大 人對他說：「我們下來是要捆綁你，把你交在 非利士 人手中。」 參孫 說：「你們要向我起誓，你們自己不殺害我。」
JUDG|15|13|他們說：「我們絕不殺你，只把你捆綁，交在 非利士 人手中。」於是他們用兩條新繩綁住 參孫 ，把他從 以坦巖 帶上去。
JUDG|15|14|參孫 到了 利希 ， 非利士 人對著他喊叫。耶和華的靈大大感動 參孫 ，他手臂上的繩子就像著火的麻一樣，綁他的繩子從他手上脫落下來。
JUDG|15|15|他找到一塊未乾的驢腮骨，就伸手拾起來，用它殺了一千人。
JUDG|15|16|參孫 說： 「用驢腮骨， 一堆又一堆 ； 用驢腮骨， 我殺了一千人。」
JUDG|15|17|說完這話，就把那腮骨從手裏拋出去。因此，那地叫作 拉末‧利希 。
JUDG|15|18|參孫 非常口渴，就求告耶和華說：「你既藉僕人的手施行這麼大的拯救，現在我要渴死，落在未受割禮的人手中嗎？」
JUDG|15|19|上帝就使 利希 的窪地裂開，從中湧出水來。 參孫 喝了，精神恢復。因此那泉名叫 隱‧哈歌利 ，直到今日它仍在 利希 。
JUDG|15|20|在 非利士 人轄制的時候， 參孫 作 以色列 的士師二十年。
JUDG|16|1|參孫 到了 迦薩 ，在那裏看見一個妓女，就與她親近。
JUDG|16|2|有人告訴 迦薩 人說：「 參孫 到這裏來了！」他們就包圍起來，整夜在城門埋伏等著他。他們整夜靜悄悄地，說：「等到天一亮我們就殺他。」
JUDG|16|3|參孫 睡到半夜，在半夜起來，抓住城門的門扇和兩個門框，把它們和門閂一起拆下來，扛在肩上，抬到 希伯崙 前面的山頂上。
JUDG|16|4|這事以後， 參孫 在 梭烈谷 愛上了一個女子，名叫 大利拉 。
JUDG|16|5|非利士 人的領袖上去，到那女子那裏，對她說：「請你哄騙 參孫 ，探出他為何有這麼大的力氣，以及我們要用甚麼方法才能勝他，將他捆綁制伏。我們就每人給你一千一百塊銀子。」
JUDG|16|6|大利拉 對 參孫 說：「請你告訴我，你為何有這麼大的力氣，要用甚麼方法才能捆綁制伏你。」
JUDG|16|7|參孫 對她說：「若用七條未乾的新繩子捆綁我，我就像平常人一樣軟弱。」
JUDG|16|8|於是 非利士 人的領袖拿了七條未乾的新繩子來，交給她，她就用繩子捆綁 參孫 。
JUDG|16|9|當時，埋伏的人正在她的內室等著。她對 參孫 說：「 參孫 ， 非利士 人來捉你了！」 參孫 就掙斷繩子，繩子如遇到火的麻線斷裂一樣。這樣，人還是不知道他的力量從哪裏來。
JUDG|16|10|大利拉 對 參孫 說：「看哪，你欺騙我，對我說謊。現在請你告訴我，要用甚麼方法才能捆綁你。」
JUDG|16|11|參孫 對她說：「若用未曾用過的新繩子捆綁我，我就像平常人一樣軟弱。」
JUDG|16|12|大利拉 就用新繩子捆綁他，對他說：「 參孫 ， 非利士 人來捉你了！」當時，埋伏的人在內室等著。 參孫 掙斷手臂上的繩子，如掙斷一條線一樣。
JUDG|16|13|大利拉 對 參孫 說：「你到現在還是欺騙我，對我說謊。請你告訴我，要用甚麼方法才能捆綁你。」 參孫 對她說：「只要用織布的線將我頭上的七條髮綹編織起來就可以了」。
JUDG|16|14|於是 大利拉 用梭子將他的髮綹釘住，對他說：「 參孫 ， 非利士 人來捉你了！」 參孫 從睡中醒來，將織布機上的梭子和織布的線一齊都拔出來了。
JUDG|16|15|大利拉 對 參孫 說：「你既不與我同心，怎麼能說『我愛你』呢？你這三次欺騙我，不告訴我，你為甚麼有這麼大的力氣。」
JUDG|16|16|大利拉 天天用話催逼他，糾纏他，他就心裏煩得要死，
JUDG|16|17|終於把心中的一切都告訴她。 參孫 對她說：「從來沒有人用剃刀剃我的頭，因為我一出母胎就歸給上帝作拿細耳人。若有人剃了我的頭髮，我的力氣就會離開我，我就像平常人一樣軟弱。」
JUDG|16|18|大利拉 見他說出了心中的一切，就派人去召 非利士 人的領袖，說：「請再上來一次，因為他已經說出了心中的一切。」於是 非利士 人的領袖手裏拿著銀子，上到她那裏。
JUDG|16|19|大利拉 哄 參孫 睡在她的膝上，叫一個人來剃掉 參孫 頭上的七條髮綹。於是 大利拉 開始制伏 參孫 ，他的力氣就離開他了。
JUDG|16|20|大利拉 說：「 參孫 ， 非利士 人來捉你了！」 參孫 從睡中醒來，說：「我要像前幾次一樣脫身而去。」他卻不知道耶和華已經離開他了。
JUDG|16|21|非利士 人逮住他，挖了他的眼睛，帶他下到 迦薩 ，用銅鏈鎖住他，叫他在監獄裏推磨。
JUDG|16|22|然而他的頭髮被剃以後，又開始長起來了。
JUDG|16|23|非利士 人的領袖聚集，要向他們的神明 大袞 獻大祭，並且慶祝，說：「我們的神明把我們的仇敵 參孫 交在我們手中了。」
JUDG|16|24|眾人看見 參孫 ，就讚美他們的神明說：「我們的神明把那毀壞我們的地、殺害我們許多人的仇敵交在我們手中了。」
JUDG|16|25|他們心裏高興的時候，就說：「叫 參孫 來，逗我們歡樂。」於是他們把 參孫 從監獄裏提出來，在他們面前戲耍。他們叫他站在兩根柱子中間。
JUDG|16|26|參孫 對牽他手的童僕說：「讓我摸摸支撐這廟宇的柱子，我要靠一靠。」
JUDG|16|27|那時廟宇內充滿男女， 非利士 人的眾領袖也都在那裏，屋頂上約有三千男女觀看 參孫 逗他們歡樂。
JUDG|16|28|參孫 求告耶和華說：「主耶和華啊，求你眷念我。上帝啊，就這一次，求你賜給我力量，使我向 非利士 人報那挖我雙眼的仇。」
JUDG|16|29|參孫 抱住中間支撐廟宇的兩根柱子，左手抱一根，右手抱一根。
JUDG|16|30|然後他說：「讓我與 非利士 人一起死吧！」他盡力彎腰，廟宇就倒塌了，壓住領袖和廟宇內的眾人。這樣， 參孫 死的時候所殺的人比活著所殺的還多。
JUDG|16|31|他的兄弟和他父親的全家都下去收他的屍首，抬上去，葬在 瑣拉 和 以實陶 中間、他父親 瑪挪亞 的墳墓裏。 參孫 作 以色列 的士師二十年。
JUDG|17|1|以法蓮 山區有一個人，名叫 米迦 。
JUDG|17|2|他對母親說：「你的一千一百塊銀子被人拿走了，為此你發咒起誓，也說給我聽。看哪，銀子在我這裏，是我拿的。」他母親說：「願我兒蒙耶和華賜福！」
JUDG|17|3|米迦 把這一千一百塊銀子還他母親。他母親說：「我把這銀子分別為聖，親手獻給耶和華，為我兒子造一尊雕刻的像，以及一尊鑄成的像。現在我把銀子交給你。」
JUDG|17|4|米迦 把銀子還他母親，他母親把二百塊銀子交給銀匠，去造一尊雕刻的像，以及一尊鑄成的像，安置在 米迦 的房子裏。
JUDG|17|5|米迦 這個人有了神堂，又造了以弗得和家中的神像，派他的一個兒子作祭司。
JUDG|17|6|那時， 以色列 中沒有王，各人照自己眼中看為對的去做。
JUDG|17|7|猶大 的 伯利恆 有一個年輕人，是 猶大 族的人。他是 利未 人，寄居在那裏。
JUDG|17|8|這人離開 猶大 的 伯利恆城 ，要找一個可住的地方。他來到 以法蓮 山區 米迦 的家，還要往前走。
JUDG|17|9|米迦 對他說：「你從哪裏來？」他說：「我從 猶大 的 伯利恆 來。我是 利未 人，要找一個可住的地方。」
JUDG|17|10|米迦 說：「你就住在我這裏吧！我以你為父為祭司，每年給你十塊銀子和一套衣服，以及生活所需的食物。」 利未 人就來了。
JUDG|17|11|利未 人願意和這人同住；他待這年輕人如自己的兒子一樣。
JUDG|17|12|米迦 授這年輕的 利未 人祭司的職任，他就住在 米迦 的家裏。
JUDG|17|13|米迦 說：「現在我知道耶和華必恩待我，因為我有 利未 人作我的祭司。」
JUDG|18|1|那時， 以色列 中沒有王。 但 支派的人還在覓地居住，因為直到那日，他們還沒有在 以色列 支派中抽籤得地為業。
JUDG|18|2|但 人從 瑣拉 和 以實陶 派本族中的五個勇士，去窺探偵察那地，對他們說：「你們去偵察那地。」他們來到 以法蓮 山區 米迦 的家中，就在那裏住宿。
JUDG|18|3|他們臨近 米迦 的家，聽出那年輕的 利未 人的口音，就繞到那裏，對他說：「誰領你到這裏來？你在這裏做甚麼？你在這裏得了甚麼？」
JUDG|18|4|他對他們說：「 米迦 如此如此待我，他雇用我，我就作了他的祭司。」
JUDG|18|5|他們對他說：「請你求問上帝，使我們知道所走的道路是否通達。」
JUDG|18|6|祭司對他們說：「你們平平安安去吧，你們所行的道路是在耶和華面前的。」
JUDG|18|7|五人就走了，來到 拉億 ，見那裏的人安居，像 西頓 人的生活一樣安寧無慮，那地無人羞辱他們，無人奪取侵略。他們離 西頓 人很遠，與世無爭 。
JUDG|18|8|五人回到 瑣拉 和 以實陶 他們的弟兄那裏。他們的弟兄對他們說：「你們怎麼了？」
JUDG|18|9|他們說：「起來，我們上去攻打他們吧！我們已經窺探了那地，看哪，那地非常好。你們還要待在這裏嗎？不要再遲延了，立刻出發去得那地為業吧！
JUDG|18|10|你們去，必來到安居的百姓和兩邊遼闊的地。上帝已將那地方交在你們手中了；那裏不缺地上的任何東西。」
JUDG|18|11|於是 但 族的六百人，各帶兵器，從 瑣拉 和 以實陶 出發，
JUDG|18|12|上到 猶大 的 基列‧耶琳 ，在那裏安營。因此那地方名叫 瑪哈尼‧但 ，直到今日。看哪，它在 基列‧耶琳 的西邊。
JUDG|18|13|他們從那裏往 以法蓮 山區去，來到 米迦 的家。
JUDG|18|14|先前窺探 拉億 地的五個人對他們的弟兄說：「你們知道嗎？這些屋子裏有以弗得和家中的神像，以及一尊雕刻的像與一尊鑄成的像。現在你們要知道該怎麼做。」
JUDG|18|15|五人轉身，進入 米迦 的家，來到那年輕 利未 人的房間，向他問安。
JUDG|18|16|六百 但 人各帶兵器，站在門口。
JUDG|18|17|那窺探這地的五個人上前去，進入裏面，拿走雕刻的像、以弗得、家中的神像，以及鑄成的像。祭司和帶兵器的六百人一同站在門口。
JUDG|18|18|當五個人進入 米迦 的家，拿走雕刻的像、以弗得、家中的神像，以及鑄成的像，祭司對他們說：「你們做甚麼呢？」
JUDG|18|19|他們對他說：「不要作聲，用手摀口，跟我們去吧！我們必以你為父為祭司。你作一家的祭司好呢？還是作 以色列 一支派一族的祭司好呢？」
JUDG|18|20|祭司心裏歡喜，拿著以弗得和家中的神像，以及雕刻的像，跟這些百姓走了。
JUDG|18|21|他們轉身離開那裏，把孩子、牲畜、財物安排在前頭。
JUDG|18|22|他們離了 米迦 的家已遠， 米迦 家附近的鄰居被召來，追趕 但 人。
JUDG|18|23|他們呼叫 但 人， 但 人回頭對 米迦 說：「你召集這許多人來做甚麼呢？」
JUDG|18|24|米迦 說：「你們把我所造的神像，還有祭司，都帶走了，我還有甚麼呢？你怎麼還對我說『你在做甚麼』呢？」
JUDG|18|25|但 人對 米迦 說：「你不要讓我們再聽見你的聲音，恐怕這群惱怒成性的人會攻擊你們，你和你的全家就會喪命。」
JUDG|18|26|但 人仍走他們的路。 米迦 見他們的勢力比自己強，就轉身回家去了。
JUDG|18|27|但 人把 米迦 造的神像和他的祭司帶走，來到 拉億 安寧無慮的百姓那裏，用刀殺了他們，放火燒了那城。
JUDG|18|28|沒有人來搭救，因為這城離 西頓 很遠，他們又與世無爭；這城在靠近 伯‧利合 的平原。 但 人建造這城，在那裏居住，
JUDG|18|29|並照著他們祖先 以色列 之子 但 的名字，給這城起名叫 但 。原先這城名叫 拉億 。
JUDG|18|30|但 人為自己設立了那雕刻的像。 摩西 的孫子， 革舜 的兒子 約拿單 和他的子孫作 但 支派的祭司，直到那地遭擄掠的日子。
JUDG|18|31|上帝的家在 示羅 多少日子， 但 人為自己設立 米迦 所雕刻的像也在 但 多少日子。
JUDG|19|1|當 以色列 中沒有王的時候，有一個 利未 人寄居 以法蓮 山區的邊界，他娶了一個 猶大伯利恆 的女子為妾。
JUDG|19|2|這妾對丈夫生氣 ，離開丈夫，回到 猶大伯利恆 的父家，在那裏住了四個月。
JUDG|19|3|她的丈夫起來，帶著一個僕人、兩匹驢跟著她去，要用好話勸她回來。女子就帶丈夫進到父親家裏。女子的父親看見了他，就歡歡喜喜地迎接他。
JUDG|19|4|這岳父，就是女子的父親，留他住了三天。他們在那裏吃喝，住宿。
JUDG|19|5|第四日，他們清早起來， 利未 人起身要走，女子的父親對女婿說：「先吃點東西，加添心力，然後你們才走。」
JUDG|19|6|於是二人坐下，一同吃喝。女子的父親對那人說：「請你答應再住一夜，使你的心舒暢。」
JUDG|19|7|那人起身要走，他岳父挽留他，他就留下，在那裏又住了一夜。
JUDG|19|8|第五日，他清早起來要走，女子的父親說：「來，請加添心力，留到太陽偏西吧。」於是二人一同再吃。
JUDG|19|9|那人同他的妾和僕人起身要走，但他岳父，就是女子的父親，對他說：「看哪，太陽下山，天快晚了，你們再住一夜吧。看哪，太陽偏西了，就在這裏住宿，使你的心舒暢，明天你們一早起來上路，回你的帳棚去。」
JUDG|19|10|那人不願再住一夜，就備上兩匹驢，帶著他的妾起身走了，來到 耶布斯 的對面， 耶布斯 就是 耶路撒冷 。
JUDG|19|11|將近 耶布斯 的時候，太陽快下山了，僕人對主人說：「來吧，我們進這 耶布斯 人的城，在這裏住宿。」
JUDG|19|12|主人對他說：「我們不可進入外邦人的城，那不是 以色列 人的地方，我們越過這裏到 基比亞 去吧。」
JUDG|19|13|他又對僕人說：「來，讓我們到 基比亞 或 拉瑪 的一個地方住宿。」
JUDG|19|14|於是他們越過那裏往前走，將到 便雅憫 的 基比亞 的時候，太陽已經下山了。
JUDG|19|15|他們進入 基比亞 要在那裏住宿。他來坐在城裏的廣場上，但沒有人接待他們到家裏住宿。
JUDG|19|16|看哪，晚上有一個老人從田間做工回來。他是 以法蓮 山區的人，寄居在 基比亞 ；那地方的人是 便雅憫 人。
JUDG|19|17|老人舉目看見那過路的人在城裏的廣場上，就說：「你從哪裏來？要到哪裏去？」
JUDG|19|18|他對他說：「我們從 猶大 的 伯利恆 過來，要到 以法蓮 山區的邊界去。我是那裏的人，去了 猶大 的 伯利恆 ，現在要到耶和華的家去，卻沒有人接待我到他的家。
JUDG|19|19|其實我有飼料草料可以餵驢，我和你的使女，以及與我們在一起的僕人都有餅有酒，甚麼都不缺。」
JUDG|19|20|老人說：「願你平安！你所需用的我都會給你們，只是不可在廣場上過夜。」
JUDG|19|21|於是老人領他到家裏，餵上驢。他們洗了腳，就吃喝起來。
JUDG|19|22|他們心裏歡樂的時候，看哪，城中的無賴圍住房子，連連叩門，對老人，這家的主人說：「把那進你家的人帶出來，我們要與他交合。」
JUDG|19|23|這家的主人出來對他們說：「弟兄們，不要做這樣的惡事。這人既然進了我的家，你們就不要做這樣可恥的事。
JUDG|19|24|看哪，我有個女兒還是處女，還有這人的妾，我把她們領出來任由你們污辱她們，就照你們看為好的對待她們吧！但對這人你們不要做這樣可恥的事。」
JUDG|19|25|那些人卻不肯聽從他。那人抓住他的妾，把她拉出去給他們。他們強姦了她，整夜凌辱她，直到早晨，天色快亮才放她走。
JUDG|19|26|到了早晨，婦人回來，仆倒在留她主人住宿的那人的家門前，直到天亮。
JUDG|19|27|早晨，她的主人起來開了門，出去要上路。看哪，那婦人，他的妾倒在屋子門前，雙手搭在門檻上。
JUDG|19|28|他對婦人說：「起來，我們走吧！」婦人卻沒有回應。那人就將她馱在驢上，起身回自己的地方去了。
JUDG|19|29|到了家裏，他拿刀，抓住他的妾，把她的屍身切成十二塊，分送到 以色列 全境。
JUDG|19|30|凡看見的人都說：「自從 以色列 人離開 埃及 地上來，直到今日，像這樣的事還沒有發生過，也沒有見過。大家應當想一想，商討一下再說。」
JUDG|20|1|於是 以色列 眾人從 但 到 別是巴 ，以及從 基列 地出來，如同一人，聚集在 米斯巴 耶和華那裏。
JUDG|20|2|以色列 各支派中眾百姓的領袖，都站在上帝百姓的會中。拿刀的步兵共有四十萬。
JUDG|20|3|便雅憫 人聽見 以色列 人上了 米斯巴 。 以色列 人說：「請說，這惡事是怎麼發生的呢？」
JUDG|20|4|那 利未 人，就是被害婦人的丈夫，回答說：「我和我的妾來到 便雅憫 的 基比亞 住宿。
JUDG|20|5|基比亞 人夜間起來攻擊我，包圍我住的屋子。他們想要殺我，並把我的妾污辱致死。
JUDG|20|6|我把我的妾切成塊，分送到 以色列 得為業的全地，因為 基比亞 人在 以色列 中做了邪惡可恥的事。
JUDG|20|7|看哪，你們大家， 以色列 人哪，在此提出你們的建議和對策吧！」
JUDG|20|8|眾百姓都起來如同一人，說：「我們誰也不回自己的帳棚，誰也不回自己的家去！
JUDG|20|9|現在，我們要這樣對付 基比亞 ，照所抽的籤去攻打他們。
JUDG|20|10|我們要在 以色列 各支派中，一百人選十人，一千人選一百人，一萬人選一千人，為那到 便雅憫 的 迦巴 去的士兵運糧；因為 基比亞 在 以色列 中行了可恥的事。」
JUDG|20|11|於是 以色列 眾人彼此聯合如同一人，聚集攻擊那城。
JUDG|20|12|以色列 眾支派派人去，問 便雅憫 支派的各家說：「你們中間怎麼做了這樣的惡事呢？
JUDG|20|13|現在你們要把 基比亞 的那些無賴交出來，我們好處死他們，從 以色列 中除掉這惡。」 便雅憫 人卻不肯聽從他們弟兄 以色列 人的話。
JUDG|20|14|便雅憫 人從各城聚集到 基比亞 ，出來要與 以色列 人打仗。
JUDG|20|15|那日， 便雅憫 人從各城裏徵召了拿刀的士兵，共有二萬六千，另外還從 基比亞 居民中徵召七百個精兵。
JUDG|20|16|全軍中有特選的七百個精兵，都是慣用左手的，個個能用機弦甩石，毫髮不差。
JUDG|20|17|以色列 人，除了 便雅憫 之外，共徵召了四十萬拿刀的，個個都是戰士。
JUDG|20|18|以色列 人起來，上到 伯特利 去求問上帝說：「我們中間誰當首先上去與 便雅憫 人爭戰呢？」耶和華說：「 猶大 先上去。」
JUDG|20|19|以色列 人早晨起來，對著 基比亞 安營。
JUDG|20|20|以色列 人出來與 便雅憫 人打仗， 以色列 人在 基比亞 對著他們擺陣。
JUDG|20|21|便雅憫 人從 基比亞 出來，當日把 以色列 中二萬二千人殺倒在地。
JUDG|20|22|以色列 人的士兵鼓起勇氣，在第一日擺陣的地方又擺陣。
JUDG|20|23|因 以色列 人上去，在耶和華面前哀哭，直到晚上。他們求問耶和華說：「我可以再出兵與我弟兄 便雅憫 人打仗嗎？」耶和華說：「可以上去攻打他們。」
JUDG|20|24|第二日， 以色列 人就上前攻擊 便雅憫 人。
JUDG|20|25|便雅憫 人也在第二日從 基比亞 出來與他們交戰，又把 以色列 人一萬八千個拿刀的士兵殺倒在地。
JUDG|20|26|以色列 眾人和全體士兵上到 伯特利 ，坐在耶和華面前哭泣。那日，他們禁食直到晚上，又在耶和華面前獻燔祭和平安祭。
JUDG|20|27|以色列 人去求問耶和華；那時，上帝的約櫃在那裏。
JUDG|20|28|那時， 亞倫 的孫子， 以利亞撒 的兒子 非尼哈 侍立在約櫃前。他們說：「我可以再出去與我弟兄 便雅憫 人打仗嗎？還是停戰呢？」耶和華說：「你們可以上去，因為明日我必把他交在你手中。」
JUDG|20|29|以色列 在 基比亞 的四圍設下埋伏。
JUDG|20|30|第三日， 以色列 人又上去攻擊 便雅憫 人，在 基比亞 前擺陣，與前兩次一樣。
JUDG|20|31|便雅憫 人也出來迎敵，就被引誘出城外。在田間的兩條路上，一條通往 伯特利 ，一條通往 基比亞 ，他們像前兩次一樣，動手殺了約三十個 以色列 人。
JUDG|20|32|便雅憫 人說：「他們仍像以前一樣敗在我們面前。」但 以色列 人說：「讓我們逃跑，引誘他們離開城到路上來。」
JUDG|20|33|以色列 眾人都起來，在 巴力‧他瑪 擺陣， 以色列 的伏兵從 馬利‧迦巴 埋伏的地方衝上前去。
JUDG|20|34|全 以色列 中的一萬精兵來到 基比亞 前，戰爭十分激烈。 便雅憫 人卻不知道災禍臨近了。
JUDG|20|35|耶和華在 以色列 面前擊打 便雅憫 。那日， 以色列 人殲滅二萬五千一百個 便雅憫 人，都是拿刀的士兵。
JUDG|20|36|便雅憫 人看到自己戰敗了。 以色列 人因為信任在 基比亞 前所設的伏兵，就在 便雅憫 人面前假裝撤退。
JUDG|20|37|伏兵迅速闖進 基比亞 ；他們繼續前進，用刀殺死全城的人。
JUDG|20|38|以色列 人預先與伏兵約定在城內放火，以上騰的煙為信號。
JUDG|20|39|以色列 人從陣上撤退， 便雅憫 人動手殺死 以色列 人，約有三十個，就說：「他們仍像以前一樣敗在我們面前。」
JUDG|20|40|當煙如柱一般從城中上騰的時候， 便雅憫 人回頭，看哪，全城已經濃煙沖天了。
JUDG|20|41|以色列 人又轉身回來， 便雅憫 人就很驚惶，因為看見災禍臨到自己了。
JUDG|20|42|他們在 以色列 人面前轉身往曠野逃跑，戰況對他們不利，那從城裏出來的也去夾攻，殺滅他們。
JUDG|20|43|以色列 人圍攻 便雅憫 人，追趕他們，在他們歇腳之處，直到向日出方向的 基比亞 的對面，踐踏他們。
JUDG|20|44|便雅憫 人倒下的有一萬八千名，這些全都是勇士。
JUDG|20|45|其餘的人轉身往曠野逃跑，到 臨門巖 去。 以色列 人在路上殺了五千人，如拾穗一樣，緊追他們直到 基頓 ，又殺了二千人。
JUDG|20|46|那日 便雅憫 人倒下的有二萬五千名，這些全都是拿刀的勇士。
JUDG|20|47|有六百人轉身往曠野逃跑，到了 臨門巖 ，在 臨門巖 住了四個月。
JUDG|20|48|以色列 人又轉回去攻擊 便雅憫 人，凡經過的各城，其中的人和牲畜都用刀殺了，又放火燒了所經過的一切城鎮。
JUDG|21|1|以色列 人在 米斯巴 曾起誓說：「我們中誰都不把女兒嫁給 便雅憫 人。」
JUDG|21|2|以色列 人來到 伯特利 ，坐在那裏直到晚上，在上帝面前放聲大哭，
JUDG|21|3|說：「耶和華－ 以色列 的上帝啊，為何 以色列 中會發生這樣的事，使 以色列 今日缺了一個支派呢？」
JUDG|21|4|次日，百姓清早起來，在那裏築了一座壇，獻燔祭和平安祭。
JUDG|21|5|以色列 人說：「 以色列 各支派中，誰沒有同會眾一起上到耶和華那裏呢？」因為 以色列 人曾起重誓說：「凡不上 米斯巴 到耶和華那裏的，必被處死。」
JUDG|21|6|以色列 人憐憫他們的弟兄 便雅憫 ，說：「如今 以色列 中斷絕一個支派了。
JUDG|21|7|我們既然向耶和華起誓說，必不把我們的女兒嫁給 便雅憫 人，現在我們該怎麼辦，使他們剩下的人可以娶妻呢？」
JUDG|21|8|他們又說：「 以色列 支派中誰沒有上 米斯巴 到耶和華那裏呢？」看哪， 基列 的 雅比 沒有一人進營到會眾那裏，
JUDG|21|9|百姓被數點的時候，看哪， 基列 的 雅比 居民沒有一人在那裏。
JUDG|21|10|會眾就派一萬二千名大勇士，吩咐他們說：「你們去用刀把 基列 的 雅比 居民連婦女帶孩子都殺了。
JUDG|21|11|這是你們當做的事：要把所有男人和曾與男人同房共寢的女人全都殺了。」
JUDG|21|12|他們在 基列 的 雅比 居民中，找到四百個未曾與男人同房共寢的處女，就帶她們到 迦南 地的 示羅 營裏。
JUDG|21|13|全會眾派人到 臨門巖 的 便雅憫 人那裏，與他們講和。
JUDG|21|14|當時 便雅憫 人回來了， 以色列 人就把所留下， 基列 的 雅比 活著的女子嫁給他們，可是還是不夠。
JUDG|21|15|百姓憐憫 便雅憫 人，因為耶和華使 以色列 支派中有一個缺口。
JUDG|21|16|會眾中的長老說：「 便雅憫 中的女子既然都除滅了，我們該怎麼辦，使剩下的人可以娶妻呢？」
JUDG|21|17|他們又說：「 便雅憫 逃脫的人應當有地業，免得 以色列 中的一個支派被塗去。
JUDG|21|18|只是我們不能把自己的女兒嫁給他們。」因為 以色列 人曾起誓說：「把女兒嫁給 便雅憫 人的必受詛咒。」
JUDG|21|19|他們又說：「看哪，一年一度耶和華的節期正在 示羅 舉行。」 示羅 位於 利波拿 的南邊， 伯特利 的北邊，從 伯特利 往 示劍 大路的東邊。
JUDG|21|20|他們吩咐 便雅憫 人說：「你們去，躲在葡萄園中，
JUDG|21|21|觀看；看哪，若 示羅 的女子出來跳舞，你們就從葡萄園出來，各人從 示羅 的女子中搶一個為妻，然後到 便雅憫 地去。
JUDG|21|22|他們的父親或兄弟若來與我們爭論，我們就對他們說：『請看我們的情面恩待這些人吧！因為我們在戰爭的時候沒有給他們任何人留下女子為妻。這次也不是你們給他們的，若是你們給的，就算有罪了。』」
JUDG|21|23|於是 便雅憫 人就照樣做了，按照他們的人數，把從跳舞女子中搶來的娶為妻子，帶回自己的地業，重建城鎮，居住在其中。
JUDG|21|24|那時 以色列 人離開那裏，各自回到自己的支派、宗族；他們從那裏起行，各自回到自己的地業去了。
JUDG|21|25|那時， 以色列 中沒有王，各人照自己眼中看為對的去做。
