REV|1|1|Откровение Иисуса Христа, которое дал Ему Бог, чтобы показать рабам Своим, чему надлежит быть вскоре. И Он показал, послав [оное] через Ангела Своего рабу Своему Иоанну,
REV|1|2|который свидетельствовал слово Божие и свидетельство Иисуса Христа и что он видел.
REV|1|3|Блажен читающий и слушающие слова пророчества сего и соблюдающие написанное в нем; ибо время близко.
REV|1|4|Иоанн семи церквам, находящимся в Асии: благодать вам и мир от Того, Который есть и был и грядет, и от семи духов, находящихся перед престолом Его,
REV|1|5|и от Иисуса Христа, Который есть свидетель верный, первенец из мертвых и владыка царей земных. Ему, возлюбившему нас и омывшему нас от грехов наших Кровию Своею
REV|1|6|и соделавшему нас царями и священниками Богу и Отцу Своему, слава и держава во веки веков, аминь.
REV|1|7|Се, грядет с облаками, и узрит Его всякое око и те, которые пронзили Его; и возрыдают пред Ним все племена земные. Ей, аминь.
REV|1|8|Я есмь Альфа и Омега, начало и конец, говорит Господь, Который есть и был и грядет, Вседержитель.
REV|1|9|Я, Иоанн, брат ваш и соучастник в скорби и в царствии и в терпении Иисуса Христа, был на острове, называемом Патмос, за слово Божие и за свидетельство Иисуса Христа.
REV|1|10|Я был в духе в день воскресный, и слышал позади себя громкий голос, как бы трубный, который говорил: Я есмь Альфа и Омега, Первый и Последний;
REV|1|11|то, что видишь, напиши в книгу и пошли церквам, находящимся в Асии: в Ефес, и в Смирну, и в Пергам, и в Фиатиру, и в Сардис, и в Филадельфию, и в Лаодикию.
REV|1|12|Я обратился, чтобы увидеть, чей голос, говоривший со мною; и обратившись, увидел семь золотых светильников
REV|1|13|и, посреди семи светильников, подобного Сыну Человеческому, облеченного в подир и по персям опоясанного золотым поясом:
REV|1|14|глава Его и волосы белы, как белая волна, как снег; и очи Его, как пламень огненный;
REV|1|15|и ноги Его подобны халколивану, как раскаленные в печи, и голос Его, как шум вод многих.
REV|1|16|Он держал в деснице Своей семь звезд, и из уст Его выходил острый с обеих сторон меч; и лице Его, как солнце, сияющее в силе своей.
REV|1|17|И когда я увидел Его, то пал к ногам Его, как мертвый. И Он положил на меня десницу Свою и сказал мне: не бойся; Я есмь Первый и Последний,
REV|1|18|и живый; и был мертв, и се, жив во веки веков, аминь; и имею ключи ада и смерти.
REV|1|19|Итак напиши, что ты видел, и что есть, и что будет после сего.
REV|1|20|Тайна семи звезд, которые ты видел в деснице Моей, и семи золотых светильников [есть сия]: семь звезд суть Ангелы семи церквей; а семь светильников, которые ты видел, суть семь церквей.
REV|2|1|Ангелу Ефесской церкви напиши: так говорит Держащий семь звезд в деснице Своей, Ходящий посреди семи золотых светильников:
REV|2|2|знаю дела твои, и труд твой, и терпение твое, и то, что ты не можешь сносить развратных, и испытал тех, которые называют себя апостолами, а они не таковы, и нашел, что они лжецы;
REV|2|3|ты много переносил и имеешь терпение, и для имени Моего трудился и не изнемогал.
REV|2|4|Но имею против тебя то, что ты оставил первую любовь твою.
REV|2|5|Итак вспомни, откуда ты ниспал, и покайся, и твори прежние дела; а если не так, скоро приду к тебе, и сдвину светильник твой с места его, если не покаешься.
REV|2|6|Впрочем то в тебе [хорошо], что ты ненавидишь дела Николаитов, которые и Я ненавижу.
REV|2|7|Имеющий ухо да слышит, что Дух говорит церквам: побеждающему дам вкушать от древа жизни, которое посреди рая Божия.
REV|2|8|И Ангелу Смирнской церкви напиши: так говорит Первый и Последний, Который был мертв, и се, жив:
REV|2|9|Знаю твои дела, и скорбь, и нищету (впрочем ты богат), и злословие от тех, которые говорят о себе, что они Иудеи, а они не таковы, но сборище сатанинское.
REV|2|10|Не бойся ничего, что тебе надобно будет претерпеть. Вот, диавол будет ввергать из среды вас в темницу, чтобы искусить вас, и будете иметь скорбь дней десять. Будь верен до смерти, и дам тебе венец жизни.
REV|2|11|Имеющий ухо (слышать) да слышит, что Дух говорит церквам: побеждающий не потерпит вреда от второй смерти.
REV|2|12|И Ангелу Пергамской церкви напиши: так говорит Имеющий острый с обеих сторон меч:
REV|2|13|знаю твои дела, и что ты живешь там, где престол сатаны, и что содержишь имя Мое, и не отрекся от веры Моей даже в те дни, в которые у вас, где живет сатана, умерщвлен верный свидетель Мой Антипа.
REV|2|14|Но имею немного против тебя, потому что есть у тебя там держащиеся учения Валаама, который научил Валака ввести в соблазн сынов Израилевых, чтобы они ели идоложертвенное и любодействовали.
REV|2|15|Так и у тебя есть держащиеся учения Николаитов, которое Я ненавижу.
REV|2|16|Покайся; а если не так, скоро приду к тебе и сражусь с ними мечом уст Моих.
REV|2|17|Имеющий ухо (слышать) да слышит, что Дух говорит церквам: побеждающему дам вкушать сокровенную манну, и дам ему белый камень и на камне написанное новое имя, которого никто не знает, кроме того, кто получает.
REV|2|18|И Ангелу Фиатирской церкви напиши: так говорит Сын Божий, у Которого очи, как пламень огненный, и ноги подобны халколивану:
REV|2|19|знаю твои дела и любовь, и служение, и веру, и терпение твое, и то, что последние дела твои больше первых.
REV|2|20|Но имею немного против тебя, потому что ты попускаешь жене Иезавели, называющей себя пророчицею, учить и вводить в заблуждение рабов Моих, любодействовать и есть идоложертвенное.
REV|2|21|Я дал ей время покаяться в любодеянии ее, но она не покаялась.
REV|2|22|Вот, Я повергаю ее на одр и любодействующих с нею в великую скорбь, если не покаются в делах своих.
REV|2|23|И детей ее поражу смертью, и уразумеют все церкви, что Я есмь испытующий сердца и внутренности; и воздам каждому из вас по делам вашим.
REV|2|24|Вам же и прочим, находящимся в Фиатире, которые не держат сего учения и которые не знают так называемых глубин сатанинских, сказываю, что не наложу на вас иного бремени;
REV|2|25|только то, что имеете, держите, пока приду.
REV|2|26|Кто побеждает и соблюдает дела Мои до конца, тому дам власть над язычниками,
REV|2|27|и будет пасти их жезлом железным; как сосуды глиняные, они сокрушатся, как и Я получил [власть] от Отца Моего;
REV|2|28|и дам ему звезду утреннюю.
REV|2|29|Имеющий ухо (слышать) да слышит, что Дух говорит церквам.
REV|3|1|И Ангелу Сардийской церкви напиши: так говорит Имеющий семь духов Божиих и семь звезд: знаю твои дела; ты носишь имя, будто жив, но ты мертв.
REV|3|2|Бодрствуй и утверждай прочее близкое к смерти; ибо Я не нахожу, чтобы дела твои были совершенны пред Богом Моим.
REV|3|3|Вспомни, что ты принял и слышал, и храни и покайся. Если же не будешь бодрствовать, то Я найду на тебя, как тать, и ты не узнаешь, в который час найду на тебя.
REV|3|4|Впрочем у тебя в Сардисе есть несколько человек, которые не осквернили одежд своих, и будут ходить со Мною в белых [одеждах], ибо они достойны.
REV|3|5|Побеждающий облечется в белые одежды; и не изглажу имени его из книги жизни, и исповедаю имя его пред Отцем Моим и пред Ангелами Его.
REV|3|6|Имеющий ухо да слышит, что Дух говорит церквам.
REV|3|7|И Ангелу Филадельфийской церкви напиши: так говорит Святый, Истинный, имеющий ключ Давидов, Который отворяет – и никто не затворит, затворяет – и никто не отворит:
REV|3|8|знаю твои дела; вот, Я отворил перед тобою дверь, и никто не может затворить ее; ты не много имеешь силы, и сохранил слово Мое, и не отрекся имени Моего.
REV|3|9|Вот, Я сделаю, что из сатанинского сборища, из тех, которые говорят о себе, что они Иудеи, но не суть таковы, а лгут, – вот, Я сделаю то, что они придут и поклонятся пред ногами твоими, и познают, что Я возлюбил тебя.
REV|3|10|И как ты сохранил слово терпения Моего, то и Я сохраню тебя от годины искушения, которая придет на всю вселенную, чтобы испытать живущих на земле.
REV|3|11|Се, гряду скоро; держи, что имеешь, дабы кто не восхитил венца твоего.
REV|3|12|Побеждающего сделаю столпом в храме Бога Моего, и он уже не выйдет вон; и напишу на нем имя Бога Моего и имя града Бога Моего, нового Иерусалима, нисходящего с неба от Бога Моего, и имя Мое новое.
REV|3|13|Имеющий ухо да слышит, что Дух говорит церквам.
REV|3|14|И Ангелу Лаодикийской церкви напиши: так говорит Аминь, свидетель верный и истинный, начало создания Божия:
REV|3|15|знаю твои дела; ты ни холоден, ни горяч; о, если бы ты был холоден, или горяч!
REV|3|16|Но, как ты тепл, а не горяч и не холоден, то извергну тебя из уст Моих.
REV|3|17|Ибо ты говоришь: "я богат, разбогател и ни в чем не имею нужды"; а не знаешь, что ты несчастен, и жалок, и нищ, и слеп, и наг.
REV|3|18|Советую тебе купить у Меня золото, огнем очищенное, чтобы тебе обогатиться, и белую одежду, чтобы одеться и чтобы не видна была срамота наготы твоей, и глазною мазью помажь глаза твои, чтобы видеть.
REV|3|19|Кого Я люблю, тех обличаю и наказываю. Итак будь ревностен и покайся.
REV|3|20|Се, стою у двери и стучу: если кто услышит голос Мой и отворит дверь, войду к нему, и буду вечерять с ним, и он со Мною.
REV|3|21|Побеждающему дам сесть со Мною на престоле Моем, как и Я победил и сел с Отцем Моим на престоле Его.
REV|3|22|Имеющий ухо да слышит, что Дух говорит церквам.
REV|4|1|После сего я взглянул, и вот, дверь отверста на небе, и прежний голос, который я слышал как бы звук трубы, говоривший со мною, сказал: взойди сюда, и покажу тебе, чему надлежит быть после сего.
REV|4|2|И тотчас я был в духе; и вот, престол стоял на небе, и на престоле был Сидящий;
REV|4|3|и Сей Сидящий видом был подобен камню яспису и сардису; и радуга вокруг престола, видом подобная смарагду.
REV|4|4|И вокруг престола двадцать четыре престола; а на престолах видел я сидевших двадцать четыре старца, которые облечены были в белые одежды и имели на головах своих золотые венцы.
REV|4|5|И от престола исходили молнии и громы и гласы, и семь светильников огненных горели перед престолом, которые суть семь духов Божиих;
REV|4|6|и перед престолом море стеклянное, подобное кристаллу; и посреди престола и вокруг престола четыре животных, исполненных очей спереди и сзади.
REV|4|7|И первое животное было подобно льву, и второе животное подобно тельцу, и третье животное имело лице, как человек, и четвертое животное подобно орлу летящему.
REV|4|8|И каждое из четырех животных имело по шести крыл вокруг, а внутри они исполнены очей; и ни днем, ни ночью не имеют покоя, взывая: свят, свят, свят Господь Бог Вседержитель, Который был, есть и грядет.
REV|4|9|И когда животные воздают славу и честь и благодарение Сидящему на престоле, Живущему во веки веков,
REV|4|10|тогда двадцать четыре старца падают пред Сидящим на престоле, и поклоняются Живущему во веки веков, и полагают венцы свои перед престолом, говоря:
REV|4|11|достоин Ты, Господи, приять славу и честь и силу: ибо Ты сотворил все, и [все] по Твоей воле существует и сотворено.
REV|5|1|И видел я в деснице у Сидящего на престоле книгу, написанную внутри и отвне, запечатанную семью печатями.
REV|5|2|И видел я Ангела сильного, провозглашающего громким голосом: кто достоин раскрыть сию книгу и снять печати ее?
REV|5|3|И никто не мог, ни на небе, ни на земле, ни под землею, раскрыть сию книгу, ни посмотреть в нее.
REV|5|4|И я много плакал о том, что никого не нашлось достойного раскрыть и читать сию книгу, и даже посмотреть в нее.
REV|5|5|И один из старцев сказал мне: не плачь; вот, лев от колена Иудина, корень Давидов, победил, [и может] раскрыть сию книгу и снять семь печатей ее.
REV|5|6|И я взглянул, и вот, посреди престола и четырех животных и посреди старцев стоял Агнец как бы закланный, имеющий семь рогов и семь очей, которые суть семь духов Божиих, посланных во всю землю.
REV|5|7|И Он пришел и взял книгу из десницы Сидящего на престоле.
REV|5|8|И когда он взял книгу, тогда четыре животных и двадцать четыре старца пали пред Агнцем, имея каждый гусли и золотые чаши, полные фимиама, которые суть молитвы святых.
REV|5|9|И поют новую песнь, говоря: достоин Ты взять книгу и снять с нее печати, ибо Ты был заклан, и Кровию Своею искупил нас Богу из всякого колена и языка, и народа и племени,
REV|5|10|и соделал нас царями и священниками Богу нашему; и мы будем царствовать на земле.
REV|5|11|И я видел, и слышал голос многих Ангелов вокруг престола и животных и старцев, и число их было тьмы тем и тысячи тысяч,
REV|5|12|которые говорили громким голосом: достоин Агнец закланный принять силу и богатство, и премудрость и крепость, и честь и славу и благословение.
REV|5|13|И всякое создание, находящееся на небе и на земле, и под землею, и на море, и все, что в них, слышал я, говорило: Сидящему на престоле и Агнцу благословение и честь, и слава и держава во веки веков.
REV|5|14|И четыре животных говорили: аминь. И двадцать четыре старца пали и поклонились Живущему во веки веков.
REV|6|1|И я видел, что Агнец снял первую из семи печатей, и я услышал одно из четырех животных, говорящее как бы громовым голосом: иди и смотри.
REV|6|2|Я взглянул, и вот, конь белый, и на нем всадник, имеющий лук, и дан был ему венец; и вышел он [как] победоносный, и чтобы победить.
REV|6|3|И когда он снял вторую печать, я слышал второе животное, говорящее: иди и смотри.
REV|6|4|И вышел другой конь, рыжий; и сидящему на нем дано взять мир с земли, и чтобы убивали друг друга; и дан ему большой меч.
REV|6|5|И когда Он снял третью печать, я слышал третье животное, говорящее: иди и смотри. Я взглянул, и вот, конь вороной, и на нем всадник, имеющий меру в руке своей.
REV|6|6|И слышал я голос посреди четырех животных, говорящий: хиникс пшеницы за динарий, и три хиникса ячменя за динарий; елея же и вина не повреждай.
REV|6|7|И когда Он снял четвертую печать, я слышал голос четвертого животного, говорящий: иди и смотри.
REV|6|8|И я взглянул, и вот, конь бледный, и на нем всадник, которому имя "смерть"; и ад следовал за ним; и дана ему власть над четвертою частью земли – умерщвлять мечом и голодом, и мором и зверями земными.
REV|6|9|И когда Он снял пятую печать, я увидел под жертвенником души убиенных за слово Божие и за свидетельство, которое они имели.
REV|6|10|И возопили они громким голосом, говоря: доколе, Владыка Святый и Истинный, не судишь и не мстишь живущим на земле за кровь нашу?
REV|6|11|И даны были каждому из них одежды белые, и сказано им, чтобы они успокоились еще на малое время, пока и сотрудники их и братья их, которые будут убиты, как и они, дополнят число.
REV|6|12|И когда Он снял шестую печать, я взглянул, и вот, произошло великое землетрясение, и солнце стало мрачно как власяница, и луна сделалась как кровь.
REV|6|13|И звезды небесные пали на землю, как смоковница, потрясаемая сильным ветром, роняет незрелые смоквы свои.
REV|6|14|И небо скрылось, свившись как свиток; и всякая гора и остров двинулись с мест своих.
REV|6|15|И цари земные, и вельможи, и богатые, и тысяченачальники, и сильные, и всякий раб, и всякий свободный скрылись в пещеры и в ущелья гор,
REV|6|16|и говорят горам и камням: падите на нас и сокройте нас от лица Сидящего на престоле и от гнева Агнца;
REV|6|17|ибо пришел великий день гнева Его, и кто может устоять?
REV|7|1|И после сего видел я четырех Ангелов, стоящих на четырех углах земли, держащих четыре ветра земли, чтобы не дул ветер ни на землю, ни на море, ни на какое дерево.
REV|7|2|И видел я иного Ангела, восходящего от востока солнца и имеющего печать Бога живаго. И воскликнул он громким голосом к четырем Ангелам, которым дано вредить земле и морю, говоря:
REV|7|3|не делайте вреда ни земле, ни морю, ни деревам, доколе не положим печати на челах рабов Бога нашего.
REV|7|4|И я слышал число запечатленных: запечатленных было сто сорок четыре тысячи из всех колен сынов Израилевых.
REV|7|5|Из колена Иудина запечатлено двенадцать тысяч; из колена Рувимова запечатлено двенадцать тысяч; из колена Гадова запечатлено двенадцать тысяч;
REV|7|6|из колена Асирова запечатлено двенадцать тысяч; из колена Неффалимова запечатлено двенадцать тысяч; из колена Манассиина запечатлено двенадцать тысяч;
REV|7|7|из колена Симеонова запечатлено двенадцать тысяч; из колена Левиина запечатлено двенадцать тысяч; из колена Иссахарова запечатлено двенадцать тысяч;
REV|7|8|из колена Завулонова запечатлено двенадцать тысяч; из колена Иосифова запечатлено двенадцать тысяч; из колена Вениаминова запечатлено двенадцать тысяч.
REV|7|9|После сего взглянул я, и вот, великое множество людей, которого никто не мог перечесть, из всех племен и колен, и народов и языков, стояло пред престолом и пред Агнцем в белых одеждах и с пальмовыми ветвями в руках своих.
REV|7|10|И восклицали громким голосом, говоря: спасение Богу нашему, сидящему на престоле, и Агнцу!
REV|7|11|И все Ангелы стояли вокруг престола и старцев и четырех животных, и пали перед престолом на лица свои, и поклонились Богу,
REV|7|12|говоря: аминь! благословение и слава, и премудрость и благодарение, и честь и сила и крепость Богу нашему во веки веков! Аминь.
REV|7|13|И, начав речь, один из старцев спросил меня: сии облеченные в белые одежды кто, и откуда пришли?
REV|7|14|Я сказал ему: ты знаешь, господин. И он сказал мне: это те, которые пришли от великой скорби; они омыли одежды свои и убелили одежды свои Кровию Агнца.
REV|7|15|За это они пребывают [ныне] перед престолом Бога и служат Ему день и ночь в храме Его, и Сидящий на престоле будет обитать в них.
REV|7|16|Они не будут уже ни алкать, ни жаждать, и не будет палить их солнце и никакой зной:
REV|7|17|ибо Агнец, Который среди престола, будет пасти их и водить их на живые источники вод; и отрет Бог всякую слезу с очей их.
REV|8|1|И когда Он снял седьмую печать, сделалось безмолвие на небе, как бы на полчаса.
REV|8|2|И я видел семь Ангелов, которые стояли пред Богом; и дано им семь труб.
REV|8|3|И пришел иной Ангел, и стал перед жертвенником, держа золотую кадильницу; и дано было ему множество фимиама, чтобы он с молитвами всех святых возложил его на золотой жертвенник, который перед престолом.
REV|8|4|И вознесся дым фимиама с молитвами святых от руки Ангела пред Бога.
REV|8|5|И взял Ангел кадильницу, и наполнил ее огнем с жертвенника, и поверг на землю: и произошли голоса и громы, и молнии и землетрясение.
REV|8|6|И семь Ангелов, имеющие семь труб, приготовились трубить.
REV|8|7|Первый Ангел вострубил, и сделались град и огонь, смешанные с кровью, и пали на землю; и третья часть дерев сгорела, и вся трава зеленая сгорела.
REV|8|8|Второй Ангел вострубил, и как бы большая гора, пылающая огнем, низверглась в море; и третья часть моря сделалась кровью,
REV|8|9|и умерла третья часть одушевленных тварей, живущих в море, и третья часть судов погибла.
REV|8|10|Третий ангел вострубил, и упала с неба большая звезда, горящая подобно светильнику, и пала на третью часть рек и на источники вод.
REV|8|11|Имя сей звезде "полынь"; и третья часть вод сделалась полынью, и многие из людей умерли от вод, потому что они стали горьки.
REV|8|12|Четвертый Ангел вострубил, и поражена была третья часть солнца и третья часть луны и третья часть звезд, так что затмилась третья часть их, и третья часть дня не светла была – так, как и ночи.
REV|8|13|И видел я и слышал одного Ангела, летящего посреди неба и говорящего громким голосом: горе, горе, горе живущим на земле от остальных трубных голосов трех Ангелов, которые будут трубить!
REV|9|1|Пятый Ангел вострубил, и я увидел звезду, падшую с неба на землю, и дан был ей ключ от кладязя бездны.
REV|9|2|Она отворила кладязь бездны, и вышел дым из кладязя, как дым из большой печи; и помрачилось солнце и воздух от дыма из кладязя.
REV|9|3|И из дыма вышла саранча на землю, и дана была ей власть, какую имеют земные скорпионы.
REV|9|4|И сказано было ей, чтобы не делала вреда траве земной, и никакой зелени, и никакому дереву, а только одним людям, которые не имеют печати Божией на челах своих.
REV|9|5|И дано ей не убивать их, а только мучить пять месяцев; и мучение от нее подобно мучению от скорпиона, когда ужалит человека.
REV|9|6|В те дни люди будут искать смерти, но не найдут ее; пожелают умереть, но смерть убежит от них.
REV|9|7|По виду своему саранча была подобна коням, приготовленным на войну; и на головах у ней как бы венцы, похожие на золотые, лица же ее – как лица человеческие;
REV|9|8|и волосы у ней – как волосы у женщин, а зубы у ней были, как у львов.
REV|9|9|На ней были брони, как бы брони железные, а шум от крыльев ее – как стук от колесниц, когда множество коней бежит на войну;
REV|9|10|у ней были хвосты, как у скорпионов, и в хвостах ее были жала; власть же ее была – вредить людям пять месяцев.
REV|9|11|Царем над собою она имела ангела бездны; имя ему по–еврейски Аваддон, а по–гречески Аполлион.
REV|9|12|Одно горе прошло; вот, идут за ним еще два горя.
REV|9|13|Шестой Ангел вострубил, и я услышал один голос от четырех рогов золотого жертвенника, стоящего пред Богом,
REV|9|14|говоривший шестому Ангелу, имевшему трубу: освободи четырех Ангелов, связанных при великой реке Евфрате.
REV|9|15|И освобождены были четыре Ангела, приготовленные на час и день, и месяц и год, для того, чтобы умертвить третью часть людей.
REV|9|16|Число конного войска было две тьмы тем; и я слышал число его.
REV|9|17|Так видел я в видении коней и на них всадников, которые имели на себе брони огненные, гиацинтовые и серные; головы у коней – как головы у львов, и изо рта их выходил огонь, дым и сера.
REV|9|18|От этих трех язв, от огня, дыма и серы, выходящих изо рта их, умерла третья часть людей;
REV|9|19|ибо сила коней заключалась во рту их и в хвостах их; а хвосты их были подобны змеям, и имели головы, и ими они вредили.
REV|9|20|Прочие же люди, которые не умерли от этих язв, не раскаялись в делах рук своих, так чтобы не поклоняться бесам и золотым, серебряным, медным, каменным и деревянным идолам, которые не могут ни видеть, ни слышать, ни ходить.
REV|9|21|И не раскаялись они в убийствах своих, ни в чародействах своих, ни в блудодеянии своем, ни в воровстве своем.
REV|10|1|И видел я другого Ангела сильного, сходящего с неба, облеченного облаком; над головою его была радуга, и лице его как солнце, и ноги его как столпы огненные,
REV|10|2|в руке у него была книжка раскрытая. И поставил он правую ногу свою на море, а левую на землю,
REV|10|3|и воскликнул громким голосом, как рыкает лев; и когда он воскликнул, тогда семь громов проговорили голосами своими.
REV|10|4|И когда семь громов проговорили голосами своими, я хотел было писать; но услышал голос с неба, говорящий мне: скрой, что говорили семь громов, и не пиши сего.
REV|10|5|И Ангел, которого я видел стоящим на море и на земле, поднял руку свою к небу
REV|10|6|и клялся Живущим во веки веков, Который сотворил небо и все, что на нем, землю и все, что на ней, и море и все, что в нем, что времени уже не будет;
REV|10|7|но в те дни, когда возгласит седьмой Ангел, когда он вострубит, совершится тайна Божия, как Он благовествовал рабам Своим пророкам.
REV|10|8|И голос, который я слышал с неба, опять стал говорить со мною, и сказал: пойди, возьми раскрытую книжку из руки Ангела, стоящего на море и на земле.
REV|10|9|И я пошел к Ангелу, и сказал ему: дай мне книжку. Он сказал мне: возьми и съешь ее; она будет горька во чреве твоем, но в устах твоих будет сладка, как мед.
REV|10|10|И взял я книжку из руки Ангела, и съел ее; и она в устах моих была сладка, как мед; когда же съел ее, то горько стало во чреве моем.
REV|10|11|И сказал он мне: тебе надлежит опять пророчествовать о народах и племенах, и языках и царях многих.
REV|11|1|И дана мне трость, подобная жезлу, и сказано: встань и измерь храм Божий и жертвенник, и поклоняющихся в нем.
REV|11|2|А внешний двор храма исключи и не измеряй его, ибо он дан язычникам: они будут попирать святый город сорок два месяца.
REV|11|3|И дам двум свидетелям Моим, и они будут пророчествовать тысячу двести шестьдесят дней, будучи облечены во вретище.
REV|11|4|Это суть две маслины и два светильника, стоящие пред Богом земли.
REV|11|5|И если кто захочет их обидеть, то огонь выйдет из уст их и пожрет врагов их; если кто захочет их обидеть, тому надлежит быть убиту.
REV|11|6|Они имеют власть затворить небо, чтобы не шел дождь на землю во дни пророчествования их, и имеют власть над водами, превращать их в кровь, и поражать землю всякою язвою, когда только захотят.
REV|11|7|И когда кончат они свидетельство свое, зверь, выходящий из бездны, сразится с ними, и победит их, и убьет их,
REV|11|8|и трупы их оставит на улице великого города, который духовно называется Содом и Египет, где и Господь наш распят.
REV|11|9|И [многие] из народов и колен, и языков и племен будут смотреть на трупы их три дня с половиною, и не позволят положить трупы их во гробы.
REV|11|10|И живущие на земле будут радоваться сему и веселиться, и пошлют дары друг другу, потому что два пророка сии мучили живущих на земле.
REV|11|11|Но после трех дней с половиною вошел в них дух жизни от Бога, и они оба стали на ноги свои; и великий страх напал на тех, которые смотрели на них.
REV|11|12|И услышали они с неба громкий голос, говоривший им: взойдите сюда. И они взошли на небо на облаке; и смотрели на них враги их.
REV|11|13|И в тот же час произошло великое землетрясение, и десятая часть города пала, и погибло при землетрясении семь тысяч имен человеческих; и прочие объяты были страхом и воздали славу Богу небесному.
REV|11|14|Второе горе прошло; вот, идет скоро третье горе.
REV|11|15|И седьмой Ангел вострубил, и раздались на небе громкие голоса, говорящие: царство мира соделалось [царством] Господа нашего и Христа Его, и будет царствовать во веки веков.
REV|11|16|И двадцать четыре старца, сидящие пред Богом на престолах своих, пали на лица свои и поклонились Богу,
REV|11|17|говоря: благодарим Тебя, Господи Боже Вседержитель, Который еси и был и грядешь, что ты приял силу Твою великую и воцарился.
REV|11|18|И рассвирепели язычники; и пришел гнев Твой и время судить мертвых и дать возмездие рабам Твоим, пророкам и святым и боящимся имени Твоего, малым и великим, и погубить губивших землю.
REV|11|19|И отверзся храм Божий на небе, и явился ковчег завета Его в храме Его; и произошли молнии и голоса, и громы и землетрясение и великий град.
REV|12|1|И явилось на небе великое знамение: жена, облеченная в солнце; под ногами ее луна, и на главе ее венец из двенадцати звезд.
REV|12|2|Она имела во чреве, и кричала от болей и мук рождения.
REV|12|3|И другое знамение явилось на небе: вот, большой красный дракон с семью головами и десятью рогами, и на головах его семь диадим.
REV|12|4|Хвост его увлек с неба третью часть звезд и поверг их на землю. Дракон сей стал перед женою, которой надлежало родить, дабы, когда она родит, пожрать ее младенца.
REV|12|5|И родила она младенца мужеского пола, которому надлежит пасти все народы жезлом железным; и восхищено было дитя ее к Богу и престолу Его.
REV|12|6|А жена убежала в пустыню, где приготовлено было для нее место от Бога, чтобы питали ее там тысячу двести шестьдесят дней.
REV|12|7|И произошла на небе война: Михаил и Ангелы его воевали против дракона, и дракон и ангелы его воевали [против них],
REV|12|8|но не устояли, и не нашлось уже для них места на небе.
REV|12|9|И низвержен был великий дракон, древний змий, называемый диаволом и сатаною, обольщающий всю вселенную, низвержен на землю, и ангелы его низвержены с ним.
REV|12|10|И услышал я громкий голос, говорящий на небе: ныне настало спасение и сила и царство Бога нашего и власть Христа Его, потому что низвержен клеветник братий наших, клеветавший на них пред Богом нашим день и ночь.
REV|12|11|Они победили его кровию Агнца и словом свидетельства своего, и не возлюбили души своей даже до смерти.
REV|12|12|Итак веселитесь, небеса и обитающие на них! Горе живущим на земле и на море! потому что к вам сошел диавол в сильной ярости, зная, что немного ему остается времени.
REV|12|13|Когда же дракон увидел, что низвержен на землю, начал преследовать жену, которая родила младенца мужеского пола.
REV|12|14|И даны были жене два крыла большого орла, чтобы она летела в пустыню в свое место от лица змия и там питалась в продолжение времени, времен и полвремени.
REV|12|15|И пустил змий из пасти своей вслед жены воду как реку, дабы увлечь ее рекою.
REV|12|16|Но земля помогла жене, и разверзла земля уста свои, и поглотила реку, которую пустил дракон из пасти своей.
REV|12|17|И рассвирепел дракон на жену, и пошел, чтобы вступить в брань с прочими от семени ее, сохраняющими заповеди Божии и имеющими свидетельство Иисуса Христа.
REV|13|1|И стал я на песке морском, и увидел выходящего из моря зверя с семью головами и десятью рогами: на рогах его было десять диадим, а на головах его имена богохульные.
REV|13|2|Зверь, которого я видел, был подобен барсу; ноги у него – как у медведя, а пасть у него – как пасть у льва; и дал ему дракон силу свою и престол свой и великую власть.
REV|13|3|И видел я, что одна из голов его как бы смертельно была ранена, но эта смертельная рана исцелела. И дивилась вся земля, следя за зверем, и поклонились дракону, который дал власть зверю,
REV|13|4|и поклонились зверю, говоря: кто подобен зверю сему? и кто может сразиться с ним?
REV|13|5|И даны были ему уста, говорящие гордо и богохульно, и дана ему власть действовать сорок два месяца.
REV|13|6|И отверз он уста свои для хулы на Бога, чтобы хулить имя Его, и жилище Его, и живущих на небе.
REV|13|7|И дано было ему вести войну со святыми и победить их; и дана была ему власть над всяким коленом и народом, и языком и племенем.
REV|13|8|И поклонятся ему все живущие на земле, которых имена не написаны в книге жизни у Агнца, закланного от создания мира.
REV|13|9|Кто имеет ухо, да слышит.
REV|13|10|Кто ведет в плен, тот сам пойдет в плен; кто мечом убивает, тому самому надлежит быть убиту мечом. Здесь терпение и вера святых.
REV|13|11|И увидел я другого зверя, выходящего из земли; он имел два рога, подобные агнчим, и говорил как дракон.
REV|13|12|Он действует перед ним со всею властью первого зверя и заставляет всю землю и живущих на ней поклоняться первому зверю, у которого смертельная рана исцелела;
REV|13|13|и творит великие знамения, так что и огонь низводит с неба на землю перед людьми.
REV|13|14|И чудесами, которые дано было ему творить перед зверем, он обольщает живущих на земле, говоря живущим на земле, чтобы они сделали образ зверя, который имеет рану от меча и жив.
REV|13|15|И дано ему было вложить дух в образ зверя, чтобы образ зверя и говорил и действовал так, чтобы убиваем был всякий, кто не будет поклоняться образу зверя.
REV|13|16|И он сделает то, что всем, малым и великим, богатым и нищим, свободным и рабам, положено будет начертание на правую руку их или на чело их,
REV|13|17|и что никому нельзя будет ни покупать, ни продавать, кроме того, кто имеет это начертание, или имя зверя, или число имени его.
REV|13|18|Здесь мудрость. Кто имеет ум, тот сочти число зверя, ибо это число человеческое; число его шестьсот шестьдесят шесть.
REV|14|1|И взглянул я, и вот, Агнец стоит на горе Сионе, и с Ним сто сорок четыре тысячи, у которых имя Отца Его написано на челах.
REV|14|2|И услышал я голос с неба, как шум от множества вод и как звук сильного грома; и услышал голос как бы гуслистов, играющих на гуслях своих.
REV|14|3|Они поют как бы новую песнь пред престолом и пред четырьмя животными и старцами; и никто не мог научиться сей песни, кроме сих ста сорока четырех тысяч, искупленных от земли.
REV|14|4|Это те, которые не осквернились с женами, ибо они девственники; это те, которые следуют за Агнцем, куда бы Он ни пошел. Они искуплены из людей, как первенцу Богу и Агнцу,
REV|14|5|и в устах их нет лукавства; они непорочны пред престолом Божиим.
REV|14|6|И увидел я другого Ангела, летящего по средине неба, который имел вечное Евангелие, чтобы благовествовать живущим на земле и всякому племени и колену, и языку и народу;
REV|14|7|и говорил он громким голосом: убойтесь Бога и воздайте Ему славу, ибо наступил час суда Его, и поклонитесь Сотворившему небо и землю, и море и источники вод.
REV|14|8|И другой Ангел следовал за ним, говоря: пал, пал Вавилон, город великий, потому что он яростным вином блуда своего напоил все народы.
REV|14|9|И третий Ангел последовал за ними, говоря громким голосом: кто поклоняется зверю и образу его и принимает начертание на чело свое, или на руку свою,
REV|14|10|тот будет пить вино ярости Божией, вино цельное, приготовленное в чаше гнева Его, и будет мучим в огне и сере пред святыми Ангелами и пред Агнцем;
REV|14|11|и дым мучения их будет восходить во веки веков, и не будут иметь покоя ни днем, ни ночью поклоняющиеся зверю и образу его и принимающие начертание имени его.
REV|14|12|Здесь терпение святых, соблюдающих заповеди Божии и веру в Иисуса.
REV|14|13|И услышал я голос с неба, говорящий мне: напиши: отныне блаженны мертвые, умирающие в Господе; ей, говорит Дух, они успокоятся от трудов своих, и дела их идут вслед за ними.
REV|14|14|И взглянул я, и вот светлое облако, и на облаке сидит подобный Сыну Человеческому; на голове его золотой венец, и в руке его острый серп.
REV|14|15|И вышел другой Ангел из храма и воскликнул громким голосом к сидящему на облаке: пусти серп твой и пожни, потому что пришло время жатвы, ибо жатва на земле созрела.
REV|14|16|И поверг сидящий на облаке серп свой на землю, и земля была пожата.
REV|14|17|И другой Ангел вышел из храма, находящегося на небе, также с острым серпом.
REV|14|18|И иной Ангел, имеющий власть над огнем, вышел от жертвенника и с великим криком воскликнул к имеющему острый серп, говоря: пусти острый серп твой и обрежь гроздья винограда на земле, потому что созрели на нем ягоды.
REV|14|19|И поверг Ангел серп свой на землю, и обрезал виноград на земле, и бросил в великое точило гнева Божия.
REV|14|20|И истоптаны [ягоды] в точиле за городом, и потекла кровь из точила даже до узд конских, на тысячу шестьсот стадий.
REV|15|1|И увидел я иное знамение на небе, великое и чудное: семь Ангелов, имеющих семь последних язв, которыми оканчивалась ярость Божия.
REV|15|2|И видел я как бы стеклянное море, смешанное с огнем; и победившие зверя и образ его, и начертание его и число имени его, стоят на этом стеклянном море, держа гусли Божии,
REV|15|3|и поют песнь Моисея, раба Божия, и песнь Агнца, говоря: велики и чудны дела Твои, Господи Боже Вседержитель! Праведны и истинны пути Твои, Царь святых!
REV|15|4|Кто не убоится Тебя, Господи, и не прославит имени Твоего? ибо Ты един свят. Все народы придут и поклонятся пред Тобою, ибо открылись суды Твои.
REV|15|5|И после сего я взглянул, и вот, отверзся храм скинии свидетельства на небе.
REV|15|6|И вышли из храма семь Ангелов, имеющие семь язв, облеченные в чистую и светлую льняную одежду и опоясанные по персям золотыми поясами.
REV|15|7|И одно из четырех животных дало семи Ангелам семь золотых чаш, наполненных гневом Бога, живущего во веки веков.
REV|15|8|И наполнился храм дымом от славы Божией и от силы Его, и никто не мог войти в храм, доколе не окончились семь язв семи Ангелов.
REV|16|1|И услышал я из храма громкий голос, говорящий семи Ангелам: идите и вылейте семь чаш гнева Божия на землю.
REV|16|2|Пошел первый Ангел и вылил чашу свою на землю: и сделались жестокие и отвратительные гнойные раны на людях, имеющих начертание зверя и поклоняющихся образу его.
REV|16|3|Второй Ангел вылил чашу свою в море: и сделалась кровь, как бы мертвеца, и все одушевленное умерло в море.
REV|16|4|Третий Ангел вылил чашу свою в реки и источники вод: и сделалась кровь.
REV|16|5|И услышал я Ангела вод, который говорил: праведен Ты, Господи, Который еси и был, и свят, потому что так судил;
REV|16|6|за то, что они пролили кровь святых и пророков, Ты дал им пить кровь: они достойны того.
REV|16|7|И услышал я другого от жертвенника говорящего: ей, Господи Боже Вседержитель, истинны и праведны суды Твои.
REV|16|8|Четвертый Ангел вылил чашу свою на солнце: и дано было ему жечь людей огнем.
REV|16|9|И жег людей сильный зной, и они хулили имя Бога, имеющего власть над сими язвами, и не вразумились, чтобы воздать Ему славу.
REV|16|10|Пятый Ангел вылил чашу свою на престол зверя: и сделалось царство его мрачно, и они кусали языки свои от страдания,
REV|16|11|и хулили Бога небесного от страданий своих и язв своих; и не раскаялись в делах своих.
REV|16|12|Шестой Ангел вылил чашу свою в великую реку Евфрат: и высохла в ней вода, чтобы готов был путь царям от восхода солнечного.
REV|16|13|И видел я [выходящих] из уст дракона и из уст зверя и из уст лжепророка трех духов нечистых, подобных жабам:
REV|16|14|это – бесовские духи, творящие знамения; они выходят к царям земли всей вселенной, чтобы собрать их на брань в оный великий день Бога Вседержителя.
REV|16|15|Се, иду как тать: блажен бодрствующий и хранящий одежду свою, чтобы не ходить ему нагим и чтобы не увидели срамоты его.
REV|16|16|И он собрал их на место, называемое по–еврейски Армагеддон.
REV|16|17|Седьмой Ангел вылил чашу свою на воздух: и из храма небесного от престола раздался громкий голос, говорящий: совершилось!
REV|16|18|И произошли молнии, громы и голоса, и сделалось великое землетрясение, какого не бывало с тех пор, как люди на земле. Такое землетрясение! Так великое!
REV|16|19|И город великий распался на три части, и города языческие пали, и Вавилон великий воспомянут пред Богом, чтобы дать ему чашу вина ярости гнева Его.
REV|16|20|И всякий остров убежал, и гор не стало;
REV|16|21|и град, величиною в талант, пал с неба на людей; и хулили люди Бога за язвы от града, потому что язва от него была весьма тяжкая.
REV|17|1|И пришел один из семи Ангелов, имеющих семь чаш, и, говоря со мною, сказал мне: подойди, я покажу тебе суд над великою блудницею, сидящею на водах многих;
REV|17|2|с нею блудодействовали цари земные, и вином ее блудодеяния упивались живущие на земле.
REV|17|3|И повел меня в духе в пустыню; и я увидел жену, сидящую на звере багряном, преисполненном именами богохульными, с семью головами и десятью рогами.
REV|17|4|И жена облечена была в порфиру и багряницу, украшена золотом, драгоценными камнями и жемчугом, и держала золотую чашу в руке своей, наполненную мерзостями и нечистотою блудодейства ее;
REV|17|5|и на челе ее написано имя: тайна, Вавилон великий, мать блудницам и мерзостям земным.
REV|17|6|Я видел, что жена упоена была кровью святых и кровью свидетелей Иисусовых, и видя ее, дивился удивлением великим.
REV|17|7|И сказал мне Ангел: что ты дивишься? я скажу тебе тайну жены сей и зверя, носящего ее, имеющего семь голов и десять рогов.
REV|17|8|Зверь, которого ты видел, был, и нет его, и выйдет из бездны, и пойдет в погибель; и удивятся те из живущих на земле, имена которых не вписаны в книгу жизни от начала мира, видя, что зверь был, и нет его, и явится.
REV|17|9|Здесь ум, имеющий мудрость. Семь голов суть семь гор, на которых сидит жена,
REV|17|10|и семь царей, из которых пять пали, один есть, а другой еще не пришел, и когда придет, не долго ему быть.
REV|17|11|И зверь, который был и которого нет, есть восьмой, и из числа семи, и пойдет в погибель.
REV|17|12|И десять рогов, которые ты видел, суть десять царей, которые еще не получили царства, но примут власть со зверем, как цари, на один час.
REV|17|13|Они имеют одни мысли и передадут силу и власть свою зверю.
REV|17|14|Они будут вести брань с Агнцем, и Агнец победит их; ибо Он есть Господь господствующих и Царь царей, и те, которые с Ним, суть званые и избранные и верные.
REV|17|15|И говорит мне: воды, которые ты видел, где сидит блудница, суть люди и народы, и племена и языки.
REV|17|16|И десять рогов, которые ты видел на звере, сии возненавидят блудницу, и разорят ее, и обнажат, и плоть ее съедят, и сожгут ее в огне;
REV|17|17|потому что Бог положил им на сердце – исполнить волю Его, исполнить одну волю, и отдать царство их зверю, доколе не исполнятся слова Божии.
REV|17|18|Жена же, которую ты видел, есть великий город, царствующий над земными царями.
REV|18|1|После сего я увидел иного Ангела, сходящего с неба и имеющего власть великую; земля осветилась от славы его.
REV|18|2|И воскликнул он сильно, громким голосом говоря: пал, пал Вавилон, великая [блудница], сделался жилищем бесов и пристанищем всякому нечистому духу, пристанищем всякой нечистой и отвратительной птице; ибо яростным вином блудодеяния своего она напоила все народы,
REV|18|3|и цари земные любодействовали с нею, и купцы земные разбогатели от великой роскоши ее.
REV|18|4|И услышал я иной голос с неба, говорящий: выйди от нее, народ Мой, чтобы не участвовать вам в грехах ее и не подвергнуться язвам ее;
REV|18|5|ибо грехи ее дошли до неба, и Бог воспомянул неправды ее.
REV|18|6|Воздайте ей так, как и она воздала вам, и вдвое воздайте ей по делам ее; в чаше, в которой она приготовляла вам вино, приготовьте ей вдвое.
REV|18|7|Сколько славилась она и роскошествовала, столько воздайте ей мучений и горестей. Ибо она говорит в сердце своем: "сижу царицею, я не вдова и не увижу горести!"
REV|18|8|За то в один день придут на нее казни, смерть и плач и голод, и будет сожжена огнем, потому что силен Господь Бог, судящий ее.
REV|18|9|И восплачут и возрыдают о ней цари земные, блудодействовавшие и роскошествовавшие с нею, когда увидят дым от пожара ее,
REV|18|10|стоя издали от страха мучений ее [и] говоря: горе, горе [тебе], великий город Вавилон, город крепкий! ибо в один час пришел суд твой.
REV|18|11|И купцы земные восплачут и возрыдают о ней, потому что товаров их никто уже не покупает,
REV|18|12|товаров золотых и серебряных, и камней драгоценных и жемчуга, и виссона и порфиры, и шелка и багряницы, и всякого благовонного дерева, и всяких изделий из слоновой кости, и всяких изделий из дорогих дерев, из меди и железа и мрамора,
REV|18|13|корицы и фимиама, и мира и ладана, и вина и елея, и муки и пшеницы, и скота и овец, и коней и колесниц, и тел и душ человеческих.
REV|18|14|И плодов, угодных для души твоей, не стало у тебя, и все тучное и блистательное удалилось от тебя; ты уже не найдешь его.
REV|18|15|Торговавшие всем сим, обогатившиеся от нее, станут вдали от страха мучений ее, плача и рыдая
REV|18|16|и говоря: горе, горе [тебе], великий город, одетый в виссон и порфиру и багряницу, украшенный золотом и камнями драгоценными и жемчугом,
REV|18|17|ибо в один час погибло такое богатство! И все кормчие, и все плывущие на кораблях, и все корабельщики, и все торгующие на море стали вдали
REV|18|18|и, видя дым от пожара ее, возопили, говоря: какой город подобен городу великому!
REV|18|19|И посыпали пеплом головы свои, и вопили, плача и рыдая: горе, горе [тебе], город великий, драгоценностями которого обогатились все, имеющие корабли на море, ибо опустел в один час!
REV|18|20|Веселись о сем, небо и святые Апостолы и пророки; ибо совершил Бог суд ваш над ним.
REV|18|21|И один сильный Ангел взял камень, подобный большому жернову, и поверг в море, говоря: с таким стремлением повержен будет Вавилон, великий город, и уже не будет его.
REV|18|22|И голоса играющих на гуслях, и поющих, и играющих на свирелях, и трубящих трубами в тебе уже не слышно будет; не будет уже в тебе никакого художника, никакого художества, и шума от жерновов не слышно уже будет в тебе;
REV|18|23|и свет светильника уже не появится в тебе; и голоса жениха и невесты не будет уже слышно в тебе: ибо купцы твои были вельможи земли, и волшебством твоим введены в заблуждение все народы.
REV|18|24|И в нем найдена кровь пророков и святых и всех убитых на земле.
REV|19|1|После сего я услышал на небе громкий голос как бы многочисленного народа, который говорил: аллилуия! спасение и слава, и честь и сила Господу нашему!
REV|19|2|Ибо истинны и праведны суды Его: потому что Он осудил ту великую любодейцу, которая растлила землю любодейством своим, и взыскал кровь рабов Своих от руки ее.
REV|19|3|И вторично сказали: аллилуия! И дым ее восходил во веки веков.
REV|19|4|Тогда двадцать четыре старца и четыре животных пали и поклонились Богу, сидящему на престоле, говоря: аминь! аллилуия!
REV|19|5|И голос от престола исшел, говорящий: хвалите Бога нашего, все рабы Его и боящиеся Его, малые и великие.
REV|19|6|И слышал я как бы голос многочисленного народа, как бы шум вод многих, как бы голос громов сильных, говорящих: аллилуия! ибо воцарился Господь Бог Вседержитель.
REV|19|7|Возрадуемся и возвеселимся и воздадим Ему славу; ибо наступил брак Агнца, и жена Его приготовила себя.
REV|19|8|И дано было ей облечься в виссон чистый и светлый; виссон же есть праведность святых.
REV|19|9|И сказал мне [Ангел]: напиши: блаженны званые на брачную вечерю Агнца. И сказал мне: сии суть истинные слова Божии.
REV|19|10|Я пал к ногам его, чтобы поклониться ему; но он сказал мне: смотри, не делай сего; я сослужитель тебе и братьям твоим, имеющим свидетельство Иисусово; Богу поклонись; ибо свидетельство Иисусово есть дух пророчества.
REV|19|11|И увидел я отверстое небо, и вот конь белый, и сидящий на нем называется Верный и Истинный, Который праведно судит и воинствует.
REV|19|12|Очи у Него как пламень огненный, и на голове Его много диадим. [Он] имел имя написанное, которого никто не знал, кроме Его Самого.
REV|19|13|[Он был] облечен в одежду, обагренную кровью. Имя Ему: "Слово Божие".
REV|19|14|И воинства небесные следовали за Ним на конях белых, облеченные в виссон белый и чистый.
REV|19|15|Из уст же Его исходит острый меч, чтобы им поражать народы. Он пасет их жезлом железным; Он топчет точило вина ярости и гнева Бога Вседержителя.
REV|19|16|На одежде и на бедре Его написано имя: "Царь царей и Господь господствующих".
REV|19|17|И увидел я одного Ангела, стоящего на солнце; и он воскликнул громким голосом, говоря всем птицам, летающим по средине неба: летите, собирайтесь на великую вечерю Божию,
REV|19|18|чтобы пожрать трупы царей, трупы сильных, трупы тысяченачальников, трупы коней и сидящих на них, трупы всех свободных и рабов, и малых и великих.
REV|19|19|И увидел я зверя и царей земных и воинства их, собранные, чтобы сразиться с Сидящим на коне и с воинством Его.
REV|19|20|И схвачен был зверь и с ним лжепророк, производивший чудеса пред ним, которыми он обольстил принявших начертание зверя и поклоняющихся его изображению: оба живые брошены в озеро огненное, горящее серою;
REV|19|21|а прочие убиты мечом Сидящего на коне, исходящим из уст Его, и все птицы напитались их трупами.
REV|20|1|И увидел я Ангела, сходящего с неба, который имел ключ от бездны и большую цепь в руке своей.
REV|20|2|Он взял дракона, змия древнего, который есть диавол и сатана, и сковал его на тысячу лет,
REV|20|3|и низверг его в бездну, и заключил его, и положил над ним печать, дабы не прельщал уже народы, доколе не окончится тысяча лет; после же сего ему должно быть освобожденным на малое время.
REV|20|4|И увидел я престолы и сидящих на них, которым дано было судить, и души обезглавленных за свидетельство Иисуса и за слово Божие, которые не поклонились зверю, ни образу его, и не приняли начертания на чело свое и на руку свою. Они ожили и царствовали со Христом тысячу лет.
REV|20|5|Прочие же из умерших не ожили, доколе не окончится тысяча лет. Это – первое воскресение.
REV|20|6|Блажен и свят имеющий участие в воскресении первом: над ними смерть вторая не имеет власти, но они будут священниками Бога и Христа и будут царствовать с Ним тысячу лет.
REV|20|7|Когда же окончится тысяча лет, сатана будет освобожден из темницы своей и выйдет обольщать народы, находящиеся на четырех углах земли, Гога и Магога, и собирать их на брань; число их как песок морской.
REV|20|8|И вышли на широту земли, и окружили стан святых и город возлюбленный.
REV|20|9|И ниспал огонь с неба от Бога и пожрал их;
REV|20|10|а диавол, прельщавший их, ввержен в озеро огненное и серное, где зверь и лжепророк, и будут мучиться день и ночь во веки веков.
REV|20|11|И увидел я великий белый престол и Сидящего на нем, от лица Которого бежало небо и земля, и не нашлось им места.
REV|20|12|И увидел я мертвых, малых и великих, стоящих пред Богом, и книги раскрыты были, и иная книга раскрыта, которая есть книга жизни; и судимы были мертвые по написанному в книгах, сообразно с делами своими.
REV|20|13|Тогда отдало море мертвых, бывших в нем, и смерть и ад отдали мертвых, которые были в них; и судим был каждый по делам своим.
REV|20|14|И смерть и ад повержены в озеро огненное. Это смерть вторая.
REV|20|15|И кто не был записан в книге жизни, тот был брошен в озеро огненное.
REV|21|1|И увидел я новое небо и новую землю, ибо прежнее небо и прежняя земля миновали, и моря уже нет.
REV|21|2|И я, Иоанн, увидел святый город Иерусалим, новый, сходящий от Бога с неба, приготовленный как невеста, украшенная для мужа своего.
REV|21|3|И услышал я громкий голос с неба, говорящий: се, скиния Бога с человеками, и Он будет обитать с ними; они будут Его народом, и Сам Бог с ними будет Богом их.
REV|21|4|И отрет Бог всякую слезу с очей их, и смерти не будет уже; ни плача, ни вопля, ни болезни уже не будет, ибо прежнее прошло.
REV|21|5|И сказал Сидящий на престоле: се, творю все новое. И говорит мне: напиши; ибо слова сии истинны и верны.
REV|21|6|И сказал мне: совершилось! Я есмь Альфа и Омега, начало и конец; жаждущему дам даром от источника воды живой.
REV|21|7|Побеждающий наследует все, и буду ему Богом, и он будет Мне сыном.
REV|21|8|Боязливых же и неверных, и скверных и убийц, и любодеев и чародеев, и идолослужителей и всех лжецов участь в озере, горящем огнем и серою. Это смерть вторая.
REV|21|9|И пришел ко мне один из семи Ангелов, у которых было семь чаш, наполненных семью последними язвами, и сказал мне: пойди, я покажу тебе жену, невесту Агнца.
REV|21|10|И вознес меня в духе на великую и высокую гору, и показал мне великий город, святый Иерусалим, который нисходил с неба от Бога.
REV|21|11|Он имеет славу Божию. Светило его подобно драгоценнейшему камню, как бы камню яспису кристалловидному.
REV|21|12|Он имеет большую и высокую стену, имеет двенадцать ворот и на них двенадцать Ангелов; на воротах написаны имена двенадцати колен сынов Израилевых:
REV|21|13|с востока трое ворот, с севера трое ворот, с юга трое ворот, с запада трое ворот.
REV|21|14|Стена города имеет двенадцать оснований, и на них имена двенадцати Апостолов Агнца.
REV|21|15|Говоривший со мною имел золотую трость для измерения города и ворот его и стены его.
REV|21|16|Город расположен четвероугольником, и длина его такая же, как и широта. И измерил он город тростью на двенадцать тысяч стадий; длина и широта и высота его равны.
REV|21|17|И стену его измерил во сто сорок четыре локтя, мерою человеческою, какова мера и Ангела.
REV|21|18|Стена его построена из ясписа, а город был чистое золото, подобен чистому стеклу.
REV|21|19|Основания стены города украшены всякими драгоценными камнями: основание первое яспис, второе сапфир, третье халкидон, четвертое смарагд,
REV|21|20|пятое сардоникс, шестое сердолик, седьмое хризолит, восьмое вирилл, девятое топаз, десятое хризопрас, одиннадцатое гиацинт, двенадцатое аметист.
REV|21|21|А двенадцать ворот – двенадцать жемчужин: каждые ворота были из одной жемчужины. Улица города – чистое золото, как прозрачное стекло.
REV|21|22|Храма же я не видел в нем, ибо Господь Бог Вседержитель – храм его, и Агнец.
REV|21|23|И город не имеет нужды ни в солнце, ни в луне для освещения своего, ибо слава Божия осветила его, и светильник его – Агнец.
REV|21|24|Спасенные народы будут ходить во свете его, и цари земные принесут в него славу и честь свою.
REV|21|25|Ворота его не будут запираться днем; а ночи там не будет.
REV|21|26|И принесут в него славу и честь народов.
REV|21|27|И не войдет в него ничто нечистое и никто преданный мерзости и лжи, а только те, которые написаны у Агнца в книге жизни.
REV|22|1|И показал мне чистую реку воды жизни, светлую, как кристалл, исходящую от престола Бога и Агнца.
REV|22|2|Среди улицы его, и по ту и по другую сторону реки, древо жизни, двенадцать [раз] приносящее плоды, дающее на каждый месяц плод свой; и листья дерева – для исцеления народов.
REV|22|3|И ничего уже не будет проклятого; но престол Бога и Агнца будет в нем, и рабы Его будут служить Ему.
REV|22|4|И узрят лице Его, и имя Его будет на челах их.
REV|22|5|И ночи не будет там, и не будут иметь нужды ни в светильнике, ни в свете солнечном, ибо Господь Бог освещает их; и будут царствовать во веки веков.
REV|22|6|И сказал мне: сии слова верны и истинны; и Господь Бог святых пророков послал Ангела Своего показать рабам Своим то, чему надлежит быть вскоре.
REV|22|7|Се, гряду скоро: блажен соблюдающий слова пророчества книги сей.
REV|22|8|Я, Иоанн, видел и слышал сие. Когда же услышал и увидел, пал к ногам Ангела, показывающего мне сие, чтобы поклониться [ему];
REV|22|9|но он сказал мне: смотри, не делай сего; ибо я сослужитель тебе и братьям твоим пророкам и соблюдающим слова книги сей; Богу поклонись.
REV|22|10|И сказал мне: не запечатывай слов пророчества книги сей; ибо время близко.
REV|22|11|Неправедный пусть еще делает неправду; нечистый пусть еще сквернится; праведный да творит правду еще, и святый да освящается еще.
REV|22|12|Се, гряду скоро, и возмездие Мое со Мною, чтобы воздать каждому по делам его.
REV|22|13|Я есмь Альфа и Омега, начало и конец, Первый и Последний.
REV|22|14|Блаженны те, которые соблюдают заповеди Его, чтобы иметь им право на древо жизни и войти в город воротами.
REV|22|15|А вне – псы и чародеи, и любодеи, и убийцы, и идолослужители, и всякий любящий и делающий неправду.
REV|22|16|Я, Иисус, послал Ангела Моего засвидетельствовать вам сие в церквах. Я есмь корень и потомок Давида, звезда светлая и утренняя.
REV|22|17|И Дух и невеста говорят: прииди! И слышавший да скажет прииди! Жаждущий пусть приходит, и желающий пусть берет воду жизни даром.
REV|22|18|И я также свидетельствую всякому слышащему слова пророчества книги сей: если кто приложит что к ним, на того наложит Бог язвы, о которых написано в книге сей;
REV|22|19|и если кто отнимет что от слов книги пророчества сего, у того отнимет Бог участие в книге жизни и в святом граде и в том, что написано в книге сей.
REV|22|20|Свидетельствующий сие говорит: ей, гряду скоро! Аминь. Ей, гряди, Господи Иисусе!
REV|22|21|Благодать Господа нашего Иисуса Христа со всеми вами. Аминь.
