2THESS|1|1|Paul, Silvanus, and Timothy, To the church of the Thessalonians in God our Father and the Lord Jesus Christ:
2THESS|1|2|Grace to you and peace from God our Father and the Lord Jesus Christ.
2THESS|1|3|We ought always to give thanks to God for you, brothers, as is right, because your faith is growing abundantly, and the love of every one of you for one another is increasing.
2THESS|1|4|Therefore we ourselves boast about you in the churches of God for your steadfastness and faith in all your persecutions and in the afflictions that you are enduring.
2THESS|1|5|This is evidence of the righteous judgment of God, that you may be considered worthy of the kingdom of God, for which you are also suffering-
2THESS|1|6|since indeed God considers it just to repay with affliction those who afflict you,
2THESS|1|7|and to grant relief to you who are afflicted as well as to us, when the Lord Jesus is revealed from heaven with his mighty angels
2THESS|1|8|in flaming fire, inflicting vengeance on those who do not know God and on those who do not obey the gospel of our Lord Jesus.
2THESS|1|9|They will suffer the punishment of eternal destruction, away from the presence of the Lord and from the glory of his might,
2THESS|1|10|when he comes on that day to be glorified in his saints, and to be marveled at among all who have believed, because our testimony to you was believed.
2THESS|1|11|To this end we always pray for you, that our God may make you worthy of his calling and may fulfill every resolve for good and every work of faith by his power,
2THESS|1|12|so that the name of our Lord Jesus may be glorified in you, and you in him, according to the grace of our God and the Lord Jesus Christ.
2THESS|2|1|Now concerning the coming of our Lord Jesus Christ and our being gathered together to him, we ask you, brothers,
2THESS|2|2|not to be quickly shaken in mind or alarmed, either by a spirit or a spoken word, or a letter seeming to be from us, to the effect that the day of the Lord has come.
2THESS|2|3|Let no one deceive you in any way. For that day will not come, unless the rebellion comes first, and the man of lawlessness is revealed, the son of destruction,
2THESS|2|4|who opposes and exalts himself against every so-called god or object of worship, so that he takes his seat in the temple of God, proclaiming himself to be God.
2THESS|2|5|Do you not remember that when I was still with you I told you these things?
2THESS|2|6|And you know what is restraining him now so that he may be revealed in his time.
2THESS|2|7|For the mystery of lawlessness is already at work. Only he who now restrains it will do so until he is out of the way.
2THESS|2|8|And then the lawless one will be revealed, whom the Lord Jesus will kill with the breath of his mouth and bring to nothing by the appearance of his coming.
2THESS|2|9|The coming of the lawless one is by the activity of Satan with all power and false signs and wonders,
2THESS|2|10|and with all wicked deception for those who are perishing, because they refused to love the truth and so be saved.
2THESS|2|11|Therefore God sends them a strong delusion, so that they may believe what is false,
2THESS|2|12|in order that all may be condemned who did not believe the truth but had pleasure in unrighteousness.
2THESS|2|13|But we ought always to give thanks to God for you, brothers beloved by the Lord, because God chose you as the first fruits to be saved, through sanctification by the Spirit and belief in the truth.
2THESS|2|14|To this he called you through our gospel, so that you may obtain the glory of our Lord Jesus Christ.
2THESS|2|15|So then, brothers, stand firm and hold to the traditions that you were taught by us, either by our spoken word or by our letter.
2THESS|2|16|Now may our Lord Jesus Christ himself, and God our Father, who loved us and gave us eternal comfort and good hope through grace,
2THESS|2|17|comfort your hearts and establish them in every good work and word.
2THESS|3|1|Finally, brothers, pray for us, that the word of the Lord may speed ahead and be honored, as happened among you,
2THESS|3|2|and that we may be delivered from wicked and evil men. For not all have faith.
2THESS|3|3|But the Lord is faithful. He will establish you and guard you against the evil one.
2THESS|3|4|And we have confidence in the Lord about you, that you are doing and will do the things that we command.
2THESS|3|5|May the Lord direct your hearts to the love of God and to the steadfastness of Christ.
2THESS|3|6|Now we command you, brothers, in the name of our Lord Jesus Christ, that you keep away from any brother who is walking in idleness and not in accord with the tradition that you received from us.
2THESS|3|7|For you yourselves know how you ought to imitate us, because we were not idle when we were with you,
2THESS|3|8|nor did we eat anyone's bread without paying for it, but with toil and labor we worked night and day, that we might not be a burden to any of you.
2THESS|3|9|It was not because we do not have that right, but to give you in ourselves an example to imitate.
2THESS|3|10|For even when we were with you, we would give you this command: If anyone is not willing to work, let him not eat.
2THESS|3|11|For we hear that some among you walk in idleness, not busy at work, but busybodies.
2THESS|3|12|Now such persons we command and encourage in the Lord Jesus Christ to do their work quietly and to earn their own living.
2THESS|3|13|As for you, brothers, do not grow weary in doing good.
2THESS|3|14|If anyone does not obey what we say in this letter, take note of that person, and have nothing to do with him, that he may be ashamed.
2THESS|3|15|Do not regard him as an enemy, but warn him as a brother.
2THESS|3|16|Now may the Lord of peace himself give you peace at all times in every way. The Lord be with you all.
2THESS|3|17|I, Paul, write this greeting with my own hand. This is the sign of genuineness in every letter of mine; it is the way I write.
2THESS|3|18|The grace of our Lord Jesus Christ be with you all.
