1CHR|1|1|亚当 ， 塞特 ， 以挪士 ，
1CHR|1|2|该南 ， 玛勒列 ， 雅列 ，
1CHR|1|3|以诺 ， 玛土撒拉 ， 拉麦 ，
1CHR|1|4|挪亚 ， 闪 ， 含 ， 雅弗 。
1CHR|1|5|雅弗 的儿子是 歌篾 、 玛各 、 玛代 、 雅完 、 土巴 、 米设 和 提拉 。
1CHR|1|6|歌篾 的儿子是 亚实基拿 、 低法 和 陀迦玛 。
1CHR|1|7|雅完 的儿子是 以利沙 、 他施 、 基提 和 罗单 人 。
1CHR|1|8|含 的儿子是 古实 、 麦西 、 弗 和 迦南 。
1CHR|1|9|古实 的儿子是 西巴 、 哈腓拉 、 撒弗他 、 拉玛 和 撒弗提迦 。 拉玛 的儿子是 示巴 和 底但 。
1CHR|1|10|古实 又生 宁录 ，他是地上第一个勇士。
1CHR|1|11|麦西 生 路低 人、 亚拿米 人、 利哈比 人、 拿弗土希 人、
1CHR|1|12|帕斯鲁细 人、 迦斯路希 人和 迦斐托 人； 非利士 人是从 迦斐托 人 出来的。
1CHR|1|13|迦南 生了长子 西顿 ，又生 赫
1CHR|1|14|和 耶布斯 人、 亚摩利 人、 革迦撒 人、
1CHR|1|15|希未 人、 亚基 人、 西尼 人、
1CHR|1|16|亚瓦底 人、 洗玛利 人和 哈马 人。
1CHR|1|17|闪 的儿子是 以拦 、 亚述 、 亚法撒 、 路德 、 亚兰 、 乌斯 、 户勒 、 基帖 和 米设 。
1CHR|1|18|亚法撒 生 沙拉 ； 沙拉 生 希伯 。
1CHR|1|19|希伯 生了两个儿子：一个名叫 法勒 ，因为那时人分地居住； 法勒 的兄弟名叫 约坍 。
1CHR|1|20|约坍 生 亚摩答 、 沙列 、 哈萨玛非 、 耶拉 、
1CHR|1|21|哈多兰 、 乌萨 、 德拉 、
1CHR|1|22|以巴录 、 亚比玛利 、 示巴 、
1CHR|1|23|阿斐 、 哈腓拉 和 约巴 。这些都是 约坍 的儿子。
1CHR|1|24|闪 ， 亚法撒 ， 沙拉 ，
1CHR|1|25|希伯 ， 法勒 ， 拉吴 ，
1CHR|1|26|西鹿 ， 拿鹤 ， 他拉 ，
1CHR|1|27|亚伯兰 ， 亚伯兰 就是 亚伯拉罕 。
1CHR|1|28|亚伯拉罕 的儿子是 以撒 和 以实玛利 。
1CHR|1|29|以实玛利 的后代如下： 以实玛利 的长子是 尼拜约 ，又有 基达 、 亚德别 、 米比衫 、
1CHR|1|30|米施玛 、 度玛 、 玛撒 、 哈大 、 提玛 、
1CHR|1|31|伊突 、 拿非施 和 基底玛 。这些都是 以实玛利 的儿子。
1CHR|1|32|亚伯拉罕 的妾 基土拉 所生的儿子，就是 心兰 、 约珊 、 米但 、 米甸 、 伊施巴 和 书亚 。 约珊 的儿子是 示巴 和 底但 。
1CHR|1|33|米甸 的儿子是 以法 、 以弗 、 哈诺 、 亚比大 和 以勒大 。这些都是 基土拉 的子孙。
1CHR|1|34|亚伯拉罕 生 以撒 ； 以撒 的儿子是 以扫 和 以色列 。
1CHR|1|35|以扫 的儿子是 以利法 、 流珥 、 耶乌施 、 雅兰 和 可拉 。
1CHR|1|36|以利法 的儿子是 提幔 、 阿抹 、 洗玻 、 迦坦 、 基纳斯 、 亭纳 和 亚玛力 。
1CHR|1|37|流珥 的儿子是 拿哈 、 谢拉 、 沙玛 和 米撒 。
1CHR|1|38|西珥 的儿子是 罗坍 、 朔巴 、 祭便 、 亚拿 、 底顺 、 以察 和 底珊 。
1CHR|1|39|罗坍 的儿子是 何利 和 荷幔 ； 罗坍 的妹妹是 亭纳 。
1CHR|1|40|朔巴 的儿子是 亚勒文 、 玛拿辖 、 以巴录 、 示非 和 阿南 。 祭便 的儿子是 爱亚 和 亚拿 。
1CHR|1|41|亚拿 的儿子是 底顺 。 底顺 的儿子是 哈默兰 、 伊是班 、 益兰 和 基兰 。
1CHR|1|42|以察 的儿子是 辟罕 、 撒番 ，和 亚干 。 底珊 的儿子是 乌斯 和 亚兰 。
1CHR|1|43|以色列 人未有君王治理之前，这些是在 以东 地作王的。有 比珥 的儿子 比拉 ，他的城名叫 亭哈巴 。
1CHR|1|44|比拉 死了， 波斯拉 人 谢拉 的儿子 约巴 接续他作王。
1CHR|1|45|约巴 死了， 提幔 人之地的 户珊 接续他作王。
1CHR|1|46|户珊 死了， 比达 的儿子 哈达 接续他作王， 哈达 曾在 摩押 地击败 米甸 人，他的城名叫 亚未得 。
1CHR|1|47|哈达 死了， 玛士利加 人 桑拉 接续他作王。
1CHR|1|48|桑拉 死了， 大河 边的 利河伯 人 扫罗 接续他作王。
1CHR|1|49|扫罗 死了， 亚革波 的儿子 巴勒．哈南 接续他作王。
1CHR|1|50|巴勒．哈南 死了， 哈达 接续他作王，他的城名叫 巴伊 。他的妻子名叫 米希她别 ，是 米．萨合 的孙女， 玛特列 的女儿。
1CHR|1|51|哈达 死了。 以东 的族长有： 亭纳 族长、 亚勒瓦 族长、 耶帖 族长、
1CHR|1|52|阿何利巴玛 族长、 以拉 族长、 比嫩 族长、
1CHR|1|53|基纳斯 族长、 提幔 族长、 米比萨 族长、
1CHR|1|54|玛基叠 族长、 以兰 族长。这些都是 以东 的族长。
1CHR|2|1|以色列 的儿子是 吕便 、 西缅 、 利未 、 犹大 、 以萨迦 、 西布伦 、
1CHR|2|2|但 、 约瑟 、 便雅悯 、 拿弗他利 、 迦得 和 亚设 。
1CHR|2|3|犹大 的儿子是 珥 、 俄南 和 示拉 ，这三人是 迦南 女子 拔．书亚 所生的。 犹大 的长子 珥 在耶和华眼中看为恶，耶和华就杀死了他。
1CHR|2|4|犹大 的媳妇 她玛 为 犹大 生了 法勒斯 和 谢拉 。 犹大 共有五个儿子。
1CHR|2|5|法勒斯 的儿子是 希斯仑 和 哈母勒 。
1CHR|2|6|谢拉 的儿子是 心利 、 以探 、 希幔 、 甲各 和 大拉 ，共五人。
1CHR|2|7|迦米 的儿子是 亚迦 ，他在当灭的物上犯了罪，连累了 以色列 人。
1CHR|2|8|以探 的儿子是 亚撒利雅 。
1CHR|2|9|希斯仑 所生的儿子是 耶拉篾 、 兰 和 基路拜 。
1CHR|2|10|兰 生 亚米拿达 ； 亚米拿达 生 拿顺 ， 拿顺 是 犹大 人的领袖。
1CHR|2|11|拿顺 生 撒门 ； 撒门 生 波阿斯 ；
1CHR|2|12|波阿斯 生 俄备得 ； 俄备得 生 耶西 ；
1CHR|2|13|耶西 生长子 以利押 ，次子 亚比拿达 ，三子 示米亚 ，
1CHR|2|14|四子 拿坦业 ，五子 拉代 ，
1CHR|2|15|六子 阿鲜 ，七子 大卫 。
1CHR|2|16|他们的姊妹是 洗鲁雅 和 亚比该 。 洗鲁雅 的儿子是 亚比筛 、 约押 和 亚撒黑 ，共三人。
1CHR|2|17|亚比该 生 亚玛撒 ； 亚玛撒 的父亲是 以实玛利 人 益帖 。
1CHR|2|18|希斯仑 的儿子 迦勒 娶 阿苏巴 和 耶略 为妻， 阿苏巴 的儿子是 耶设 、 朔罢 和 押墩 。
1CHR|2|19|阿苏巴 死了， 迦勒 又娶 以法她 ，生了 户珥 。
1CHR|2|20|户珥 生 乌利 ； 乌利 生 比撒列 。
1CHR|2|21|后来， 希斯仑 六十岁时娶了 基列 的父亲 玛吉 的女儿，与她同房； 玛吉 的女儿为他生了 西割 ；
1CHR|2|22|西割 生 睚珥 。 睚珥 在 基列 地有二十三座城。
1CHR|2|23|后来 基述 和 亚兰 夺了 哈倭特．睚珥 ，以及 基纳 和所属的乡镇 ，共六十个。这些城镇的人全都是 基列 的父亲 玛吉 的子孙。
1CHR|2|24|希斯仑 在 迦勒．以法他 死后，他的妻子 亚比雅 为他生了 提哥亚 的父亲 亚施户 。
1CHR|2|25|希斯仑 的长子 耶拉篾 的儿子有长子 兰 、 布拿 、 阿连 、 阿鲜 和 亚希雅 。
1CHR|2|26|耶拉篾 又娶一妻名叫 亚她拉 ，是 阿南 的母亲。
1CHR|2|27|耶拉篾 的长子 兰 的儿子有 玛斯 、 雅悯 和 以结 。
1CHR|2|28|阿南 的儿子是 沙买 和 雅大 。 沙买 的儿子是 拿答 和 亚比述 。
1CHR|2|29|亚比述 的妻子名叫 亚比孩 ，为他生了 亚办 和 摩利 。
1CHR|2|30|拿答 的儿子是 西列 和 亚遍 ； 西列 死了，没有儿子。
1CHR|2|31|亚遍 的儿子是 以示 ； 以示 的儿子是 示珊 ； 示珊 的儿子是 亚来 。
1CHR|2|32|沙买 的兄弟 雅大 的儿子是 益帖 和 约拿单 ； 益帖 死了，没有儿子。
1CHR|2|33|约拿单 的儿子是 比勒 和 撒萨 。这些都是 耶拉篾 的子孙。
1CHR|2|34|示珊 没有儿子，只有女儿。 示珊 有一个仆人名叫 耶哈 ，是 埃及 人。
1CHR|2|35|示珊 把女儿嫁给仆人 耶哈 ，她为他生了 亚太 。
1CHR|2|36|亚太 生 拿单 ； 拿单 生 撒拔 ；
1CHR|2|37|撒拔 生 以弗拉 ； 以弗拉 生 俄备得 ；
1CHR|2|38|俄备得 生 耶户 ； 耶户 生 亚撒利雅 ；
1CHR|2|39|亚撒利雅 生 希利斯 ； 希利斯 生 以利亚萨 ；
1CHR|2|40|以利亚萨 生 西斯买 ； 西斯买 生 沙龙 ；
1CHR|2|41|沙龙 生 耶加米雅 ； 耶加米雅 生 以利沙玛 。
1CHR|2|42|耶拉篾 的兄弟 迦勒 的众儿子：长子是 米沙 ， 米沙 是 西弗 的父亲，还有 希伯伦 的父亲 玛利沙 的众儿子。
1CHR|2|43|希伯伦 的儿子是 可拉 、 他普亚 、 利肯 和 示玛 。
1CHR|2|44|示玛 生 拉含 ，是 约干 之祖。 利肯 生 沙买 。
1CHR|2|45|沙买 的儿子是 玛云 ； 玛云 是 伯．夙 的父亲。
1CHR|2|46|迦勒 的妾 以法 生 哈兰 、 摩撒 和 迦谢 ； 哈兰 生 迦卸 。
1CHR|2|47|雅代 的儿子是 利健 、 约坦 、 基珊 、 毗力 、 以法 和 沙亚弗 。
1CHR|2|48|迦勒 的妾 玛迦 生 示别 和 特哈拿 ，
1CHR|2|49|又生 麦玛拿 的父亲 沙亚弗 ，又生 抹比拿 和 基比亚 的父亲 示法 。 迦勒 的女儿是 押撒 。
1CHR|2|50|这些都是 迦勒 的子孙。 以法她 的长子 户珥 的子孙： 基列．耶琳 之祖 朔巴 ，
1CHR|2|51|伯利恒 之祖 萨玛 ， 伯．迦得 之祖 哈勒 。
1CHR|2|52|基列．耶琳 之祖 朔巴 的子孙是 哈罗以 和一半的 米努哈 人 。
1CHR|2|53|基列．耶琳 的宗族有 以帖 人、 布特 人、 舒玛 人、 密来 人，又从这些宗族生出 琐拉 人和 以实陶 人。
1CHR|2|54|萨玛 的子孙有 伯利恒 人、 尼陀法 人、 亚他绿．伯．约押 人、一半的 玛拿哈 人、 琐利 人。
1CHR|2|55|住 雅比斯 的文士的宗族有 特拉 人、 示米押 人和 苏甲 人。这些都是 利甲 家之祖 哈末 所生的 基尼 人。
1CHR|3|1|大卫 在 希伯仑 所生的儿子如下：长子 暗嫩 是 耶斯列 人 亚希暖 生的。次子 但以利 是 迦密 人 亚比该 生的。
1CHR|3|2|三子 押沙龙 是 基述 王 达买 的女儿 玛迦 生的。四子 亚多尼雅 是 哈及 生的。
1CHR|3|3|五子 示法提雅 是 亚比她 生的。六子 以特念 是 大卫 的妻子 以格拉 生的。
1CHR|3|4|这六人都是 大卫 在 希伯仑 生的。 大卫 在 希伯仑 作王七年六个月，在 耶路撒冷 作王三十三年。
1CHR|3|5|大卫 在 耶路撒冷 所生的儿子是 示米亚 、 朔罢 、 拿单 和 所罗门 。这四人是 亚米利 的女儿 拔．书亚 生的。
1CHR|3|6|还有 益辖 、 以利沙玛 、 以利法列 、
1CHR|3|7|挪迦 、 尼斐 、 雅非亚 、
1CHR|3|8|以利沙玛 、 以利雅大 、 以利法列 ，共九人。
1CHR|3|9|这些全都是 大卫 的儿子，妃嫔的儿子不在其内； 她玛 是他们的妹妹。
1CHR|3|10|所罗门 的后裔如下： 罗波安 ，他的儿子 亚比雅 ，他的儿子 亚撒 ，他的儿子 约沙法 ，
1CHR|3|11|他的儿子 约兰 ，他的儿子 亚哈谢 ，他的儿子 约阿施 ，
1CHR|3|12|他的儿子 亚玛谢 ，他的儿子 亚撒利雅 ，他的儿子 约坦 ；
1CHR|3|13|他的儿子 亚哈斯 ，他的儿子 希西家 ，他的儿子 玛拿西 ，
1CHR|3|14|他的儿子 亚们 ，他的儿子 约西亚 ，
1CHR|3|15|他的长子 约哈难 ，次子 约雅敬 ，三子 西底家 ，四子 沙龙 。
1CHR|3|16|约雅敬 的后裔：他的儿子 耶哥尼雅 ，他的儿子 西底家 。
1CHR|3|17|被掳的 耶哥尼雅 的后裔如下：他的儿子 撒拉铁 、
1CHR|3|18|玛基兰 、 毗大雅 、 示拿萨 、 耶加米 、 何沙玛 和 尼大比雅 。
1CHR|3|19|毗大雅 的儿子是 所罗巴伯 和 示每 。 所罗巴伯 的儿子是 米书兰 和 哈拿尼雅 ， 示罗密 是他们的妹妹；
1CHR|3|20|还有 哈舒巴 、 阿黑 、 比利家 、 哈撒底 、 于沙．希悉 ，共五人。
1CHR|3|21|哈拿尼雅 的儿子是 毗拉提 和 耶筛亚 。还有 利法雅 的众儿子， 亚珥难 的众儿子， 俄巴底亚 的众儿子， 示迦尼 的众儿子。
1CHR|3|22|示迦尼 的后裔： 示玛雅 ， 示玛雅 的儿子 哈突 、 以甲 、 巴利亚 、 尼利雅 、 沙法 ，共六人。
1CHR|3|23|尼利雅 的儿子是 以利约乃 、 希西家 、 亚斯利干 ，共三人。
1CHR|3|24|以利约乃 的儿子是 何大雅 、 以利亚实 、 毗莱雅 、 阿谷 、 约哈难 、 第莱雅 、 阿拿尼 ，共七人。
1CHR|4|1|犹大 的儿子是 法勒斯 、 希斯仑 、 迦米 、 户珥 和 朔巴 。
1CHR|4|2|朔巴 的儿子 利亚雅 生 雅哈 ； 雅哈 生 亚户买 和 拉哈 。这些是 琐拉 人的宗族。
1CHR|4|3|以坦 之祖 是 耶斯列 、 伊施玛 和 伊得巴 ；他们的妹妹名叫 哈悉勒玻尼 。
1CHR|4|4|基多 之祖是 毗努伊勒 。 户沙 之祖是 以谢珥 。这些都是 伯利恒 之祖， 以法她 的长子 户珥 的后裔。
1CHR|4|5|提哥亚 的父亲 亚施户 有两个妻子， 希拉 和 拿拉 。
1CHR|4|6|拿拉 为 亚施户 生 亚户撒 、 希弗 、 提米尼 和 哈辖斯他利 。这些都是 拿拉 的儿子。
1CHR|4|7|希拉 生的是 洗列 、 琐辖 和 伊提南 。
1CHR|4|8|哥斯 生 亚诺 、 琐比巴 和 哈仑 的儿子 亚哈黑 的宗族。
1CHR|4|9|雅比斯 比他众兄弟更尊贵，他母亲给他起名叫 雅比斯 ，意思说：“我生他甚是痛苦。”
1CHR|4|10|雅比斯 求告 以色列 的上帝说：“甚愿你赐福与我，扩张我的疆界，你的手常与我同在，保佑我不遭患难，不受艰苦。”上帝就应允他所求的。
1CHR|4|11|书哈 的兄弟 基绿 生 米黑 ， 米黑 是 伊施屯 的父亲。
1CHR|4|12|伊施屯 生 伯拉巴 、 巴西亚 和 珥．拿辖 之祖 提欣拿 。这些都是 利迦 人。
1CHR|4|13|基纳斯 的儿子是 俄陀聂 和 西莱雅 。 俄陀聂 的儿子是 哈塔 。
1CHR|4|14|悯挪太 生 俄弗拉 ； 西莱雅 生 革．夏纳欣 之祖 约押 。他们都是工匠。
1CHR|4|15|耶孚尼 的儿子 迦勒 的后裔： 以路 、 以拉 和 拿安 。 以拉 的儿子是 基纳斯 。
1CHR|4|16|耶哈利勒 的儿子是 西弗 、 西法 、 提利 和 亚撒列 。
1CHR|4|17|以斯拉 的儿子是 益帖 、 米列 、 以弗 和 雅伦 。 米列 所娶法老的女儿 比提雅 的后裔如下：她怀了 米利暗 、 沙买 ，和 以实提摩 之祖 益巴 。 米列 的 犹大 妻子生 基多 之祖 雅列 ， 梭哥 之祖 希伯 ，和 撒挪亚 之祖 耶古铁 。
1CHR|4|18|
1CHR|4|19|拿含 的妹妹， 荷第雅 的妻子所生的是 达利亚 ， 迦米 人 基伊拉 和 玛迦 人 以实提摩 的祖先。
1CHR|4|20|示门 的儿子是 暗嫩 、 林拿 、 便．哈南 和 提伦 。 以示 的儿子是 梭黑 和 便．梭黑 。
1CHR|4|21|犹大 的儿子 示拉 的后裔： 利迦 之祖 珥 ， 玛利沙 之祖 拉大 ，和住在 伯．亚实比 织细麻布的各宗族。
1CHR|4|22|还有 约敬 、 哥西巴 人、 约阿施 ，和那在 摩押 娶妻，回到 利恒 的 萨拉 。这都是古时的记载。
1CHR|4|23|这些人都是陶匠，是 尼他应 和 基底拉 的居民。他们住在王那里，为王做工。
1CHR|4|24|西缅 的后裔如下： 尼母利 、 雅悯 、 雅立 、 谢拉 和 扫罗 ；
1CHR|4|25|他的儿子 沙龙 ，他的儿子 米比衫 ，他的儿子 米施玛 ；
1CHR|4|26|米施玛 的后裔：他的儿子 哈母利 ，他的儿子 撒刻 ，他的儿子 示每 。
1CHR|4|27|示每 有十六个儿子和六个女儿，但他兄弟的儿女不多，他们各家族也不如 犹大 族那样人丁兴旺。
1CHR|4|28|西缅 人住在 别是巴 、 摩拉大 、 哈萨．书亚 、
1CHR|4|29|辟拉 、 以森 、 陀腊 、
1CHR|4|30|彼土利 、 何珥玛 、 洗革拉 、
1CHR|4|31|伯．玛加博 、 哈萨．苏撒 、 伯．比利 和 沙拉音 ，这些城镇直到 大卫 作王的时候都是属 西缅 人的；
1CHR|4|32|还有所属的村庄 以坦 、 亚因 、 临门 、 陀健 、 亚珊 ，共五个城镇；
1CHR|4|33|连同环绕这些城镇的一切乡村，直到 巴力 。这是他们的住处，他们都有家谱。
1CHR|4|34|还有 米所巴 、 雅米勒 、 亚玛谢 的儿子 约沙 、
1CHR|4|35|约珥 ，和 亚薛 的曾孙， 西莱雅 的孙子， 约示比 的儿子 耶户 。
1CHR|4|36|还有 以利约乃 、 雅哥巴 、 约朔海 、 亚帅雅 、 亚底业 、 耶西篾 、 比拿雅 、
1CHR|4|37|细撒 ； 细撒 是 示非 的儿子， 示非 是 亚龙 的儿子， 亚龙 是 耶大雅 的儿子， 耶大雅 是 申利 的儿子， 申利 是 示玛雅 的儿子。
1CHR|4|38|以上所记的人名都是作族长的，他们父系的家属大量增加。
1CHR|4|39|他们往平原东边 基多口 去，寻找牧放羊群的草场，
1CHR|4|40|找到了肥沃优美的草场，又宽阔又平静安宁之地；从前住那里的是 含 族的人。
1CHR|4|41|以上纪录上有名的人，在 犹大 王 希西家 的日子，来攻击 含 族人的帐棚和那里所有的 米乌尼 人，把他们灭尽，就住在他们的地方，直到今日，因为那里有草场可以牧放羊群。
1CHR|4|42|这些 西缅 人中有五百人上 西珥山 ，率领他们的是 以示 的儿子 毗拉提 、 尼利雅 、 利法雅 和 乌薛 。
1CHR|4|43|他们杀了 亚玛力 剩下的残存之民，就住在那里，直到今日。
1CHR|5|1|以色列 的长子 吕便 的后裔。 吕便 玷污了父亲的床，他长子的名分就归了 以色列 的儿子 约瑟 的后裔；因此，家谱就不按出生顺序登录。
1CHR|5|2|虽然 犹大 比他兄弟强盛，君王也从他而出，然而长子的名分却归 约瑟 。
1CHR|5|3|以色列 长子 吕便 的后裔如下： 哈诺 、 法路 、 希斯伦 和 迦米 。
1CHR|5|4|约珥 的后裔：他的儿子 示玛雅 ，他的儿子 歌革 ，他的儿子 示每 ，
1CHR|5|5|他的儿子 米迦 ，他的儿子 利亚雅 ，他的儿子 巴力 ，
1CHR|5|6|他的儿子 备拉 ；这 备拉 作 吕便 支派的领袖，被 亚述 王 提革拉．毗列色 掳去。
1CHR|5|7|他的弟兄照着宗族，按着家谱作族长的是 耶利 、 撒迦利雅 、
1CHR|5|8|比拉 ； 比拉 是 亚撒 的儿子， 亚撒 是 示玛 的儿子， 示玛 是 约珥 的儿子； 约珥 住在 亚罗珥 ，直到 尼波 和 巴力．免 。
1CHR|5|9|他也住在东边，直到 幼发拉底河 这边的旷野边界，因为他们在 基列 地牲畜增多。
1CHR|5|10|扫罗 年间，他们与 夏甲 人争战， 夏甲 人倒在他们手下，他们就在 基列 东边的全地，住在 夏甲 人的帐棚里。
1CHR|5|11|迦得 的后裔在 吕便 对面，住在 巴珊 地，延伸到 撒迦 ：
1CHR|5|12|有作族长的 约珥 ，有作副族长的 沙番 ，还有 雅乃 和住在 巴珊 的 沙法 。
1CHR|5|13|按着家族，他们的弟兄是 米迦勒 、 米书兰 、 示巴 、 约赖 、 雅干 、 细亚 和 希伯 ，共七人。
1CHR|5|14|这些都是 亚比孩 的儿子； 亚比孩 是 户利 的儿子， 户利 是 耶罗亚 的儿子， 耶罗亚 是 基列 的儿子， 基列 是 米迦勒 的儿子， 米迦勒 是 耶示筛 的儿子， 耶示筛 是 耶哈多 的儿子， 耶哈多 是 布斯 的儿子；
1CHR|5|15|古尼 的孙子， 押比叠 的儿子 亚希 是他们的族长。
1CHR|5|16|他们住在 基列 、 巴珊 和所属的乡镇，以及 沙仑 一切的郊野，直到四围的交界。
1CHR|5|17|这些人在 犹大 王 约坦 和 以色列 王 耶罗波安 年间，都载入家谱。
1CHR|5|18|吕便 人、 迦得 人和 玛拿西 半支派的人，能拿盾牌和刀剑、拉弓、出征善战的勇士共有四万四千七百六十名。
1CHR|5|19|他们与 夏甲 人、 伊突 人、 拿非施 人、 挪答 人打仗。
1CHR|5|20|他们在打仗的时候得了上帝的帮助， 夏甲 人和所有跟随 夏甲 人的人都交在他们手中；因为他们在阵上呼求上帝，倚赖他，他就应允他们。
1CHR|5|21|他们掳掠了 夏甲 人的牲畜，有五万匹骆驼，二十五万只羊，二千匹驴，又有十万人；
1CHR|5|22|被杀仆倒的很多，因为这战争是出乎上帝。他们就住在 夏甲 人的地上，直到被掳的时候。
1CHR|5|23|玛拿西 半支派的人住在那地，从 巴珊 延到 巴力．黑门 、 示尼珥 和 黑门山 ，他们人数增多 。
1CHR|5|24|他们的族长如下： 以弗 、 以示 、 以利业 、 亚斯列 、 耶利米 、 何达威雅 和 雅叠 ；他们都是大能的勇士，有名的人，是作族长的。
1CHR|5|25|但他们得罪了他们列祖的上帝，随从当地百姓的神明而行淫，这百姓就是上帝在他们面前所除灭的。
1CHR|5|26|因此， 以色列 的上帝激发 亚述 王 普勒 ，就是 亚述 王 提革拉．毗列色 的心，他掳掠了 吕便 人、 迦得 人、 玛拿西 半支派的人，把他们带到 哈腊 、 哈博 、 哈拉 与 歌散河 边，直到今日。
1CHR|6|1|利未 的后裔： 革顺 、 哥辖 和 米拉利 。
1CHR|6|2|哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 和 乌薛 。
1CHR|6|3|暗兰 的儿女是 亚伦 、 摩西 和 米利暗 。 亚伦 的儿子是 拿答 、 亚比户 、 以利亚撒 和 以他玛 。
1CHR|6|4|以利亚撒 生 非尼哈 ； 非尼哈 生 亚比书 ；
1CHR|6|5|亚比书 生 布基 ； 布基 生 乌西 ；
1CHR|6|6|乌西 生 西拉希雅 ； 西拉希雅 生 米拉约 ；
1CHR|6|7|米拉约 生 亚玛利雅 ； 亚玛利雅 生 亚希突 ；
1CHR|6|8|亚希突 生 撒督 ； 撒督 生 亚希玛斯 ；
1CHR|6|9|亚希玛斯 生 亚撒利雅 ； 亚撒利雅 生 约哈难 ；
1CHR|6|10|约哈难 生 亚撒利雅 ， 亚撒利雅 在 所罗门 建造的 耶路撒冷 殿中担任祭司的职分；
1CHR|6|11|亚撒利雅 生 亚玛利雅 ； 亚玛利雅 生 亚希突 ；
1CHR|6|12|亚希突 生 撒督 ； 撒督 生 沙龙 ；
1CHR|6|13|沙龙 生 希勒家 ； 希勒家 生 亚撒利雅 ；
1CHR|6|14|亚撒利雅 生 西莱雅 ； 西莱雅 生 约萨答 。
1CHR|6|15|当耶和华藉 尼布甲尼撒 的手掳掠 犹大 和 耶路撒冷 的时候， 约萨答 也被掳去。
1CHR|6|16|利未 的后裔： 革顺 、 哥辖 和 米拉利 。
1CHR|6|17|革顺 的儿子名叫 立尼 和 示每 。
1CHR|6|18|哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 和 乌薛 。
1CHR|6|19|米拉利 的儿子是 抹利 和 母示 。这是按着父系所分 利未 人的宗族。
1CHR|6|20|属 革顺 的：他的儿子 立尼 ，他的儿子 雅哈 ，他的儿子 薪玛 ，
1CHR|6|21|他的儿子 约亚 ，他的儿子 易多 ，他的儿子 谢拉 ，他的儿子 耶特赖 。
1CHR|6|22|哥辖 的后裔：他的儿子 亚米拿达 ，他的儿子 可拉 ，他的儿子 亚惜 ，
1CHR|6|23|他的儿子 以利加拿 ，他的儿子 以比雅撒 ，他的儿子 亚惜 ，
1CHR|6|24|他的儿子 他哈 ，他的儿子 乌列 ，他的儿子 乌西雅 ，他的儿子 少罗 。
1CHR|6|25|以利加拿 的儿子是 亚玛赛 、 亚希摩 、
1CHR|6|26|以利加拿 。 以利加拿 的后裔：他的儿子 琐菲 ，他的儿子 拿哈 ，
1CHR|6|27|他的儿子 以利押 ，他的儿子 耶罗罕 ，他的儿子 以利加拿 ，他的儿子 撒母耳 。
1CHR|6|28|撒母耳 的儿子是长子 约珥 和次子 亚比亚 。
1CHR|6|29|米拉利 的后裔： 抹利 ，他的儿子 立尼 ，他的儿子 示每 ，他的儿子 乌撒 ，
1CHR|6|30|他的儿子 示米亚 ，他的儿子 哈基雅 ，他的儿子 亚帅雅 。
1CHR|6|31|这些是约柜安设之后， 大卫 派在耶和华殿中管理歌唱事奉的人。
1CHR|6|32|他们在会幕前负责歌唱的事奉，及至 所罗门 在 耶路撒冷 建造了耶和华的殿，他们就按着班次供职。
1CHR|6|33|供职的人和他们的子孙如下： 哥辖 的子孙中有歌唱的 希幔 ； 希幔 是 约珥 的儿子， 约珥 是 撒母耳 的儿子，
1CHR|6|34|撒母耳 是 以利加拿 的儿子， 以利加拿 是 耶罗罕 的儿子， 耶罗罕 是 以利业 的儿子， 以利业 是 陀亚 的儿子，
1CHR|6|35|陀亚 是 苏弗 的儿子， 苏弗 是 以利加拿 的儿子， 以利加拿 是 玛哈 的儿子， 玛哈 是 亚玛赛 的儿子，
1CHR|6|36|亚玛赛 是 以利加拿 的儿子， 以利加拿 是 约珥 的儿子， 约珥 是 亚撒利雅 的儿子， 亚撒利雅 是 西番雅 的儿子，
1CHR|6|37|西番雅 是 他哈 的儿子， 他哈 是 亚惜 的儿子， 亚惜 是 以比雅撒 的儿子， 以比雅撒 是 可拉 的儿子，
1CHR|6|38|可拉 是 以斯哈 的儿子， 以斯哈 是 哥辖 的儿子， 哥辖 是 利未 的儿子， 利未 是 以色列 的儿子。
1CHR|6|39|希幔 的弟兄 亚萨 在 希幔 的右边供职； 亚萨 是 比利家 的儿子， 比利家 是 示米亚 的儿子，
1CHR|6|40|示米亚 是 米迦勒 的儿子， 米迦勒 是 巴西雅 的儿子， 巴西雅 是 玛基雅 的儿子，
1CHR|6|41|玛基雅 是 伊特尼 的儿子， 伊特尼 是 谢拉 的儿子， 谢拉 是 亚大雅 的儿子，
1CHR|6|42|亚大雅 是 以探 的儿子， 以探 是 薪玛 的儿子， 薪玛 是 示每 的儿子，
1CHR|6|43|示每 是 雅哈 的儿子， 雅哈 是 革顺 的儿子， 革顺 是 利未 的儿子。
1CHR|6|44|他们的弟兄 米拉利 的子孙，在他们左边供职的有 以探 ； 以探 是 基示 的儿子， 基示 是 亚伯底 的儿子， 亚伯底 是 玛鹿 的儿子，
1CHR|6|45|玛鹿 是 哈沙比雅 的儿子， 哈沙比雅 是 亚玛谢 的儿子， 亚玛谢 是 希勒家 的儿子，
1CHR|6|46|希勒家 是 暗西 的儿子， 暗西 是 巴尼 的儿子， 巴尼 是 沙麦 的儿子，
1CHR|6|47|沙麦 是 末力 的儿子， 末力 是 母示 的儿子， 母示 是 米拉利 的儿子， 米拉利 是 利未 的儿子。
1CHR|6|48|他们的弟兄 利未 人也被派办理上帝殿中帐幕的一切事务。
1CHR|6|49|亚伦 和他的子孙在燔祭坛和香坛上献祭烧香，办理至圣所一切的事，为 以色列 赎罪，正如上帝仆人 摩西 所吩咐的一切。
1CHR|6|50|亚伦 的后裔如下：他的儿子 以利亚撒 ，他的儿子 非尼哈 ，他的儿子 亚比书 ，
1CHR|6|51|他的儿子 布基 ，他的儿子 乌西 ，他的儿子 西拉希雅 ，
1CHR|6|52|他的儿子 米拉约 ，他的儿子 亚玛利雅 ，他的儿子 亚希突 ，
1CHR|6|53|他的儿子 撒督 ，他的儿子 亚希玛斯 。
1CHR|6|54|他们的住处按着境内的营寨如下： 亚伦 的子孙 哥辖 族先抽签得地，
1CHR|6|55|得了 犹大 地的 希伯仑 和四围的郊野；
1CHR|6|56|只是这城的田地和所属的村庄都为 耶孚尼 的儿子 迦勒 所得。
1CHR|6|57|亚伦 的子孙所得逃城如下： 希伯仑 、 立拿 与其郊野、 雅提珥 、 以实提莫 与其郊野、
1CHR|6|58|希仑 与其郊野、 底璧 与其郊野、
1CHR|6|59|亚珊 与其郊野、 伯．示麦 与其郊野。
1CHR|6|60|他们也从 便雅悯 支派中得了 迦巴 与其郊野、 阿勒篾 与其郊野、 亚拿突 与其郊野。他们宗族所得的城共十三座。
1CHR|6|61|哥辖 族其余的人抽签，按支派的宗族，从半个支派，就是 玛拿西 半支派中得了十座城。
1CHR|6|62|革顺 族按着宗族，从 以萨迦 支派、 亚设 支派、 拿弗他利 支派、 巴珊 内的 玛拿西 支派中，得了十三座城。
1CHR|6|63|米拉利 族按着宗族抽签，从 吕便 支派、 迦得 支派、 西布伦 支派中，得了十二座城。
1CHR|6|64|以色列 人把这些城与其郊野给了 利未 人。
1CHR|6|65|以色列 人用抽签的方式，从 犹大 人、 西缅 人、 便雅悯 人三支派中，把以上提到名字的城给了他们。
1CHR|6|66|哥辖 子孙中有几个宗族从 以法莲 支派中也得了城镇作为他们的区域。
1CHR|6|67|他们在 以法莲 山区所得的逃城： 示剑 与其郊野、 基色 与其郊野、
1CHR|6|68|约缅 与其郊野、 伯．和仑 与其郊野、
1CHR|6|69|亚雅仑 与其郊野、 迦特．临门 与其郊野。
1CHR|6|70|哥辖 其余的子孙从 玛拿西 半支派中得了 亚乃 与其郊野、 比连 与其郊野。
1CHR|6|71|革顺 子孙从 玛拿西 半支派中得了 巴珊 的 哥兰 与其郊野、 亚斯她录 与其郊野；
1CHR|6|72|从 以萨迦 支派中得了 基低斯 与其郊野、 大比拉 与其郊野、
1CHR|6|73|拉末 与其郊野、 亚年 与其郊野；
1CHR|6|74|从 亚设 支派中得了 玛沙 与其郊野、 押顿 与其郊野、
1CHR|6|75|户割 与其郊野、 利合 与其郊野；
1CHR|6|76|从 拿弗他利 支派中得了 加利利 的 基低斯 与其郊野、 哈们 与其郊野、 基列亭 与其郊野。
1CHR|6|77|米拉利 其余的子孙从 西布伦 支派中得了 临摩挪 与其郊野、 他泊 与其郊野；
1CHR|6|78|又在 耶利哥 的 约旦河 东，从 吕便 支派中得了旷野的 比悉 与其郊野、 雅杂 与其郊野，
1CHR|6|79|基底莫 与其郊野、 米法押 与其郊野；
1CHR|6|80|又从 迦得 支派中得了 基列 的 拉末 与其郊野、 玛哈念 与其郊野、
1CHR|6|81|希实本 与其郊野、 雅谢 与其郊野。
1CHR|7|1|以萨迦 的后裔： 陀拉 、 普瓦 、 雅述 和 伸仑 ，共四人。
1CHR|7|2|陀拉 的后裔： 乌西 、 利法雅 、 耶勒 、 雅买 、 易伯散 和 示母利 ，都是 陀拉 的族长，在他们世代中是大能的勇士。到 大卫 年间，他们的人数共有二万二千六百名。
1CHR|7|3|乌西 的后裔： 伊斯拉希 ， 伊斯拉希 的儿子 米迦勒 、 俄巴底亚 、 约珥 和 伊示雅 ，共五人，全都是族长。
1CHR|7|4|他们所率领的，按着家谱，照着父家，可作战的军队共有三万六千人，因为他们的妻子和儿子众多。
1CHR|7|5|他们的弟兄在 以萨迦 各族中的大能勇士，登记在家谱中的全部共有八万七千人。
1CHR|7|6|便雅悯 ： 比拉 、 比结 和 耶叠 ，共三人。
1CHR|7|7|比拉 的儿子： 以斯本 、 乌西 、 乌薛 、 耶利末 和 以利 ，共五人，都是族长，是大能的勇士。登记在家谱中的人共有二万二千零三十四人。
1CHR|7|8|比结 的儿子： 细米拉 、 约阿施 、 以利以谢 、 以利约乃 、 暗利 、 耶列末 、 亚比雅 、 亚拿突 和 亚拉篾 ；这些全都是 比结 的儿子。
1CHR|7|9|登记在家谱中，按家谱的族长，大能的勇士，共有二万零二百人。
1CHR|7|10|耶叠 的后裔： 比勒罕 ， 比勒罕 的儿子 耶乌施 、 便雅悯 、 以笏 、 基拿拿 、 细坦 、 他施 和 亚希沙哈 。
1CHR|7|11|这些全都是 耶叠 的后裔，都是族长，是大能的勇士，能上阵打仗的共有一万七千二百人。
1CHR|7|12|还有 以珥 的儿子 书品 和 户品 ，以及 亚黑 的儿子 户伸 。
1CHR|7|13|拿弗他利 的后裔： 雅薛 、 沽尼 、 耶色 和 沙龙 ，都是 辟拉 的子孙。
1CHR|7|14|玛拿西 的儿子 亚斯烈 是他的妾 亚兰 女子所生的；她又生了 玛吉 ，是 基列 的父亲。
1CHR|7|15|玛吉 为 户品 和 书品 各娶了一妻，他的姊妹名叫 玛迦 。第二个名叫 西罗非哈 ； 西罗非哈 只有女儿。
1CHR|7|16|玛吉 的妻子 玛迦 生了一个儿子， 玛迦 给他起名叫 毗利施 。 毗利施 的弟弟名叫 示利施 ； 示利施 的儿子是 乌兰 和 利金 。
1CHR|7|17|乌兰 的儿子是 比但 。这些都是 基列 的子孙； 基列 是 玛吉 的儿子， 玛吉 是 玛拿西 的儿子。
1CHR|7|18|基列 的妹妹 哈摩利吉 生了 伊施荷 、 亚比以谢 和 玛拉 。
1CHR|7|19|示米大 的儿子是 亚现 、 示剑 、 利克希 和 阿尼安 。
1CHR|7|20|以法莲 的后裔： 书提拉 ，他的儿子 比列 ，他的儿子 他哈 ，他的儿子 以拉大 ，他的儿子 他哈 ，
1CHR|7|21|他的儿子 撒拔 ，他的儿子 书提拉 。 以法莲 又生 以谢 和 以列 ；这二人因为下去夺取 迦特 人的牲畜，被本地的 迦特 人杀了。
1CHR|7|22|他们的父亲 以法莲 为他们悲哀了多日，他的兄弟都来安慰他。
1CHR|7|23|以法莲 与妻子同房，妻子怀孕生了一子， 以法莲 因为家里遭祸，就给这儿子起名叫 比利亚 。
1CHR|7|24|他的女儿名叫 舍伊拉 ， 舍伊拉 建筑了 上伯．和仑 、 下伯．和仑 和 乌羡．舍伊拉 。
1CHR|7|25|他的儿子 利法 和 利悉 ，他的儿子 他拉 ，他的儿子 他罕 ，
1CHR|7|26|他的儿子 拉但 ，他的儿子 亚米忽 ，他的儿子 以利沙玛 ，
1CHR|7|27|他的儿子 嫩 ，他的儿子 约书亚 。
1CHR|7|28|以法莲 人的地业和住处是 伯特利 和所属的乡镇，东边 拿兰 ，西边 基色 和所属的乡镇， 示剑 和所属的乡镇，直到 艾雅 和所属的乡镇；
1CHR|7|29|还有靠近 玛拿西 人的边界， 伯．善 和所属的乡镇， 他纳 和所属的乡镇， 米吉多 和所属的乡镇， 多珥 和所属的乡镇。 以色列 儿子 约瑟 的子孙住在这些地方。
1CHR|7|30|亚设 的后裔： 音拿 、 亦施瓦 、 亦施韦 和 比利亚 ，还有他们的妹妹 西拉 。
1CHR|7|31|比利亚 的儿子是 希别 和 玛结 ； 玛结 是 比撒威 的父亲。
1CHR|7|32|希别 生 雅弗勒 、 朔默 、 何坦 和他们的妹妹 书雅 。
1CHR|7|33|雅弗勒 的儿子是 巴萨 、 宾哈 和 亚施法 ；这些都是 雅弗勒 的儿子。
1CHR|7|34|朔默 的儿子是 亚希 、 罗迦 、 耶户巴 和 亚兰 。
1CHR|7|35|朔默 的兄弟 希连 的儿子是 琐法 、 音那 、 示利斯 和 亚抹 。
1CHR|7|36|琐法 的儿子是 书亚 、 哈尼弗 、 书阿勒 、 比利 、 音拉 、
1CHR|7|37|比悉 、 河得 、 珊玛 、 施沙 、 益兰 和 比拉 。
1CHR|7|38|益帖 的儿子是 耶孚尼 、 毗斯巴 和 亚拉 。
1CHR|7|39|乌拉 的儿子是 亚拉 、 汉尼业 和 利写 。
1CHR|7|40|这些全都是 亚设 的子孙，都是族长，是精壮大能的勇士，也是领袖中的领袖。登记在家谱中，能上阵打仗的共有二万六千人。
1CHR|8|1|便雅悯 生长子 比拉 ，次子 亚实别 ，三子 亚哈拉 ，
1CHR|8|2|四子 挪哈 ，五子 拉法 。
1CHR|8|3|比拉 的儿子是 亚大 、 基拉 、 亚比忽 、
1CHR|8|4|亚比书 、 乃幔 、 亚何亚 、
1CHR|8|5|基拉 、 示孚汛 和 户兰 。
1CHR|8|6|以忽 的后裔如下，他们是 迦巴 居民的族长，曾被掳到 玛拿辖 ：
1CHR|8|7|乃幔 、 亚希亚 、 基拉 ；他掳了他们，又生了 乌撒 和 亚希忽 。
1CHR|8|8|沙哈连 休了两个妻子 户伸 和 巴拉 之后，在 摩押 地生了儿子。
1CHR|8|9|他与妻子 贺得 生了 约巴 、 洗比雅 、 米沙 、 玛拉干 、
1CHR|8|10|耶乌斯 、 沙迦 和 米玛 ；这些是他的儿子，都是族长。
1CHR|8|11|户伸 为他生了 亚比突 和 以利巴力 。
1CHR|8|12|以利巴力 的儿子是 希伯 、 米珊 和 沙麦 ； 沙麦 建立 阿挪 、 罗德 和所属的乡镇。
1CHR|8|13|比利亚 和 示玛 是 亚雅仑 居民的族长，他们驱逐了 迦特 的居民。
1CHR|8|14|亚希约 、 沙煞 、 耶列末 、
1CHR|8|15|西巴第雅 、 亚拉得 、 亚得 、
1CHR|8|16|米迦勒 、 伊施巴 和 约哈 都是 比利亚 的儿子。
1CHR|8|17|西巴第雅 、 米书兰 、 希西基 、 希伯 、
1CHR|8|18|伊施米莱 、 伊斯利亚 和 约巴 都是 以利巴力 的儿子。
1CHR|8|19|雅金 、 细基利 、 撒底 、
1CHR|8|20|以利乃 、 洗勒太 、 以利业 、
1CHR|8|21|亚大雅 、 比拉雅 和 申拉 都是 示每 的儿子。
1CHR|8|22|伊施班 、 希伯 、 以利业 、
1CHR|8|23|亚伯顿 、 细基利 、 哈难 、
1CHR|8|24|哈拿尼雅 、 以拦 、 安陀提雅 、
1CHR|8|25|伊弗底雅 、 毗努伊勒 都是 沙煞 的儿子。
1CHR|8|26|珊示莱 、 示哈利 、 亚他利雅 、
1CHR|8|27|雅利西 、 以利亚 和 细基利 都是 耶罗罕 的儿子。
1CHR|8|28|这些人按照他们的家谱都是族长，是领袖，都住在 耶路撒冷 。
1CHR|8|29|在 基遍 住的有 基遍 的父亲 耶利 ，他的妻子名叫 玛迦 ；
1CHR|8|30|他的长子是 亚伯顿 ，还有 苏珥 、 基士 、 巴力 、 拿答 、
1CHR|8|31|基多 、 亚希约 和 撒迦 。
1CHR|8|32|米基罗 生 示米暗 。这些人在他们弟兄的对面，和他们的弟兄同住在 耶路撒冷 。
1CHR|8|33|尼珥 生 基士 ； 基士 生 扫罗 ； 扫罗 生 约拿单 、 麦基．舒亚 、 亚比拿达 和 伊施巴力 。
1CHR|8|34|约拿单 的儿子是 米力．巴力 ； 米力．巴力 生 米迦 。
1CHR|8|35|米迦 的儿子是 毗敦 、 米勒 、 他利亚 和 亚哈斯 ；
1CHR|8|36|亚哈斯 生 耶何阿达 ； 耶何阿达 生 亚拉篾 、 亚斯玛威 和 心利 ； 心利 生 摩撒 ；
1CHR|8|37|摩撒 生 比尼亚 ； 比尼亚 的儿子是 拉法 ， 拉法 的儿子是 以利亚萨 ， 以利亚萨 的儿子是 亚悉 。
1CHR|8|38|亚悉 有六个儿子，他们的名字是 亚斯利干 、 波基路 、 以实玛利 、 示亚利雅 、 俄巴底雅 和 哈难 ；这些全都是 亚悉 的儿子。
1CHR|8|39|亚悉 兄弟 以设 的儿子：长子是 乌兰 ，次子是 耶乌施 ，三子是 以利法列 。
1CHR|8|40|乌兰 的儿子都是大能的勇士，是弓箭手，他们有许多的子孙，共一百五十名，都是 便雅悯 人。
1CHR|9|1|以色列 众人按家谱登记，看哪，都写在《以色列诸王记》上。 犹大 人因背叛被掳到 巴比伦 。
1CHR|9|2|从 巴比伦 先回来，住在自己地业城镇中的有 以色列 人、祭司、 利未 人和殿役。
1CHR|9|3|住在 耶路撒冷 的有 犹大 人、 便雅悯 人、 以法莲 人和 玛拿西 人：
1CHR|9|4|犹大 儿子 法勒斯 的子孙中有 乌太 ， 乌太 是 亚米忽 的儿子， 亚米忽 是 暗利 的儿子， 暗利 是 音利 的儿子， 音利 是 巴尼 的儿子；
1CHR|9|5|示罗 人中有长子 亚帅雅 和他的众儿子；
1CHR|9|6|谢拉 的子孙中有 耶乌利 和他的弟兄，共六百九十人；
1CHR|9|7|便雅悯 人中有 哈西努亚 的曾孙， 何达威雅 的孙子， 米书兰 的儿子 撒路 ；
1CHR|9|8|又有 耶罗罕 的儿子 伊比内雅 ； 米基立 的孙子， 乌西 的儿子 以拉 ； 伊比尼雅 的曾孙， 流珥 的孙子， 示法提雅 的儿子 米书兰 ；
1CHR|9|9|和他们的弟兄，按着家谱登记，共有九百五十六名；这些人都是族长。
1CHR|9|10|祭司中有 耶大雅 、 耶何雅立 、 雅斤 ，
1CHR|9|11|还有管理上帝殿的 亚撒利雅 ， 亚撒利雅 是 希勒家 的儿子， 希勒家 是 米书兰 的儿子， 米书兰 是 撒督 的儿子， 撒督 是 米拉约 的儿子， 米拉约 是 亚希突 的儿子。
1CHR|9|12|还有 玛基雅 的曾孙， 巴施户珥 的孙子， 耶罗罕 的儿子 亚大雅 ；又有 玛赛 ， 玛赛 是 亚第业 的儿子， 亚第业 是 雅希细拉 的儿子， 雅希细拉 是 米书兰 的儿子， 米书兰 是 米实利密 的儿子， 米实利密 是 音麦 的儿子。
1CHR|9|13|他们和他们的弟兄都是族长，共有一千七百六十人，都善于做上帝殿的事工。
1CHR|9|14|利未 人 米拉利 的子孙中有 哈沙比雅 的曾孙， 押利甘 的孙子， 哈述 的儿子 示玛雅 ；
1CHR|9|15|有 拔巴甲 、 黑勒施 、 加拉 和 亚萨 的曾孙， 细基利 的孙子， 米迦 的儿子 玛探雅 ；
1CHR|9|16|又有 耶杜顿 的曾孙， 加拉 的孙子， 示玛雅 的儿子 俄巴底 ，还有 以利加拿 的孙子， 亚撒 的儿子 比利家 。他们都住在 尼陀法 人的村庄。
1CHR|9|17|守卫是 沙龙 、 亚谷 、 达们 、 亚希幔 和他们的弟兄； 沙龙 是领袖。
1CHR|9|18|从前这些人看守朝东的王门，如今是 利未 人营中的守卫。
1CHR|9|19|可拉 的曾孙， 以比雅撒 的孙子， 可利 的儿子 沙龙 ，和他父家的弟兄 可拉 人管理事务，看守会幕的门。他们的祖宗曾管理耶和华的军营，把守营的入口。
1CHR|9|20|从前 以利亚撒 的儿子 非尼哈 管理他们，耶和华也与他同在。
1CHR|9|21|米施利米雅 的儿子 撒迦利雅 是看守会幕门口的。
1CHR|9|22|被选作门口守卫的总共有二百一十二名。他们在自己的村庄，按着家谱登记，是 大卫 和 撒母耳 先见所派担当这受托之职任的。
1CHR|9|23|他们和他们的子孙看守耶和华殿的门，就是会幕的门口。
1CHR|9|24|在东西南北，四方 都有守卫。
1CHR|9|25|他们的弟兄住在村庄，每七日来与他们换班。
1CHR|9|26|这些守卫的四个领袖都是 利未 人，各有受托的职任，看守上帝殿的房间和宝库。
1CHR|9|27|他们住在上帝殿的四围，受托看守圣殿，负责每日早晨开门。
1CHR|9|28|利未 人中有人管理所使用的器皿，拿出拿入都按数目点算。
1CHR|9|29|又有人管理器具和圣所一切的器皿，以及细面、酒、油、乳香和香料。
1CHR|9|30|祭司的子孙中有人用香料做膏油。
1CHR|9|31|利未 人 玛他提雅 是 可拉 族 沙龙 的长子，他受托做烤饼。
1CHR|9|32|他们弟兄 哥辖 子孙中，有人负责每安息日排列供饼。
1CHR|9|33|歌唱的有 利未 人的族长，住在殿的房间，昼夜供职，不做别样的工。
1CHR|9|34|以上都是 利未 人的族长，按各世系作领袖，他们都住在 耶路撒冷 。
1CHR|9|35|在 基遍 住的有 基遍 的父亲 耶利 ，他的妻子名叫 玛迦 ；
1CHR|9|36|他的长子是 亚伯顿 ，还有 苏珥 、 基士 、 巴力 、 尼珥 、 拿答 、
1CHR|9|37|基多 、 亚希约 、 撒迦利雅 和 米基罗 。
1CHR|9|38|米基罗 生 示米暗 。这些人在他们弟兄的对面，和他们的弟兄同住在 耶路撒冷 。
1CHR|9|39|尼珥 生 基士 ； 基士 生 扫罗 ； 扫罗 生 约拿单 、 麦基．舒亚 、 亚比拿达 和 伊施巴力 。
1CHR|9|40|约拿单 的儿子是 米力．巴力 ； 米力．巴力 生 米迦 。
1CHR|9|41|米迦 的儿子是 毗敦 、 米勒 、 他利亚 和 亚哈斯 。
1CHR|9|42|亚哈斯 生 雅拉 ； 雅拉 生 亚拉篾 、 亚斯玛威 和 心利 ； 心利 生 摩撒 ；
1CHR|9|43|摩撒 生 比尼亚 ； 比尼亚 的儿子是 利法雅 ， 利法雅 的儿子是 以利亚萨 ， 以利亚萨 的儿子是 亚悉 。
1CHR|9|44|亚悉 有六个儿子，他们的名字是 亚斯利干 、 波基路 、 以实玛利 、 示亚利雅 、 俄巴底雅 和 哈难 ；这些都是 亚悉 的儿子。
1CHR|10|1|非利士 人攻打 以色列 。 以色列 人在 非利士 人面前逃跑，很多人 在 基利波山 被杀仆倒。
1CHR|10|2|非利士 人紧追 扫罗 和他的儿子，杀了 扫罗 的儿子 约拿单 、 亚比拿达 、 麦基．舒亚 。
1CHR|10|3|攻击 扫罗 的战事激烈， 扫罗 被弓箭手射中，被他们射伤。
1CHR|10|4|扫罗 吩咐拿他兵器的人说：“你拔出刀来，把我刺死，免得那些未受割礼的人来凌辱我。”但拿兵器的人非常惧怕，不肯刺他。于是 扫罗 拿起刀来，伏在刀上。
1CHR|10|5|拿兵器的人见 扫罗 已死，也伏在刀上死了。
1CHR|10|6|这样， 扫罗 和他三个儿子，以及他的全家都一起阵亡了。
1CHR|10|7|住平原的 以色列 众人见 以色列 军兵 逃跑， 扫罗 和他儿子都死了，就弃城逃跑。 非利士 人前来，占据了他们的城。
1CHR|10|8|次日， 非利士 人来剥那些被杀之人的衣服，看见 扫罗 和他儿子仆倒在 基利波山 。
1CHR|10|9|他们剥了他的军装，拿着他的首级和盔甲，派人到 非利士 人之地的四境，报信给他们的偶像和百姓。
1CHR|10|10|他们将 扫罗 的盔甲放在他们神明的庙里，把他的首级钉在 大衮 庙中。
1CHR|10|11|基列 的 雅比 居民听见 非利士 人向 扫罗 所行的一切事，
1CHR|10|12|他们中间所有的勇士就起身，把 扫罗 和他儿子的尸身送到 雅比 ，把他们的尸骨葬在 雅比 的橡树下，禁食七日。
1CHR|10|13|这样， 扫罗 为了他的不忠死了；因为他干犯耶和华，没有遵守耶和华的话，又因他求问招魂的妇人，
1CHR|10|14|不求问耶和华，所以耶和华使他被杀，把王国给了 耶西 的儿子 大卫 。
1CHR|11|1|以色列 众人聚集到 希伯仑 见 大卫 ，说：“看哪，我们是你的骨肉。
1CHR|11|2|从前 扫罗 作王的时候，率领 以色列 人出入的是你；耶和华－你的上帝也曾对你说：‘你必牧养我的百姓 以色列 ，你必作我百姓 以色列 的君王。’”
1CHR|11|3|于是 以色列 的众长老都来到 希伯仑 见王。 大卫 在 希伯仑 ，在耶和华面前与他们立约，他们就膏 大卫 作 以色列 的王，正如耶和华藉 撒母耳 所说的话。
1CHR|11|4|大卫 和 以色列 众人到了 耶路撒冷 ，就是 耶布斯 ；那时 耶布斯 人住在那里。
1CHR|11|5|耶布斯 人对 大卫 说：“你必不能进到这里。”然而 大卫 攻取了 锡安 的堡垒，就是 大卫 的城。
1CHR|11|6|大卫 说：“谁先攻打 耶布斯 人，必作领袖，作元帅。” 洗鲁雅 的儿子 约押 先上去，就作了领袖。
1CHR|11|7|大卫 住在堡垒里，所以那堡垒叫作 大卫城 。
1CHR|11|8|大卫 又从 米罗 起，四围建筑城墙，其余的由 约押 修建。
1CHR|11|9|大卫 日见强大，万军之耶和华与他同在。
1CHR|11|10|以下是跟随 大卫 勇士的领袖；他们奋勇帮助他得到国度，并照着耶和华吩咐 以色列 的话，与 以色列 众人一同立他作王。
1CHR|11|11|大卫 勇士的名单如下： 哈革摩尼 的儿子 雅朔班 ，他是军官的统领 ，曾一次举枪杀了三百人。
1CHR|11|12|其次是 亚何亚 人 朵多 的儿子 以利亚撒 ，他是三个勇士里的一个。
1CHR|11|13|他从前与 大卫 在 巴斯．大悯 ， 非利士 人聚集要打仗。那里有一块长满大麦的田。百姓在 非利士 人面前逃跑，
1CHR|11|14|他们 却站在那块田的中间，防守那田，击败了 非利士 人。耶和华大获全胜。
1CHR|11|15|三十个领袖中的三个人下到磐石那里，进了 亚杜兰洞 见 大卫 ； 非利士 的军队在 利乏音谷 安营。
1CHR|11|16|那时 大卫 在山寨， 非利士 人的驻军在 伯利恒 。
1CHR|11|17|大卫 渴想着说：“但愿有人从 伯利恒 城门旁的井里打水来给我喝！”
1CHR|11|18|这三个勇士就闯过 非利士 人的军营，从 伯利恒 城门旁的井里打水，拿来给 大卫 喝。 大卫 却不肯喝，将水浇在耶和华面前，
1CHR|11|19|说：“我的上帝啊，我绝不做这事！这些人冒死去打水，这水是他们用生命换来的，我怎能喝他们的血呢？” 大卫 不肯喝这水。这是三个勇士所做的事。
1CHR|11|20|约押 的兄弟 亚比筛 是这三个 勇士的领袖；他曾举枪杀了三百人，就在三个勇士中得了名。
1CHR|11|21|他在这三个勇士里比其他两个更有名望，所以作他们的领袖，只是不及前三个勇士。
1CHR|11|22|耶何耶大 的儿子 比拿雅 是来自 甲薛 的勇士，曾行了大事。他杀了 摩押 人 亚利伊勒 的两个儿子，又在下雪的时候下到坑里去，杀了一只狮子。
1CHR|11|23|他又杀了一个身高五肘的 埃及 人； 埃及 人手里拿着枪，枪杆粗如织布机的轴。 比拿雅 只拿着棍子下到他那里去，从 埃及 人手里夺过枪来，用那枪杀死了他。
1CHR|11|24|这些是 耶何耶大 的儿子 比拿雅 所做的事，就在三个勇士里得了名。
1CHR|11|25|看哪，他比那三十个勇士更有名望，只是不及前三个勇士。 大卫 立他作护卫长。
1CHR|11|26|军中的勇士有 约押 的兄弟 亚撒黑 ， 伯利恒 人 朵多 的儿子 伊勒哈难 ，
1CHR|11|27|哈律 人 沙玛 ， 比伦 人 希利斯 ，
1CHR|11|28|提哥亚 人 益吉 的儿子 以拉 ， 亚拿突 人 亚比以谢 ，
1CHR|11|29|户沙 人 西比该 ， 亚何亚 人 以来 ，
1CHR|11|30|尼陀法 人 玛哈莱 ， 尼陀法 人 巴拿 的儿子 希立 ，
1CHR|11|31|便雅悯 族 基比亚 人 利拜 的儿子 以太 ， 比拉顿 人 比拿雅 ，
1CHR|11|32|迦实溪 人 户莱 ， 亚拉巴 人 亚比 ，
1CHR|11|33|巴路米 人 押斯玛弗 ， 沙本 人 以利雅哈巴 ，
1CHR|11|34|基孙 人 哈深 的众儿子， 哈拉 人 沙基 的儿子 约拿单 ，
1CHR|11|35|哈拉 人 沙甲 的儿子 亚希暗 ， 吾珥 的儿子 以利法勒 ，
1CHR|11|36|米基拉 人 希弗 ， 比伦 人 亚希雅 ，
1CHR|11|37|迦密 人 希斯罗 ， 伊斯拜 的儿子 拿莱 ，
1CHR|11|38|拿单 的兄弟 约珥 ， 哈基利 的儿子 弥伯哈 ，
1CHR|11|39|亚扪 人 洗勒 ， 比录 人 拿哈莱 ，他是给 洗鲁雅 的儿子 约押 拿兵器的，
1CHR|11|40|以帖 人 以拉 ， 以帖 人 迦立 ，
1CHR|11|41|赫 人 乌利亚 ， 亚莱 的儿子 撒拔 ，
1CHR|11|42|吕便 人 示撒 的儿子 亚第拿 ，是 吕便 支派中的一个领袖，率领三十人，
1CHR|11|43|玛迦 的儿子 哈难 ， 弥特尼 人 约沙法 ，
1CHR|11|44|亚施他拉 人 乌西亚 ， 亚罗珥 人 何坦 的儿子 沙玛 和 耶利 ，
1CHR|11|45|提洗 人 申利 的儿子 耶叠 和他的兄弟 约哈 ，
1CHR|11|46|玛哈未 人 以利业 ， 伊利拿安 的儿子 耶利拜 和 约沙未雅 ， 摩押 人 伊特玛 、
1CHR|11|47|以利业 、 俄备得 ，以及 米琐八 人 雅西业 。
1CHR|12|1|以下是 大卫 因 基士 的儿子 扫罗 的缘故被放逐到 洗革拉 的时候，到他那里帮助他打仗的勇士；
1CHR|12|2|他们是弓箭手，能左右甩石，开弓射箭，都是 便雅悯 人 扫罗 同族的弟兄：
1CHR|12|3|为首的是 亚希以谢 ，其次是 约阿施 ，都是 基比亚 人 示玛 的儿子。还有 亚斯玛威 的儿子 耶薛 和 毗力 ， 比拉迦 ， 亚拿突 人 耶户 ，
1CHR|12|4|基遍 人 以实买雅 ，他在三十人中是勇士，管理这三十人，又有 耶利米 ， 雅哈悉 ， 约哈难 ， 基底拉 人 约撒拔 ，
1CHR|12|5|伊利乌赛 ， 耶利末 ， 比亚利雅 ， 示玛利雅 ， 哈律弗 人 示法提雅 ，
1CHR|12|6|可拉 人 以利加拿 、 耶西亚 、 亚萨列 、 约以谢 、 雅朔班 ，
1CHR|12|7|基多 人 耶罗罕 的儿子 犹拉 和 西巴第雅 。
1CHR|12|8|迦得 人中有人到旷野的山寨投奔 大卫 ，都是大能的勇士，能拿盾牌和枪的战士。他们的面貌好像狮子，敏捷如山上的鹿。
1CHR|12|9|第一 以薛 ，第二 俄巴底雅 ，第三 以利押 ，
1CHR|12|10|第四 弥施玛拿 ，第五 耶利米 ，
1CHR|12|11|第六 亚太 ，第七 以利业 ，
1CHR|12|12|第八 约哈难 ，第九 以利萨巴 ，
1CHR|12|13|第十 耶利米 ，第十一 末巴奈 。
1CHR|12|14|这些都是 迦得 人中的军官，小的能抵一百人，大的能抵一千人 。
1CHR|12|15|正月， 约旦河 水涨过两岸的时候，他们过河，使所有住河谷的人东奔西逃。
1CHR|12|16|便雅悯 人和 犹大 人中有人来到山寨 大卫 那里。
1CHR|12|17|大卫 出去迎接他们，回答他们说：“你们若和平地来帮助我，我的心就与你们契合；但你们若把我这双手无辜的人卖给敌人，愿我们列祖的上帝察看责罚。”
1CHR|12|18|那时军官 的领袖 亚玛撒 受灵的感动说： “ 大卫 啊，我们归向你！ 耶西 的儿子啊，我们帮助你！ 愿你平平安安， 愿帮助你的也都平安！ 因为你的上帝帮助你。” 大卫 就收留他们，派他们作军官。
1CHR|12|19|大卫 从前与 非利士 人同去，要与 扫罗 争战，有些 玛拿西 人来投奔 大卫 。其实他们并没有帮助 非利士 人，因为 非利士 人的领袖商议，打发他回去，说：“恐怕 大卫 拿我们的首级去向他的主人 扫罗 投诚。”
1CHR|12|20|大卫 往 洗革拉 去的时候，有 玛拿西 人的千夫长 押拿 、 约撒拔 、 耶叠 、 米迦勒 、 约撒拔 、 以利户 、 洗勒太 都来投奔他。
1CHR|12|21|他们帮助 大卫 攻击敌军；因为他们都是大能的勇士，又作军官。
1CHR|12|22|那时天天有人来帮助 大卫 ，以致成了强大的军队，如上帝的军队一样。
1CHR|12|23|以下是来到 希伯仑 见 大卫 ，要照耶和华的话把 扫罗 的国位归给 大卫 的武装士兵的数目：
1CHR|12|24|犹大 人，拿盾牌和枪的武装战士有六千八百人。
1CHR|12|25|西缅 人中，能上阵的大能勇士有七千一百人。
1CHR|12|26|利未 人中，有四千六百人。
1CHR|12|27|耶何耶大 是 亚伦 家的领袖，跟从他的有三千七百人。
1CHR|12|28|还有大能的青年勇士 撒督 ，同他本族的二十二个军官。
1CHR|12|29|便雅悯 人中， 扫罗 同族的弟兄也有三千人；直到现在他们大部分仍然效忠 扫罗 家。
1CHR|12|30|以法莲 人中，在本族中著名的大能勇士有二万零八百人。
1CHR|12|31|玛拿西 半支派，册上有名来拥立 大卫 作王的，有一万八千人。
1CHR|12|32|以萨迦 人中，通达时务，知道 以色列 所当行，同族弟兄也都听从他们命令的族长有二百人。
1CHR|12|33|西布伦 中，能上阵用各样作战的兵器、不生二心帮助打仗的有五万人。
1CHR|12|34|拿弗他利 中，有一千个军官；跟从他们、拿盾牌和枪的有三万七千人。
1CHR|12|35|但 人中，能摆阵的有二万八千六百人。
1CHR|12|36|亚设 中，能上阵打仗的有四万人。
1CHR|12|37|约旦河 东的 吕便 人、 迦得 人、 玛拿西 半支派，拿各样兵器打仗的有十二万人。
1CHR|12|38|以上都是能列队上阵的战士，他们都全心来到 希伯仑 ，要拥立 大卫 作全 以色列 的王。 以色列 其余的人也都一心要拥立 大卫 作王。
1CHR|12|39|他们在那里三日，与 大卫 一同吃喝，因为他们同族的弟兄已经为他们预备好了。
1CHR|12|40|他们附近的人，以及 以萨迦 、 西布伦 、 拿弗他利 人，都将食物，许多面饼、无花果饼、干葡萄、酒、油，用驴、骆驼、骡子、牛驮来，又带了许多的牛和羊来，因为在 以色列 中充满了欢乐。
1CHR|13|1|大卫 与千夫长、百夫长，以及所有的领袖商议。
1CHR|13|2|大卫 对 以色列 全会众说：“你们若以为好，见这事是出于耶和华－我们的上帝，我们就派人到远近各处去见仍留在 以色列 各地我们的弟兄，以及住在有郊野之城的祭司和 利未 人，使他们都到我们这里来聚集。
1CHR|13|3|我们要把上帝的约柜接到这里来；因为在 扫罗 年间，我们没有去寻求约柜 。”
1CHR|13|4|全会众都说可以这么做，因这事在众百姓眼中都看为好。
1CHR|13|5|于是， 大卫 把 以色列 众人从 埃及 的 西曷河 直到 哈马口 都召集了来，要从 基列．耶琳 将上帝的约柜接来。
1CHR|13|6|大卫 率领 以色列 众人上到 巴拉 ，就是属 犹大 的 基列．耶琳 ，要将耶和华上帝的约柜从那里接上来，他坐在二基路伯之上，这约柜是以他的名来命名的。
1CHR|13|7|他们将上帝的约柜从 亚比拿达 的家里抬出来，放在新车上，由 乌撒 和 亚希约 赶车。
1CHR|13|8|大卫 和 以色列 众人在上帝面前随着诗歌、琴、瑟、鼓、钹、号，极力跳舞。
1CHR|13|9|到了 基顿 的禾场，因为牛失前蹄 ， 乌撒 就伸手扶住约柜。
1CHR|13|10|耶和华的怒气向 乌撒 发作，因他伸手扶住约柜而击杀他，他就死在那里，在上帝面前。
1CHR|13|11|大卫 因耶和华突然冲出撞死 乌撒 就生气，称那地方为 毗列斯．乌撒 ，直到今日。
1CHR|13|12|那日， 大卫 惧怕上帝，说：“我怎能将上帝的约柜接到我这里来呢？”
1CHR|13|13|于是 大卫 不将约柜接进 大卫城 他自己的地方，却转送到 迦特 人 俄别．以东 的家中。
1CHR|13|14|上帝的约柜停在 俄别．以东 家中三个月，耶和华赐福给 俄别．以东 的家和他一切所有的。
1CHR|14|1|推罗 王 希兰 派使者把香柏木运到 大卫 那里，又派石匠和木匠给 大卫 建造宫殿。
1CHR|14|2|大卫 知道耶和华坚立他作 以色列 王，又为自己百姓 以色列 的缘故，使他的国兴盛。
1CHR|14|3|大卫 在 耶路撒冷 又立后妃，又生儿女。
1CHR|14|4|在 耶路撒冷 所生的孩子名字是 沙母亚 、 朔罢 、 拿单 、 所罗门 、
1CHR|14|5|益辖 、 以利书亚 、 以法列 、
1CHR|14|6|挪迦 、 尼斐 、 雅非亚 、
1CHR|14|7|以利沙玛 、 比利雅大 、 以利法列 。
1CHR|14|8|非利士 人听见 大卫 受膏作全 以色列 的王， 非利士 众人就上来寻索 大卫 。 大卫 听见了，就出去迎敌。
1CHR|14|9|非利士 人来了，侵犯 利乏音谷 。
1CHR|14|10|大卫 求问上帝说：“我可以上去攻打 非利士 人吗？你将他们交在我手里吗？”耶和华对他说：“你可以上去，我必将他们交在你手里。”
1CHR|14|11|非利士 人上到 巴力．毗拉心 ， 大卫 在那里击败他们。 大卫 说：“上帝藉我的手冲破敌人，如水冲破一样。”因此那地方称为 巴力．毗拉心 。
1CHR|14|12|非利士 人把神像抛弃在那里， 大卫 吩咐人用火焚烧了。
1CHR|14|13|非利士 人又侵犯 利乏音谷 。
1CHR|14|14|大卫 再求问上帝。上帝对他说：“不要从他们后头追上去，要绕道离开他们，从桑树林对面攻打他们。
1CHR|14|15|你听见桑树梢上有脚步的声音，那时你就要出战，因为上帝已经出去，在你前头攻打 非利士 人的军队了。”
1CHR|14|16|大卫 就遵照上帝所吩咐的去做，攻打 非利士 人的军队，从 基遍 直到 基色 。
1CHR|14|17|于是 大卫 的名传扬到万邦，耶和华使万国都惧怕他。
1CHR|15|1|大卫 在 大卫城 为自己建造宫殿，又为上帝的约柜预备地方，支搭帐幕。
1CHR|15|2|那时 大卫 说：“除了 利未 人之外，无人可抬上帝的约柜，因为耶和华拣选他们抬上帝的约柜，永远事奉他。”
1CHR|15|3|大卫 召集 以色列 众人到 耶路撒冷 ，要将耶和华的约柜接到他所预备的地方。
1CHR|15|4|大卫 又召集 亚伦 的子孙和 利未 人：
1CHR|15|5|哥辖 子孙中有领袖 乌列 和他的弟兄一百二十人，
1CHR|15|6|米拉利 子孙中有领袖 亚帅雅 和他的弟兄二百二十人，
1CHR|15|7|革顺 子孙中有领袖 约珥 和他的弟兄一百三十人，
1CHR|15|8|以利撒反 子孙中有领袖 示玛雅 和他的弟兄二百人，
1CHR|15|9|希伯伦 子孙中有领袖 以利业 和他的弟兄八十人，
1CHR|15|10|乌薛 子孙中有领袖 亚米拿达 和他的弟兄一百一十二人。
1CHR|15|11|大卫 召来 撒督 和 亚比亚他 二位祭司，以及 利未 人 乌列 、 亚帅雅 、 约珥 、 示玛雅 、 以利业 、 亚米拿达 ，
1CHR|15|12|对他们说：“你们是 利未 人的族长，你们和你们的弟兄应当使自己分别为圣，好将耶和华－ 以色列 上帝的约柜接到我所预备的地方。
1CHR|15|13|因为你们上一次没有抬这约柜，并且我们没有按规矩求问耶和华－我们的上帝，所以他冲出来攻击我们。”
1CHR|15|14|于是祭司和 利未 人使自己分别为圣，将耶和华－ 以色列 上帝的约柜接上来。
1CHR|15|15|利未 子孙用杠，把上帝的约柜抬在肩上，正如 摩西 按照耶和华的话所吩咐的。
1CHR|15|16|大卫 吩咐 利未 人的领袖派他们歌唱的弟兄用琴瑟和钹的乐器奏乐，欢欢喜喜地大声歌颂。
1CHR|15|17|于是 利未 人派 约珥 的儿子 希幔 和他弟兄中 比利家 的儿子 亚萨 ，以及他们同族弟兄 米拉利 子孙里 古沙雅 的儿子 以探 。
1CHR|15|18|其次还有跟随他们的弟兄 撒迦利雅 、 便．雅薛 、 示米拉末 、 耶歇 、 乌尼 、 以利押 、 比拿雅 、 玛西雅 、 玛他提雅 、 以利斐利户 、 弥克尼雅 ，以及门口的守卫 俄别．以东 和 耶利 。
1CHR|15|19|歌唱的 希幔 、 亚萨 和 以探 ，敲铜钹，声音响亮；
1CHR|15|20|撒迦利雅 、 雅薛 、 示米拉末 、 耶歇 、 乌尼 、 以利押 、 玛西雅 、 比拿雅 鼓瑟，调用女音；
1CHR|15|21|玛他提雅 、 以利斐利户 、 弥克尼雅 、 俄别．以东 、 耶利 、 亚撒西雅 用琴指挥，调用第八。
1CHR|15|22|基拿尼雅 是 利未 人圣咏团的领袖，又教导人唱歌，因为他精通此事。
1CHR|15|23|比利家 和 以利加拿 是约柜的守卫。
1CHR|15|24|示巴尼 、 约沙法 、 拿坦业 、 亚玛赛 、 撒迦利雅 、 比拿亚 、 以利以谢 众祭司在上帝的约柜前吹号。 俄别．以东 和 耶希亚 也是约柜的守卫。
1CHR|15|25|于是， 大卫 和 以色列 的长老，以及千夫长都去，欢欢喜喜地将耶和华的约柜从 俄别．以东 家中接上来。
1CHR|15|26|上帝赐恩给抬耶和华约柜的 利未 人，他们就献上七头公牛，七只公羊。
1CHR|15|27|大卫 和所有抬约柜的 利未 人，以及圣咏团的领袖 基拿尼雅 和歌唱的人，都穿着细麻布外袍； 大卫 另外穿着细麻布以弗得。
1CHR|15|28|这样， 以色列 众人欢呼、吹角、吹号、敲钹、鼓瑟、弹琴，声音响亮，将耶和华的约柜接上来。
1CHR|15|29|耶和华的约柜进 大卫城 的时候， 扫罗 的女儿 米甲 从窗户里往外观看，见 大卫 王踊跃跳舞，心里就轻视他。
1CHR|16|1|众人将上帝的约柜请进去，安放在 大卫 为它搭的帐幕中，就在上帝面前献燔祭和平安祭。
1CHR|16|2|大卫 献完了燔祭和平安祭，就奉耶和华的名祝福百姓，
1CHR|16|3|并且分给每一个 以色列 人，无论男女，每人一个饼，一个枣子饼 ，一个葡萄饼。
1CHR|16|4|大卫 派几个 利未 人在耶和华的约柜前事奉，颂扬，称谢，赞美耶和华－ 以色列 的上帝：
1CHR|16|5|为首的是 亚萨 ，其次是 撒迦利雅 、 耶利 、 示米拉末 、 耶歇 、 玛他提雅 、 以利押 、 比拿雅 、 俄别．以东 、 耶利 ；他们鼓瑟弹琴， 亚萨 敲钹，声音响亮；
1CHR|16|6|比拿雅 和 雅哈悉 二位祭司常在上帝的约柜前吹号。
1CHR|16|7|那日， 大卫 初次指派 亚萨 和他的弟兄称谢耶和华。
1CHR|16|8|你们要称谢耶和华，求告他的名， 在万民中传扬他的作为！
1CHR|16|9|要向他唱诗，向他歌颂， 述说他一切奇妙的作为！
1CHR|16|10|要夸耀他的圣名！ 愿寻求耶和华的人心中欢喜！
1CHR|16|11|要寻求耶和华与他的能力， 时常寻求他的面。
1CHR|16|12|他仆人 以色列 的后裔， 他所拣选 雅各 的子孙哪， 要记念他奇妙的作为和他的奇事， 并他口中的判语。
1CHR|16|13|
1CHR|16|14|他是耶和华－我们的上帝， 全地都有他的判断。
1CHR|16|15|要记念他的约，直到永远； 记念他吩咐的话，直到千代，
1CHR|16|16|就是他与 亚伯拉罕 所立的约， 向 以撒 所起的誓。
1CHR|16|17|他将这约向 雅各 定为律例， 向 以色列 定为永远的约，
1CHR|16|18|说：“我必将 迦南 地赐给你， 作你们应得的产业。”
1CHR|16|19|当时，你们人丁有限， 数目稀少，在那地寄居。
1CHR|16|20|他们从这邦游到那邦， 从这国去到另一民族。
1CHR|16|21|他不容人欺负他们， 为他们的缘故责备君王：
1CHR|16|22|“不可伤害我的受膏者， 也不可恶待我的先知。”
1CHR|16|23|全地都要向耶和华歌唱！ 天天传扬他的救恩！
1CHR|16|24|在列国中述说他的荣耀！ 在万民中述说他的奇事！
1CHR|16|25|因耶和华本为大，当受极大的赞美； 他在万神之上，当受敬畏。
1CHR|16|26|因万民的神明都属虚无； 惟独耶和华创造诸天。
1CHR|16|27|有尊荣和威严在他面前， 有能力和喜乐在他自己的地方。
1CHR|16|28|民中的万族啊，要将荣耀、能力归给耶和华， 都归给耶和华！
1CHR|16|29|要将耶和华的名所当得的荣耀归给他， 拿供物来献在他面前； 当敬拜神圣荣耀的耶和华 。
1CHR|16|30|全地都要在他面前战抖！ 世界坚定，不得动摇。
1CHR|16|31|愿天欢喜，愿地快乐！ 愿人在列国中说： “耶和华作王了！”
1CHR|16|32|愿海和其中所充满的澎湃！ 愿田和其中所有的都欢乐！
1CHR|16|33|那时，林中的树木都要在耶和华面前欢呼， 因为他来要审判全地。
1CHR|16|34|你们要称谢耶和华，因他本为善， 他的慈爱永远长存！
1CHR|16|35|你们要说： “拯救我们的上帝啊，求你拯救我们， 聚集我们，救我们脱离列国， 我们好颂扬你的圣名， 以赞美你为夸胜。
1CHR|16|36|耶和华－ 以色列 的上帝是应当称颂的， 从亘古直到永远。” 全体百姓都说：“阿们！”并且赞美耶和华。
1CHR|16|37|大卫 把 亚萨 和他的弟兄留在耶和华的约柜那里，经常在约柜前事奉，天天尽本分供职，
1CHR|16|38|又有 俄别．以东 和他的弟兄六十八人； 耶杜顿 的儿子 俄别．以东 ，以及 何萨 作门口的守卫。
1CHR|16|39|还有 撒督 祭司和他弟兄众祭司在 基遍 的丘坛、耶和华的帐幕前，
1CHR|16|40|在燔祭坛上，每日早晚，照着写在耶和华律法书上所吩咐 以色列 的，经常献燔祭给耶和华。
1CHR|16|41|与他们一同的还有 希幔 、 耶杜顿 ，和其余被选、名字录在册上的，为要称谢耶和华，因他的慈爱永远长存。
1CHR|16|42|希幔 、 耶杜顿 同他们吹号、敲钹，声音响亮，并用其他乐器配合，歌颂上帝。 耶杜顿 的子孙作门口的守卫。
1CHR|16|43|于是众百姓各自回家， 大卫 也回去为家人祝福。
1CHR|17|1|大卫 住在自己宫中，对 拿单 先知说：“看哪，我住在香柏木的宫中，耶和华的约柜却在幔子里。”
1CHR|17|2|拿单 对 大卫 说：“你可以完全照你的心意去做，因为上帝与你同在。”
1CHR|17|3|当夜上帝的话临到 拿单 ，说：
1CHR|17|4|“你去对我仆人 大卫 说：‘耶和华如此说：你不可建造殿宇给我居住。
1CHR|17|5|自从我领 以色列 人上来，直到今日，我未曾住过殿宇；我从这会幕到那会幕，从这帐幕到那帐幕 。
1CHR|17|6|凡我同 以色列 人所走的地方，我何曾向 以色列 的一个士师，就是我吩咐牧养我百姓的，说过这话：你们为何不给我建造香柏木的殿宇呢？’
1CHR|17|7|现在，你要对我仆人 大卫 这样说：‘万军之耶和华如此说：我从羊圈中将你召来，叫你不再牧放羊群，立你作我百姓 以色列 的君王。
1CHR|17|8|你无论往哪里去，我都与你同在，剪除你所有的仇敌。我必使你得大名，好像世上伟人的名一样。
1CHR|17|9|我必为我百姓 以色列 选定一个地方，栽植他们，使他们住自己的地方，不再受搅扰；凶恶之子也不再像从前那样扰乱他们，
1CHR|17|10|并不像我命令士师治理我百姓 以色列 的日子。我必制伏你所有的仇敌，并且我应许你 ，耶和华必为你建立家室。
1CHR|17|11|当你寿数满足归你祖先的时候，我必使你的后裔，你自己的儿子接续你；我也必坚定他的国。
1CHR|17|12|他必为我建造殿宇，我必坚定他的王位，直到永远。
1CHR|17|13|我要作他的父，他要作我的子；我必不使我的慈爱离开他，像离开在你以前的那位一样。
1CHR|17|14|我要永远坚立他在我的家和我的国里；他的王位也必坚定，直到永远。’”
1CHR|17|15|拿单 就按这一切话，照这一切异象告诉 大卫 。
1CHR|17|16|于是 大卫 王进去，坐在耶和华面前，说：“耶和华上帝啊，我是谁，我的家算什么，你竟带领我到这地步呢？
1CHR|17|17|上帝啊，这在你眼中还看为小，你又说到你仆人的家将来的情况。耶和华上帝啊，你看顾我好像看顾尊贵的人。
1CHR|17|18|你加于仆人的尊荣， 大卫 还有什么可以对你说呢？你是知道你仆人的。
1CHR|17|19|耶和华啊，因你仆人的缘故，也照着你的心意，你行这一切大事，为了显明这一切伟大的事。
1CHR|17|20|耶和华啊，照我们耳中一切所听见的，没有可比你的，除你以外再没有上帝。
1CHR|17|21|世上有何国能比你的百姓 以色列 呢？上帝亲自去救赎世上的一国 ，作自己的子民，又行大而可畏的事，显出你的大名，在你从 埃及 赎出来的子民面前驱逐了列国。
1CHR|17|22|你使你的百姓 以色列 作你的子民，直到永远；你－耶和华也作他们的上帝。
1CHR|17|23|现在，耶和华啊，你所应许仆人和仆人家的话，求你坚定，直到永远；求你照你所说的而行。
1CHR|17|24|愿你的名永远坚立，被尊为大，人要说：‘万军之耶和华－ 以色列 的上帝，是 以色列 的上帝。’这样，你仆人 大卫 的家必在你面前坚立。
1CHR|17|25|我的上帝啊，因你启示你的仆人，要为他建立家室，所以仆人大胆在你面前祈祷。
1CHR|17|26|现在，耶和华啊，惟有你是上帝！你应许将这福气赐给仆人。
1CHR|17|27|现在，你喜悦赐福给仆人的家，可以永存在你面前。耶和华啊，因你已经赐福，还要赐福到永远。”
1CHR|18|1|此后， 大卫 攻打 非利士 人，制伏了他们，从 非利士 人手中夺取了 迦特 和所属的乡镇。
1CHR|18|2|他又攻打 摩押 ， 摩押 人就臣服 大卫 ，向他进贡。
1CHR|18|3|琐巴 王 哈大底谢 往 幼发拉底河 去，要巩固自己的国权。 大卫 攻打他，直到 哈马 ，
1CHR|18|4|夺了他的战车一千，俘掳了骑兵七千人，步兵二万人。 大卫 把所有战马的蹄筋砍断，只留下一百辆战车。
1CHR|18|5|大马士革 的 亚兰 人来帮助 琐巴 王 哈大底谢 ， 大卫 杀了 亚兰 人二万二千。
1CHR|18|6|于是 大卫 在 大马士革 的 亚兰 地设立军营 ， 亚兰 人就臣服 大卫 ，向他进贡。 大卫 无论往哪里去，耶和华都使他得胜。
1CHR|18|7|大卫 夺了 哈大底谢 臣仆拥有的金盾牌，带到 耶路撒冷 。
1CHR|18|8|大卫 又从 哈大底谢 的 提巴 和 均 二城夺取了许多的铜；后来 所罗门 用这些铜制造铜海、铜柱和铜器。
1CHR|18|9|哈马 王 陀乌 听见 大卫 击败 琐巴 王 哈大底谢 的全军，
1CHR|18|10|就派他儿子 哈多兰 到 大卫 王那里，向他请安，为他祝福，因他与 哈大底谢 争战，并且击败了他；原来 哈大底谢 与 陀乌 常常争战。 哈多兰 带了金银铜的各样器皿来。
1CHR|18|11|大卫 王把这些器皿，以及从各国夺来的金银，就是从 以东 、 摩押 、 亚扪 人、 非利士 人、 亚玛力 所夺来的，都分别为圣献给耶和华。
1CHR|18|12|洗鲁雅 的儿子 亚比筛 在 盐谷 击杀了一万八千 以东 人。
1CHR|18|13|大卫 在 以东 设立军营， 以东 人就都臣服他。 大卫 无论往哪里去，耶和华都使他得胜。
1CHR|18|14|大卫 作全 以色列 的王，又向众百姓秉公行义。
1CHR|18|15|洗鲁雅 的儿子 约押 作元帅； 亚希律 的儿子 约沙法 作史官；
1CHR|18|16|亚希突 的儿子 撒督 和 亚比亚他 的儿子 亚希米勒 作祭司； 沙威沙 作书记；
1CHR|18|17|耶何耶大 的儿子 比拿雅 管辖 基利提 人和 比利提 人。 大卫 的众儿子都在王的左右作领袖。
1CHR|19|1|此后， 亚扪 人的王 拿辖 死了，他儿子接续他作王。
1CHR|19|2|大卫 说：“ 哈嫩 的父亲 拿辖 怎样向我施恩，我也要怎样向 哈嫩 施恩。”于是 大卫 派使者为他的父亲安慰他。 大卫 的臣仆到了 亚扪 人的境内来见 哈嫩 ，要安慰他。
1CHR|19|3|但 亚扪 人的领袖对 哈嫩 说：“ 大卫 派人来安慰你，你看他是要尊敬你父亲吗？他的臣仆来见你，不是为了要窥探侦察，而倾覆这地吗？”
1CHR|19|4|哈嫩 就抓住 大卫 的臣仆，剃去他们的胡须，又割断他们下半截的衣服，露出臀部，然后放了他们。
1CHR|19|5|他们走了，有人把臣仆所遭遇的事告诉 大卫 ，他就派人去迎接他们，因为这些人觉得很羞耻。王说：“可以住在 耶利哥 ，等到胡须长出来再回来。”
1CHR|19|6|亚扪 人看到 大卫 憎恶他们， 哈嫩 和 亚扪 人就派人拿一千他连得银子，从 美索不达米亚 、 亚兰．玛迦 、 琐巴 雇用战车和骑兵。
1CHR|19|7|他们雇了三万二千辆战车，以及 玛迦 王和他的军兵；这些部队来安营在 米底巴 前。 亚扪 人也从他们的城里出来，聚集预备作战。
1CHR|19|8|大卫 听见了，就派 约押 和所有勇猛的军队出去。
1CHR|19|9|亚扪 人出来，在城门前摆阵，前来的诸王另在郊野摆阵。
1CHR|19|10|约押 看见战阵对着他前后摆列，就把从 以色列 所有精兵中挑选出来的，摆阵迎战 亚兰 人。
1CHR|19|11|他把其余的兵交在他兄弟 亚比筛 手里，他们就摆阵迎战 亚扪 人。
1CHR|19|12|约押 说：“ 亚兰 人若强过我，你就来帮助我； 亚扪 人若强过你，我就去帮助你。
1CHR|19|13|你要刚强，我们要为自己的百姓，为我们上帝的城镇奋勇。愿耶和华照他所看为好的去做！”
1CHR|19|14|于是， 约押 和跟随他的士兵前进攻打 亚兰 人； 亚兰 人在他面前逃跑。
1CHR|19|15|亚扪 人见 亚兰 人逃跑，他们也在 约押 的兄弟 亚比筛 面前逃跑进城。 约押 就回 耶路撒冷 去了。
1CHR|19|16|亚兰 人见自己被 以色列 打败，就派使者把 大河 那边的 亚兰 人调来，由 哈大底谢 的将军 朔法 在他们前面率领。
1CHR|19|17|有人告诉 大卫 ，他就聚集 以色列 众人过 约旦河 ，来到 亚兰 人那里，迎着他们摆阵。 大卫 摆阵攻击 亚兰 人， 亚兰 人就与他打仗。
1CHR|19|18|亚兰 人在 以色列 人面前逃跑。 大卫 杀了 亚兰 七千辆战车的士兵，四万步兵，又杀死 亚兰 的将军 朔法 。
1CHR|19|19|哈大底谢 的臣仆见自己被 以色列 打败，就与 大卫 讲和，臣服他。于是 亚兰 人不愿再帮助 亚扪 人了。
1CHR|20|1|到了年初，诸王出征的时候， 约押 率领军兵蹂躏 亚扪 人的地，前来围攻 拉巴 ； 大卫 仍住在 耶路撒冷 。 约押 攻打 拉巴 ，把它毁坏。
1CHR|20|2|大卫 夺了 米勒公 所戴的冠冕，其上的金子重一他连得，又嵌着宝石。这冠冕就戴在 大卫 头上。 大卫 又从城里夺了许多财物，
1CHR|20|3|把城里的百姓拉出来，放在锯下，或铁耙下，或斧 的下面； 大卫 待 亚扪 各城的居民都是如此。于是， 大卫 和全军都回 耶路撒冷 去了。
1CHR|20|4|后来， 以色列 人在 基色 与 非利士 人打仗。 户沙 人 西比该 杀了巨人族的后裔 细派 ， 非利士 人就被制伏了。
1CHR|20|5|他们又与 非利士 人打仗。 睚珥 的儿子 伊勒哈难 杀了 迦特 人 歌利亚 的兄弟 拉哈米 ；这人的枪杆粗如织布机的轴。
1CHR|20|6|又有一次，他们在 迦特 打仗。那里有一个身材高大的人，手指脚趾都是六根，共有二十四根；他也是巨人族的后裔。
1CHR|20|7|他向 以色列 骂阵， 大卫 的哥哥 示米亚 的儿子 约拿单 就杀了他。
1CHR|20|8|这些人是 迦特 巨人族的后裔，都仆倒在 大卫 和他仆人的手下。
1CHR|21|1|撒但起来攻击 以色列 ，激起 大卫 数点以色列人。
1CHR|21|2|大卫 对 约押 和百姓的领袖说：“去，数点 以色列 人，从 别是巴 直到 但 ，回来告诉我，我好知道他们的数目。”
1CHR|21|3|约押 说：“愿耶和华使他的百姓比现在加增百倍。我主我王啊，他们不都是我主的仆人吗？我主为何吩咐行这事，为何使 以色列 陷入罪里呢？”
1CHR|21|4|但王坚持他对 约押 的命令。 约押 就出去，来回走遍 以色列 ，然后回到 耶路撒冷 。
1CHR|21|5|约押 向 大卫 报告百姓的总数：全 以色列 拿刀的有一百一十万人； 犹大 拿刀的有四十七万人。
1CHR|21|6|惟有 利未 人和 便雅悯 人没有算在其中，因为 约押 厌恶王的这命令。
1CHR|21|7|这件事在上帝眼中看为恶，上帝就降灾给 以色列 。
1CHR|21|8|大卫 对上帝说：“我做这事大大有罪了。现在求你除掉仆人的罪孽，因为我所做的非常愚昧。”
1CHR|21|9|耶和华吩咐 迦得 ， 大卫 的先见，说：
1CHR|21|10|“你去告诉 大卫 说：‘耶和华如此说：我列出三样灾祸给你，随你选择一样，我好降与你。’”
1CHR|21|11|于是， 迦得 来到 大卫 那里，对他说：“耶和华如此说：‘你可以随意选择：
1CHR|21|12|三年的饥荒，或败在敌人面前，被敌人的刀追杀三个月，或在国中三日有耶和华的刀，就是瘟疫，让耶和华的使者在 以色列 全境施行毁灭呢？’现在你要想一想，我怎样去回覆那差我来的。”
1CHR|21|13|大卫 对 迦得 说：“我很为难。我宁愿落在耶和华的手里，因为他有丰盛的怜悯；我不愿落在人的手里。”
1CHR|21|14|于是，耶和华降瘟疫给 以色列 ， 以色列 中死了七万人。
1CHR|21|15|上帝派遣使者去毁灭 耶路撒冷 ，刚要毁灭的时候，耶和华看见就改变心意，不降这灾了。他吩咐那灭城的天使说：“够了，住手吧！”耶和华的使者正站在 耶布斯 人 阿珥楠 的禾场那里。
1CHR|21|16|大卫 举目，看见耶和华的使者站在天和地之间，手里有拔出来的刀，伸在 耶路撒冷 以上。 大卫 和长老都披上麻布，脸伏于地。
1CHR|21|17|大卫 向上帝说：“吩咐数点百姓的不是我吗？是我犯了罪，行了大恶，但这群羊做了什么呢？耶和华－我的上帝啊，愿你的手攻击我和我的父家，不要降瘟疫给你的百姓。”
1CHR|21|18|耶和华的使者吩咐 迦得 去告诉 大卫 ，叫他上去，在 耶布斯 人 阿珥楠 的禾场上为耶和华立一座坛。
1CHR|21|19|大卫 就照着 迦得 奉耶和华名所说的话上去。
1CHR|21|20|阿珥楠 回头看见天使，跟他在一起的四个儿子都藏起来了， 阿珥楠 继续打麦子。
1CHR|21|21|大卫 到了 阿珥楠 那里， 阿珥楠 观看，看见 大卫 ，就从禾场上出去，脸伏于地，向他下拜。
1CHR|21|22|大卫 对 阿珥楠 说：“你把这禾场的地方给我，照着十足的价钱卖给我，我好在其上为耶和华筑一座坛，使瘟疫在百姓中停止。”
1CHR|21|23|阿珥楠 对 大卫 说：“请用这禾场吧，愿我主我王照你眼中看为好的去做。看，我提供牛作燔祭，打粮的器具作柴，麦子作素祭，这一切我全都提供。”
1CHR|21|24|大卫 王对 阿珥楠 说：“不，我一定要按十足的价钱买；因我不能用你的东西献给耶和华，也不能用白得之物献为燔祭。”
1CHR|21|25|于是 大卫 为那个地方付了六百舍客勒重的金子给 阿珥楠 。
1CHR|21|26|大卫 在那里为耶和华筑了一座坛，献燔祭和平安祭，求告耶和华。耶和华就应允他，使火从天降在燔祭坛上。
1CHR|21|27|耶和华吩咐使者，他就收刀入鞘。
1CHR|21|28|那时， 大卫 见耶和华在 耶布斯 人 阿珥楠 的禾场上应允了他，就在那里献祭。
1CHR|21|29|摩西 在旷野所造之耶和华的帐幕和燔祭坛，当时都在 基遍 的丘坛，
1CHR|21|30|只是 大卫 不能前去求问上帝，因为他惧怕耶和华使者的刀。
1CHR|22|1|大卫 说：“这是耶和华上帝的殿，这是 以色列 献燔祭的坛。”
1CHR|22|2|大卫 吩咐人召集住 以色列 地的寄居者，又派石匠凿石头，要建造上帝的殿。
1CHR|22|3|大卫 预备许多铁，要做门上的钉子和钩子，又预备许多铜，多得无法可秤；
1CHR|22|4|还有无数的香柏木，因为 西顿 人和 推罗 人给 大卫 运了许多香柏木来。
1CHR|22|5|大卫 说：“我儿子 所罗门 还年幼脆弱，要为耶和华建造的殿宇必须高大辉煌，使名声荣耀传遍万国，所以我要为殿预备。”于是， 大卫 在未死之前预备了许多材料。
1CHR|22|6|大卫 召了他儿子 所罗门 来，吩咐他为耶和华－ 以色列 的上帝建造殿宇。
1CHR|22|7|大卫 对 所罗门 说：“我儿啊，我心里本想为耶和华－我上帝的名建造殿宇，
1CHR|22|8|可是耶和华的话临到我说：‘你流了许多的血，打了多次大仗；你不可为我的名建造殿宇，因为你在我面前使许多血流在地上。
1CHR|22|9|看哪，你要生一个儿子，他必成为安宁的人；我必使他得享安宁，不被四围仇敌扰乱。他的名字要叫 所罗门 ，在他的日子，我必使 以色列 平安康泰。
1CHR|22|10|他必为我的名建造殿宇。他要作我的子，我要作他的父。我必坚定他国度的王位，使他治理 以色列 ，直到永远。’
1CHR|22|11|我儿啊，现今愿耶和华与你同在，使你亨通，建造耶和华－你上帝的殿，正如他指着你所说的。
1CHR|22|12|但愿耶和华赐你聪明智慧，好按着他吩咐你的去治理 以色列 ，遵行耶和华－你上帝的律法。
1CHR|22|13|那时候，你若谨守遵行耶和华藉 摩西 吩咐 以色列 的律例典章，就得亨通。你当刚强壮胆，不要惧怕，也不要惊惶。
1CHR|22|14|看哪，我辛苦地为耶和华的殿预备了十万他连得金子，一百万他连得银子，铜和铁多得无法可秤；我也预备了木头、石头，你还可以增添。
1CHR|22|15|你有许多工匠，就是石匠、木匠，和一切能做各样工的巧匠，
1CHR|22|16|以及无数的金银铜铁。你当起来做工，愿耶和华与你同在。”
1CHR|22|17|大卫 又吩咐 以色列 的众官长帮助他儿子 所罗门 ：
1CHR|22|18|“耶和华－你们的上帝不是与你们同在吗？他不是使你们四围都平安吗？因他已将这地的居民交在我手中，这地已在耶和华与他百姓面前制伏了。
1CHR|22|19|现在你们应当立定心意，寻求耶和华－你们的上帝。你们当起来建造耶和华上帝的圣所，好将耶和华的约柜和上帝神圣的器皿都搬进为耶和华的名建造的殿里。”
1CHR|23|1|大卫 年纪老迈，日子满足，就立他儿子 所罗门 作 以色列 的王。
1CHR|23|2|大卫 召集 以色列 的众领袖、祭司和 利未 人。
1CHR|23|3|利未 人三十岁以上的都被数点，他们男丁的数目共有三万八千；
1CHR|23|4|其中有二万四千人管理耶和华殿的事务，有六千人作官长和审判官，
1CHR|23|5|有四千人作门口的守卫，又有四千人颂赞耶和华，用 大卫 造的乐器来颂赞。
1CHR|23|6|大卫 把 利未 人 革顺 、 哥辖 、 米拉利 的子孙分了班次。
1CHR|23|7|属 革顺 的有 拉但 和 示每 。
1CHR|23|8|拉但 的长子是 耶歇 ，还有 西坦 和 约珥 ，共三人。
1CHR|23|9|示每 的儿子是 示罗密 、 哈薛 、 哈兰 三人。这是 拉但 族的族长。
1CHR|23|10|示每 的儿子是 雅哈 、 细拿 、 耶乌施 、 比利亚 ，这四人是 示每 的儿子。
1CHR|23|11|雅哈 是长子， 细撒 是次子。但 耶乌施 和 比利亚 的子孙不多，所以算为一族。
1CHR|23|12|哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 、 乌薛 ，共四人。
1CHR|23|13|暗兰 的儿子是 亚伦 和 摩西 。 亚伦 被分别出来，把至圣之物分别为圣，使他和他的子孙在耶和华面前烧香、事奉他，奉他的名祝福，直到永远。
1CHR|23|14|至于神人 摩西 ，他的子孙记名在 利未 支派下。
1CHR|23|15|摩西 的儿子是 革舜 和 以利以谢 。
1CHR|23|16|革舜 的儿子，长子是 细布业 ；
1CHR|23|17|以利以谢 的儿子，长子是 利哈比雅 。 以利以谢 没有别的儿子，但 利哈比雅 的子孙很多。
1CHR|23|18|以斯哈 的儿子，长子是 示罗密 。
1CHR|23|19|希伯伦 的儿子，长子是 耶利雅 ，次子是 亚玛利亚 ，三子是 雅哈悉 ，四子是 耶加面 。
1CHR|23|20|乌薛 的儿子，长子是 米迦 ，次子是 耶西雅 。
1CHR|23|21|米拉利 的儿子是 抹利 和 母示 。 抹利 的儿子是 以利亚撒 和 基士 。
1CHR|23|22|以利亚撒 死了，没有儿子，只有女儿，他们本族 基士 的几个儿子娶了她们为妻。
1CHR|23|23|母示 的儿子是 末力 、 以得 、 耶列末 ，共三人。
1CHR|23|24|以上是 利未 子孙作族长的，按着父系、照着男丁的数目，二十岁以上登记的，都办理耶和华殿的事务。
1CHR|23|25|大卫 说：“耶和华－ 以色列 的上帝已经使他的百姓得享安宁，他永远住在 耶路撒冷 。
1CHR|23|26|因此， 利未 人不必再抬帐幕和其中所使用的一切器皿了。”
1CHR|23|27|照着 大卫 临终的话， 利未 人二十岁以上的都被数点。
1CHR|23|28|他们的职务是作 亚伦 子孙的帮手，在耶和华的殿事奉，照管院子和屋子，洁净一切圣物，办理上帝殿的事务。
1CHR|23|29|他们负责预备供饼、素祭的细面和无酵薄饼，或用盘烤，或用油调和的祭物，确认其数量和大小。
1CHR|23|30|每日早晚、安息日、初一，以及节期，按数照例，经常献燔祭给耶和华的时候，他们站立称谢赞美耶和华。
1CHR|23|31|
1CHR|23|32|他们照管会幕和圣所，服事他们的弟兄 亚伦 的子孙，办理耶和华殿的事务。
1CHR|24|1|亚伦 子孙的班次如下： 亚伦 的儿子是 拿答 、 亚比户 、 以利亚撒 、 以他玛 。
1CHR|24|2|拿答 和 亚比户 死在他们父亲之先，没有留下儿子；因此， 以利亚撒 和 以他玛 担任祭司的职分。
1CHR|24|3|大卫 和 以利亚撒 的子孙 撒督 ，以及 以他玛 的子孙 亚希米勒 ，把他们按照任务分成班次，
1CHR|24|4|发现 以利亚撒 子孙中作领袖的，比 以他玛 子孙中作领袖的更多，就分班如下： 以利亚撒 的子孙中有十六个族长， 以他玛 的子孙中有八个族长。
1CHR|24|5|他们抽签分配，彼此一样。在圣所和上帝面前作领袖的有 以利亚撒 的子孙，也有 以他玛 的子孙。
1CHR|24|6|作书记的 利未 人 拿坦业 的儿子 示玛雅 在王和领袖，与 撒督 祭司、 亚比亚他 的儿子 亚希米勒 ，以及祭司和 利未 人的族长面前记录他们的名字；在 以利亚撒 的子孙中取一族，在 以他玛 的子孙中也取一族。
1CHR|24|7|抽签的时候，第一签抽到的是 耶何雅立 ，第二是 耶大雅 ，
1CHR|24|8|第三是 哈琳 ，第四是 梭琳 ，
1CHR|24|9|第五是 玛基雅 ，第六是 米雅民 ，
1CHR|24|10|第七是 哈歌斯 ，第八是 亚比雅 ，
1CHR|24|11|第九是 耶书亚 ，第十是 示迦尼 ，
1CHR|24|12|第十一是 以利亚实 ，第十二是 雅金 ，
1CHR|24|13|第十三是 胡巴 ，第十四是 耶是比押 ，
1CHR|24|14|第十五是 璧迦 ，第十六是 音麦 ，
1CHR|24|15|第十七是 希悉 ，第十八是 哈辟悉 ，
1CHR|24|16|第十九是 毗他希雅 ，第二十是 以西结 ，
1CHR|24|17|第二十一是 雅斤 ，第二十二是 迦末 ，
1CHR|24|18|第二十三是 第来雅 ，第二十四是 玛西亚 。
1CHR|24|19|这就是他们事奉的班次，要照耶和华－ 以色列 的上帝藉他们祖宗 亚伦 所吩咐的条例，进入耶和华的殿办理事务。
1CHR|24|20|利未 其余的子孙如下： 暗兰 的子孙中有 书巴业 ； 书巴业 的子孙中有 耶希底亚 。
1CHR|24|21|属 利哈比雅 ， 利哈比雅 的儿子中有长子 伊示雅 。
1CHR|24|22|属 以斯哈 人的有 示罗摩 ； 示罗摩 的子孙中有 雅哈 。
1CHR|24|23|希伯伦 的儿子中有长子 耶利雅 ，次子 亚玛利亚 ，三子 雅哈悉 ，四子 耶加面 。
1CHR|24|24|乌薛 的子孙中有 米迦 ； 米迦 的子孙中有 沙密 。
1CHR|24|25|米迦 的兄弟是 伊示雅 ； 伊示雅 的子孙中有 撒迦利雅 。
1CHR|24|26|米拉利 的儿子是 抹利 和 母示 ； 雅西雅 的子孙中有 比挪 ；
1CHR|24|27|米拉利 的子孙中有属 雅西雅 的 比挪 、 朔含 、 撒刻 、 伊比利 。
1CHR|24|28|属 抹利 的有 以利亚撒 ； 以利亚撒 没有儿子。
1CHR|24|29|属 基士 ， 基士 的子孙中有 耶拉篾 。
1CHR|24|30|母示 的儿子是 末力 、 以得 、 耶利末 。按着宗族，这些都是 利未 的子孙。
1CHR|24|31|他们在 大卫 王和 撒督 ，以及 亚希米勒 与祭司和 利未 人的族长面前也抽签，正如他们弟兄 亚伦 的子孙一样。各族的族长与最年轻的兄弟都一样。
1CHR|25|1|大卫 和事奉团队的众领袖分派 亚萨 、 希幔 ，以及 耶杜顿 的子孙唱歌 ，以弹琴、鼓瑟、敲钹伴奏。他们供职的人数如下：
1CHR|25|2|亚萨 的儿子 撒刻 、 约瑟 、 尼探雅 、 亚萨利拉 ， 亚萨 的儿子都在 亚萨 的指导下，遵王的指示唱歌。
1CHR|25|3|属 耶杜顿 ， 耶杜顿 的儿子 基大利 、 西利 、 耶筛亚 、 示每 、 哈沙比雅 、 玛他提雅 共六人，都在他们父亲 耶杜顿 的指导下唱歌，以弹琴伴奏，称谢，颂赞耶和华。
1CHR|25|4|属 希幔 ， 希幔 的儿子是 布基雅 、 玛探雅 、 乌薛 、 细布业 、 耶利末 、 哈拿尼雅 、 哈拿尼 、 以利亚他 、 基大利提 、 罗幔提．以谢 、 约施比加沙 、 玛罗提 、 何提 、 玛哈秀 。
1CHR|25|5|这些都是 希幔 的儿子； 希幔 奉上帝之命作王的先见，吹角颂赞。上帝赐给 希幔 十四个儿子，三个女儿，
1CHR|25|6|他们都在父亲的指导下，在耶和华的殿唱歌，以敲钹、弹琴、鼓瑟伴奏，遵从王的指示，在上帝的殿里事奉。 亚萨 、 耶杜顿 、 希幔 ，
1CHR|25|7|他们和他们的弟兄学习颂赞耶和华，精通者的数目共有二百八十八人。
1CHR|25|8|这些人无论大小，为师的、为徒的，都一同抽签分了班次。
1CHR|25|9|抽签的时候，第一签抽到的是 亚萨 的儿子 约瑟 。第二是 基大利 ；他和他兄弟，以及儿子共十二人。
1CHR|25|10|第三是 撒刻 ，他儿子和他兄弟共十二人。
1CHR|25|11|第四是 伊洗利 ，他儿子和他兄弟共十二人。
1CHR|25|12|第五是 尼探雅 ，他儿子和他兄弟共十二人。
1CHR|25|13|第六是 布基雅 ，他儿子和他兄弟共十二人。
1CHR|25|14|第七是 耶萨利拉 ，他儿子和他兄弟共十二人。
1CHR|25|15|第八是 耶筛亚 ，他儿子和他兄弟共十二人。
1CHR|25|16|第九是 玛探雅 ，他儿子和他兄弟共十二人。
1CHR|25|17|第十是 示每 ，他儿子和他兄弟共十二人。
1CHR|25|18|第十一是 亚萨烈 ，他儿子和他兄弟共十二人。
1CHR|25|19|第十二是 哈沙比雅 ，他儿子和他兄弟共十二人。
1CHR|25|20|第十三是 书巴业 ，他儿子和他兄弟共十二人。
1CHR|25|21|第十四是 玛他提雅 ，他儿子和他兄弟共十二人。
1CHR|25|22|第十五是 耶列末 ，他儿子和他兄弟共十二人。
1CHR|25|23|第十六是 哈拿尼雅 ，他儿子和他兄弟共十二人。
1CHR|25|24|第十七是 约施比加沙 ，他儿子和他兄弟共十二人。
1CHR|25|25|第十八是 哈拿尼 ，他儿子和他兄弟共十二人。
1CHR|25|26|第十九是 玛罗提 ，他儿子和他兄弟共十二人。
1CHR|25|27|第二十是 以利亚他 ，他儿子和他兄弟共十二人。
1CHR|25|28|第二十一是 何提 ，他儿子和他兄弟共十二人。
1CHR|25|29|第二十二是 基大利提 ，他儿子和他兄弟共十二人。
1CHR|25|30|第二十三是 玛哈秀 ，他儿子和他兄弟共十二人。
1CHR|25|31|第二十四是 罗幔提．以谢 ，他儿子和他兄弟共十二人。
1CHR|26|1|门口守卫的班次如下： 可拉 族 以比雅撒 的子孙中，有 可利 的儿子 米施利米雅 。
1CHR|26|2|米施利米雅 的长子是 撒迦利亚 ，次子是 耶叠 ，三子是 西巴第雅 ，四子是 耶提聂 ，
1CHR|26|3|五子是 以拦 ，六子是 约哈难 ，七子是 以利约乃 。
1CHR|26|4|俄别．以东 的长子是 示玛雅 ，次子是 约萨拔 ，三子是 约亚 ，四子是 沙甲 ，五子是 拿坦业 ，
1CHR|26|5|六子是 亚米利 ，七子是 以萨迦 ，八子是 毗乌利太 ，因为上帝赐福给 俄别．以东 。
1CHR|26|6|他的儿子 示玛雅 生了几个儿子，都是大能的勇士，管理父亲的家。
1CHR|26|7|示玛雅 的儿子是 俄得尼 、 利法益 、 俄备得 、 以利萨巴 。 以利萨巴 的兄弟 以利户 和 西玛迦 是能人。
1CHR|26|8|这些都是 俄别．以东 的子孙，他们和他们的儿子，以及兄弟，都是善于办事的能人。属 俄别．以东 的共六十二人。
1CHR|26|9|米施利米雅 的儿子和兄弟都是能人，共十八人。
1CHR|26|10|米拉利 子孙中的 何萨 有几个儿子：为首的是 申利 ；他原不是长子，是他父亲立他为首的，
1CHR|26|11|次子是 希勒家 ，三子是 底巴利雅 ，四子是 撒迦利亚 。 何萨 的儿子和兄弟共十三人。
1CHR|26|12|这些是门口守卫的班次，各随他们的班长，与他们的兄弟一同在耶和华殿里按班供职。
1CHR|26|13|他们无论大小，都按着父系抽签，分守各门。
1CHR|26|14|抽到东门的是 示利米雅 ；他的儿子 撒迦利亚 是精明的谋士，抽到北门。
1CHR|26|15|俄别．以东 守南门，他的儿子守仓库。
1CHR|26|16|书聘 与 何萨 守西门，在靠近 沙利基 门、通往上去的街道上，守卫与守卫相对。
1CHR|26|17|东门有六个 利未 人 ，北门每日有四人，南门每日有四人，库房有两人轮流替换。
1CHR|26|18|至于走廊，在西面街道上有四人，在走廊上有两人。
1CHR|26|19|以上是 可拉 子孙和 米拉利 子孙门口守卫的班次。
1CHR|26|20|利未 人中有 亚希雅 管理上帝殿的库房和圣物的库房。
1CHR|26|21|拉但 子孙中， 革顺 族属 拉但 、作族长的是 革顺 族属 拉但 的 耶希伊利 。
1CHR|26|22|耶希伊利 的儿子 西坦 和他兄弟 约珥 管理耶和华殿的库房。
1CHR|26|23|暗兰 人、 以斯哈 人、 希伯伦 人、 乌薛 人也有职务。
1CHR|26|24|摩西 的孙子， 革舜 的儿子 细布业 管理库房。
1CHR|26|25|还有他的弟兄： 以利以谢 ， 以利以谢 的儿子 利哈比雅 ， 利哈比雅 的儿子 耶筛亚 ， 耶筛亚 的儿子 约兰 ， 约兰 的儿子 细基利 ， 细基利 的儿子 示罗密 。
1CHR|26|26|这 示罗密 和他的兄弟管理一切库房的圣物，就是 大卫 王和众族长、千夫长、百夫长，以及军官所分别为圣之物。
1CHR|26|27|他们把打仗时夺取的一些财物分别为圣，用来修造耶和华的殿。
1CHR|26|28|凡 撒母耳 先见、 基士 的儿子 扫罗 、 尼珥 的儿子 押尼珥 、 洗鲁雅 的儿子 约押 分别为圣的，一切分别为圣之物都归 示罗密 和他的兄弟掌管。
1CHR|26|29|以斯哈 人有 基拿尼雅 和他众儿子作官长和审判官，管理 以色列 对外的事务。
1CHR|26|30|希伯伦 人有 哈沙比雅 和他弟兄一千七百人，都是能人，在 约旦河 西监督 以色列 人，办理耶和华的一切工作和王的事务。
1CHR|26|31|希伯伦 人中有 耶利雅 作族长。 大卫 作王第四十年在各族各家从事寻访，在 基列 的 雅谢 ，从这族中发现大能的勇士。
1CHR|26|32|耶利雅 的弟兄有二千七百人，都是能人，又是族长； 大卫 王派他们在 吕便 人、 迦得 人、 玛拿西 半支派中管理上帝和王的一切事务。
1CHR|27|1|以色列 人的族长、千夫长、百夫长和官长都分配班次，每班二万四千人，整年按月轮流出入，按班次服事王。
1CHR|27|2|正月第一班的班长是 撒巴第业 的儿子 雅朔班 ；他班内有二万四千人。
1CHR|27|3|他是 法勒斯 的后裔，统管正月军队所有的官长。
1CHR|27|4|二月的班长是 亚何亚 人 朵代 ，他的班有总长 密基罗 ；他班内有二万四千人。
1CHR|27|5|三月第三班的班长是 耶何耶大 祭司长的儿子 比拿雅 ；他班内有二万四千人。
1CHR|27|6|这 比拿雅 是那三十人中的勇士，管理那三十人；他班内又有他儿子 暗米萨拔 。
1CHR|27|7|四月第四班的班长是 约押 的兄弟 亚撒黑 。接续他的是他儿子 西巴第雅 ；他班内有二万四千人。
1CHR|27|8|五月第五班的班长是 伊斯拉 人 珊合 ；他班内有二万四千人。
1CHR|27|9|六月第六班的班长是 提哥亚 人 益吉 的儿子 以拉 ；他班内有二万四千人。
1CHR|27|10|七月第七班的班长是 以法莲 族 比伦 人 希利斯 ；他班内有二万四千人。
1CHR|27|11|八月第八班的班长是 谢拉 族 户沙 人 西比该 ；他班内有二万四千人。
1CHR|27|12|九月第九班的班长是 便雅悯 族 亚拿突 人 亚比以谢 ；他班内有二万四千人。
1CHR|27|13|十月第十班的班长是 谢拉 族 尼陀法 人 玛哈莱 ；他班内有二万四千人。
1CHR|27|14|十一月第十一班的班长是 以法莲 族 比拉顿 人 比拿雅 ；他班内有二万四千人。
1CHR|27|15|十二月第十二班的班长是 俄陀聂 族 尼陀法 人 黑玳 ；他班内有二万四千人。
1CHR|27|16|管理 以色列 众支派的如下：管 吕便 人的是 细基利 的儿子 以利以谢 ；管 西缅 人的是 玛迦 的儿子 示法提雅 ；
1CHR|27|17|管 利未 的是 基摩利 的儿子 哈沙比雅 ；管 亚伦 子孙的是 撒督 ；
1CHR|27|18|管 犹大 的是 大卫 的一个哥哥 以利户 ；管 以萨迦 的是 米迦勒 的儿子 暗利 ；
1CHR|27|19|管 西布伦 的是 俄巴第雅 的儿子 伊施玛雅 ；管 拿弗他利 的是 亚斯列 的儿子 耶利摩 ；
1CHR|27|20|管 以法莲 的是 阿撒细雅 的儿子 何细亚 ；管 玛拿西 半支派的是 毗大雅 的儿子 约珥 ；
1CHR|27|21|管 基列 地 玛拿西 半支派的是 撒迦利亚 的儿子 易多 ；管 便雅悯 的是 押尼珥 的儿子 雅西业 ；
1CHR|27|22|管 但 的是 耶罗罕 的儿子 亚萨列 。以上是 以色列 众支派的领袖。
1CHR|27|23|以色列 人二十岁以下的， 大卫 没有记其数目；因耶和华曾应许，必加增 以色列 人如天上的星那样多。
1CHR|27|24|洗鲁雅 的儿子 约押 开始数点，却还没有数完。为了这事，烈怒临到 以色列 ，数点的数目也没有写在《大卫王记》上。
1CHR|27|25|管理王的库房的是 亚叠 的儿子 押斯马威 。管理田野、城镇、村庄、堡垒之仓库的是 乌西雅 的儿子 约拿单 。
1CHR|27|26|管理耕田种地的是 基绿 的儿子 以斯利 。
1CHR|27|27|管理葡萄园的是 拉玛 人 示每 。管理葡萄园酒窖的是 实弗米 人 撒巴底 。
1CHR|27|28|管理 谢非拉 橄榄树和桑树的是 基第利 人 巴勒．哈南 。管理油库的是 约阿施 。
1CHR|27|29|管理 沙仑 牧放牛群的是 沙仑 人 施提莱 。管理山谷牧养牛群的是 亚第莱 的儿子 沙法 。
1CHR|27|30|管理骆驼群的是 以实玛利 人 阿比勒 。管理驴群的是 米仑 人 耶希底亚 。管理羊群的是 夏甲 人 雅悉 。
1CHR|27|31|这些都是为 大卫 王管理产业的领袖。
1CHR|27|32|大卫 的叔父 约拿单 作谋士；这人有智慧，又作书记。 哈摩尼 的儿子 耶歇 陪伴王的众儿子。
1CHR|27|33|亚希多弗 作王的谋士。 亚基 人 户筛 作王的顾问。
1CHR|27|34|亚希多弗 之后，有 比拿雅 的儿子 耶何耶大 ，以及 亚比亚他 接续他。 约押 作王的元帅。
1CHR|28|1|大卫 召集 以色列 所有的领袖，各支派的领袖、轮班服事王的官长、千夫长、百夫长、掌管王和王子一切产业牲畜的、宫廷官员、勇士，和所有大能的勇士，都到 耶路撒冷 来。
1CHR|28|2|大卫 王站起来，说：“我的弟兄，我的百姓啊，请听我说！我心里本想建造殿宇，安放耶和华的约柜，作为我们上帝的脚凳，并且我已经预备了建造的材料。
1CHR|28|3|只是上帝对我说：‘你不可为我的名建造殿宇，因你是战士，流了人的血。’
1CHR|28|4|然而，耶和华－ 以色列 的上帝在我父的全家拣选我作 以色列 的王，直到永远。因他拣选 犹大 为领袖，在 犹大 家中拣选我父家，在我父的众儿子里喜悦我，立我作全 以色列 的王。
1CHR|28|5|耶和华赐我许多儿子，在我儿子中拣选我儿子 所罗门 坐耶和华国度的王位，治理 以色列 。
1CHR|28|6|耶和华对我说：‘你儿子 所罗门 必建造我的殿和院宇，因为我拣选他作我的子，我也必作他的父。
1CHR|28|7|他若恒久遵行我的诫命典章如今日一样，我就必坚定他的国，直到永远。’
1CHR|28|8|现今在 以色列 众人眼前，在耶和华的会中，在我们上帝的垂听下，你们务要遵行并寻求耶和华－你们上帝的一切诫命，如此你们就可以承受这美地，并留给你们的子孙，永远为业。
1CHR|28|9|“我儿 所罗门 哪，你当认识耶和华－你父的上帝，全心乐意地事奉他，因为耶和华鉴察众人的心，知道一切心思意念。你若寻求他，他必使你寻见；你若离弃他，他必永远丢弃你。
1CHR|28|10|现在你当谨慎，因耶和华拣选你建造殿宇作为圣所。你当刚强去做。”
1CHR|28|11|大卫 指示他儿子 所罗门 有关殿的走廊、屋子、库房、楼房、内殿和柜盖 之处的样式，
1CHR|28|12|被灵感动所得的一切样式：耶和华殿的院子、周围一切的房屋、上帝殿的库房和圣物库房；
1CHR|28|13|祭司和 利未 人的班次，耶和华殿里各样事奉的工作，耶和华殿里一切事奉用的器皿，
1CHR|28|14|以及各样事奉所用金器的重量，和各样事奉所用银器的重量，
1CHR|28|15|金灯台和金灯的重量，按每一个灯台和灯的重量；银灯台和银灯的重量，按每一个灯台和灯的重量，都按照每一个灯台的用途；
1CHR|28|16|每张供饼桌子的金子重量，和银桌子的银子重量，
1CHR|28|17|纯金的肉叉子、盘子，和壶的重量，金碗，按每个金碗的重量，和银碗，按每个银碗的重量，
1CHR|28|18|纯金香坛的重量，金基路伯座车的样式，基路伯张开翅膀，遮盖耶和华的约柜。
1CHR|28|19|大卫 说：“这一切，所有工作的样式，是耶和华用手写的文件使我明白的。”
1CHR|28|20|大卫 又对他儿子 所罗门 说：“你当刚强壮胆去做！不要惧怕，也不要惊惶，因为耶和华上帝，我的上帝与你同在。他必不撇下你，也不丢弃你，直到耶和华殿的工作都完毕。
1CHR|28|21|看哪，有祭司和 利未 人的班次，为要办理上帝殿各样的事务，又有擅长做各样事务的人，乐意在各样工作上帮助你，并且领袖和众百姓也都听从你的一切命令。”
1CHR|29|1|大卫 王对全会众说：“我儿子 所罗门 是上帝特选的，还年幼脆弱，但这工程浩大，因这殿不是为人，而是为耶和华上帝建造的。
1CHR|29|2|我为我上帝的殿已经尽力，预备金子做金器，银子做银器，铜做铜器，铁做铁器，木做木器，还有红玛瑙、可镶嵌的宝石、彩石、各样的宝石和许多大理石。
1CHR|29|3|此外，因我爱慕我上帝的殿，在预备建造圣殿的一切材料之外，又将我自己积蓄的金银献给我上帝的殿，
1CHR|29|4|就是三千他连得 俄斐 金子、七千他连得纯银，用来贴殿的墙；
1CHR|29|5|金子做金器，银子做银器，并藉工匠的手做一切的工。今日有谁愿意将自己献给耶和华呢？”
1CHR|29|6|于是，众族长和 以色列 各支派的领袖、千夫长、百夫长，以及监管王工作的官长，都乐意奉献。
1CHR|29|7|他们为上帝殿的工程献上五千他连得又一万达利克 金子，一万他连得银子，一万八千他连得铜，十万他连得铁。
1CHR|29|8|凡有宝石的都送入耶和华殿的库房，由 革顺 人 耶歇 的手管理。
1CHR|29|9|因这些人全心乐意献给耶和华，百姓就欢喜， 大卫 王也大大欢喜。
1CHR|29|10|大卫 在全会众眼前称颂耶和华； 大卫 说：“耶和华－ 以色列 的上帝，我们的父，你是应当称颂的，直到永永远远！
1CHR|29|11|耶和华啊，尊大、能力、荣耀、胜利、威严都是你的；天上地下的一切都是你的；耶和华啊，国度是你的，并且你为至高，为万有之首。
1CHR|29|12|丰富尊荣都从你而来，你也治理万物。在你手里有大能大力，你的手使人尊大强盛。
1CHR|29|13|我们的上帝啊，现在我们称谢你，赞美你荣耀之名！
1CHR|29|14|“我算什么，我的百姓算什么，竟然能够如此乐意奉献？因为万物都从你而来，我们把从你的手得来的献给你。
1CHR|29|15|我们在你面前是客旅，是寄居的，与我们的列祖一样。我们在世的日子如影子，没有盼望。
1CHR|29|16|耶和华－我们的上帝啊，我们预备这许多材料，要为你的圣名建造殿宇，都是从你的手而来，都是属你的。
1CHR|29|17|我的上帝啊，我知道你察验人心，喜悦正直；我以正直的心乐意献上这一切。现在我欢喜见你的百姓在此乐意奉献给你。
1CHR|29|18|耶和华－我们列祖 亚伯拉罕 、 以撒 、 以色列 的上帝啊，求你使你的百姓心中常存这样的心思意念，坚定他们的心归向你，
1CHR|29|19|又求你赐我儿子 所罗门 全心遵守你的命令、法度、律例，成就这一切的事，用我所预备的建造殿宇。”
1CHR|29|20|大卫 对全会众说：“你们应当称颂耶和华－你们的上帝。”于是全会众称颂耶和华－他们列祖的上帝，低头向耶和华和王下拜。
1CHR|29|21|次日，他们向耶和华献平安祭和燔祭，献一千头公牛，一千只公绵羊，一千只羔羊，以及同献的浇酒祭，并为 以色列 众人献许多的祭。
1CHR|29|22|那日，他们在耶和华面前吃喝，大大欢乐。 他们再次立 大卫 的儿子 所罗门 作王，膏他归耶和华作君王，又膏 撒督 作祭司。
1CHR|29|23|于是 所罗门 坐在耶和华所赐的王位上，接续他父亲 大卫 作王；他万事亨通，全 以色列 都听从他。
1CHR|29|24|众领袖和勇士，以及 大卫 王的众儿子，都顺服 所罗门 王。
1CHR|29|25|耶和华使 所罗门 在 以色列 众人眼前非常尊大，赐他君王的威严，胜过他以前任何一位 以色列 王。
1CHR|29|26|耶西 的儿子 大卫 作全 以色列 的王。
1CHR|29|27|他作 以色列 王的时期共四十年：在 希伯仑 作王七年，在 耶路撒冷 作王三十三年。
1CHR|29|28|他死的时候年纪老迈，日子满足，享尽荣华富贵。他的儿子 所罗门 接续他作王。
1CHR|29|29|大卫 王自始至终的事迹，看哪，都写在 撒母耳 先见的书上、 拿单 先知的书上和 迦得 先见的书上，
1CHR|29|30|包括他治国的一切和他英勇的事迹，以及他和 以色列 与世上列国所经历的事。
