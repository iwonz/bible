SONG|1|1|Соломонова Пісня над піснями.
SONG|1|2|Нехай він цілує мене поцілунками уст своїх, бо ліпші кохання твої від вина!
SONG|1|3|На запах оливи твої запашні, твоє ймення неначе олива розлита, тому діви кохають тебе!
SONG|1|4|Потягни ти мене за собою, біжім! Цар впровадив мене у палати свої, ми радіти та тішитись будемо тобою, згадаємо кохання твої, від вина приємніші, поправді кохають тебе!
SONG|1|5|Дочки єрусалимські, я чорна та гарна, немов ті намети кедарські, мов занавіси Соломонові!
SONG|1|6|Не дивіться на те, що смуглявенька я, бож сонце мене опалило, сини неньки моєї на мене розгнівалися, настановили мене сторожити виноградники, та свого виноградника власного не встерегла я!...
SONG|1|7|Скажи ж мені ти, кого покохала душа моя: Де ти пасеш? Де даєш ти спочити у спеку отарі? Пощо біля стад твоїх друзів я буду, немов та причинна?
SONG|1|8|Якщо ти не знаєш цього, вродливіша посеред жінок, то вийди собі за слідами отари, і випасуй при шатрах пастуших козлятка свої.
SONG|1|9|Я тебе прирівняв до лошиці в возах фараонових, о моя ти подруженько!
SONG|1|10|Гарні щічки твої поміж шнурами перел, а шийка твоя між разками намиста!
SONG|1|11|Ланцюжки золоті ми поробимо тобі разом із срібними кульками!
SONG|1|12|Доки цар при своєму столі, то мій нард видає свої пахощі.
SONG|1|13|Мій коханий для мене мов китиця мирри: спочиває між персами в мене!
SONG|1|14|Мій коханий для мене мов кипрове гроно в ен-ґедських садах-виноградах!
SONG|1|15|Яка ти прекрасна, моя ти подруженько, яка ти хороша! Твої очі немов голубині!
SONG|1|16|Який ти прекрасний, о мій ти коханий, який ти приємний! а ложе нам зелень!
SONG|1|17|Бруси наших домів то кедрини, стелі в нас кипариси!
SONG|2|1|Я саронська троянда, я долинна лілея!
SONG|2|2|Як лілея між тереном, так подруга моя поміж дівами!
SONG|2|3|Як та яблуня між лісовими деревами, так мій коханий поміж юнаками, його тіні жадала й сиділа я в ній, і його плід для мого піднебіння солодкий!
SONG|2|4|Він впровадив мене до винярні, а прапор його надо мною кохання!
SONG|2|5|Підкріпіте мене виноградовим печивом, освіжіть мене яблуками, бо я хвора з кохання!
SONG|2|6|Ліва рука його під головою моєю, правиця ж його пригортає мене!...
SONG|2|7|Заклинаю я вас, дочки єрусалимські, газелями чи польовими оленями, щоб ви не сполохали, й щоб не збудили кохання, аж доки йому до вподоби!...
SONG|2|8|Голос мого коханого!... Ось він іде, ось він скаче горами, по пагірках вистрибує...
SONG|2|9|Мій коханий подібний до сарни чи до молодого оленя. Он стоїть він у нас за стіною, зазирає у вікна, заглядає у ґрати...
SONG|2|10|Мій коханий озвався й промовив до мене: Уставай же, подруго моя, моя красна, й до мене ходи!
SONG|2|11|Бо оце проминула пора дощова, дощ ущух, перейшов собі він.
SONG|2|12|Показались квітки на землі, пора соловейка настала, і голос горлиці в нашому краї лунає!
SONG|2|13|Фіґа випустила свої ранні плоди, і розцвілі виноградини пахощі видали. Уставай же, подруго моя, моя красна, й до мене ходи!
SONG|2|14|Голубко моя у розщілинах скельних, у бескіднім сховку, дай побачити мені твоє личко, дай почути мені голосок твій, бо голос твій милий, а личко твоє уродливе!
SONG|2|15|Ловіть нам лисиці, лисинята маленькі, що ушкоджують нам виноградники, виноградники ж наші у цвіті!
SONG|2|16|Мій коханий він мій, я ж його, він пасе між лілеями!
SONG|2|17|Поки день прохолоду навіє, а тіні втечуть, вернись, мій коханий, стань подібний до сарни чи до молодого оленя в пахучих горах!
SONG|3|1|По ночах на ложі своїм я шукала того, кого покохала душа моя... Шукала його, та його не знайшла...
SONG|3|2|Хай устану й нехай я пройдуся по місті, хай на вулицях та на майданах того пошукаю, кого покохала душа моя! Шукала його, та його не знайшла...
SONG|3|3|Спіткали мене сторожі, що по місті проходять... Чи не бачили часом того, кого покохала душа моя?
SONG|3|4|Небагато пройшла я від них, та й знайшла я того, кого покохала душа моя: схопила його, й не пустила його, аж поки його не ввела у дім неньки своєї, та в кімнату тієї, що в утробі носила мене!...
SONG|3|5|Заклинаю я вас, дочки єрусалимські, газелями чи польовими оленями, щоб ви не сполохали, щоб не збудили кохання, аж доки йому до вподоби!...
SONG|3|6|Хто вона, що виходить із пустині, немов стовпи диму, окурена миррою й ладаном, всілякими пахощами продавця?
SONG|3|7|Ось ложе його, Соломонове, шістдесят лицарів навколо нього, із лицарів славних Ізраїлевих!
SONG|3|8|Усі вони мають меча, усі вправні в бою, кожен має свого меча при своєму стегні проти страху нічного.
SONG|3|9|Ноші зробив собі цар Соломон із ливанських дерев:
SONG|3|10|стовпці їхні зробив він із срібла, а їхне опертя золоте, пурпурове сидіння, їхня середина вистелена коханням дочок єрусалимських!...
SONG|3|11|Підіть і побачте, о дочки сіонські, царя Соломона в вінку, що ним мати його увінчала його в день весілля його та в день радости серця його!
SONG|4|1|Яка ти прекрасна, моя ти подруженько, яка ти хороша! Твої оченятка, немов ті голубки, глядять з-за серпанку твого! Твої коси немов стадо кіз, що хвилями сходять з гори Гілеадської!
SONG|4|2|Твої зубки немов та отара овець пообстриганих, що з купелю вийшли, що котять близнята, і між ними немає неплідної...
SONG|4|3|Твої губки немов кармазинова нитка, твої устонька красні, мов частина гранатного яблука скроня твоя за серпанком твоїм!
SONG|4|4|Твоя шия немов та Давидова башта, на зброю збудована: тисяча щитів повішена в ній, усе щити лицарів!
SONG|4|5|Два перса твої мов ті двоє близнят молодих у газелі, що випасуються між лілеями...
SONG|4|6|Поки день прохолоду навіє, а тіні втечуть, піду я собі на ту миррину гору й на пагірок ладану...
SONG|4|7|Уся ти прекрасна, моя ти подруженько, і плями нема на тобі!
SONG|4|8|Зо мною з Лівану, моя наречена, зо мною з Лівану ти підеш! Споглянеш з вершини Амани, з вершини Сеніру й Гермону, з леговища левів, з леопардових гір.
SONG|4|9|Забрала ти серце мені, моя сестро, моя наречена, забрала ти серце мені самим очком своїм, разочком одненьким намиста свого!...
SONG|4|10|Яке любе кохання твоє, о сестрице моя, наречена! Скільки ліпше кохання твоє за вино, а запашність олив твоїх за всі пахощі!...
SONG|4|11|Уста твої крапають мед щільниковий, моя наречена, мед і молоко під твоїм язичком, а пахощ одежі твоєї як ліванські ті пахощі!
SONG|4|12|Замкнений садок то сестриця моя, наречена моя замкнений садок, джерело запечатане...
SONG|4|13|Лоно твоє сад гранатових яблук з плодом досконалим, кипри із нардами,
SONG|4|14|нард і шафран, пахуча тростина й кориця з усіма деревами ладану, мирра й алое зо всіма найзапашнішими пахощами,
SONG|4|15|ти джерело садкове, криниця живої води, та тієї, що плине з Ливану!...
SONG|4|16|Прокинься, о вітре з півночі, і прилинь, вітре з полудня, повій на садок мій: нехай потечуть його пахощі! Хай коханий мій прийде до саду свого, і нехай споживе плід найкращий його!...
SONG|5|1|Прийшов я до саду свого, о сестро моя, наречена! Збираю я мирру свою із бальзамом своїм, споживаю свого стільника разом із медом своїм, п'ю вино я своє зо своїм молоком!... Споживайте, співдрузі, пийте до схочу, кохані!
SONG|5|2|Я сплю, моє ж серце чуває... Ось голос мого коханого!... Стукає... Відчини мені, сестро моя, о моя ти подруженько, голубко моя, моя чиста, бо росою покрилася вся моя голова, мої кучері краплями ночі!...
SONG|5|3|Зняла я одежу свою, як знову її надягну? Помила я ніжки свої, як же їх занечищу?...
SONG|5|4|Мій коханий простяг свою руку крізь отвір, і нутро моє схвилювалось від нього!...
SONG|5|5|Встала я відчинити своєму коханому, а з рук моїх капала мирра, і мирра текла на засувки замка з моїх пальців...
SONG|5|6|Відчинила своєму коханому, а коханий мій зник, відійшов!... Душі не ставало в мені, як він говорив... Я шукала його, та його не знайшла... Я гукала його, та він не відізвався до мене...
SONG|5|7|Стріли мене сторожі, що ходять по місті, набили мене, завдали мені рани... Здерли з мене моє покривало, сторожі міських мурів!
SONG|5|8|Заклинаю я вас, дочки єрусалимські, як мого коханого стрінете ви, що йому повісте? Що я хвора з кохання!
SONG|5|9|Чим коханий твій кращий від інших коханих, вродливіша з жінок? Чим коханий твій кращий від інших коханих, що так заклинаєш ти нас?
SONG|5|10|Коханий мій білий й рум'яний, визначніший він від десяти тисяч інших...
SONG|5|11|Голова його щиреє золото, його кучері пальмове віття, чорні, як ворон...
SONG|5|12|Його очі немов голубки над джерелами водними, у молоці повимивані, що над повним струмком посідали!
SONG|5|13|Його личка як грядка бальзаму, немов квітники запашні! Його губи лілеї, з яких капає мирра текуча!
SONG|5|14|Його руки стовпці золоті, повисаджувані хризолітом, а лоно його твір мистецький з слонової кости, покритий сапфірами!
SONG|5|15|Його стегна стовпи мармурові, поставлені на золотії підстави! Його вигляд немов той Ливан, він юнак як ті кедри!
SONG|5|16|Уста його солодощі, і він увесь пожадання... Оце мій коханий, й оце мій дружок, дочки єрусалимські!
SONG|6|1|Куди твій коханий пішов, о найвродливіша з жінок? Куди спрямував твій коханий? Бо ми пошукаємо його із тобою.
SONG|6|2|Мій коханий пішов до садочка свого, в квітники запашні, щоб пасти в садках і збирати лілеї.
SONG|6|3|Я належу своєму коханому, а мені мій коханий, що пасе між лілеями!
SONG|6|4|Ти прекрасна, моя ти подруженько, мов та Тірца, ти хороша, як Єрусалим, ти грізна, як війська з прапорами!
SONG|6|5|Відверни ти свої оченята від мене, бо вони непокоять мене! Твої коси немов стадо кіз, що хвилями сходять з того Гілеаду!
SONG|6|6|Твої зуби немов та отара овець, що з купелю вийшли, що котять близнята, і між ними немає неплідної!
SONG|6|7|Мов частина гранатного яблука скроня твоя за серпанком твоїм!
SONG|6|8|Шістдесят є цариць, і вісімдесят є наложниць, а дівчатам немає числа,
SONG|6|9|та єдина вона ця голубка моя, моя чиста! У неньки своєї вона одиначка, обрана вона у своєї родительки! Як бачили дочки Сіону її, то щасливою звали її, цариці й наложниці то вихваляли її:
SONG|6|10|Хто це така, що вона виглядає, немов та досвітня зоря, прекрасна, як місяць, як сонце ясна, як полки з прапорами грізна?
SONG|6|11|Зійшла я в оріховий сад, щоб поглянути на пуп'яночки при потоці, щоб побачити там, чи зацвів виноград, чи гранатові яблуні порозцвітали?
SONG|6|12|І не зчулася я, як мене посадила душа моя між колесниці моєї дружини бояр...
SONG|6|13|(7-1) Вернися, вернись, Суламітко! Вернися, вернися, нехай ми на тебе надивимось! Чого вам дивитися на Суламітку, немов би на танець військовий?
SONG|7|1|(7-2) Хороші які стали ноги твої в черевичках, князівно моя! Заокруглення стегон твоїх мов намисто, руками мистецькими виточене!
SONG|7|2|(7-3) Твоє лоно немов круглоточена чаша, в якій не забракне вина запашного! Твій живіт сніп пшениці, оточений тими лілеями!
SONG|7|3|(7-4) Два перса твої немов двоє сарняток близнят!
SONG|7|4|(7-5) Твоя шия як башта із кости слонової, твої очі озерця в Хешбоні при брамі того Бат-Рабіму, в тебе ніс немов башта ливанська, що дивиться все в бік Дамаску!
SONG|7|5|(7-6) Голівка твоя на тобі мов Кармел, а коса на голівці твоїй немов пурпур, полонений цар тими кучерями!
SONG|7|6|(7-7) Яка ти прекрасна й приємна яка, о кохання в розкошах!
SONG|7|7|(7-8) Став подібний до пальми твій стан, твої ж перса до грон виноградних!
SONG|7|8|(7-9) Я подумав: виберуся на цю пальму, схоплюся за віття її, і нехай стануть перса твої, немов виноградні ті грона, а пахощ дихання твого як яблука!...
SONG|7|9|(7-10) А уста твої як найліпше вино: простує воно до мого коханого, чинить промовистими й уста сплячих!
SONG|7|10|(7-11) Я належу своєму коханому, а його пожадання до мене!
SONG|7|11|(7-12) Ходи ж, мій коханий, та вийдемо в поле, переночуємо в селах!
SONG|7|12|(7-13) Устанемо рано, й ходім у сади-виногради, подивимося, чи зацвів виноград, чи квітки розцвілись, чи гранатові яблуні порозцвітали?... Там кохання своє тобі дам!
SONG|7|13|(7-14) Видадуть пах мандрагори, при наших же входах всілякі коштовні плоди, нові та старі, що я їх заховала для тебе, коханий ти мій!
SONG|8|1|О, коли б ти мені був за брата, що перса ссав в нені моєї, коли б стріла тебе я на вулиці, цілувала б тебе, і ніхто мені не докоряв би!
SONG|8|2|Повела б я тебе й привела б у дім нені своєї: ти навчав би мене, я б тебе напоїла вином запашним, соком гранатових яблук своїх!
SONG|8|3|Ліва рука його під головою моєю, правиця ж його пригортає мене!...
SONG|8|4|Заклинаю я вас, дочки єрусалимські, нащо б сполохали, й нащо б збудили кохання, аж доки йому до вподоби!
SONG|8|5|Хто вона, що виходить із пустині, спираючися на свого коханого? Під яблунею я збудила тебе, там повила тебе мати твоя, там тебе повила твоя породителька!
SONG|8|6|Поклади ти мене, як печатку на серце своє, як печать на рамено своє, бо сильне кохання, як смерть, заздрощі непереможні, немов той шеол, його жар жар огню, воно полум'я Господа!
SONG|8|7|Води великі не зможуть згасити кохання, ані ріки його не заллють! Коли б хто давав за кохання маєток увесь свого дому, то ним погордили б зовсім!...
SONG|8|8|Є сестра в нас мала, й перс у неї нема ще. Що зробимо нашій сестричці в той день, коли сватати будуть її?
SONG|8|9|Якщо вона мур, забороло із срібла збудуємо на ній, а якщо вона двері обкладемо кедровою дошкою їх...
SONG|8|10|Я мур, мої ж перса як башти, тоді я була в його очах мов та, яка спокій провадить...
SONG|8|11|Виноградника мав Соломон у Баал-Гамоні, виноградника він віддавав сторожам, щоб кожен приносив за плід його тисячу срібла.
SONG|8|12|Але мій виноградник, що маю його, при мені! Тобі, Соломоне, хай буде та тисяча, а сторожам його плоду дві сотні!
SONG|8|13|О ти, що сидиш у садках, друзі твої прислухаються до твого голосу: дай почути його і мені!
SONG|8|14|Утікай, мій коханий, і станься подібний до сарни собі, чи до молодого оленя у бальзамових горах!
