2KGS|1|1|After Ahab's death, Moab rebelled against Israel.
2KGS|1|2|Now Ahaziah had fallen through the lattice of his upper room in Samaria and injured himself. So he sent messengers, saying to them, "Go and consult Baal-Zebub, the god of Ekron, to see if I will recover from this injury."
2KGS|1|3|But the angel of the LORD said to Elijah the Tishbite, "Go up and meet the messengers of the king of Samaria and ask them, 'Is it because there is no God in Israel that you are going off to consult Baal-Zebub, the god of Ekron?'
2KGS|1|4|Therefore this is what the LORD says: 'You will not leave the bed you are lying on. You will certainly die!'" So Elijah went.
2KGS|1|5|When the messengers returned to the king, he asked them, "Why have you come back?"
2KGS|1|6|"A man came to meet us," they replied. "And he said to us, 'Go back to the king who sent you and tell him, "This is what the LORD says: Is it because there is no God in Israel that you are sending men to consult Baal-Zebub, the god of Ekron? Therefore you will not leave the bed you are lying on. You will certainly die!"'"
2KGS|1|7|The king asked them, "What kind of man was it who came to meet you and told you this?"
2KGS|1|8|They replied, "He was a man with a garment of hair and with a leather belt around his waist." The king said, "That was Elijah the Tishbite."
2KGS|1|9|Then he sent to Elijah a captain with his company of fifty men. The captain went up to Elijah, who was sitting on the top of a hill, and said to him, "Man of God, the king says, 'Come down!'"
2KGS|1|10|Elijah answered the captain, "If I am a man of God, may fire come down from heaven and consume you and your fifty men!" Then fire fell from heaven and consumed the captain and his men.
2KGS|1|11|At this the king sent to Elijah another captain with his fifty men. The captain said to him, "Man of God, this is what the king says, 'Come down at once!'"
2KGS|1|12|"If I am a man of God," Elijah replied, "may fire come down from heaven and consume you and your fifty men!" Then the fire of God fell from heaven and consumed him and his fifty men.
2KGS|1|13|So the king sent a third captain with his fifty men. This third captain went up and fell on his knees before Elijah. "Man of God," he begged, "please have respect for my life and the lives of these fifty men, your servants!
2KGS|1|14|See, fire has fallen from heaven and consumed the first two captains and all their men. But now have respect for my life!"
2KGS|1|15|The angel of the LORD said to Elijah, "Go down with him; do not be afraid of him." So Elijah got up and went down with him to the king.
2KGS|1|16|He told the king, "This is what the LORD says: Is it because there is no God in Israel for you to consult that you have sent messengers to consult Baal-Zebub, the god of Ekron? Because you have done this, you will never leave the bed you are lying on. You will certainly die!"
2KGS|1|17|So he died, according to the word of the LORD that Elijah had spoken. Because Ahaziah had no son, Joram succeeded him as king in the second year of Jehoram son of Jehoshaphat king of Judah.
2KGS|1|18|As for all the other events of Ahaziah's reign, and what he did, are they not written in the book of the annals of the kings of Israel?
2KGS|2|1|When the LORD was about to take Elijah up to heaven in a whirlwind, Elijah and Elisha were on their way from Gilgal.
2KGS|2|2|Elijah said to Elisha, "Stay here; the LORD has sent me to Bethel." But Elisha said, "As surely as the LORD lives and as you live, I will not leave you." So they went down to Bethel.
2KGS|2|3|The company of the prophets at Bethel came out to Elisha and asked, "Do you know that the LORD is going to take your master from you today?Yes, I know," Elisha replied, "but do not speak of it."
2KGS|2|4|Then Elijah said to him, "Stay here, Elisha; the LORD has sent me to Jericho." And he replied, "As surely as the LORD lives and as you live, I will not leave you." So they went to Jericho.
2KGS|2|5|The company of the prophets at Jericho went up to Elisha and asked him, "Do you know that the LORD is going to take your master from you today?Yes, I know," he replied, "but do not speak of it."
2KGS|2|6|Then Elijah said to him, "Stay here; the LORD has sent me to the Jordan." And he replied, "As surely as the LORD lives and as you live, I will not leave you." So the two of them walked on.
2KGS|2|7|Fifty men of the company of the prophets went and stood at a distance, facing the place where Elijah and Elisha had stopped at the Jordan.
2KGS|2|8|Elijah took his cloak, rolled it up and struck the water with it. The water divided to the right and to the left, and the two of them crossed over on dry ground.
2KGS|2|9|When they had crossed, Elijah said to Elisha, "Tell me, what can I do for you before I am taken from you?Let me inherit a double portion of your spirit," Elisha replied.
2KGS|2|10|"You have asked a difficult thing," Elijah said, "yet if you see me when I am taken from you, it will be yours-otherwise not."
2KGS|2|11|As they were walking along and talking together, suddenly a chariot of fire and horses of fire appeared and separated the two of them, and Elijah went up to heaven in a whirlwind.
2KGS|2|12|Elisha saw this and cried out, "My father! My father! The chariots and horsemen of Israel!" And Elisha saw him no more. Then he took hold of his own clothes and tore them apart.
2KGS|2|13|He picked up the cloak that had fallen from Elijah and went back and stood on the bank of the Jordan.
2KGS|2|14|Then he took the cloak that had fallen from him and struck the water with it. "Where now is the LORD, the God of Elijah?" he asked. When he struck the water, it divided to the right and to the left, and he crossed over.
2KGS|2|15|The company of the prophets from Jericho, who were watching, said, "The spirit of Elijah is resting on Elisha." And they went to meet him and bowed to the ground before him.
2KGS|2|16|"Look," they said, "we your servants have fifty able men. Let them go and look for your master. Perhaps the Spirit of the LORD has picked him up and set him down on some mountain or in some valley.No," Elisha replied, "do not send them."
2KGS|2|17|But they persisted until he was too ashamed to refuse. So he said, "Send them." And they sent fifty men, who searched for three days but did not find him.
2KGS|2|18|When they returned to Elisha, who was staying in Jericho, he said to them, "Didn't I tell you not to go?"
2KGS|2|19|The men of the city said to Elisha, "Look, our lord, this town is well situated, as you can see, but the water is bad and the land is unproductive."
2KGS|2|20|"Bring me a new bowl," he said, "and put salt in it." So they brought it to him.
2KGS|2|21|Then he went out to the spring and threw the salt into it, saying, "This is what the LORD says: 'I have healed this water. Never again will it cause death or make the land unproductive.'"
2KGS|2|22|And the water has remained wholesome to this day, according to the word Elisha had spoken.
2KGS|2|23|From there Elisha went up to Bethel. As he was walking along the road, some youths came out of the town and jeered at him. "Go on up, you baldhead!" they said. "Go on up, you baldhead!"
2KGS|2|24|He turned around, looked at them and called down a curse on them in the name of the LORD. Then two bears came out of the woods and mauled forty-two of the youths.
2KGS|2|25|And he went on to Mount Carmel and from there returned to Samaria.
2KGS|3|1|Joram son of Ahab became king of Israel in Samaria in the eighteenth year of Jehoshaphat king of Judah, and he reigned twelve years.
2KGS|3|2|He did evil in the eyes of the LORD, but not as his father and mother had done. He got rid of the sacred stone of Baal that his father had made.
2KGS|3|3|Nevertheless he clung to the sins of Jeroboam son of Nebat, which he had caused Israel to commit; he did not turn away from them.
2KGS|3|4|Now Mesha king of Moab raised sheep, and he had to supply the king of Israel with a hundred thousand lambs and with the wool of a hundred thousand rams.
2KGS|3|5|But after Ahab died, the king of Moab rebelled against the king of Israel.
2KGS|3|6|So at that time King Joram set out from Samaria and mobilized all Israel.
2KGS|3|7|He also sent this message to Jehoshaphat king of Judah: "The king of Moab has rebelled against me. Will you go with me to fight against Moab?I will go with you," he replied. "I am as you are, my people as your people, my horses as your horses."
2KGS|3|8|"By what route shall we attack?" he asked. "Through the Desert of Edom," he answered.
2KGS|3|9|So the king of Israel set out with the king of Judah and the king of Edom. After a roundabout march of seven days, the army had no more water for themselves or for the animals with them.
2KGS|3|10|"What!" exclaimed the king of Israel. "Has the LORD called us three kings together only to hand us over to Moab?"
2KGS|3|11|But Jehoshaphat asked, "Is there no prophet of the LORD here, that we may inquire of the LORD through him?" An officer of the king of Israel answered, "Elisha son of Shaphat is here. He used to pour water on the hands of Elijah. "
2KGS|3|12|Jehoshaphat said, "The word of the LORD is with him." So the king of Israel and Jehoshaphat and the king of Edom went down to him.
2KGS|3|13|Elisha said to the king of Israel, "What do we have to do with each other? Go to the prophets of your father and the prophets of your mother.No," the king of Israel answered, "because it was the LORD who called us three kings together to hand us over to Moab."
2KGS|3|14|Elisha said, "As surely as the LORD Almighty lives, whom I serve, if I did not have respect for the presence of Jehoshaphat king of Judah, I would not look at you or even notice you.
2KGS|3|15|But now bring me a harpist." While the harpist was playing, the hand of the LORD came upon Elisha
2KGS|3|16|and he said, "This is what the LORD says: Make this valley full of ditches.
2KGS|3|17|For this is what the LORD says: You will see neither wind nor rain, yet this valley will be filled with water, and you, your cattle and your other animals will drink.
2KGS|3|18|This is an easy thing in the eyes of the LORD; he will also hand Moab over to you.
2KGS|3|19|You will overthrow every fortified city and every major town. You will cut down every good tree, stop up all the springs, and ruin every good field with stones."
2KGS|3|20|The next morning, about the time for offering the sacrifice, there it was-water flowing from the direction of Edom! And the land was filled with water.
2KGS|3|21|Now all the Moabites had heard that the kings had come to fight against them; so every man, young and old, who could bear arms was called up and stationed on the border.
2KGS|3|22|When they got up early in the morning, the sun was shining on the water. To the Moabites across the way, the water looked red-like blood.
2KGS|3|23|"That's blood!" they said. "Those kings must have fought and slaughtered each other. Now to the plunder, Moab!"
2KGS|3|24|But when the Moabites came to the camp of Israel, the Israelites rose up and fought them until they fled. And the Israelites invaded the land and slaughtered the Moabites.
2KGS|3|25|They destroyed the towns, and each man threw a stone on every good field until it was covered. They stopped up all the springs and cut down every good tree. Only Kir Hareseth was left with its stones in place, but men armed with slings surrounded it and attacked it as well.
2KGS|3|26|When the king of Moab saw that the battle had gone against him, he took with him seven hundred swordsmen to break through to the king of Edom, but they failed.
2KGS|3|27|Then he took his firstborn son, who was to succeed him as king, and offered him as a sacrifice on the city wall. The fury against Israel was great; they withdrew and returned to their own land.
2KGS|4|1|The wife of a man from the company of the prophets cried out to Elisha, "Your servant my husband is dead, and you know that he revered the LORD. But now his creditor is coming to take my two boys as his slaves."
2KGS|4|2|Elisha replied to her, "How can I help you? Tell me, what do you have in your house?Your servant has nothing there at all," she said, "except a little oil."
2KGS|4|3|Elisha said, "Go around and ask all your neighbors for empty jars. Don't ask for just a few.
2KGS|4|4|Then go inside and shut the door behind you and your sons. Pour oil into all the jars, and as each is filled, put it to one side."
2KGS|4|5|She left him and afterward shut the door behind her and her sons. They brought the jars to her and she kept pouring.
2KGS|4|6|When all the jars were full, she said to her son, "Bring me another one." But he replied, "There is not a jar left." Then the oil stopped flowing.
2KGS|4|7|She went and told the man of God, and he said, "Go, sell the oil and pay your debts. You and your sons can live on what is left."
2KGS|4|8|One day Elisha went to Shunem. And a well-to-do woman was there, who urged him to stay for a meal. So whenever he came by, he stopped there to eat.
2KGS|4|9|She said to her husband, "I know that this man who often comes our way is a holy man of God.
2KGS|4|10|Let's make a small room on the roof and put in it a bed and a table, a chair and a lamp for him. Then he can stay there whenever he comes to us."
2KGS|4|11|One day when Elisha came, he went up to his room and lay down there.
2KGS|4|12|He said to his servant Gehazi, "Call the Shunammite." So he called her, and she stood before him.
2KGS|4|13|Elisha said to him, "Tell her, 'You have gone to all this trouble for us. Now what can be done for you? Can we speak on your behalf to the king or the commander of the army?'" She replied, "I have a home among my own people."
2KGS|4|14|"What can be done for her?" Elisha asked. Gehazi said, "Well, she has no son and her husband is old."
2KGS|4|15|Then Elisha said, "Call her." So he called her, and she stood in the doorway.
2KGS|4|16|"About this time next year," Elisha said, "you will hold a son in your arms.No, my lord," she objected. "Don't mislead your servant, O man of God!"
2KGS|4|17|But the woman became pregnant, and the next year about that same time she gave birth to a son, just as Elisha had told her.
2KGS|4|18|The child grew, and one day he went out to his father, who was with the reapers.
2KGS|4|19|"My head! My head!" he said to his father. His father told a servant, "Carry him to his mother."
2KGS|4|20|After the servant had lifted him up and carried him to his mother, the boy sat on her lap until noon, and then he died.
2KGS|4|21|She went up and laid him on the bed of the man of God, then shut the door and went out.
2KGS|4|22|She called her husband and said, "Please send me one of the servants and a donkey so I can go to the man of God quickly and return."
2KGS|4|23|"Why go to him today?" he asked. "It's not the New Moon or the Sabbath.It's all right," she said.
2KGS|4|24|She saddled the donkey and said to her servant, "Lead on; don't slow down for me unless I tell you."
2KGS|4|25|So she set out and came to the man of God at Mount Carmel. When he saw her in the distance, the man of God said to his servant Gehazi, "Look! There's the Shunammite!
2KGS|4|26|Run to meet her and ask her, 'Are you all right? Is your husband all right? Is your child all right?' Everything is all right," she said.
2KGS|4|27|When she reached the man of God at the mountain, she took hold of his feet. Gehazi came over to push her away, but the man of God said, "Leave her alone! She is in bitter distress, but the LORD has hidden it from me and has not told me why."
2KGS|4|28|"Did I ask you for a son, my lord?" she said. "Didn't I tell you, 'Don't raise my hopes'?"
2KGS|4|29|Elisha said to Gehazi, "Tuck your cloak into your belt, take my staff in your hand and run. If you meet anyone, do not greet him, and if anyone greets you, do not answer. Lay my staff on the boy's face."
2KGS|4|30|But the child's mother said, "As surely as the LORD lives and as you live, I will not leave you." So he got up and followed her.
2KGS|4|31|Gehazi went on ahead and laid the staff on the boy's face, but there was no sound or response. So Gehazi went back to meet Elisha and told him, "The boy has not awakened."
2KGS|4|32|When Elisha reached the house, there was the boy lying dead on his couch.
2KGS|4|33|He went in, shut the door on the two of them and prayed to the LORD.
2KGS|4|34|Then he got on the bed and lay upon the boy, mouth to mouth, eyes to eyes, hands to hands. As he stretched himself out upon him, the boy's body grew warm.
2KGS|4|35|Elisha turned away and walked back and forth in the room and then got on the bed and stretched out upon him once more. The boy sneezed seven times and opened his eyes.
2KGS|4|36|Elisha summoned Gehazi and said, "Call the Shunammite." And he did. When she came, he said, "Take your son."
2KGS|4|37|She came in, fell at his feet and bowed to the ground. Then she took her son and went out.
2KGS|4|38|Elisha returned to Gilgal and there was a famine in that region. While the company of the prophets was meeting with him, he said to his servant, "Put on the large pot and cook some stew for these men."
2KGS|4|39|One of them went out into the fields to gather herbs and found a wild vine. He gathered some of its gourds and filled the fold of his cloak. When he returned, he cut them up into the pot of stew, though no one knew what they were.
2KGS|4|40|The stew was poured out for the men, but as they began to eat it, they cried out, "O man of God, there is death in the pot!" And they could not eat it.
2KGS|4|41|Elisha said, "Get some flour." He put it into the pot and said, "Serve it to the people to eat." And there was nothing harmful in the pot.
2KGS|4|42|A man came from Baal Shalishah, bringing the man of God twenty loaves of barley bread baked from the first ripe grain, along with some heads of new grain. "Give it to the people to eat," Elisha said.
2KGS|4|43|"How can I set this before a hundred men?" his servant asked. But Elisha answered, "Give it to the people to eat. For this is what the LORD says: 'They will eat and have some left over.'"
2KGS|4|44|Then he set it before them, and they ate and had some left over, according to the word of the LORD.
2KGS|5|1|Now Naaman was commander of the army of the king of Aram. He was a great man in the sight of his master and highly regarded, because through him the LORD had given victory to Aram. He was a valiant soldier, but he had leprosy.
2KGS|5|2|Now bands from Aram had gone out and had taken captive a young girl from Israel, and she served Naaman's wife.
2KGS|5|3|She said to her mistress, "If only my master would see the prophet who is in Samaria! He would cure him of his leprosy."
2KGS|5|4|Naaman went to his master and told him what the girl from Israel had said.
2KGS|5|5|"By all means, go," the king of Aram replied. "I will send a letter to the king of Israel." So Naaman left, taking with him ten talents of silver, six thousand shekels of gold and ten sets of clothing.
2KGS|5|6|The letter that he took to the king of Israel read: "With this letter I am sending my servant Naaman to you so that you may cure him of his leprosy."
2KGS|5|7|As soon as the king of Israel read the letter, he tore his robes and said, "Am I God? Can I kill and bring back to life? Why does this fellow send someone to me to be cured of his leprosy? See how he is trying to pick a quarrel with me!"
2KGS|5|8|When Elisha the man of God heard that the king of Israel had torn his robes, he sent him this message: "Why have you torn your robes? Have the man come to me and he will know that there is a prophet in Israel."
2KGS|5|9|So Naaman went with his horses and chariots and stopped at the door of Elisha's house.
2KGS|5|10|Elisha sent a messenger to say to him, "Go, wash yourself seven times in the Jordan, and your flesh will be restored and you will be cleansed."
2KGS|5|11|But Naaman went away angry and said, "I thought that he would surely come out to me and stand and call on the name of the LORD his God, wave his hand over the spot and cure me of my leprosy.
2KGS|5|12|Are not Abana and Pharpar, the rivers of Damascus, better than any of the waters of Israel? Couldn't I wash in them and be cleansed?" So he turned and went off in a rage.
2KGS|5|13|Naaman's servants went to him and said, "My father, if the prophet had told you to do some great thing, would you not have done it? How much more, then, when he tells you, 'Wash and be cleansed'!"
2KGS|5|14|So he went down and dipped himself in the Jordan seven times, as the man of God had told him, and his flesh was restored and became clean like that of a young boy.
2KGS|5|15|Then Naaman and all his attendants went back to the man of God. He stood before him and said, "Now I know that there is no God in all the world except in Israel. Please accept now a gift from your servant."
2KGS|5|16|The prophet answered, "As surely as the LORD lives, whom I serve, I will not accept a thing." And even though Naaman urged him, he refused.
2KGS|5|17|"If you will not," said Naaman, "please let me, your servant, be given as much earth as a pair of mules can carry, for your servant will never again make burnt offerings and sacrifices to any other god but the LORD.
2KGS|5|18|But may the LORD forgive your servant for this one thing: When my master enters the temple of Rimmon to bow down and he is leaning on my arm and I bow there also-when I bow down in the temple of Rimmon, may the LORD forgive your servant for this."
2KGS|5|19|"Go in peace," Elisha said. After Naaman had traveled some distance,
2KGS|5|20|Gehazi, the servant of Elisha the man of God, said to himself, "My master was too easy on Naaman, this Aramean, by not accepting from him what he brought. As surely as the LORD lives, I will run after him and get something from him."
2KGS|5|21|So Gehazi hurried after Naaman. When Naaman saw him running toward him, he got down from the chariot to meet him. "Is everything all right?" he asked.
2KGS|5|22|"Everything is all right," Gehazi answered. "My master sent me to say, 'Two young men from the company of the prophets have just come to me from the hill country of Ephraim. Please give them a talent of silver and two sets of clothing.'"
2KGS|5|23|"By all means, take two talents," said Naaman. He urged Gehazi to accept them, and then tied up the two talents of silver in two bags, with two sets of clothing. He gave them to two of his servants, and they carried them ahead of Gehazi.
2KGS|5|24|When Gehazi came to the hill, he took the things from the servants and put them away in the house. He sent the men away and they left.
2KGS|5|25|Then he went in and stood before his master Elisha. "Where have you been, Gehazi?" Elisha asked. "Your servant didn't go anywhere," Gehazi answered.
2KGS|5|26|But Elisha said to him, "Was not my spirit with you when the man got down from his chariot to meet you? Is this the time to take money, or to accept clothes, olive groves, vineyards, flocks, herds, or menservants and maidservants?
2KGS|5|27|Naaman's leprosy will cling to you and to your descendants forever." Then Gehazi went from Elisha's presence and he was leprous, as white as snow.
2KGS|6|1|The company of the prophets said to Elisha, "Look, the place where we meet with you is too small for us.
2KGS|6|2|Let us go to the Jordan, where each of us can get a pole; and let us build a place there for us to live." And he said, "Go."
2KGS|6|3|Then one of them said, "Won't you please come with your servants?I will," Elisha replied.
2KGS|6|4|And he went with them. They went to the Jordan and began to cut down trees.
2KGS|6|5|As one of them was cutting down a tree, the iron axhead fell into the water. "Oh, my lord," he cried out, "it was borrowed!"
2KGS|6|6|The man of God asked, "Where did it fall?" When he showed him the place, Elisha cut a stick and threw it there, and made the iron float.
2KGS|6|7|"Lift it out," he said. Then the man reached out his hand and took it.
2KGS|6|8|Now the king of Aram was at war with Israel. After conferring with his officers, he said, "I will set up my camp in such and such a place."
2KGS|6|9|The man of God sent word to the king of Israel: "Beware of passing that place, because the Arameans are going down there."
2KGS|6|10|So the king of Israel checked on the place indicated by the man of God. Time and again Elisha warned the king, so that he was on his guard in such places.
2KGS|6|11|This enraged the king of Aram. He summoned his officers and demanded of them, "Will you not tell me which of us is on the side of the king of Israel?"
2KGS|6|12|"None of us, my lord the king," said one of his officers, "but Elisha, the prophet who is in Israel, tells the king of Israel the very words you speak in your bedroom."
2KGS|6|13|"Go, find out where he is," the king ordered, "so I can send men and capture him." The report came back: "He is in Dothan."
2KGS|6|14|Then he sent horses and chariots and a strong force there. They went by night and surrounded the city.
2KGS|6|15|When the servant of the man of God got up and went out early the next morning, an army with horses and chariots had surrounded the city. "Oh, my lord, what shall we do?" the servant asked.
2KGS|6|16|"Don't be afraid," the prophet answered. "Those who are with us are more than those who are with them."
2KGS|6|17|And Elisha prayed, "O LORD, open his eyes so he may see." Then the LORD opened the servant's eyes, and he looked and saw the hills full of horses and chariots of fire all around Elisha.
2KGS|6|18|As the enemy came down toward him, Elisha prayed to the LORD, "Strike these people with blindness." So he struck them with blindness, as Elisha had asked.
2KGS|6|19|Elisha told them, "This is not the road and this is not the city. Follow me, and I will lead you to the man you are looking for." And he led them to Samaria.
2KGS|6|20|After they entered the city, Elisha said, "LORD, open the eyes of these men so they can see." Then the LORD opened their eyes and they looked, and there they were, inside Samaria.
2KGS|6|21|When the king of Israel saw them, he asked Elisha, "Shall I kill them, my father? Shall I kill them?"
2KGS|6|22|"Do not kill them," he answered. "Would you kill men you have captured with your own sword or bow? Set food and water before them so that they may eat and drink and then go back to their master."
2KGS|6|23|So he prepared a great feast for them, and after they had finished eating and drinking, he sent them away, and they returned to their master. So the bands from Aram stopped raiding Israel's territory.
2KGS|6|24|Some time later, Ben-Hadad king of Aram mobilized his entire army and marched up and laid siege to Samaria.
2KGS|6|25|There was a great famine in the city; the siege lasted so long that a donkey's head sold for eighty shekels of silver, and a quarter of a cab of seed pods for five shekels.
2KGS|6|26|As the king of Israel was passing by on the wall, a woman cried to him, "Help me, my lord the king!"
2KGS|6|27|The king replied, "If the LORD does not help you, where can I get help for you? From the threshing floor? From the winepress?"
2KGS|6|28|Then he asked her, "What's the matter?" She answered, "This woman said to me, 'Give up your son so we may eat him today, and tomorrow we'll eat my son.'
2KGS|6|29|So we cooked my son and ate him. The next day I said to her, 'Give up your son so we may eat him,' but she had hidden him."
2KGS|6|30|When the king heard the woman's words, he tore his robes. As he went along the wall, the people looked, and there, underneath, he had sackcloth on his body.
2KGS|6|31|He said, "May God deal with me, be it ever so severely, if the head of Elisha son of Shaphat remains on his shoulders today!"
2KGS|6|32|Now Elisha was sitting in his house, and the elders were sitting with him. The king sent a messenger ahead, but before he arrived, Elisha said to the elders, "Don't you see how this murderer is sending someone to cut off my head? Look, when the messenger comes, shut the door and hold it shut against him. Is not the sound of his master's footsteps behind him?"
2KGS|6|33|While he was still talking to them, the messenger came down to him. And the king said, "This disaster is from the LORD. Why should I wait for the LORD any longer?"
2KGS|7|1|Elisha said, "Hear the word of the LORD. This is what the LORD says: About this time tomorrow, a seah of flour will sell for a shekel and two seahs of barley for a shekel at the gate of Samaria."
2KGS|7|2|The officer on whose arm the king was leaning said to the man of God, "Look, even if the LORD should open the floodgates of the heavens, could this happen?You will see it with your own eyes," answered Elisha, "but you will not eat any of it!"
2KGS|7|3|Now there were four men with leprosy at the entrance of the city gate. They said to each other, "Why stay here until we die?
2KGS|7|4|If we say, 'We'll go into the city'-the famine is there, and we will die. And if we stay here, we will die. So let's go over to the camp of the Arameans and surrender. If they spare us, we live; if they kill us, then we die."
2KGS|7|5|At dusk they got up and went to the camp of the Arameans. When they reached the edge of the camp, not a man was there,
2KGS|7|6|for the Lord had caused the Arameans to hear the sound of chariots and horses and a great army, so that they said to one another, "Look, the king of Israel has hired the Hittite and Egyptian kings to attack us!"
2KGS|7|7|So they got up and fled in the dusk and abandoned their tents and their horses and donkeys. They left the camp as it was and ran for their lives.
2KGS|7|8|The men who had leprosy reached the edge of the camp and entered one of the tents. They ate and drank, and carried away silver, gold and clothes, and went off and hid them. They returned and entered another tent and took some things from it and hid them also.
2KGS|7|9|Then they said to each other, "We're not doing right. This is a day of good news and we are keeping it to ourselves. If we wait until daylight, punishment will overtake us. Let's go at once and report this to the royal palace."
2KGS|7|10|So they went and called out to the city gatekeepers and told them, "We went into the Aramean camp and not a man was there-not a sound of anyone-only tethered horses and donkeys, and the tents left just as they were."
2KGS|7|11|The gatekeepers shouted the news, and it was reported within the palace.
2KGS|7|12|The king got up in the night and said to his officers, "I will tell you what the Arameans have done to us. They know we are starving; so they have left the camp to hide in the countryside, thinking, 'They will surely come out, and then we will take them alive and get into the city.'"
2KGS|7|13|One of his officers answered, "Have some men take five of the horses that are left in the city. Their plight will be like that of all the Israelites left here-yes, they will only be like all these Israelites who are doomed. So let us send them to find out what happened."
2KGS|7|14|So they selected two chariots with their horses, and the king sent them after the Aramean army. He commanded the drivers, "Go and find out what has happened."
2KGS|7|15|They followed them as far as the Jordan, and they found the whole road strewn with the clothing and equipment the Arameans had thrown away in their headlong flight. So the messengers returned and reported to the king.
2KGS|7|16|Then the people went out and plundered the camp of the Arameans. So a seah of flour sold for a shekel, and two seahs of barley sold for a shekel, as the LORD had said.
2KGS|7|17|Now the king had put the officer on whose arm he leaned in charge of the gate, and the people trampled him in the gateway, and he died, just as the man of God had foretold when the king came down to his house.
2KGS|7|18|It happened as the man of God had said to the king: "About this time tomorrow, a seah of flour will sell for a shekel and two seahs of barley for a shekel at the gate of Samaria."
2KGS|7|19|The officer had said to the man of God, "Look, even if the LORD should open the floodgates of the heavens, could this happen?" The man of God had replied, "You will see it with your own eyes, but you will not eat any of it!"
2KGS|7|20|And that is exactly what happened to him, for the people trampled him in the gateway, and he died.
2KGS|8|1|Now Elisha had said to the woman whose son he had restored to life, "Go away with your family and stay for a while wherever you can, because the LORD has decreed a famine in the land that will last seven years."
2KGS|8|2|The woman proceeded to do as the man of God said. She and her family went away and stayed in the land of the Philistines seven years.
2KGS|8|3|At the end of the seven years she came back from the land of the Philistines and went to the king to beg for her house and land.
2KGS|8|4|The king was talking to Gehazi, the servant of the man of God, and had said, "Tell me about all the great things Elisha has done."
2KGS|8|5|Just as Gehazi was telling the king how Elisha had restored the dead to life, the woman whose son Elisha had brought back to life came to beg the king for her house and land. Gehazi said, "This is the woman, my lord the king, and this is her son whom Elisha restored to life."
2KGS|8|6|The king asked the woman about it, and she told him. Then he assigned an official to her case and said to him, "Give back everything that belonged to her, including all the income from her land from the day she left the country until now."
2KGS|8|7|Elisha went to Damascus, and Ben-Hadad king of Aram was ill. When the king was told, "The man of God has come all the way up here,"
2KGS|8|8|he said to Hazael, "Take a gift with you and go to meet the man of God. Consult the LORD through him; ask him, 'Will I recover from this illness?'"
2KGS|8|9|Hazael went to meet Elisha, taking with him as a gift forty camel-loads of all the finest wares of Damascus. He went in and stood before him, and said, "Your son Ben-Hadad king of Aram has sent me to ask, 'Will I recover from this illness?'"
2KGS|8|10|Elisha answered, "Go and say to him, 'You will certainly recover'; but the LORD has revealed to me that he will in fact die."
2KGS|8|11|He stared at him with a fixed gaze until Hazael felt ashamed. Then the man of God began to weep.
2KGS|8|12|"Why is my lord weeping?" asked Hazael. "Because I know the harm you will do to the Israelites," he answered. "You will set fire to their fortified places, kill their young men with the sword, dash their little children to the ground, and rip open their pregnant women."
2KGS|8|13|Hazael said, "How could your servant, a mere dog, accomplish such a feat?The LORD has shown me that you will become king of Aram," answered Elisha.
2KGS|8|14|Then Hazael left Elisha and returned to his master. When Ben-Hadad asked, "What did Elisha say to you?" Hazael replied, "He told me that you would certainly recover."
2KGS|8|15|But the next day he took a thick cloth, soaked it in water and spread it over the king's face, so that he died. Then Hazael succeeded him as king.
2KGS|8|16|In the fifth year of Joram son of Ahab king of Israel, when Jehoshaphat was king of Judah, Jehoram son of Jehoshaphat began his reign as king of Judah.
2KGS|8|17|He was thirty-two years old when he became king, and he reigned in Jerusalem eight years.
2KGS|8|18|He walked in the ways of the kings of Israel, as the house of Ahab had done, for he married a daughter of Ahab. He did evil in the eyes of the LORD.
2KGS|8|19|Nevertheless, for the sake of his servant David, the LORD was not willing to destroy Judah. He had promised to maintain a lamp for David and his descendants forever.
2KGS|8|20|In the time of Jehoram, Edom rebelled against Judah and set up its own king.
2KGS|8|21|So Jehoram went to Zair with all his chariots. The Edomites surrounded him and his chariot commanders, but he rose up and broke through by night; his army, however, fled back home.
2KGS|8|22|To this day Edom has been in rebellion against Judah. Libnah revolted at the same time.
2KGS|8|23|As for the other events of Jehoram's reign, and all he did, are they not written in the book of the annals of the kings of Judah?
2KGS|8|24|Jehoram rested with his fathers and was buried with them in the City of David. And Ahaziah his son succeeded him as king.
2KGS|8|25|In the twelfth year of Joram son of Ahab king of Israel, Ahaziah son of Jehoram king of Judah began to reign.
2KGS|8|26|Ahaziah was twenty-two years old when he became king, and he reigned in Jerusalem one year. His mother's name was Athaliah, a granddaughter of Omri king of Israel.
2KGS|8|27|He walked in the ways of the house of Ahab and did evil in the eyes of the LORD, as the house of Ahab had done, for he was related by marriage to Ahab's family.
2KGS|8|28|Ahaziah went with Joram son of Ahab to war against Hazael king of Aram at Ramoth Gilead. The Arameans wounded Joram;
2KGS|8|29|so King Joram returned to Jezreel to recover from the wounds the Arameans had inflicted on him at Ramoth in his battle with Hazael king of Aram. Then Ahaziah son of Jehoram king of Judah went down to Jezreel to see Joram son of Ahab, because he had been wounded.
2KGS|9|1|The prophet Elisha summoned a man from the company of the prophets and said to him, "Tuck your cloak into your belt, take this flask of oil with you and go to Ramoth Gilead.
2KGS|9|2|When you get there, look for Jehu son of Jehoshaphat, the son of Nimshi. Go to him, get him away from his companions and take him into an inner room.
2KGS|9|3|Then take the flask and pour the oil on his head and declare, 'This is what the LORD says: I anoint you king over Israel.' Then open the door and run; don't delay!"
2KGS|9|4|So the young man, the prophet, went to Ramoth Gilead.
2KGS|9|5|When he arrived, he found the army officers sitting together. "I have a message for you, commander," he said. "For which of us?" asked Jehu. "For you, commander," he replied.
2KGS|9|6|Jehu got up and went into the house. Then the prophet poured the oil on Jehu's head and declared, "This is what the LORD, the God of Israel, says: 'I anoint you king over the LORD's people Israel.
2KGS|9|7|You are to destroy the house of Ahab your master, and I will avenge the blood of my servants the prophets and the blood of all the LORD's servants shed by Jezebel.
2KGS|9|8|The whole house of Ahab will perish. I will cut off from Ahab every last male in Israel-slave or free.
2KGS|9|9|I will make the house of Ahab like the house of Jeroboam son of Nebat and like the house of Baasha son of Ahijah.
2KGS|9|10|As for Jezebel, dogs will devour her on the plot of ground at Jezreel, and no one will bury her.'" Then he opened the door and ran.
2KGS|9|11|When Jehu went out to his fellow officers, one of them asked him, "Is everything all right? Why did this madman come to you?You know the man and the sort of things he says," Jehu replied.
2KGS|9|12|"That's not true!" they said. "Tell us." Jehu said, "Here is what he told me: 'This is what the LORD says: I anoint you king over Israel.'"
2KGS|9|13|They hurried and took their cloaks and spread them under him on the bare steps. Then they blew the trumpet and shouted, "Jehu is king!"
2KGS|9|14|So Jehu son of Jehoshaphat, the son of Nimshi, conspired against Joram. (Now Joram and all Israel had been defending Ramoth Gilead against Hazael king of Aram,
2KGS|9|15|but King Joram had returned to Jezreel to recover from the wounds the Arameans had inflicted on him in the battle with Hazael king of Aram.) Jehu said, "If this is the way you feel, don't let anyone slip out of the city to go and tell the news in Jezreel."
2KGS|9|16|Then he got into his chariot and rode to Jezreel, because Joram was resting there and Ahaziah king of Judah had gone down to see him.
2KGS|9|17|When the lookout standing on the tower in Jezreel saw Jehu's troops approaching, he called out, "I see some troops coming.Get a horseman," Joram ordered. "Send him to meet them and ask, 'Do you come in peace?'"
2KGS|9|18|The horseman rode off to meet Jehu and said, "This is what the king says: 'Do you come in peace?' What do you have to do with peace?" Jehu replied. "Fall in behind me." The lookout reported, "The messenger has reached them, but he isn't coming back."
2KGS|9|19|So the king sent out a second horseman. When he came to them he said, "This is what the king says: 'Do you come in peace?'" Jehu replied, "What do you have to do with peace? Fall in behind me."
2KGS|9|20|The lookout reported, "He has reached them, but he isn't coming back either. The driving is like that of Jehu son of Nimshi-he drives like a madman."
2KGS|9|21|"Hitch up my chariot," Joram ordered. And when it was hitched up, Joram king of Israel and Ahaziah king of Judah rode out, each in his own chariot, to meet Jehu. They met him at the plot of ground that had belonged to Naboth the Jezreelite.
2KGS|9|22|When Joram saw Jehu he asked, "Have you come in peace, Jehu?How can there be peace," Jehu replied, "as long as all the idolatry and witchcraft of your mother Jezebel abound?"
2KGS|9|23|Joram turned about and fled, calling out to Ahaziah, "Treachery, Ahaziah!"
2KGS|9|24|Then Jehu drew his bow and shot Joram between the shoulders. The arrow pierced his heart and he slumped down in his chariot.
2KGS|9|25|Jehu said to Bidkar, his chariot officer, "Pick him up and throw him on the field that belonged to Naboth the Jezreelite. Remember how you and I were riding together in chariots behind Ahab his father when the LORD made this prophecy about him:
2KGS|9|26|'Yesterday I saw the blood of Naboth and the blood of his sons, declares the LORD, and I will surely make you pay for it on this plot of ground, declares the LORD.' Now then, pick him up and throw him on that plot, in accordance with the word of the LORD."
2KGS|9|27|When Ahaziah king of Judah saw what had happened, he fled up the road to Beth Haggan. Jehu chased him, shouting, "Kill him too!" They wounded him in his chariot on the way up to Gur near Ibleam, but he escaped to Megiddo and died there.
2KGS|9|28|His servants took him by chariot to Jerusalem and buried him with his fathers in his tomb in the City of David.
2KGS|9|29|(In the eleventh year of Joram son of Ahab, Ahaziah had become king of Judah.)
2KGS|9|30|Then Jehu went to Jezreel. When Jezebel heard about it, she painted her eyes, arranged her hair and looked out of a window.
2KGS|9|31|As Jehu entered the gate, she asked, "Have you come in peace, Zimri, you murderer of your master?"
2KGS|9|32|He looked up at the window and called out, "Who is on my side? Who?" Two or three eunuchs looked down at him.
2KGS|9|33|"Throw her down!" Jehu said. So they threw her down, and some of her blood spattered the wall and the horses as they trampled her underfoot.
2KGS|9|34|Jehu went in and ate and drank. "Take care of that cursed woman," he said, "and bury her, for she was a king's daughter."
2KGS|9|35|But when they went out to bury her, they found nothing except her skull, her feet and her hands.
2KGS|9|36|They went back and told Jehu, who said, "This is the word of the LORD that he spoke through his servant Elijah the Tishbite: On the plot of ground at Jezreel dogs will devour Jezebel's flesh.
2KGS|9|37|Jezebel's body will be like refuse on the ground in the plot at Jezreel, so that no one will be able to say, 'This is Jezebel.'"
2KGS|10|1|Now there were in Samaria seventy sons of the house of Ahab. So Jehu wrote letters and sent them to Samaria: to the officials of Jezreel, to the elders and to the guardians of Ahab's children. He said,
2KGS|10|2|"As soon as this letter reaches you, since your master's sons are with you and you have chariots and horses, a fortified city and weapons,
2KGS|10|3|choose the best and most worthy of your master's sons and set him on his father's throne. Then fight for your master's house."
2KGS|10|4|But they were terrified and said, "If two kings could not resist him, how can we?"
2KGS|10|5|So the palace administrator, the city governor, the elders and the guardians sent this message to Jehu: "We are your servants and we will do anything you say. We will not appoint anyone as king; you do whatever you think best."
2KGS|10|6|Then Jehu wrote them a second letter, saying, "If you are on my side and will obey me, take the heads of your master's sons and come to me in Jezreel by this time tomorrow." Now the royal princes, seventy of them, were with the leading men of the city, who were rearing them.
2KGS|10|7|When the letter arrived, these men took the princes and slaughtered all seventy of them. They put their heads in baskets and sent them to Jehu in Jezreel.
2KGS|10|8|When the messenger arrived, he told Jehu, "They have brought the heads of the princes." Then Jehu ordered, "Put them in two piles at the entrance of the city gate until morning."
2KGS|10|9|The next morning Jehu went out. He stood before all the people and said, "You are innocent. It was I who conspired against my master and killed him, but who killed all these?
2KGS|10|10|Know then, that not a word the LORD has spoken against the house of Ahab will fail. The LORD has done what he promised through his servant Elijah."
2KGS|10|11|So Jehu killed everyone in Jezreel who remained of the house of Ahab, as well as all his chief men, his close friends and his priests, leaving him no survivor.
2KGS|10|12|Jehu then set out and went toward Samaria. At Beth Eked of the Shepherds,
2KGS|10|13|he met some relatives of Ahaziah king of Judah and asked, "Who are you?" They said, "We are relatives of Ahaziah, and we have come down to greet the families of the king and of the queen mother."
2KGS|10|14|"Take them alive!" he ordered. So they took them alive and slaughtered them by the well of Beth Eked-forty-two men. He left no survivor.
2KGS|10|15|After he left there, he came upon Jehonadab son of Recab, who was on his way to meet him. Jehu greeted him and said, "Are you in accord with me, as I am with you?I am," Jehonadab answered. "If so," said Jehu, "give me your hand." So he did, and Jehu helped him up into the chariot.
2KGS|10|16|Jehu said, "Come with me and see my zeal for the LORD." Then he had him ride along in his chariot.
2KGS|10|17|When Jehu came to Samaria, he killed all who were left there of Ahab's family; he destroyed them, according to the word of the LORD spoken to Elijah.
2KGS|10|18|Then Jehu brought all the people together and said to them, "Ahab served Baal a little; Jehu will serve him much.
2KGS|10|19|Now summon all the prophets of Baal, all his ministers and all his priests. See that no one is missing, because I am going to hold a great sacrifice for Baal. Anyone who fails to come will no longer live." But Jehu was acting deceptively in order to destroy the ministers of Baal.
2KGS|10|20|Jehu said, "Call an assembly in honor of Baal." So they proclaimed it.
2KGS|10|21|Then he sent word throughout Israel, and all the ministers of Baal came; not one stayed away. They crowded into the temple of Baal until it was full from one end to the other.
2KGS|10|22|And Jehu said to the keeper of the wardrobe, "Bring robes for all the ministers of Baal." So he brought out robes for them.
2KGS|10|23|Then Jehu and Jehonadab son of Recab went into the temple of Baal. Jehu said to the ministers of Baal, "Look around and see that no servants of the LORD are here with you-only ministers of Baal."
2KGS|10|24|So they went in to make sacrifices and burnt offerings. Now Jehu had posted eighty men outside with this warning: "If one of you lets any of the men I am placing in your hands escape, it will be your life for his life."
2KGS|10|25|As soon as Jehu had finished making the burnt offering, he ordered the guards and officers: "Go in and kill them; let no one escape." So they cut them down with the sword. The guards and officers threw the bodies out and then entered the inner shrine of the temple of Baal.
2KGS|10|26|They brought the sacred stone out of the temple of Baal and burned it.
2KGS|10|27|They demolished the sacred stone of Baal and tore down the temple of Baal, and people have used it for a latrine to this day.
2KGS|10|28|So Jehu destroyed Baal worship in Israel.
2KGS|10|29|However, he did not turn away from the sins of Jeroboam son of Nebat, which he had caused Israel to commit-the worship of the golden calves at Bethel and Dan.
2KGS|10|30|The LORD said to Jehu, "Because you have done well in accomplishing what is right in my eyes and have done to the house of Ahab all I had in mind to do, your descendants will sit on the throne of Israel to the fourth generation."
2KGS|10|31|Yet Jehu was not careful to keep the law of the LORD, the God of Israel, with all his heart. He did not turn away from the sins of Jeroboam, which he had caused Israel to commit.
2KGS|10|32|In those days the LORD began to reduce the size of Israel. Hazael overpowered the Israelites throughout their territory
2KGS|10|33|east of the Jordan in all the land of Gilead (the region of Gad, Reuben and Manasseh), from Aroer by the Arnon Gorge through Gilead to Bashan.
2KGS|10|34|As for the other events of Jehu's reign, all he did, and all his achievements, are they not written in the book of the annals of the kings of Israel?
2KGS|10|35|Jehu rested with his fathers and was buried in Samaria. And Jehoahaz his son succeeded him as king.
2KGS|10|36|The time that Jehu reigned over Israel in Samaria was twenty-eight years.
2KGS|11|1|When Athaliah the mother of Ahaziah saw that her son was dead, she proceeded to destroy the whole royal family.
2KGS|11|2|But Jehosheba, the daughter of King Jehoram and sister of Ahaziah, took Joash son of Ahaziah and stole him away from among the royal princes, who were about to be murdered. She put him and his nurse in a bedroom to hide him from Athaliah; so he was not killed.
2KGS|11|3|He remained hidden with his nurse at the temple of the LORD for six years while Athaliah ruled the land.
2KGS|11|4|In the seventh year Jehoiada sent for the commanders of units of a hundred, the Carites and the guards and had them brought to him at the temple of the LORD. He made a covenant with them and put them under oath at the temple of the LORD. Then he showed them the king's son.
2KGS|11|5|He commanded them, saying, "This is what you are to do: You who are in the three companies that are going on duty on the Sabbath-a third of you guarding the royal palace,
2KGS|11|6|a third at the Sur Gate, and a third at the gate behind the guard, who take turns guarding the temple-
2KGS|11|7|and you who are in the other two companies that normally go off Sabbath duty are all to guard the temple for the king.
2KGS|11|8|Station yourselves around the king, each man with his weapon in his hand. Anyone who approaches your ranks must be put to death. Stay close to the king wherever he goes."
2KGS|11|9|The commanders of units of a hundred did just as Jehoiada the priest ordered. Each one took his men-those who were going on duty on the Sabbath and those who were going off duty-and came to Jehoiada the priest.
2KGS|11|10|Then he gave the commanders the spears and shields that had belonged to King David and that were in the temple of the LORD.
2KGS|11|11|The guards, each with his weapon in his hand, stationed themselves around the king-near the altar and the temple, from the south side to the north side of the temple.
2KGS|11|12|Jehoiada brought out the king's son and put the crown on him; he presented him with a copy of the covenant and proclaimed him king. They anointed him, and the people clapped their hands and shouted, "Long live the king!"
2KGS|11|13|When Athaliah heard the noise made by the guards and the people, she went to the people at the temple of the LORD.
2KGS|11|14|She looked and there was the king, standing by the pillar, as the custom was. The officers and the trumpeters were beside the king, and all the people of the land were rejoicing and blowing trumpets. Then Athaliah tore her robes and called out, "Treason! Treason!"
2KGS|11|15|Jehoiada the priest ordered the commanders of units of a hundred, who were in charge of the troops: "Bring her out between the ranks and put to the sword anyone who follows her." For the priest had said, "She must not be put to death in the temple of the LORD."
2KGS|11|16|So they seized her as she reached the place where the horses enter the palace grounds, and there she was put to death.
2KGS|11|17|Jehoiada then made a covenant between the LORD and the king and people that they would be the LORD's people. He also made a covenant between the king and the people.
2KGS|11|18|All the people of the land went to the temple of Baal and tore it down. They smashed the altars and idols to pieces and killed Mattan the priest of Baal in front of the altars. Then Jehoiada the priest posted guards at the temple of the LORD.
2KGS|11|19|He took with him the commanders of hundreds, the Carites, the guards and all the people of the land, and together they brought the king down from the temple of the LORD and went into the palace, entering by way of the gate of the guards. The king then took his place on the royal throne,
2KGS|11|20|and all the people of the land rejoiced. And the city was quiet, because Athaliah had been slain with the sword at the palace.
2KGS|11|21|Joash was seven years old when he began to reign.
2KGS|12|1|In the seventh year of Jehu, Joash became king, and he reigned in Jerusalem forty years. His mother's name was Zibiah; she was from Beersheba.
2KGS|12|2|Joash did what was right in the eyes of the LORD all the years Jehoiada the priest instructed him.
2KGS|12|3|The high places, however, were not removed; the people continued to offer sacrifices and burn incense there.
2KGS|12|4|Joash said to the priests, "Collect all the money that is brought as sacred offerings to the temple of the LORD -the money collected in the census, the money received from personal vows and the money brought voluntarily to the temple.
2KGS|12|5|Let every priest receive the money from one of the treasurers, and let it be used to repair whatever damage is found in the temple."
2KGS|12|6|But by the twenty-third year of King Joash the priests still had not repaired the temple.
2KGS|12|7|Therefore King Joash summoned Jehoiada the priest and the other priests and asked them, "Why aren't you repairing the damage done to the temple? Take no more money from your treasurers, but hand it over for repairing the temple."
2KGS|12|8|The priests agreed that they would not collect any more money from the people and that they would not repair the temple themselves.
2KGS|12|9|Jehoiada the priest took a chest and bored a hole in its lid. He placed it beside the altar, on the right side as one enters the temple of the LORD. The priests who guarded the entrance put into the chest all the money that was brought to the temple of the LORD.
2KGS|12|10|Whenever they saw that there was a large amount of money in the chest, the royal secretary and the high priest came, counted the money that had been brought into the temple of the LORD and put it into bags.
2KGS|12|11|When the amount had been determined, they gave the money to the men appointed to supervise the work on the temple. With it they paid those who worked on the temple of the LORD -the carpenters and builders,
2KGS|12|12|the masons and stonecutters. They purchased timber and dressed stone for the repair of the temple of the LORD, and met all the other expenses of restoring the temple.
2KGS|12|13|The money brought into the temple was not spent for making silver basins, wick trimmers, sprinkling bowls, trumpets or any other articles of gold or silver for the temple of the LORD;
2KGS|12|14|it was paid to the workmen, who used it to repair the temple.
2KGS|12|15|They did not require an accounting from those to whom they gave the money to pay the workers, because they acted with complete honesty.
2KGS|12|16|The money from the guilt offerings and sin offerings was not brought into the temple of the LORD; it belonged to the priests.
2KGS|12|17|About this time Hazael king of Aram went up and attacked Gath and captured it. Then he turned to attack Jerusalem.
2KGS|12|18|But Joash king of Judah took all the sacred objects dedicated by his fathers-Jehoshaphat, Jehoram and Ahaziah, the kings of Judah-and the gifts he himself had dedicated and all the gold found in the treasuries of the temple of the LORD and of the royal palace, and he sent them to Hazael king of Aram, who then withdrew from Jerusalem.
2KGS|12|19|As for the other events of the reign of Joash, and all he did, are they not written in the book of the annals of the kings of Judah?
2KGS|12|20|His officials conspired against him and assassinated him at Beth Millo, on the road down to Silla.
2KGS|12|21|The officials who murdered him were Jozabad son of Shimeath and Jehozabad son of Shomer. He died and was buried with his fathers in the City of David. And Amaziah his son succeeded him as king.
2KGS|13|1|In the twenty-third year of Joash son of Ahaziah king of Judah, Jehoahaz son of Jehu became king of Israel in Samaria, and he reigned seventeen years.
2KGS|13|2|He did evil in the eyes of the LORD by following the sins of Jeroboam son of Nebat, which he had caused Israel to commit, and he did not turn away from them.
2KGS|13|3|So the LORD's anger burned against Israel, and for a long time he kept them under the power of Hazael king of Aram and Ben-Hadad his son.
2KGS|13|4|Then Jehoahaz sought the LORD's favor, and the LORD listened to him, for he saw how severely the king of Aram was oppressing Israel.
2KGS|13|5|The LORD provided a deliverer for Israel, and they escaped from the power of Aram. So the Israelites lived in their own homes as they had before.
2KGS|13|6|But they did not turn away from the sins of the house of Jeroboam, which he had caused Israel to commit; they continued in them. Also, the Asherah pole remained standing in Samaria.
2KGS|13|7|Nothing had been left of the army of Jehoahaz except fifty horsemen, ten chariots and ten thousand foot soldiers, for the king of Aram had destroyed the rest and made them like the dust at threshing time.
2KGS|13|8|As for the other events of the reign of Jehoahaz, all he did and his achievements, are they not written in the book of the annals of the kings of Israel?
2KGS|13|9|Jehoahaz rested with his fathers and was buried in Samaria. And Jehoash his son succeeded him as king.
2KGS|13|10|In the thirty-seventh year of Joash king of Judah, Jehoash son of Jehoahaz became king of Israel in Samaria, and he reigned sixteen years.
2KGS|13|11|He did evil in the eyes of the LORD and did not turn away from any of the sins of Jeroboam son of Nebat, which he had caused Israel to commit; he continued in them.
2KGS|13|12|As for the other events of the reign of Jehoash, all he did and his achievements, including his war against Amaziah king of Judah, are they not written in the book of the annals of the kings of Israel?
2KGS|13|13|Jehoash rested with his fathers, and Jeroboam succeeded him on the throne. Jehoash was buried in Samaria with the kings of Israel.
2KGS|13|14|Now Elisha was suffering from the illness from which he died. Jehoash king of Israel went down to see him and wept over him. "My father! My father!" he cried. "The chariots and horsemen of Israel!"
2KGS|13|15|Elisha said, "Get a bow and some arrows," and he did so.
2KGS|13|16|"Take the bow in your hands," he said to the king of Israel. When he had taken it, Elisha put his hands on the king's hands.
2KGS|13|17|"Open the east window," he said, and he opened it. "Shoot!" Elisha said, and he shot. "The LORD's arrow of victory, the arrow of victory over Aram!" Elisha declared. "You will completely destroy the Arameans at Aphek."
2KGS|13|18|Then he said, "Take the arrows," and the king took them. Elisha told him, "Strike the ground." He struck it three times and stopped.
2KGS|13|19|The man of God was angry with him and said, "You should have struck the ground five or six times; then you would have defeated Aram and completely destroyed it. But now you will defeat it only three times."
2KGS|13|20|Elisha died and was buried. Now Moabite raiders used to enter the country every spring.
2KGS|13|21|Once while some Israelites were burying a man, suddenly they saw a band of raiders; so they threw the man's body into Elisha's tomb. When the body touched Elisha's bones, the man came to life and stood up on his feet.
2KGS|13|22|Hazael king of Aram oppressed Israel throughout the reign of Jehoahaz.
2KGS|13|23|But the LORD was gracious to them and had compassion and showed concern for them because of his covenant with Abraham, Isaac and Jacob. To this day he has been unwilling to destroy them or banish them from his presence.
2KGS|13|24|Hazael king of Aram died, and Ben-Hadad his son succeeded him as king.
2KGS|13|25|Then Jehoash son of Jehoahaz recaptured from Ben-Hadad son of Hazael the towns he had taken in battle from his father Jehoahaz. Three times Jehoash defeated him, and so he recovered the Israelite towns.
2KGS|14|1|In the second year of Jehoash son of Jehoahaz king of Israel, Amaziah son of Joash king of Judah began to reign.
2KGS|14|2|He was twenty-five years old when he became king, and he reigned in Jerusalem twenty-nine years. His mother's name was Jehoaddin; she was from Jerusalem.
2KGS|14|3|He did what was right in the eyes of the LORD, but not as his father David had done. In everything he followed the example of his father Joash.
2KGS|14|4|The high places, however, were not removed; the people continued to offer sacrifices and burn incense there.
2KGS|14|5|After the kingdom was firmly in his grasp, he executed the officials who had murdered his father the king.
2KGS|14|6|Yet he did not put the sons of the assassins to death, in accordance with what is written in the Book of the Law of Moses where the LORD commanded: "Fathers shall not be put to death for their children, nor children put to death for their fathers; each is to die for his own sins."
2KGS|14|7|He was the one who defeated ten thousand Edomites in the Valley of Salt and captured Sela in battle, calling it Joktheel, the name it has to this day.
2KGS|14|8|Then Amaziah sent messengers to Jehoash son of Jehoahaz, the son of Jehu, king of Israel, with the challenge: "Come, meet me face to face."
2KGS|14|9|But Jehoash king of Israel replied to Amaziah king of Judah: "A thistle in Lebanon sent a message to a cedar in Lebanon, 'Give your daughter to my son in marriage.' Then a wild beast in Lebanon came along and trampled the thistle underfoot.
2KGS|14|10|You have indeed defeated Edom and now you are arrogant. Glory in your victory, but stay at home! Why ask for trouble and cause your own downfall and that of Judah also?"
2KGS|14|11|Amaziah, however, would not listen, so Jehoash king of Israel attacked. He and Amaziah king of Judah faced each other at Beth Shemesh in Judah.
2KGS|14|12|Judah was routed by Israel, and every man fled to his home.
2KGS|14|13|Jehoash king of Israel captured Amaziah king of Judah, the son of Joash, the son of Ahaziah, at Beth Shemesh. Then Jehoash went to Jerusalem and broke down the wall of Jerusalem from the Ephraim Gate to the Corner Gate-a section about six hundred feet long.
2KGS|14|14|He took all the gold and silver and all the articles found in the temple of the LORD and in the treasuries of the royal palace. He also took hostages and returned to Samaria.
2KGS|14|15|As for the other events of the reign of Jehoash, what he did and his achievements, including his war against Amaziah king of Judah, are they not written in the book of the annals of the kings of Israel?
2KGS|14|16|Jehoash rested with his fathers and was buried in Samaria with the kings of Israel. And Jeroboam his son succeeded him as king.
2KGS|14|17|Amaziah son of Joash king of Judah lived for fifteen years after the death of Jehoash son of Jehoahaz king of Israel.
2KGS|14|18|As for the other events of Amaziah's reign, are they not written in the book of the annals of the kings of Judah?
2KGS|14|19|They conspired against him in Jerusalem, and he fled to Lachish, but they sent men after him to Lachish and killed him there.
2KGS|14|20|He was brought back by horse and was buried in Jerusalem with his fathers, in the City of David.
2KGS|14|21|Then all the people of Judah took Azariah, who was sixteen years old, and made him king in place of his father Amaziah.
2KGS|14|22|He was the one who rebuilt Elath and restored it to Judah after Amaziah rested with his fathers.
2KGS|14|23|In the fifteenth year of Amaziah son of Joash king of Judah, Jeroboam son of Jehoash king of Israel became king in Samaria, and he reigned forty-one years.
2KGS|14|24|He did evil in the eyes of the LORD and did not turn away from any of the sins of Jeroboam son of Nebat, which he had caused Israel to commit.
2KGS|14|25|He was the one who restored the boundaries of Israel from Lebo Hamath to the Sea of the Arabah, in accordance with the word of the LORD, the God of Israel, spoken through his servant Jonah son of Amittai, the prophet from Gath Hepher.
2KGS|14|26|The LORD had seen how bitterly everyone in Israel, whether slave or free, was suffering; there was no one to help them.
2KGS|14|27|And since the LORD had not said he would blot out the name of Israel from under heaven, he saved them by the hand of Jeroboam son of Jehoash.
2KGS|14|28|As for the other events of Jeroboam's reign, all he did, and his military achievements, including how he recovered for Israel both Damascus and Hamath, which had belonged to Yaudi, are they not written in the book of the annals of the kings of Israel?
2KGS|14|29|Jeroboam rested with his fathers, the kings of Israel. And Zechariah his son succeeded him as king.
2KGS|15|1|In the twenty-seventh year of Jeroboam king of Israel, Azariah son of Amaziah king of Judah began to reign.
2KGS|15|2|He was sixteen years old when he became king, and he reigned in Jerusalem fifty-two years. His mother's name was Jecoliah; she was from Jerusalem.
2KGS|15|3|He did what was right in the eyes of the LORD, just as his father Amaziah had done.
2KGS|15|4|The high places, however, were not removed; the people continued to offer sacrifices and burn incense there.
2KGS|15|5|The LORD afflicted the king with leprosy until the day he died, and he lived in a separate house. Jotham the king's son had charge of the palace and governed the people of the land.
2KGS|15|6|As for the other events of Azariah's reign, and all he did, are they not written in the book of the annals of the kings of Judah?
2KGS|15|7|Azariah rested with his fathers and was buried near them in the City of David. And Jotham his son succeeded him as king.
2KGS|15|8|In the thirty-eighth year of Azariah king of Judah, Zechariah son of Jeroboam became king of Israel in Samaria, and he reigned six months.
2KGS|15|9|He did evil in the eyes of the LORD, as his fathers had done. He did not turn away from the sins of Jeroboam son of Nebat, which he had caused Israel to commit.
2KGS|15|10|Shallum son of Jabesh conspired against Zechariah. He attacked him in front of the people, assassinated him and succeeded him as king.
2KGS|15|11|The other events of Zechariah's reign are written in the book of the annals of the kings of Israel.
2KGS|15|12|So the word of the LORD spoken to Jehu was fulfilled: "Your descendants will sit on the throne of Israel to the fourth generation."
2KGS|15|13|Shallum son of Jabesh became king in the thirty-ninth year of Uzziah king of Judah, and he reigned in Samaria one month.
2KGS|15|14|Then Menahem son of Gadi went from Tirzah up to Samaria. He attacked Shallum son of Jabesh in Samaria, assassinated him and succeeded him as king.
2KGS|15|15|The other events of Shallum's reign, and the conspiracy he led, are written in the book of the annals of the kings of Israel.
2KGS|15|16|At that time Menahem, starting out from Tirzah, attacked Tiphsah and everyone in the city and its vicinity, because they refused to open their gates. He sacked Tiphsah and ripped open all the pregnant women.
2KGS|15|17|In the thirty-ninth year of Azariah king of Judah, Menahem son of Gadi became king of Israel, and he reigned in Samaria ten years.
2KGS|15|18|He did evil in the eyes of the LORD. During his entire reign he did not turn away from the sins of Jeroboam son of Nebat, which he had caused Israel to commit.
2KGS|15|19|Then Pul king of Assyria invaded the land, and Menahem gave him a thousand talents of silver to gain his support and strengthen his own hold on the kingdom.
2KGS|15|20|Menahem exacted this money from Israel. Every wealthy man had to contribute fifty shekels of silver to be given to the king of Assyria. So the king of Assyria withdrew and stayed in the land no longer.
2KGS|15|21|As for the other events of Menahem's reign, and all he did, are they not written in the book of the annals of the kings of Israel?
2KGS|15|22|Menahem rested with his fathers. And Pekahiah his son succeeded him as king.
2KGS|15|23|In the fiftieth year of Azariah king of Judah, Pekahiah son of Menahem became king of Israel in Samaria, and he reigned two years.
2KGS|15|24|Pekahiah did evil in the eyes of the LORD. He did not turn away from the sins of Jeroboam son of Nebat, which he had caused Israel to commit.
2KGS|15|25|One of his chief officers, Pekah son of Remaliah, conspired against him. Taking fifty men of Gilead with him, he assassinated Pekahiah, along with Argob and Arieh, in the citadel of the royal palace at Samaria. So Pekah killed Pekahiah and succeeded him as king.
2KGS|15|26|The other events of Pekahiah's reign, and all he did, are written in the book of the annals of the kings of Israel.
2KGS|15|27|In the fifty-second year of Azariah king of Judah, Pekah son of Remaliah became king of Israel in Samaria, and he reigned twenty years.
2KGS|15|28|He did evil in the eyes of the LORD. He did not turn away from the sins of Jeroboam son of Nebat, which he had caused Israel to commit.
2KGS|15|29|In the time of Pekah king of Israel, Tiglath-Pileser king of Assyria came and took Ijon, Abel Beth Maacah, Janoah, Kedesh and Hazor. He took Gilead and Galilee, including all the land of Naphtali, and deported the people to Assyria.
2KGS|15|30|Then Hoshea son of Elah conspired against Pekah son of Remaliah. He attacked and assassinated him, and then succeeded him as king in the twentieth year of Jotham son of Uzziah.
2KGS|15|31|As for the other events of Pekah's reign, and all he did, are they not written in the book of the annals of the kings of Israel?
2KGS|15|32|In the second year of Pekah son of Remaliah king of Israel, Jotham son of Uzziah king of Judah began to reign.
2KGS|15|33|He was twenty-five years old when he became king, and he reigned in Jerusalem sixteen years. His mother's name was Jerusha daughter of Zadok.
2KGS|15|34|He did what was right in the eyes of the LORD, just as his father Uzziah had done.
2KGS|15|35|The high places, however, were not removed; the people continued to offer sacrifices and burn incense there. Jotham rebuilt the Upper Gate of the temple of the LORD.
2KGS|15|36|As for the other events of Jotham's reign, and what he did, are they not written in the book of the annals of the kings of Judah?
2KGS|15|37|(In those days the LORD began to send Rezin king of Aram and Pekah son of Remaliah against Judah.)
2KGS|15|38|Jotham rested with his fathers and was buried with them in the City of David, the city of his father. And Ahaz his son succeeded him as king.
2KGS|16|1|In the seventeenth year of Pekah son of Remaliah, Ahaz son of Jotham king of Judah began to reign.
2KGS|16|2|Ahaz was twenty years old when he became king, and he reigned in Jerusalem sixteen years. Unlike David his father, he did not do what was right in the eyes of the LORD his God.
2KGS|16|3|He walked in the ways of the kings of Israel and even sacrificed his son in the fire, following the detestable ways of the nations the LORD had driven out before the Israelites.
2KGS|16|4|He offered sacrifices and burned incense at the high places, on the hilltops and under every spreading tree.
2KGS|16|5|Then Rezin king of Aram and Pekah son of Remaliah king of Israel marched up to fight against Jerusalem and besieged Ahaz, but they could not overpower him.
2KGS|16|6|At that time, Rezin king of Aram recovered Elath for Aram by driving out the men of Judah. Edomites then moved into Elath and have lived there to this day.
2KGS|16|7|Ahaz sent messengers to say to Tiglath-Pileser king of Assyria, "I am your servant and vassal. Come up and save me out of the hand of the king of Aram and of the king of Israel, who are attacking me."
2KGS|16|8|And Ahaz took the silver and gold found in the temple of the LORD and in the treasuries of the royal palace and sent it as a gift to the king of Assyria.
2KGS|16|9|The king of Assyria complied by attacking Damascus and capturing it. He deported its inhabitants to Kir and put Rezin to death.
2KGS|16|10|Then King Ahaz went to Damascus to meet Tiglath-Pileser king of Assyria. He saw an altar in Damascus and sent to Uriah the priest a sketch of the altar, with detailed plans for its construction.
2KGS|16|11|So Uriah the priest built an altar in accordance with all the plans that King Ahaz had sent from Damascus and finished it before King Ahaz returned.
2KGS|16|12|When the king came back from Damascus and saw the altar, he approached it and presented offerings on it.
2KGS|16|13|He offered up his burnt offering and grain offering, poured out his drink offering, and sprinkled the blood of his fellowship offerings on the altar.
2KGS|16|14|The bronze altar that stood before the LORD he brought from the front of the temple-from between the new altar and the temple of the LORD -and put it on the north side of the new altar.
2KGS|16|15|King Ahaz then gave these orders to Uriah the priest: "On the large new altar, offer the morning burnt offering and the evening grain offering, the king's burnt offering and his grain offering, and the burnt offering of all the people of the land, and their grain offering and their drink offering. Sprinkle on the altar all the blood of the burnt offerings and sacrifices. But I will use the bronze altar for seeking guidance."
2KGS|16|16|And Uriah the priest did just as King Ahaz had ordered.
2KGS|16|17|King Ahaz took away the side panels and removed the basins from the movable stands. He removed the Sea from the bronze bulls that supported it and set it on a stone base.
2KGS|16|18|He took away the Sabbath canopy that had been built at the temple and removed the royal entryway outside the temple of the LORD, in deference to the king of Assyria.
2KGS|16|19|As for the other events of the reign of Ahaz, and what he did, are they not written in the book of the annals of the kings of Judah?
2KGS|16|20|Ahaz rested with his fathers and was buried with them in the City of David. And Hezekiah his son succeeded him as king.
2KGS|17|1|In the twelfth year of Ahaz king of Judah, Hoshea son of Elah became king of Israel in Samaria, and he reigned nine years.
2KGS|17|2|He did evil in the eyes of the LORD, but not like the kings of Israel who preceded him.
2KGS|17|3|Shalmaneser king of Assyria came up to attack Hoshea, who had been Shalmaneser's vassal and had paid him tribute.
2KGS|17|4|But the king of Assyria discovered that Hoshea was a traitor, for he had sent envoys to So king of Egypt, and he no longer paid tribute to the king of Assyria, as he had done year by year. Therefore Shalmaneser seized him and put him in prison.
2KGS|17|5|The king of Assyria invaded the entire land, marched against Samaria and laid siege to it for three years.
2KGS|17|6|In the ninth year of Hoshea, the king of Assyria captured Samaria and deported the Israelites to Assyria. He settled them in Halah, in Gozan on the Habor River and in the towns of the Medes.
2KGS|17|7|All this took place because the Israelites had sinned against the LORD their God, who had brought them up out of Egypt from under the power of Pharaoh king of Egypt. They worshiped other gods
2KGS|17|8|and followed the practices of the nations the LORD had driven out before them, as well as the practices that the kings of Israel had introduced.
2KGS|17|9|The Israelites secretly did things against the LORD their God that were not right. From watchtower to fortified city they built themselves high places in all their towns.
2KGS|17|10|They set up sacred stones and Asherah poles on every high hill and under every spreading tree.
2KGS|17|11|At every high place they burned incense, as the nations whom the LORD had driven out before them had done. They did wicked things that provoked the LORD to anger.
2KGS|17|12|They worshiped idols, though the LORD had said, "You shall not do this."
2KGS|17|13|The LORD warned Israel and Judah through all his prophets and seers: "Turn from your evil ways. Observe my commands and decrees, in accordance with the entire Law that I commanded your fathers to obey and that I delivered to you through my servants the prophets."
2KGS|17|14|But they would not listen and were as stiff-necked as their fathers, who did not trust in the LORD their God.
2KGS|17|15|They rejected his decrees and the covenant he had made with their fathers and the warnings he had given them. They followed worthless idols and themselves became worthless. They imitated the nations around them although the LORD had ordered them, "Do not do as they do," and they did the things the LORD had forbidden them to do.
2KGS|17|16|They forsook all the commands of the LORD their God and made for themselves two idols cast in the shape of calves, and an Asherah pole. They bowed down to all the starry hosts, and they worshiped Baal.
2KGS|17|17|They sacrificed their sons and daughters in the fire. They practiced divination and sorcery and sold themselves to do evil in the eyes of the LORD, provoking him to anger.
2KGS|17|18|So the LORD was very angry with Israel and removed them from his presence. Only the tribe of Judah was left,
2KGS|17|19|and even Judah did not keep the commands of the LORD their God. They followed the practices Israel had introduced.
2KGS|17|20|Therefore the LORD rejected all the people of Israel; he afflicted them and gave them into the hands of plunderers, until he thrust them from his presence.
2KGS|17|21|When he tore Israel away from the house of David, they made Jeroboam son of Nebat their king. Jeroboam enticed Israel away from following the LORD and caused them to commit a great sin.
2KGS|17|22|The Israelites persisted in all the sins of Jeroboam and did not turn away from them
2KGS|17|23|until the LORD removed them from his presence, as he had warned through all his servants the prophets. So the people of Israel were taken from their homeland into exile in Assyria, and they are still there.
2KGS|17|24|The king of Assyria brought people from Babylon, Cuthah, Avva, Hamath and Sepharvaim and settled them in the towns of Samaria to replace the Israelites. They took over Samaria and lived in its towns.
2KGS|17|25|When they first lived there, they did not worship the LORD; so he sent lions among them and they killed some of the people.
2KGS|17|26|It was reported to the king of Assyria: "The people you deported and resettled in the towns of Samaria do not know what the god of that country requires. He has sent lions among them, which are killing them off, because the people do not know what he requires."
2KGS|17|27|Then the king of Assyria gave this order: "Have one of the priests you took captive from Samaria go back to live there and teach the people what the god of the land requires."
2KGS|17|28|So one of the priests who had been exiled from Samaria came to live in Bethel and taught them how to worship the LORD.
2KGS|17|29|Nevertheless, each national group made its own gods in the several towns where they settled, and set them up in the shrines the people of Samaria had made at the high places.
2KGS|17|30|The men from Babylon made Succoth Benoth, the men from Cuthah made Nergal, and the men from Hamath made Ashima;
2KGS|17|31|the Avvites made Nibhaz and Tartak, and the Sepharvites burned their children in the fire as sacrifices to Adrammelech and Anammelech, the gods of Sepharvaim.
2KGS|17|32|They worshiped the LORD, but they also appointed all sorts of their own people to officiate for them as priests in the shrines at the high places.
2KGS|17|33|They worshiped the LORD, but they also served their own gods in accordance with the customs of the nations from which they had been brought.
2KGS|17|34|To this day they persist in their former practices. They neither worship the LORD nor adhere to the decrees and ordinances, the laws and commands that the LORD gave the descendants of Jacob, whom he named Israel.
2KGS|17|35|When the LORD made a covenant with the Israelites, he commanded them: "Do not worship any other gods or bow down to them, serve them or sacrifice to them.
2KGS|17|36|But the LORD, who brought you up out of Egypt with mighty power and outstretched arm, is the one you must worship. To him you shall bow down and to him offer sacrifices.
2KGS|17|37|You must always be careful to keep the decrees and ordinances, the laws and commands he wrote for you. Do not worship other gods.
2KGS|17|38|Do not forget the covenant I have made with you, and do not worship other gods.
2KGS|17|39|Rather, worship the LORD your God; it is he who will deliver you from the hand of all your enemies."
2KGS|17|40|They would not listen, however, but persisted in their former practices.
2KGS|17|41|Even while these people were worshiping the LORD, they were serving their idols. To this day their children and grandchildren continue to do as their fathers did.
2KGS|18|1|In the third year of Hoshea son of Elah king of Israel, Hezekiah son of Ahaz king of Judah began to reign.
2KGS|18|2|He was twenty-five years old when he became king, and he reigned in Jerusalem twenty-nine years. His mother's name was Abijah daughter of Zechariah.
2KGS|18|3|He did what was right in the eyes of the LORD, just as his father David had done.
2KGS|18|4|He removed the high places, smashed the sacred stones and cut down the Asherah poles. He broke into pieces the bronze snake Moses had made, for up to that time the Israelites had been burning incense to it. (It was called Nehushtan. )
2KGS|18|5|Hezekiah trusted in the LORD, the God of Israel. There was no one like him among all the kings of Judah, either before him or after him.
2KGS|18|6|He held fast to the LORD and did not cease to follow him; he kept the commands the LORD had given Moses.
2KGS|18|7|And the LORD was with him; he was successful in whatever he undertook. He rebelled against the king of Assyria and did not serve him.
2KGS|18|8|From watchtower to fortified city, he defeated the Philistines, as far as Gaza and its territory.
2KGS|18|9|In King Hezekiah's fourth year, which was the seventh year of Hoshea son of Elah king of Israel, Shalmaneser king of Assyria marched against Samaria and laid siege to it.
2KGS|18|10|At the end of three years the Assyrians took it. So Samaria was captured in Hezekiah's sixth year, which was the ninth year of Hoshea king of Israel.
2KGS|18|11|The king of Assyria deported Israel to Assyria and settled them in Halah, in Gozan on the Habor River and in towns of the Medes.
2KGS|18|12|This happened because they had not obeyed the LORD their God, but had violated his covenant-all that Moses the servant of the LORD commanded. They neither listened to the commands nor carried them out.
2KGS|18|13|In the fourteenth year of King Hezekiah's reign, Sennacherib king of Assyria attacked all the fortified cities of Judah and captured them.
2KGS|18|14|So Hezekiah king of Judah sent this message to the king of Assyria at Lachish: "I have done wrong. Withdraw from me, and I will pay whatever you demand of me." The king of Assyria exacted from Hezekiah king of Judah three hundred talents of silver and thirty talents of gold.
2KGS|18|15|So Hezekiah gave him all the silver that was found in the temple of the LORD and in the treasuries of the royal palace.
2KGS|18|16|At this time Hezekiah king of Judah stripped off the gold with which he had covered the doors and doorposts of the temple of the LORD, and gave it to the king of Assyria.
2KGS|18|17|The king of Assyria sent his supreme commander, his chief officer and his field commander with a large army, from Lachish to King Hezekiah at Jerusalem. They came up to Jerusalem and stopped at the aqueduct of the Upper Pool, on the road to the Washerman's Field.
2KGS|18|18|They called for the king; and Eliakim son of Hilkiah the palace administrator, Shebna the secretary, and Joah son of Asaph the recorder went out to them.
2KGS|18|19|The field commander said to them, "Tell Hezekiah: "'This is what the great king, the king of Assyria, says: On what are you basing this confidence of yours?
2KGS|18|20|You say you have strategy and military strength-but you speak only empty words. On whom are you depending, that you rebel against me?
2KGS|18|21|Look now, you are depending on Egypt, that splintered reed of a staff, which pierces a man's hand and wounds him if he leans on it! Such is Pharaoh king of Egypt to all who depend on him.
2KGS|18|22|And if you say to me, "We are depending on the LORD our God"-isn't he the one whose high places and altars Hezekiah removed, saying to Judah and Jerusalem, "You must worship before this altar in Jerusalem"?
2KGS|18|23|"'Come now, make a bargain with my master, the king of Assyria: I will give you two thousand horses-if you can put riders on them!
2KGS|18|24|How can you repulse one officer of the least of my master's officials, even though you are depending on Egypt for chariots and horsemen?
2KGS|18|25|Furthermore, have I come to attack and destroy this place without word from the LORD? The LORD himself told me to march against this country and destroy it.'"
2KGS|18|26|Then Eliakim son of Hilkiah, and Shebna and Joah said to the field commander, "Please speak to your servants in Aramaic, since we understand it. Don't speak to us in Hebrew in the hearing of the people on the wall."
2KGS|18|27|But the commander replied, "Was it only to your master and you that my master sent me to say these things, and not to the men sitting on the wall-who, like you, will have to eat their own filth and drink their own urine?"
2KGS|18|28|Then the commander stood and called out in Hebrew: "Hear the word of the great king, the king of Assyria!
2KGS|18|29|This is what the king says: Do not let Hezekiah deceive you. He cannot deliver you from my hand.
2KGS|18|30|Do not let Hezekiah persuade you to trust in the LORD when he says, 'The LORD will surely deliver us; this city will not be given into the hand of the king of Assyria.'
2KGS|18|31|"Do not listen to Hezekiah. This is what the king of Assyria says: Make peace with me and come out to me. Then every one of you will eat from his own vine and fig tree and drink water from his own cistern,
2KGS|18|32|until I come and take you to a land like your own, a land of grain and new wine, a land of bread and vineyards, a land of olive trees and honey. Choose life and not death! "Do not listen to Hezekiah, for he is misleading you when he says, 'The LORD will deliver us.'
2KGS|18|33|Has the god of any nation ever delivered his land from the hand of the king of Assyria?
2KGS|18|34|Where are the gods of Hamath and Arpad? Where are the gods of Sepharvaim, Hena and Ivvah? Have they rescued Samaria from my hand?
2KGS|18|35|Who of all the gods of these countries has been able to save his land from me? How then can the LORD deliver Jerusalem from my hand?"
2KGS|18|36|But the people remained silent and said nothing in reply, because the king had commanded, "Do not answer him."
2KGS|18|37|Then Eliakim son of Hilkiah the palace administrator, Shebna the secretary and Joah son of Asaph the recorder went to Hezekiah, with their clothes torn, and told him what the field commander had said.
2KGS|19|1|When King Hezekiah heard this, he tore his clothes and put on sackcloth and went into the temple of the LORD.
2KGS|19|2|He sent Eliakim the palace administrator, Shebna the secretary and the leading priests, all wearing sackcloth, to the prophet Isaiah son of Amoz.
2KGS|19|3|They told him, "This is what Hezekiah says: This day is a day of distress and rebuke and disgrace, as when children come to the point of birth and there is no strength to deliver them.
2KGS|19|4|It may be that the LORD your God will hear all the words of the field commander, whom his master, the king of Assyria, has sent to ridicule the living God, and that he will rebuke him for the words the LORD your God has heard. Therefore pray for the remnant that still survives."
2KGS|19|5|When King Hezekiah's officials came to Isaiah,
2KGS|19|6|Isaiah said to them, "Tell your master, 'This is what the LORD says: Do not be afraid of what you have heard-those words with which the underlings of the king of Assyria have blasphemed me.
2KGS|19|7|Listen! I am going to put such a spirit in him that when he hears a certain report, he will return to his own country, and there I will have him cut down with the sword.'"
2KGS|19|8|When the field commander heard that the king of Assyria had left Lachish, he withdrew and found the king fighting against Libnah.
2KGS|19|9|Now Sennacherib received a report that Tirhakah, the Cushite king of Egypt, was marching out to fight against him. So he again sent messengers to Hezekiah with this word:
2KGS|19|10|"Say to Hezekiah king of Judah: Do not let the god you depend on deceive you when he says, 'Jerusalem will not be handed over to the king of Assyria.'
2KGS|19|11|Surely you have heard what the kings of Assyria have done to all the countries, destroying them completely. And will you be delivered?
2KGS|19|12|Did the gods of the nations that were destroyed by my forefathers deliver them: the gods of Gozan, Haran, Rezeph and the people of Eden who were in Tel Assar?
2KGS|19|13|Where is the king of Hamath, the king of Arpad, the king of the city of Sepharvaim, or of Hena or Ivvah?"
2KGS|19|14|Hezekiah received the letter from the messengers and read it. Then he went up to the temple of the LORD and spread it out before the LORD.
2KGS|19|15|And Hezekiah prayed to the LORD: "O LORD, God of Israel, enthroned between the cherubim, you alone are God over all the kingdoms of the earth. You have made heaven and earth.
2KGS|19|16|Give ear, O LORD, and hear; open your eyes, O LORD, and see; listen to the words Sennacherib has sent to insult the living God.
2KGS|19|17|"It is true, O LORD, that the Assyrian kings have laid waste these nations and their lands.
2KGS|19|18|They have thrown their gods into the fire and destroyed them, for they were not gods but only wood and stone, fashioned by men's hands.
2KGS|19|19|Now, O LORD our God, deliver us from his hand, so that all kingdoms on earth may know that you alone, O LORD, are God."
2KGS|19|20|Then Isaiah son of Amoz sent a message to Hezekiah: "This is what the LORD, the God of Israel, says: I have heard your prayer concerning Sennacherib king of Assyria.
2KGS|19|21|This is the word that the LORD has spoken against him: "'The Virgin Daughter of Zion despises you and mocks you. The Daughter of Jerusalem tosses her head as you flee.
2KGS|19|22|Who is it you have insulted and blasphemed? Against whom have you raised your voice and lifted your eyes in pride? Against the Holy One of Israel!
2KGS|19|23|By your messengers you have heaped insults on the Lord. And you have said, "With my many chariots I have ascended the heights of the mountains, the utmost heights of Lebanon. I have cut down its tallest cedars, the choicest of its pines. I have reached its remotest parts, the finest of its forests.
2KGS|19|24|I have dug wells in foreign lands and drunk the water there. With the soles of my feet I have dried up all the streams of Egypt."
2KGS|19|25|"'Have you not heard? Long ago I ordained it. In days of old I planned it; now I have brought it to pass, that you have turned fortified cities into piles of stone.
2KGS|19|26|Their people, drained of power, are dismayed and put to shame. They are like plants in the field, like tender green shoots, like grass sprouting on the roof, scorched before it grows up.
2KGS|19|27|"'But I know where you stay and when you come and go and how you rage against me.
2KGS|19|28|Because you rage against me and your insolence has reached my ears, I will put my hook in your nose and my bit in your mouth, and I will make you return by the way you came.'
2KGS|19|29|"This will be the sign for you, O Hezekiah: "This year you will eat what grows by itself, and the second year what springs from that. But in the third year sow and reap, plant vineyards and eat their fruit.
2KGS|19|30|Once more a remnant of the house of Judah will take root below and bear fruit above.
2KGS|19|31|For out of Jerusalem will come a remnant, and out of Mount Zion a band of survivors. The zeal of the LORD Almighty will accomplish this.
2KGS|19|32|"Therefore this is what the LORD says concerning the king of Assyria: "He will not enter this city or shoot an arrow here. He will not come before it with shield or build a siege ramp against it.
2KGS|19|33|By the way that he came he will return; he will not enter this city, declares the LORD.
2KGS|19|34|I will defend this city and save it, for my sake and for the sake of David my servant."
2KGS|19|35|That night the angel of the LORD went out and put to death a hundred and eighty-five thousand men in the Assyrian camp. When the people got up the next morning-there were all the dead bodies!
2KGS|19|36|So Sennacherib king of Assyria broke camp and withdrew. He returned to Nineveh and stayed there.
2KGS|19|37|One day, while he was worshiping in the temple of his god Nisroch, his sons Adrammelech and Sharezer cut him down with the sword, and they escaped to the land of Ararat. And Esarhaddon his son succeeded him as king.
2KGS|20|1|In those days Hezekiah became ill and was at the point of death. The prophet Isaiah son of Amoz went to him and said, "This is what the LORD says: Put your house in order, because you are going to die; you will not recover."
2KGS|20|2|Hezekiah turned his face to the wall and prayed to the LORD,
2KGS|20|3|"Remember, O LORD, how I have walked before you faithfully and with wholehearted devotion and have done what is good in your eyes." And Hezekiah wept bitterly.
2KGS|20|4|Before Isaiah had left the middle court, the word of the LORD came to him:
2KGS|20|5|"Go back and tell Hezekiah, the leader of my people, 'This is what the LORD, the God of your father David, says: I have heard your prayer and seen your tears; I will heal you. On the third day from now you will go up to the temple of the LORD.
2KGS|20|6|I will add fifteen years to your life. And I will deliver you and this city from the hand of the king of Assyria. I will defend this city for my sake and for the sake of my servant David.'"
2KGS|20|7|Then Isaiah said, "Prepare a poultice of figs." They did so and applied it to the boil, and he recovered.
2KGS|20|8|Hezekiah had asked Isaiah, "What will be the sign that the LORD will heal me and that I will go up to the temple of the LORD on the third day from now?"
2KGS|20|9|Isaiah answered, "This is the LORD's sign to you that the LORD will do what he has promised: Shall the shadow go forward ten steps, or shall it go back ten steps?"
2KGS|20|10|"It is a simple matter for the shadow to go forward ten steps," said Hezekiah. "Rather, have it go back ten steps."
2KGS|20|11|Then the prophet Isaiah called upon the LORD, and the LORD made the shadow go back the ten steps it had gone down on the stairway of Ahaz.
2KGS|20|12|At that time Merodach-Baladan son of Baladan king of Babylon sent Hezekiah letters and a gift, because he had heard of Hezekiah's illness.
2KGS|20|13|Hezekiah received the messengers and showed them all that was in his storehouses-the silver, the gold, the spices and the fine oil-his armory and everything found among his treasures. There was nothing in his palace or in all his kingdom that Hezekiah did not show them.
2KGS|20|14|Then Isaiah the prophet went to King Hezekiah and asked, "What did those men say, and where did they come from?From a distant land," Hezekiah replied. "They came from Babylon."
2KGS|20|15|The prophet asked, "What did they see in your palace?They saw everything in my palace," Hezekiah said. "There is nothing among my treasures that I did not show them."
2KGS|20|16|Then Isaiah said to Hezekiah, "Hear the word of the LORD:
2KGS|20|17|The time will surely come when everything in your palace, and all that your fathers have stored up until this day, will be carried off to Babylon. Nothing will be left, says the LORD.
2KGS|20|18|And some of your descendants, your own flesh and blood, that will be born to you, will be taken away, and they will become eunuchs in the palace of the king of Babylon."
2KGS|20|19|"The word of the LORD you have spoken is good," Hezekiah replied. For he thought, "Will there not be peace and security in my lifetime?"
2KGS|20|20|As for the other events of Hezekiah's reign, all his achievements and how he made the pool and the tunnel by which he brought water into the city, are they not written in the book of the annals of the kings of Judah?
2KGS|20|21|Hezekiah rested with his fathers. And Manasseh his son succeeded him as king.
2KGS|21|1|Manasseh was twelve years old when he became king, and he reigned in Jerusalem fifty-five years. His mother's name was Hephzibah.
2KGS|21|2|He did evil in the eyes of the LORD, following the detestable practices of the nations the LORD had driven out before the Israelites.
2KGS|21|3|He rebuilt the high places his father Hezekiah had destroyed; he also erected altars to Baal and made an Asherah pole, as Ahab king of Israel had done. He bowed down to all the starry hosts and worshiped them.
2KGS|21|4|He built altars in the temple of the LORD, of which the LORD had said, "In Jerusalem I will put my Name."
2KGS|21|5|In both courts of the temple of the LORD, he built altars to all the starry hosts.
2KGS|21|6|He sacrificed his own son in the fire, practiced sorcery and divination, and consulted mediums and spiritists. He did much evil in the eyes of the LORD, provoking him to anger.
2KGS|21|7|He took the carved Asherah pole he had made and put it in the temple, of which the LORD had said to David and to his son Solomon, "In this temple and in Jerusalem, which I have chosen out of all the tribes of Israel, I will put my Name forever.
2KGS|21|8|I will not again make the feet of the Israelites wander from the land I gave their forefathers, if only they will be careful to do everything I commanded them and will keep the whole Law that my servant Moses gave them."
2KGS|21|9|But the people did not listen. Manasseh led them astray, so that they did more evil than the nations the LORD had destroyed before the Israelites.
2KGS|21|10|The LORD said through his servants the prophets:
2KGS|21|11|"Manasseh king of Judah has committed these detestable sins. He has done more evil than the Amorites who preceded him and has led Judah into sin with his idols.
2KGS|21|12|Therefore this is what the LORD, the God of Israel, says: I am going to bring such disaster on Jerusalem and Judah that the ears of everyone who hears of it will tingle.
2KGS|21|13|I will stretch out over Jerusalem the measuring line used against Samaria and the plumb line used against the house of Ahab. I will wipe out Jerusalem as one wipes a dish, wiping it and turning it upside down.
2KGS|21|14|I will forsake the remnant of my inheritance and hand them over to their enemies. They will be looted and plundered by all their foes,
2KGS|21|15|because they have done evil in my eyes and have provoked me to anger from the day their forefathers came out of Egypt until this day."
2KGS|21|16|Moreover, Manasseh also shed so much innocent blood that he filled Jerusalem from end to end-besides the sin that he had caused Judah to commit, so that they did evil in the eyes of the LORD.
2KGS|21|17|As for the other events of Manasseh's reign, and all he did, including the sin he committed, are they not written in the book of the annals of the kings of Judah?
2KGS|21|18|Manasseh rested with his fathers and was buried in his palace garden, the garden of Uzza. And Amon his son succeeded him as king.
2KGS|21|19|Amon was twenty-two years old when he became king, and he reigned in Jerusalem two years. His mother's name was Meshullemeth daughter of Haruz; she was from Jotbah.
2KGS|21|20|He did evil in the eyes of the LORD, as his father Manasseh had done.
2KGS|21|21|He walked in all the ways of his father; he worshiped the idols his father had worshiped, and bowed down to them.
2KGS|21|22|He forsook the LORD, the God of his fathers, and did not walk in the way of the LORD.
2KGS|21|23|Amon's officials conspired against him and assassinated the king in his palace.
2KGS|21|24|Then the people of the land killed all who had plotted against King Amon, and they made Josiah his son king in his place.
2KGS|21|25|As for the other events of Amon's reign, and what he did, are they not written in the book of the annals of the kings of Judah?
2KGS|21|26|He was buried in his grave in the garden of Uzza. And Josiah his son succeeded him as king.
2KGS|22|1|Josiah was eight years old when he became king, and he reigned in Jerusalem thirty-one years. His mother's name was Jedidah daughter of Adaiah; she was from Bozkath.
2KGS|22|2|He did what was right in the eyes of the LORD and walked in all the ways of his father David, not turning aside to the right or to the left.
2KGS|22|3|In the eighteenth year of his reign, King Josiah sent the secretary, Shaphan son of Azaliah, the son of Meshullam, to the temple of the LORD. He said:
2KGS|22|4|"Go up to Hilkiah the high priest and have him get ready the money that has been brought into the temple of the LORD, which the doorkeepers have collected from the people.
2KGS|22|5|Have them entrust it to the men appointed to supervise the work on the temple. And have these men pay the workers who repair the temple of the LORD -
2KGS|22|6|the carpenters, the builders and the masons. Also have them purchase timber and dressed stone to repair the temple.
2KGS|22|7|But they need not account for the money entrusted to them, because they are acting faithfully."
2KGS|22|8|Hilkiah the high priest said to Shaphan the secretary, "I have found the Book of the Law in the temple of the LORD." He gave it to Shaphan, who read it.
2KGS|22|9|Then Shaphan the secretary went to the king and reported to him: "Your officials have paid out the money that was in the temple of the LORD and have entrusted it to the workers and supervisors at the temple."
2KGS|22|10|Then Shaphan the secretary informed the king, "Hilkiah the priest has given me a book." And Shaphan read from it in the presence of the king.
2KGS|22|11|When the king heard the words of the Book of the Law, he tore his robes.
2KGS|22|12|He gave these orders to Hilkiah the priest, Ahikam son of Shaphan, Acbor son of Micaiah, Shaphan the secretary and Asaiah the king's attendant:
2KGS|22|13|"Go and inquire of the LORD for me and for the people and for all Judah about what is written in this book that has been found. Great is the LORD's anger that burns against us because our fathers have not obeyed the words of this book; they have not acted in accordance with all that is written there concerning us."
2KGS|22|14|Hilkiah the priest, Ahikam, Acbor, Shaphan and Asaiah went to speak to the prophetess Huldah, who was the wife of Shallum son of Tikvah, the son of Harhas, keeper of the wardrobe. She lived in Jerusalem, in the Second District.
2KGS|22|15|She said to them, "This is what the LORD, the God of Israel, says: Tell the man who sent you to me,
2KGS|22|16|'This is what the LORD says: I am going to bring disaster on this place and its people, according to everything written in the book the king of Judah has read.
2KGS|22|17|Because they have forsaken me and burned incense to other gods and provoked me to anger by all the idols their hands have made, my anger will burn against this place and will not be quenched.'
2KGS|22|18|Tell the king of Judah, who sent you to inquire of the LORD, 'This is what the LORD, the God of Israel, says concerning the words you heard:
2KGS|22|19|Because your heart was responsive and you humbled yourself before the LORD when you heard what I have spoken against this place and its people, that they would become accursed and laid waste, and because you tore your robes and wept in my presence, I have heard you, declares the LORD.
2KGS|22|20|Therefore I will gather you to your fathers, and you will be buried in peace. Your eyes will not see all the disaster I am going to bring on this place.'" So they took her answer back to the king.
2KGS|23|1|Then the king called together all the elders of Judah and Jerusalem.
2KGS|23|2|He went up to the temple of the LORD with the men of Judah, the people of Jerusalem, the priests and the prophets-all the people from the least to the greatest. He read in their hearing all the words of the Book of the Covenant, which had been found in the temple of the LORD.
2KGS|23|3|The king stood by the pillar and renewed the covenant in the presence of the LORD -to follow the LORD and keep his commands, regulations and decrees with all his heart and all his soul, thus confirming the words of the covenant written in this book. Then all the people pledged themselves to the covenant.
2KGS|23|4|The king ordered Hilkiah the high priest, the priests next in rank and the doorkeepers to remove from the temple of the LORD all the articles made for Baal and Asherah and all the starry hosts. He burned them outside Jerusalem in the fields of the Kidron Valley and took the ashes to Bethel.
2KGS|23|5|He did away with the pagan priests appointed by the kings of Judah to burn incense on the high places of the towns of Judah and on those around Jerusalem-those who burned incense to Baal, to the sun and moon, to the constellations and to all the starry hosts.
2KGS|23|6|He took the Asherah pole from the temple of the LORD to the Kidron Valley outside Jerusalem and burned it there. He ground it to powder and scattered the dust over the graves of the common people.
2KGS|23|7|He also tore down the quarters of the male shrine prostitutes, which were in the temple of the LORD and where women did weaving for Asherah.
2KGS|23|8|Josiah brought all the priests from the towns of Judah and desecrated the high places, from Geba to Beersheba, where the priests had burned incense. He broke down the shrines at the gates-at the entrance to the Gate of Joshua, the city governor, which is on the left of the city gate.
2KGS|23|9|Although the priests of the high places did not serve at the altar of the LORD in Jerusalem, they ate unleavened bread with their fellow priests.
2KGS|23|10|He desecrated Topheth, which was in the Valley of Ben Hinnom, so no one could use it to sacrifice his son or daughter in the fire to Molech.
2KGS|23|11|He removed from the entrance to the temple of the LORD the horses that the kings of Judah had dedicated to the sun. They were in the court near the room of an official named Nathan-Melech. Josiah then burned the chariots dedicated to the sun.
2KGS|23|12|He pulled down the altars the kings of Judah had erected on the roof near the upper room of Ahaz, and the altars Manasseh had built in the two courts of the temple of the LORD. He removed them from there, smashed them to pieces and threw the rubble into the Kidron Valley.
2KGS|23|13|The king also desecrated the high places that were east of Jerusalem on the south of the Hill of Corruption-the ones Solomon king of Israel had built for Ashtoreth the vile goddess of the Sidonians, for Chemosh the vile god of Moab, and for Molech the detestable god of the people of Ammon.
2KGS|23|14|Josiah smashed the sacred stones and cut down the Asherah poles and covered the sites with human bones.
2KGS|23|15|Even the altar at Bethel, the high place made by Jeroboam son of Nebat, who had caused Israel to sin-even that altar and high place he demolished. He burned the high place and ground it to powder, and burned the Asherah pole also.
2KGS|23|16|Then Josiah looked around, and when he saw the tombs that were there on the hillside, he had the bones removed from them and burned on the altar to defile it, in accordance with the word of the LORD proclaimed by the man of God who foretold these things.
2KGS|23|17|The king asked, "What is that tombstone I see?" The men of the city said, "It marks the tomb of the man of God who came from Judah and pronounced against the altar of Bethel the very things you have done to it."
2KGS|23|18|"Leave it alone," he said. "Don't let anyone disturb his bones." So they spared his bones and those of the prophet who had come from Samaria.
2KGS|23|19|Just as he had done at Bethel, Josiah removed and defiled all the shrines at the high places that the kings of Israel had built in the towns of Samaria that had provoked the LORD to anger.
2KGS|23|20|Josiah slaughtered all the priests of those high places on the altars and burned human bones on them. Then he went back to Jerusalem.
2KGS|23|21|The king gave this order to all the people: "Celebrate the Passover to the LORD your God, as it is written in this Book of the Covenant."
2KGS|23|22|Not since the days of the judges who led Israel, nor throughout the days of the kings of Israel and the kings of Judah, had any such Passover been observed.
2KGS|23|23|But in the eighteenth year of King Josiah, this Passover was celebrated to the LORD in Jerusalem.
2KGS|23|24|Furthermore, Josiah got rid of the mediums and spiritists, the household gods, the idols and all the other detestable things seen in Judah and Jerusalem. This he did to fulfill the requirements of the law written in the book that Hilkiah the priest had discovered in the temple of the LORD.
2KGS|23|25|Neither before nor after Josiah was there a king like him who turned to the LORD as he did-with all his heart and with all his soul and with all his strength, in accordance with all the Law of Moses.
2KGS|23|26|Nevertheless, the LORD did not turn away from the heat of his fierce anger, which burned against Judah because of all that Manasseh had done to provoke him to anger.
2KGS|23|27|So the LORD said, "I will remove Judah also from my presence as I removed Israel, and I will reject Jerusalem, the city I chose, and this temple, about which I said, 'There shall my Name be.'"
2KGS|23|28|As for the other events of Josiah's reign, and all he did, are they not written in the book of the annals of the kings of Judah?
2KGS|23|29|While Josiah was king, Pharaoh Neco king of Egypt went up to the Euphrates River to help the king of Assyria. King Josiah marched out to meet him in battle, but Neco faced him and killed him at Megiddo.
2KGS|23|30|Josiah's servants brought his body in a chariot from Megiddo to Jerusalem and buried him in his own tomb. And the people of the land took Jehoahaz son of Josiah and anointed him and made him king in place of his father.
2KGS|23|31|Jehoahaz was twenty-three years old when he became king, and he reigned in Jerusalem three months. His mother's name was Hamutal daughter of Jeremiah; she was from Libnah.
2KGS|23|32|He did evil in the eyes of the LORD, just as his fathers had done.
2KGS|23|33|Pharaoh Neco put him in chains at Riblah in the land of Hamath so that he might not reign in Jerusalem, and he imposed on Judah a levy of a hundred talents of silver and a talent of gold.
2KGS|23|34|Pharaoh Neco made Eliakim son of Josiah king in place of his father Josiah and changed Eliakim's name to Jehoiakim. But he took Jehoahaz and carried him off to Egypt, and there he died.
2KGS|23|35|Jehoiakim paid Pharaoh Neco the silver and gold he demanded. In order to do so, he taxed the land and exacted the silver and gold from the people of the land according to their assessments.
2KGS|23|36|Jehoiakim was twenty-five years old when he became king, and he reigned in Jerusalem eleven years. His mother's name was Zebidah daughter of Pedaiah; she was from Rumah.
2KGS|23|37|And he did evil in the eyes of the LORD, just as his fathers had done.
2KGS|24|1|During Jehoiakim's reign, Nebuchadnezzar king of Babylon invaded the land, and Jehoiakim became his vassal for three years. But then he changed his mind and rebelled against Nebuchadnezzar.
2KGS|24|2|The LORD sent Babylonian, Aramean, Moabite and Ammonite raiders against him. He sent them to destroy Judah, in accordance with the word of the LORD proclaimed by his servants the prophets.
2KGS|24|3|Surely these things happened to Judah according to the LORD's command, in order to remove them from his presence because of the sins of Manasseh and all he had done,
2KGS|24|4|including the shedding of innocent blood. For he had filled Jerusalem with innocent blood, and the LORD was not willing to forgive.
2KGS|24|5|As for the other events of Jehoiakim's reign, and all he did, are they not written in the book of the annals of the kings of Judah?
2KGS|24|6|Jehoiakim rested with his fathers. And Jehoiachin his son succeeded him as king.
2KGS|24|7|The king of Egypt did not march out from his own country again, because the king of Babylon had taken all his territory, from the Wadi of Egypt to the Euphrates River.
2KGS|24|8|Jehoiachin was eighteen years old when he became king, and he reigned in Jerusalem three months. His mother's name was Nehushta daughter of Elnathan; she was from Jerusalem.
2KGS|24|9|He did evil in the eyes of the LORD, just as his father had done.
2KGS|24|10|At that time the officers of Nebuchadnezzar king of Babylon advanced on Jerusalem and laid siege to it,
2KGS|24|11|and Nebuchadnezzar himself came up to the city while his officers were besieging it.
2KGS|24|12|Jehoiachin king of Judah, his mother, his attendants, his nobles and his officials all surrendered to him. In the eighth year of the reign of the king of Babylon, he took Jehoiachin prisoner.
2KGS|24|13|As the LORD had declared, Nebuchadnezzar removed all the treasures from the temple of the LORD and from the royal palace, and took away all the gold articles that Solomon king of Israel had made for the temple of the LORD.
2KGS|24|14|He carried into exile all Jerusalem: all the officers and fighting men, and all the craftsmen and artisans-a total of ten thousand. Only the poorest people of the land were left.
2KGS|24|15|Nebuchadnezzar took Jehoiachin captive to Babylon. He also took from Jerusalem to Babylon the king's mother, his wives, his officials and the leading men of the land.
2KGS|24|16|The king of Babylon also deported to Babylon the entire force of seven thousand fighting men, strong and fit for war, and a thousand craftsmen and artisans.
2KGS|24|17|He made Mattaniah, Jehoiachin's uncle, king in his place and changed his name to Zedekiah.
2KGS|24|18|Zedekiah was twenty-one years old when he became king, and he reigned in Jerusalem eleven years. His mother's name was Hamutal daughter of Jeremiah; she was from Libnah.
2KGS|24|19|He did evil in the eyes of the LORD, just as Jehoiakim had done.
2KGS|24|20|It was because of the LORD's anger that all this happened to Jerusalem and Judah, and in the end he thrust them from his presence. Now Zedekiah rebelled against the king of Babylon.
2KGS|25|1|So in the ninth year of Zedekiah's reign, on the tenth day of the tenth month, Nebuchadnezzar king of Babylon marched against Jerusalem with his whole army. He encamped outside the city and built siege works all around it.
2KGS|25|2|The city was kept under siege until the eleventh year of King Zedekiah.
2KGS|25|3|By the ninth day of the fourth month the famine in the city had become so severe that there was no food for the people to eat.
2KGS|25|4|Then the city wall was broken through, and the whole army fled at night through the gate between the two walls near the king's garden, though the Babylonians were surrounding the city. They fled toward the Arabah,
2KGS|25|5|but the Babylonian army pursued the king and overtook him in the plains of Jericho. All his soldiers were separated from him and scattered,
2KGS|25|6|and he was captured. He was taken to the king of Babylon at Riblah, where sentence was pronounced on him.
2KGS|25|7|They killed the sons of Zedekiah before his eyes. Then they put out his eyes, bound him with bronze shackles and took him to Babylon.
2KGS|25|8|On the seventh day of the fifth month, in the nineteenth year of Nebuchadnezzar king of Babylon, Nebuzaradan commander of the imperial guard, an official of the king of Babylon, came to Jerusalem.
2KGS|25|9|He set fire to the temple of the LORD, the royal palace and all the houses of Jerusalem. Every important building he burned down.
2KGS|25|10|The whole Babylonian army, under the commander of the imperial guard, broke down the walls around Jerusalem.
2KGS|25|11|Nebuzaradan the commander of the guard carried into exile the people who remained in the city, along with the rest of the populace and those who had gone over to the king of Babylon.
2KGS|25|12|But the commander left behind some of the poorest people of the land to work the vineyards and fields.
2KGS|25|13|The Babylonians broke up the bronze pillars, the movable stands and the bronze Sea that were at the temple of the LORD and they carried the bronze to Babylon.
2KGS|25|14|They also took away the pots, shovels, wick trimmers, dishes and all the bronze articles used in the temple service.
2KGS|25|15|The commander of the imperial guard took away the censers and sprinkling bowls-all that were made of pure gold or silver.
2KGS|25|16|The bronze from the two pillars, the Sea and the movable stands, which Solomon had made for the temple of the LORD, was more than could be weighed.
2KGS|25|17|Each pillar was twenty-seven feet high. The bronze capital on top of one pillar was four and a half feet high and was decorated with a network and pomegranates of bronze all around. The other pillar, with its network, was similar.
2KGS|25|18|The commander of the guard took as prisoners Seraiah the chief priest, Zephaniah the priest next in rank and the three doorkeepers.
2KGS|25|19|Of those still in the city, he took the officer in charge of the fighting men and five royal advisers. He also took the secretary who was chief officer in charge of conscripting the people of the land and sixty of his men who were found in the city.
2KGS|25|20|Nebuzaradan the commander took them all and brought them to the king of Babylon at Riblah.
2KGS|25|21|There at Riblah, in the land of Hamath, the king had them executed. So Judah went into captivity, away from her land.
2KGS|25|22|Nebuchadnezzar king of Babylon appointed Gedaliah son of Ahikam, the son of Shaphan, to be over the people he had left behind in Judah.
2KGS|25|23|When all the army officers and their men heard that the king of Babylon had appointed Gedaliah as governor, they came to Gedaliah at Mizpah-Ishmael son of Nethaniah, Johanan son of Kareah, Seraiah son of Tanhumeth the Netophathite, Jaazaniah the son of the Maacathite, and their men.
2KGS|25|24|Gedaliah took an oath to reassure them and their men. "Do not be afraid of the Babylonian officials," he said. "Settle down in the land and serve the king of Babylon, and it will go well with you."
2KGS|25|25|In the seventh month, however, Ishmael son of Nethaniah, the son of Elishama, who was of royal blood, came with ten men and assassinated Gedaliah and also the men of Judah and the Babylonians who were with him at Mizpah.
2KGS|25|26|At this, all the people from the least to the greatest, together with the army officers, fled to Egypt for fear of the Babylonians.
2KGS|25|27|In the thirty-seventh year of the exile of Jehoiachin king of Judah, in the year Evil-Merodach became king of Babylon, he released Jehoiachin from prison on the twenty-seventh day of the twelfth month.
2KGS|25|28|He spoke kindly to him and gave him a seat of honor higher than those of the other kings who were with him in Babylon.
2KGS|25|29|So Jehoiachin put aside his prison clothes and for the rest of his life ate regularly at the king's table.
2KGS|25|30|Day by day the king gave Jehoiachin a regular allowance as long as he lived.
