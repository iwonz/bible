RUTH|1|1|В те дни, когда управляли судьи, случился голод на земле. И пошел один человек из Вифлеема Иудейского со своею женою и двумя сыновьями своими жить на полях Моавитских.
RUTH|1|2|Имя человека того Елимелех, имя жены его Ноеминь, а имена двух сынов его Махлон и Хилеон; [они были] Ефрафяне из Вифлеема Иудейского. И пришли они на поля Моавитские и остались там.
RUTH|1|3|И умер Елимелех, муж Ноемини, и осталась она с двумя сыновьями своими.
RUTH|1|4|Они взяли себе жен из Моавитянок, имя одной Орфа, а имя другой Руфь, и жили там около десяти лет.
RUTH|1|5|Но потом и оба [сына ее], Махлон и Хилеон, умерли, и осталась та женщина после обоих своих сыновей и после мужа своего.
RUTH|1|6|И встала она со снохами своими и пошла обратно с полей Моавитских, ибо услышала на полях Моавитских, что Бог посетил народ Свой и дал им хлеб.
RUTH|1|7|И вышла она из того места, в котором жила, и обе снохи ее с нею. Когда они шли по дороге, возвращаясь в землю Иудейскую,
RUTH|1|8|Ноеминь сказала двум снохам своим: пойдите, возвратитесь каждая в дом матери своей; да сотворит Господь с вами милость, как вы поступали с умершими и со мною!
RUTH|1|9|да даст вам Господь, чтобы вы нашли пристанище каждая в доме своего мужа! И поцеловала их. Но они подняли вопль и плакали
RUTH|1|10|и сказали: нет, мы с тобою возвратимся к народу твоему.
RUTH|1|11|Ноеминь же сказала: возвратитесь, дочери мои; зачем вам идти со мною? Разве еще есть у меня сыновья в моем чреве, которые были бы вам мужьями?
RUTH|1|12|Возвратитесь, дочери мои, пойдите, ибо я уже стара, чтоб быть замужем. Да если б я и сказала: "есть мне еще надежда", и даже если бы я сию же ночь была с мужем и потом родила сыновей, –
RUTH|1|13|то можно ли вам ждать, пока они выросли бы? можно ли вам медлить и не выходить замуж? Нет, дочери мои, я весьма сокрушаюсь о вас, ибо рука Господня постигла меня.
RUTH|1|14|Они подняли вопль и опять стали плакать. И Орфа простилась со свекровью своею, а Руфь осталась с нею.
RUTH|1|15|[Ноеминь] сказала [Руфи]: вот, невестка твоя возвратилась к народу своему и к своим богам; возвратись и ты вслед за невесткою твоею.
RUTH|1|16|Но Руфь сказала: не принуждай меня оставить тебя и возвратиться от тебя; но куда ты пойдешь, туда и я пойду, и где ты жить будешь, там и я буду жить; народ твой будет моим народом, и твой Бог – моим Богом;
RUTH|1|17|и где ты умрешь, там и я умру и погребена буду; пусть то и то сделает мне Господь, и еще больше сделает; смерть одна разлучит меня с тобою.
RUTH|1|18|[Ноеминь], видя, что она твердо решилась идти с нею, перестала уговаривать ее.
RUTH|1|19|И шли обе они, доколе не пришли в Вифлеем. Когда пришли они в Вифлеем, весь город пришел в движение от них, и говорили: это Ноеминь?
RUTH|1|20|Она сказала им: не называйте меня Ноеминью, а называйте меня Марою, потому что Вседержитель послал мне великую горесть;
RUTH|1|21|я вышла отсюда с достатком, а возвратил меня Господь с пустыми руками; зачем называть меня Ноеминью, когда Господь заставил меня страдать, и Вседержитель послал мне несчастье?
RUTH|1|22|И возвратилась Ноеминь, и с нею сноха ее Руфь Моавитянка, пришедшая с полей Моавитских, и пришли они в Вифлеем в начале жатвы ячменя.
RUTH|2|1|У Ноемини был родственник по мужу ее, человек весьма знатный, из племени Елимелехова, имя ему Вооз.
RUTH|2|2|И сказала Руфь Моавитянка Ноемини: пойду я на поле и буду подбирать колосья по следам того, у кого найду благоволение. Она сказала ей: пойди, дочь моя.
RUTH|2|3|Она пошла, и пришла, и подбирала в поле [колосья] позади жнецов. И случилось, что та часть поля принадлежала Воозу, который из племени Елимелехова.
RUTH|2|4|И вот, Вооз пришел из Вифлеема и сказал жнецам: Господь с вами! Они сказали ему: да благословит тебя Господь!
RUTH|2|5|И сказал Вооз слуге своему, приставленному к жнецам: чья это молодая женщина?
RUTH|2|6|Слуга, приставленный к жнецам, отвечал и сказал: эта молодая женщина – Моавитянка, пришедшая с Ноеминью с полей Моавитских;
RUTH|2|7|она сказала: "буду я подбирать и собирать между снопами позади жнецов"; и пришла, и находится [здесь] с самого утра доселе; мало бывает она дома.
RUTH|2|8|И сказал Вооз Руфи: послушай, дочь моя, не ходи подбирать на другом поле и не переходи отсюда, но будь здесь с моими служанками;
RUTH|2|9|пусть в глазах твоих будет то поле, где они жнут, и ходи за ними; вот, я приказал слугам моим не трогать тебя; когда захочешь пить, иди к сосудам и пей, откуда черпают слуги мои.
RUTH|2|10|Она пала на лице свое и поклонилась до земли и сказала ему: чем снискала я в глазах твоих милость, что ты принимаешь меня, хотя я и чужеземка?
RUTH|2|11|Вооз отвечал и сказал ей: мне сказано все, что сделала ты для свекрови своей по смерти мужа твоего, что ты оставила твоего отца и твою мать и твою родину и пришла к народу, которого ты не знала вчера и третьего дня;
RUTH|2|12|да воздаст Господь за это дело твое, и да будет тебе полная награда от Господа Бога Израилева, к Которому ты пришла, чтоб успокоиться под Его крылами!
RUTH|2|13|Она сказала: да буду я в милости пред очами твоими, господин мой! Ты утешил меня и говорил по сердцу рабы твоей, между тем как я не стою ни одной из рабынь твоих.
RUTH|2|14|И сказал ей Вооз: время обеда; приди сюда и ешь хлеб и обмакивай кусок твой в уксус. И села она возле жнецов. Он подал ей хлеба; она ела, наелась, и еще осталось.
RUTH|2|15|И встала, чтобы подбирать. Вооз дал приказ слугам своим, сказав: пусть подбирает она и между снопами, и не обижайте ее;
RUTH|2|16|да и от снопов откидывайте ей и оставляйте, пусть она подбирает, и не браните ее.
RUTH|2|17|Так подбирала она на поле до вечера и вымолотила собранное, и вышло около ефы ячменя.
RUTH|2|18|Взяв это, она пошла в город, и свекровь ее увидела, что она набрала. И вынула [Руфь из пазухи своей] и дала ей то, что оставила, наевшись сама.
RUTH|2|19|И сказала ей свекровь ее: где ты собирала сегодня и где работала? да будет благословен принявший тебя! [Руфь]! объявила свекрови своей, у кого она работала, и сказала: человеку тому, у которого я сегодня работала, имя Вооз.
RUTH|2|20|И сказала Ноеминь снохе своей: благословен он от Господа за то, что не лишил милости своей ни живых, ни мертвых! И сказала ей Ноеминь: человек этот близок к нам; он из наших родственников.
RUTH|2|21|Руфь Моавитянка сказала: он даже сказал мне: будь с моими служанками, доколе не докончат они жатвы моей.
RUTH|2|22|И сказала Ноеминь снохе своей Руфи: хорошо, дочь моя, что ты будешь ходить со служанками его, и не будут оскорблять тебя на другом поле.
RUTH|2|23|Так была она со служанками Воозовыми и подбирала [колосья], доколе не кончилась жатва ячменя и жатва пшеницы, и жила у свекрови своей.
RUTH|3|1|И сказала ей Ноеминь, свекровь ее: дочь моя, не поискать ли тебе пристанища, чтобы тебе хорошо было?
RUTH|3|2|Вот, Вооз, со служанками которого ты была, родственник наш; вот, он в эту ночь веет на гумне ячмень;
RUTH|3|3|умойся, помажься, надень на себя [нарядные] одежды твои и пойди на гумно, но не показывайся ему, доколе не кончит есть и пить;
RUTH|3|4|когда же он ляжет спать, узнай место, где он ляжет; тогда придешь и откроешь у ног его и ляжешь; он скажет тебе, что тебе делать.
RUTH|3|5|[Руфь] сказала ей: сделаю все, что ты сказала мне.
RUTH|3|6|И пошла на гумно и сделала все так, как приказывала ей свекровь ее.
RUTH|3|7|Вооз наелся и напился, и развеселил сердце свое, и пошел [и лег] спать подле скирда. И она пришла тихонько, открыла у ног его и легла.
RUTH|3|8|В полночь он содрогнулся, приподнялся, и вот, у ног его лежит женщина.
RUTH|3|9|И сказал [ей Вооз]: кто ты? Она сказала: я Руфь, раба твоя, простри крыло твое на рабу твою, ибо ты родственник.
RUTH|3|10|[Вооз] сказал: благословенна ты от Господа, дочь моя! это последнее твое доброе дело сделала ты еще лучше прежнего, что ты не пошла искать молодых людей, ни бедных, ни богатых;
RUTH|3|11|итак, дочь моя, не бойся, я сделаю тебе все, что ты сказала; ибо у всех ворот народа моего знают, что ты женщина добродетельная;
RUTH|3|12|хотя и правда, что я родственник, но есть еще родственник ближе меня;
RUTH|3|13|переночуй эту ночь; завтра же, если он примет тебя, то хорошо, пусть примет; а если он не захочет принять тебя, то я приму; жив Господь! Спи до утра.
RUTH|3|14|И спала она у ног его до утра и встала прежде, нежели могли они распознать друг друга. И сказал Вооз: пусть не знают, что женщина приходила на гумно.
RUTH|3|15|И сказал ей: подай верхнюю одежду, которая на тебе, подержи ее. Она держала, и он отмерил [ей] шесть мер ячменя, и положил на нее, и пошел в город.
RUTH|3|16|А [Руфь] пришла к свекрови своей. Та сказала [ей]: что, дочь моя? Она пересказала ей все, что сделал ей человек тот.
RUTH|3|17|И сказала [ей]: эти шесть мер ячменя он дал мне и сказал мне: не ходи к свекрови своей с пустыми руками.
RUTH|3|18|Та сказала: подожди, дочь моя, доколе не узнаешь, чем кончится дело; ибо человек тот не останется в покое, не кончив сегодня дела.
RUTH|4|1|Вооз вышел к воротам и сидел там. И вот, идет мимо родственник, о котором говорил Вооз. И сказал ему [Вооз]: зайди сюда и сядь здесь. Тот зашел и сел.
RUTH|4|2|[Вооз] взял десять человек из старейшин города и сказал: сядьте здесь. И они сели.
RUTH|4|3|И сказал [Вооз] родственнику: Ноеминь, возвратившаяся с полей Моавитских, продает часть поля, принадлежащую брату нашему Елимелеху;
RUTH|4|4|я решился довести до ушей твоих и сказать: купи при сидящих здесь и при старейшинах народа моего; если хочешь выкупить, выкупай; а если не хочешь выкупить, скажи мне, и я буду знать; ибо кроме тебя некому выкупить; а по тебе я. Тот сказал: я выкупаю.
RUTH|4|5|Вооз сказал: когда ты купишь поле у Ноемини, то должен купить и у Руфи Моавитянки, жены умершего, и должен взять ее в замужество, чтобы восстановить имя умершего в уделе его.
RUTH|4|6|И сказал тот родственник: не могу я взять ее себе, чтобы не расстроить своего удела; прими ее ты, ибо я не могу принять.
RUTH|4|7|Прежде такой был [обычай] у Израиля при выкупе и при мене для подтверждения какого–либо дела: один снимал сапог свой и давал другому, и это было свидетельством у Израиля.
RUTH|4|8|И сказал тот родственник Воозу: купи себе. И снял сапог свой.
RUTH|4|9|И сказал Вооз старейшинам и всему народу: вы теперь свидетели тому, что я покупаю у Ноемини все Елимелехово и все Хилеоново и Махлоново;
RUTH|4|10|также и Руфь Моавитянку, жену Махлонову, беру себе в жену, чтоб оставить имя умершего в уделе его, и чтобы не исчезло имя умершего между братьями его и у ворот местопребывания его: вы сегодня свидетели тому.
RUTH|4|11|И сказал весь народ, который при воротах, и старейшины: мы свидетели; да соделает Господь жену, входящую в дом твой, как Рахиль и как Лию, которые обе устроили дом Израилев; приобретай богатство в Ефрафе, и да славится имя твое в Вифлееме;
RUTH|4|12|и да будет дом твой, как дом Фареса, которого родила Фамарь Иуде, от того семени, которое даст тебе Господь от этой молодой женщины.
RUTH|4|13|И взял Вооз Руфь, и она сделалась его женою. И вошел он к ней, и Господь дал ей беременность, и она родила сына.
RUTH|4|14|И говорили женщины Ноемини: благословен Господь, что Он не оставил тебя ныне без наследника! И да будет славно имя его в Израиле!
RUTH|4|15|Он будет тебе отрадою и питателем в старости твоей, ибо его родила сноха твоя, которая любит тебя, которая для тебя лучше семи сыновей.
RUTH|4|16|И взяла Ноеминь дитя сие, и носила его в объятиях своих, и была ему нянькою.
RUTH|4|17|Соседки нарекли ему имя и говорили: "у Ноемини родился сын", и нарекли ему имя: Овид. Он отец Иессея, отца Давидова.
RUTH|4|18|И вот род Фаресов: Фарес родил Есрома;
RUTH|4|19|Есром родил Арама; Арам родил Аминадава;
RUTH|4|20|Аминадав родил Наассона; Наассон родил Салмона;
RUTH|4|21|Салмон родил Вооза; Вооз родил Овида;
RUTH|4|22|Овид родил Иессея; Иессей родил Давида.
