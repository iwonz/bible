ROM|1|1|Paulus servus Christi Iesu, vo catus apostolus, segregatus in evangelium Dei,
ROM|1|2|quod ante promiserat per prophetas suos in Scripturis sanctis
ROM|1|3|de Filio suo, qui factus est ex semine David secundum carnem,
ROM|1|4|qui constitutus est Filius Dei in virtute secundum Spiritum sanctificationis ex resurrectione mortuorum, Iesu Christo Domino nostro,
ROM|1|5|per quem accepimus gratiam et apostolatum ad oboeditionem fidei in omnibus gentibus pro nomine eius,
ROM|1|6|in quibus estis et vos vocati Iesu Christi,
ROM|1|7|omnibus, qui sunt Romae dilectis Dei, vocatis sanctis: gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
ROM|1|8|Primum quidem gratias ago Deo meo per Iesum Christum pro omnibus vobis, quia fides vestra annuntiatur in universo mundo;
ROM|1|9|testis enim mihi est Deus, cui servio in spiritu meo in evangelio Filii eius, quomodo sine intermissione memoriam vestri faciam
ROM|1|10|semper in orationibus meis obsecrans, si quo modo tandem aliquando prosperum iter habeam in voluntate Dei veniendi ad vos.
ROM|1|11|Desidero enim videre vos, ut aliquid impertiar gratiae vobis spiritalis ad confirmandos vos,
ROM|1|12|id est una vobiscum consolari per eam, quae invicem est, fidem vestram atque meam.
ROM|1|13|Nolo autem vos ignorare, fratres, quia saepe proposui venire ad vos et prohibitus sum usque adhuc, ut aliquem fructum habeam et in vobis, sicut et in ceteris gentibus.
ROM|1|14|Graecis ac barbaris, sapientibus et insipientibus debitor sum.
ROM|1|15|Itaque, quod in me est, promptus sum et vobis, qui Romae estis, evangelizare.
ROM|1|16|Non enim erubesco evangelium: virtus enim Dei est in salutem omni credenti, Iudaeo primum et Graeco.
ROM|1|17|Iustitia enim Dei in eo revelatur ex fide in fidem, sicut scriptum est: Iustus autem ex fide vivet ".
ROM|1|18|Revelatur enim ira Dei de caelo super omnem impietatem et iniustitiam hominum, qui veritatem in iniustitia detinent,
ROM|1|19|quia, quod noscibile est Dei, manifestum est in illis; Deus enim illis manifestavit.
ROM|1|20|Invisibilia enim ipsius a creatura mundi per ea, quae facta sunt, intellecta conspiciuntur, sempiterna eius et virtus et divinitas, ut sint inexcusabiles;
ROM|1|21|quia, cum cognovissent Deum, non sicut Deum glorificaverunt aut gratias egerunt, sed evanuerunt in cogitationibus suis, et obscuratum est insipiens cor eorum.
ROM|1|22|Dicentes se esse sapientes, stulti facti sunt,
ROM|1|23|et mutaverunt gloriam incorruptibilis Dei in similitudinem imaginis corruptibilis hominis et volucrum et quadrupedum et serpentium.
ROM|1|24|Propter quod tradidit illos Deus in concupiscentiis cordis eorum in immunditiam, ut ignominia afficiant corpora sua in semetipsis,
ROM|1|25|qui commutaverunt veritatem Dei in mendacio et coluerunt et servierunt creaturae potius quam Creatori, qui est benedictus in saecula. Amen.
ROM|1|26|Propterea tradidit illos Deus in passiones ignominiae. Nam et feminae eorum immutaverunt naturalem usum in eum, qui est contra naturam;
ROM|1|27|similiter et masculi, relicto naturali usu feminae, exarserunt in desideriis suis in invicem, masculi in masculos turpitudinem operantes et mercedem, quam oportuit, erroris sui in semetipsis recipientes.
ROM|1|28|Et sicut non probaverunt Deum habere in notitia, tradidit eos Deus in reprobum sensum, ut faciant, quae non conveniunt,
ROM|1|29|repletos omni iniquitate, malitia, avaritia, nequitia, plenos invidia, homicidio, contentione, dolo, malignitate, susurrones,
ROM|1|30|detractores, Deo odibiles, contumeliosos, superbos, elatos, inventores malorum, parentibus non oboedientes,
ROM|1|31|insipientes, incompositos, sine affectione, sine misericordia.
ROM|1|32|Qui cum iudicium Dei cognovissent, quoniam qui talia agunt, digni sunt morte, non solum ea faciunt, sed et consentiunt facientibus.
ROM|2|1|Propter quod inexcusabilis es, o homo omnis, qui iudicas. In quo enim iudicas alterum, teipsum condemnas; eadem enim agis, qui iudicas.
ROM|2|2|Scimus enim quoniam iudicium Dei est secundum veritatem in eos, qui talia agunt.
ROM|2|3|Existimas autem hoc, o homo, qui iudicas eos, qui talia agunt, et facis ea, quia tu effugies iudicium Dei?
ROM|2|4|An divitias benignitatis eius et patientiae et longanimitatis contemnis, ignorans quoniam benignitas Dei ad paenitentiam te adducit?
ROM|2|5|Secundum duritiam autem tuam et impaenitens cor thesaurizas tibi iram in die irae et revelationis iusti iudicii Dei,
ROM|2|6|qui reddet unicuique secundum opera eius:
ROM|2|7|his quidem, qui secundum patientiam boni operis gloriam et honorem et incorruptionem quaerunt, vitam aeternam;
ROM|2|8|his autem, qui ex contentione et non oboediunt veritati, oboediunt autem iniquitati, ira et indignatio.
ROM|2|9|Tribulatio et angustia in omnem animam hominis operantis malum, Iudaei primum et Graeci;
ROM|2|10|gloria autem et honor et pax omni operanti bonum, Iudaeo primum et Graeco.
ROM|2|11|Non est enim personarum acceptio apud Deum!
ROM|2|12|Quicumque enim sine lege peccaverunt, sine lege et peribunt; et, quicumque in lege peccaverunt, per legem iudicabuntur.
ROM|2|13|Non enim auditores legis iusti sunt apud Deum, sed factores legis iustificabuntur.
ROM|2|14|Cum enim gentes, quae legem non habent, naturaliter, quae legis sunt, faciunt, eiusmodi legem non habentes ipsi sibi sunt lex;
ROM|2|15|qui ostendunt opus legis scriptum in cordibus suis, testimonium simul reddente illis conscientia ipsorum, et inter se invicem cogitationibus accusantibus aut etiam defendentibus,
ROM|2|16|in die, cum iudicabit Deus occulta hominum secundum evangelium meum per Christum Iesum.
ROM|2|17|Si autem tu Iudaeus cognominaris et requiescis in lege et gloriaris in Deo,
ROM|2|18|et nosti Voluntatem et discernis potiora instructus per legem,
ROM|2|19|et confidis teipsum ducem esse caecorum, lumen eorum, qui in tenebris sunt,
ROM|2|20|eruditorem insipientium, magistrum infantium, habentem formam scientiae et veritatis in lege.
ROM|2|21|Qui ergo alium doces, teipsum non doces? Qui praedicas non furandum, furaris?
ROM|2|22|Qui dicis non moechandum, moecharis? Qui abominaris idola, templa spolias?
ROM|2|23|Qui in lege gloriaris, per praevaricationem legis Deum inhonoras?
ROM|2|24|" Nomen enim Dei propter vos blasphematur inter gentes ", sicut scriptum est.
ROM|2|25|Circumcisio quidem prodest, si legem observes; si autem praevaricator legis sis, circumcisio tua praeputium facta est.
ROM|2|26|Si igitur praeputium iustitias legis custodiat, nonne praeputium illius in circumcisionem reputabitur?
ROM|2|27|Et iudicabit, quod ex natura est praeputium legem consummans, te, qui per litteram et circumcisionem praevaricator legis es.
ROM|2|28|Non enim qui manifesto Iudaeus est, neque quae manifesto in carne circumcisio,
ROM|2|29|sed qui in abscondito Iudaeus est, et circumcisio cordis in spiritu non littera, cuius laus non ex hominibus sed ex Deo est.
ROM|3|1|Quid ergo amplius est Iudaeo, aut quae utilitas circumcisionis?
ROM|3|2|Multum per omnem modum. Primum quidem, quia credita sunt illis eloquia Dei.
ROM|3|3|Quid enim, si quidam non crediderunt? Numquid incredulitas illorum fidem Dei evacuabit?
ROM|3|4|Absit! Exstet autem Deus verax, omnis autem homo mendax, sicut scriptum est: " Ut iustificeris in sermonibus tuis et vincas cum iudicaris ".
ROM|3|5|Si autem iniustitia nostra iustitiam Dei commendat, quid dicemus? Numquid iniustus Deus, qui infert iram? Secundum hominem dico.
ROM|3|6|Absit! Alioquin quomodo iudicabit Deus mundum?
ROM|3|7|Si enim veritas Dei in meo mendacio abundavit in gloriam ipsius, quid adhuc et ego tamquam peccator iudicor?
ROM|3|8|Et non, sicut blasphemamur, et sicut aiunt quidam nos dicere: " Faciamus mala, ut veniant bona "? Quorum damnatio iusta est.
ROM|3|9|Quid igitur? Praecellimus eos? Nequaquam! Antea enim causati sumus Iudaeos et Graecos omnes sub peccato esse,
ROM|3|10|sicut scriptum est: Non est iustus quisquam,
ROM|3|11|non est intellegens, non est requirens Deum.
ROM|3|12|Omnes declinaverunt, simul inutiles facti sunt;non est qui faciat bonum, non est usque ad unum.
ROM|3|13|Sepulcrum patens est guttur eorum,linguis suis dolose agebant,venenum aspidum sub labiis eorum,
ROM|3|14|quorum os maledictione et amaritudine plenum est;
ROM|3|15|veloces pedes eorum ad effundendum sanguinem,
ROM|3|16|contritio et infelicitas in viis eorum,
ROM|3|17|et viam pacis non cognoverunt.
ROM|3|18|Non est timor Dei ante oculos eorum ".
ROM|3|19|Scimus autem quoniam, quaecumque lex loquitur, his, qui in lege sunt, loquitur, ut omne os obstruatur, et obnoxius fiat omnis mundus Deo;
ROM|3|20|quia ex operibus legis non iustificabitur omnis caro coram illo, per legem enim cognitio peccati.
ROM|3|21|Nunc autem sine lege iustitia Dei manifestata est, testificata a Lege et Prophetis,
ROM|3|22|iustitia autem Dei per fidem Iesu Christi, in omnes, qui credunt. Non enim est distinctio:
ROM|3|23|omnes enim peccaverunt et egent gloria Dei,
ROM|3|24|iustificati gratis per gratiam ipsius per redemptionem, quae est in Christo Iesu;
ROM|3|25|quem proposuit Deus propitiatorium per fidem in sanguine ipsius ad ostensionem iustitiae suae, cum praetermisisset praecedentia delicta
ROM|3|26|in sustentatione Dei, ad ostensionem iustitiae eius in hoc tempore, ut sit ipse iustus et iustificans eum, qui ex fide est Iesu.
ROM|3|27|Ubi est ergo gloriatio? Exclusa est. Per quam legem? Operum? Non, sed per legem fidei.
ROM|3|28|Arbitramur enim iustificari hominem per fidem sine operibus legis.
ROM|3|29|An Iudaeorum Deus tantum? Nonne et gentium? Immo et gentium,
ROM|3|30|quoniam quidem unus Deus, qui iustificabit circumcisionem ex fide et praeputium per fidem.
ROM|3|31|Legem ergo destruimus per fidem? Absit, sed legem statuimus.
ROM|4|1|Quid ergo dicemus invenisse Abraham progenitorem no strum secundum carnem?
ROM|4|2|Si enim Abraham ex operibus iustificatus est, habet gloriam sed non apud Deum.
ROM|4|3|Quid enim Scriptura dicit? " Credidit autem Abraham Deo, et reputatum est illi ad iustitiam ".
ROM|4|4|Ei autem, qui operatur, merces non reputatur secundum gratiam sed secundum debitum;
ROM|4|5|ei vero, qui non operatur, sed credit in eum, qui iustificat impium, reputatur fides eius ad iustitiam,
ROM|4|6|sicut et David dicit beatitudinem hominis, cui Deus reputat iustitiam sine operibus:
ROM|4|7|" Beati, quorum remissae sunt iniquitates,et quorum tecta sunt peccata.
ROM|4|8|Beatus vir, cui non imputabit Dominus peccatum ".
ROM|4|9|Beatitudo ergo haec in circumcisione an etiam in praeputio? Dicimus enim: " Reputata est Abrahae fides ad iustitiam ".
ROM|4|10|Quomodo ergo reputata est? In circumcisione an in praeputio? Non in circumcisione sed in praeputio:
ROM|4|11|et signum accepit circumcisionis, signaculum iustitiae fidei, quae fuit in praeputio, ut esset pater omnium credentium per praeputium, ut reputetur illis iustitia,
ROM|4|12|et pater circumcisionis his non tantum, qui ex circumcisione sunt, sed et qui sectantur vestigia eius, quae fuit in praeputio, fidei patris nostri Abrahae.
ROM|4|13|Non enim per legem promissio Abrahae aut semini eius, ut heres esset mundi, sed per iustitiam fidei;
ROM|4|14|si enim qui ex lege heredes sunt, exinanita est fides, et abolita est promissio.
ROM|4|15|Lex enim iram operatur; ubi autem non est lex, nec praevaricatio.
ROM|4|16|Ideo ex fide, ut secundum gratiam, ut firma sit promissio omni semini, non ei, qui ex lege est solum, sed et ei, qui ex fide est Abrahae - qui est pater omnium nostrum,
ROM|4|17|sicut scriptum est: " Patrem multarum gentium posui te " C, ante Deum, cui credidit, qui vivificat mortuos et vocat ea, quae non sunt, quasi sint;
ROM|4|18|qui contra spem in spe credidit, ut fieret pater multarum gentium, secundum quod dictum est: " Sic erit semen tuum ".
ROM|4|19|Et non infirmatus fide consideravit corpus suum iam emortuum, cum fere centum annorum esset, et emortuam vulvam Sarae;
ROM|4|20|in repromissione autem Dei non haesitavit diffidentia, sed confortatus est fide, dans gloriam Deo,
ROM|4|21|et plenissime sciens quia, quod promisit, potens est et facere.
ROM|4|22|Ideo et reputatum est illi ad iustitiam.
ROM|4|23|Non est autem scriptum tantum propter ipsum: reputatum est illi,
ROM|4|24|sed et propter nos, quibus reputabitur, credentibus in eum, qui suscitavit Iesum Dominum nostrum a mortuis,
ROM|4|25|qui traditus est propter delicta nostra et suscitatus est propter iustificationem nostram.
ROM|5|1|Iustificati igitur ex fide, pacem habemus ad Deum per Domi num nostrum Iesum Christum,
ROM|5|2|per quem et accessum habemus fide in gratiam istam, in qua stamus et gloriamur in spe gloriae Dei.
ROM|5|3|Non solum autem, sed et gloriamur in tribulationibus, scientes quod tribulatio patientiam operatur,
ROM|5|4|patientia autem probationem, probatio vero spem;
ROM|5|5|spes autem non confundit, quia caritas Dei diffusa est in cordibus nostris per Spiritum Sanctum, qui datus est nobis.
ROM|5|6|Adhuc enim Christus, cum adhuc infirmi essemus, secundum tempus pro impiis mortuus est.
ROM|5|7|Vix enim pro iusto quis moritur; nam pro bono forsitan quis et audeat mori.
ROM|5|8|Commendat autem suam caritatem Deus in nos, quoniam, cum adhuc peccatores essemus, Christus pro nobis mortuus est.
ROM|5|9|Multo igitur magis iustificati nunc in sanguine ipsius, salvi erimus ab ira per ipsum!
ROM|5|10|Si enim, cum inimici essemus, reconciliati sumus Deo per mortem Filii eius, multo magis reconciliati salvi erimus in vita ipsius;
ROM|5|11|non solum autem, sed et gloriamur in Deo per Dominum nostrum Iesum Christum, per quem nunc reconciliationem accepimus.
ROM|5|12|Propterea, sicut per unum hominem peccatum in hunc mundum intravit, et per peccatum mors, et ita in omnes homines mors pertransiit, eo quod omnes peccaverunt.
ROM|5|13|Usque ad legem enim peccatum erat in mundo; peccatum autem non imputatur, cum lex non est,
ROM|5|14|sed regnavit mors ab Adam usque ad Moysen etiam in eos, qui non peccaverunt in similitudine praevaricationis Adae, qui est figura futuri.
ROM|5|15|Sed non sicut delictum, ita et donum; si enim unius delicto multi mortui sunt, multo magis gratia Dei et donum in gratia unius hominis Iesu Christi in multos abundavit.
ROM|5|16|Et non sicut per unum, qui peccavit, ita et donum; nam iudicium ex uno in condemnationem, gratia autem ex multis delictis in iustificationem.
ROM|5|17|Si enim unius delicto mors regnavit per unum, multo magis, qui abundantiam gratiae et donationis iustitiae accipiunt, in vita regnabunt per unum Iesum Christum.
ROM|5|18|Igitur sicut per unius delictum in omnes homines in condemnationem, sic et per unius iustitiam in omnes homines in iustificationem vitae;
ROM|5|19|sicut enim per inoboedientiam unius hominis peccatores constituti sunt multi, ita et per unius oboeditionem iusti constituentur multi.
ROM|5|20|Lex autem subintravit, ut abundaret delictum; ubi autem abundavit peccatum, superabundavit gratia,
ROM|5|21|ut sicut regnavit peccatum in morte, ita et gratia regnet per iustitiam in vitam aeternam per Iesum Christum Dominum nostrum.
ROM|6|1|Quid ergo dicemus? Perma nebimus in peccato, ut gratia abundet?
ROM|6|2|Absit! Qui enim mortui sumus peccato, quomodo adhuc vivemus in illo?
ROM|6|3|An ignoratis quia, quicumque baptizati sumus in Christum Iesum, in mortem ipsius baptizati sumus?
ROM|6|4|Consepulti ergo sumus cum illo per baptismum in mortem, ut quemadmodum suscitatus est Christus a mortuis per gloriam Patris, ita et nos in novitate vitae ambulemus.
ROM|6|5|Si enim complantati facti sumus similitudini mortis eius, sed et resurrectionis erimus;
ROM|6|6|hoc scientes quia vetus homo noster simul crucifixus est, ut destruatur corpus peccati, ut ultra non serviamus peccato.
ROM|6|7|Qui enim mortuus est, iustificatus est a peccato.
ROM|6|8|Si autem mortui sumus cum Christo, credimus quia simul etiam vivemus cum eo;
ROM|6|9|scientes quod Christus suscitatus ex mortuis iam non moritur, mors illi ultra non dominatur.
ROM|6|10|Quod enim mortuus est, peccato mortuus est semel; quod autem vivit, vivit Deo.
ROM|6|11|Ita et vos existimate vos mortuos quidem esse peccato, viventes autem Deo in Christo Iesu.
ROM|6|12|Non ergo regnet peccatum in vestro mortali corpore, ut oboediatis concupiscentiis eius,
ROM|6|13|neque exhibeatis membra vestra arma iniustitiae peccato, sed exhibete vos Deo tamquam ex mortuis viventes et membra vestra arma iustitiae Deo.
ROM|6|14|Peccatum enim vobis non dominabitur; non enim sub lege estis sed sub gratia.
ROM|6|15|Quid ergo? Peccabimus, quoniam non sumus sub lege sed sub gratia? Absit!
ROM|6|16|Nescitis quoniam, cui exhibetis vos servos ad oboedientiam, servi estis eius, cui oboeditis, sive peccati ad mortem, sive oboeditionis ad iustitiam?
ROM|6|17|Gratias autem Deo quod fuistis servi peccati, oboedistis autem ex corde in eam formam doctrinae, in quam traditi estis,
ROM|6|18|liberati autem a peccato servi facti estis iustitiae.
ROM|6|19|Humanum dico propter infirmitatem carnis vestrae. Sicut enim exhibuistis membra vestra servientia immunditiae et iniquitati ad iniquitatem, ita nunc exhibete membra vestra servientia iustitiae ad sanctificationem.
ROM|6|20|Cum enim servi essetis peccati, liberi eratis iustitiae.
ROM|6|21|Quem ergo fructum habebatis tunc, in quibus nunc erubescitis? Nam finis illorum mors!
ROM|6|22|Nunc vero liberati a peccato, servi autem facti Deo, habetis fructum vestrum in sanctificationem, finem vero vitam aeternam!
ROM|6|23|Stipendia enim peccati mors, donum autem Dei vita aeterna in Christo Iesu Domino nostro.
ROM|7|1|An ignoratis, fratres - scienti bus enim legem loquor - quia lex in homine dominatur, quanto tempore vivit?
ROM|7|2|Nam quae sub viro est mulier, viventi viro alligata est lege; si autem mortuus fuerit vir, soluta est a lege viri.
ROM|7|3|Igitur, vivente viro, vocabitur adultera, si fuerit alterius viri; si autem mortuus fuerit vir, libera est a lege, ut non sit adultera, si fuerit alterius viri.
ROM|7|4|Itaque, fratres mei, et vos mortificati estis legi per corpus Christi, ut sitis alterius, eius qui ex mortuis suscitatus est, ut fructificaremus Deo.
ROM|7|5|Cum enim essemus in carne, passiones peccatorum, quae per legem sunt, operabantur in membris nostris, ut fructificarent morti;
ROM|7|6|nunc autem soluti sumus a lege, mortui ei, in qua detinebamur, ita ut serviamus in novitate Spiritus et non in vetustate litterae.
ROM|7|7|Quid ergo dicemus? Lex peccatum est? Absit! Sed peccatum non cognovi, nisi per legem; nam concupiscentiam nescirem, nisi lex diceret: " Non concupisces ".
ROM|7|8|Occasione autem accepta, peccatum per mandatum operatum est in me omnem concupiscentiam; sine lege enim peccatum mortuum erat.
ROM|7|9|Ego autem vivebam sine lege aliquando; sed, cum venisset mandatum, peccatum revixit,
ROM|7|10|ego autem mortuus sum; et inventum est mihi mandatum, quod erat ad vitam, hoc esse ad mortem;
ROM|7|11|nam peccatum, occasione accepta, per mandatum seduxit me et per illud occidit.
ROM|7|12|Itaque lex quidem sancta, et mandatum sanctum et iustum et bonum.
ROM|7|13|Quod ergo bonum est, mihi factum est mors? Absit! Sed peccatum, ut appareat peccatum, per bonum mihi operatum est mortem; ut fiat supra modum peccans peccatum per mandatum.
ROM|7|14|Scimus enim quod lex spiritalis est; ego autem carnalis sum, venumdatus sub peccato.
ROM|7|15|Quod enim operor, non intellego; non enim, quod volo, hoc ago, sed quod odi, illud facio.
ROM|7|16|Si autem, quod nolo, illud facio, consentio legi quoniam bona.
ROM|7|17|Nunc autem iam non ego operor illud, sed, quod habitat in me, peccatum.
ROM|7|18|Scio enim quia non habitat in me, hoc est in carne mea, bonum; nam velle adiacet mihi, operari autem bonum, non!
ROM|7|19|Non enim, quod volo bonum, facio, sed, quod nolo malum, hoc ago.
ROM|7|20|Si autem, quod nolo, illud facio, iam non ego operor illud, sed, quod habitat in me, peccatum.
ROM|7|21|Invenio igitur hanc legem volenti mihi facere bonum, quoniam mihi malum adiacet.
ROM|7|22|Condelector enim legi Dei secundum interiorem hominem;
ROM|7|23|video autem aliam legem in membris meis repugnantem legi mentis meae et captivantem me in lege peccati, quae est in membris meis.
ROM|7|24|Infelix ego homo! Quis me liberabit de corpore mortis huius?
ROM|7|25|Gratias autem Deo per Iesum Christum Dominum nostrum! Igitur ego ipse mente servio legi Dei, carne autem legi peccati.
ROM|8|1|Nihil ergo nunc damnationis est his, qui sunt in Christo Iesu;
ROM|8|2|lex enim Spiritus vitae in Christo Iesu liberavit te a lege peccati et mortis.
ROM|8|3|Nam, quod impossibile erat legi, in quo infirmabatur per carnem, Deus Filium suum mittens in similitudine carnis peccati et pro peccato, damnavit peccatum in carne,
ROM|8|4|ut iustitia legis impleretur in nobis, qui non secundum carnem ambulamus sed secundum Spiritum.
ROM|8|5|Qui enim secundum carnem sunt, quae carnis sunt, sapiunt; qui vero secundum Spiritum, quae sunt Spiritus.
ROM|8|6|Nam sapientia carnis mors, sapientia autem Spiritus vita et pax;
ROM|8|7|quoniam sapientia carnis inimicitia est in Deum, legi enim Dei non subicitur nec enim potest.
ROM|8|8|Qui autem in carne sunt, Deo placere non possunt.
ROM|8|9|Vos autem in carne non estis sed in Spiritu, si tamen Spiritus Dei habitat in vobis. Si quis autem Spiritum Christi non habet, hic non est eius.
ROM|8|10|Si autem Christus in vobis est, corpus quidem mortuum est propter peccatum, Spiritus vero vita propter iustitiam.
ROM|8|11|Quod si Spiritus eius, qui suscitavit Iesum a mortuis, habitat in vobis, qui suscitavit Christum a mortuis vivificabit et mortalia corpora vestra per inhabitantem Spiritum suum in vobis.
ROM|8|12|Ergo, fratres, debitores sumus non carni, ut secundum carnem vivamus.
ROM|8|13|Si enim secundum carnem vixeritis, moriemini; si autem Spiritu opera corporis mortificatis, vivetis.
ROM|8|14|Quicumque enim Spiritu Dei aguntur, hi filii Dei sunt.
ROM|8|15|Non enim accepistis spiritum servitutis iterum in timorem, sed accepistis Spiritum adoptionis filiorum, in quo clamamus: " Abba, Pater!.
ROM|8|16|Ipse Spiritus testimonium reddit una cum spiritu nostro, quod sumus filii Dei.
ROM|8|17|Si autem filii, et heredes: heredes quidem Dei, coheredes autem Christi, si tamen compatimur, ut et conglorificemur.
ROM|8|18|Existimo enim quod non sunt condignae passiones huius temporis ad futuram gloriam, quae revelanda est in nobis.
ROM|8|19|Nam exspectatio creaturae revelationem filiorum Dei exspectat;
ROM|8|20|vanitati enim creatura subiecta est, non volens sed propter eum, qui subiecit, in spem,
ROM|8|21|quia et ipsa creatura liberabitur a servitute corruptionis in libertatem gloriae filiorum Dei.
ROM|8|22|Scimus enim quod omnis creatura congemiscit et comparturit usque adhuc;
ROM|8|23|non solum autem, sed et nos ipsi primitias Spiritus habentes, et ipsi intra nos gemimus adoptionem filiorum exspectantes, redemptionem corporis nostri.
ROM|8|24|Spe enim salvi facti sumus; spes autem, quae videtur, non est spes; nam, quod videt, quis sperat?
ROM|8|25|Si autem, quod non videmus, speramus, per patientiam exspectamus.
ROM|8|26|Similiter autem et Spiritus adiuvat infirmitatem nostram; nam quid oremus, sicut oportet, nescimus, sed ipse Spiritus interpellat gemitibus inenarrabilibus;
ROM|8|27|qui autem scrutatur corda, scit quid desideret Spiritus, quia secundum Deum postulat pro sanctis.
ROM|8|28|Scimus autem quoniam diligentibus Deum omnia cooperantur in bonum, his, qui secundum propositum vocati sunt.
ROM|8|29|Nam, quos praescivit, et praedestinavit conformes fieri imaginis Filii eius, ut sit ipse primogenitus in multis fratribus;
ROM|8|30|quos autem praedestinavit, hos et vocavit; et quos vocavit, hos et iustificavit; quos autem iustificavit, illos et glorificavit.
ROM|8|31|Quid ergo dicemus ad haec? Si Deus pro nobis, quis contra nos?
ROM|8|32|Qui Filio suo non pepercit, sed pro nobis omnibus tradidit illum, quomodo non etiam cum illo omnia nobis donabit?
ROM|8|33|Quis accusabit adversus electos Dei? Deus, qui iustificat?
ROM|8|34|Quis est qui condemnet? Christus Iesus, qui mortuus est, immo qui suscitatus est, qui et est ad dexteram Dei, qui etiam interpellat pro nobis?
ROM|8|35|Quis nos separabit a caritate Christi? Tribulatio an angustia an persecutio an fames an nuditas an periculum an gladius?
ROM|8|36|Sicut scriptum est: Propter te mortificamur tota die,aestimati sumus ut oves occisionis ".
ROM|8|37|Sed in his omnibus supervincimus per eum, qui dilexit nos.
ROM|8|38|Certus sum enim quia neque mors neque vita neque angeli neque principatus neque instantia neque futura neque virtutes
ROM|8|39|neque altitudo neque profundum neque alia quaelibet creatura poterit nos separare a caritate Dei, quae est in Christo Iesu Domino nostro.
ROM|9|1|Veritatem dico in Christo, non mentior, testimonium mihi per hibente conscientia mea in Spiritu Sancto,
ROM|9|2|quoniam tristitia est mihi magna, et continuus dolor cordi meo.
ROM|9|3|Optarem enim ipse ego anathema esse a Christo pro fratribus meis, cognatis meis secundum carnem,
ROM|9|4|qui sunt Israelitae, quorum adoptio est filiorum et gloria et testamenta et legislatio et cultus et promissiones,
ROM|9|5|quorum sunt patres, et ex quibus Christus secundum carnem: qui est super omnia Deus benedictus in saecula. Amen.
ROM|9|6|Non autem quod exciderit verbum Dei. Non enim omnes, qui ex Israel, hi sunt Israel;
ROM|9|7|neque quia semen sunt Abrahae, omnes filii, sed: " In Isaac vocabitur tibi semen ".
ROM|9|8|Id est, non qui filii carnis, hi filii Dei, sed qui filii sunt promissionis, aestimantur semen;
ROM|9|9|promissionis enim verbum hoc est: " Secundum hoc tempus veniam, et erit Sarae filius ".
ROM|9|10|Non solum autem, sed et Rebecca ex uno concubitum habens, Isaac patre nostro;
ROM|9|11|cum enim nondum nati fuissent aut aliquid egissent bonum aut malum, ut secundum electionem propositum Dei maneret,
ROM|9|12|non ex operibus sed ex vocante dictum est ei: " Maior serviet minori ";
ROM|9|13|sicut scriptum est: " Iacob dilexi, Esau autem odio habui ".
ROM|9|14|Quid ergo dicemus? Numquid iniustitia apud Deum? Absit!
ROM|9|15|Moysi enim dicit: " Miserebor, cuius misereor, et misericordiam praestabo, cui misericordiam praesto ".
ROM|9|16|Igitur non volentis neque currentis sed miserentis Dei.
ROM|9|17|Dicit enim Scriptura pharaoni: " In hoc ipsum excitavi te, ut ostendam in te virtutem meam, et ut annuntietur nomen meum in universa terra ".
ROM|9|18|Ergo, cuius vult, miseretur et, quem vult, indurat.
ROM|9|19|Dices itaque mihi: " Quid ergo adhuc queritur? Voluntati enim eius quis restitit? ".
ROM|9|20|O homo, sed tu quis es, qui respondeas Deo? Numquid dicet figmentum ei, qui se finxit: " Quid me fecisti sic? ".
ROM|9|21|An non habet potestatem figulus luti ex eadem massa facere aliud quidem vas in honorem, aliud vero in ignominiam?
ROM|9|22|Quod si volens Deus ostendere iram et notam facere potentiam suam, sustinuit in multa patientia vasa irae aptata in interitum;
ROM|9|23|et ut ostenderet divitias gloriae suae in vasa misericordiae, quae praeparavit in gloriam,
ROM|9|24|quos et vocavit nos non solum ex Iudaeis sed etiam ex gentibus?
ROM|9|25|Sicut et in Osee dicit: Vocabo Non plebem meam Plebem meamet Non dilectam Dilectam.
ROM|9|26|Et erit: in loco, ubi dictum est eis:Non plebs mea vos",ibi vocabuntur Filii Dei vivi ".
ROM|9|27|Isaias autem clamat pro Israel: " Si fuerit numerus filiorum Israel tamquam arena maris, reliquiae salvae fient.
ROM|9|28|Verbum enim consummans et brevians faciet Dominus super terram ".
ROM|9|29|Et sicut praedixit Isaias: Nisi Dominus Sabaoth reliquisset nobis semen,sicut Sodoma facti essemuset sicut Gomorra similes fuissemus ".
ROM|9|30|Quid ergo dicemus? Quod gentes, quae non sectabantur iustitiam, apprehenderunt iustitiam, iustitiam autem, quae ex fide est;
ROM|9|31|Israel vero sectans legem iustitiae in legem non pervenit.
ROM|9|32|Quare? Quia non ex fide sed quasi ex operibus; offenderunt in lapidem offensionis,
ROM|9|33|sicut scriptum est: Ecce pono in Sion lapidem offensionis et petram scandali;et, qui credit in eo, non confundetur ".
ROM|10|1|Fratres, voluntas quidem cordis mei et obsecratio ad Deum pro illis in salutem.
ROM|10|2|Testimonium enim perhibeo illis quod aemulationem Dei habent sed non secundum scientiam;
ROM|10|3|ignorantes enim Dei iustitiam et suam iustitiam quaerentes statuere, iustitiae Dei non sunt subiecti;
ROM|10|4|finis enim legis Christus ad iustitiam omni credenti.
ROM|10|5|Moyses enim scribit de iustitia, quae ex lege est: " Qui fecerit homo, vivet in eis ".
ROM|10|6|Quae autem ex fide est iustitia, sic dicit: " Ne dixeris in corde tuo: Quis ascendet in caelum?", id est Christum deducere;
ROM|10|7|aut: " Quis descendet in abyssum? ", hoc est Christum ex mortuis revocare.
ROM|10|8|Sed quid dicit? " Prope te est verbum, in ore tuo et in corde tuo "; hoc est verbum fidei, quod praedicamus.
ROM|10|9|Quia si confitearis in ore tuo: " Dominum Iesum! ", et in corde tuo credideris quod Deus illum excitavit ex mortuis, salvus eris.
ROM|10|10|Corde enim creditur ad iustitiam, ore autem confessio fit in salutem.
ROM|10|11|Dicit enim Scriptura: Omnis, qui credit in illo, non confundetur ".
ROM|10|12|Non enim est distinctio Iudaei et Graeci, nam idem Dominus omnium, dives in omnes, qui invocant illum:
ROM|10|13|Omnis enim, quicumque invocaverit nomen Domini, salvus erit.
ROM|10|14|Quomodo ergo invocabunt, in quem non crediderunt? Aut quomodo credent ei, quem non audierunt? Quomodo autem audient sine praedicante?
ROM|10|15|Quomodo vero praedicabunt nisi mittantur? Sicut scriptum est: Quam speciosi pedes evangelizantium bona ".
ROM|10|16|Sed non omnes oboedierunt evangelio; Isaias enim dicit: Domine, quis credidit auditui nostro? ".
ROM|10|17|Ergo fides ex auditu, auditus autem per verbum Christi.
ROM|10|18|Sed dico: Numquid non audierunt? Quin immo,in omnem terram exiit sonus eorum,et in fines orbis terrae verba eorum.
ROM|10|19|Sed dico: Numquid Israel non cognovit? Primus Moyses dicit: Ego ad aemulationem vos adducam per Non gentem:per gentem insipientem ad iram vos provocabo ".
ROM|10|20|Isaias autem audet et dicit: " Inventus sum in non quaerentibus me; palam apparui his, qui me non interrogabant ".
ROM|10|21|Ad Israel autem dicit: " Tota die expandi manus meas ad populum non credentem et contradicentem ".
ROM|11|1|Dico ergo: Numquid repulit Deus populum suum? Absit! Nam et ego Israelita sum, ex semine Abraham, tribu Beniamin.
ROM|11|2|Non reppulit Deus plebem suam, quam praescivit. An nescitis in Elia quid dicit Scriptura? Quemadmodum interpellat Deum adversus Israel:
ROM|11|3|" Domine, prophetas tuos occiderunt, altaria tua suffoderunt, et ego relictus sum solus, et quaerunt animam meam ".
ROM|11|4|Sed quid dicit illi responsum divinum? Reliqui mihi septem milia virorum, qui non curvaverunt genu Baal ".
ROM|11|5|Sic ergo et in hoc tempore reliquiae secundum electionem gratiae factae sunt.
ROM|11|6|Si autem gratia, iam non ex operibus, alioquin gratia iam non est gratia.
ROM|11|7|Quid ergo? Quod quaerit Israel, hoc non est consecutus, electio autem consecuta est; ceteri vero excaecati sunt,
ROM|11|8|sicut scriptum est: Dedit illis Deus spiritum soporis,oculos, ut non videant,et aures, ut non audiant,usque in hodiernum diem ".
ROM|11|9|Et David dicit: Fiat mensa eorum in laqueum et in captionemet in scandalum et in retributionem illis.
ROM|11|10|Obscurentur oculi eorum, ne videant,et dorsum illorum semper incurva! ".
ROM|11|11|Dico ergo: Numquid sic offenderunt, ut caderent? Absit! Sed illorum casu salus gentibus, ut illi ad aemulationem adducantur.
ROM|11|12|Quod si casus illorum divitiae sunt mundi, et deminutio eorum divitiae gentium, quanto magis plenitudo eorum!
ROM|11|13|Vobis autem dico gentibus: Quantum quidem ego sum gentium apostolus, ministerium meum honorifico,
ROM|11|14|si quo modo ad aemulandum provocem carnem meam et salvos faciam aliquos ex illis.
ROM|11|15|Si enim amissio eorum reconciliatio est mundi, quae assumptio, nisi vita ex mortuis?
ROM|11|16|Quod si primitiae sanctae sunt, et massa; et si radix sancta, et rami.
ROM|11|17|Quod si aliqui ex ramis fracti sunt, tu autem, cum oleaster esses, insertus es in illis et consocius radicis pinguedinis olivae factus es,
ROM|11|18|noli gloriari adversus ramos; quod si gloriaris, non tu radicem portas, sed radix te.
ROM|11|19|Dices ergo: " Fracti sunt rami, ut ego inserar ".
ROM|11|20|Bene; incredulitate fracti sunt, tu autem fide stas. Noli altum sapere, sed time:
ROM|11|21|si enim Deus naturalibus ramis non pepercit, ne forte nec tibi parcat.
ROM|11|22|Vide ergo bonitatem et severitatem Dei: in eos quidem, qui ceciderunt, severitatem; in te autem bonitatem Dei, si permanseris in bonitate, alioquin et tu excideris.
ROM|11|23|Sed et illi, si non permanserint in incredulitate, inserentur; potens est enim Deus iterum inserere illos!
ROM|11|24|Nam si tu ex naturali excisus es oleastro et contra naturam insertus es in bonam olivam, quanto magis hi, qui secundum naturam sunt, inserentur suae olivae.
ROM|11|25|Nolo enim vos ignorare, fratres, mysterium hoc, ut non sitis vobis ipsis sapientes, quia caecitas ex parte contigit in Israel, donec plenitudo gentium intraret,
ROM|11|26|et sic omnis Israel salvus fiet, sicut scriptum est: Veniet ex Sion, qui eripiat,avertet impietates ab Iacob;
ROM|11|27|et hoc illis a me testamentum,cum abstulero peccata eorum ".
ROM|11|28|Secundum evangelium quidem inimici propter vos, secundum electionem autem carissimi propter patres;
ROM|11|29|sine paenitentia enim sunt dona et vocatio Dei!
ROM|11|30|Sicut enim aliquando vos non credidistis Deo, nunc autem misericordiam consecuti estis propter illorum incredulitatem,
ROM|11|31|ita et isti nunc non crediderunt propter vestram misericordiam, ut et ipsi nunc misericordiam consequantur.
ROM|11|32|Conclusit enim Deus omnes in incredulitatem, ut omnium misereatur!
ROM|11|33|O altitudo divitiarum et sapientiae et scientiae Dei! Quam incomprehensibilia sunt iudicia eius, et investigabiles viae eius!
ROM|11|34|Quis enim cognovit sensum Domini?Aut quis consiliarius eius fuit?
ROM|11|35|Aut quis prior dedit illi,et retribuetur ei?
ROM|11|36|Quoniam ex ipso et per ipsum et in ipsum omnia. Ipsi gloria in saecula. Amen.
ROM|12|1|Obsecro itaque vos, fratres, per misericordiam Dei, ut exhibeatis corpora vestra hostiam viventem, sanctam, Deo placentem, rationabile obsequium vestrum;
ROM|12|2|et nolite conformari huic saeculo, sed transformamini renovatione mentis, ut probetis quid sit voluntas Dei, quid bonum et bene placens et perfectum.
ROM|12|3|Dico enim per gratiam, quae data est mihi, omnibus, qui sunt inter vos, non altius sapere quam oportet sapere, sed sapere ad sobrietatem, unicuique sicut Deus divisit mensuram fidei.
ROM|12|4|Sicut enim in uno corpore multa membra habemus, omnia autem membra non eundem actum habent,
ROM|12|5|ita multi unum corpus sumus in Christo, singuli autem alter alterius membra.
ROM|12|6|Habentes autem donationes secundum gratiam, quae data est nobis, differentes: sive prophetiam, secundum rationem fidei;
ROM|12|7|sive ministerium, in ministrando; sive qui docet, in doctrina;
ROM|12|8|sive qui exhortatur, in exhortando; qui tribuit, in simplicitate; qui praeest, in sollicitudine; qui miseretur, in hilaritate.
ROM|12|9|Dilectio sine simulatione. Odientes malum, adhaerentes bono;
ROM|12|10|caritate fraternitatis invicem diligentes, honore invicem praevenientes,
ROM|12|11|sollicitudine non pigri, spiritu ferventes, Domino servientes,
ROM|12|12|spe gaudentes, in tribulatione patientes, orationi instantes,
ROM|12|13|necessitatibus sanctorum communicantes, hospitalitatem sectantes.
ROM|12|14|Benedicite persequentibus; benedicite et nolite maledicere!
ROM|12|15|Gaudere cum gaudentibus, flere cum flentibus.
ROM|12|16|Idipsum invicem sentientes, non alta sapientes, sed humilibus consentientes. Nolite esse prudentes apud vosmetipsos.
ROM|12|17|Nulli malum pro malo reddentes; providentes bona coram omnibus hominibus;
ROM|12|18|si fieri potest, quod ex vobis est, cum omnibus hominibus pacem habentes;
ROM|12|19|non vosmetipsos vindicantes, carissimi, sed date locum irae, scriptum est enim: " Mihi vindicta, ego retribuam ", dicit Dominus.
ROM|12|20|Sed si esurierit inimicus tuus, ciba illum; si sitit, potum da illi. Hoc enim faciens, carbones ignis congeres super caput eius.
ROM|12|21|Noli vinci a malo, sed vince in bono malum.
ROM|13|1|Omnis anima potestatibus sublimioribus subdita sit. Non est enim potestas nisi a Deo; quae autem sunt, a Deo ordinatae sunt.
ROM|13|2|Itaque, qui resistit potestati, Dei ordinationi resistit; qui autem resistunt ipsi, sibi damnationem acquirent.
ROM|13|3|Nam principes non sunt timori bono operi sed malo. Vis autem non timere potestatem? Bonum fac, et habebis laudem ex illa;
ROM|13|4|Dei enim ministra est tibi in bonum. Si autem malum feceris, time; non enim sine causa gladium portat; Dei enim ministra est, vindex in iram ei, qui malum agit.
ROM|13|5|Ideo necesse est subditos esse, non solum propter iram sed et propter conscientiam.
ROM|13|6|Ideo enim et tributa praestatis; ministri enim Dei sunt in hoc ipsum instantes.
ROM|13|7|Reddite omnibus debita: cui tributum tributum, cui vectigal vectigal, cui timorem timorem, cui honorem honorem.
ROM|13|8|Nemini quidquam debeatis, nisi ut invicem diligatis: qui enim diligit proximum, legem implevit.
ROM|13|9|Nam: Non adulterabis, Non occides, Non furaberis, Non concupisces, et si quod est aliud mandatum, in hoc verbo recapitulatur: Diliges proximum tuum tamquam teipsum.
ROM|13|10|Dilectio proximo malum non operatur; plenitudo ergo legis est dilectio.
ROM|13|11|Et hoc scientes tempus, quia hora est iam vos de somno surgere; nunc enim propior est nobis salus quam cum credidimus.
ROM|13|12|Nox processit, dies autem appropiavit. Abiciamus ergo opera tenebrarum et induamur arma lucis.
ROM|13|13|Sicut in die honeste ambulemus: non in comissationibus et ebrietatibus, non in cubilibus et impudicitiis, non in contentione et aemulatione;
ROM|13|14|sed induite Dominum Iesum Christum et carnis curam ne feceritis in concupiscentiis.
ROM|14|1|Infirmum autem in fide assumite, non in disceptatio nibus cogitationum.
ROM|14|2|Alius enim credit manducare omnia; qui autem infirmus est, holus manducat.
ROM|14|3|Is qui manducat, non manducantem non spernat; et, qui non manducat, manducantem non iudicet, Deus enim illum assumpsit.
ROM|14|4|Tu quis es, qui iudices alienum servum? Suo domino stat aut cadit; stabit autem, potens est enim Dominus statuere illum.
ROM|14|5|Nam alius iudicat inter diem et diem, alius iudicat omnem diem; unusquisque in suo sensu abundet.
ROM|14|6|Qui sapit diem, Domino sapit; et, qui manducat, Domino manducat, gratias enim agit Deo; et, qui non manducat, Domino non manducat et gratias agit Deo.
ROM|14|7|Nemo enim nostrum sibi vivit, et nemo sibi moritur;
ROM|14|8|sive enim vivimus, Domino vivimus, sive morimur, Domino morimur. Sive ergo vivimus, sive morimur, Domini sumus.
ROM|14|9|In hoc enim Christus et mortuus est et vixit, ut et mortuorum et vivorum dominetur.
ROM|14|10|Tu autem, quid iudicas fratrem tuum? Aut tu, quare spernis fratrem tuum? Omnes enim stabimus ante tribunal Dei;
ROM|14|11|scriptum est enim: Vivo ego, dicit Dominus,mihi flectetur omne genu,et omnis lingua confitebitur Deo ".
ROM|14|12|Itaque unusquisque nostrum pro se rationem reddet Deo.
ROM|14|13|Non ergo amplius invicem iudicemus, sed hoc iudicate magis, ne ponatis offendiculum fratri vel scandalum.
ROM|14|14|Scio et certus sum in Domino Iesu, quia nihil commune per seipsum, nisi ei, qui existimat quid commune esse, illi commune est.
ROM|14|15|Si enim propter cibum frater tuus contristatur, iam non secundum caritatem ambulas. Noli cibo tuo illum perdere, pro quo Christus mortuus est!
ROM|14|16|Non ergo blasphemetur bonum vestrum!
ROM|14|17|Non est enim regnum Dei esca et potus, sed iustitia et pax et gaudium in Spiritu Sancto;
ROM|14|18|qui enim in hoc servit Christo, placet Deo et probatus est hominibus.
ROM|14|19|Itaque, quae pacis sunt, sectemur et quae aedificationis sunt in invicem.
ROM|14|20|Noli propter escam destruere opus Dei! Omnia quidem munda sunt, sed malum est homini, qui per offendiculum manducat.
ROM|14|21|Bonum est non manducare carnem et non bibere vinum neque id, in quo frater tuus offendit.
ROM|14|22|Tu, quam fidem habes, penes temetipsum habe coram Deo. Beatus, qui non iudicat semetipsum in eo quod probat.
ROM|14|23|Qui autem discernit si manducaverit, damnatus est, quia non ex fide; omne autem, quod non ex fide, peccatum est.
ROM|15|1|Debemus autem nos fir miores imbecillitates infir morum sustinere et non nobis placere.
ROM|15|2|Unusquisque nostrum proximo placeat in bonum ad aedificationem;
ROM|15|3|etenim Christus non sibi placuit, sed sicut scriptum est: " Improperia improperantium tibi ceciderunt super me ".
ROM|15|4|Quaecumque enim antea scripta sunt, ad nostram doctrinam scripta sunt, ut per patientiam et consolationem Scripturarum spem habeamus.
ROM|15|5|Deus autem patientiae et solacii det vobis idipsum sapere in alterutrum secundum Christum Iesum,
ROM|15|6|ut unanimes uno ore glorificetis Deum et Patrem Domini nostri Iesu Christi.
ROM|15|7|Propter quod suscipite invicem, sicut et Christus suscepit vos, in gloriam Dei.
ROM|15|8|Dico enim Christum ministrum fuisse circumcisionis propter veritatem Dei ad confirmandas promissiones patrum;
ROM|15|9|gentes autem propter misericordiam glorificare Deum, sicut scriptum est: Propter hoc confitebor tibi in gentibus et nomini tuo cantabo ".
ROM|15|10|Et iterum dicit: " Laetamini, gentes, cum plebe eius ".
ROM|15|11|Et iterum: Laudate, omnes gentes, Dominum,et magnificent eum omnes populi ".
ROM|15|12|Et rursus Isaias ait: Erit radix Iesse,et qui exsurget regere gentes:in eo gentes sperabunt ".
ROM|15|13|Deus autem spei repleat vos omni gaudio et pace in credendo, ut abundetis in spe in virtute Spiritus Sancti.
ROM|15|14|Certus sum autem, fratres mei, et ego ipse de vobis, quoniam et ipsi pleni estis bonitate, repleti omni scientia, ita ut possitis et alterutrum monere.
ROM|15|15|Audacius autem scripsi vobis ex parte, tamquam in memoriam vos reducens propter gratiam, quae data est mihi a Deo,
ROM|15|16|ut sim minister Christi Iesu ad gentes, consecrans evangelium Dei, ut fiat oblatio gentium accepta, sanctificata in Spiritu Sancto.
ROM|15|17|Habeo igitur gloriationem in Christo Iesu ad Deum;
ROM|15|18|non enim audebo aliquid loqui eorum, quae per me non effecit Christus in oboedientiam gentium, verbo et factis,
ROM|15|19|in virtute signorum et prodigiorum, in virtute Spiritus, ita ut ab Ierusalem et per circuitum usque in Illyricum repleverim evangelium Christi,
ROM|15|20|sic autem contendens praedicare evangelium, non ubi nominatus est Christus, ne super alienum fundamentum aedificarem,
ROM|15|21|sed sicut scriptum est: Quibus non est annuntiatum de eo, videbunt;et, qui non audierunt, intellegent ".
ROM|15|22|Propter quod et impediebar plurimum venire ad vos;
ROM|15|23|nunc vero ulterius locum non habens in his regionibus, cupiditatem autem habens veniendi ad vos ex multis iam annis,
ROM|15|24|cum in Hispaniam proficisci coepero, spero enim quod praeteriens videam vos et a vobis deducar illuc, si vobis primum ex parte fruitus fuero.
ROM|15|25|Nunc autem proficiscor in Ierusalem ministrare sanctis;
ROM|15|26|probaverunt enim Macedonia et Achaia communicationem aliquam facere in pauperes sanctorum, qui sunt in Ierusalem.
ROM|15|27|Placuit enim eis, et debitores sunt eorum; nam si spiritalibus eorum communicaverunt gentes, debent et in carnalibus ministrare eis.
ROM|15|28|Hoc igitur cum consummavero et assignavero eis fructum hunc, proficiscar per vos in Hispaniam;
ROM|15|29|scio autem quoniam veniens ad vos, in abundantia benedictionis Christi veniam.
ROM|15|30|Obsecro autem vos, fratres, per Dominum nostrum Iesum Christum et per caritatem Spiritus, ut concertemini mecum in orationibus pro me ad Deum,
ROM|15|31|ut liberer ab infidelibus, qui sunt in Iudaea, et ministerium meum pro Ierusalem acceptum sit sanctis,
ROM|15|32|ut veniens ad vos in gaudio per voluntatem Dei refrigerer vobiscum.
ROM|15|33|Deus autem pacis sit cum omnibus vobis. Amen.
ROM|16|1|Commendo autem vobis Phoebem sororem nostram, quae est ministra ecclesiae, quae est Cenchreis,
ROM|16|2|ut eam suscipiatis in Domino digne sanctis et assistatis ei in quocumque negotio vestri indiguerit; etenim ipsa astitit multis et mihi ipsi.
ROM|16|3|Salutate Priscam et Aquilam adiutores meos in Christo Iesu,
ROM|16|4|qui pro anima mea suas cervices supposuerunt, quibus non solus ego gratias ago sed et cunctae ecclesiae gentium;
ROM|16|5|et domesticam eorum ecclesiam.Salutate Epaenetum dilectum mihi, primitias Asiae in Christo.
ROM|16|6|Salutate Mariam, quae multum laboravit in vobis.
ROM|16|7|Salutate Andronicum et Iuniam cognatos meos et concaptivos meos, qui sunt nobiles in apostolis, qui et ante me fuerunt in Christo.
ROM|16|8|Salutate Ampliatum dilectissimum mihi in Domino.
ROM|16|9|Salutate Urbanum adiutorem nostrum in Christo et Stachyn dilectum meum.
ROM|16|10|Salutate Apellem probatum in Christo. Salutate eos, qui sunt ex Aristobuli.
ROM|16|11|Salutate Herodionem cognatum meum. Salutate eos, qui sunt ex Narcissi, qui sunt in Domino.
ROM|16|12|Salutate Tryphaenam et Tryphosam, quae laborant in Domino. Salutate Persidam carissimam, quae multum laboravit in Domino.
ROM|16|13|Salutate Rufum electum in Domino et matrem eius et meam.
ROM|16|14|Salutate Asyncritum, Phlegonta, Hermen, Patrobam, Hermam et, qui cum eis sunt, fratres.
ROM|16|15|Salutate Philologum et Iuliam, Nereum et sororem eius et Olympam et omnes, qui cum eis sunt, sanctos.
ROM|16|16|Salutate invicem in osculo sancto. Salutant vos omnes ecclesiae Christi.
ROM|16|17|Rogo autem vos, fratres, ut observetis eos, qui dissensiones et offendicula praeter doctrinam, quam vos didicistis, faciunt, et declinate ab illis;
ROM|16|18|huiusmodi enim Domino nostro Christo non serviunt sed suo ventri, et per dulces sermones et benedictiones seducunt corda innocentium.
ROM|16|19|Vestra enim oboedientia ad omnes pervenit; gaudeo igitur in vobis, sed volo vos sapientes esse in bono et simplices in malo.
ROM|16|20|Deus autem pacis conteret Satanam sub pedibus vestris velociter.Gratia Domini nostri Iesu vobiscum.
ROM|16|21|Salutat vos Timotheus adiutor meus et Lucius et Iason et Sosipater cognati mei.
ROM|16|22|Saluto vos ego Tertius, qui scripsi epistulam in Domino.
ROM|16|23|Salutat vos Gaius hospes meus et universae ecclesiae. Salutat vos Erastus arcarius civitatis et Quartus frater.
ROM|16|24|()
ROM|16|25|Ei autem, qui potens est vos confirmare iuxta evangelium meum et praedicationem Iesu Christi secundum revelationem mysterii temporibus aeternis taciti,
ROM|16|26|manifestati autem nunc, et per scripturas Prophetarum secundum praeceptum aeterni Dei ad oboeditionem fidei in cunctis gentibus patefacti,
ROM|16|27|soli sapienti Deo per Iesum Christum, cui gloria in saecula. Amen.
