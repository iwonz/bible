MIC|1|1|verbum Domini quod factum est ad Micham Morasthiten in diebus Ioatham Ahaz Ezechiae regum Iuda quod vidit super Samariam et Hierusalem
MIC|1|2|audite populi omnes et adtendat terra et plenitudo eius et sit Dominus Deus vobis in testem Dominus de templo sancto suo
MIC|1|3|quia ecce Dominus egreditur de loco suo et descendet et calcabit super excelsa terrae
MIC|1|4|et consumentur montes subtus eum et valles scindentur sicut cera a facie ignis sicut aquae quae decurrunt in praeceps
MIC|1|5|in scelere Iacob omne istud et in peccatis domus Israhel quod scelus Iacob nonne Samaria et quae excelsa Iudae nonne Hierusalem
MIC|1|6|et ponam Samariam quasi acervum lapidum in agro cum plantatur vinea et detraham in vallem lapides eius et fundamenta eius revelabo
MIC|1|7|et omnia sculptilia eius concidentur et omnes mercedes eius conburentur igni et omnia idola eius ponam in perditionem quia de mercedibus meretricis congregata sunt et usque ad mercedem meretricis revertentur
MIC|1|8|super hoc plangam et ululabo vadam spoliatus et nudus faciam planctum velut draconum et luctum quasi strutionum
MIC|1|9|quia desperata est plaga eius quia venit usque ad Iudam tetigit portam populi mei usque ad Hierusalem
MIC|1|10|in Geth nolite adnuntiare lacrimis ne ploretis in domo Pulveris pulvere vos conspergite
MIC|1|11|et transite vobis habitatio Pulchra confusa ignominia non est egressa quae habitat in Exitu planctum domus Vicinae accipiet ex vobis quae stetit sibimet
MIC|1|12|quia infirmata est in bonum quae habitat in Amaritudinibus quia descendit malum a Domino in portam Hierusalem
MIC|1|13|tumultus quadrigae stuporis habitanti Lachis principium peccati est filiae Sion quia in te inventa sunt scelera Israhel
MIC|1|14|propterea dabit emissarios super hereditatem Geth domus Mendacii in deceptionem regibus Israhel
MIC|1|15|adhuc heredem adducam tibi quae habitas in Maresa usque Adollam veniet gloria Israhel
MIC|1|16|decalvare et tondere super filios deliciarum tuarum dilata calvitium tuum sicut aquila quoniam captivi ducti sunt ex te
MIC|2|1|vae qui cogitatis inutile et operamini malum in cubilibus vestris in luce matutina faciunt illud quoniam contra Deum est manus eorum
MIC|2|2|et concupierunt agros et violenter tulerunt et domos rapuerunt et calumniabantur virum et domum eius virum et hereditatem eius
MIC|2|3|idcirco haec dicit Dominus ecce ego cogito super familiam istam malum unde non auferetis colla vestra et non ambulabitis superbi quoniam tempus pessimum est
MIC|2|4|in die illa sumetur super vos parabola et cantabitur canticum cum suavitate dicentium depopulatione vastati sumus pars populi mei commutata est quomodo recedet a me cum revertatur qui regiones nostras dividat
MIC|2|5|propter hoc non erit tibi mittens funiculum sortis in coetu Domini
MIC|2|6|ne loquamini loquentes non stillabit super istos non conprehendet confusio
MIC|2|7|dicit domus Iacob numquid adbreviatus est spiritus Domini aut tales sunt cogitationes eius nonne verba mea bona sunt cum eo qui recte graditur
MIC|2|8|et e contrario populus meus in adversarium consurrexit desuper tunica pallium sustulistis eos qui transiebant simpliciter convertistis in bellum
MIC|2|9|mulieres populi mei eiecistis de domo deliciarum suarum a parvulis earum tulistis laudem meam in perpetuum
MIC|2|10|surgite et ite quia non habetis hic requiem propter inmunditiam eius corrumpetur putredine pessima
MIC|2|11|utinam non essem vir habens spiritum et mendacium potius loquerer stillabo tibi in vinum et in ebrietatem et erit super quem stillatur populus iste
MIC|2|12|congregatione congregabo Iacob totum te in unum conducam reliquias Israhel pariter ponam illum quasi gregem in ovili quasi pecus in medio caularum tumultuabuntur a multitudine hominum
MIC|2|13|ascendet enim pandens iter ante eos divident et transibunt portam et egredientur per eam et transibit rex eorum coram eis et Dominus in capite eorum
MIC|3|1|et dixi audite principes Iacob et duces domus Israhel numquid non vestrum est scire iudicium
MIC|3|2|qui odio habetis bonum et diligitis malum qui violenter tollitis pelles eorum desuper eos et carnem eorum desuper ossibus eorum
MIC|3|3|qui comederunt carnem populi mei et pellem eorum desuper excoriaverunt et ossa eorum confregerunt et conciderunt sicut in lebete et quasi carnem in medio ollae
MIC|3|4|tunc clamabunt ad Dominum et non exaudiet eos et abscondet faciem suam ab eis in tempore illo sicut nequiter egerunt in adinventionibus suis
MIC|3|5|haec dicit Dominus super prophetas qui seducunt populum meum qui mordent dentibus suis et praedicant pacem et si quis non dederit in ore eorum quippiam sanctificant super eum proelium
MIC|3|6|propterea nox vobis pro visione erit et tenebrae vobis pro divinatione et occumbet sol super prophetas et obtenebrabitur super eos dies
MIC|3|7|et confundentur qui vident visiones et confundentur divini et operient vultus suos omnes quia non est responsum Dei
MIC|3|8|verumtamen ego repletus sum fortitudine spiritus Domini iudicio et virtute ut adnuntiem Iacob scelus suum et Israhel peccatum suum
MIC|3|9|audite haec principes domus Iacob et iudices domus Israhel qui abominamini iudicium et omnia recta pervertitis
MIC|3|10|qui aedificatis Sion in sanguinibus et Hierusalem in iniquitate
MIC|3|11|principes eius in muneribus iudicabant et sacerdotes eius in mercede docebant et prophetae eius in pecunia divinabant et super Dominum requiescebant dicentes numquid non Dominus in medio nostrum non venient super nos mala
MIC|3|12|propter hoc causa vestri Sion quasi ager arabitur et Hierusalem quasi acervus lapidum erit et mons templi in excelsa silvarum
MIC|4|1|et in novissimo dierum erit mons domus Domini praeparatus in vertice montium et sublimis super colles et fluent ad eum populi
MIC|4|2|et properabunt gentes multae et dicent venite ascendamus ad montem Domini et ad domum Dei Iacob et docebit nos de viis suis et ibimus in semitis eius quia de Sion egredietur lex et verbum Domini de Hierusalem
MIC|4|3|et iudicabit inter populos multos et corripiet gentes fortes usque in longinquum et concident gladios suos in vomeres et hastas suas in ligones non sumet gens adversus gentem gladium et non discent ultra belligerare
MIC|4|4|et sedebit vir subtus vineam suam et subtus ficum suam et non erit qui deterreat quia os Domini exercituum locutum est
MIC|4|5|quia omnes populi ambulabunt unusquisque in nomine dei sui nos autem ambulabimus in nomine Domini Dei nostri in aeternum et ultra
MIC|4|6|in die illa dicit Dominus congregabo claudicantem et eam quam eieceram colligam et quam adflixeram
MIC|4|7|et ponam claudicantem in reliquias et eam quae laboraverat in gentem robustam et regnabit Dominus super eos in monte Sion ex hoc nunc et usque in aeternum
MIC|4|8|et tu turris Gregis nebulosa filiae Sion usque ad te veniet et veniet potestas prima regnum filiae Hierusalem
MIC|4|9|nunc quare maerore contraheris numquid rex non est tibi aut consiliarius tuus periit quia conprehendit te dolor sicut parturientem
MIC|4|10|dole et satage filia Sion quasi parturiens quia nunc egredieris de civitate et habitabis in regione et venies usque ad Babylonem ibi liberaberis ibi redimet te Dominus de manu inimicorum tuorum
MIC|4|11|et nunc congregatae sunt super te gentes multae quae dicunt lapidetur et aspiciat in Sion oculus noster
MIC|4|12|ipsi autem non cognoverunt cogitationes Domini et non intellexerunt consilium eius quia congregavit eos quasi faenum areae
MIC|4|13|surge et tritura filia Sion quia cornu tuum ponam ferreum et ungulas tuas ponam aereas et comminues populos multos et interficiam Domino rapinas eorum et fortitudinem eorum Domino universae terrae
MIC|5|1|nunc vastaberis filia latronis obsidionem posuerunt super nos in virga percutient maxillam iudicis Israhel
MIC|5|2|et tu Bethleem Ephrata parvulus es in milibus Iuda ex te mihi egredietur qui sit dominator in Israhel et egressus eius ab initio a diebus aeternitatis
MIC|5|3|propter hoc dabit eos usque ad tempus in quo parturiens pariet reliquiae fratrum eius convertentur ad filios Israhel
MIC|5|4|et stabit et pascet in fortitudine Domini in sublimitate nominis Domini Dei sui et convertentur quia nunc magnificabitur usque ad terminos terrae
MIC|5|5|et erit iste pax Assyrius cum venerit in terram nostram et quando calcaverit in domibus nostris et suscitabimus super eum septem pastores et octo primates homines
MIC|5|6|et pascent terram Assur in gladio et terram Nemrod in lanceis eius et liberabit ab Assur cum venerit in terram nostram et cum calcaverit in finibus nostris
MIC|5|7|et erunt reliquiae Iacob in medio populorum multorum quasi ros a Domino et quasi stillae super herbam quae non expectat virum et non praestolatur filios hominum
MIC|5|8|et erunt reliquiae Iacob in gentibus in medio populorum multorum quasi leo in iumentis silvarum et quasi catulus leonis in gregibus pecorum qui cum transierit et conculcaverit et ceperit non est qui eruat
MIC|5|9|exaltabitur manus tua super hostes tuos et omnes inimici tui interibunt
MIC|5|10|et erit in die illa dicit Dominus auferam equos tuos de medio tui et disperdam quadrigas tuas
MIC|5|11|et perdam civitates terrae tuae et destruam omnes munitiones tuas et auferam maleficia de manu tua et divinationes non erunt in te
MIC|5|12|et perire faciam sculptilia tua et statuas tuas de medio tui et non adorabis ultra opera manuum tuarum
MIC|5|13|et evellam lucos tuos de medio tui et conteram civitates tuas
MIC|5|14|et faciam in furore et in indignatione ultionem in omnibus gentibus quae non audierunt
MIC|6|1|audite quae Dominus loquitur surge contende iudicio adversum montes et audiant colles vocem tuam
MIC|6|2|audiant montes iudicium Domini et fortia fundamenta terrae quia iudicium Domini cum populo suo et cum Israhel diiudicabitur
MIC|6|3|populus meus quid feci tibi et quid molestus fui tibi responde mihi
MIC|6|4|quia eduxi te de terra Aegypti et de domo servientium liberavi te et misi ante faciem tuam Mosen et Aaron et Mariam
MIC|6|5|populus meus memento quaeso quid cogitaverit Balac rex Moab et quid responderit ei Balaam filius Beor de Setthim usque ad Galgalam ut cognosceret iustitias Domini
MIC|6|6|quid dignum offeram Domino curvem genu Deo excelso numquid offeram ei holocaustomata et vitulos anniculos
MIC|6|7|numquid placari potest Dominus in milibus arietum aut in multis milibus hircorum pinguium numquid dabo primogenitum meum pro scelere meo fructum ventris mei pro peccato animae meae
MIC|6|8|indicabo tibi o homo quid sit bonum et quid Dominus quaerat a te utique facere iudicium et diligere misericordiam et sollicitum ambulare cum Deo tuo
MIC|6|9|vox Domini ad civitatem clamat et salus erit timentibus nomen tuum audite tribus et quis adprobabit illud
MIC|6|10|adhuc ignis in domo impii thesauri iniquitatis et mensura minor irae plena
MIC|6|11|numquid iustificabo stateram impiam et saccelli pondera dolosa
MIC|6|12|in quibus divites eius repleti sunt iniquitate et habitantes in ea loquebantur mendacium et lingua eorum fraudulenta in ore eorum
MIC|6|13|et ego ergo coepi percutere te perditione super peccatis tuis
MIC|6|14|tu comedes et non saturaberis et humiliatio tua in medio tui et adprehendes et non salvabis et quos salvaveris in gladium dabo
MIC|6|15|tu seminabis et non metes tu calcabis olivam et non ungueris oleo et mustum et non bibes vinum
MIC|6|16|et custodisti praecepta Omri et omne opus domus Achab et ambulasti in voluntatibus eorum ut darem te in perditionem et habitantes in ea in sibilum et obprobrium populi mei portabitis
MIC|7|1|vae mihi quia factus sum sicut qui colligit in autumno racemos vindemiae non est botrus ad comedendum praecoquas ficus desideravit anima mea
MIC|7|2|periit sanctus de terra et rectus in hominibus non est omnes in sanguine insidiantur vir fratrem suum venatur ad mortem
MIC|7|3|malum manuum suarum dicunt bonum princeps postulat et iudex in reddendo est et magnus locutus est desiderium animae suae et conturbaverunt eam
MIC|7|4|qui optimus in eis est quasi paliurus et qui rectus quasi spina de sepe dies speculationis tuae visitatio tua venit nunc erit vastitas eorum
MIC|7|5|nolite credere amico et nolite confidere in duce ab ea quae dormit in sinu tuo custodi claustra oris tui
MIC|7|6|quia filius contumeliam facit patri filia consurgit adversus matrem suam nurus contra socrum suam inimici hominis domestici eius
MIC|7|7|ego autem ad Dominum aspiciam expectabo Deum salvatorem meum audiet me Deus meus
MIC|7|8|ne laeteris inimica mea super me quia cecidi consurgam cum sedero in tenebris Dominus lux mea est
MIC|7|9|iram Domini portabo quoniam peccavi ei donec iudicet causam meam et faciat iudicium meum educet me in lucem videbo in iustitiam eius
MIC|7|10|et aspiciet inimica mea et operietur confusione quae dicit ad me ubi est Dominus Deus tuus oculi mei videbunt in eam nunc erit in conculcationem ut lutum platearum
MIC|7|11|dies ut aedificentur maceriae tuae in die illa longe fiet lex
MIC|7|12|in die illa et usque ad te veniet Assur et usque ad civitates munitas et a civitatibus munitis usque ad flumen et ad mare de mari et ad montem de monte
MIC|7|13|et erit terra in desolationem propter habitatores suos et propter fructum cogitationum eorum
MIC|7|14|pasce populum tuum in virga tua gregem hereditatis tuae habitantes solos in saltu in medio Carmeli pascentur Basan et Galaad iuxta dies antiquos
MIC|7|15|secundum dies egressionis tuae de terra Aegypti ostendam ei mirabilia
MIC|7|16|videbunt gentes et confundentur super omni fortitudine sua ponent manus super os aures eorum surdae erunt
MIC|7|17|lingent pulverem sicut serpens velut reptilia terrae proturbabuntur de aedibus suis Dominum Deum nostrum desiderabunt et timebunt te
MIC|7|18|quis Deus similis tui qui aufers iniquitatem et transis peccatum reliquiarum hereditatis tuae non inmittet ultra furorem suum quoniam volens misericordiam est
MIC|7|19|revertetur et miserebitur nostri deponet iniquitates nostras et proiciet in profundum maris omnia peccata nostra
MIC|7|20|dabis veritatem Iacob misericordiam Abraham quae iurasti patribus nostris a diebus antiquis
