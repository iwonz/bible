2TIM|1|1|Павел, волею Божиею Апостол Иисуса Христа, по обетованию жизни во Христе Иисусе,
2TIM|1|2|Тимофею, возлюбленному сыну: благодать, милость, мир от Бога Отца и Христа Иисуса, Господа нашего.
2TIM|1|3|Благодарю Бога, Которому служу от прародителей с чистою совестью, что непрестанно вспоминаю о тебе в молитвах моих днем и ночью,
2TIM|1|4|и желаю видеть тебя, вспоминая о слезах твоих, дабы мне исполниться радости,
2TIM|1|5|приводя на память нелицемерную веру твою, которая прежде обитала в бабке твоей Лоиде и матери твоей Евнике; уверен, что она и в тебе.
2TIM|1|6|По сей причине напоминаю тебе возгревать дар Божий, который в тебе через мое рукоположение;
2TIM|1|7|ибо дал нам Бог духа не боязни, но силы и любви и целомудрия.
2TIM|1|8|Итак, не стыдись свидетельства Господа нашего Иисуса Христа, ни меня, узника Его; но страдай с благовестием Христовым силою Бога,
2TIM|1|9|спасшего нас и призвавшего званием святым, не по делам нашим, но по Своему изволению и благодати, данной нам во Христе Иисусе прежде вековых времен,
2TIM|1|10|открывшейся же ныне явлением Спасителя нашего Иисуса Христа, разрушившего смерть и явившего жизнь и нетление через благовестие,
2TIM|1|11|для которого я поставлен проповедником и Апостолом и учителем язычников.
2TIM|1|12|По сей причине я и страдаю так; но не стыжусь. Ибо я знаю, в Кого уверовал, и уверен, что Он силен сохранить залог мой на оный день.
2TIM|1|13|Держись образца здравого учения, которое ты слышал от меня, с верою и любовью во Христе Иисусе.
2TIM|1|14|Храни добрый залог Духом Святым, живущим в нас.
2TIM|1|15|Ты знаешь, что все Асийские оставили меня; в числе их Фигелл и Ермоген.
2TIM|1|16|Да даст Господь милость дому Онисифора за то, что он многократно покоил меня и не стыдился уз моих,
2TIM|1|17|но, быв в Риме, с великим тщанием искал меня и нашел.
2TIM|1|18|Да даст ему Господь обрести милость у Господа в оный день; а сколько он служил мне в Ефесе, ты лучше знаешь.
2TIM|2|1|Итак укрепляйся, сын мой, в благодати Христом Иисусом,
2TIM|2|2|и что слышал от меня при многих свидетелях, то передай верным людям, которые были бы способны и других научить.
2TIM|2|3|Итак переноси страдания, как добрый воин Иисуса Христа.
2TIM|2|4|Никакой воин не связывает себя делами житейскими, чтобы угодить военачальнику.
2TIM|2|5|Если же кто и подвизается, не увенчивается, если незаконно будет подвизаться.
2TIM|2|6|Трудящемуся земледельцу первому должно вкусить от плодов.
2TIM|2|7|Разумей, что я говорю. Да даст тебе Господь разумение во всем.
2TIM|2|8|Помни Господа Иисуса Христа от семени Давидова, воскресшего из мертвых, по благовествованию моему,
2TIM|2|9|за которое я страдаю даже до уз, как злодей; но для слова Божия нет уз.
2TIM|2|10|Посему я все терплю ради избранных, дабы и они получили спасение во Христе Иисусе с вечною славою.
2TIM|2|11|Верно слово: если мы с Ним умерли, то с Ним и оживем;
2TIM|2|12|если терпим, то с Ним и царствовать будем; если отречемся, и Он отречется от нас;
2TIM|2|13|если мы неверны, Он пребывает верен, ибо Себя отречься не может.
2TIM|2|14|Сие напоминай, заклиная пред Господом не вступать в словопрения, что нимало не служит к пользе, а к расстройству слушающих.
2TIM|2|15|Старайся представить себя Богу достойным, делателем неукоризненным, верно преподающим слово истины.
2TIM|2|16|А непотребного пустословия удаляйся; ибо они еще более будут преуспевать в нечестии,
2TIM|2|17|и слово их, как рак, будет распространяться. Таковы Именей и Филит,
2TIM|2|18|которые отступили от истины, говоря, что воскресение уже было, и разрушают в некоторых веру.
2TIM|2|19|Но твердое основание Божие стоит, имея печать сию: "познал Господь Своих"; и: "да отступит от неправды всякий, исповедующий имя Господа".
2TIM|2|20|А в большом доме есть сосуды не только золотые и серебряные, но и деревянные и глиняные; и одни в почетном, а другие в низком употреблении.
2TIM|2|21|Итак, кто будет чист от сего, тот будет сосудом в чести, освященным и благопотребным Владыке, годным на всякое доброе дело.
2TIM|2|22|Юношеских похотей убегай, а держись правды, веры, любви, мира со всеми призывающими Господа от чистого сердца.
2TIM|2|23|От глупых и невежественных состязаний уклоняйся, зная, что они рождают ссоры;
2TIM|2|24|рабу же Господа не должно ссориться, но быть приветливым ко всем, учительным, незлобивым,
2TIM|2|25|с кротостью наставлять противников, не даст ли им Бог покаяния к познанию истины,
2TIM|2|26|чтобы они освободились от сети диавола, который уловил их в свою волю.
2TIM|3|1|Знай же, что в последние дни наступят времена тяжкие.
2TIM|3|2|Ибо люди будут самолюбивы, сребролюбивы, горды, надменны, злоречивы, родителям непокорны, неблагодарны, нечестивы, недружелюбны,
2TIM|3|3|непримирительны, клеветники, невоздержны, жестоки, не любящие добра,
2TIM|3|4|предатели, наглы, напыщенны, более сластолюбивы, нежели боголюбивы,
2TIM|3|5|имеющие вид благочестия, силы же его отрекшиеся. Таковых удаляйся.
2TIM|3|6|К сим принадлежат те, которые вкрадываются в домы и обольщают женщин, утопающих во грехах, водимых различными похотями,
2TIM|3|7|всегда учащихся и никогда не могущих дойти до познания истины.
2TIM|3|8|Как Ианний и Иамврий противились Моисею, так и сии противятся истине, люди, развращенные умом, невежды в вере.
2TIM|3|9|Но они не много успеют; ибо их безумие обнаружится перед всеми, как и с теми случилось.
2TIM|3|10|А ты последовал мне в учении, житии, расположении, вере, великодушии, любви, терпении,
2TIM|3|11|в гонениях, страданиях, постигших меня в Антиохии, Иконии, Листрах; каковые гонения я перенес, и от всех избавил меня Господь.
2TIM|3|12|Да и все, желающие жить благочестиво во Христе Иисусе, будут гонимы.
2TIM|3|13|Злые же люди и обманщики будут преуспевать во зле, вводя в заблуждение и заблуждаясь.
2TIM|3|14|А ты пребывай в том, чему научен и что тебе вверено, зная, кем ты научен.
2TIM|3|15|Притом же ты из детства знаешь священные писания, которые могут умудрить тебя во спасение верою во Христа Иисуса.
2TIM|3|16|Все Писание богодухновенно и полезно для научения, для обличения, для исправления, для наставления в праведности,
2TIM|3|17|да будет совершен Божий человек, ко всякому доброму делу приготовлен.
2TIM|4|1|Итак заклинаю тебя пред Богом и Господом нашим Иисусом Христом, Который будет судить живых и мертвых в явление Его и Царствие Его:
2TIM|4|2|проповедуй слово, настой во время и не во время, обличай, запрещай, увещевай со всяким долготерпением и назиданием.
2TIM|4|3|Ибо будет время, когда здравого учения принимать не будут, но по своим прихотям будут избирать себе учителей, которые льстили бы слуху;
2TIM|4|4|и от истины отвратят слух и обратятся к басням.
2TIM|4|5|Но ты будь бдителен во всем, переноси скорби, совершай дело благовестника, исполняй служение твое.
2TIM|4|6|Ибо я уже становлюсь жертвою, и время моего отшествия настало.
2TIM|4|7|Подвигом добрым я подвизался, течение совершил, веру сохранил;
2TIM|4|8|а теперь готовится мне венец правды, который даст мне Господь, праведный Судия, в день оный; и не только мне, но и всем, возлюбившим явление Его.
2TIM|4|9|Постарайся придти ко мне скоро.
2TIM|4|10|Ибо Димас оставил меня, возлюбив нынешний век, и пошел в Фессалонику, Крискент в Галатию, Тит в Далматию; один Лука со мною.
2TIM|4|11|Марка возьми и приведи с собою, ибо он мне нужен для служения.
2TIM|4|12|Тихика я послал в Ефес.
2TIM|4|13|Когда пойдешь, принеси фелонь, который я оставил в Троаде у Карпа, и книги, особенно кожаные.
2TIM|4|14|Александр медник много сделал мне зла. Да воздаст ему Господь по делам его!
2TIM|4|15|Берегись его и ты, ибо он сильно противился нашим словам.
2TIM|4|16|При первом моем ответе никого не было со мною, но все меня оставили. Да не вменится им!
2TIM|4|17|Господь же предстал мне и укрепил меня, дабы через меня утвердилось благовестие и услышали все язычники; и я избавился из львиных челюстей.
2TIM|4|18|И избавит меня Господь от всякого злого дела и сохранит для Своего Небесного Царства, Ему слава во веки веков. Аминь.
2TIM|4|19|Приветствуй Прискиллу и Акилу и дом Онисифоров.
2TIM|4|20|Ераст остался в Коринфе; Трофима же я оставил больного в Милите.
2TIM|4|21|Постарайся придти до зимы. Приветствуют тебя Еввул, и Пуд, и Лин, и Клавдия, и все братия.
2TIM|4|22|Господь Иисус Христос со духом твоим. Благодать с вами. Аминь.
