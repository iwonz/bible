TITUS|1|1|Paul, a servant of God and an apostle of Jesus Christ, for the sake of the faith of God's elect and their knowledge of the truth, which accords with godliness,
TITUS|1|2|in hope of eternal life, which God, who never lies, promised before the ages began
TITUS|1|3|and at the proper time manifested in his word through the preaching with which I have been entrusted by the command of God our Savior;
TITUS|1|4|To Titus, my true child in a common faith: Grace and peace from God the Father and Christ Jesus our Savior.
TITUS|1|5|This is why I left you in Crete, so that you might put what remained into order, and appoint elders in every town as I directed you-
TITUS|1|6|if anyone is above reproach, the husband of one wife, and his children are believers and not open to the charge of debauchery or insubordination.
TITUS|1|7|For an overseer, as God's steward, must be above reproach. He must not be arrogant or quick-tempered or a drunkard or violent or greedy for gain,
TITUS|1|8|but hospitable, a lover of good, self-controlled, upright, holy, and disciplined.
TITUS|1|9|He must hold firm to the trustworthy word as taught, so that he may be able to give instruction in sound doctrine and also to rebuke those who contradict it.
TITUS|1|10|For there are many who are insubordinate, empty talkers and deceivers, especially those of the circumcision party.
TITUS|1|11|They must be silenced, since they are upsetting whole families by teaching for shameful gain what they ought not to teach.
TITUS|1|12|One of the Cretans, a prophet of their own, said, "Cretans are always liars, evil beasts, lazy gluttons."
TITUS|1|13|This testimony is true. Therefore rebuke them sharply, that they may be sound in the faith,
TITUS|1|14|not devoting themselves to Jewish myths and the commands of people who turn away from the truth.
TITUS|1|15|To the pure, all things are pure, but to the defiled and unbelieving, nothing is pure; but both their minds and their consciences are defiled.
TITUS|1|16|They profess to know God, but they deny him by their works. They are detestable, disobedient, unfit for any good work.
TITUS|2|1|But as for you, teach what accords with sound doctrine.
TITUS|2|2|Older men are to be sober-minded, dignified, self-controlled, sound in faith, in love, and in steadfastness.
TITUS|2|3|Older women likewise are to be reverent in behavior, not slanderers or slaves to much wine. They are to teach what is good,
TITUS|2|4|and so train the young women to love their husbands and children,
TITUS|2|5|to be self-controlled, pure, working at home, kind, and submissive to their own husbands, that the word of God may not be reviled.
TITUS|2|6|Likewise, urge the younger men to be self-controlled.
TITUS|2|7|Show yourself in all respects to be a model of good works, and in your teaching show integrity, dignity,
TITUS|2|8|and sound speech that cannot be condemned, so that an opponent may be put to shame, having nothing evil to say about us.
TITUS|2|9|Slaves are to be submissive to their own masters in everything; they are to be well-pleasing, not argumentative,
TITUS|2|10|not pilfering, but showing all good faith, so that in everything they may adorn the doctrine of God our Savior.
TITUS|2|11|For the grace of God has appeared, bringing salvation for all people,
TITUS|2|12|training us to renounce ungodliness and worldly passions, and to live self-controlled, upright, and godly lives in the present age,
TITUS|2|13|waiting for our blessed hope, the appearing of the glory of our great God and Savior Jesus Christ,
TITUS|2|14|who gave himself for us to redeem us from all lawlessness and to purify for himself a people for his own possession who are zealous for good works.
TITUS|2|15|Declare these things; exhort and rebuke with all authority. Let no one disregard you.
TITUS|3|1|Remind them to be submissive to rulers and authorities, to be obedient, to be ready for every good work,
TITUS|3|2|to speak evil of no one, to avoid quarreling, to be gentle, and to show perfect courtesy toward all people.
TITUS|3|3|For we ourselves were once foolish, disobedient, led astray, slaves to various passions and pleasures, passing our days in malice and envy, hated by others and hating one another.
TITUS|3|4|But when the goodness and loving kindness of God our Savior appeared,
TITUS|3|5|he saved us, not because of works done by us in righteousness, but according to his own mercy, by the washing of regeneration and renewal of the Holy Spirit,
TITUS|3|6|whom he poured out on us richly through Jesus Christ our Savior,
TITUS|3|7|so that being justified by his grace we might become heirs according to the hope of eternal life.
TITUS|3|8|The saying is trustworthy, and I want you to insist on these things, so that those who have believed in God may be careful to devote themselves to good works. These things are excellent and profitable for people.
TITUS|3|9|But avoid foolish controversies, genealogies, dissensions, and quarrels about the law, for they are unprofitable and worthless.
TITUS|3|10|As for a person who stirs up division, after warning him once and then twice, have nothing more to do with him,
TITUS|3|11|knowing that such a person is warped and sinful; he is self-condemned.
TITUS|3|12|When I send Artemas or Tychicus to you, do your best to come to me at Nicopolis, for I have decided to spend the winter there.
TITUS|3|13|Do your best to speed Zenas the lawyer and Apollos on their way; see that they lack nothing.
TITUS|3|14|And let our people learn to devote themselves to good works, so as to help cases of urgent need, and not be unfruitful.
TITUS|3|15|All who are with me send greetings to you. Greet those who love us in the faith. Grace be with you all.
