LUKE|1|1|Как уже многие начали составлять повествования о совершенно известных между нами событиях,
LUKE|1|2|как передали нам то бывшие с самого начала очевидцами и служителями Слова,
LUKE|1|3|то рассудилось и мне, по тщательном исследовании всего сначала, по порядку описать тебе, достопочтенный Феофил,
LUKE|1|4|чтобы ты узнал твердое основание того учения, в котором был наставлен.
LUKE|1|5|Во дни Ирода, царя Иудейского, был священник из Авиевой чреды, именем Захария, и жена его из рода Ааронова, имя ей Елисавета.
LUKE|1|6|Оба они были праведны пред Богом, поступая по всем заповедям и уставам Господним беспорочно.
LUKE|1|7|У них не было детей, ибо Елисавета была неплодна, и оба были уже в летах преклонных.
LUKE|1|8|Однажды, когда он в порядке своей чреды служил пред Богом,
LUKE|1|9|по жребию, как обыкновенно было у священников, досталось ему войти в храм Господень для каждения,
LUKE|1|10|а все множество народа молилось вне во время каждения, –
LUKE|1|11|тогда явился ему Ангел Господень, стоя по правую сторону жертвенника кадильного.
LUKE|1|12|Захария, увидев его, смутился, и страх напал на него.
LUKE|1|13|Ангел же сказал ему: не бойся, Захария, ибо услышана молитва твоя, и жена твоя Елисавета родит тебе сына, и наречешь ему имя: Иоанн;
LUKE|1|14|и будет тебе радость и веселие, и многие о рождении его возрадуются,
LUKE|1|15|ибо он будет велик пред Господом; не будет пить вина и сикера, и Духа Святаго исполнится еще от чрева матери своей;
LUKE|1|16|и многих из сынов Израилевых обратит к Господу Богу их;
LUKE|1|17|и предъидет пред Ним в духе и силе Илии, чтобы возвратить сердца отцов детям, и непокоривым образ мыслей праведников, дабы представить Господу народ приготовленный.
LUKE|1|18|И сказал Захария Ангелу: по чему я узнаю это? ибо я стар, и жена моя в летах преклонных.
LUKE|1|19|Ангел сказал ему в ответ: я Гавриил, предстоящий пред Богом, и послан говорить с тобою и благовестить тебе сие;
LUKE|1|20|и вот, ты будешь молчать и не будешь иметь возможности говорить до того дня, как это сбудется, за то, что ты не поверил словам моим, которые сбудутся в свое время.
LUKE|1|21|Между тем народ ожидал Захарию и дивился, что он медлит в храме.
LUKE|1|22|Он же, выйдя, не мог говорить к ним; и они поняли, что он видел видение в храме; и он объяснялся с ними знаками, и оставался нем.
LUKE|1|23|А когда окончились дни службы его, возвратился в дом свой.
LUKE|1|24|После сих дней зачала Елисавета, жена его, и таилась пять месяцев и говорила:
LUKE|1|25|так сотворил мне Господь во дни сии, в которые призрел на меня, чтобы снять с меня поношение между людьми.
LUKE|1|26|В шестой же месяц послан был Ангел Гавриил от Бога в город Галилейский, называемый Назарет,
LUKE|1|27|к Деве, обрученной мужу, именем Иосифу, из дома Давидова; имя же Деве: Мария.
LUKE|1|28|Ангел, войдя к Ней, сказал: радуйся, Благодатная! Господь с Тобою; благословенна Ты между женами.
LUKE|1|29|Она же, увидев его, смутилась от слов его и размышляла, что бы это было за приветствие.
LUKE|1|30|И сказал Ей Ангел: не бойся, Мария, ибо Ты обрела благодать у Бога;
LUKE|1|31|и вот, зачнешь во чреве, и родишь Сына, и наречешь Ему имя: Иисус.
LUKE|1|32|Он будет велик и наречется Сыном Всевышнего, и даст Ему Господь Бог престол Давида, отца Его;
LUKE|1|33|и будет царствовать над домом Иакова во веки, и Царству Его не будет конца.
LUKE|1|34|Мария же сказала Ангелу: как будет это, когда Я мужа не знаю?
LUKE|1|35|Ангел сказал Ей в ответ: Дух Святый найдет на Тебя, и сила Всевышнего осенит Тебя; посему и рождаемое Святое наречется Сыном Божиим.
LUKE|1|36|Вот и Елисавета, родственница Твоя, называемая неплодною, и она зачала сына в старости своей, и ей уже шестой месяц,
LUKE|1|37|ибо у Бога не останется бессильным никакое слово.
LUKE|1|38|Тогда Мария сказала: се, Раба Господня; да будет Мне по слову твоему. И отошел от Нее Ангел.
LUKE|1|39|Встав же Мария во дни сии, с поспешностью пошла в нагорную страну, в город Иудин,
LUKE|1|40|и вошла в дом Захарии, и приветствовала Елисавету.
LUKE|1|41|Когда Елисавета услышала приветствие Марии, взыграл младенец во чреве ее; и Елисавета исполнилась Святаго Духа,
LUKE|1|42|и воскликнула громким голосом, и сказала: благословенна Ты между женами, и благословен плод чрева Твоего!
LUKE|1|43|И откуда это мне, что пришла Матерь Господа моего ко мне?
LUKE|1|44|Ибо когда голос приветствия Твоего дошел до слуха моего, взыграл младенец радостно во чреве моем.
LUKE|1|45|И блаженна Уверовавшая, потому что совершится сказанное Ей от Господа.
LUKE|1|46|И сказала Мария: величит душа Моя Господа,
LUKE|1|47|и возрадовался дух Мой о Боге, Спасителе Моем,
LUKE|1|48|что призрел Он на смирение Рабы Своей, ибо отныне будут ублажать Меня все роды;
LUKE|1|49|что сотворил Мне величие Сильный, и свято имя Его;
LUKE|1|50|и милость Его в роды родов к боящимся Его;
LUKE|1|51|явил силу мышцы Своей; рассеял надменных помышлениями сердца их;
LUKE|1|52|низложил сильных с престолов, и вознес смиренных;
LUKE|1|53|алчущих исполнил благ, и богатящихся отпустил ни с чем;
LUKE|1|54|воспринял Израиля, отрока Своего, воспомянув милость,
LUKE|1|55|как говорил отцам нашим, к Аврааму и семени его до века.
LUKE|1|56|Пребыла же Мария с нею около трех месяцев, и возвратилась в дом свой.
LUKE|1|57|Елисавете же настало время родить, и она родила сына.
LUKE|1|58|И услышали соседи и родственники ее, что возвеличил Господь милость Свою над нею, и радовались с нею.
LUKE|1|59|В восьмой день пришли обрезать младенца и хотели назвать его, по имени отца его, Захариею.
LUKE|1|60|На это мать его сказала: нет, а назвать его Иоанном.
LUKE|1|61|И сказали ей: никого нет в родстве твоем, кто назывался бы сим именем.
LUKE|1|62|И спрашивали знаками у отца его, как бы он хотел назвать его.
LUKE|1|63|Он потребовал дощечку и написал: Иоанн имя ему. И все удивились.
LUKE|1|64|И тотчас разрешились уста его и язык его, и он стал говорить, благословляя Бога.
LUKE|1|65|И был страх на всех живущих вокруг них; и рассказывали обо всем этом по всей нагорной стране Иудейской.
LUKE|1|66|Все слышавшие положили это на сердце своем и говорили: что будет младенец сей? И рука Господня была с ним.
LUKE|1|67|И Захария, отец его, исполнился Святаго Духа и пророчествовал, говоря:
LUKE|1|68|благословен Господь Бог Израилев, что посетил народ Свой и сотворил избавление ему,
LUKE|1|69|и воздвиг рог спасения нам в дому Давида, отрока Своего,
LUKE|1|70|как возвестил устами бывших от века святых пророков Своих,
LUKE|1|71|что спасет нас от врагов наших и от руки всех ненавидящих нас;
LUKE|1|72|сотворит милость с отцами нашими и помянет святой завет Свой,
LUKE|1|73|клятву, которою клялся Он Аврааму, отцу нашему, дать нам,
LUKE|1|74|небоязненно, по избавлении от руки врагов наших,
LUKE|1|75|служить Ему в святости и правде пред Ним, во все дни жизни нашей.
LUKE|1|76|И ты, младенец, наречешься пророком Всевышнего, ибо предъидешь пред лицем Господа приготовить пути Ему,
LUKE|1|77|дать уразуметь народу Его спасение в прощении грехов их,
LUKE|1|78|по благоутробному милосердию Бога нашего, которым посетил нас Восток свыше,
LUKE|1|79|просветить сидящих во тьме и тени смертной, направить ноги наши на путь мира.
LUKE|1|80|Младенец же возрастал и укреплялся духом, и был в пустынях до дня явления своего Израилю.
LUKE|2|1|В те дни вышло от кесаря Августа повеление сделать перепись по всей земле.
LUKE|2|2|Эта перепись была первая в правление Квириния Сириею.
LUKE|2|3|И пошли все записываться, каждый в свой город.
LUKE|2|4|Пошел также и Иосиф из Галилеи, из города Назарета, в Иудею, в город Давидов, называемый Вифлеем, потому что он был из дома и рода Давидова,
LUKE|2|5|записаться с Мариею, обрученною ему женою, которая была беременна.
LUKE|2|6|Когда же они были там, наступило время родить Ей;
LUKE|2|7|и родила Сына своего Первенца, и спеленала Его, и положила Его в ясли, потому что не было им места в гостинице.
LUKE|2|8|В той стране были на поле пастухи, которые содержали ночную стражу у стада своего.
LUKE|2|9|Вдруг предстал им Ангел Господень, и слава Господня осияла их; и убоялись страхом великим.
LUKE|2|10|И сказал им Ангел: не бойтесь; я возвещаю вам великую радость, которая будет всем людям:
LUKE|2|11|ибо ныне родился вам в городе Давидовом Спаситель, Который есть Христос Господь;
LUKE|2|12|и вот вам знак: вы найдете Младенца в пеленах, лежащего в яслях.
LUKE|2|13|И внезапно явилось с Ангелом многочисленное воинство небесное, славящее Бога и взывающее:
LUKE|2|14|слава в вышних Богу, и на земле мир, в человеках благоволение!
LUKE|2|15|Когда Ангелы отошли от них на небо, пастухи сказали друг другу: пойдем в Вифлеем и посмотрим, что там случилось, о чем возвестил нам Господь.
LUKE|2|16|И, поспешив, пришли и нашли Марию и Иосифа, и Младенца, лежащего в яслях.
LUKE|2|17|Увидев же, рассказали о том, что было возвещено им о Младенце Сем.
LUKE|2|18|И все слышавшие дивились тому, что рассказывали им пастухи.
LUKE|2|19|А Мария сохраняла все слова сии, слагая в сердце Своем.
LUKE|2|20|И возвратились пастухи, славя и хваля Бога за все то, что слышали и видели, как им сказано было.
LUKE|2|21|По прошествии восьми дней, когда надлежало обрезать [Младенца], дали Ему имя Иисус, нареченное Ангелом прежде зачатия Его во чреве.
LUKE|2|22|А когда исполнились дни очищения их по закону Моисееву, принесли Его в Иерусалим, чтобы представить пред Господа,
LUKE|2|23|как предписано в законе Господнем, чтобы всякий младенец мужеского пола, разверзающий ложесна, был посвящен Господу,
LUKE|2|24|и чтобы принести в жертву, по реченному в законе Господнем, две горлицы или двух птенцов голубиных.
LUKE|2|25|Тогда был в Иерусалиме человек, именем Симеон. Он был муж праведный и благочестивый, чающий утешения Израилева; и Дух Святый был на нем.
LUKE|2|26|Ему было предсказано Духом Святым, что он не увидит смерти, доколе не увидит Христа Господня.
LUKE|2|27|И пришел он по вдохновению в храм. И, когда родители принесли Младенца Иисуса, чтобы совершить над Ним законный обряд,
LUKE|2|28|он взял Его на руки, благословил Бога и сказал:
LUKE|2|29|Ныне отпускаешь раба Твоего, Владыко, по слову Твоему, с миром,
LUKE|2|30|ибо видели очи мои спасение Твое,
LUKE|2|31|которое Ты уготовал пред лицем всех народов,
LUKE|2|32|свет к просвещению язычников и славу народа Твоего Израиля.
LUKE|2|33|Иосиф же и Матерь Его дивились сказанному о Нем.
LUKE|2|34|И благословил их Симеон и сказал Марии, Матери Его: се, лежит Сей на падение и на восстание многих в Израиле и в предмет пререканий, –
LUKE|2|35|и Тебе Самой оружие пройдет душу, – да откроются помышления многих сердец.
LUKE|2|36|Тут была также Анна пророчица, дочь Фануилова, от колена Асирова, достигшая глубокой старости, прожив с мужем от девства своего семь лет,
LUKE|2|37|вдова лет восьмидесяти четырех, которая не отходила от храма, постом и молитвою служа Богу день и ночь.
LUKE|2|38|И она в то время, подойдя, славила Господа и говорила о Нем всем, ожидавшим избавления в Иерусалиме.
LUKE|2|39|И когда они совершили все по закону Господню, возвратились в Галилею, в город свой Назарет.
LUKE|2|40|Младенец же возрастал и укреплялся духом, исполняясь премудрости, и благодать Божия была на Нем.
LUKE|2|41|Каждый год родители Его ходили в Иерусалим на праздник Пасхи.
LUKE|2|42|И когда Он был двенадцати лет, пришли они также по обычаю в Иерусалим на праздник.
LUKE|2|43|Когда же, по окончании дней [праздника], возвращались, остался Отрок Иисус в Иерусалиме; и не заметили того Иосиф и Матерь Его,
LUKE|2|44|но думали, что Он идет с другими. Пройдя же дневной путь, стали искать Его между родственниками и знакомыми
LUKE|2|45|и, не найдя Его, возвратились в Иерусалим, ища Его.
LUKE|2|46|Через три дня нашли Его в храме, сидящего посреди учителей, слушающего их и спрашивающего их;
LUKE|2|47|все слушавшие Его дивились разуму и ответам Его.
LUKE|2|48|И, увидев Его, удивились; и Матерь Его сказала Ему: Чадо! что Ты сделал с нами? Вот, отец Твой и Я с великою скорбью искали Тебя.
LUKE|2|49|Он сказал им: зачем было вам искать Меня? или вы не знали, что Мне должно быть в том, что принадлежит Отцу Моему?
LUKE|2|50|Но они не поняли сказанных Им слов.
LUKE|2|51|И Он пошел с ними и пришел в Назарет; и был в повиновении у них. И Матерь Его сохраняла все слова сии в сердце Своем.
LUKE|2|52|Иисус же преуспевал в премудрости и возрасте и в любви у Бога и человеков.
LUKE|3|1|В пятнадцатый же год правления Тиверия кесаря, когда Понтий Пилат начальствовал в Иудее, Ирод был четвертовластником в Галилее, Филипп, брат его, четвертовластником в Итурее и Трахонитской области, а Лисаний четвертовластником в Авилинее,
LUKE|3|2|при первосвященниках Анне и Каиафе, был глагол Божий к Иоанну, сыну Захарии, в пустыне.
LUKE|3|3|И он проходил по всей окрестной стране Иорданской, проповедуя крещение покаяния для прощения грехов,
LUKE|3|4|как написано в книге слов пророка Исаии, который говорит: глас вопиющего в пустыне: приготовьте путь Господу, прямыми сделайте стези Ему;
LUKE|3|5|всякий дол да наполнится, и всякая гора и холм да понизятся, кривизны выпрямятся и неровные пути сделаются гладкими;
LUKE|3|6|и узрит всякая плоть спасение Божие.
LUKE|3|7|[Иоанн] приходившему креститься от него народу говорил: порождения ехиднины! кто внушил вам бежать от будущего гнева?
LUKE|3|8|Сотворите же достойные плоды покаяния и не думайте говорить в себе: отец у нас Авраам, ибо говорю вам, что Бог может из камней сих воздвигнуть детей Аврааму.
LUKE|3|9|Уже и секира при корне дерев лежит: всякое дерево, не приносящее доброго плода, срубают и бросают в огонь.
LUKE|3|10|И спрашивал его народ: что же нам делать?
LUKE|3|11|Он сказал им в ответ: у кого две одежды, тот дай неимущему, и у кого есть пища, делай то же.
LUKE|3|12|Пришли и мытари креститься, и сказали ему: учитель! что нам делать?
LUKE|3|13|Он отвечал им: ничего не требуйте более определенного вам.
LUKE|3|14|Спрашивали его также и воины: а нам что делать? И сказал им: никого не обижайте, не клевещите, и довольствуйтесь своим жалованьем.
LUKE|3|15|Когда же народ был в ожидании, и все помышляли в сердцах своих об Иоанне, не Христос ли он, –
LUKE|3|16|Иоанн всем отвечал: я крещу вас водою, но идет Сильнейший меня, у Которого я недостоин развязать ремень обуви; Он будет крестить вас Духом Святым и огнем.
LUKE|3|17|Лопата Его в руке Его, и Он очистит гумно Свое и соберет пшеницу в житницу Свою, а солому сожжет огнем неугасимым.
LUKE|3|18|Многое и другое благовествовал он народу, поучая его.
LUKE|3|19|Ирод же четвертовластник, обличаемый от него за Иродиаду, жену брата своего, и за все, что сделал Ирод худого,
LUKE|3|20|прибавил ко всему прочему и то, что заключил Иоанна в темницу.
LUKE|3|21|Когда же крестился весь народ, и Иисус, крестившись, молился: отверзлось небо,
LUKE|3|22|и Дух Святый нисшел на Него в телесном виде, как голубь, и был глас с небес, глаголющий: Ты Сын Мой Возлюбленный; в Тебе Мое благоволение!
LUKE|3|23|Иисус, начиная [Свое служение], был лет тридцати, и был, как думали, Сын Иосифов, Илиев,
LUKE|3|24|Матфатов, Левиин, Мелхиев, Ианнаев, Иосифов,
LUKE|3|25|Маттафиев, Амосов, Наумов, Еслимов, Наггеев,
LUKE|3|26|Маафов, Маттафиев, Семеиев, Иосифов, Иудин,
LUKE|3|27|Иоаннанов, Рисаев, Зоровавелев, Салафиилев, Нириев,
LUKE|3|28|Мелхиев, Аддиев, Косамов, Елмодамов, Иров,
LUKE|3|29|Иосиев, Елиезеров, Иоримов, Матфатов, Левиин,
LUKE|3|30|Симеонов, Иудин, Иосифов, Ионанов, Елиакимов,
LUKE|3|31|Мелеаев, Маинанов, Маттафаев, Нафанов, Давидов,
LUKE|3|32|Иессеев, Овидов, Воозов, Салмонов, Наассонов,
LUKE|3|33|Аминадавов, Арамов, Есромов, Фаресов, Иудин,
LUKE|3|34|Иаковлев, Исааков, Авраамов, Фаррин, Нахоров,
LUKE|3|35|Серухов, Рагавов, Фалеков, Еверов, Салин,
LUKE|3|36|Каинанов, Арфаксадов, Симов, Ноев, Ламехов,
LUKE|3|37|Мафусалов, Енохов, Иаредов, Малелеилов, Каинанов,
LUKE|3|38|Еносов, Сифов, Адамов, Божий.
LUKE|4|1|Иисус, исполненный Духа Святаго, возвратился от Иордана и поведен был Духом в пустыню.
LUKE|4|2|Там сорок дней Он был искушаем от диавола и ничего не ел в эти дни, а по прошествии их напоследок взалкал.
LUKE|4|3|И сказал Ему диавол: если Ты Сын Божий, то вели этому камню сделаться хлебом.
LUKE|4|4|Иисус сказал ему в ответ: написано, что не хлебом одним будет жить человек, но всяким словом Божиим.
LUKE|4|5|И, возведя Его на высокую гору, диавол показал Ему все царства вселенной во мгновение времени,
LUKE|4|6|и сказал Ему диавол: Тебе дам власть над всеми сими [царствами] и славу их, ибо она предана мне, и я, кому хочу, даю ее;
LUKE|4|7|итак, если Ты поклонишься мне, то все будет Твое.
LUKE|4|8|Иисус сказал ему в ответ: отойди от Меня, сатана; написано: Господу Богу твоему поклоняйся, и Ему одному служи.
LUKE|4|9|И повел Его в Иерусалим, и поставил Его на крыле храма, и сказал Ему: если Ты Сын Божий, бросься отсюда вниз,
LUKE|4|10|ибо написано: Ангелам Своим заповедает о Тебе сохранить Тебя;
LUKE|4|11|и на руках понесут Тебя, да не преткнешься о камень ногою Твоею.
LUKE|4|12|Иисус сказал ему в ответ: сказано: не искушай Господа Бога твоего.
LUKE|4|13|И, окончив все искушение, диавол отошел от Него до времени.
LUKE|4|14|И возвратился Иисус в силе духа в Галилею; и разнеслась молва о Нем по всей окрестной стране.
LUKE|4|15|Он учил в синагогах их, и от всех был прославляем.
LUKE|4|16|И пришел в Назарет, где был воспитан, и вошел, по обыкновению Своему, в день субботний в синагогу, и встал читать.
LUKE|4|17|Ему подали книгу пророка Исаии; и Он, раскрыв книгу, нашел место, где было написано:
LUKE|4|18|Дух Господень на Мне; ибо Он помазал Меня благовествовать нищим, и послал Меня исцелять сокрушенных сердцем, проповедывать пленным освобождение, слепым прозрение, отпустить измученных на свободу,
LUKE|4|19|проповедывать лето Господне благоприятное.
LUKE|4|20|И, закрыв книгу и отдав служителю, сел; и глаза всех в синагоге были устремлены на Него.
LUKE|4|21|И Он начал говорить им: ныне исполнилось писание сие, слышанное вами.
LUKE|4|22|И все засвидетельствовали Ему это, и дивились словам благодати, исходившим из уст Его, и говорили: не Иосифов ли это сын?
LUKE|4|23|Он сказал им: конечно, вы скажете Мне присловие: врач! исцели Самого Себя; сделай и здесь, в Твоем отечестве, то, что, мы слышали, было в Капернауме.
LUKE|4|24|И сказал: истинно говорю вам: никакой пророк не принимается в своем отечестве.
LUKE|4|25|Поистине говорю вам: много вдов было в Израиле во дни Илии, когда заключено было небо три года и шесть месяцев, так что сделался большой голод по всей земле,
LUKE|4|26|и ни к одной из них не был послан Илия, а только ко вдове в Сарепту Сидонскую;
LUKE|4|27|много также было прокаженных в Израиле при пророке Елисее, и ни один из них не очистился, кроме Неемана Сириянина.
LUKE|4|28|Услышав это, все в синагоге исполнились ярости
LUKE|4|29|и, встав, выгнали Его вон из города и повели на вершину горы, на которой город их был построен, чтобы свергнуть Его;
LUKE|4|30|но Он, пройдя посреди них, удалился.
LUKE|4|31|И пришел в Капернаум, город Галилейский, и учил их в дни субботние.
LUKE|4|32|И дивились учению Его, ибо слово Его было со властью.
LUKE|4|33|Был в синагоге человек, имевший нечистого духа бесовского, и он закричал громким голосом:
LUKE|4|34|оставь; что Тебе до нас, Иисус Назарянин? Ты пришел погубить нас; знаю Тебя, кто Ты, Святый Божий.
LUKE|4|35|Иисус запретил ему, сказав: замолчи и выйди из него. И бес, повергнув его посреди [синагоги], вышел из него, нимало не повредив ему.
LUKE|4|36|И напал на всех ужас, и рассуждали между собою: что это значит, что Он со властью и силою повелевает нечистым духам, и они выходят?
LUKE|4|37|И разнесся слух о Нем по всем окрестным местам.
LUKE|4|38|Выйдя из синагоги, Он вошел в дом Симона; теща же Симонова была одержима сильною горячкою; и просили Его о ней.
LUKE|4|39|Подойдя к ней, Он запретил горячке; и оставила ее. Она тотчас встала и служила им.
LUKE|4|40|При захождении же солнца все, имевшие больных различными болезнями, приводили их к Нему и Он, возлагая на каждого из них руки, исцелял их.
LUKE|4|41|Выходили также и бесы из многих с криком и говорили: Ты Христос, Сын Божий. А Он запрещал им сказывать, что они знают, что Он Христос.
LUKE|4|42|Когда же настал день, Он, выйдя [из дома], пошел в пустынное место, и народ искал Его и, придя к Нему, удерживал Его, чтобы не уходил от них.
LUKE|4|43|Но Он сказал им: и другим городам благовествовать Я должен Царствие Божие, ибо на то Я послан.
LUKE|4|44|И проповедывал в синагогах галилейских.
LUKE|5|1|Однажды, когда народ теснился к Нему, чтобы слышать слово Божие, а Он стоял у озера Геннисаретского,
LUKE|5|2|увидел Он две лодки, стоящие на озере; а рыболовы, выйдя из них, вымывали сети.
LUKE|5|3|Войдя в одну лодку, которая была Симонова, Он просил его отплыть несколько от берега и, сев, учил народ из лодки.
LUKE|5|4|Когда же перестал учить, сказал Симону: отплыви на глубину и закиньте сети свои для лова.
LUKE|5|5|Симон сказал Ему в ответ: Наставник! мы трудились всю ночь и ничего не поймали, но по слову Твоему закину сеть.
LUKE|5|6|Сделав это, они поймали великое множество рыбы, и даже сеть у них прорывалась.
LUKE|5|7|И дали знак товарищам, находившимся на другой лодке, чтобы пришли помочь им; и пришли, и наполнили обе лодки, так что они начинали тонуть.
LUKE|5|8|Увидев это, Симон Петр припал к коленям Иисуса и сказал: выйди от меня, Господи! потому что я человек грешный.
LUKE|5|9|Ибо ужас объял его и всех, бывших с ним, от этого лова рыб, ими пойманных;
LUKE|5|10|также и Иакова и Иоанна, сыновей Зеведеевых, бывших товарищами Симону. И сказал Симону Иисус: не бойся; отныне будешь ловить человеков.
LUKE|5|11|И, вытащив обе лодки на берег, оставили все и последовали за Ним.
LUKE|5|12|Когда Иисус был в одном городе, пришел человек весь в проказе и, увидев Иисуса, пал ниц, умоляя Его и говоря: Господи! если хочешь, можешь меня очистить.
LUKE|5|13|Он простер руку, прикоснулся к нему и сказал: хочу, очистись. И тотчас проказа сошла с него.
LUKE|5|14|И Он повелел ему никому не сказывать, а пойти показаться священнику и принести [жертву] за очищение свое, как повелел Моисей, во свидетельство им.
LUKE|5|15|Но тем более распространялась молва о Нем, и великое множество народа стекалось к Нему слушать и врачеваться у Него от болезней своих.
LUKE|5|16|Но Он уходил в пустынные места и молился.
LUKE|5|17|В один день, когда Он учил, и сидели тут фарисеи и законоучители, пришедшие из всех мест Галилеи и Иудеи и из Иерусалима, и сила Господня являлась в исцелении [больных], –
LUKE|5|18|вот, принесли некоторые на постели человека, который был расслаблен, и старались внести его [в дом] и положить перед Иисусом;
LUKE|5|19|и, не найдя, где пронести его за многолюдством, влезли на верх дома и сквозь кровлю спустили его с постелью на средину пред Иисуса.
LUKE|5|20|И Он, видя веру их, сказал человеку тому: прощаются тебе грехи твои.
LUKE|5|21|Книжники и фарисеи начали рассуждать, говоря: кто это, который богохульствует? кто может прощать грехи, кроме одного Бога?
LUKE|5|22|Иисус, уразумев помышления их, сказал им в ответ: что вы помышляете в сердцах ваших?
LUKE|5|23|Что легче сказать: прощаются тебе грехи твои, или сказать: встань и ходи?
LUKE|5|24|Но чтобы вы знали, что Сын Человеческий имеет власть на земле прощать грехи, – сказал Он расслабленному: тебе говорю: встань, возьми постель твою и иди в дом твой.
LUKE|5|25|И он тотчас встал перед ними, взял, на чем лежал, и пошел в дом свой, славя Бога.
LUKE|5|26|И ужас объял всех, и славили Бога и, быв исполнены страха, говорили: чудные дела видели мы ныне.
LUKE|5|27|После сего [Иисус] вышел и увидел мытаря, именем Левия, сидящего у сбора пошлин, и говорит ему: следуй за Мною.
LUKE|5|28|И он, оставив все, встал и последовал за Ним.
LUKE|5|29|И сделал для Него Левий в доме своем большое угощение; и там было множество мытарей и других, которые возлежали с ними.
LUKE|5|30|Книжники же и фарисеи роптали и говорили ученикам Его: зачем вы едите и пьете с мытарями и грешниками?
LUKE|5|31|Иисус же сказал им в ответ: не здоровые имеют нужду во враче, но больные;
LUKE|5|32|Я пришел призвать не праведников, а грешников к покаянию.
LUKE|5|33|Они же сказали Ему: почему ученики Иоанновы постятся часто и молитвы творят, также и фарисейские, а Твои едят и пьют?
LUKE|5|34|Он сказал им: можете ли заставить сынов чертога брачного поститься, когда с ними жених?
LUKE|5|35|Но придут дни, когда отнимется у них жених, и тогда будут поститься в те дни.
LUKE|5|36|При сем сказал им притчу: никто не приставляет заплаты к ветхой одежде, отодрав от новой одежды; а иначе и новую раздерет, и к старой не подойдет заплата от новой.
LUKE|5|37|И никто не вливает молодого вина в мехи ветхие; а иначе молодое вино прорвет мехи, и само вытечет, и мехи пропадут;
LUKE|5|38|но молодое вино должно вливать в мехи новые; тогда сбережется и то и другое.
LUKE|5|39|И никто, пив старое [вино], не захочет тотчас молодого, ибо говорит: старое лучше.
LUKE|6|1|В субботу, первую по втором дне Пасхи, случилось Ему проходить засеянными полями, и ученики Его срывали колосья и ели, растирая руками.
LUKE|6|2|Некоторые же из фарисеев сказали им: зачем вы делаете то, чего не должно делать в субботы?
LUKE|6|3|Иисус сказал им в ответ: разве вы не читали, что сделал Давид, когда взалкал сам и бывшие с ним?
LUKE|6|4|Как он вошел в дом Божий, взял хлебы предложения, которых не должно было есть никому, кроме одних священников, и ел, и дал бывшим с ним?
LUKE|6|5|И сказал им: Сын Человеческий есть господин и субботы.
LUKE|6|6|Случилось же и в другую субботу войти Ему в синагогу и учить. Там был человек, у которого правая рука была сухая.
LUKE|6|7|Книжники же и фарисеи наблюдали за Ним, не исцелит ли в субботу, чтобы найти обвинение против Него.
LUKE|6|8|Но Он, зная помышления их, сказал человеку, имеющему сухую руку: встань и выступи на средину. И он встал и выступил.
LUKE|6|9|Тогда сказал им Иисус: спрошу Я вас: что должно делать в субботу? добро, или зло? спасти душу, или погубить? Они молчали.
LUKE|6|10|И, посмотрев на всех их, сказал тому человеку: протяни руку твою. Он так и сделал; и стала рука его здорова, как другая.
LUKE|6|11|Они же пришли в бешенство и говорили между собою, что бы им сделать с Иисусом.
LUKE|6|12|В те дни взошел Он на гору помолиться и пробыл всю ночь в молитве к Богу.
LUKE|6|13|Когда же настал день, призвал учеников Своих и избрал из них двенадцать, которых и наименовал Апостолами:
LUKE|6|14|Симона, которого и назвал Петром, и Андрея, брата его, Иакова и Иоанна, Филиппа и Варфоломея,
LUKE|6|15|Матфея и Фому, Иакова Алфеева и Симона, прозываемого Зилотом,
LUKE|6|16|Иуду Иаковлева и Иуду Искариота, который потом сделался предателем.
LUKE|6|17|И, сойдя с ними, стал Он на ровном месте, и множество учеников Его, и много народа из всей Иудеи и Иерусалима и приморских мест Тирских и Сидонских,
LUKE|6|18|которые пришли послушать Его и исцелиться от болезней своих, также и страждущие от нечистых духов; и исцелялись.
LUKE|6|19|И весь народ искал прикасаться к Нему, потому что от Него исходила сила и исцеляла всех.
LUKE|6|20|И Он, возведя очи Свои на учеников Своих, говорил: Блаженны нищие духом, ибо ваше есть Царствие Божие.
LUKE|6|21|Блаженны алчущие ныне, ибо насытитесь. Блаженны плачущие ныне, ибо воссмеетесь.
LUKE|6|22|Блаженны вы, когда возненавидят вас люди и когда отлучат вас, и будут поносить, и пронесут имя ваше, как бесчестное, за Сына Человеческого.
LUKE|6|23|Возрадуйтесь в тот день и возвеселитесь, ибо велика вам награда на небесах. Так поступали с пророками отцы их.
LUKE|6|24|Напротив, горе вам, богатые! ибо вы уже получили свое утешение.
LUKE|6|25|Горе вам, пресыщенные ныне! ибо взалчете. Горе вам, смеющиеся ныне! ибо восплачете и возрыдаете.
LUKE|6|26|Горе вам, когда все люди будут говорить о вас хорошо! ибо так поступали с лжепророками отцы их.
LUKE|6|27|Но вам, слушающим, говорю: любите врагов ваших, благотворите ненавидящим вас,
LUKE|6|28|благословляйте проклинающих вас и молитесь за обижающих вас.
LUKE|6|29|Ударившему тебя по щеке подставь и другую, и отнимающему у тебя верхнюю одежду не препятствуй взять и рубашку.
LUKE|6|30|Всякому, просящему у тебя, давай, и от взявшего твое не требуй назад.
LUKE|6|31|И как хотите, чтобы с вами поступали люди, так и вы поступайте с ними.
LUKE|6|32|И если любите любящих вас, какая вам за то благодарность? ибо и грешники любящих их любят.
LUKE|6|33|И если делаете добро тем, которые вам делают добро, какая вам за то благодарность? ибо и грешники то же делают.
LUKE|6|34|И если взаймы даете тем, от которых надеетесь получить обратно, какая вам за то благодарность? ибо и грешники дают взаймы грешникам, чтобы получить обратно столько же.
LUKE|6|35|Но вы любите врагов ваших, и благотворите, и взаймы давайте, не ожидая ничего; и будет вам награда великая, и будете сынами Всевышнего; ибо Он благ и к неблагодарным и злым.
LUKE|6|36|Итак, будьте милосерды, как и Отец ваш милосерд.
LUKE|6|37|Не судите, и не будете судимы; не осуждайте, и не будете осуждены; прощайте, и прощены будете;
LUKE|6|38|давайте, и дастся вам: мерою доброю, утрясенною, нагнетенною и переполненною отсыплют вам в лоно ваше; ибо, какою мерою мерите, такою же отмерится и вам.
LUKE|6|39|Сказал также им притчу: может ли слепой водить слепого? не оба ли упадут в яму?
LUKE|6|40|Ученик не бывает выше своего учителя; но, и усовершенствовавшись, будет всякий, как учитель его.
LUKE|6|41|Что ты смотришь на сучок в глазе брата твоего, а бревна в твоем глазе не чувствуешь?
LUKE|6|42|Или, как можешь сказать брату твоему: брат! дай, я выну сучок из глаза твоего, когда сам не видишь бревна в твоем глазе? Лицемер! вынь прежде бревно из твоего глаза, и тогда увидишь, как вынуть сучок из глаза брата твоего.
LUKE|6|43|Нет доброго дерева, которое приносило бы худой плод; и нет худого дерева, которое приносило бы плод добрый,
LUKE|6|44|ибо всякое дерево познается по плоду своему, потому что не собирают смокв с терновника и не снимают винограда с кустарника.
LUKE|6|45|Добрый человек из доброго сокровища сердца своего выносит доброе, а злой человек из злого сокровища сердца своего выносит злое, ибо от избытка сердца говорят уста его.
LUKE|6|46|Что вы зовете Меня: Господи! Господи! – и не делаете того, что Я говорю?
LUKE|6|47|Всякий, приходящий ко Мне и слушающий слова Мои и исполняющий их, скажу вам, кому подобен.
LUKE|6|48|Он подобен человеку, строящему дом, который копал, углубился и положил основание на камне; почему, когда случилось наводнение и вода наперла на этот дом, то не могла поколебать его, потому что он основан был на камне.
LUKE|6|49|А слушающий и неисполняющий подобен человеку, построившему дом на земле без основания, который, когда наперла на него вода, тотчас обрушился; и разрушение дома сего было великое.
LUKE|7|1|Когда Он окончил все слова Свои к слушавшему народу, то вошел в Капернаум.
LUKE|7|2|У одного сотника слуга, которым он дорожил, был болен при смерти.
LUKE|7|3|Услышав об Иисусе, он послал к Нему Иудейских старейшин просить Его, чтобы пришел исцелить слугу его.
LUKE|7|4|И они, придя к Иисусу, просили Его убедительно, говоря: он достоин, чтобы Ты сделал для него это,
LUKE|7|5|ибо он любит народ наш и построил нам синагогу.
LUKE|7|6|Иисус пошел с ними. И когда Он недалеко уже был от дома, сотник прислал к Нему друзей сказать Ему: не трудись, Господи! ибо я недостоин, чтобы Ты вошел под кров мой;
LUKE|7|7|потому и себя самого не почел я достойным придти к Тебе; но скажи слово, и выздоровеет слуга мой.
LUKE|7|8|Ибо я и подвластный человек, но, имея у себя в подчинении воинов, говорю одному: пойди, и идет; и другому: приди, и приходит; и слуге моему: сделай то, и делает.
LUKE|7|9|Услышав сие, Иисус удивился ему и, обратившись, сказал идущему за Ним народу: сказываю вам, что и в Израиле не нашел Я такой веры.
LUKE|7|10|Посланные, возвратившись в дом, нашли больного слугу выздоровевшим.
LUKE|7|11|После сего Иисус пошел в город, называемый Наин; и с Ним шли многие из учеников Его и множество народа.
LUKE|7|12|Когда же Он приблизился к городским воротам, тут выносили умершего, единственного сына у матери, а она была вдова; и много народа шло с нею из города.
LUKE|7|13|Увидев ее, Господь сжалился над нею и сказал ей: не плачь.
LUKE|7|14|И, подойдя, прикоснулся к одру; несшие остановились, и Он сказал: юноша! тебе говорю, встань!
LUKE|7|15|Мертвый, поднявшись, сел и стал говорить; и отдал его [Иисус] матери его.
LUKE|7|16|И всех объял страх, и славили Бога, говоря: великий пророк восстал между нами, и Бог посетил народ Свой.
LUKE|7|17|Такое мнение о Нем распространилось по всей Иудее и по всей окрестности.
LUKE|7|18|И возвестили Иоанну ученики его о всем том.
LUKE|7|19|Иоанн, призвав двоих из учеников своих, послал к Иисусу спросить: Ты ли Тот, Который должен придти, или ожидать нам другого?
LUKE|7|20|Они, придя к [Иисусу], сказали: Иоанн Креститель послал нас к Тебе спросить: Ты ли Тот, Которому должно придти, или другого ожидать нам?
LUKE|7|21|А в это время Он многих исцелил от болезней и недугов и от злых духов, и многим слепым даровал зрение.
LUKE|7|22|И сказал им Иисус в ответ: пойдите, скажите Иоанну, что вы видели и слышали: слепые прозревают, хромые ходят, прокаженные очищаются, глухие слышат, мертвые воскресают, нищие благовествуют;
LUKE|7|23|и блажен, кто не соблазнится о Мне!
LUKE|7|24|По отшествии же посланных Иоанном, начал говорить к народу об Иоанне: что смотреть ходили вы в пустыню? трость ли, ветром колеблемую?
LUKE|7|25|Что же смотреть ходили вы? человека ли, одетого в мягкие одежды? Но одевающиеся пышно и роскошно живущие находятся при дворах царских.
LUKE|7|26|Что же смотреть ходили вы? пророка ли? Да, говорю вам, и больше пророка.
LUKE|7|27|Сей есть, о котором написано: вот, Я посылаю Ангела Моего пред лицем Твоим, который приготовит путь Твой пред Тобою.
LUKE|7|28|Ибо говорю вам: из рожденных женами нет ни одного пророка больше Иоанна Крестителя; но меньший в Царствии Божием больше его.
LUKE|7|29|И весь народ, слушавший [Его], и мытари воздали славу Богу, крестившись крещением Иоанновым;
LUKE|7|30|а фарисеи и законники отвергли волю Божию о себе, не крестившись от него.
LUKE|7|31|Тогда Господь сказал: с кем сравню людей рода сего? и кому они подобны?
LUKE|7|32|Они подобны детям, которые сидят на улице, кличут друг друга и говорят: мы играли вам на свирели, и вы не плясали; мы пели вам плачевные песни, и вы не плакали.
LUKE|7|33|Ибо пришел Иоанн Креститель: ни хлеба не ест, ни вина не пьет; и говорите: в нем бес.
LUKE|7|34|Пришел Сын Человеческий: ест и пьет; и говорите: вот человек, который любит есть и пить вино, друг мытарям и грешникам.
LUKE|7|35|И оправдана премудрость всеми чадами ее.
LUKE|7|36|Некто из фарисеев просил Его вкусить с ним пищи; и Он, войдя в дом фарисея, возлег.
LUKE|7|37|И вот, женщина того города, которая была грешница, узнав, что Он возлежит в доме фарисея, принесла алавастровый сосуд с миром
LUKE|7|38|и, став позади у ног Его и плача, начала обливать ноги Его слезами и отирать волосами головы своей, и целовала ноги Его, и мазала миром.
LUKE|7|39|Видя это, фарисей, пригласивший Его, сказал сам в себе: если бы Он был пророк, то знал бы, кто и какая женщина прикасается к Нему, ибо она грешница.
LUKE|7|40|Обратившись к нему, Иисус сказал: Симон! Я имею нечто сказать тебе. Он говорит: скажи, Учитель.
LUKE|7|41|Иисус сказал: у одного заимодавца было два должника: один должен был пятьсот динариев, а другой пятьдесят,
LUKE|7|42|но как они не имели чем заплатить, он простил обоим. Скажи же, который из них более возлюбит его?
LUKE|7|43|Симон отвечал: думаю, тот, которому более простил. Он сказал ему: правильно ты рассудил.
LUKE|7|44|И, обратившись к женщине, сказал Симону: видишь ли ты эту женщину? Я пришел в дом твой, и ты воды Мне на ноги не дал, а она слезами облила Мне ноги и волосами головы своей отерла;
LUKE|7|45|ты целования Мне не дал, а она, с тех пор как Я пришел, не перестает целовать у Меня ноги;
LUKE|7|46|ты головы Мне маслом не помазал, а она миром помазала Мне ноги.
LUKE|7|47|А потому сказываю тебе: прощаются грехи ее многие за то, что она возлюбила много, а кому мало прощается, тот мало любит.
LUKE|7|48|Ей же сказал: прощаются тебе грехи.
LUKE|7|49|И возлежавшие с Ним начали говорить про себя: кто это, что и грехи прощает?
LUKE|7|50|Он же сказал женщине: вера твоя спасла тебя, иди с миром.
LUKE|8|1|После сего Он проходил по городам и селениям, проповедуя и благовествуя Царствие Божие, и с Ним двенадцать,
LUKE|8|2|и некоторые женщины, которых Он исцелил от злых духов и болезней: Мария, называемая Магдалиною, из которой вышли семь бесов,
LUKE|8|3|и Иоанна, жена Хузы, домоправителя Иродова, и Сусанна, и многие другие, которые служили Ему имением своим.
LUKE|8|4|Когда же собралось множество народа, и из всех городов жители сходились к Нему, Он начал говорить притчею:
LUKE|8|5|вышел сеятель сеять семя свое, и когда он сеял, иное упало при дороге и было потоптано, и птицы небесные поклевали его;
LUKE|8|6|а иное упало на камень и, взойдя, засохло, потому что не имело влаги;
LUKE|8|7|а иное упало между тернием, и выросло терние и заглушило его;
LUKE|8|8|а иное упало на добрую землю и, взойдя, принесло плод сторичный. Сказав сие, возгласил: кто имеет уши слышать, да слышит!
LUKE|8|9|Ученики же Его спросили у Него: что бы значила притча сия?
LUKE|8|10|Он сказал: вам дано знать тайны Царствия Божия, а прочим в притчах, так что они видя не видят и слыша не разумеют.
LUKE|8|11|Вот что значит притча сия: семя есть слово Божие;
LUKE|8|12|а упавшее при пути, это суть слушающие, к которым потом приходит диавол и уносит слово из сердца их, чтобы они не уверовали и не спаслись;
LUKE|8|13|а упавшее на камень, это те, которые, когда услышат слово, с радостью принимают, но которые не имеют корня, и временем веруют, а во время искушения отпадают;
LUKE|8|14|а упавшее в терние, это те, которые слушают слово, но, отходя, заботами, богатством и наслаждениями житейскими подавляются и не приносят плода;
LUKE|8|15|а упавшее на добрую землю, это те, которые, услышав слово, хранят его в добром и чистом сердце и приносят плод в терпении. Сказав это, Он возгласил: кто имеет уши слышать, да слышит!
LUKE|8|16|Никто, зажегши свечу, не покрывает ее сосудом, или не ставит под кровать, а ставит на подсвечник, чтобы входящие видели свет.
LUKE|8|17|Ибо нет ничего тайного, что не сделалось бы явным, ни сокровенного, что не сделалось бы известным и не обнаружилось бы.
LUKE|8|18|Итак, наблюдайте, как вы слушаете: ибо, кто имеет, тому дано будет, а кто не имеет, у того отнимется и то, что он думает иметь.
LUKE|8|19|И пришли к Нему Матерь и братья Его, и не могли подойти к Нему по причине народа.
LUKE|8|20|И дали знать Ему: Матерь и братья Твои стоят вне, желая видеть Тебя.
LUKE|8|21|Он сказал им в ответ: матерь Моя и братья Мои суть слушающие слово Божие и исполняющие его.
LUKE|8|22|В один день Он вошел с учениками Своими в лодку и сказал им: переправимся на ту сторону озера. И отправились.
LUKE|8|23|Во время плавания их Он заснул. На озере поднялся бурный ветер, и заливало их [волнами], и они были в опасности.
LUKE|8|24|И, подойдя, разбудили Его и сказали: Наставник! Наставник! погибаем. Но Он, встав, запретил ветру и волнению воды; и перестали, и сделалась тишина.
LUKE|8|25|Тогда Он сказал им: где вера ваша? Они же в страхе и удивлении говорили друг другу: кто же это, что и ветрам повелевает и воде, и повинуются Ему?
LUKE|8|26|И приплыли в страну Гадаринскую, лежащую против Галилеи.
LUKE|8|27|Когда же вышел Он на берег, встретил Его один человек из города, одержимый бесами с давнего времени, и в одежду не одевавшийся, и живший не в доме, а в гробах.
LUKE|8|28|Он, увидев Иисуса, вскричал, пал пред Ним и громким голосом сказал: что Тебе до меня, Иисус, Сын Бога Всевышнего? умоляю Тебя, не мучь меня.
LUKE|8|29|Ибо [Иисус] повелел нечистому духу выйти из сего человека, потому что он долгое время мучил его, так что его связывали цепями и узами, сберегая его; но он разрывал узы и был гоним бесом в пустыни.
LUKE|8|30|Иисус спросил его: как тебе имя? Он сказал: легион, – потому что много бесов вошло в него.
LUKE|8|31|И они просили Иисуса, чтобы не повелел им идти в бездну.
LUKE|8|32|Тут же на горе паслось большое стадо свиней; и [бесы] просили Его, чтобы позволил им войти в них. Он позволил им.
LUKE|8|33|Бесы, выйдя из человека, вошли в свиней, и бросилось стадо с крутизны в озеро и потонуло.
LUKE|8|34|Пастухи, видя происшедшее, побежали и рассказали в городе и в селениях.
LUKE|8|35|И вышли видеть происшедшее; и, придя к Иисусу, нашли человека, из которого вышли бесы, сидящего у ног Иисуса, одетого и в здравом уме; и ужаснулись.
LUKE|8|36|Видевшие же рассказали им, как исцелился бесновавшийся.
LUKE|8|37|И просил Его весь народ Гадаринской окрестности удалиться от них, потому что они объяты были великим страхом. Он вошел в лодку и возвратился.
LUKE|8|38|Человек же, из которого вышли бесы, просил Его, чтобы быть с Ним. Но Иисус отпустил его, сказав:
LUKE|8|39|возвратись в дом твой и расскажи, что сотворил тебе Бог. Он пошел и проповедывал по всему городу, что сотворил ему Иисус.
LUKE|8|40|Когда же возвратился Иисус, народ принял Его, потому что все ожидали Его.
LUKE|8|41|И вот, пришел человек, именем Иаир, который был начальником синагоги; и, пав к ногам Иисуса, просил Его войти к нему в дом,
LUKE|8|42|потому что у него была одна дочь, лет двенадцати, и та была при смерти. Когда же Он шел, народ теснил Его.
LUKE|8|43|И женщина, страдавшая кровотечением двенадцать лет, которая, издержав на врачей все имение, ни одним не могла быть вылечена,
LUKE|8|44|подойдя сзади, коснулась края одежды Его; и тотчас течение крови у ней остановилось.
LUKE|8|45|И сказал Иисус: кто прикоснулся ко Мне? Когда же все отрицались, Петр сказал и бывшие с Ним: Наставник! народ окружает Тебя и теснит, – и Ты говоришь: кто прикоснулся ко Мне?
LUKE|8|46|Но Иисус сказал: прикоснулся ко Мне некто, ибо Я чувствовал силу, исшедшую из Меня.
LUKE|8|47|Женщина, видя, что она не утаилась, с трепетом подошла и, пав пред Ним, объявила Ему перед всем народом, по какой причине прикоснулась к Нему и как тотчас исцелилась.
LUKE|8|48|Он сказал ей: дерзай, дщерь! вера твоя спасла тебя; иди с миром.
LUKE|8|49|Когда Он еще говорил это, приходит некто из дома начальника синагоги и говорит ему: дочь твоя умерла; не утруждай Учителя.
LUKE|8|50|Но Иисус, услышав это, сказал ему: не бойся, только веруй, и спасена будет.
LUKE|8|51|Придя же в дом, не позволил войти никому, кроме Петра, Иоанна и Иакова, и отца девицы, и матери.
LUKE|8|52|Все плакали и рыдали о ней. Но Он сказал: не плачьте; она не умерла, но спит.
LUKE|8|53|И смеялись над Ним, зная, что она умерла.
LUKE|8|54|Он же, выслав всех вон и взяв ее за руку, возгласил: девица! встань.
LUKE|8|55|И возвратился дух ее; она тотчас встала, и Он велел дать ей есть.
LUKE|8|56|И удивились родители ее. Он же повелел им не сказывать никому о происшедшем.
LUKE|9|1|Созвав же двенадцать, дал силу и власть над всеми бесами и врачевать от болезней,
LUKE|9|2|и послал их проповедывать Царствие Божие и исцелять больных.
LUKE|9|3|И сказал им: ничего не берите на дорогу: ни посоха, ни сумы, ни хлеба, ни серебра, и не имейте по две одежды;
LUKE|9|4|и в какой дом войдете, там оставайтесь и оттуда отправляйтесь [в] [путь].
LUKE|9|5|А если где не примут вас, то, выходя из того города, отрясите и прах от ног ваших во свидетельство на них.
LUKE|9|6|Они пошли и проходили по селениям, благовествуя и исцеляя повсюду.
LUKE|9|7|Услышал Ирод четвертовластник о всем, что делал [Иисус], и недоумевал: ибо одни говорили, что это Иоанн восстал из мертвых;
LUKE|9|8|другие, что Илия явился, а иные, что один из древних пророков воскрес.
LUKE|9|9|И сказал Ирод: Иоанна я обезглавил; кто же Этот, о Котором я слышу такое? И искал увидеть Его.
LUKE|9|10|Апостолы, возвратившись, рассказали Ему, что они сделали; и Он, взяв их с Собою, удалился особо в пустое место, близ города, называемого Вифсаидою.
LUKE|9|11|Но народ, узнав, пошел за Ним; и Он, приняв их, беседовал с ними о Царствии Божием и требовавших исцеления исцелял.
LUKE|9|12|День же начал склоняться к вечеру. И, приступив к Нему, двенадцать говорили Ему: отпусти народ, чтобы они пошли в окрестные селения и деревни ночевать и достали пищи; потому что мы здесь в пустом месте.
LUKE|9|13|Но Он сказал им: вы дайте им есть. Они сказали: у нас нет более пяти хлебов и двух рыб; разве нам пойти купить пищи для всех сих людей?
LUKE|9|14|Ибо их было около пяти тысяч человек. Но Он сказал ученикам Своим: рассадите их рядами по пятидесяти.
LUKE|9|15|И сделали так, и рассадили всех.
LUKE|9|16|Он же, взяв пять хлебов и две рыбы и воззрев на небо, благословил их, преломил и дал ученикам, чтобы раздать народу.
LUKE|9|17|И ели, и насытились все; и оставшихся у них кусков набрано двенадцать коробов.
LUKE|9|18|В одно время, когда Он молился в уединенном месте, и ученики были с Ним, Он спросил их: за кого почитает Меня народ?
LUKE|9|19|Они сказали в ответ: за Иоанна Крестителя, а иные за Илию; другие же [говорят], что один из древних пророков воскрес.
LUKE|9|20|Он же спросил их: а вы за кого почитаете Меня? Отвечал Петр: за Христа Божия.
LUKE|9|21|Но Он строго приказал им никому не говорить о сем,
LUKE|9|22|сказав, что Сыну Человеческому должно много пострадать, и быть отвержену старейшинами, первосвященниками и книжниками, и быть убиту, и в третий день воскреснуть.
LUKE|9|23|Ко всем же сказал: если кто хочет идти за Мною, отвергнись себя, и возьми крест свой, и следуй за Мною.
LUKE|9|24|Ибо кто хочет душу свою сберечь, тот потеряет ее; а кто потеряет душу свою ради Меня, тот сбережет ее.
LUKE|9|25|Ибо что пользы человеку приобрести весь мир, а себя самого погубить или повредить себе?
LUKE|9|26|Ибо кто постыдится Меня и Моих слов, того Сын Человеческий постыдится, когда приидет во славе Своей и Отца и святых Ангелов.
LUKE|9|27|Говорю же вам истинно: есть некоторые из стоящих здесь, которые не вкусят смерти, как уже увидят Царствие Божие.
LUKE|9|28|После сих слов, дней через восемь, взяв Петра, Иоанна и Иакова, взошел Он на гору помолиться.
LUKE|9|29|И когда молился, вид лица Его изменился, и одежда Его сделалась белою, блистающею.
LUKE|9|30|И вот, два мужа беседовали с Ним, которые были Моисей и Илия;
LUKE|9|31|явившись во славе, они говорили об исходе Его, который Ему надлежало совершить в Иерусалиме.
LUKE|9|32|Петр же и бывшие с ним отягчены были сном; но, пробудившись, увидели славу Его и двух мужей, стоявших с Ним.
LUKE|9|33|И когда они отходили от Него, сказал Петр Иисусу: Наставник! хорошо нам здесь быть; сделаем три кущи: одну Тебе, одну Моисею и одну Илии, – не зная, что говорил.
LUKE|9|34|Когда же он говорил это, явилось облако и осенило их; и устрашились, когда вошли в облако.
LUKE|9|35|И был из облака глас, глаголющий: Сей есть Сын Мой Возлюбленный, Его слушайте.
LUKE|9|36|Когда был глас сей, остался Иисус один. И они умолчали, и никому не говорили в те дни о том, что видели.
LUKE|9|37|В следующий же день, когда они сошли с горы, встретило Его много народа.
LUKE|9|38|Вдруг некто из народа воскликнул: Учитель! умоляю Тебя взглянуть на сына моего, он один у меня:
LUKE|9|39|его схватывает дух, и он внезапно вскрикивает, и терзает его, так что он испускает пену; и насилу отступает от него, измучив его.
LUKE|9|40|Я просил учеников Твоих изгнать его, и они не могли.
LUKE|9|41|Иисус же, отвечая, сказал: о, род неверный и развращенный! доколе буду с вами и буду терпеть вас? приведи сюда сына твоего.
LUKE|9|42|Когда же тот еще шел, бес поверг его и стал бить; но Иисус запретил нечистому духу, и исцелил отрока, и отдал его отцу его.
LUKE|9|43|И все удивлялись величию Божию. Когда же все дивились всему, что творил Иисус, Он сказал ученикам Своим:
LUKE|9|44|вложите вы себе в уши слова сии: Сын Человеческий будет предан в руки человеческие.
LUKE|9|45|Но они не поняли слова сего, и оно было закрыто от них, так что они не постигли его, а спросить Его о сем слове боялись.
LUKE|9|46|Пришла же им мысль: кто бы из них был больше?
LUKE|9|47|Иисус же, видя помышление сердца их, взяв дитя, поставил его пред Собою
LUKE|9|48|и сказал им: кто примет сие дитя во имя Мое, тот Меня принимает; а кто примет Меня, тот принимает Пославшего Меня; ибо кто из вас меньше всех, тот будет велик.
LUKE|9|49|При сем Иоанн сказал: Наставник! мы видели человека, именем Твоим изгоняющего бесов, и запретили ему, потому что он не ходит с нами.
LUKE|9|50|Иисус сказал ему: не запрещайте, ибо кто не против вас, тот за вас.
LUKE|9|51|Когда же приближались дни взятия Его [от мира], Он восхотел идти в Иерусалим;
LUKE|9|52|и послал вестников пред лицем Своим; и они пошли и вошли в селение Самарянское; чтобы приготовить для Него;
LUKE|9|53|но [там] не приняли Его, потому что Он имел вид путешествующего в Иерусалим.
LUKE|9|54|Видя то, ученики Его, Иаков и Иоанн, сказали: Господи! хочешь ли, мы скажем, чтобы огонь сошел с неба и истребил их, как и Илия сделал?
LUKE|9|55|Но Он, обратившись к ним, запретил им и сказал: не знаете, какого вы духа;
LUKE|9|56|ибо Сын Человеческий пришел не губить души человеческие, а спасать. И пошли в другое селение.
LUKE|9|57|Случилось, что когда они были в пути, некто сказал Ему: Господи! я пойду за Тобою, куда бы Ты ни пошел.
LUKE|9|58|Иисус сказал ему: лисицы имеют норы, и птицы небесные – гнезда; а Сын Человеческий не имеет, где приклонить голову.
LUKE|9|59|А другому сказал: следуй за Мною. Тот сказал: Господи! позволь мне прежде пойти и похоронить отца моего.
LUKE|9|60|Но Иисус сказал ему: предоставь мертвым погребать своих мертвецов, а ты иди, благовествуй Царствие Божие.
LUKE|9|61|Еще другой сказал: я пойду за Тобою, Господи! но прежде позволь мне проститься с домашними моими.
LUKE|9|62|Но Иисус сказал ему: никто, возложивший руку свою на плуг и озирающийся назад, не благонадежен для Царствия Божия.
LUKE|10|1|После сего избрал Господь и других семьдесят [учеников], и послал их по два пред лицем Своим во всякий город и место, куда Сам хотел идти,
LUKE|10|2|и сказал им: жатвы много, а делателей мало; итак, молите Господина жатвы, чтобы выслал делателей на жатву Свою.
LUKE|10|3|Идите! Я посылаю вас, как агнцев среди волков.
LUKE|10|4|Не берите ни мешка, ни сумы, ни обуви, и никого на дороге не приветствуйте.
LUKE|10|5|В какой дом войдете, сперва говорите: мир дому сему;
LUKE|10|6|и если будет там сын мира, то почиет на нем мир ваш, а если нет, то к вам возвратится.
LUKE|10|7|В доме же том оставайтесь, ешьте и пейте, что у них есть, ибо трудящийся достоин награды за труды свои; не переходите из дома в дом.
LUKE|10|8|И если придете в какой город и примут вас, ешьте, что вам предложат,
LUKE|10|9|и исцеляйте находящихся в нем больных, и говорите им: приблизилось к вам Царствие Божие.
LUKE|10|10|Если же придете в какой город и не примут вас, то, выйдя на улицу, скажите:
LUKE|10|11|и прах, прилипший к нам от вашего города, отрясаем вам; однако же знайте, что приблизилось к вам Царствие Божие.
LUKE|10|12|Сказываю вам, что Содому в день оный будет отраднее, нежели городу тому.
LUKE|10|13|Горе тебе, Хоразин! горе тебе, Вифсаида! ибо если бы в Тире и Сидоне явлены были силы, явленные в вас, то давно бы они, сидя во вретище и пепле, покаялись;
LUKE|10|14|но и Тиру и Сидону отраднее будет на суде, нежели вам.
LUKE|10|15|И ты, Капернаум, до неба вознесшийся, до ада низвергнешься.
LUKE|10|16|Слушающий вас Меня слушает, и отвергающийся вас Меня отвергается; а отвергающийся Меня отвергается Пославшего Меня.
LUKE|10|17|Семьдесят [учеников] возвратились с радостью и говорили: Господи! и бесы повинуются нам о имени Твоем.
LUKE|10|18|Он же сказал им: Я видел сатану, спадшего с неба, как молнию;
LUKE|10|19|се, даю вам власть наступать на змей и скорпионов и на всю силу вражью, и ничто не повредит вам;
LUKE|10|20|однакож тому не радуйтесь, что духи вам повинуются, но радуйтесь тому, что имена ваши написаны на небесах.
LUKE|10|21|В тот час возрадовался духом Иисус и сказал: славлю Тебя, Отче, Господи неба и земли, что Ты утаил сие от мудрых и разумных и открыл младенцам. Ей, Отче! Ибо таково было Твое благоволение.
LUKE|10|22|И, обратившись к ученикам, сказал: все предано Мне Отцем Моим; и кто есть Сын, не знает никто, кроме Отца, и кто есть Отец, [не знает] [никто], кроме Сына, и кому Сын хочет открыть.
LUKE|10|23|И, обратившись к ученикам, сказал им особо: блаженны очи, видящие то, что вы видите!
LUKE|10|24|ибо сказываю вам, что многие пророки и цари желали видеть, что вы видите, и не видели, и слышать, что вы слышите, и не слышали.
LUKE|10|25|И вот, один законник встал и, искушая Его, сказал: Учитель! что мне делать, чтобы наследовать жизнь вечную?
LUKE|10|26|Он же сказал ему: в законе что написано? как читаешь?
LUKE|10|27|Он сказал в ответ: возлюби Господа Бога твоего всем сердцем твоим, и всею душею твоею, и всею крепостию твоею, и всем разумением твоим, и ближнего твоего, как самого себя.
LUKE|10|28|[Иисус] сказал ему: правильно ты отвечал; так поступай, и будешь жить.
LUKE|10|29|Но он, желая оправдать себя, сказал Иисусу: а кто мой ближний?
LUKE|10|30|На это сказал Иисус: некоторый человек шел из Иерусалима в Иерихон и попался разбойникам, которые сняли с него одежду, изранили его и ушли, оставив его едва живым.
LUKE|10|31|По случаю один священник шел тою дорогою и, увидев его, прошел мимо.
LUKE|10|32|Также и левит, быв на том месте, подошел, посмотрел и прошел мимо.
LUKE|10|33|Самарянин же некто, проезжая, нашел на него и, увидев его, сжалился
LUKE|10|34|и, подойдя, перевязал ему раны, возливая масло и вино; и, посадив его на своего осла, привез его в гостиницу и позаботился о нем;
LUKE|10|35|а на другой день, отъезжая, вынул два динария, дал содержателю гостиницы и сказал ему: позаботься о нем; и если издержишь что более, я, когда возвращусь, отдам тебе.
LUKE|10|36|Кто из этих троих, думаешь ты, был ближний попавшемуся разбойникам?
LUKE|10|37|Он сказал: оказавший ему милость. Тогда Иисус сказал ему: иди, и ты поступай так же.
LUKE|10|38|В продолжение пути их пришел Он в одно селение; здесь женщина, именем Марфа, приняла Его в дом свой;
LUKE|10|39|у нее была сестра, именем Мария, которая села у ног Иисуса и слушала слово Его.
LUKE|10|40|Марфа же заботилась о большом угощении и, подойдя, сказала: Господи! или Тебе нужды нет, что сестра моя одну меня оставила служить? скажи ей, чтобы помогла мне.
LUKE|10|41|Иисус же сказал ей в ответ: Марфа! Марфа! ты заботишься и суетишься о многом,
LUKE|10|42|а одно только нужно; Мария же избрала благую часть, которая не отнимется у нее.
LUKE|11|1|Случилось, что когда Он в одном месте молился, и перестал, один из учеников Его сказал Ему: Господи! научи нас молиться, как и Иоанн научил учеников своих.
LUKE|11|2|Он сказал им: когда молитесь, говорите: Отче наш, сущий на небесах! да святится имя Твое; да приидет Царствие Твое; да будет воля Твоя и на земле, как на небе;
LUKE|11|3|хлеб наш насущный подавай нам на каждый день;
LUKE|11|4|и прости нам грехи наши, ибо и мы прощаем всякому должнику нашему; и не введи нас в искушение, но избавь нас от лукавого.
LUKE|11|5|И сказал им: [положим, что] кто–нибудь из вас, имея друга, придет к нему в полночь и скажет ему: друг! дай мне взаймы три хлеба,
LUKE|11|6|ибо друг мой с дороги зашел ко мне, и мне нечего предложить ему;
LUKE|11|7|а тот изнутри скажет ему в ответ: не беспокой меня, двери уже заперты, и дети мои со мною на постели; не могу встать и дать тебе.
LUKE|11|8|Если, говорю вам, он не встанет и не даст ему по дружбе с ним, то по неотступности его, встав, даст ему, сколько просит.
LUKE|11|9|И Я скажу вам: просите, и дано будет вам; ищите, и найдете; стучите, и отворят вам,
LUKE|11|10|ибо всякий просящий получает, и ищущий находит, и стучащему отворят.
LUKE|11|11|Какой из вас отец, [когда] сын попросит у него хлеба, подаст ему камень? или, [когда попросит] рыбы, подаст ему змею вместо рыбы?
LUKE|11|12|Или, если попросит яйца, подаст ему скорпиона?
LUKE|11|13|Итак, если вы, будучи злы, умеете даяния благие давать детям вашим, тем более Отец Небесный даст Духа Святаго просящим у Него.
LUKE|11|14|Однажды изгнал Он беса, который был нем; и когда бес вышел, немой стал говорить; и народ удивился.
LUKE|11|15|Некоторые же из них говорили: Он изгоняет бесов силою веельзевула, князя бесовского.
LUKE|11|16|А другие, искушая, требовали от Него знамения с неба.
LUKE|11|17|Но Он, зная помышления их, сказал им: всякое царство, разделившееся само в себе, опустеет, и дом, [разделившийся] сам в себе, падет;
LUKE|11|18|если же и сатана разделится сам в себе, то как устоит царство его? а вы говорите, что Я силою веельзевула изгоняю бесов;
LUKE|11|19|и если Я силою веельзевула изгоняю бесов, то сыновья ваши чьею силою изгоняют их? Посему они будут вам судьями.
LUKE|11|20|Если же Я перстом Божиим изгоняю бесов, то, конечно, достигло до вас Царствие Божие.
LUKE|11|21|Когда сильный с оружием охраняет свой дом, тогда в безопасности его имение;
LUKE|11|22|когда же сильнейший его нападет на него и победит его, тогда возьмет все оружие его, на которое он надеялся, и разделит похищенное у него.
LUKE|11|23|Кто не со Мною, тот против Меня; и кто не собирает со Мною, тот расточает.
LUKE|11|24|Когда нечистый дух выйдет из человека, то ходит по безводным местам, ища покоя, и, не находя, говорит: возвращусь в дом мой, откуда вышел;
LUKE|11|25|и, придя, находит его выметенным и убранным;
LUKE|11|26|тогда идет и берет с собою семь других духов, злейших себя, и, войдя, живут там, – и бывает для человека того последнее хуже первого.
LUKE|11|27|Когда же Он говорил это, одна женщина, возвысив голос из народа, сказала Ему: блаженно чрево, носившее Тебя, и сосцы, Тебя питавшие!
LUKE|11|28|А Он сказал: блаженны слышащие слово Божие и соблюдающие его.
LUKE|11|29|Когда же народ стал сходиться во множестве, Он начал говорить: род сей лукав, он ищет знамения, и знамение не дастся ему, кроме знамения Ионы пророка;
LUKE|11|30|ибо как Иона был знамением для Ниневитян, так будет и Сын Человеческий для рода сего.
LUKE|11|31|Царица южная восстанет на суд с людьми рода сего и осудит их, ибо она приходила от пределов земли послушать мудрости Соломоновой; и вот, здесь больше Соломона.
LUKE|11|32|Ниневитяне восстанут на суд с родом сим и осудят его, ибо они покаялись от проповеди Иониной, и вот, здесь больше Ионы.
LUKE|11|33|Никто, зажегши свечу, не ставит ее в сокровенном месте, ни под сосудом, но на подсвечнике, чтобы входящие видели свет.
LUKE|11|34|Светильник тела есть око; итак, если око твое будет чисто, то и все тело твое будет светло; а если оно будет худо, то и тело твое будет темно.
LUKE|11|35|Итак, смотри: свет, который в тебе, не есть ли тьма?
LUKE|11|36|Если же тело твое все светло и не имеет ни одной темной части, то будет светло все так, как бы светильник освещал тебя сиянием.
LUKE|11|37|Когда Он говорил это, один фарисей просил Его к себе обедать. Он пришел и возлег.
LUKE|11|38|Фарисей же удивился, увидев, что Он не умыл [рук] перед обедом.
LUKE|11|39|Но Господь сказал ему: ныне вы, фарисеи, внешность чаши и блюда очищаете, а внутренность ваша исполнена хищения и лукавства.
LUKE|11|40|Неразумные! не Тот же ли, Кто сотворил внешнее, сотворил и внутреннее?
LUKE|11|41|Подавайте лучше милостыню из того, что у вас есть, тогда все будет у вас чисто.
LUKE|11|42|Но горе вам, фарисеям, что даете десятину с мяты, руты и всяких овощей, и нерадите о суде и любви Божией: сие надлежало делать, и того не оставлять.
LUKE|11|43|Горе вам, фарисеям, что любите председания в синагогах и приветствия в народных собраниях.
LUKE|11|44|Горе вам, книжники и фарисеи, лицемеры, что вы – как гробы скрытые, над которыми люди ходят и не знают того.
LUKE|11|45|На это некто из законников сказал Ему: Учитель! говоря это, Ты и нас обижаешь.
LUKE|11|46|Но Он сказал: и вам, законникам, горе, что налагаете на людей бремена неудобоносимые, а сами и одним перстом своим не дотрагиваетесь до них.
LUKE|11|47|Горе вам, что строите гробницы пророкам, которых избили отцы ваши:
LUKE|11|48|сим вы свидетельствуете о делах отцов ваших и соглашаетесь с ними, ибо они избили пророков, а вы строите им гробницы.
LUKE|11|49|Потому и премудрость Божия сказала: пошлю к ним пророков и Апостолов, и из них одних убьют, а других изгонят,
LUKE|11|50|да взыщется от рода сего кровь всех пророков, пролитая от создания мира,
LUKE|11|51|от крови Авеля до крови Захарии, убитого между жертвенником и храмом. Ей, говорю вам, взыщется от рода сего.
LUKE|11|52|Горе вам, законникам, что вы взяли ключ разумения: сами не вошли, и входящим воспрепятствовали.
LUKE|11|53|Когда Он говорил им это, книжники и фарисеи начали сильно приступать к Нему, вынуждая у Него ответы на многое,
LUKE|11|54|подыскиваясь под Него и стараясь уловить что–нибудь из уст Его, чтобы обвинить Его.
LUKE|12|1|Между тем, когда собрались тысячи народа, так что теснили друг друга, Он начал говорить сперва ученикам Своим: берегитесь закваски фарисейской, которая есть лицемерие.
LUKE|12|2|Нет ничего сокровенного, что не открылось бы, и тайного, чего не узнали бы.
LUKE|12|3|Посему, что вы сказали в темноте, то услышится во свете; и что говорили на ухо внутри дома, то будет провозглашено на кровлях.
LUKE|12|4|Говорю же вам, друзьям Моим: не бойтесь убивающих тело и потом не могущих ничего более сделать;
LUKE|12|5|но скажу вам, кого бояться: бойтесь того, кто, по убиении, может ввергнуть в геенну: ей, говорю вам, того бойтесь.
LUKE|12|6|Не пять ли малых птиц продаются за два ассария? и ни одна из них не забыта у Бога.
LUKE|12|7|А у вас и волосы на голове все сочтены. Итак не бойтесь: вы дороже многих малых птиц.
LUKE|12|8|Сказываю же вам: всякого, кто исповедает Меня пред человеками, и Сын Человеческий исповедает пред Ангелами Божиими;
LUKE|12|9|а кто отвергнется Меня пред человеками, тот отвержен будет пред Ангелами Божиими.
LUKE|12|10|И всякому, кто скажет слово на Сына Человеческого, прощено будет; а кто скажет хулу на Святаго Духа, тому не простится.
LUKE|12|11|Когда же приведут вас в синагоги, к начальствам и властям, не заботьтесь, как или что отвечать, или что говорить,
LUKE|12|12|ибо Святый Дух научит вас в тот час, что должно говорить.
LUKE|12|13|Некто из народа сказал Ему: Учитель! скажи брату моему, чтобы он разделил со мною наследство.
LUKE|12|14|Он же сказал человеку тому: кто поставил Меня судить или делить вас?
LUKE|12|15|При этом сказал им: смотрите, берегитесь любостяжания, ибо жизнь человека не зависит от изобилия его имения.
LUKE|12|16|И сказал им притчу: у одного богатого человека был хороший урожай в поле;
LUKE|12|17|и он рассуждал сам с собою: что мне делать? некуда мне собрать плодов моих?
LUKE|12|18|И сказал: вот что сделаю: сломаю житницы мои и построю большие, и соберу туда весь хлеб мой и все добро мое,
LUKE|12|19|и скажу душе моей: душа! много добра лежит у тебя на многие годы: покойся, ешь, пей, веселись.
LUKE|12|20|Но Бог сказал ему: безумный! в сию ночь душу твою возьмут у тебя; кому же достанется то, что ты заготовил?
LUKE|12|21|Так [бывает с тем], кто собирает сокровища для себя, а не в Бога богатеет.
LUKE|12|22|И сказал ученикам Своим: посему говорю вам, – не заботьтесь для души вашей, что вам есть, ни для тела, во что одеться:
LUKE|12|23|душа больше пищи, и тело – одежды.
LUKE|12|24|Посмотрите на воронов: они не сеют, не жнут; нет у них ни хранилищ, ни житниц, и Бог питает их; сколько же вы лучше птиц?
LUKE|12|25|Да и кто из вас, заботясь, может прибавить себе роста хотя на один локоть?
LUKE|12|26|Итак, если и малейшего сделать не можете, что заботитесь о прочем?
LUKE|12|27|Посмотрите на лилии, как они растут: не трудятся, не прядут; но говорю вам, что и Соломон во всей славе своей не одевался так, как всякая из них.
LUKE|12|28|Если же траву на поле, которая сегодня есть, а завтра будет брошена в печь, Бог так одевает, то кольми паче вас, маловеры!
LUKE|12|29|Итак, не ищите, что вам есть, или что пить, и не беспокойтесь,
LUKE|12|30|потому что всего этого ищут люди мира сего; ваш же Отец знает, что вы имеете нужду в том;
LUKE|12|31|наипаче ищите Царствия Божия, и это все приложится вам.
LUKE|12|32|Не бойся, малое стадо! ибо Отец ваш благоволил дать вам Царство.
LUKE|12|33|Продавайте имения ваши и давайте милостыню. Приготовляйте себе влагалища не ветшающие, сокровище неоскудевающее на небесах, куда вор не приближается и где моль не съедает,
LUKE|12|34|ибо где сокровище ваше, там и сердце ваше будет.
LUKE|12|35|Да будут чресла ваши препоясаны и светильники горящи.
LUKE|12|36|И вы будьте подобны людям, ожидающим возвращения господина своего с брака, дабы, когда придет и постучит, тотчас отворить ему.
LUKE|12|37|Блаженны рабы те, которых господин, придя, найдет бодрствующими; истинно говорю вам, он препояшется и посадит их, и, подходя, станет служить им.
LUKE|12|38|И если придет во вторую стражу, и в третью стражу придет, и найдет их так, то блаженны рабы те.
LUKE|12|39|Вы знаете, что если бы ведал хозяин дома, в который час придет вор, то бодрствовал бы и не допустил бы подкопать дом свой.
LUKE|12|40|Будьте же и вы готовы, ибо, в который час не думаете, приидет Сын Человеческий.
LUKE|12|41|Тогда сказал Ему Петр: Господи! к нам ли притчу сию говоришь, или и ко всем?
LUKE|12|42|Господь же сказал: кто верный и благоразумный домоправитель, которого господин поставил над слугами своими раздавать им в свое время меру хлеба?
LUKE|12|43|Блажен раб тот, которого господин его, придя, найдет поступающим так.
LUKE|12|44|Истинно говорю вам, что над всем имением своим поставит его.
LUKE|12|45|Если же раб тот скажет в сердце своем: не скоро придет господин мой, и начнет бить слуг и служанок, есть и пить и напиваться, –
LUKE|12|46|то придет господин раба того в день, в который он не ожидает, и в час, в который не думает, и рассечет его, и подвергнет его одной участи с неверными.
LUKE|12|47|Раб же тот, который знал волю господина своего, и не был готов, и не делал по воле его, бит будет много;
LUKE|12|48|а который не знал, и сделал достойное наказания, бит будет меньше. И от всякого, кому дано много, много и потребуется, и кому много вверено, с того больше взыщут.
LUKE|12|49|Огонь пришел Я низвести на землю, и как желал бы, чтобы он уже возгорелся!
LUKE|12|50|Крещением должен Я креститься; и как Я томлюсь, пока сие совершится!
LUKE|12|51|Думаете ли вы, что Я пришел дать мир земле? Нет, говорю вам, но разделение;
LUKE|12|52|ибо отныне пятеро в одном доме станут разделяться, трое против двух, и двое против трех:
LUKE|12|53|отец будет против сына, и сын против отца; мать против дочери, и дочь против матери; свекровь против невестки своей, и невестка против свекрови своей.
LUKE|12|54|Сказал же и народу: когда вы видите облако, поднимающееся с запада, тотчас говорите: дождь будет, и бывает так;
LUKE|12|55|и когда дует южный ветер, говорите: зной будет, и бывает.
LUKE|12|56|Лицемеры! лице земли и неба распознавать умеете, как же времени сего не узнаете?
LUKE|12|57|Зачем же вы и по самим себе не судите, чему быть должно?
LUKE|12|58|Когда ты идешь с соперником своим к начальству, то на дороге постарайся освободиться от него, чтобы он не привел тебя к судье, а судья не отдал тебя истязателю, а истязатель не вверг тебя в темницу;
LUKE|12|59|Сказываю тебе: не выйдешь оттуда, пока не отдашь и последней полушки.
LUKE|13|1|В это время пришли некоторые и рассказали Ему о Галилеянах, которых кровь Пилат смешал с жертвами их.
LUKE|13|2|Иисус сказал им на это: думаете ли вы, что эти Галилеяне были грешнее всех Галилеян, что так пострадали?
LUKE|13|3|Нет, говорю вам, но, если не покаетесь, все так же погибнете.
LUKE|13|4|Или думаете ли, что те восемнадцать человек, на которых упала башня Силоамская и побила их, виновнее были всех, живущих в Иерусалиме?
LUKE|13|5|Нет, говорю вам, но, если не покаетесь, все так же погибнете.
LUKE|13|6|И сказал сию притчу: некто имел в винограднике своем посаженную смоковницу, и пришел искать плода на ней, и не нашел;
LUKE|13|7|и сказал виноградарю: вот, я третий год прихожу искать плода на этой смоковнице и не нахожу; сруби ее: на что она и землю занимает?
LUKE|13|8|Но он сказал ему в ответ: господин! оставь ее и на этот год, пока я окопаю ее и обложу навозом, –
LUKE|13|9|не принесет ли плода; если же нет, то в следующий [год] срубишь ее.
LUKE|13|10|В одной из синагог учил Он в субботу.
LUKE|13|11|Там была женщина, восемнадцать лет имевшая духа немощи: она была скорчена и не могла выпрямиться.
LUKE|13|12|Иисус, увидев ее, подозвал и сказал ей: женщина! ты освобождаешься от недуга твоего.
LUKE|13|13|И возложил на нее руки, и она тотчас выпрямилась и стала славить Бога.
LUKE|13|14|При этом начальник синагоги, негодуя, что Иисус исцелил в субботу, сказал народу: есть шесть дней, в которые должно делать; в те и приходите исцеляться, а не в день субботний.
LUKE|13|15|Господь сказал ему в ответ: лицемер! не отвязывает ли каждый из вас вола своего или осла от яслей в субботу и не ведет ли поить?
LUKE|13|16|сию же дочь Авраамову, которую связал сатана вот уже восемнадцать лет, не надлежало ли освободить от уз сих в день субботний?
LUKE|13|17|И когда говорил Он это, все противившиеся Ему стыдились; и весь народ радовался о всех славных делах Его.
LUKE|13|18|Он же сказал: чему подобно Царствие Божие? и чему уподоблю его?
LUKE|13|19|Оно подобно зерну горчичному, которое, взяв, человек посадил в саду своем; и выросло, и стало большим деревом, и птицы небесные укрывались в ветвях его.
LUKE|13|20|Еще сказал: чему уподоблю Царствие Божие?
LUKE|13|21|Оно подобно закваске, которую женщина, взяв, положила в три меры муки, доколе не вскисло все.
LUKE|13|22|И проходил по городам и селениям, уча и направляя путь к Иерусалиму.
LUKE|13|23|Некто сказал Ему: Господи! неужели мало спасающихся? Он же сказал им:
LUKE|13|24|подвизайтесь войти сквозь тесные врата, ибо, сказываю вам, многие поищут войти, и не возмогут.
LUKE|13|25|Когда хозяин дома встанет и затворит двери, тогда вы, стоя вне, станете стучать в двери и говорить: Господи! Господи! отвори нам; но Он скажет вам в ответ: не знаю вас, откуда вы.
LUKE|13|26|Тогда станете говорить: мы ели и пили пред Тобою, и на улицах наших учил Ты.
LUKE|13|27|Но Он скажет: говорю вам: не знаю вас, откуда вы; отойдите от Меня все делатели неправды.
LUKE|13|28|Там будет плач и скрежет зубов, когда увидите Авраама, Исаака и Иакова и всех пророков в Царствии Божием, а себя изгоняемыми вон.
LUKE|13|29|И придут от востока и запада, и севера и юга, и возлягут в Царствии Божием.
LUKE|13|30|И вот, есть последние, которые будут первыми, и есть первые, которые будут последними.
LUKE|13|31|В тот день пришли некоторые из фарисеев и говорили Ему: выйди и удались отсюда, ибо Ирод хочет убить Тебя.
LUKE|13|32|И сказал им: пойдите, скажите этой лисице: се, изгоняю бесов и совершаю исцеления сегодня и завтра, и в третий [день] кончу;
LUKE|13|33|а впрочем, Мне должно ходить сегодня, завтра и в последующий день, потому что не бывает, чтобы пророк погиб вне Иерусалима.
LUKE|13|34|Иерусалим! Иерусалим! избивающий пророков и камнями побивающий посланных к тебе! сколько раз хотел Я собрать чад твоих, как птица птенцов своих под крылья, и вы не захотели!
LUKE|13|35|Се, оставляется вам дом ваш пуст. Сказываю же вам, что вы не увидите Меня, пока не придет время, когда скажете: благословен Грядый во имя Господне!
LUKE|14|1|Случилось Ему в субботу придти в дом одного из начальников фарисейских вкусить хлеба, и они наблюдали за Ним.
LUKE|14|2|И вот, предстал пред Него человек, страждущий водяною болезнью.
LUKE|14|3|По сему случаю Иисус спросил законников и фарисеев: позволительно ли врачевать в субботу?
LUKE|14|4|Они молчали. И, прикоснувшись, исцелил его и отпустил.
LUKE|14|5|При сем сказал им: если у кого из вас осел или вол упадет в колодезь, не тотчас ли вытащит его и в субботу?
LUKE|14|6|И не могли отвечать Ему на это.
LUKE|14|7|Замечая же, как званые выбирали первые места, сказал им притчу:
LUKE|14|8|когда ты будешь позван кем на брак, не садись на первое место, чтобы не случился кто из званых им почетнее тебя,
LUKE|14|9|и звавший тебя и его, подойдя, не сказал бы тебе: уступи ему место; и тогда со стыдом должен будешь занять последнее место.
LUKE|14|10|Но когда зван будешь, придя, садись на последнее место, чтобы звавший тебя, подойдя, сказал: друг! пересядь выше; тогда будет тебе честь пред сидящими с тобою,
LUKE|14|11|ибо всякий возвышающий сам себя унижен будет, а унижающий себя возвысится.
LUKE|14|12|Сказал же и позвавшему Его: когда делаешь обед или ужин, не зови друзей твоих, ни братьев твоих, ни родственников твоих, ни соседей богатых, чтобы и они тебя когда не позвали, и не получил ты воздаяния.
LUKE|14|13|Но, когда делаешь пир, зови нищих, увечных, хромых, слепых,
LUKE|14|14|и блажен будешь, что они не могут воздать тебе, ибо воздастся тебе в воскресение праведных.
LUKE|14|15|Услышав это, некто из возлежащих с Ним сказал Ему: блажен, кто вкусит хлеба в Царствии Божием!
LUKE|14|16|Он же сказал ему: один человек сделал большой ужин и звал многих,
LUKE|14|17|и когда наступило время ужина, послал раба своего сказать званым: идите, ибо уже все готово.
LUKE|14|18|И начали все, как бы сговорившись, извиняться. Первый сказал ему: я купил землю и мне нужно пойти посмотреть ее; прошу тебя, извини меня.
LUKE|14|19|Другой сказал: я купил пять пар волов и иду испытать их; прошу тебя, извини меня.
LUKE|14|20|Третий сказал: я женился и потому не могу придти.
LUKE|14|21|И, возвратившись, раб тот донес о сем господину своему. Тогда, разгневавшись, хозяин дома сказал рабу своему: пойди скорее по улицам и переулкам города и приведи сюда нищих, увечных, хромых и слепых.
LUKE|14|22|И сказал раб: господин! исполнено, как приказал ты, и еще есть место.
LUKE|14|23|Господин сказал рабу: пойди по дорогам и изгородям и убеди придти, чтобы наполнился дом мой.
LUKE|14|24|Ибо сказываю вам, что никто из тех званых не вкусит моего ужина, ибо много званых, но мало избранных.
LUKE|14|25|С Ним шло множество народа; и Он, обратившись, сказал им:
LUKE|14|26|если кто приходит ко Мне и не возненавидит отца своего и матери, и жены и детей, и братьев и сестер, а притом и самой жизни своей, тот не может быть Моим учеником;
LUKE|14|27|и кто не несет креста своего и идет за Мною, не может быть Моим учеником.
LUKE|14|28|Ибо кто из вас, желая построить башню, не сядет прежде и не вычислит издержек, имеет ли он, что нужно для совершения ее,
LUKE|14|29|дабы, когда положит основание и не возможет совершить, все видящие не стали смеяться над ним,
LUKE|14|30|говоря: этот человек начал строить и не мог окончить?
LUKE|14|31|Или какой царь, идя на войну против другого царя, не сядет и не посоветуется прежде, силен ли он с десятью тысячами противостать идущему на него с двадцатью тысячами?
LUKE|14|32|Иначе, пока тот еще далеко, он пошлет к нему посольство просить о мире.
LUKE|14|33|Так всякий из вас, кто не отрешится от всего, что имеет, не может быть Моим учеником.
LUKE|14|34|Соль – добрая вещь; но если соль потеряет силу, чем исправить ее?
LUKE|14|35|ни в землю, ни в навоз не годится; вон выбрасывают ее. Кто имеет уши слышать, да слышит!
LUKE|15|1|Приближались к Нему все мытари и грешники слушать Его.
LUKE|15|2|Фарисеи же и книжники роптали, говоря: Он принимает грешников и ест с ними.
LUKE|15|3|Но Он сказал им следующую притчу:
LUKE|15|4|кто из вас, имея сто овец и потеряв одну из них, не оставит девяноста девяти в пустыне и не пойдет за пропавшею, пока не найдет ее?
LUKE|15|5|А найдя, возьмет ее на плечи свои с радостью
LUKE|15|6|и, придя домой, созовет друзей и соседей и скажет им: порадуйтесь со мною: я нашел мою пропавшую овцу.
LUKE|15|7|Сказываю вам, что так на небесах более радости будет об одном грешнике кающемся, нежели о девяноста девяти праведниках, не имеющих нужды в покаянии.
LUKE|15|8|Или какая женщина, имея десять драхм, если потеряет одну драхму, не зажжет свечи и не станет мести комнату и искать тщательно, пока не найдет,
LUKE|15|9|а найдя, созовет подруг и соседок и скажет: порадуйтесь со мною: я нашла потерянную драхму.
LUKE|15|10|Так, говорю вам, бывает радость у Ангелов Божиих и об одном грешнике кающемся.
LUKE|15|11|Еще сказал: у некоторого человека было два сына;
LUKE|15|12|и сказал младший из них отцу: отче! дай мне следующую [мне] часть имения. И [отец] разделил им имение.
LUKE|15|13|По прошествии немногих дней младший сын, собрав все, пошел в дальнюю сторону и там расточил имение свое, живя распутно.
LUKE|15|14|Когда же он прожил все, настал великий голод в той стране, и он начал нуждаться;
LUKE|15|15|и пошел, пристал к одному из жителей страны той, а тот послал его на поля свои пасти свиней;
LUKE|15|16|и он рад был наполнить чрево свое рожками, которые ели свиньи, но никто не давал ему.
LUKE|15|17|Придя же в себя, сказал: сколько наемников у отца моего избыточествуют хлебом, а я умираю от голода;
LUKE|15|18|встану, пойду к отцу моему и скажу ему: отче! я согрешил против неба и пред тобою
LUKE|15|19|и уже недостоин называться сыном твоим; прими меня в число наемников твоих.
LUKE|15|20|Встал и пошел к отцу своему. И когда он был еще далеко, увидел его отец его и сжалился; и, побежав, пал ему на шею и целовал его.
LUKE|15|21|Сын же сказал ему: отче! я согрешил против неба и пред тобою и уже недостоин называться сыном твоим.
LUKE|15|22|А отец сказал рабам своим: принесите лучшую одежду и оденьте его, и дайте перстень на руку его и обувь на ноги;
LUKE|15|23|и приведите откормленного теленка, и заколите; станем есть и веселиться!
LUKE|15|24|ибо этот сын мой был мертв и ожил, пропадал и нашелся. И начали веселиться.
LUKE|15|25|Старший же сын его был на поле; и возвращаясь, когда приблизился к дому, услышал пение и ликование;
LUKE|15|26|и, призвав одного из слуг, спросил: что это такое?
LUKE|15|27|Он сказал ему: брат твой пришел, и отец твой заколол откормленного теленка, потому что принял его здоровым.
LUKE|15|28|Он осердился и не хотел войти. Отец же его, выйдя, звал его.
LUKE|15|29|Но он сказал в ответ отцу: вот, я столько лет служу тебе и никогда не преступал приказания твоего, но ты никогда не дал мне и козленка, чтобы мне повеселиться с друзьями моими;
LUKE|15|30|а когда этот сын твой, расточивший имение свое с блудницами, пришел, ты заколол для него откормленного теленка.
LUKE|15|31|Он же сказал ему: сын мой! ты всегда со мною, и все мое твое,
LUKE|15|32|а о том надобно было радоваться и веселиться, что брат твой сей был мертв и ожил, пропадал и нашелся.
LUKE|16|1|Сказал же и к ученикам Своим: один человек был богат и имел управителя, на которого донесено было ему, что расточает имение его;
LUKE|16|2|и, призвав его, сказал ему: что это я слышу о тебе? дай отчет в управлении твоем, ибо ты не можешь более управлять.
LUKE|16|3|Тогда управитель сказал сам в себе: что мне делать? господин мой отнимает у меня управление домом; копать не могу, просить стыжусь;
LUKE|16|4|знаю, что сделать, чтобы приняли меня в домы свои, когда отставлен буду от управления домом.
LUKE|16|5|И, призвав должников господина своего, каждого порознь, сказал первому: сколько ты должен господину моему?
LUKE|16|6|Он сказал: сто мер масла. И сказал ему: возьми твою расписку и садись скорее, напиши: пятьдесят.
LUKE|16|7|Потом другому сказал: а ты сколько должен? Он отвечал: сто мер пшеницы. И сказал ему: возьми твою расписку и напиши: восемьдесят.
LUKE|16|8|И похвалил господин управителя неверного, что догадливо поступил; ибо сыны века сего догадливее сынов света в своем роде.
LUKE|16|9|И Я говорю вам: приобретайте себе друзей богатством неправедным, чтобы они, когда обнищаете, приняли вас в вечные обители.
LUKE|16|10|Верный в малом и во многом верен, а неверный в малом неверен и во многом.
LUKE|16|11|Итак, если вы в неправедном богатстве не были верны, кто поверит вам истинное?
LUKE|16|12|И если в чужом не были верны, кто даст вам ваше?
LUKE|16|13|Никакой слуга не может служить двум господам, ибо или одного будет ненавидеть, а другого любить, или одному станет усердствовать, а о другом нерадеть. Не можете служить Богу и маммоне.
LUKE|16|14|Слышали все это и фарисеи, которые были сребролюбивы, и они смеялись над Ним.
LUKE|16|15|Он сказал им: вы выказываете себя праведниками пред людьми, но Бог знает сердца ваши, ибо что высоко у людей, то мерзость пред Богом.
LUKE|16|16|Закон и пророки до Иоанна; с сего времени Царствие Божие благовествуется, и всякий усилием входит в него.
LUKE|16|17|Но скорее небо и земля прейдут, нежели одна черта из закона пропадет.
LUKE|16|18|Всякий, разводящийся с женою своею и женящийся на другой, прелюбодействует, и всякий, женящийся на разведенной с мужем, прелюбодействует.
LUKE|16|19|Некоторый человек был богат, одевался в порфиру и виссон и каждый день пиршествовал блистательно.
LUKE|16|20|Был также некоторый нищий, именем Лазарь, который лежал у ворот его в струпьях
LUKE|16|21|и желал напитаться крошками, падающими со стола богача, и псы, приходя, лизали струпья его.
LUKE|16|22|Умер нищий и отнесен был Ангелами на лоно Авраамово. Умер и богач, и похоронили его.
LUKE|16|23|И в аде, будучи в муках, он поднял глаза свои, увидел вдали Авраама и Лазаря на лоне его
LUKE|16|24|и, возопив, сказал: отче Аврааме! умилосердись надо мною и пошли Лазаря, чтобы омочил конец перста своего в воде и прохладил язык мой, ибо я мучаюсь в пламени сем.
LUKE|16|25|Но Авраам сказал: чадо! вспомни, что ты получил уже доброе твое в жизни твоей, а Лазарь – злое; ныне же он здесь утешается, а ты страдаешь;
LUKE|16|26|и сверх всего того между нами и вами утверждена великая пропасть, так что хотящие перейти отсюда к вам не могут, также и оттуда к нам не переходят.
LUKE|16|27|Тогда сказал он: так прошу тебя, отче, пошли его в дом отца моего,
LUKE|16|28|ибо у меня пять братьев; пусть он засвидетельствует им, чтобы и они не пришли в это место мучения.
LUKE|16|29|Авраам сказал ему: у них есть Моисей и пророки; пусть слушают их.
LUKE|16|30|Он же сказал: нет, отче Аврааме, но если кто из мертвых придет к ним, покаются.
LUKE|16|31|Тогда [Авраам] сказал ему: если Моисея и пророков не слушают, то если бы кто и из мертвых воскрес, не поверят.
LUKE|17|1|Сказал также [Иисус] ученикам: невозможно не придти соблазнам, но горе тому, через кого они приходят;
LUKE|17|2|лучше было бы ему, если бы мельничный жернов повесили ему на шею и бросили его в море, нежели чтобы он соблазнил одного из малых сих.
LUKE|17|3|Наблюдайте за собою. Если же согрешит против тебя брат твой, выговори ему; и если покается, прости ему;
LUKE|17|4|и если семь раз в день согрешит против тебя и семь раз в день обратится, и скажет: каюсь, – прости ему.
LUKE|17|5|И сказали Апостолы Господу: умножь в нас веру.
LUKE|17|6|Господь сказал: если бы вы имели веру с зерно горчичное и сказали смоковнице сей: исторгнись и пересадись в море, то она послушалась бы вас.
LUKE|17|7|Кто из вас, имея раба пашущего или пасущего, по возвращении его с поля, скажет ему: пойди скорее, садись за стол?
LUKE|17|8|Напротив, не скажет ли ему: приготовь мне поужинать и, подпоясавшись, служи мне, пока буду есть и пить, и потом ешь и пей сам?
LUKE|17|9|Станет ли он благодарить раба сего за то, что он исполнил приказание? Не думаю.
LUKE|17|10|Так и вы, когда исполните все повеленное вам, говорите: мы рабы ничего не стоящие, потому что сделали, что должны были сделать.
LUKE|17|11|Идя в Иерусалим, Он проходил между Самариею и Галилеею.
LUKE|17|12|И когда входил Он в одно селение, встретили Его десять человек прокаженных, которые остановились вдали
LUKE|17|13|и громким голосом говорили: Иисус Наставник! помилуй нас.
LUKE|17|14|Увидев [их], Он сказал им: пойдите, покажитесь священникам. И когда они шли, очистились.
LUKE|17|15|Один же из них, видя, что исцелен, возвратился, громким голосом прославляя Бога,
LUKE|17|16|и пал ниц к ногам Его, благодаря Его; и это был Самарянин.
LUKE|17|17|Тогда Иисус сказал: не десять ли очистились? где же девять?
LUKE|17|18|как они не возвратились воздать славу Богу, кроме сего иноплеменника?
LUKE|17|19|И сказал ему: встань, иди; вера твоя спасла тебя.
LUKE|17|20|Быв же спрошен фарисеями, когда придет Царствие Божие, отвечал им: не придет Царствие Божие приметным образом,
LUKE|17|21|и не скажут: вот, оно здесь, или: вот, там. Ибо вот, Царствие Божие внутрь вас есть.
LUKE|17|22|Сказал также ученикам: придут дни, когда пожелаете видеть хотя один из дней Сына Человеческого, и не увидите;
LUKE|17|23|и скажут вам: вот, здесь, или: вот, там, – не ходите и не гоняйтесь,
LUKE|17|24|ибо, как молния, сверкнувшая от одного края неба, блистает до другого края неба, так будет Сын Человеческий в день Свой.
LUKE|17|25|Но прежде надлежит Ему много пострадать и быть отвержену родом сим.
LUKE|17|26|И как было во дни Ноя, так будет и во дни Сына Человеческого:
LUKE|17|27|ели, пили, женились, выходили замуж, до того дня, как вошел Ной в ковчег, и пришел потоп и погубил всех.
LUKE|17|28|Так же, как было и во дни Лота: ели, пили, покупали, продавали, садили, строили;
LUKE|17|29|но в день, в который Лот вышел из Содома, пролился с неба дождь огненный и серный и истребил всех;
LUKE|17|30|так будет и в тот день, когда Сын Человеческий явится.
LUKE|17|31|В тот день, кто будет на кровле, а вещи его в доме, тот не сходи взять их; и кто будет на поле, также не обращайся назад.
LUKE|17|32|Вспоминайте жену Лотову.
LUKE|17|33|Кто станет сберегать душу свою, тот погубит ее; а кто погубит ее, тот оживит ее.
LUKE|17|34|Сказываю вам: в ту ночь будут двое на одной постели: один возьмется, а другой оставится;
LUKE|17|35|две будут молоть вместе: одна возьмется, а другая оставится;
LUKE|17|36|двое будут на поле: один возьмется, а другой оставится.
LUKE|17|37|На это сказали Ему: где, Господи? Он же сказал им: где труп, там соберутся и орлы.
LUKE|18|1|Сказал также им притчу о том, что должно всегда молиться и не унывать,
LUKE|18|2|говоря: в одном городе был судья, который Бога не боялся и людей не стыдился.
LUKE|18|3|В том же городе была одна вдова, и она, приходя к нему, говорила: защити меня от соперника моего.
LUKE|18|4|Но он долгое время не хотел. А после сказал сам в себе: хотя я и Бога не боюсь и людей не стыжусь,
LUKE|18|5|но, как эта вдова не дает мне покоя, защищу ее, чтобы она не приходила больше докучать мне.
LUKE|18|6|И сказал Господь: слышите, что говорит судья неправедный?
LUKE|18|7|Бог ли не защитит избранных Своих, вопиющих к Нему день и ночь, хотя и медлит защищать их?
LUKE|18|8|сказываю вам, что подаст им защиту вскоре. Но Сын Человеческий, придя, найдет ли веру на земле?
LUKE|18|9|Сказал также к некоторым, которые уверены были о себе, что они праведны, и уничижали других, следующую притчу:
LUKE|18|10|два человека вошли в храм помолиться: один фарисей, а другой мытарь.
LUKE|18|11|Фарисей, став, молился сам в себе так: Боже! благодарю Тебя, что я не таков, как прочие люди, грабители, обидчики, прелюбодеи, или как этот мытарь:
LUKE|18|12|пощусь два раза в неделю, даю десятую часть из всего, что приобретаю.
LUKE|18|13|Мытарь же, стоя вдали, не смел даже поднять глаз на небо; но, ударяя себя в грудь, говорил: Боже! будь милостив ко мне грешнику!
LUKE|18|14|Сказываю вам, что сей пошел оправданным в дом свой более, нежели тот: ибо всякий, возвышающий сам себя, унижен будет, а унижающий себя возвысится.
LUKE|18|15|Приносили к Нему и младенцев, чтобы Он прикоснулся к ним; ученики же, видя то, возбраняли им.
LUKE|18|16|Но Иисус, подозвав их, сказал: пустите детей приходить ко Мне и не возбраняйте им, ибо таковых есть Царствие Божие.
LUKE|18|17|Истинно говорю вам: кто не примет Царствия Божия, как дитя, тот не войдет в него.
LUKE|18|18|И спросил Его некто из начальствующих: Учитель благий! что мне делать, чтобы наследовать жизнь вечную?
LUKE|18|19|Иисус сказал ему: что ты называешь Меня благим? никто не благ, как только один Бог;
LUKE|18|20|знаешь заповеди: не прелюбодействуй, не убивай, не кради, не лжесвидетельствуй, почитай отца твоего и матерь твою.
LUKE|18|21|Он же сказал: все это сохранил я от юности моей.
LUKE|18|22|Услышав это, Иисус сказал ему: еще одного недостает тебе: все, что имеешь, продай и раздай нищим, и будешь иметь сокровище на небесах, и приходи, следуй за Мною.
LUKE|18|23|Он же, услышав сие, опечалился, потому что был очень богат.
LUKE|18|24|Иисус, видя, что он опечалился, сказал: как трудно имеющим богатство войти в Царствие Божие!
LUKE|18|25|ибо удобнее верблюду пройти сквозь игольные уши, нежели богатому войти в Царствие Божие.
LUKE|18|26|Слышавшие сие сказали: кто же может спастись?
LUKE|18|27|Но Он сказал: невозможное человекам возможно Богу.
LUKE|18|28|Петр же сказал: вот, мы оставили все и последовали за Тобою.
LUKE|18|29|Он сказал им: истинно говорю вам: нет никого, кто оставил бы дом, или родителей, или братьев, или сестер, или жену, или детей для Царствия Божия,
LUKE|18|30|и не получил бы гораздо более в сие время, и в век будущий жизни вечной.
LUKE|18|31|Отозвав же двенадцать учеников Своих, сказал им: вот, мы восходим в Иерусалим, и совершится все, написанное через пророков о Сыне Человеческом,
LUKE|18|32|ибо предадут Его язычникам, и поругаются над Ним, и оскорбят Его, и оплюют Его,
LUKE|18|33|и будут бить, и убьют Его: и в третий день воскреснет.
LUKE|18|34|Но они ничего из этого не поняли; слова сии были для них сокровенны, и они не разумели сказанного.
LUKE|18|35|Когда же подходил Он к Иерихону, один слепой сидел у дороги, прося милостыни,
LUKE|18|36|и, услышав, что мимо него проходит народ, спросил: что это такое?
LUKE|18|37|Ему сказали, что Иисус Назорей идет.
LUKE|18|38|Тогда он закричал: Иисус, Сын Давидов! помилуй меня.
LUKE|18|39|Шедшие впереди заставляли его молчать; но он еще громче кричал: Сын Давидов! помилуй меня.
LUKE|18|40|Иисус, остановившись, велел привести его к Себе: и, когда тот подошел к Нему, спросил его:
LUKE|18|41|чего ты хочешь от Меня? Он сказал: Господи! чтобы мне прозреть.
LUKE|18|42|Иисус сказал ему: прозри! вера твоя спасла тебя.
LUKE|18|43|И он тотчас прозрел и пошел за Ним, славя Бога; и весь народ, видя это, воздал хвалу Богу.
LUKE|19|1|Потом [Иисус] вошел в Иерихон и проходил через него.
LUKE|19|2|И вот, некто, именем Закхей, начальник мытарей и человек богатый,
LUKE|19|3|искал видеть Иисуса, кто Он, но не мог за народом, потому что мал был ростом,
LUKE|19|4|и, забежав вперед, взлез на смоковницу, чтобы увидеть Его, потому что Ему надлежало проходить мимо нее.
LUKE|19|5|Иисус, когда пришел на это место, взглянув, увидел его и сказал ему: Закхей! сойди скорее, ибо сегодня надобно Мне быть у тебя в доме.
LUKE|19|6|И он поспешно сошел и принял Его с радостью.
LUKE|19|7|И все, видя то, начали роптать, и говорили, что Он зашел к грешному человеку;
LUKE|19|8|Закхей же, став, сказал Господу: Господи! половину имения моего я отдам нищим, и, если кого чем обидел, воздам вчетверо.
LUKE|19|9|Иисус сказал ему: ныне пришло спасение дому сему, потому что и он сын Авраама,
LUKE|19|10|ибо Сын Человеческий пришел взыскать и спасти погибшее.
LUKE|19|11|Когда же они слушали это, присовокупил притчу: ибо Он был близ Иерусалима, и они думали, что скоро должно открыться Царствие Божие.
LUKE|19|12|Итак сказал: некоторый человек высокого рода отправлялся в дальнюю страну, чтобы получить себе царство и возвратиться;
LUKE|19|13|призвав же десять рабов своих, дал им десять мин и сказал им: употребляйте их в оборот, пока я возвращусь.
LUKE|19|14|Но граждане ненавидели его и отправили вслед за ним посольство, сказав: не хотим, чтобы он царствовал над нами.
LUKE|19|15|И когда возвратился, получив царство, велел призвать к себе рабов тех, которым дал серебро, чтобы узнать, кто что приобрел.
LUKE|19|16|Пришел первый и сказал: господин! мина твоя принесла десять мин.
LUKE|19|17|И сказал ему: хорошо, добрый раб! за то, что ты в малом был верен, возьми в управление десять городов.
LUKE|19|18|Пришел второй и сказал: господин! мина твоя принесла пять мин.
LUKE|19|19|Сказал и этому: и ты будь над пятью городами.
LUKE|19|20|Пришел третий и сказал: господин! вот твоя мина, которую я хранил, завернув в платок,
LUKE|19|21|ибо я боялся тебя, потому что ты человек жестокий: берешь, чего не клал, и жнешь, чего не сеял.
LUKE|19|22|[Господин] сказал ему: твоими устами буду судить тебя, лукавый раб! ты знал, что я человек жестокий, беру, чего не клал, и жну, чего не сеял;
LUKE|19|23|для чего же ты не отдал серебра моего в оборот, чтобы я, придя, получил его с прибылью?
LUKE|19|24|И сказал предстоящим: возьмите у него мину и дайте имеющему десять мин.
LUKE|19|25|И сказали ему: господин! у него есть десять мин.
LUKE|19|26|Сказываю вам, что всякому имеющему дано будет, а у неимеющего отнимется и то, что имеет;
LUKE|19|27|врагов же моих тех, которые не хотели, чтобы я царствовал над ними, приведите сюда и избейте предо мною.
LUKE|19|28|Сказав это, Он пошел далее, восходя в Иерусалим.
LUKE|19|29|И когда приблизился к Виффагии и Вифании, к горе, называемой Елеонскою, послал двух учеников Своих,
LUKE|19|30|сказав: пойдите в противолежащее селение; войдя в него, найдете молодого осла привязанного, на которого никто из людей никогда не садился; отвязав его, приведите;
LUKE|19|31|и если кто спросит вас: зачем отвязываете? скажите ему так: он надобен Господу.
LUKE|19|32|Посланные пошли и нашли, как Он сказал им.
LUKE|19|33|Когда же они отвязывали молодого осла, хозяева его сказали им: зачем отвязываете осленка?
LUKE|19|34|Они отвечали: он надобен Господу.
LUKE|19|35|И привели его к Иисусу, и, накинув одежды свои на осленка, посадили на него Иисуса.
LUKE|19|36|И, когда Он ехал, постилали одежды свои по дороге.
LUKE|19|37|А когда Он приблизился к спуску с горы Елеонской, все множество учеников начало в радости велегласно славить Бога за все чудеса, какие видели они,
LUKE|19|38|говоря: благословен Царь, грядущий во имя Господне! мир на небесах и слава в вышних!
LUKE|19|39|И некоторые фарисеи из среды народа сказали Ему: Учитель! запрети ученикам Твоим.
LUKE|19|40|Но Он сказал им в ответ: сказываю вам, что если они умолкнут, то камни возопиют.
LUKE|19|41|И когда приблизился к городу, то, смотря на него, заплакал о нем
LUKE|19|42|и сказал: о, если бы и ты хотя в сей твой день узнал, что служит к миру твоему! Но это сокрыто ныне от глаз твоих,
LUKE|19|43|ибо придут на тебя дни, когда враги твои обложат тебя окопами и окружат тебя, и стеснят тебя отовсюду,
LUKE|19|44|и разорят тебя, и побьют детей твоих в тебе, и не оставят в тебе камня на камне за то, что ты не узнал времени посещения твоего.
LUKE|19|45|И, войдя в храм, начал выгонять продающих в нем и покупающих,
LUKE|19|46|говоря им: написано: дом Мой есть дом молитвы, а вы сделали его вертепом разбойников.
LUKE|19|47|И учил каждый день в храме. Первосвященники же и книжники и старейшины народа искали погубить Его,
LUKE|19|48|и не находили, что бы сделать с Ним; потому что весь народ неотступно слушал Его.
LUKE|20|1|В один из тех дней, когда Он учил народ в храме и благовествовал, приступили первосвященники и книжники со старейшинами,
LUKE|20|2|и сказали Ему: скажи нам, какою властью Ты это делаешь, или кто дал Тебе власть сию?
LUKE|20|3|Он сказал им в ответ: спрошу и Я вас об одном, и скажите Мне:
LUKE|20|4|крещение Иоанново с небес было, или от человеков?
LUKE|20|5|Они же, рассуждая между собою, говорили: если скажем: с небес, то скажет: почему же вы не поверили ему?
LUKE|20|6|а если скажем: от человеков, то весь народ побьет нас камнями, ибо он уверен, что Иоанн есть пророк.
LUKE|20|7|И отвечали: не знаем откуда.
LUKE|20|8|Иисус сказал им: и Я не скажу вам, какою властью это делаю.
LUKE|20|9|И начал Он говорить к народу притчу сию: один человек насадил виноградник и отдал его виноградарям, и отлучился на долгое время;
LUKE|20|10|и в свое время послал к виноградарям раба, чтобы они дали ему плодов из виноградника; но виноградари, прибив его, отослали ни с чем.
LUKE|20|11|Еще послал другого раба; но они и этого, прибив и обругав, отослали ни с чем.
LUKE|20|12|И еще послал третьего; но они и того, изранив, выгнали.
LUKE|20|13|Тогда сказал господин виноградника: что мне делать? Пошлю сына моего возлюбленного; может быть, увидев его, постыдятся.
LUKE|20|14|Но виноградари, увидев его, рассуждали между собою, говоря: это наследник; пойдем, убьем его, и наследство его будет наше.
LUKE|20|15|И, выведя его вон из виноградника, убили. Что же сделает с ними господин виноградника?
LUKE|20|16|Придет и погубит виноградарей тех, и отдаст виноградник другим. Слышавшие же это сказали: да не будет!
LUKE|20|17|Но Он, взглянув на них, сказал: что значит сие написанное: камень, который отвергли строители, тот самый сделался главою угла?
LUKE|20|18|Всякий, кто упадет на тот камень, разобьется, а на кого он упадет, того раздавит.
LUKE|20|19|И искали в это время первосвященники и книжники, чтобы наложить на Него руки, но побоялись народа, ибо поняли, что о них сказал Он эту притчу.
LUKE|20|20|И, наблюдая за Ним, подослали лукавых людей, которые, притворившись благочестивыми, уловили бы Его в каком–либо слове, чтобы предать Его начальству и власти правителя.
LUKE|20|21|И они спросили Его: Учитель! мы знаем, что Ты правдиво говоришь и учишь и не смотришь на лице, но истинно пути Божию учишь;
LUKE|20|22|позволительно ли нам давать подать кесарю, или нет?
LUKE|20|23|Он же, уразумев лукавство их, сказал им: что вы Меня искушаете?
LUKE|20|24|Покажите Мне динарий: чье на нем изображение и надпись? Они отвечали: кесаревы.
LUKE|20|25|Он сказал им: итак, отдавайте кесарево кесарю, а Божие Богу.
LUKE|20|26|И не могли уловить Его в слове перед народом, и, удивившись ответу Его, замолчали.
LUKE|20|27|Тогда пришли некоторые из саддукеев, отвергающих воскресение, и спросили Его:
LUKE|20|28|Учитель! Моисей написал нам, что если у кого умрет брат, имевший жену, и умрет бездетным, то брат его должен взять его жену и восставить семя брату своему.
LUKE|20|29|Было семь братьев, первый, взяв жену, умер бездетным;
LUKE|20|30|взял ту жену второй, и тот умер бездетным;
LUKE|20|31|взял ее третий; также и все семеро, и умерли, не оставив детей;
LUKE|20|32|после всех умерла и жена;
LUKE|20|33|итак, в воскресение которого из них будет она женою, ибо семеро имели ее женою?
LUKE|20|34|Иисус сказал им в ответ: чада века сего женятся и выходят замуж;
LUKE|20|35|а сподобившиеся достигнуть того века и воскресения из мертвых ни женятся, ни замуж не выходят,
LUKE|20|36|и умереть уже не могут, ибо они равны Ангелам и суть сыны Божии, будучи сынами воскресения.
LUKE|20|37|А что мертвые воскреснут, и Моисей показал при купине, когда назвал Господа Богом Авраама и Богом Исаака и Богом Иакова.
LUKE|20|38|Бог же не есть [Бог] мертвых, но живых, ибо у Него все живы.
LUKE|20|39|На это некоторые из книжников сказали: Учитель! Ты хорошо сказал.
LUKE|20|40|И уже не смели спрашивать Его ни о чем. Он же сказал им:
LUKE|20|41|как говорят, что Христос есть Сын Давидов,
LUKE|20|42|а сам Давид говорит в книге псалмов: сказал Господь Господу моему: седи одесную Меня,
LUKE|20|43|доколе положу врагов Твоих в подножие ног Твоих?
LUKE|20|44|Итак, Давид Господом называет Его; как же Он Сын ему?
LUKE|20|45|И когда слушал весь народ, Он сказал ученикам Своим:
LUKE|20|46|остерегайтесь книжников, которые любят ходить в длинных одеждах и любят приветствия в народных собраниях, председания в синагогах и предвозлежания на пиршествах,
LUKE|20|47|которые поедают домы вдов и лицемерно долго молятся; они примут тем большее осуждение.
LUKE|21|1|Взглянув же, Он увидел богатых, клавших дары свои в сокровищницу;
LUKE|21|2|увидел также и бедную вдову, положившую туда две лепты,
LUKE|21|3|и сказал: истинно говорю вам, что эта бедная вдова больше всех положила;
LUKE|21|4|ибо все те от избытка своего положили в дар Богу, а она от скудости своей положила все пропитание свое, какое имела.
LUKE|21|5|И когда некоторые говорили о храме, что он украшен дорогими камнями и вкладами, Он сказал:
LUKE|21|6|придут дни, в которые из того, что вы здесь видите, не останется камня на камне; все будет разрушено.
LUKE|21|7|И спросили Его: Учитель! когда же это будет? и какой признак, когда это должно произойти?
LUKE|21|8|Он сказал: берегитесь, чтобы вас не ввели в заблуждение, ибо многие придут под именем Моим, говоря, что это Я; и это время близко: не ходите вслед их.
LUKE|21|9|Когда же услышите о войнах и смятениях, не ужасайтесь, ибо этому надлежит быть прежде; но не тотчас конец.
LUKE|21|10|Тогда сказал им: восстанет народ на народ, и царство на царство;
LUKE|21|11|будут большие землетрясения по местам, и глады, и моры, и ужасные явления, и великие знамения с неба.
LUKE|21|12|Прежде же всего того возложат на вас руки и будут гнать [вас], предавая в синагоги и в темницы, и поведут пред царей и правителей за имя Мое;
LUKE|21|13|будет же это вам для свидетельства.
LUKE|21|14|Итак положите себе на сердце не обдумывать заранее, что отвечать,
LUKE|21|15|ибо Я дам вам уста и премудрость, которой не возмогут противоречить ни противостоять все, противящиеся вам.
LUKE|21|16|Преданы также будете и родителями, и братьями, и родственниками, и друзьями, и некоторых из вас умертвят;
LUKE|21|17|и будете ненавидимы всеми за имя Мое,
LUKE|21|18|но и волос с головы вашей не пропадет, –
LUKE|21|19|терпением вашим спасайте души ваши.
LUKE|21|20|Когда же увидите Иерусалим, окруженный войсками, тогда знайте, что приблизилось запустение его:
LUKE|21|21|тогда находящиеся в Иудее да бегут в горы; и кто в городе, выходи из него; и кто в окрестностях, не входи в него,
LUKE|21|22|потому что это дни отмщения, да исполнится все написанное.
LUKE|21|23|Горе же беременным и питающим сосцами в те дни; ибо великое будет бедствие на земле и гнев на народ сей:
LUKE|21|24|и падут от острия меча, и отведутся в плен во все народы; и Иерусалим будет попираем язычниками, доколе не окончатся времена язычников.
LUKE|21|25|И будут знамения в солнце и луне и звездах, а на земле уныние народов и недоумение; и море восшумит и возмутится;
LUKE|21|26|люди будут издыхать от страха и ожидания [бедствий], грядущих на вселенную, ибо силы небесные поколеблются,
LUKE|21|27|и тогда увидят Сына Человеческого, грядущего на облаке с силою и славою великою.
LUKE|21|28|Когда же начнет это сбываться, тогда восклонитесь и поднимите головы ваши, потому что приближается избавление ваше.
LUKE|21|29|И сказал им притчу: посмотрите на смоковницу и на все деревья:
LUKE|21|30|когда они уже распускаются, то, видя это, знаете сами, что уже близко лето.
LUKE|21|31|Так, и когда вы увидите то сбывающимся, знайте, что близко Царствие Божие.
LUKE|21|32|Истинно говорю вам: не прейдет род сей, как все это будет;
LUKE|21|33|небо и земля прейдут, но слова Мои не прейдут.
LUKE|21|34|Смотрите же за собою, чтобы сердца ваши не отягчались объядением и пьянством и заботами житейскими, и чтобы день тот не постиг вас внезапно,
LUKE|21|35|ибо он, как сеть, найдет на всех живущих по всему лицу земному;
LUKE|21|36|итак бодрствуйте на всякое время и молитесь, да сподобитесь избежать всех сих будущих [бедствий] и предстать пред Сына Человеческого.
LUKE|21|37|Днем Он учил в храме, а ночи, выходя, проводил на горе, называемой Елеонскою.
LUKE|21|38|И весь народ с утра приходил к Нему в храм слушать Его.
LUKE|22|1|Приближался праздник опресноков, называемый Пасхою,
LUKE|22|2|и искали первосвященники и книжники, как бы погубить Его, потому что боялись народа.
LUKE|22|3|Вошел же сатана в Иуду, прозванного Искариотом, одного из числа двенадцати,
LUKE|22|4|и он пошел, и говорил с первосвященниками и начальниками, как Его предать им.
LUKE|22|5|Они обрадовались и согласились дать ему денег;
LUKE|22|6|и он обещал, и искал удобного времени, чтобы предать Его им не при народе.
LUKE|22|7|Настал же день опресноков, в который надлежало заколать пасхального [агнца],
LUKE|22|8|и послал [Иисус] Петра и Иоанна, сказав: пойдите, приготовьте нам есть пасху.
LUKE|22|9|Они же сказали Ему: где велишь нам приготовить?
LUKE|22|10|Он сказал им: вот, при входе вашем в город, встретится с вами человек, несущий кувшин воды; последуйте за ним в дом, в который войдет он,
LUKE|22|11|и скажите хозяину дома: Учитель говорит тебе: где комната, в которой бы Мне есть пасху с учениками Моими?
LUKE|22|12|И он покажет вам горницу большую устланную; там приготовьте.
LUKE|22|13|Они пошли, и нашли, как сказал им, и приготовили пасху.
LUKE|22|14|И когда настал час, Он возлег, и двенадцать Апостолов с Ним,
LUKE|22|15|и сказал им: очень желал Я есть с вами сию пасху прежде Моего страдания,
LUKE|22|16|ибо сказываю вам, что уже не буду есть ее, пока она не совершится в Царствии Божием.
LUKE|22|17|И, взяв чашу и благодарив, сказал: приимите ее и разделите между собою,
LUKE|22|18|ибо сказываю вам, что не буду пить от плода виноградного, доколе не придет Царствие Божие.
LUKE|22|19|И, взяв хлеб и благодарив, преломил и подал им, говоря: сие есть тело Мое, которое за вас предается; сие творите в Мое воспоминание.
LUKE|22|20|Также и чашу после вечери, говоря: сия чаша [есть] Новый Завет в Моей крови, которая за вас проливается.
LUKE|22|21|И вот, рука предающего Меня со Мною за столом;
LUKE|22|22|впрочем, Сын Человеческий идет по предназначению, но горе тому человеку, которым Он предается.
LUKE|22|23|И они начали спрашивать друг друга, кто бы из них был, который это сделает.
LUKE|22|24|Был же и спор между ними, кто из них должен почитаться большим.
LUKE|22|25|Он же сказал им: цари господствуют над народами, и владеющие ими благодетелями называются,
LUKE|22|26|а вы не так: но кто из вас больше, будь как меньший, и начальствующий – как служащий.
LUKE|22|27|Ибо кто больше: возлежащий, или служащий? не возлежащий ли? А Я посреди вас, как служащий.
LUKE|22|28|Но вы пребыли со Мною в напастях Моих,
LUKE|22|29|и Я завещаваю вам, как завещал Мне Отец Мой, Царство,
LUKE|22|30|да ядите и пиете за трапезою Моею в Царстве Моем, и сядете на престолах судить двенадцать колен Израилевых.
LUKE|22|31|И сказал Господь: Симон! Симон! се, сатана просил, чтобы сеять вас как пшеницу,
LUKE|22|32|но Я молился о тебе, чтобы не оскудела вера твоя; и ты некогда, обратившись, утверди братьев твоих.
LUKE|22|33|Он отвечал Ему: Господи! с Тобою я готов и в темницу и на смерть идти.
LUKE|22|34|Но Он сказал: говорю тебе, Петр, не пропоет петух сегодня, как ты трижды отречешься, что не знаешь Меня.
LUKE|22|35|И сказал им: когда Я посылал вас без мешка и без сумы и без обуви, имели ли вы в чем недостаток? Они отвечали: ни в чем.
LUKE|22|36|Тогда Он сказал им: но теперь, кто имеет мешок, тот возьми его, также и суму; а у кого нет, продай одежду свою и купи меч;
LUKE|22|37|ибо сказываю вам, что должно исполниться на Мне и сему написанному: и к злодеям причтен. Ибо то, что о Мне, приходит к концу.
LUKE|22|38|Они сказали: Господи! вот, здесь два меча. Он сказал им: довольно.
LUKE|22|39|И, выйдя, пошел по обыкновению на гору Елеонскую, за Ним последовали и ученики Его.
LUKE|22|40|Придя же на место, сказал им: молитесь, чтобы не впасть в искушение.
LUKE|22|41|И Сам отошел от них на вержение камня, и, преклонив колени, молился,
LUKE|22|42|говоря: Отче! о, если бы Ты благоволил пронести чашу сию мимо Меня! впрочем не Моя воля, но Твоя да будет.
LUKE|22|43|Явился же Ему Ангел с небес и укреплял Его.
LUKE|22|44|И, находясь в борении, прилежнее молился, и был пот Его, как капли крови, падающие на землю.
LUKE|22|45|Встав от молитвы, Он пришел к ученикам, и нашел их спящими от печали
LUKE|22|46|и сказал им: что вы спите? встаньте и молитесь, чтобы не впасть в искушение.
LUKE|22|47|Когда Он еще говорил это, появился народ, а впереди его шел один из двенадцати, называемый Иуда, и он подошел к Иисусу, чтобы поцеловать Его. Ибо он такой им дал знак: Кого я поцелую, Тот и есть.
LUKE|22|48|Иисус же сказал ему: Иуда! целованием ли предаешь Сына Человеческого?
LUKE|22|49|Бывшие же с Ним, видя, к чему идет дело, сказали Ему: Господи! не ударить ли нам мечом?
LUKE|22|50|И один из них ударил раба первосвященникова, и отсек ему правое ухо.
LUKE|22|51|Тогда Иисус сказал: оставьте, довольно. И, коснувшись уха его, исцелил его.
LUKE|22|52|Первосвященникам же и начальникам храма и старейшинам, собравшимся против Него, сказал Иисус: как будто на разбойника вышли вы с мечами и кольями, чтобы взять Меня?
LUKE|22|53|Каждый день бывал Я с вами в храме, и вы не поднимали на Меня рук, но теперь ваше время и власть тьмы.
LUKE|22|54|Взяв Его, повели и привели в дом первосвященника. Петр же следовал издали.
LUKE|22|55|Когда они развели огонь среди двора и сели вместе, сел и Петр между ними.
LUKE|22|56|Одна служанка, увидев его сидящего у огня и всмотревшись в него, сказала: и этот был с Ним.
LUKE|22|57|Но он отрекся от Него, сказав женщине: я не знаю Его.
LUKE|22|58|Вскоре потом другой, увидев его, сказал: и ты из них. Но Петр сказал этому человеку: нет!
LUKE|22|59|Прошло с час времени, еще некто настоятельно говорил: точно и этот был с Ним, ибо он Галилеянин.
LUKE|22|60|Но Петр сказал тому человеку: не знаю, что ты говоришь. И тотчас, когда еще говорил он, запел петух.
LUKE|22|61|Тогда Господь, обратившись, взглянул на Петра, и Петр вспомнил слово Господа, как Он сказал ему: прежде нежели пропоет петух, отречешься от Меня трижды.
LUKE|22|62|И, выйдя вон, горько заплакал.
LUKE|22|63|Люди, державшие Иисуса, ругались над Ним и били Его;
LUKE|22|64|и, закрыв Его, ударяли Его по лицу и спрашивали Его: прореки, кто ударил Тебя?
LUKE|22|65|И много иных хулений произносили против Него.
LUKE|22|66|И как настал день, собрались старейшины народа, первосвященники и книжники, и ввели Его в свой синедрион
LUKE|22|67|и сказали: Ты ли Христос? скажи нам. Он сказал им: если скажу вам, вы не поверите;
LUKE|22|68|если же и спрошу вас, не будете отвечать Мне и не отпустите [Меня];
LUKE|22|69|отныне Сын Человеческий воссядет одесную силы Божией.
LUKE|22|70|И сказали все: итак, Ты Сын Божий? Он отвечал им: вы говорите, что Я.
LUKE|22|71|Они же сказали: какое еще нужно нам свидетельство? ибо мы сами слышали из уст Его.
LUKE|23|1|И поднялось все множество их, и повели Его к Пилату,
LUKE|23|2|и начали обвинять Его, говоря: мы нашли, что Он развращает народ наш и запрещает давать подать кесарю, называя Себя Христом Царем.
LUKE|23|3|Пилат спросил Его: Ты Царь Иудейский? Он сказал ему в ответ: ты говоришь.
LUKE|23|4|Пилат сказал первосвященникам и народу: я не нахожу никакой вины в этом человеке.
LUKE|23|5|Но они настаивали, говоря, что Он возмущает народ, уча по всей Иудее, начиная от Галилеи до сего места.
LUKE|23|6|Пилат, услышав о Галилее, спросил: разве Он Галилеянин?
LUKE|23|7|И, узнав, что Он из области Иродовой, послал Его к Ироду, который в эти дни был также в Иерусалиме.
LUKE|23|8|Ирод, увидев Иисуса, очень обрадовался, ибо давно желал видеть Его, потому что много слышал о Нем, и надеялся увидеть от Него какое–нибудь чудо,
LUKE|23|9|и предлагал Ему многие вопросы, но Он ничего не отвечал ему.
LUKE|23|10|Первосвященники же и книжники стояли и усильно обвиняли Его.
LUKE|23|11|Но Ирод со своими воинами, уничижив Его и насмеявшись над Ним, одел Его в светлую одежду и отослал обратно к Пилату.
LUKE|23|12|И сделались в тот день Пилат и Ирод друзьями между собою, ибо прежде были во вражде друг с другом.
LUKE|23|13|Пилат же, созвав первосвященников и начальников и народ,
LUKE|23|14|сказал им: вы привели ко мне человека сего, как развращающего народ; и вот, я при вас исследовал и не нашел человека сего виновным ни в чем том, в чем вы обвиняете Его;
LUKE|23|15|и Ирод также, ибо я посылал Его к нему; и ничего не найдено в Нем достойного смерти;
LUKE|23|16|итак, наказав Его, отпущу.
LUKE|23|17|А ему и нужно было для праздника отпустить им одного [узника].
LUKE|23|18|Но весь народ стал кричать: смерть Ему! а отпусти нам Варавву.
LUKE|23|19|Варавва был посажен в темницу за произведенное в городе возмущение и убийство.
LUKE|23|20|Пилат снова возвысил голос, желая отпустить Иисуса.
LUKE|23|21|Но они кричали: распни, распни Его!
LUKE|23|22|Он в третий раз сказал им: какое же зло сделал Он? я ничего достойного смерти не нашел в Нем; итак, наказав Его, отпущу.
LUKE|23|23|Но они продолжали с великим криком требовать, чтобы Он был распят; и превозмог крик их и первосвященников.
LUKE|23|24|И Пилат решил быть по прошению их,
LUKE|23|25|и отпустил им посаженного за возмущение и убийство в темницу, которого они просили; а Иисуса предал в их волю.
LUKE|23|26|И когда повели Его, то, захватив некоего Симона Киринеянина, шедшего с поля, возложили на него крест, чтобы нес за Иисусом.
LUKE|23|27|И шло за Ним великое множество народа и женщин, которые плакали и рыдали о Нем.
LUKE|23|28|Иисус же, обратившись к ним, сказал: дщери Иерусалимские! не плачьте обо Мне, но плачьте о себе и о детях ваших,
LUKE|23|29|ибо приходят дни, в которые скажут: блаженны неплодные, и утробы неродившие, и сосцы непитавшие!
LUKE|23|30|тогда начнут говорить горам: падите на нас! и холмам: покройте нас!
LUKE|23|31|Ибо если с зеленеющим деревом это делают, то с сухим что будет?
LUKE|23|32|Вели с Ним на смерть и двух злодеев.
LUKE|23|33|И когда пришли на место, называемое Лобное, там распяли Его и злодеев, одного по правую, а другого по левую сторону.
LUKE|23|34|Иисус же говорил: Отче! прости им, ибо не знают, что делают. И делили одежды Его, бросая жребий.
LUKE|23|35|И стоял народ и смотрел. Насмехались же вместе с ними и начальники, говоря: других спасал; пусть спасет Себя Самого, если Он Христос, избранный Божий.
LUKE|23|36|Также и воины ругались над Ним, подходя и поднося Ему уксус
LUKE|23|37|и говоря: если Ты Царь Иудейский, спаси Себя Самого.
LUKE|23|38|И была над Ним надпись, написанная словами греческими, римскими и еврейскими: Сей есть Царь Иудейский.
LUKE|23|39|Один из повешенных злодеев злословил Его и говорил: если Ты Христос, спаси Себя и нас.
LUKE|23|40|Другой же, напротив, унимал его и говорил: или ты не боишься Бога, когда и сам осужден на то же?
LUKE|23|41|и мы [осуждены] справедливо, потому что достойное по делам нашим приняли, а Он ничего худого не сделал.
LUKE|23|42|И сказал Иисусу: помяни меня, Господи, когда приидешь в Царствие Твое!
LUKE|23|43|И сказал ему Иисус: истинно говорю тебе, ныне же будешь со Мною в раю.
LUKE|23|44|Было же около шестого часа дня, и сделалась тьма по всей земле до часа девятого:
LUKE|23|45|и померкло солнце, и завеса в храме раздралась по средине.
LUKE|23|46|Иисус, возгласив громким голосом, сказал: Отче! в руки Твои предаю дух Мой. И, сие сказав, испустил дух.
LUKE|23|47|Сотник же, видев происходившее, прославил Бога и сказал: истинно человек этот был праведник.
LUKE|23|48|И весь народ, сшедшийся на сие зрелище, видя происходившее, возвращался, бия себя в грудь.
LUKE|23|49|Все же, знавшие Его, и женщины, следовавшие за Ним из Галилеи, стояли вдали и смотрели на это.
LUKE|23|50|Тогда некто, именем Иосиф, член совета, человек добрый и правдивый,
LUKE|23|51|не участвовавший в совете и в деле их; из Аримафеи, города Иудейского, ожидавший также Царствия Божия,
LUKE|23|52|пришел к Пилату и просил тела Иисусова;
LUKE|23|53|и, сняв его, обвил плащаницею и положил его в гробе, высеченном [в скале], где еще никто не был положен.
LUKE|23|54|День тот был пятница, и наступала суббота.
LUKE|23|55|Последовали также и женщины, пришедшие с Иисусом из Галилеи, и смотрели гроб, и как полагалось тело Его;
LUKE|23|56|возвратившись же, приготовили благовония и масти; и в субботу остались в покое по заповеди.
LUKE|24|1|В первый же день недели, очень рано, неся приготовленные ароматы, пришли они ко гробу, и вместе с ними некоторые другие;
LUKE|24|2|но нашли камень отваленным от гроба.
LUKE|24|3|И, войдя, не нашли тела Господа Иисуса.
LUKE|24|4|Когда же недоумевали они о сем, вдруг предстали перед ними два мужа в одеждах блистающих.
LUKE|24|5|И когда они были в страхе и наклонили лица [свои] к земле, сказали им: что вы ищете живого между мертвыми?
LUKE|24|6|Его нет здесь: Он воскрес; вспомните, как Он говорил вам, когда был еще в Галилее,
LUKE|24|7|сказывая, что Сыну Человеческому надлежит быть предану в руки человеков грешников, и быть распяту, и в третий день воскреснуть.
LUKE|24|8|И вспомнили они слова Его;
LUKE|24|9|и, возвратившись от гроба, возвестили все это одиннадцати и всем прочим.
LUKE|24|10|То были Магдалина Мария, и Иоанна, и Мария, [мать] Иакова, и другие с ними, которые сказали о сем Апостолам.
LUKE|24|11|И показались им слова их пустыми, и не поверили им.
LUKE|24|12|Но Петр, встав, побежал ко гробу и, наклонившись, увидел только пелены лежащие, и пошел назад, дивясь сам в себе происшедшему.
LUKE|24|13|В тот же день двое из них шли в селение, отстоящее стадий на шестьдесят от Иерусалима, называемое Эммаус;
LUKE|24|14|и разговаривали между собою о всех сих событиях.
LUKE|24|15|И когда они разговаривали и рассуждали между собою, и Сам Иисус, приблизившись, пошел с ними.
LUKE|24|16|Но глаза их были удержаны, так что они не узнали Его.
LUKE|24|17|Он же сказал им: о чем это вы, идя, рассуждаете между собою, и отчего вы печальны?
LUKE|24|18|Один из них, именем Клеопа, сказал Ему в ответ: неужели Ты один из пришедших в Иерусалим не знаешь о происшедшем в нем в эти дни?
LUKE|24|19|И сказал им: о чем? Они сказали Ему: что было с Иисусом Назарянином, Который был пророк, сильный в деле и слове пред Богом и всем народом;
LUKE|24|20|как предали Его первосвященники и начальники наши для осуждения на смерть и распяли Его.
LUKE|24|21|А мы надеялись было, что Он есть Тот, Который должен избавить Израиля; но со всем тем, уже третий день ныне, как это произошло.
LUKE|24|22|Но и некоторые женщины из наших изумили нас: они были рано у гроба
LUKE|24|23|и не нашли тела Его и, придя, сказывали, что они видели и явление Ангелов, которые говорят, что Он жив.
LUKE|24|24|И пошли некоторые из наших ко гробу и нашли так, как и женщины говорили, но Его не видели.
LUKE|24|25|Тогда Он сказал им: о, несмысленные и медлительные сердцем, чтобы веровать всему, что предсказывали пророки!
LUKE|24|26|Не так ли надлежало пострадать Христу и войти в славу Свою?
LUKE|24|27|И, начав от Моисея, из всех пророков изъяснял им сказанное о Нем во всем Писании.
LUKE|24|28|И приблизились они к тому селению, в которое шли; и Он показывал им вид, что хочет идти далее.
LUKE|24|29|Но они удерживали Его, говоря: останься с нами, потому что день уже склонился к вечеру. И Он вошел и остался с ними.
LUKE|24|30|И когда Он возлежал с ними, то, взяв хлеб, благословил, преломил и подал им.
LUKE|24|31|Тогда открылись у них глаза, и они узнали Его. Но Он стал невидим для них.
LUKE|24|32|И они сказали друг другу: не горело ли в нас сердце наше, когда Он говорил нам на дороге и когда изъяснял нам Писание?
LUKE|24|33|И, встав в тот же час, возвратились в Иерусалим и нашли вместе одиннадцать [Апостолов] и бывших с ними,
LUKE|24|34|которые говорили, что Господь истинно воскрес и явился Симону.
LUKE|24|35|И они рассказывали о происшедшем на пути, и как Он был узнан ими в преломлении хлеба.
LUKE|24|36|Когда они говорили о сем, Сам Иисус стал посреди них и сказал им: мир вам.
LUKE|24|37|Они, смутившись и испугавшись, подумали, что видят духа.
LUKE|24|38|Но Он сказал им: что смущаетесь, и для чего такие мысли входят в сердца ваши?
LUKE|24|39|Посмотрите на руки Мои и на ноги Мои; это Я Сам; осяжите Меня и рассмотрите; ибо дух плоти и костей не имеет, как видите у Меня.
LUKE|24|40|И, сказав это, показал им руки и ноги.
LUKE|24|41|Когда же они от радости еще не верили и дивились, Он сказал им: есть ли у вас здесь какая пища?
LUKE|24|42|Они подали Ему часть печеной рыбы и сотового меда.
LUKE|24|43|И, взяв, ел пред ними.
LUKE|24|44|И сказал им: вот то, о чем Я вам говорил, еще быв с вами, что надлежит исполниться всему, написанному о Мне в законе Моисеевом и в пророках и псалмах.
LUKE|24|45|Тогда отверз им ум к уразумению Писаний.
LUKE|24|46|И сказал им: так написано, и так надлежало пострадать Христу, и воскреснуть из мертвых в третий день,
LUKE|24|47|и проповедану быть во имя Его покаянию и прощению грехов во всех народах, начиная с Иерусалима.
LUKE|24|48|Вы же свидетели сему.
LUKE|24|49|И Я пошлю обетование Отца Моего на вас; вы же оставайтесь в городе Иерусалиме, доколе не облечетесь силою свыше.
LUKE|24|50|И вывел их вон [из города] до Вифании и, подняв руки Свои, благословил их.
LUKE|24|51|И, когда благословлял их, стал отдаляться от них и возноситься на небо.
LUKE|24|52|Они поклонились Ему и возвратились в Иерусалим с великою радостью.
LUKE|24|53|И пребывали всегда в храме, прославляя и благословляя Бога. Аминь.
