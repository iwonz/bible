JOEL|1|1|Слово Господнє, що було до Йоіла, Петуїлового сина.
JOEL|1|2|Послухайте це, ви старші, і візьміть до вух, усі мешканці землі: чи бувало таке за днів ваших, або за днів ваших батьків?
JOEL|1|3|Оповідайте про це синам вашим, а ваші сини своїм дітям, а їхні сини поколінню наступному.
JOEL|1|4|Що лишилось по гусені, зжерла те все сарана, що ж зосталося по сарані пожер коник, а решту по конику зжерла черва.
JOEL|1|5|Пробудіться, п'яниці, і плачте й ридайте за виноградовим соком усі, хто вина напивається, бо віднятий він від уст ваших!
JOEL|1|6|Бо на Край Мій прийшов люд міцний й незчисленний, його зуби як лев'ячі зуби, а паща його як в левиці.
JOEL|1|7|Виноград Мій зробив він спустошенням, Моє ж фіґове дерево геть поламав, дощенту його оголив та й покинув, галузки його побіліли.
JOEL|1|8|Голоси, як та дівчина, веретою оперезана, за нареченим юнацтва свого.
JOEL|1|9|Жертва хлібна й жертва лита спинилася в домі Господньому, впали в жалобу священики, слуги Господні.
JOEL|1|10|Опустошене поле, упала в жалобу земля, бо спустошене збіжжя, вино молоде пересохло, зів'яла оливка.
JOEL|1|11|Засоромилися рільники, голосили були виноградарі за пшеницю й ячмінь, бо вигинуло жниво поля.
JOEL|1|12|Усох виноград, а фіґа зів'яла, гранатове дерево, й пальма та яблуня, і повсихали всі пільні дерева, бо Він висушив радість від людських синів.
JOEL|1|13|Опережіться веретою, і ридайте, священики, голосіть, слуги жертівника, входьте, ночуйте в веретах, служителі Бога мого, бо хлібна жертва і жертва та лита затримана буде від дому вашого Бога!
JOEL|1|14|Оголосіть святий піст, скличте збори, позбирайте старших, всіх мешканців землі до дому Господа, вашого Бога, і кличте до Господа.
JOEL|1|15|Горе дневі тому! Бо близький день Господній, і прийде він від Всемогутнього, мов те спустошення!
JOEL|1|16|Чи ж з-перед очей наших не відіймається їжа, з дому нашого Бога веселість та втіха?
JOEL|1|17|Покорчились зерна під своїми грудами, спорожніли комори, поруйновані клуні, бо висохло збіжжя.
JOEL|1|18|Як стогне товар, поголомшені череди, бо немає їм паші, отари спустошені!
JOEL|1|19|До тебе я кличу, о Господи, пожер бо огонь пасовища пустині, а жар попалив усі дерева на полі.
JOEL|1|20|Навіть пільна худоба прагне до Тебе, бо водні джерела посохли, огонь же пожер пасовища пустині!
JOEL|2|1|Засурміть на Сіоні в сурму, здійміть крик на святій горі Моїй! Затремтіть, всі мешканці землі, бо прийшов день Господній, бо близько вже він,
JOEL|2|2|день темноти та темряви, день хмари й імли! Як несеться досвітня зоря по горах, так народ цей великий й міцний. Такого, як він, не бувало відвіку, і по ньому не буде вже більш аж до літ з роду в рід!
JOEL|2|3|Перед ним пожирає огонь, і палахкотить за ним полум'я! Земля перед ним, як еденський садок, а за ним опустіла пустиня, і рятунку від нього нема!
JOEL|2|4|Його вигляд ніби коні, гарцюють вони, наче ті верхівці!
JOEL|2|5|Як гуркіт військових возів, вони скачуть гірськими верхів'ями, як вереск огнистого полум'я, що солому жере, наче потужний народ, що до бою поставлений.
JOEL|2|6|Народи тремтять перед ним, всі обличчя поблідли.
JOEL|2|7|Як лицарі, мчаться вони, немов вояки вибігають на мур, і кожен своєю дорогою йдуть, і з стежок своїх не позбиваються,
JOEL|2|8|не пхають вони один одного, ходять своєю дорогою битою, а коли на списа упадуть, то не зраняться.
JOEL|2|9|По місті хурчать, по мурі біжать, увіходять в доми, через вікна пролазять, як злодій.
JOEL|2|10|Трясеться земля перед ним, тремтить небо, сонце та місяць темніють, а зорі загублюють сяйво своє.
JOEL|2|11|І голос Свій видасть Господь перед військом Своїм, бо табір Його величезний, бо міцний виконавець слова Його, бо великий день Господа й вельми страшний, і хто зможе його перенести?
JOEL|2|12|Тому то тепер промовляє Господь: Верніться до Мене всім серцем своїм, і постом святим, і плачем та риданням!
JOEL|2|13|І деріть своє серце, а не свою одіж, і наверніться до Господа, вашого Бога, бо ласкавий Він та милосердний, довготерпеливий та многомилостивий, і жалкує за зло!
JOEL|2|14|Хто знає, чи Він не повернеться та не пожалує, і по Собі не залишить благословення, жертву хлібну та жертву ту литу для Господа, вашого Бога.
JOEL|2|15|Засурміть на Сіоні в сурму, оголосіть святий піст, скличте зібрання!
JOEL|2|16|Зберіте народ, оголосіть святі збори, старців згромадьте, позбирайте дітей та грудних немовлят, нехай вийде з кімнати своєї також молодий, молода ж з-під свого накриття!
JOEL|2|17|Між притвором та жертівником нехай плачуть священики, слуги Господні, хай молять вони: Змилуйся, Господи, над народом Своїм, і не видай на ганьбу спадку Свого, щоб над ним панували погани. Нащо будуть казати між народами: Де їхній Бог?
JOEL|2|18|І заздрісним стане Господь за Свій Край, і змилується над народом Своїм.
JOEL|2|19|І Господь відповів і сказав до народу Свого: Ось Я посилаю вам збіжжя й вино молоде та оливу, і насититесь нею, і більше не дам вас на наругу народам.
JOEL|2|20|А цього північного ворога віддалю Я від вас, і його в край сухий та спустошений вижену, його перед до східнього моря, його ж край до того моря заднього. І вийде злий запах його, і підійметься сморід його, бо він лихо велике чинив.
JOEL|2|21|Не бійся ти, земле, а тішся й радій, бо велике Господь учинив!
JOEL|2|22|Не бійтеся, ти пільна худобо, бо пустинні пасовиська зазеленіють, бо дерево видасть свій плід, фіґовниця та виноград свою силу дадуть.
JOEL|2|23|А ви, сіонські сини, радійте та тіштеся Господом, Богом своїм, бо вам їжі Він дасть на спасіння, і найперше зішле вам дощу, дощу раннього й пізнього.
JOEL|2|24|І токи наповняться збіжжям, чавильні ж кадки будуть переливатись вином молодим та оливою.
JOEL|2|25|І надолужу Я вам за ті роки, що пожерла була сарана, коник і черва та гусінь, Моє військо велике, що Я посилав проти вас.
JOEL|2|26|А їсти ви будете їсти й насичуватись, і хвалитимете Ім'я Господа, вашого Бога, що з вами на подив зробив, і посоромлений більше не буде народ Мій навіки!
JOEL|2|27|І пізнаєте ви, що Я серед Ізраїля, і що Я Господь, Бог ваш, і немає вже іншого, і посоромлений більше не буде народ Мій навіки!
JOEL|2|28|(3-1) І буде потому, виллю Я Духа Свого на кожне тіло, і пророкуватимуть ваші сини й ваші дочки, а вашим старим будуть снитися сни, юнаки ваші бачити будуть видіння.
JOEL|2|29|(3-2) І також на рабів та невільниць за тих днів виллю Духа Свого.
JOEL|2|30|(3-3) І дам Я ознаки на небі й землі, кров та огонь, та стовпи диму.
JOEL|2|31|(3-4) Заміниться сонце на темність, а місяць на кров перед приходом Господнього дня, великого та страшного!
JOEL|2|32|(3-5) І станеться, кожен, хто кликати буде Господнє Ім'я, той спасеться, бо на Сіонській горі та в Єрусалимі буде спасіння, як Господь говорив, та для тих позосталих, що Господь їх покличе.
JOEL|3|1|(4-1) Бо ось тими днями та часу того, коли долю Юді та Єрусалиму верну,
JOEL|3|2|(4-2) то зберу всі народи, зведу їх у долину Йосафатову, і там буду судитися з ними за народ Мій й спадщину Мою, за Ізраїля, що його розпорошили поміж народами, а Мій Край поділили.
JOEL|3|3|(4-3) І за народ Мій вони кидали жереба, і юнака за блудницю давали, а дівчину за вино продавали, і пили.
JOEL|3|4|(4-4) І що вам до Мене, Тире й Сидоне, та всі филистимські довкілля? Чи свій чин на Мені надолужите? Може хочете щось учинити Мені, то легко та скоро зверну Я ваш чин вам на голову,
JOEL|3|5|(4-5) що срібло Моє й Моє золото позабирали, а коштовні клейноди Мої в свої храми повносили...
JOEL|3|6|(4-6) А синів Юди та Єрусалиму ви грецьким синам продали, щоб їх віддалити від їхніх границь...
JOEL|3|7|(4-7) Ось Я їх позбуджую з місця того, куди їх продали, ваш чин поверну вам на голову!
JOEL|3|8|(4-8) І попродаю ваших синів та ваших дочок в руку Юдських синів, а вони віддадуть їх шев'янам, до люду далекого, бо Господь так сказав.
JOEL|3|9|(4-9) Кличте про це між народами, оголосіте святую війну, збудіте лицарство, хай сходяться, нехай підіймаються всі вояки.
JOEL|3|10|(4-10) Перекуйте свої лемеші на мечі, а ваші серпи на списи, хай навіть безсилий говорить: Я лицар!
JOEL|3|11|(4-11) Поспішіть і прийдіть, всі народи з довкілля, й зберіться, туди, Господи, спустиш лицарство Своє.
JOEL|3|12|(4-12) Нехай збудяться й зійдуть народи в долину Йосафатову, бо сяду Я там, щоб судити всі народи з довкілля.
JOEL|3|13|(4-13) Пошліть на роботу серпа, бо жниво дозріло, приходьте, зійдіть, бо чавило наповнене, кадки переливаються, бо зло їхнє розмножилось!
JOEL|3|14|(4-14) Натовпи, натовпи у вирішальній долині, бо близький день Господній у вирішальній долині.
JOEL|3|15|(4-15) Сонце та місяць стемніють, а зорі загублять свій блиск,
JOEL|3|16|(4-16) і Господь загримить із Сіону, та з Єрусалиму Свій голос подасть, і небо й земля затремтять, та Господь охорона Своєму народові, і твердиня синам Ізраїлевим!
JOEL|3|17|(4-17) І пізнаєте ви, що Я Господь, Бог ваш, Який пробуває в Сіоні, на святій Своїй горі. І станеться Єрусалим за святиню, і чужі вже не будуть ходити по ньому.
JOEL|3|18|(4-18) І станеться в день той, гори будуть кропити виноградовий сік, а підгірки стоятимуть у молоці, і всі Юдські потоки водою заб'ють, а з дому Господнього вийде джерело, і напоїть долину Шіттім.
JOEL|3|19|(4-19) Єгипет спустошенням стане, і пустинею голою стане Едом за насильство синам Юди, за те, що лили кров невинну у їхньому Краї.
JOEL|3|20|(4-20) А Юдея жити буде повіки, і Єрусалим з роду в рід,
JOEL|3|21|(4-21) і помщу за їхню кров, що за неї Я ще не помстив, і буде Господь пробувати на Сіоні!
