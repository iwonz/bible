2TIM|1|1|奉上帝旨意，按照基督耶稣里所应许的生命，作基督耶稣使徒的 保罗 ，
2TIM|1|2|写信给我亲爱的儿子 提摩太 。愿恩惠、怜悯、平安 从父上帝和我们的主基督耶稣归给你！
2TIM|1|3|我感谢上帝，就是我接续祖先用纯洁的良心所事奉的上帝，在祈祷中昼夜不停地想念你。
2TIM|1|4|我一想起你的眼泪，就急切想见你，好让我满心快乐。
2TIM|1|5|我记得你无伪的信心，这信心先存在你外祖母 罗以 和你母亲 友妮基 的心里，我深信也存在你的心里。
2TIM|1|6|为这缘故，我提醒你要把上帝藉着我按手所给你的恩赐再如火挑旺起来。
2TIM|1|7|因为上帝赐给我们的不是胆怯的心，而是刚强、仁爱、自制的心。
2TIM|1|8|所以，不要以给我们的主作见证为耻，也不要以我这为主被囚的为耻；总要靠着上帝的大能，与我为福音同受苦难。
2TIM|1|9|上帝救了我们， 以圣召召我们， 不是按我们的行为， 而是按他的旨意和恩典； 这恩典是万古之先 在基督耶稣里赐给我们的，
2TIM|1|10|但如今 藉着我们的救主基督耶稣的显现已经表明出来； 他把死废去， 藉着福音，将不朽的生命彰显出来。
2TIM|1|11|我为这福音奉派作传道，作使徒，作教师。
2TIM|1|12|为这缘故，我也受这些苦难。然而，我不以为耻，因为我知道我所信的是谁，也深信他能保全他所交托我的 ，直到那日。
2TIM|1|13|你从我听到那健全的言论，要用在基督耶稣里的信心和爱心常常守着，作为规范。
2TIM|1|14|你要靠着那住在我们里面的圣灵，牢牢守住所交托给你那美好的事。
2TIM|1|15|你知道，所有在 亚细亚 的人都离弃了我，其中有 腓吉路 和 黑摩其尼 。
2TIM|1|16|愿主怜悯 阿尼色弗 一家的人，因为他屡次令我欣慰。他不以我的铁链为耻，
2TIM|1|17|反而一到 罗马 就急切寻找我，并且找到了。
2TIM|1|18|愿主使他在那日能蒙主的怜悯。他在 以弗所 怎样多服事我，你是清楚知道的。
2TIM|2|1|我儿啊，你要在基督耶稣的恩典上刚强起来。
2TIM|2|2|你在许多见证人面前听见我所教导的，也要交托给那忠心而又能教导别人的人。
2TIM|2|3|你要和我同受苦难，作基督耶稣的精兵。
2TIM|2|4|凡当兵的，不让世务缠身，好使那招他当兵的人喜悦。
2TIM|2|5|运动员在比赛的时候，不按规则就不能得冠冕。
2TIM|2|6|勤劳的农夫理当先得粮食。
2TIM|2|7|我所说的话，你要考虑，因为主必在凡事上给你聪明。
2TIM|2|8|要记得耶稣基督，他是 大卫 的后裔，从死人中复活；这就是我所传的福音。
2TIM|2|9|我为这福音受苦难，甚至像犯人一样被捆绑，然而上帝的话没有被捆绑。
2TIM|2|10|所以，我为了选民事事忍耐，为使他们也能得到那在基督耶稣里的救恩和永远的荣耀。
2TIM|2|11|这话是可信的： 我们若与基督同死，也必与他同活；
2TIM|2|12|我们若忍耐到底，也必和他一同作王。 我们若不认他，他也必不认我们；
2TIM|2|13|我们纵然失信，他仍是可信的， 因为他不能否认自己。
2TIM|2|14|你要向众人提醒这些事，在上帝 面前嘱咐他们不可在言词上争辩；这是没有益处的，只能伤害听的人。
2TIM|2|15|你当竭力在上帝面前作一个经得起考验、无愧的工人，按着正意讲解真理的话。
2TIM|2|16|要远避世俗的空谈，因为这等空谈会使人进到更不敬虔的地步。
2TIM|2|17|他们的话如同毒疮越烂越大；其中有 许米乃 和 腓理徒 ，
2TIM|2|18|他们偏离了真理，说复活的事已过去，败坏了好些人的信心。
2TIM|2|19|然而，上帝坚固的根基屹立不移；上面有这印记说：“主认得他自己的人”，又说：“凡称呼主名的人总要离开不义。”
2TIM|2|20|大户人家不但有金器银器，也有木器瓦器；有作为贵重之用的，有作为卑贱之用的。
2TIM|2|21|人若自洁，脱离卑贱的事，必成为贵重的器皿，成为圣洁，合乎主用，预备行各样的善事。
2TIM|2|22|你要逃避年轻人的私欲，同那以纯洁的心求告主的人追求公义、信实、仁爱、和平。
2TIM|2|23|但要弃绝那愚拙无知的辩论，因为你知道这等事只会引起争辩。
2TIM|2|24|主的仆人不可争辩，只要温和待人，善于教导，恒心忍耐，
2TIM|2|25|用温柔劝导反对的人。也许上帝会给他们悔改的心能明白真理，
2TIM|2|26|让他们这些已被魔鬼掳去顺从他诡计的人能醒悟过来，脱离他的罗网。
2TIM|3|1|你该知道，末世必有艰难的日子来到。
2TIM|3|2|那时人会专爱自己，贪爱钱财，自夸，狂傲，毁谤，违背父母，忘恩负义，心不圣洁，
2TIM|3|3|没有亲情，抗拒和解，好说谗言，不能节制，性情凶暴，不爱良善，
2TIM|3|4|卖主卖友，任意妄为，自高自大，爱好宴乐，不爱上帝，
2TIM|3|5|有敬虔的外貌，却背弃了敬虔的实质，这等人你要避开。
2TIM|3|6|他们当中有人潜入别人家里，操纵无知的妇女；这些妇女被罪恶压制，被各样的私欲引诱，
2TIM|3|7|虽然常常学习，终久无法达到明白真理的地步。
2TIM|3|8|从前 雅尼 和 佯庇 怎样反对 摩西 ，这等人也怎样抵挡真理；他们的心地败坏，信仰经不起考验。
2TIM|3|9|然而，他们没有进步，因为他们的愚昧必在众人面前显露出来，像那两人一样。
2TIM|3|10|但你已经追随了我的教导、行为、志向、信心、宽容、爱心、忍耐，
2TIM|3|11|以及我在 安提阿 、 以哥念 、 路司得 所遭遇的迫害和苦难。我忍受了何等的迫害！但从这一切苦难中，主都把我救了出来。
2TIM|3|12|其实，凡立志在基督耶稣里敬虔度日的，也都将受迫害。
2TIM|3|13|只是作恶的和骗人的将变本加厉，迷惑人也被人迷惑。
2TIM|3|14|至于你，你要持守所学习的和所确信的，因为你知道是跟谁学的，
2TIM|3|15|并且知道你从小明白圣经，这圣经能使你因在基督耶稣里的信 有得救的智慧。
2TIM|3|16|圣经都是上帝所默示的 ，于教训、督责、使人归正、教导人学义都是有益的，
2TIM|3|17|叫属上帝的人得以完全，预备行各样的善事。
2TIM|4|1|我在上帝面前，并在将来审判活人死人的基督耶稣面前，凭着他的显现和他的国度郑重地劝戒你：
2TIM|4|2|务要传道；无论得时不得时总要专心，并以百般的忍耐和各样的教导责备人，警戒人，劝勉人。
2TIM|4|3|因为时候将到，那时人会厌烦健全的教导，耳朵发痒，就随心所欲地增添好些教师，
2TIM|4|4|并且掩耳不听真理，偏向无稽的传说。
2TIM|4|5|至于你，凡事要谨慎，忍受苦难，做传福音的工作，尽你的职分。
2TIM|4|6|至于我，我已经被浇献，离世的时候到了。
2TIM|4|7|那美好的仗我已经打过了，当跑的路我已经跑尽了，该信的道我已经守住了。
2TIM|4|8|从此以后，有公义的冠冕为我存留，就是按着公义审判的主到了那日要赐给我的；不但赐给我，也赐给凡爱慕他显现的人。
2TIM|4|9|你要赶紧到我这里来。
2TIM|4|10|因为 底马 贪爱现今的世界，已经离弃我，往 帖撒罗尼迦 去了； 革勒士 往 加拉太 去； 提多 往 挞马太 去；
2TIM|4|11|只有 路加 在我这里。你来的时候把 马可 带来，因为他在服事 上于我有益。
2TIM|4|12|我已经打发 推基古 往 以弗所 去。
2TIM|4|13|我在 特罗亚 留给 加布 的那件外衣，你来的时候要带来，那些书也带来，特别是那几卷羊皮的书。
2TIM|4|14|铜匠 亚历山大 多方害我；主必照他所行的报应他。
2TIM|4|15|你也要防备他，因为他极力抗拒我们的话。
2TIM|4|16|我初次上诉时，没有人前来帮助，竟都离弃了我，但愿这罪不归在他们身上。
2TIM|4|17|惟有主站在我身边，加给我力量，使我能把福音完整地传开，让所有的外邦人都听见；我也从狮子口里被救出来。
2TIM|4|18|主必救我脱离一切的凶恶，也必救我进他的天国。愿荣耀归给他，直到永永远远。阿们！
2TIM|4|19|请向 百基拉 、 亚居拉 和 阿尼色弗 一家的人问安。
2TIM|4|20|以拉都 在 哥林多 住下了。 特罗非摩 病了，我把他留在 米利都 。
2TIM|4|21|你要赶紧在冬天以前到我这里来。 友布罗 、 布田 、 利奴 、 革老底亚 和众弟兄都向你问安。
2TIM|4|22|愿主与你的灵同在！愿恩惠与你们同在！
