1TIM|1|1|奉我们的救主上帝，和我们的盼望基督耶稣的命令，作基督耶稣使徒的 保罗 ，
1TIM|1|2|写信给那因信主作我真儿子的 提摩太 。愿恩惠、怜悯、平安 从父上帝和我们主基督耶稣归给你！
1TIM|1|3|我往 马其顿 去的时候，曾劝你留在 以弗所 ，好嘱咐某些人不可传别的教义，
1TIM|1|4|也不要听从无稽的传说和冗长的家谱；这样的事只会引起争论，无助于上帝的计划，这计划是凭着信才能了解的。
1TIM|1|5|但命令的目的就是爱；这爱是出于清洁的心、无愧的良心和无伪的信心。
1TIM|1|6|有人偏离了这些而转向空谈，
1TIM|1|7|想要作律法教师，却不明白自己所讲的是什么，也不知道所主张的是什么。
1TIM|1|8|我们知道，只要人善用律法，律法是好的；
1TIM|1|9|因为知道律法不是为义人订立的，而是为不法和叛逆的，不虔诚和犯罪的，不圣洁和恋世俗的，弑父母和杀人的，
1TIM|1|10|犯淫乱和亲男色的，拐卖人口和说谎话的，并起假誓的，或是为任何违背健全教义的事订立的。
1TIM|1|11|这是按照可称颂、荣耀之上帝交托我的福音说的。
1TIM|1|12|我感谢那赐给我力量的我们的主基督耶稣，因为他认为我可信任，派我服事他。
1TIM|1|13|我从前是亵渎、迫害、侮慢上帝的人；然而我还蒙了怜悯，因为我是在不信、不明白的时候做的。
1TIM|1|14|而且我们的主的恩典格外丰盛，使我在基督耶稣里有信心和爱心。
1TIM|1|15|这话可信，值得完全接受：“基督耶稣到世上来是要拯救罪人”，而在罪人中我是个罪魁。
1TIM|1|16|然而，我蒙了怜悯，好让基督耶稣在我这罪魁身上显明他完全的忍耐，给后来信他得永生的人作榜样。
1TIM|1|17|愿尊贵、荣耀归给永世的君王，那不朽坏、看不见、独一的上帝，直到永永远远。阿们！
1TIM|1|18|我儿 提摩太 啊，我照从前指着你的预言把这命令交托你，使你能藉着这些预言打那美好的仗，
1TIM|1|19|常存信心和无愧的良心。有些人丢弃良心，在信仰上触了礁；
1TIM|1|20|其中有 许米乃 和 亚历山大 ，我已经把他们交给撒但，让他们学会不再亵渎。
1TIM|2|1|所以，我劝你，首先要为人人祈求、祷告、代求、感谢；
1TIM|2|2|为君王和一切在位的，也要如此，使我们能够敬虔端正地过平稳宁静的生活。
1TIM|2|3|这是好的，在我们的救主上帝面前可蒙悦纳。
1TIM|2|4|他愿意人人得救，并得以认识真理。
1TIM|2|5|因为只有一位上帝， 在上帝和人之间也只有一位中保， 是成为人的基督耶稣。
1TIM|2|6|他献上自己作人人的赎价； 在适当的时候这事已经证实了。
1TIM|2|7|我为此奉派作传道，作使徒，在信仰和真理上作外邦人的教师。我说的是真话，不是说谎。
1TIM|2|8|我希望男人举起圣洁的手随处祷告，不发怒，不争论。
1TIM|2|9|我也希望女人以端正、克制和合乎体统的服装打扮自己，不以编发、金饰、珍珠和名贵衣裳来打扮。
1TIM|2|10|要有善行，这才与自称为敬畏上帝的女人相称。
1TIM|2|11|女人要事事顺服地安静学习。
1TIM|2|12|我不许女人教导，也不许她管辖男人，只要安静。
1TIM|2|13|因为 亚当 先被造，然后才是 夏娃 ；
1TIM|2|14|亚当 并没有受骗，而是女人受骗，陷在过犯里。
1TIM|2|15|然而，女人若持守信心、爱心，又圣洁克制，就必藉着生产而得救。
1TIM|3|1|“若有人想望监督的职分，他是在羡慕一件好事”，这话是可信的。
1TIM|3|2|监督必须无可指责，只作一个妇人的丈夫，有节制、克己、端正，乐意接待外人，善于教导，
1TIM|3|3|不酗酒，不打人；要温和，不好斗，不贪财。
1TIM|3|4|要好好管理自己的家，使儿女顺服，凡事庄重。
1TIM|3|5|人若不知道管理自己的家，怎能照管上帝的教会呢？
1TIM|3|6|刚信主的，不可作监督，恐怕他自高自大，落在魔鬼所受的惩罚里。
1TIM|3|7|监督也必须在教外有好名声，免得被人毁谤，落在魔鬼的罗网里。
1TIM|3|8|同样，执事也必须庄重，不一口两舌，不好酒，不贪不义之财；
1TIM|3|9|要存清白的良心固守信仰的奥秘。
1TIM|3|10|这些人也要先受考验，若没有可责之处，才让他们作执事。
1TIM|3|11|同样，女执事 也必须庄重，不说闲话，有节制，凡事忠心。
1TIM|3|12|执事只作一个妇人的丈夫，要好好管儿女和自己的家。
1TIM|3|13|因为善于作执事的，为自己得到美好的地位，并且无惧地坚信在基督耶稣里的信仰。
1TIM|3|14|我希望尽快到你那里去，所以先把这些事写给你；
1TIM|3|15|倘若我延误了，你也可以知道在上帝的家中该怎样做。这家就是永生上帝的教会，真理的柱石和根基。
1TIM|3|16|敬虔的奥秘是公认为伟大的： 上帝在肉身显现， 被圣灵称义， 被天使看见， 被传于外邦， 被世人信服， 被接在荣耀里。
1TIM|4|1|圣灵明说，在末后的时期必有人离弃信仰，去听信那诱惑人的邪灵和鬼魔的教训。
1TIM|4|2|这是出于撒谎者的假冒；这些人的良心如同被热铁烙了一般。
1TIM|4|3|他们禁止嫁娶，又禁戒食物—就是上帝所造、让那信而明白真理的人存感谢的心领受的。
1TIM|4|4|上帝所造之物样样都是好的，若存感谢的心领受，没有一样是不可吃的，
1TIM|4|5|都因上帝的话和人的祈祷而成为圣洁了。
1TIM|4|6|你若把这些事提醒弟兄们，就是基督耶稣的好执事，在信仰的话语和你向来所服从的正确教义上得到了栽培。
1TIM|4|7|要弃绝那世俗的言语和老妇的无稽传说。要在敬虔上操练自己：
1TIM|4|8|因操练身体有些益处；但敬虔在各方面都有益，它有现今和未来的生命的应许。
1TIM|4|9|这话可信，值得完全接受。
1TIM|4|10|我们劳苦，努力 正是为此，因为我们的指望在乎永生的上帝。他是人人的救主，更是信徒的救主。
1TIM|4|11|你要嘱咐和教导这些事。
1TIM|4|12|不可叫人小看你年轻，总要在言语、行为、爱心、信心、清洁上，都作信徒的榜样。
1TIM|4|13|要以宣读圣经，劝勉，教导为念，直等到我来。
1TIM|4|14|不要忽略你所得的恩赐，就是从前藉着预言、在众长老按手的时候赐给你的。
1TIM|4|15|这些事你要殷勤去做，并要在这些事上专心，让众人看出你的长进来。
1TIM|4|16|要谨慎自己和自己的教导，要在这些事上恒心，因为这样做，既能救自己，又能救听你的人。
1TIM|5|1|不可严责老年人，要劝他如同父亲。要待年轻人如同弟兄，
1TIM|5|2|年老妇女如同母亲。要清清洁洁地待年轻妇女如同姊妹。
1TIM|5|3|要尊敬真正守寡的妇人。
1TIM|5|4|寡妇若有儿女，或有孙儿女，要让儿孙先在自己家中学习行孝，报答亲恩，因为这在上帝面前是可蒙悦纳的。
1TIM|5|5|独居无靠的真寡妇只仰赖上帝，昼夜不住地祈求祷告。
1TIM|5|6|但好宴乐的寡妇活着也算是死了。
1TIM|5|7|这些事，你要嘱咐她们，让她们无可指责。
1TIM|5|8|若有人不照顾亲属，尤其是自己家里的人，就是背弃信仰，还不如不信的人。
1TIM|5|9|寡妇登记，年龄必须在六十岁以上，只作一个丈夫的妻子，
1TIM|5|10|又有行善的名声，就如养育儿女，收留外人，洗圣徒的脚，救济遭难的人，竭力行各样善事。
1TIM|5|11|至于年轻的寡妇，你要拒绝登记，因为她们情欲冲动、背弃基督的时候，就想嫁人，
1TIM|5|12|她们因废弃了当初所许的愿而被定罪。
1TIM|5|13|同时，她们又学了懒惰，习惯于挨家闲逛；不但懒惰，而且说长道短，好管闲事，说些不该说的话。
1TIM|5|14|所以，我希望年轻的寡妇嫁人，生养儿女，治理家务，不让敌人有辱骂的把柄，
1TIM|5|15|因为已经有一些人转去随从撒但了。
1TIM|5|16|信主的妇女若有亲戚是寡妇，要救济她们，不可拖累教会，好使教会能救济真正无助的寡妇。
1TIM|5|17|善于督导教会的长老，尤其是勤劳讲道教导人的，应该得到加倍的敬奉。
1TIM|5|18|因为经上说：“牛在踹谷的时候，不可笼住它的嘴”；又说：“工人得工资是应当的。”
1TIM|5|19|有控告长老的案件，非有两三个证人就不要受理。
1TIM|5|20|继续犯罪的人，要在众人面前责备他，使其余的人也有所惧怕。
1TIM|5|21|我在上帝、基督耶稣和蒙拣选的天使面前嘱咐你要遵守这些话，不可存成见，做事也不可偏心。
1TIM|5|22|不可急于给人行按手礼；也不可在别人的罪上有份，要保守自己纯洁。
1TIM|5|23|为了你的胃，又常患病，不要只喝水，要稍微喝点酒。
1TIM|5|24|有些人的罪是明显的，已先受审判了；有些人的罪是随后跟着来。
1TIM|5|25|同样，善行也有明显的，就是那不明显的也不能隐藏。
1TIM|6|1|凡负轭作奴隶的，要认为自己的主人配受各样的尊敬，免得上帝的名和教导被人亵渎。
1TIM|6|2|奴隶若有信主的主人，不可因他是主内弟兄就轻看他们，更要越发服侍他们，因为得到服侍的益处的正是信徒，是蒙爱的人。 你要教导人和劝勉这些事。
1TIM|6|3|若有人传别的教义，不符合我们主耶稣基督纯正的话语与合乎敬虔的教导，
1TIM|6|4|他是自高自大，一无所知，专好争辩，擅于舌战，因而生出嫉妒、纷争、毁谤、恶意猜疑，
1TIM|6|5|和心术不正与丧失真理的人不停地争吵，以敬虔为得利的门路。
1TIM|6|6|其实，敬虔加上知足就是大利。
1TIM|6|7|因为我们没有带什么到世上来， 也不能带什么去；
1TIM|6|8|只要有衣有食， 我们就该知足。
1TIM|6|9|但那些想要发财的人就陷在诱惑、罗网和许多无知有害的欲望中，使人沉沦，以致败坏和灭亡。
1TIM|6|10|贪财是万恶之根。有人因贪恋钱财而背离信仰，用许多愁苦把自己刺透了。
1TIM|6|11|但你这属上帝的人哪，要逃避这些事；要追求公义、敬虔、信心、爱心、忍耐、温柔。
1TIM|6|12|你要为信仰打那美好的仗；要持定永生，你为此被召，也已经在许多见证人面前作了那美好的见证。
1TIM|6|13|我在那赐生命给万物的上帝面前，并在向 本丢．彼拉多 作过那美好见证的基督耶稣面前嘱咐你 ：
1TIM|6|14|要守这命令，毫不玷污，无可指责，直到我们的主耶稣基督显现。
1TIM|6|15|到了适当的时候都要显明出来： 他是那可称颂、独一的权能者， 万王之王， 万主之主，
1TIM|6|16|就是那独一不死、 住在人不能靠近的光里， 是人未曾看见，也是不能看见的。 愿尊贵和永远的权能都归给他。阿们！
1TIM|6|17|至于那些今世富足的人，你要嘱咐他们不要自高，也不要倚赖靠不住的钱财；要倚靠那厚赐万物给我们享受的上帝。
1TIM|6|18|又要嘱咐他们行善，在好事上富足，甘心施舍，乐意分享，
1TIM|6|19|为自己积存财富，而为将来打美好的根基，好使他们能把握那真正的生命。
1TIM|6|20|提摩太 啊，要持守所给你的托付。要躲避世俗的空谈和那假冒知识的矛盾言论。
1TIM|6|21|有人自称有这知识而偏离了信仰。 愿恩惠与你们同在！
