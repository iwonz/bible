JOSH|1|1|І сталося по смерті Мойсея, раба Божого, і сказав Господь до Ісуса, сина Навинового, Мойсеєвого слуги, говорячи:
JOSH|1|2|Мойсей, раб Мій, помер. А тепер уставай, перейди цей Йордан ти та ввесь народ цей до того Краю, що Я даю їм, Ізраїлевим синам.
JOSH|1|3|Кожне місце, що стопа ноги вашої ступить на ньому, Я дав вам, як Я говорив був Мойсеєві.
JOSH|1|4|Від пустині й цього Ливану й аж до Великої Річки, річки Ефрату, увесь край хіттеян, і аж до Великого моря на захід буде ваша границя.
JOSH|1|5|Не встоїть ніхто перед тобою по всі дні життя твого. Як був Я з Мойсеєм, так буду з тобою, не залишу тебе й не покину тебе.
JOSH|1|6|Будь сильний та відважний, бо ти зробиш, що народ цей посяде той Край, що Я присягнув був їхнім батькам дати їм.
JOSH|1|7|Тільки будь дуже сильний та відважний, щоб додержувати чинити за всім тим Законом, що наказав був тобі Мойсей, Мій раб, не відхилишся від нього ні праворуч, ні ліворуч, щоб щастило тобі в усьому, де ти будеш ходити.
JOSH|1|8|Нехай книга цього Закону не відійде від твоїх уст, але будеш роздумувати про неї вдень та вночі, щоб додержувати чинити все, що написано в ній, бо тоді зробиш щасливими дороги свої, і тоді буде щастити тобі.
JOSH|1|9|Чи ж не наказав Я тобі: будь сильний та відважний? Не бійся й не лякайся, бо з тобою Господь, Бог твій, у всьому, де ти будеш ходити.
JOSH|1|10|І наказав Ісус урядникам народу, говорячи:
JOSH|1|11|Перейдіть посеред табору, і накажіть народові, говорячи: Приготуйте собі поживу на дорогу, бо по трьох днях ви переходите цей Йордан, щоб увійти посісти той Край, що Господь, Бог ваш, дає вам його на спадщину.
JOSH|1|12|А Рувимовому й Ґадовому та половині племени Манасіїного Ісус сказав, говорячи:
JOSH|1|13|Пам'ятайте те слово, що вам наказав був Мойсей, раб Господній, говорячи: Господь, Бог ваш, що відпочинок дає вам, дав вам цей Край.
JOSH|1|14|Ваші жінки, діти ваші та ваша худоба зостануться в Краї, що дав вам Мойсей по той бік Йордану, а ви перейдете озброєні перед вашими братами, усі сильні військові, і допоможете їм,
JOSH|1|15|аж поки Господь не дасть відпочинку вашим братам, як вам, і посядуть і вони той Край, що Господь, Бог ваш, дає їм. І ви вернетеся до Краю вашого спадку, і посядете його, що дав вам Мойсей, раб Господній, по той бік Йордану на схід сонця.
JOSH|1|16|А вони відповіли Ісусові, говорячи: Усе, що накажеш нам, ми зробимо, і до всього, куди пошлеш нас, підемо.
JOSH|1|17|Усе так, як слухалися ми Мойсея, так будемо слухатися тебе, тільки нехай буде Господь, Бог твій, з тобою, як був Він із Мойсеєм.
JOSH|1|18|Кожен, хто буде неслухняний наказам твоїм, і не буде слухатися слів твоїх щодо всього, що накажеш йому, нехай буде вбитий. Тільки будь сильний та відважний!
JOSH|2|1|І послав Ісус, син Навинів, із Ситтіму двох таємних вивідувачів, говорячи: Ідіть, розгляньте цей Край та Єрихон. І вони пішли, і ввійшли до дому однієї блудниці, а ім'я їй Рахав. І переночували вони там.
JOSH|2|2|І було донесено єрихонському цареві, говорячи: Ось цієї ночі прийшли сюди якісь люди з Ізраїлевих синів, щоб вивідати цей Край.
JOSH|2|3|І послав єрихонський цар до Рахави, говорячи: Виведи тих людей, що до тебе прийшли, що ввійшли до твого дому, бо вони прийшли, щоб вивідати ввесь цей Край.
JOSH|2|4|А та жінка взяла двох тих людей, та й сховала їх. І сказала: Так, приходили були до мене ті люди, та я не знала, звідки вони.
JOSH|2|5|А коли замикалася брама зо смерком, то ті люди вийшли. Не знаю, куди ті люди пішли. Швидко женіться за ними, то ви доженете їх.
JOSH|2|6|А вона відвела їх на дах, та й сховала їх у жмутах льону, що були зложені в неї на даху.
JOSH|2|7|А ті люди погналися за ними йорданською дорогою аж до бродів; а браму замкнули, як тільки вийшла погоня за ними.
JOSH|2|8|І поки вони лягли спати, то вона ввійшла до них на дах,
JOSH|2|9|і сказала до тих людей: Я знаю, що Господь дав вам цей Край, і що жах перед вами напав на нас, і що всі мешканці цього Краю умлівають зо страху перед вами.
JOSH|2|10|Бо ми чули те, що Господь висушив воду Червоного моря перед вами, коли ви виходили з Єгипту, і що зробили ви обом аморейським царям, що по той бік Йордану, Сигонові та Оґові, яких ви вчинили закляттям.
JOSH|2|11|І чули ми це, і зомліло наше серце, і не стало вже духу в людини зо страху перед вами, бо Господь, Бог ваш, Він Бог на небесах угорі й на землі долі!
JOSH|2|12|А тепер присягніть мені Господом, що як я вчинила з вами милість, так зробите й ви милість з домом батька мого, і дасте мені правдивого знака.
JOSH|2|13|І зоставите при житті батька мого, і матір мою, і братів моїх, і сестер моїх, і все, що їхнє, і врятуєте наше життя від смерти.
JOSH|2|14|І сказали їй ті люди: Душа наша за вас нехай віддана буде на смерть, якщо ви не відкриєте цієї нашої справи. І буде, коли Господь передаватиме нам оцей Край, то ми вчинимо тобі милість та правду.
JOSH|2|15|І вона спустила їх шнуром через вікно, бо дім її був у стіні міського муру, і в мурі вона жила.
JOSH|2|16|І сказала вона їм: Ідіть на гору, щоб не спіткала вас погоня. І ховайтеся там три дні, аж поки не вернеться погоня, а потому підете своєю дорогою.
JOSH|2|17|І сказали до неї ті люди: Ми будемо чисті від цієї присяги тобі, що ти заприсягла нас, якщо ти не вчиниш так.
JOSH|2|18|Оце, як ми будемо входити до Краю, то ти прив'яжеш шнурка з цієї нитки червені в вікні, що ти ним нас спустила. А батька свого, і матір свою, і братів своїх, і ввесь дім свого батька збереш до себе до дому.
JOSH|2|19|І буде, усі, хто вийде з дверей твого дому назовні, кров його на голові його, а ми чисті. А всі, хто буде в домі з тобою, кров його на голові нашій, якщо наша рука буде на ньому.
JOSH|2|20|А коли ти відкриєш цю нашу справу, то ми будемо чисті від присяги тобі, якою ти заприсягла нас.
JOSH|2|21|А вона сказала: Як ви сказали, нехай буде воно так. І відпустила їх, а вони пішли. І вона прив'язала в вікні червоного суканого шнурка.
JOSH|2|22|І вони пішли, і вийшли на гору, та й сиділи там три дні, аж поки вернулася погоня. І шукала погоня по всій дорозі, та не знайшла їх.
JOSH|2|23|І повернулися ті два мужі, і зійшли з гори, і перейшли Йордан, і прийшли до Ісуса, сина Навинового, та й розповіли йому все, що їх спіткало.
JOSH|2|24|І сказали вони до Ісуса: Справді Господь дав у нашу руку всю цю землю, а всі мешканці цього Краю омліли зо страху перед нами.
JOSH|3|1|І встав Ісус рано вранці, і вони рушили з Ситтіму, та й прийшли аж до Йордану він та всі Ізраїлеві сини. І переночували вони там перше, ніж перейшли.
JOSH|3|2|І сталося по трьох днях, і перейшли урядники між табором,
JOSH|3|3|і наказали народові, говорячи: Коли ви побачите ковчега заповіту Господа, Бога вашого, та священиків-Левитів, що несуть його, то ви рушите з вашого місця, і підете за ним.
JOSH|3|4|Тільки віддаль між вами та між ним буде мірою коло двох тисяч ліктів. Не наближайтеся до нього, щоб ви знали ту дорогу, якою підете, бо ви не ходили цією дорогою ані вчора, ані позавчора.
JOSH|3|5|І сказав Ісус до народу: Освятіться, бо Господь узавтра чинитиме чуда поміж вами.
JOSH|3|6|І сказав Ісус до священиків, говорячи: Понесіть ковчега заповіту, і перейдіть Йордан перед народом. І понесли вони ковчега заповіту, і пішли перед народом.
JOSH|3|7|І сказав Господь до Ісуса: Цього дня розпічну Я звеличувати тебе на очах усього Ізраїля, який буде бачити, що як був Я з Мойсеєм, так буду з тобою.
JOSH|3|8|А ти накажеш священикам, що носять ковчега заповіту, говорячи: Коли ви ввійдете до краю води Йордану, станете в Йордані.
JOSH|3|9|І сказав Ісус до Ізраїлевих синів: Підійдіть сюди, і послухайте слів Господа, Бога вашого.
JOSH|3|10|І Ісус сказав: По цьому пізнаєте, що Бог Живий поміж вами, і конче Він вижене перед вами ханаанеянина, і хіттеянина, і хіввеянина, і періззеянина, і ґірґашеянина, і євусеянина.
JOSH|3|11|Оце ковчег заповіту Владики всієї землі переходить перед вами через Йордан.
JOSH|3|12|А тепер візьміть собі дванадцять мужів з Ізраїлевих племен, по одному мужеві на плем'я.
JOSH|3|13|І станеться, коли спиняться стопи ніг священиків, що носять ковчега Господа, Владики всієї землі, у воді Йордану, буде спинена вода, що тече зверху, і стане одним валом.
JOSH|3|14|І сталося, коли рушив народ зо своїх наметів, щоб перейти Йордан, а священики, що несли ковчега заповіту перед народом,
JOSH|3|15|і коли носії ковчегу прийшли до Йордану, а ноги священиків, що несли ковчега, занурилися в воду скраю, а Йордан був повний по всі береги свої всі дні жнив,
JOSH|3|16|то спинилась вода, що зверху текла, стала одним валом, дуже далеко від міста Адама, що збоку Цортану, а та, що текла до степу, до Солоного моря, стекла зовсім, і була відділена, а народ перейшов навпроти Єрихону.
JOSH|3|17|А священики, що несли ковчега заповіту Господнього, стали міцно на сухому посередині Йордану, і ввесь Ізраїль переходив по сухому, аж поки не скінчив переходити Йордан увесь народ.
JOSH|4|1|І сталося, як увесь народ закінчив переходити Йордан, то сказав Господь до Ісуса, говорячи:
JOSH|4|2|Візьміть собі з народу дванадцять мужів, по одному мужеві з племени.
JOSH|4|3|І накажете їм, говорячи: Винесіть звідси, із середини Йордану, із місця, де міцно стояли ноги священиків, дванадцять каменів, і перенесете їх із собою, і покладете їх на нічлігу, що в ньому будете ночувати цієї ночі.
JOSH|4|4|І покликав Ісус тих дванадцятьох мужів, що настановив з Ізраїлевих синів, по одному мужеві з племени,
JOSH|4|5|та й сказав їм Ісус: Підіть перед ковчегом Господа, Бога вашого, до середини Йордану, і підійміть собі кожен на плече своє одного каменя за числом племен Ізраїлевих синів,
JOSH|4|6|щоб то було знаком між вами, коли взавтра запитають ваші сини, говорячи: Що це в вас за каміння?
JOSH|4|7|то скажете їм, що була відділена йорданська вода перед ковчегом Господнього заповіту, коли він переходив в Йордані, була відділена йорданська вода. І будуть ті каміння за пам'ятку для Ізраїлевих синів аж навіки.
JOSH|4|8|І зробили Ізраїлеві сини так, як наказав Ісус, і понесли вони дванадцять каменів із середини Йордану, як говорив Господь до Ісуса, за числом племен Ізраїлевих синів. І перенесли їх із собою до нічлігу, та й поклали їх там.
JOSH|4|9|А інших дванадцять каменів поставив Ісус в середині Йордану на місці, де стояли ноги священиків, що несли ковчега заповіту, і вони там аж до дня цього.
JOSH|4|10|А священики, що несли ковчега, стояли в середині Йордану аж до закінчення всього, що Господь наказав був Ісусові сказати народові, згідно з усім тим, що наказав був Мойсей Ісусові. А народ квапився і переходив.
JOSH|4|11|І сталося, як увесь народ скінчив переходити, то перейшов Господній ковчег та священики перед народом.
JOSH|4|12|І перейшли Рувимові сини й сини Ґадові та половина племени Манасіїного, озброєні до бою, перед Ізраїлевими синами, як Мойсей говорив був до них.
JOSH|4|13|Коло сорока тисяч озброєних вояків перейшли перед Господнім лицем на війну до єрихонських степів.
JOSH|4|14|Того дня звеличив Господь Ісуса на очах усього Ізраїля, і стали боятися його, як боялися Мойсея по всі дні його життя.
JOSH|4|15|І сказав Господь до Ісуса, говорячи:
JOSH|4|16|Накажи священикам, що носять ковчега заповіту, і нехай вони вийдуть з Йордану.
JOSH|4|17|І наказав Ісус священикам, говорячи: Вийдіть з Йордану!
JOSH|4|18|І сталося, коли священики, що несли ковчега Господнього заповіту, вийшли з середини Йордану, а стопи ніг священиків відірвалися від нього, щоб стати на сухому, то вода Йордану вернулася на своє місце, і пішла, як учора-позавчора, по всіх його берегах.
JOSH|4|19|А народ вийшов із Йордану десятого дня першого місяця, та й таборував у Ґілґалі, на східньому боці Єрихону.
JOSH|4|20|А дванадцять тих каменів, що взяли з Йордану, Ісус поставив у Ґілґалі.
JOSH|4|21|І сказав він до Ізраїлевих синів, говорячи: Коли взавтра запитають вас ваші сини своїх батьків, говорячи: Що це за каміння?
JOSH|4|22|то познайомте ваших синів, говорячи: По сухому перейшов був Ізраїль цей Йордан,
JOSH|4|23|бо Господь, Бог ваш, висушив воду Йордану перед вами, аж поки ви не перейшли, як зробив був Господь, Бог ваш, морю Червоному, яке Він висушив перед нами, аж поки ми не перейшли,
JOSH|4|24|щоб усі народи землі пізнали руку Господню, що сильна вона, щоб боялися ви Господа, Бога вашого, по всі дні.
JOSH|5|1|І сталося, як усі аморейські царі, що по той бік Йордану на захід, і всі ханаанські царі, що над морем, почули, що Господь висушив був воду Йордану перед Ізраїлевими синами, аж поки вони перейшли, то зомліло їхнє серце, і не було вже в них духу зо страху перед Ізраїлевими синами.
JOSH|5|2|Того часу сказав Господь до Ісуса: Нароби собі камінних ножів, і пообрізуй Ізраїлевих синів знову, другий раз.
JOSH|5|3|І наробив собі Ісус камінних ножів, та й пообрізував Ізраїлевих синів при Ґів'ат-Гааралоті.
JOSH|5|4|А оце та причина, чому Ісус пообрізував: увесь народ, що вийшов був із Єгипту, чоловічої статі, усі вояки, повмирали в пустині в дорозі, коли вийшли з Єгипту.
JOSH|5|5|Бо був обрізаний увесь народ, що виходив, а всього народу, що народився в пустині в дорозі по виході з Єгипту, не обрізували.
JOSH|5|6|Бо сорок літ ходили Ізраїлеві сини в пустині, аж поки не вигинув увесь той народ, ті вояки, що вийшли були з Єгипту, що не слухалися Господнього голосу, що Господь заприсягнув був їм не показати їм того Краю, що Господь заприсягнув був їхнім батькам дати їм Край, який тече молоком та медом.
JOSH|5|7|А їхніх синів поставив замість них. Їх пообрізував Ісус, бо вони були необрізані, бо їх не обрізували в дорозі.
JOSH|5|8|І сталося, як увесь народ закінчив обрізуватися, то вони осіли в таборі на своїх місцях аж до видужання.
JOSH|5|9|І сказав Господь до Ісуса: Сьогодні Я зняв з вас єгипетську ганьбу. І назвав те місце ім'ям: Ґілґал, і так є аж до цього дня.
JOSH|5|10|І таборували Ізраїлеві сини в Ґілґалі, і справили Пасху ввечорі чотирнадцятого дня місяця на єрихонських степах.
JOSH|5|11|А назавтра по Пасці їли вони того самого дня з урожаю того Краю, опрісноки та пражене.
JOSH|5|12|І перестала падати манна з другого дня, як вони їли з урожаю того Краю, і вже більш не було Ізраїлевим синам манни, і їли вони того року з урожаю ханаанського Краю.
JOSH|5|13|І сталося, коли Ісус був при Єрихоні, то звів очі свої та й побачив, аж ось стоїть навпроти нього чоловік, а витягнений його меч у руці його. І підійшов Ісус до нього, та й сказав йому: Чи ти наш, чи наших ворогів?
JOSH|5|14|А той відказав: Ні, бо я вождь Господнього війська, тепер я прийшов. І впав Ісус на обличчя своє до землі, і вклонився, та й сказав йому: Що говорить мій пан своєму рабові?
JOSH|5|15|І сказав вождь Господнього війська до Ісуса: Скинь взуття своє з своїх ніг, бо це місце, на якому стоїш ти, святе воно! І зробив Ісус так.
JOSH|6|1|А Єрихон замкнувся, і був замкнений зо страху перед Ізраїлевими синами, ніхто не виходив і не входив.
JOSH|6|2|І сказав Господь до Ісуса: Ось, Я дав у твою руку Єрихон та царя його, сильних вояків.
JOSH|6|3|І обійдете навколо це місто, всі вояки, обхід навколо міста один раз. Так зробиш шість день.
JOSH|6|4|А сім священиків будуть нести сім сурем із баранячих рогів перед ковчегом. А сьомого дня обійдете навколо те місто сім раз, а священики засурмлять у роги.
JOSH|6|5|І станеться, коли засурмить баранячий ріг, коли ви почуєте голос тієї сурми, а ввесь народ крикне гучним криком, то мур цього міста впаде на своєму місці, а народ увійде кожен перед себе.
JOSH|6|6|І покликав Ісус, син Навинів, священиків, та й сказав до них: Несіть ковчега заповіту, а сім священиків будуть нести сім сурем із баранячих рогів перед Господнім ковчегом.
JOSH|6|7|А до народу сказав: Підіть, обійдіть навколо це місто, а озброєний піде перед Господнім ковчегом.
JOSH|6|8|І сталося, як Ісус сказав це народові, то сім священиків, що несли сім сурем із баранячих рогів, ішли та сурмили в ці сурми, а ковчег Господнього заповіту йшов за ними.
JOSH|6|9|А озброєні йшли перед священиками, що сурмили в роги, а військо заднє йшло за ковчегом. І все сурмили в сурми.
JOSH|6|10|А народові Ісус наказав, говорячи: Не будете кричати, і не дасте почути вашого голосу, і не вийде слово з ваших уст аж до дня, коли я скажу вам: Закричіть! І ви закричите.
JOSH|6|11|І Господній ковчег пішов навколо міста, обійшов один раз. І ввійшли до табору, та й ночували в таборі.
JOSH|6|12|І встав Ісус рано вранці, і понесли священики Господнього ковчега.
JOSH|6|13|А сім священиків, що несли сім сурем із баранячих рогів перед Господнім ковчегом, ішли та все сурмили в сурми, а озброєні йшли перед ними, а військо заднє йшло за Господнім ковчегом. І все сурмили в сурми.
JOSH|6|14|І обійшли навколо міста другого дня один раз, та й вернулися до табору. Так зробили шість день.
JOSH|6|15|І сталося сьомого дня, і повставали вони рано вранці, як сходила рання зоря, і обійшли навколо міста за тим приписом сім раз. Тільки того дня обійшли місто навколо сім раз.
JOSH|6|16|І сталося, коли сьомого разу засурмили священики в сурми, то Ісус сказав до народу: Закричіть, бо Господь віддав вам це місто!
JOSH|6|17|І станеться це місто закляттям, воно та все, що в ньому, для Господа. Тільки блудниця Рахав буде жити, вона та всі, хто з нею в домі, бо вона сховала була послів, яких ми посилали.
JOSH|6|18|Та тільки стережіться заклятого, щоб ви самі не стали закляттям, і не взяли з заклятого, і щоб тим не завели Ізраїлевого табору під закляття, і не довели його до нещастя.
JOSH|6|19|А все срібло та золото, і речі мідяні та залізні, це святість для Господа, воно ввійде до Господньої скарбниці.
JOSH|6|20|І закричав народ, і засурмили в сурми. І сталося, як народ почув голос сурми, і закричав народ гучним криком, то впав мур на своєму місці, а народ увійшов до міста, кожен перед себе. І здобули вони те місто.
JOSH|6|21|І зробили вони закляттям усе, що в місті, від чоловіка й аж до жінки, від юнака й аж до старого, і аж до вола, і штуки дрібної худоби, і осла, усе знищили вістрям меча.
JOSH|6|22|А до двох тих людей, що вивідували Край, Ісус сказав: Увійдіть до дому тієї жінки блудниці, і виведіть звідти ту жінку та все, що її, як ви заприсягли були їй.
JOSH|6|23|І ввійшли юнаки, вивідувачі, і вивели Рахав, і батька її, і матір її, і братів її, і все, що її, і всі роди її вивели й умістили поза Ізраїлевим табором.
JOSH|6|24|А місто та все, що в ньому, спалили огнем. Тільки срібло та золото, і речі мідяні та залізні дали до скарбниці Господнього дому.
JOSH|6|25|А блудницю Рахав, і дім її батька, і все, що її, Ісус позоставив при житті. І осіла вона серед Ізраїля, і так є аж до цього дня, бо сховала була послів, яких послав був Ісус вивідати Єрихон.
JOSH|6|26|І того часу заприсягнув Ісус, говорячи: Проклятий перед Господнім лицем кожен, хто встане й відбудує це місто Єрихон, на перворіднім своїм він заложить його, і на наймолодшім своїм поставить брами його.
JOSH|6|27|І був Господь з Ісусом, а слава його розійшлася по всім Краї.
JOSH|7|1|І спроневірилися Ізраїлеві сини в заклятому, Ахан, син Кармія, сина Завдієвого, сина Зерахового, Юдиного племени, узяв із заклятого. І запалився Господній гнів на Ізраїлевих синів.
JOSH|7|2|І послав Ісус мужів з Єрихону в Ай, що при Бет-Евені, на схід від Бет-Елу, і сказав до них, говорячи: Підіть, і вивідайте цей Край. І пішли ті мужі, і вивідали той Ай.
JOSH|7|3|І вернулися вони до Ісуса та й сказали до нього: Нехай не йде ввесь народ, коло двох тисяч люда або коло трьох тисяч люда нехай вийдуть, і поб'ють Ай. Не труди всього народу туди, бо ті вороги нечисленні.
JOSH|7|4|І пішли туди з народу коло трьох тисяч люда, та вони повтікали перед айськими людьми.
JOSH|7|5|І айські люди повибивали з них коло тридцяти й шости чоловіка, та й гнали їх з-перед брами аж до Шеварім, і розбили їх на узбіччі гори. І охляло серце народу, та й стало як вода.
JOSH|7|6|І роздер Ісус одежу свою, та й упав на обличчя своє на землю перед Господнім ковчегом, і лежав аж до вечора він та Ізраїлеві старші, і посипали порохом свою голову.
JOSH|7|7|І сказав Ісус: Ах, Владико Господи, для чого. Ти конче перепровадив цей народ через Йордан, щоб дати нас у руку амореянина, щоб вигубити нас? О, коли б ми були позосталися, і осіли по той бік Йордану!
JOSH|7|8|О, Господи! Що я скажу по тому, як Ізраїль обернув потилицю перед своїми ворогами?
JOSH|7|9|І почують ханаанеянин та всі мешканці цього Краю, і зберуться навколо на нас, і знищать ім'я наше з землі. І що Ти зробиш Своєму великому Йменню?
JOSH|7|10|І сказав Господь до Ісуса: Устань, пощо то ти падаєш на обличчя своє?
JOSH|7|11|Ізраїль згрішив, і вони переступили Мого заповіта, що Я наказав їм, і взяли з заклятого, а також крали, і обманювали, і клали поміж свої речі.
JOSH|7|12|І не зможуть Ізраїлеві сини встояти перед своїми ворогами, вони обернуть спину перед ворогами своїми, бо стали закляттям. Не буду більше з вами, якщо не вигубите заклятого з-поміж себе!
JOSH|7|13|Устань, освяти народ та й скажеш: Освятіться на завтра, бо так сказав Господь, Бог Ізраїлів: Закляте серед тебе, Ізраїлю! Ти не зможеш устояти перед своїми ворогами, аж доки ви не викинете з-поміж себе того заклятого.
JOSH|7|14|І підходьте рано вранці за вашими племенами. І станеться, те плем'я, що його виявить Господь, нехай підходить за родами; а рід, що його виявить Господь, підходитиме за домами, а дім, що його виявить Господь, підходитиме за мужчинами.
JOSH|7|15|І станеться, хто буде виявлений у заклятім, той буде спалений в огні, він та все, що його, бо переступив він заповіта Господнього, і вчинив безсоромне між Ізраїлем.
JOSH|7|16|І встав Ісус рано вранці, і привів Ізраїля за його племенами, і було виявлене Юдине плем'я.
JOSH|7|17|І привів він Юдині роди, і був виявлений рід Зархіїв. І привів він Зархіїв рід за родинами, і був виявлений Завдій.
JOSH|7|18|І привів він його дім за мужчинами, і був виявлений Ахан, син Кармія, сина Завдія, сина Зераха з Юдиного племени.
JOSH|7|19|І сказав Ісус до Ахана: Сину мій, воздай же славу для Господа, Бога Ізраїля, і признайся Йому, і подай мені, що ти зробив? Не скажи неправди передо мною!
JOSH|7|20|І відповів Ахан до Ісуса та й сказав: Дійсно, згрішив я Господеві, Богові Ізраїля, і зробив так та так.
JOSH|7|21|І побачив я в здобичі одного доброго шін'арського плаща, і дві сотні шеклів срібла, і одного золотого зливка, п'ятдесят шеклів вага його, і забажав я їх, і взяв їх. І ось вони сховані в землі в середині намету мого, а срібло під ним.
JOSH|7|22|І послав Ісус посланців, і побігли вони до намету, аж ось сховане воно в наметі, а срібло під ним.
JOSH|7|23|І забрали його з середини намету, і принесли його до Ісуса та до всіх Ізраїлевих синів, і поклали його перед Господнім лицем.
JOSH|7|24|І взяв Ісус Ахана, Зерахового сина, і те срібло, і того плаща, і того золотого зливка, і синів його, і дочок його, і вола його, і осла його, і отару його, і намета його, і все, що його, а ввесь Ізраїль із ним, та й повиводили їх до долини Ахор.
JOSH|7|25|І сказав Ісус: Нащо ти навів нещастя на нас? Нехай на тебе наведе це нещастя Господь цього дня! І вкаменували його, увесь Ізраїль, камінням. І попалили їх в огні, і вкаменували їх камінням.
JOSH|7|26|І поставили над ним велику камінну могилу, що стоїть аж до цього дня. І спинив Господь лютість гніву Свого, тому назвав ім'я того місця: Ахор, аж до цього дня.
JOSH|8|1|І сказав Господь до Ісуса: Не бійся й не лякайся, візьми з собою ввесь військовий люд, та й устань, піди на Ай. Подивися: ось дав Я в руку твою айського царя, і народ його, і місто його, і край його.
JOSH|8|2|І зробиш Аєві, і цареві його, як ти зробив Єрихонові та цареві його, тільки здобич його та худобу його заберете собі. Постав собі засідку на місто позад нього.
JOSH|8|3|І встав Ісус та ввесь військовий люд, щоб іти на Ай. І вибрав Ісус тридцять тисяч чоловіка сильних вояків, та й послав їх уночі.
JOSH|8|4|І він наказав їм, говорячи: Глядіть, чатуйте на Ай з-позад міста, не віддаляйтеся дуже від міста, і будьте всі готові.
JOSH|8|5|А я та ввесь народ, що зо мною, прийдемо до міста. І станеться, коли вийдуть навперейми нам, як перше, то ми втечемо перед ними.
JOSH|8|6|І вийдуть вони за нами, а ми відтягнемо їх від міста, бо скажуть: Вони втікають перед нами, як перше. І ми втечемо перед ними.
JOSH|8|7|А ви встанете з засідки, і здобудете те місто, і Господь, Бог ваш, дасть його вам у вашу руку.
JOSH|8|8|І станеться, як ви візьмете місто, то підпалите місто огнем, зробите за Господнім словом. Глядіть, я вам наказав.
JOSH|8|9|І послав їх Ісус, і пішли вони на засідку, та й засіли між Бет-Елом та між Аєм, із заходу від Аю. А Ісус ночував тієї ночі серед народу.
JOSH|8|10|І встав Ісус рано вранці, і переглянув народ, і пішов він та Ізраїлеві старші перед народом до Аю.
JOSH|8|11|А всі вояки, що були з ним, пішли під гору, і підійшли, і прийшли навпроти того міста, і таборували з півночі Аю, а між ним та між Аєм була долина.
JOSH|8|12|І взяв він коло п'яти тисяч чоловіка, і поставив їх як засідку між Бет-Елом та між Аєм з заходу міста.
JOSH|8|13|І розклав народ, увесь табір, що з півночі міста, а задню частину його з заходу міста. І прийшов Ісус тієї ночі на середину долини.
JOSH|8|14|І сталося, як побачив це айський цар, то люди того міста поспішили, і встали рано, і вийшли навперейми Ізраїля на бій, він та ввесь його народ, на означений час перед степ. А він не знав, що є засідка на нього з-позад міста.
JOSH|8|15|А Ісус та ввесь Ізраїль удавали, ніби побиті перед ними, і втікали дорогою на пустиню.
JOSH|8|16|А ті скликали ввесь народ, що в місті, щоб гнатися за ними. І гналися вони за Ісусом, і віддалилися від міста.
JOSH|8|17|І не полишився ніхто в Аї та в Бет-Елі, хто не погнався б за Ізраїлем. І позоставили вони місто відчиненим, та й гналися за Ізраїлем.
JOSH|8|18|І сказав Господь до Ісуса: Простягни списа, що в руці твоїй, до Аю, бо в руку твою його віддам. І простягнув Ісус списа, що в руці його, до міста.
JOSH|8|19|А засідка швидко встала зо свого місця, та й побігли, як він простягнув свою руку. І ввійшли вони до міста, і здобули його, і поквапилися та й підпалили те місто огнем.
JOSH|8|20|І обернулися айські люди позад себе, та й побачили, аж ось знявся дим міста до неба! І не було в них сили, щоб утікати ані сюди, ані туди... А народ, що втікав до пустині, обернувся на тих, хто гнався за ним.
JOSH|8|21|А Ісус та ввесь Ізраїль, як побачили, що засідка здобула те місто, і що знявся дим із міста, то вернулися, та й повбивали айських людей.
JOSH|8|22|А ті повиходили з міста навперейми них, і опинилися серед Ізраїля: ті з цього боку, а ті з того. І повбивали їх, так що не позосталося з них нікого, хто врятувався б чи втік.
JOSH|8|23|А айського царя вони схопили живого, і привели його до Ісуса.
JOSH|8|24|І сталося, як покінчив Ізраїль забивати всіх айських мешканців на полі, у пустині, що гнали їх по ній, і попадали вони від вістря меча аж до останнього, то вернувся ввесь Ізраїль до Аю, і перебили його вістрям меча.
JOSH|8|25|І було всіх, що впали того дня, від чоловіка й аж до жінки, дванадцять тисяч, усі айські мешканці.
JOSH|8|26|А Ісус не опускав своєї руки, що витягнув зо списом, аж поки не вчинив закляттям усіх айських мешканців.
JOSH|8|27|Тільки худобу та здобич того міста позабирав собі Ізраїль за словом Господа, що наказав був Ісусові.
JOSH|8|28|І спалив Ісус Ай, і поклав його вічною руїною, пусткою, і так є аж до цього дня.
JOSH|8|29|А айського царя повісив на дереві аж до вечірнього часу. А коли сонце заходило, Ісус наказав, і зняли його трупа з того дерева та й кинули його до входу брами міста. І накидали над ним велику камінну могилу, що стоїть аж до цього дня.
JOSH|8|30|Тоді Ісус збудував жертівника для Господа, Бога Ізраїлевого, на горі Евал,
JOSH|8|31|як наказав був Мойсей, раб Господній, Ізраїлевим синам, як написано в книзі Мойсеєвого Закону, жертівника з цілого каміння, що над ними не підіймали заліза. І принесли на ньому цілопалення для Господа, і приносили мирні жертви.
JOSH|8|32|І він написав там на тих каміннях відписа Мойсеєвого Закону, що той написав перед Ізраїлевими синами.
JOSH|8|33|А ввесь Ізраїль, і старші його, і урядники, і судді його, стояли з цього й з того боку ковчегу навпроти священиків-Левитів, що носять ковчега Господнього заповіту, як приходько, так і тубілець, половина його навпроти гори Ґарізім, а половина його навпроти гори Евал, як наказав був Мойсей, раб Господній, благословляти Ізраїлів народ найперше.
JOSH|8|34|А потім він читав усі слова того Закону, благословення та прокляття, усе так, як написано в Законі.
JOSH|8|35|Не було слова зо всього, що наказав був Мойсей, чого не читав би Ісус перед усіма зборами Ізраїля, і жінок, і дітей, і приходька, що ходить серед них.
JOSH|9|1|І сталося, коли це почули всі царі, що по той бік Йордану, на горі та на поділлі, та на всім березі Великого моря навпроти Ливану: хіттеянин, і амореянин, ханаанеянин, періззеянин, хіввеянин і євусеянин,
JOSH|9|2|то вони зібралися разом, щоб однодушно воювати проти Ісуса та проти Ізраїля.
JOSH|9|3|А мешканці Ґів'ону почули, що Ісус зробив Єрихонові та Аєві,
JOSH|9|4|то зробили й вони хитрість. І пішли вони, і забезпечились живністю на дорогу, і взяли повитирані мішки для ослів своїх, і бурдюки для вина повитирані, і потріскані, і пов'язані,
JOSH|9|5|і взуття повитиране та полатане на їхніх ногах, і одежа на них поношена, а ввесь хліб їхньої поживи на дорогу був сухий, запліснілий.
JOSH|9|6|І пішли вони до Ісуса, до табору в Ґілґалі, та й сказали до нього та до мужів Ізраїлевих: Ми прийшли з далекого краю, а ви тепер складіть з нами умову.
JOSH|9|7|І сказали Ізраїлеві мужі до хіввеян: Може ви сидите поблизу нас, то як ми складемо з вами умову?
JOSH|9|8|І сказали вони до Ісуса: Ми твої раби. А Ісус сказав до них: Хто ви та звідки приходите?
JOSH|9|9|І вони сказали йому: З дуже далекого краю прийшли твої раби до Ймення Господа, Бога твого, бо ми чули чутку про Нього, і все, що Він зробив був в Єгипті,
JOSH|9|10|і все, що Він зробив двом аморейським царям, що по той бік Йордану, Сигонові, цареві хешбонському, та Оґові, цареві башанському, що в Аштароті.
JOSH|9|11|І сказали до нас наші старші та всі мешканці нашого краю, говорячи: Візьміть у свою руку поживу на дорогу, і йдіть навпроти них та й скажете їм: Ми ваші раби, а тепер складіть із нами умову.
JOSH|9|12|Оце наш хліб: теплим ми забезпечилися ним у поживу на дорогу з наших домів у день нашого виходу, щоб іти до вас, а тепер ось він висох і став запліснілий.
JOSH|9|13|А ці бурдюки вина, що понаповнювали ми нові, ось подерлися! А ось одежа наша та взуття наше повитиралося від цієї дуже далекої дороги.
JOSH|9|14|І взяли люди з їхньої поживи на дорогу, а Господніх уст не питали.
JOSH|9|15|І вчинив їм Ісус мир, і склав з ними умову, щоб зоставити їх при житті, і присягнули їм начальники громади.
JOSH|9|16|І сталося по трьох днях по тому, як склали з ними умову, то почули, що близькі вони до нього, і сидять вони поміж ними.
JOSH|9|17|І рушили Ізраїлеві сини, і третього дня прибули до їхніх міст. А їхні міста: Ґів'он, і Кефіра, і Беерот, і Кір'ят-Єарім.
JOSH|9|18|І не повбивали їх Ізраїлеві сини, бо начальники громади присягли були їм Господом, Богом Ізраїля. І нарікала вся громада на начальників.
JOSH|9|19|І сказали всі начальники до всієї громади: Ми присягнули їм Господом, Богом Ізраїля, а тепер ми не можемо доторкнутися до них.
JOSH|9|20|Оце зробімо їм, позоставимо їх при житті, і не буде на нас гніву за присягу, що ми присягнули їм.
JOSH|9|21|І сказали до них начальники: Нехай вони живуть. І стали вони рубати дрова та носити воду для всієї громади, як говорили їм начальники.
JOSH|9|22|І покликав їх Ісус, і промовляв до них, говорячи: Чому ви обманили нас, говорячи: Ми дуже далекі від вас, а ви ось сидите серед нас?
JOSH|9|23|А тепер ви прокляті, і не переведеться з-посеред вас раб, і рубачі дров, і носії води для дому Бога мого.
JOSH|9|24|А вони відповіли Ісусові та й сказали: Бо справді виявлено рабам твоїм, що Господь, Бог твій, наказав Мойсеєві, Своєму рабові, дати вам увесь цей Край, і вигубити всіх мешканців цієї землі перед вами. І ми дуже налякалися за своє життя зо страху перед вами, і зробили оцю річ.
JOSH|9|25|А тепер ми оце в руці твоїй: як добре, і як справедливо в очах твоїх учинити нам, учини.
JOSH|9|26|І він зробив їм так, і врятував їх від руки Ізраїлевих синів, і не повбивали їх.
JOSH|9|27|І дав їх Ісус того дня за рубачів дров та за носіїв води для громади й для Господнього жертівника, і так є аж до цього дня, до місця, яке він вибере.
JOSH|10|1|І сталося, як почув єрусалимський цар Адоні-Цедек, що Ісус здобув Ай та вчинив його закляттям, і що як зробив Єрихонові й цареві його, так зробив Аєві та цареві його, і що мешканці Ґів'ону склали мир з Ізраїлем та були серед них,
JOSH|10|2|то дуже налякалися, бо Ґів'он місто велике, як одне з міст царських, і що він більший за Ай, а всі люди його лицарі.
JOSH|10|3|І послав єрусалимський цар Адоні-Цедек до хевронського царя Гогама, і до ярмутського царя Пір'ама, і до лахіського царя Яфії, і до еґлонського царя Девіра, говорячи:
JOSH|10|4|Прийдіть до мене, і допоможіть мені, і ми поб'ємо Ґів'она, бо він замирив з Ісусом та з Ізраїлевими синами.
JOSH|10|5|І вони зібралися, і пішли п'ять аморейських царів: цар єрусалимський, цар хевронський, цар ярмутський, цар лахіський, цар еґлонський, вони та всі табори їхні, і розтаборувалися при Ґів'оні, і воювали проти них.
JOSH|10|6|І послали ґів'онські люди до Ісуса та до табору в Ґілґал, говорячи: Не стримуй своєї руки від своїх рабів! Прийди до нас скоро, і спаси нас та допоможи нам, бо зібралися на нас усі аморейські царі, що замешкують гори.
JOSH|10|7|І рушив Ісус із Ґілґалу, він та з ним усі вояки й військові лицарі.
JOSH|10|8|І сказав Господь до Ісуса: Не бійся їх, бо Я віддав їх у твою руку, ніхто з них не встоїть перед тобою.
JOSH|10|9|І прибув до них Ісус зненацька, цілу ніч ішов із Ґілґалу.
JOSH|10|10|І Господь навів на них замішання перед Ізраїлем, і побив їх великою поразкою в Ґів'оні. І він гнав їх дорогою входу до Бет-Хорону, і бив їх аж до Азеки та аж до Маккеди.
JOSH|10|11|І сталося, коли вони втікали перед Ізраїлем і були на сході від Бет-Хорону, то Господь кидав на них із неба велике каміння аж до Азеки, і вони вмирали. Тих, що повмирали від градового каміння, було більше від тих, що Ізраїлеві сини повбивали мечем.
JOSH|10|12|Тоді Ісус говорив Господеві того дня, коли Господь дав амореянина перед Ізраїлевих синів, та й сказав на очах Ізраїля: Стань, сонце, в Ґів'оні, а ти, місяцю, ув айялонській долині!
JOSH|10|13|І сонце затрималося, а місяць спинився, аж поки народ відімстився своїм ворогам. Чи це не написане в книзі Праведного? І сонце стало на половині неба, і не поспішалося заходити майже цілий день.
JOSH|10|14|І не було такого, як день той, ані перед ним, ані по ньому, щоб Господь так слухав людського голосу, бо Господь воював для Ізраїля.
JOSH|10|15|І вернувся Ісус, а з ним увесь Ізраїль до табору в Ґілґал.
JOSH|10|16|А ті п'ять царів повтікали, та й сховалися в печері в Маккеді.
JOSH|10|17|І було донесено Ісусові й сказано: Знайдені ті п'ять царів, сховані в печері в Маккеді.
JOSH|10|18|А Ісус відказав: Приваліть велике каміння на отвір печери, і призначте до неї людей, щоб їх стерегти.
JOSH|10|19|А ви не стійте, женіться за своїми ворогами, і понищте їхні задні стежі, і не давайте їм входити до їхніх міст, бо Господь, Бог ваш, віддав їх у вашу руку.
JOSH|10|20|І сталося, як завдав їм Ісус та Ізраїлеві сини дуже велику поразку, так, що прийшов їм кінець, а врятовані повтікали від них, і повходили до твердинних міст,
JOSH|10|21|то ввесь народ у спокої вернувся до табору до Ісуса в Маккеді, і ніхто не поворушив язика свого проти кого з Ізраїлевих синів!
JOSH|10|22|І сказав Ісус: Відчиніть отвір печери, і приведіть до мене з печери тих п'ятьох царів.
JOSH|10|23|І вони зробили так, і вивели до нього з печери тих п'ятьох царів: царя єрусалимського, царя хевронського, царя ярмутського, царя лахіського, царя еґлонського.
JOSH|10|24|І сталося, як привели тих царів до Ісуса, то Ісус закликав усіх Ізраїлевих людей, і сказав військовим начальникам, що йшли з ним: Підійдіть, поставте свої ноги на шиї цих царів. І вони попідходили, і поставили свої ноги на їхні шиї.
JOSH|10|25|І сказав до них Ісус: Не бійтеся й не лякайтеся, будьте сильні та відважні, бо Господь зробить так усім вашим ворогам, із якими ви воюєте.
JOSH|10|26|А по цьому Ісус бив їх, і повбивав їх, і повісив їх на п'ятьох деревах. І висіли вони на тих деревах аж до вечора.
JOSH|10|27|І сталося на час заходу сонця, Ісус наказав, і поздіймали їх із дерев, і повкидали їх до печери, де вони були поховалися, і понакладали велике каміння на отвір печери, де воно аж до цього дня.
JOSH|10|28|А Маккеду Ісус здобув того дня, і побив вістрям меча її та царя її, учинив закляттям їх та кожну особу, хто був у ній, не позоставив жодного врятованого в ній. І зробив він її цареві те саме, що зробив був цареві єрихонському.
JOSH|10|29|А Ісус та ввесь Ізраїль із ним перейшов з Маккеди до Лівни, та й воював проти Лівни.
JOSH|10|30|І дав Господь в Ізраїлеву руку також її та царя її, і він побив вістрям меча її та кожну особу, що в ній, не позоставив жодного врятованого в ній. І зробив він цареві її, як зробив був цареві єрихонському.
JOSH|10|31|І перейшов Ісус та ввесь Ізраїль із ним із Лівни до Лахішу, і таборував при ньому та воював проти нього.
JOSH|10|32|І дав Господь в Ізраїлеву руку Лахіш, і здобув він його другого дня, і побив вістрям меча його та кожну особу, що в ньому, усе так, як зробив був Лівні.
JOSH|10|33|Тоді прийшов ґезерський цар Горам допомогти Лахішу, та Ісус побив його й народ його, так що не позоставив жодного в ньому.
JOSH|10|34|І перейшов Ісус та ввесь Ізраїль із ним з Лахішу до Еґлону, і таборували при ньому та воювали з ним.
JOSH|10|35|І здобули його того дня, і побили його вістрям меча, а кожну особу, що в ньому, того дня зробили закляттям, усе так, як зробив був Лахішу.
JOSH|10|36|І пішов Ісус та ввесь Ізраїль із ним з Еґлону до Хеврону, і воював із ним.
JOSH|10|37|І здобув його, і побив вістрям меча його та царя його, і всі міста його, і кожну особу, що в ньому, не позоставив жодного врятованого, усе так, як зробив був Еґлонові. І зробив закляттям його та кожну особу, що в ньому була.
JOSH|10|38|І вернувся Ісус та ввесь Ізраїль із ним до Девіру, і воював із ним.
JOSH|10|39|І він здобув його, і царя його, і всі міста його, і повбивали їх вістрям меча, та й зробив закляттям кожну душу, що в ньому, не позоставив жодного врятованого, як зробив був Хевронові, так зробив Девірові та цареві його, і як зробив був Лівні та цареві її.
JOSH|10|40|І побив Ісус увесь Край: гору, і Неґев і Шефелу, і узбіччя, і всіх їхніх царів, не зоставив жодного врятованого, а кожну особу зробив закляттям, як наказав був Господь, Бог Ізраїлів.
JOSH|10|41|І бив їх Ісус від Кадеш-Барнеа та аж до Аззи, і ввесь ґошенський край, і аж до Ґів'ону.
JOSH|10|42|А всіх тих царів та їхній край Ісус здобув одним разом, бо Господь, Бог Ізраїлів, воював для Ізраїля.
JOSH|10|43|І вернувся Ісус та ввесь Ізраїль із ним до табору в Ґілґал.
JOSH|11|1|І сталося, як почув це хацорський цар Явін, то послав до мадонського царя Йовава, і до царя шімронського, і до царя ахшафського,
JOSH|11|2|і до царів, що з півночі на горі та в степу на південь Кінроту, і в Шефелі, і на верхах Дори з заходу,
JOSH|11|3|ханаанеянин зо сходу та з заходу, а амореянин, і хіттеянин, і періззеянин, і євусеянин, а хіввеянин під Гермоном, у краї Міцпи.
JOSH|11|4|І вийшли вони та всі їхні табори з ними, народ, численний кількістю, як пісок, що на березі моря, і коней та колесниць дуже багато.
JOSH|11|5|І змовилися всі ці царі, і прийшли й таборували разом при озері Мером, щоб воювати з Ізраїлем.
JOSH|11|6|І сказав Господь до Ісуса: Не бійся їх, бо взавтра коло цього часу Я покладу їх усіх трупами перед Ізраїлем; їхнім коням попідрізуєш жили ніг, а їхні колесниці попалиш в огні.
JOSH|11|7|І вийшов на них зненацька Ісус та всі вояки з ним при озері Мером, та й напали на них.
JOSH|11|8|І дав їх Господь в Ізраїлеву руку, і вони повбивали їх, і гнали їх аж до Великого Сидону, і аж до Місрефот-Маїму, і аж до долини Міцпи на схід, і повибивали їх, так що не зоставили їм жодного врятованого.
JOSH|11|9|І зробив їм Ісус, як сказав йому Господь: їхнім коням попідрізував жили, а їхні колесниці попалив ув огні.
JOSH|11|10|І вернувся Ісус того часу, і здобув Хацор, а його царя вбив мечем, бо Хацор перед тим був головою всіх тих царств.
JOSH|11|11|І вони повбивали вістрям меча кожну особу, що в ньому, зробили їх закляттям, не позосталася жодна душа, а Хацора спалив огнем.
JOSH|11|12|А всі царські міста та всіх їхніх царів Ісус здобув, та й повбивав їх вістрям меча, зробив їх закляттям, як наказав був Мойсей, раб Господній.
JOSH|11|13|Тільки всі міста, що стоять на згір'ях своїх, не спалив їх Ізраїль, крім Хацору, одного його спалив Ісус.
JOSH|11|14|А всю здобич тих міст та худобу Ізраїлеві сини забрали собі; тільки кожну людину побили вістрям меча, аж поки вони не вигубили їх, не позоставили жодної душі.
JOSH|11|15|Як Господь наказав був Мойсеєві, Своєму рабові, так Мойсей наказав Ісусові, і так зробив Ісус, не занехав ані слова зо всього, що Господь наказав був Мойсеєві.
JOSH|11|16|І взяв Ісус ввесь той Край: гори Юди і ввесь Неґев, і ввесь ґошенський край, і Шефелу, і Араву, і гори Ізраїлеві, і їхню надморську низину,
JOSH|11|17|від гори Халак, що тягнеться до Сеїру, і аж до Баал-Ґаду в ливанській долині під горою Гермон. А всіх їхніх царів він забрав, і бив їх, і повбивав їх.
JOSH|11|18|Довгий час провадив Ісус війну зо всіма тими царями.
JOSH|11|19|Не було міста, що склало б мир з Ізраїлевими синами, окрім хіввеянина, ґів'онських мешканців, усе взяли війною.
JOSH|11|20|Бо від Господа було, щоб зробити запеклим їхнє серце на війну проти Ізраїля, щоб учинити їх закляттям, щоб не було для них милости, але щоб вигубити їх, як Господь наказав був Мойсеєві.
JOSH|11|21|І прийшов Ісус того часу, і вигубив велетнів із гори, з Хеврону, з Девіру, з Анаву, і з усіх Юдських гір, і з усіх Ізраїлевих гір, разом з їхніми містами Ісус зробив їх закляттям.
JOSH|11|22|Не позоставив велетня в краї Ізраїлевих синів, вони позостали тільки в Аззі, в Ґаті та в Ашдоді.
JOSH|11|23|І взяв Ісус увесь Край, усе так, як говорив був Господь до Мойсея. І Ісус дав його Ізраїлеві на спадок, за їхнім поділом на їхні племена. А Край заспокоївся від війни.
JOSH|12|1|А оце царі того Краю, яких побили Ізраїлеві сини, і посіли їхній Край по тім боці Йордану на схід сонця, від арнонського потоку аж до гори Гермон, та ввесь степ на схід:
JOSH|12|2|Сигон, цар аморейський, що сидів у Хешбоні, що панував від Ароеру, що над берегом арнонського потоку, і середина потоку, і половина Ґілеаду, і аж до потоку Яббоку, границі синів Аммонових,
JOSH|12|3|і степ аж до озера Кінроту на схід, і аж до степового моря, моря Солоного на схід, дорогою на Бет-Гаєшімот, і від Теману під узбіччями Пісґі.
JOSH|12|4|І границя Оґа, царя башанського, із остатку рефаїв, що сидів в Аштароті, і в Едреї,
JOSH|12|5|і що панував на горі Гермон, і на Салха, і на всім Башані аж до границі ґешурейської та маахатейської, і половина Ґілеаду, границя Сигона, царя хешбонського.
JOSH|12|6|Мойсей, раб Господній, та Ізраїлеві сини повбивали їх. І дав його Мойсей раб Господній, на спадок Рувимовому та Ґадовому та половині племени Манасіїного.
JOSH|12|7|А оце царі того Краю, що повбивав Ісус та Ізраїлеві сини по той бік Йордану на захід від Баал-Ґаду в ливанській долині аж до гори Халак, що підіймається до Сеїру, і Ісус віддав її Ізраїлевим племенам на спадок за їхнім поділом,
JOSH|12|8|на горі, і в Шефілі, і в Араві, і на узбіччі, і в пустині, і на півдні, хіттеянина, амореянина, і ханаанеянина, періззеянина, хіввеянина й євусеянина:
JOSH|12|9|цар єрихонський один, цар гайський, що з боку Бет-Елу, один,
JOSH|12|10|цар єрусалимський один, цар хевронський один,
JOSH|12|11|цар ярмутський один, цар лахіський один,
JOSH|12|12|цар єґлонський один, цар ґезерський один,
JOSH|12|13|цар девірський один, цар ґедерський один,
JOSH|12|14|цар хоремський один, цар арадський один,
JOSH|12|15|цар лівенський один, цар адулламський один,
JOSH|12|16|цар маккедський один, цар бет-елський один,
JOSH|12|17|цар таппуахський один, цар хеферський один,
JOSH|12|18|цар афекський один, цар шаронський один,
JOSH|12|19|цар мадонський один, цар хацорський один,
JOSH|12|20|цар шімронський один, цар ахшафський один,
JOSH|12|21|цар таанахський один, цар меґіддівський один,
JOSH|12|22|цар кедеський один, цар йокнеамський при Кармелі один,
JOSH|12|23|цар дорський при Нафат-Дорі один, цар ґоїмський при Ґілґалі один,
JOSH|12|24|цар тірцький один. Усіх царів тридцять і один.
JOSH|13|1|А Ісус постарівся й увійшов у дні. І сказав Господь до нього: Ти постарівся та ввійшов у дні, а Краю позостається ще дуже багато, щоб посісти його.
JOSH|13|2|Оце позосталий Край: усі округи филистимські, і ввесь Ґешурей,
JOSH|13|3|від Шіхору, що навпроти Єгипту, і аж до границі Екрону на північ, що до ханаанеянина залічений, п'ять филистимських князів: аззатський, ашдодський, ашкелонський, ґаттійський і екронський, та аввеї.
JOSH|13|4|Від півдня вся ханаанська земля та Меара, що сидонська, аж до Афеки, аж до аморейської границі,
JOSH|13|5|і ґівлейська земля, і ввесь Ливан на схід сонця від Баал-Ґаду під горою Гермон аж до входу до Хамату.
JOSH|13|6|Усіх мешканців гір від Ливану аж до Місрефот-Маїму, усіх сидонян, Я повиганяю їх перед Ізраїлевими синами. Тільки поділи її жеребком на спадок Ізраїлеві, як Я наказав був тобі.
JOSH|13|7|А тепер поділи цей Край на спадок дев'яти племенам та половині племени Манасіїному.
JOSH|13|8|Разом із ним Рувимові та Ґадові взяли свій спадок що дав їм Мойсей по той бік Йордану на схід, як дав їм Мойсей, раб Господній,
JOSH|13|9|від Ароеру, що на березі арнонського потоку, і місто, що серед тієї долини, і вся медевська рівнина аж до Дівону,
JOSH|13|10|і всі міста Сигона, царя аморейського, що царював у Хешбоні, аж до границі Аммонових синів,
JOSH|13|11|і Ґілеад, і границя ґешурейська та маахейська, і вся гора Гермон, і ввесь Башан аж до Салхи,
JOSH|13|12|усе царство Оґа в Башані, що царював в Аштароті та в Едреї, він позостався з останку рефаїв, а Мойсей повбивав їх та повиганяв їх.
JOSH|13|13|І не вигнали Ізраїлеві сини ґешуреянина, і маахатеянина, і сидів Ґешур та Маахат серед Ізраїля, і так є аж до цього дня.
JOSH|13|14|Тільки Левієвому племені не дав він спадку, огняні жертви Господа, Бога Ізраїля, то спадок його, як Я говорив був йому.
JOSH|13|15|І дав Мойсей племені Рувимових синів спадок за їхніми родами.
JOSH|13|16|І була їм границя від Ароеру, що на березі арнонського потоку, і місто, що серед тієї долини, і вся рівнина при Медеві,
JOSH|13|17|Хешбон і всі міста його, що на рівнині, Дівон, і Бамот-Баал, і Бет-Баал-Меон,
JOSH|13|18|і Ягца, і Кедемот, і Мефаат,
JOSH|13|19|і Кір'ятаїм, і Сівма, і Церет-Гашшахар на горі Емеку,
JOSH|13|20|і Бет-Пеор, і узбіччя Пісґі, і Бет-Гаєшімот,
JOSH|13|21|і всі міста рівнини, і все царство Сигона, царя аморейського, що царював у Хешбоні, що Мойсей убив його та мідіянських начальників: Евія, і Рекема, і Цура, і Хура, і Реву, сигонових князів, мешканців того краю.
JOSH|13|22|А Валаама, Беорового сина, чарівника, Ізраїлеві сини забили мечем серед інших, яких вони побили.
JOSH|13|23|І була границя Рувимових синів: Йордан і границя. Це спадок Рувимових синів за їхніми родами, їхні міста та їхні оселі.
JOSH|13|24|І дав Мойсей Ґадовому племені, синам Ґада за їхніми родами,
JOSH|13|25|і була їм границя: Язер, і всі ґілеадські міста, і половина краю аммонових синів аж до Ароеру, що навпроти Рабби,
JOSH|13|26|А з Хешбону аж до Рамат Гамміцпі й Бетоніму, а від Маханаїму аж до границі Девіру,
JOSH|13|27|і в долині Бет-Гараму, і Бет-Німра, і Суккот, і Цафон, останок царства Сигона, царя хешбонського, Йордан і границя аж до кінця озера Кіннерет по тім боці Йордану на схід.
JOSH|13|28|Це спадок Ґадових синів за їхніми родами, міста та їхні оселі.
JOSH|13|29|І дав Мойсей половині племени Манасіїного, і воно було половині племени Манасіїних синів за їхніми родами.
JOSH|13|30|І була їхня границя від Манахаїму, увесь Башан, усе царство Оґа, царя башанського, і всі села Яіру, що в Башані, шістдесят міст.
JOSH|13|31|А половина Ґілеаду, і Аштарот, і Едрея, міста Оґового царства в Башані, синам Махіра, Манасіїного сина, половині синів Махіра за їхніми родами.
JOSH|13|32|Оце те, що Мойсей дав на спадок в моавських степах по тім боці Йордану на схід.
JOSH|13|33|А Левієвому племені Мойсей не дав спадку, Господь, Бог Ізраїлів, Він їхній спадок, як говорив їм.
JOSH|14|1|А оце те, що посіли Ізраїлеві сини в ханаанському Краї, що дали їм на спадок священик Елеазар, і Ісус, син Навинів, та голови батьків племен Ізраїлевих синів.
JOSH|14|2|Жеребком приділили їхній спадок, як наказав був Господь через Мойсея, дев'яти племенам і половині племени.
JOSH|14|3|Бо дав Мойсей насліддя двох племен, та половини племени по той бік Йордану, а Левитам спадку не дав серед них.
JOSH|14|4|Бо Йосипових синів було двоє поколінь, Манасія та Єфрем, а Левитам не дали спадку в Краю, а тільки міста на оселення та їхні пасовиська для їхньої худоби та для їхнього маєтку.
JOSH|14|5|Як наказав був Господь Мойсеєві, так зробили Ізраїлеві сини, та й поділили Край.
JOSH|14|6|І підійшли Юдині сини до Ісуса в Ґілґалі, та й сказав до нього Калев, син Єфуннеїв, кеназзеянин: Ти знаєш те слово, що Господь говорив до Мойсея, Божого чоловіка, про мене та про тебе в Кадеш-Барнеа.
JOSH|14|7|Я був віку сорока літ, коли Мойсей, раб Господній, посилав мене з Кадеш-Барнеа вивідати той Край. І я доклав йому справу, як було в серці моїм.
JOSH|14|8|А мої браття, що ходили зо мною, знесилили були серце народу, а я обставав за Господом, Богом моїм.
JOSH|14|9|І присягнув Мойсей того дня, говорячи: Поправді кажу, той Край, що нога твоя ходила в ньому, буде на спадок тобі та синам твоїм аж навіки, бо ти обставав за Господом, Богом моїм.
JOSH|14|10|А тепер оце Господь позоставив мене при житті, як говорив. Оце сорок і п'ять літ відтоді, як Господь говорив був це слово Мойсеєві, коли Ізраїль ходив у пустині. А тепер ось я віку восьмидесяти й п'яти літ.
JOSH|14|11|Сьогодні я ще сильний, як того дня, коли Мойсей посилав мене, яка сила моя тоді, така сила моя й тепер, щоб воювати, і виходити, і приходити.
JOSH|14|12|А тепер дай же мені цей гористий край, про який Господь говорив того дня, бо ти чув того дня, що там велетні та великі укріплені міста. Може Господь буде зо мною, і я повиганяю їх, як говорив був Господь.
JOSH|14|13|І поблагословив його Ісус, і дав Калевові, синові Єфуннеєвому, Хеврон за спадок.
JOSH|14|14|Тому став Хеврон Калевові, синові Єфуннеєвому, кеназзеянинові, за спадок, і так є аж до цього дня, за те, що він обставав за Господом, Богом Ізраїля.
JOSH|14|15|А ім'я Хеврону давніше було Кір'ят-Арба, що між велетнів був найбільший чоловік. А Край заспокоївся від війни.
JOSH|15|1|І був жеребок для племени Юдиних синів за їхніми родами: до едомської границі пустиня Цін, на південь від теманського краю.
JOSH|15|2|І була їм південна границя від кінця Солоного моря, від затоки, зверненої на південь.
JOSH|15|3|І йде вона на південь від Маале-Акраббіму, і переходить до Ціну, і підіймається з півдня, від Кадеш-Барнеа й переходить до Хецрону, і підіймається до Аддару й обертається до Кар до Каркаї.
JOSH|15|4|І переходить вона до Адмону, і йде до єгипетського потоку, і границя закінчується на захід. Це буде для вас південна границя.
JOSH|15|5|А границя на схід Солоне море аж до кінця Йордану. А границя у бік півночі: від морської затоки з кінця Йордану,
JOSH|15|6|і підіймається границя до Бет-Хоґли й переходить на північ від Бет-Гаарови; і підіймається та границя до Евен-Боган-Бен-Рувена.
JOSH|15|7|І підіймається та границя від ахорської долини, а на півночі звертається до Ґілґалу, що навпроти Маале-Адумміму, що на південь від потоку. І переходить та границя до Ме-Ен-Шемешу, і закінчується при Ен-Роґелі.
JOSH|15|8|І підіймається та границя до Ґе-Бен-Гінному побіч євусеянина з півдня, це Єрусалим. І підіймається та границя до верхів'я гори, що навпроти Ґе-Гінному на захід, що в кінці Емек-Рефаіму на північ.
JOSH|15|9|І біжить та границя від верхів'я гори до джерела Ме-Нефтоаху, і йде до міст гори Ефрону; і біжить та границя до Баали, це Кір'ят-Єарім.
JOSH|15|10|І обертається та границя з Баали на захід до гори Сеїр, і переходить до плеча гори Єарім з півночі, це Кесалон; і сходить до Бет-Шемешу й переходить до Тімни.
JOSH|15|11|І йде та границя по край Екрону на північ, і біжить та границя до Шіккарону, і переходить до гори Баали, і йде до Явнеїлу. І границя закінчується при заході.
JOSH|15|12|А західня границя до Великого моря. А границя ця границя Юдиних синів навколо за їхніми родами.
JOSH|15|13|А Калеву, синові Єфуннеєвому, він дав частку серед Юдиних синів, за Господнім наказом до Ісуса, Кір'ят-Арби, батька велетнів, воно Хеврон.
JOSH|15|14|І Калев повиганяв звідти трьох велетнів: Шешая, і Ахімана, і Талмая, уроджених велетнів.
JOSH|15|15|І пішов він звідти до девірських мешканців, а ім'я Девіра давніше Кір'ят-Сефер.
JOSH|15|16|І сказав Калев: Хто поб'є Кір'ят-Сефер та здобуде його, то дам йому дочку мою Ахсу за жінку.
JOSH|15|17|І здобув його Отніїл, син Кеназів, брат Калевів. І він дав йому свою дочку Ахсу за жінку.
JOSH|15|18|І сталося, коли вона відходила, то намовила його жадати поля від її батька. І зійшла вона з осла, а Калев сказав їй: Що тобі?
JOSH|15|19|І вона сказала: Дай мені дар благословення! Бо ти дав мені землю суху, то даси мені це й водні джерела. І він дав їй Ґуллот горішній та Ґуллот долішній.
JOSH|15|20|Оце спадок племени Юдиних синів за їхніми родами.
JOSH|15|21|І були ті міста від краю племени Юдиних синів до едомської границі на півдні: Кавцеїл, і Едер, і Яґур,
JOSH|15|22|і Кіна, і Дімона, і Ад'ада,
JOSH|15|23|і Кедеш, і Хацор, і Їтнан,
JOSH|15|24|Зіф, і Телем, і Беалот,
JOSH|15|25|і Хацор-Хадатта, і Керійот-Хецрон, це Хацор,
JOSH|15|26|Амам, і Шема, і Молада,
JOSH|15|27|і Хацор-Ґадда, і Хешмон, і Бет-Пелет,
JOSH|15|28|і Хацар-Шуал, і Беер-Шева, і Бізйотея,
JOSH|15|29|Баала, і Ійїм, і Ецем,
JOSH|15|30|і Елтолад, і Хесіл, і Хорма,
JOSH|15|31|і Ціклаґ, і Мадманна, і Сансанна,
JOSH|15|32|і Леваот, і Шілхім, і Аїн, і Ріммон. Усіх міст двадцять і дев'ять та їхні оселі.
JOSH|15|33|На Шефалі: Ештаол, і Цор'а, і Ашна,
JOSH|15|34|і Заноах, і Ен-Ґаннім, Таппуах і Гаенам,
JOSH|15|35|Ярмут, і Адуллам, Сохо й Азека,
JOSH|15|36|і Шаараїм, і Адітаїм, і Ґедера, і Ґедеротаїм, чотирнадцять міст та їхні оселі.
JOSH|15|37|Ценан, і Хадаша, і Міґдал-Ґад,
JOSH|15|38|і Діл'ан, і Міцпе, і Йоктеїл,
JOSH|15|39|Лахіш, і Боцкат, і Еґлон,
JOSH|15|40|і Каббон, і Лахмас, і Кітліш,
JOSH|15|41|і Ґедерот, Бет-Даґон, і Наама, і Маккеда, шістнадцять міст та їхні оселі.
JOSH|15|42|Лівна, і Етер, і Ашан,
JOSH|15|43|і Ївтах, і Ашна, і Неців,
JOSH|15|44|і Кеіла, і Ахзів, і Мареша, дев'ять міст та їхні оселі.
JOSH|15|45|Екрон і підлеглі міста його та оселі його.
JOSH|15|46|Від Екрону й до моря усе, що при Ашдоді та їхні оселі.
JOSH|15|47|Ашдод, підлеглі міста його та оселі його; Азза, підлеглі міста її та оселі її до єгипетського потоку, і море Велике, і границя.
JOSH|15|48|І на горах: Шамір, і Яттір, і Сохо,
JOSH|15|49|і Данна, і Кір'ят-Санна, він Девір,
JOSH|15|50|і Анав, і Ештемо, і Анім,
JOSH|15|51|і Ґошен, і Холон, і Ґіло, одинадцять міст та їхні оселі.
JOSH|15|52|Арав, і Дума, і Еш'ан,
JOSH|15|53|і Янім, і Бет-Таппуах, і Афека,
JOSH|15|54|і Хумта, і Кір'ят-Арба, це Хеврон, і Ціор, дев'ять міст та їхні оселі.
JOSH|15|55|Маон, Кармел, і Зіф, і Юта,
JOSH|15|56|Їзреїл, і Йокдеам, і Заноах,
JOSH|15|57|Каїн, Ґів'а, і Тімна, десять міст та їхні оселі.
JOSH|15|58|Халхул, Бет-Цур, і Ґедор,
JOSH|15|59|і Маарат, і Бет-Анот, і Елтекон, шість міст та їхні оселі.
JOSH|15|60|Кір'ят-Баал, він Кір'ят-Єарім, і Рабба, двоє міст та їхні оселі.
JOSH|15|61|На пустині: Бет-Гаарава, Міддін, і Сехаха,
JOSH|15|62|і Нівшан, і Ір-Гаммелах, і Ен-Ґеді, шість міст та їхні оселі.
JOSH|15|63|А євусеян, мешканців Єрусалиму, Юдини сини не могли їх вигнати, і осів Євусеянин із Юдиними синами в Єрусалимі, і так є аж до цього дня,
JOSH|16|1|І вийшов жеребок для Йосипових синів: від єрихонського Йордану до єрихонської води на схід пустиня, що тягнеться від Єрихону по горі до Бет-Елу.
JOSH|16|2|І виходить вона з Бет-Елу до Луз, і переходить до границі Арки до Атароту,
JOSH|16|3|і сходить на захід до границі яфлетської, аж до границі Бет-Хорону долішнього, і аж до Ґезеру, і закінчується при морі.
JOSH|16|4|І посіли це Йосипові сини, Манасія та Єфрем.
JOSH|16|5|І була границя Єфремових синів за їхніми родами, а границя їхнього спадку на схід була: Атрот-Аддар аж до горішнього Бет-Хорону.
JOSH|16|6|І виходить та границя до Міхметату з півночі, і повертається границя на схід до Таанат-Шіло, та й переходить його зо сходу до Яноаху.
JOSH|16|7|І сходить вона з Яноаху до Атароту та до Наари, і дотикає Єрихону, і виходить до Йордану.
JOSH|16|8|А з Таппуаху границя йде на захід до потоку Кана, та й закінчується при морі. Це спадок племени Єфремових синів за їхніми родами.
JOSH|16|9|І міста, відділені для Єфремових синів, були серед спадку Манасіїних синів, усі ті міста та їхні оселі.
JOSH|16|10|Та не вигнали вони ханаанеянина, що сидів у Ґезері. І сидів ханаанеянин посеред Єфрема і так є аж до цього дня, і давав данину працею.
JOSH|17|1|І вийшов жеребок для Манасіїного племени, бо він первенець Йосипів, Махірові, Манасіїному первенцеві, Ґілеадовому батькові, бо він був вояк, то був йому Ґілеад та Башан.
JOSH|17|2|І було для позосталих Манасіїних синів за їхніми родами: синам Авіезера, і синам Хелека, і синам Азріїла, і синам Шехема, і синам Хефера, і синам Шеміда. Оце сини Манасії, Йосипового сина, мужі, за їхніми родами.
JOSH|17|3|А в Целофхада, сина Хефера, сина Ґілеада, сина Махіра, сина Манасіїного, не було в нього синів, а тільки дочки. А оце імена його дочок: Махла, і Ноа, і Хоґла, Мілка та Тірца.
JOSH|17|4|І прийшли вони до священика Елеазара, і до Ісуса, Навинового сина, та перед начальників, говорячи: Господь наказав був Мойсеєві дати нам спадок серед наших братів. І дав їм на Господній наказ спадок серед братів їхнього батька.
JOSH|17|5|І випало для Манасії десять наділів, окрім землі Ґілеаду та Башану, що по той бік Йордану,
JOSH|17|6|бо Манасіїні дочки посіли спадок серед синів його, а ґілеадський край був для позосталих Манасіїних синів.
JOSH|17|7|І була Манасіїна границя від Ашер-Гамміхметату, що навпроти Сигему, і йде та границя на південь до мешканців Ен-Таппуаху.
JOSH|17|8|Для Манасії був край Таппуах, а місто Таппуах при Манасіїній границі для Єфремових синів.
JOSH|17|9|І сходить та границя до потоку Кана, на південь від потоку. Ці міста Єфремові серед Манасіїних міст. А границя Манасії від півночі до потоку, а кінчалася при морі.
JOSH|17|10|На південь Єфремове, а на північ Манасіїне, а границею того було море. А в Асирі вони стикалися з півночі, а в Іссахарі зо сходу.
JOSH|17|11|І було для Манасії в Іссахарі та в Асирі: Бет-Шеан та його залежні міста, і Ївлеам та його залежні міста, і мешканці Доару та його залежні міста, і мешканці Таанаху та його залежні міста, і мешканці Меґіддо та його залежні міста, три верховини.
JOSH|17|12|Та Манасіїні сини не могли повиганяти мешканців цих міст, і ханаанеянин продовжував сидіти в тому краї.
JOSH|17|13|І сталося, коли Ізраїлеві сини стали сильні, то дали ханаанеянина на данину, а вигнати не вигнали його.
JOSH|17|14|І говорили Йосипові сини з Ісусом, кажучи: Чому ти дав мені на спадок один жеребок та наділ один, а я ж народ численний, бо до цього часу благословив мене Господь.
JOSH|17|15|І сказав до них Ісус: Якщо ти народ численний, то піди до лісу, та й повикорчовуєш собі там у краї періззеянина та рефаїв, бо Єфремова гора стала тісна для тебе.
JOSH|17|16|І сказали Йосипові сини: Не вистачить нам тієї гори, та й залізна колесниця в кожного ханаанеянина, що сидить у долині, як у того, що в Бет-Шеані та в його залежних містах, так і в того, що в долині Ізреельській.
JOSH|17|17|І сказав Ісус до Йосипового дому, до Єфрема та до Манасії, говорячи: Ти численний народ, і в тебе сила велика, не буде тобі один жеребок,
JOSH|17|18|але буде тобі гористий край; а що там ліс, то викорчуй його, і будуть тобі й його кінці. Бо ти виженеш ханаанеянина, хоч у нього колесниці залізні, хоч він сильний.
JOSH|18|1|І була зібрана вся громада Ізраїлевих синів до Шіло, і вони помістили там скинію заповіту, а перед ними був здобутий Край.
JOSH|18|2|І позоставалося серед Ізраїлевих синів сім племен, що не поділили ще спадку свого.
JOSH|18|3|І сказав Ісус до Ізраїлевих синів: Аж доки ви будете лінуватися піти посісти той Край, що дав вам Господь, Бог ваших батьків?
JOSH|18|4|Дайте від себе по три мужі на плем'я, і я пошлю їх. І вони встануть, і будуть ходити по Краю, і опишуть його за їхнім спадком, та й прийдуть до мене.
JOSH|18|5|І вони поділять його собі на сім частин. Юда стане на своїй границі з півдня, а Йосипів дім стане на своїй границі з півночі.
JOSH|18|6|А ви опишете той Край, сім частин, і принесете описа мені сюди, а я кину вам жеребка тут перед лицем Господа, Бога нашого.
JOSH|18|7|А Левитам нема частки поміж вами, бо священнодіяння Господнє спадщина його. А Ґад, і Рувим, та половина Манасіїного племени взяли свій спадок по той бік Йордану на схід, що дав їм Мойсей, раб Господній.
JOSH|18|8|І встали ті мужі й пішли. А Ісус наказав тим, що пішли описувати Край, говорячи: Ідіть і походіть по Краю, і опишіть його, та й вертайтеся до мене. А я кину вам жеребка тут перед Господнім лицем у Шіло.
JOSH|18|9|І пішли ті мужі, і перейшли по Краю, та й описали його за містами на сім частин у книжці. І прийшли вони до Ісуса до табору в Шіло.
JOSH|18|10|І кинув їм Ісус жеребка в Шіло перед Господнім лицем. І поділив там Ісус Край для Ізраїлевих синів за їхніми поділами.
JOSH|18|11|І вийшов жеребок для племени Веніяминових синів за їхніми родами, і вийшла границя їхнього жеребка між синами Юдиними та між синами Йосиповими.
JOSH|18|12|І була їм границя на північну сторону від Йордану. І підіймається та границя до краю Єрихону з півночі, і підіймається на гору на захід, і закінчується при пустині Бет-Евен.
JOSH|18|13|А звідти переходить та границя до Лузу, до краю Лузу на південь, це Бет-Ел. І сходить та границя до Атрот-Аддару на гору, що з півдня до долішнього Бет-Хорону.
JOSH|18|14|І тягнеться та границя, і повертається на західній бік, на південь від гори, що навпроти Бет-Хорону на південь, і закінчується при Кір'ят-Баалі, це Кір'ят-Єарім, місті Юдиних синів. Це західня сторона.
JOSH|18|15|А південна сторона від кінця Кір'ят-Єаріму. І виходить та границя на захід, і виходить до джерела Ме-Нефтоаху.
JOSH|18|16|І сходить та границя до кінця гори, що навпроти Ґе-Бен-Гіннома, що в долині Рефаїм на північ. І сходить Ґе-Гінном побіч євусеянина на південь, і сходить до Ен-Роґелу,
JOSH|18|17|і тягнеться вона з півночі, і виходить до Ен-Шемешу, і виходить до Ґелілоту, що навпроти Маале-Адуммім. І сходить вона до Евен-Боган-Бен-Реувену.
JOSH|18|18|І переходить побіч навпроти Арави на північ, та й сходить до Арави.
JOSH|18|19|І переходить та границя побіч Бет-Хоґли на північ, і закінчується границя при затоці Солоного моря на північ, до кінця Йордану з півдня. Це границя південна.
JOSH|18|20|А Йордан граничить його зо східньої сторони. Це спадок Веніяминових синів за границями його навколо, за родами його.
JOSH|18|21|І були міста для племени Веніяминових синів за їхніми родами: Єрихон, і Бет-Хоґла, і Емек-Кеціц,
JOSH|18|22|і Бет-Гаарава, і Цемараїм, і Бет-Ел,
JOSH|18|23|і Аввім, і Пара, і Офра,
JOSH|18|24|і Кефар-Гааммоні, і Офні, і Ґева, дванадцять міст та їхні оселі.
JOSH|18|25|Ґів'он, і Рама, і Беерот,
JOSH|18|26|і Міцпе, і Кефіра, і Моца,
JOSH|18|27|і Рекем, і Їрпеїл, і Пар'ала,
JOSH|18|28|і Цела, Елеф, і Євусі, воно Єрусалим, Ґів'ат, Кір'ят-Єарім, чотирнадцять міст та їхні оселі. Це спадок Веніяминових синів за їхніми родами.
JOSH|19|1|А другий жеребок вийшов Симеонові, племені Симеонових синів за їхніми родами. І був їхній спадок серед спадку Юдиних синів.
JOSH|19|2|І був їм у спадку: Беер-Шева, і Молада,
JOSH|19|3|і Хацар-Шуал, і Бала, і Ецем,
JOSH|19|4|і Елтолад, і Бетул, і Хорма,
JOSH|19|5|і Ціклаґ, і Бет-Гаммаркавот, і Хацар-Суса,
JOSH|19|6|і Бет-Леваот, і Шарухен, тринадцять міст та їхні оселі.
JOSH|19|7|Аїн, Ріммон, і Етер, і Ашан, чотири місті та їхні оселі.
JOSH|19|8|А всі оселі, що навколо тих міст аж до Баалат-Беер-Рамат-Неґеву, це спадок племени Симеонових синів за їхніми родами.
JOSH|19|9|З наділу Юдиних синів спадок синів Симеонових, бо наділ Юдиних синів був численніший від них. І посіли Симеонові сини в середині їхнього спадку.
JOSH|19|10|А третій жеребок вийшов Завулоновим синам за їхніми родами, і була границя їхнього спадку аж до Саріду.
JOSH|19|11|І підіймається їхня границя до Яму та Мар'али, і стикається з Даббешетом, і стикається з потоком, що навпроти Йокнеаму,
JOSH|19|12|і вертається з Саріду на схід, до сходу сонця, на границю Кіслот-Фавору, і виходить до Доврату, і підіймається до Яфія.
JOSH|19|13|А звідти переходить на схід, на схід до Ґат-Хеферу, Ет-Каціну, до Ріммон-Гамметоару, до Неї.
JOSH|19|14|І повертається його границя з півночі Ханнатону, і закінчується при Ґе-Їфтах-Елі.
JOSH|19|15|І Каттат, і Нагалал, і Шімрон, і Їд'ала, і Віфлеєм, дванадцять міст та їхні оселі.
JOSH|19|16|Це спадок Завулонових синів за їхніми родами, оці міста та їхні оселі.
JOSH|19|17|Четвертий жеребок вийшов Іссахарові, Іссахаровим синам за їхніми родами.
JOSH|19|18|І була їхня границя: їзреел, і Кесуллот, і Шунем,
JOSH|19|19|і Хафараїм, і Шіон, і Анахарат,
JOSH|19|20|і Раббіт, і Кішйон, Евес,
JOSH|19|21|і Ремет, і Ен-Ґаннім, і Ен-Хадда, і Бет-Паццец.
JOSH|19|22|І дотикається та границя до Фавору, і Шахаціми, і Бет-Шемету, і їхня границя закінчується при Йордані, шістнадцять міст та їхні оселі.
JOSH|19|23|Оце спадок племени Іссахарових синів за їхніми родами, міста та їхні оселі.
JOSH|19|24|А п'ятий жеребок вийшов племені Асирових синів за їхніми родами.
JOSH|19|25|І була їхня границя: Хелкат, і Халі, і Бетен, і Ахшат,
JOSH|19|26|і Алламмелех, і Ам'ад, і Міш'ал, і дотикається Кармелю на захід та Шіхор-Лівнату,
JOSH|19|27|і вертається на схід сонця до Бет-Даґону, і дотикається Завулона та Ґе-Їфтах-Елу, на північ Бет-Гаемеку та Ніелу, і виходить до Кавулу зліва.
JOSH|19|28|І Еврон, і Рехов, і Хаммон, і Кана аж до Сидону Великого.
JOSH|19|29|І вертається та границя до Рами та аж до міста Мівцар-Цору, і вертається границя до Хоси, і закінчується при заході від околиці Ахзіву,
JOSH|19|30|і Умма, і Афек, і Рехов, двадцять і двоє міст та їхні оселі.
JOSH|19|31|Оце спадок племени Асирових синів за їхніми родами, ті міста та їхні оселі.
JOSH|19|32|Синам Нефталимовим вийшов шостий жеребок, для синів Нефталимових за їхніми родами.
JOSH|19|33|І була їхня границя: від Хелефу, від Елону при Цаананнімі, і Адамі Ганнекев, і Явнеїл аж до Лаккуму, і кінчалася вона при Йордані.
JOSH|19|34|І повертається та границя на захід до Ашнот-Фавору, і виходить звідти до Хуккоку та дотикається Завулона з полудня, а Асира дотикається з заходу, а Юди при Йордані на схід сонця.
JOSH|19|35|А міста твердинні: Ціддім, Цер, і Хаммат, Раккат і Кіннерет,
JOSH|19|36|і Адама, і Рама, І Хацор,
JOSH|19|37|і Кедеш, і Едреї, і Ен-Хасор,
JOSH|19|38|і Їр'он, і Міґдал-Ел, Хорем, і Бет-Анат, і Бет-Шамеш, дев'ятнадцять міст та їхні оселі.
JOSH|19|39|Оце спадок племени синів Нефталимових за їхніми родами, міста та їхні оселі.
JOSH|19|40|А племені Данових синів за їхніми родами вийшов сьомий жеребок.
JOSH|19|41|І була границя їхнього насліддя: Цор'а, і Ештаол, і Ір-Шемеш,
JOSH|19|42|і Шаалаббін, і Айялон, і Їтла,
JOSH|19|43|і Елон, і Тімната, і Екрон,
JOSH|19|44|і Елтеке, і Ґіббетон, і Баалат,
JOSH|19|45|і Єгуд, і Бене-Берак, і Ґат-Ріммон,
JOSH|19|46|і Ме-Яркон, і Раккон із границею навпроти Яфи.
JOSH|19|47|І вийшла границя Данових синів від них. А Данові сини пішли й воювали з Лешемом, і здобули його, і побили вістрям меча, і посіли його, та й осілися в ньому. І вони назвали Лешему ім'я: Дан, як ім'я їхнього батька Дана.
JOSH|19|48|Оце спадок племени Данових синів за їхніми родами, ті міста та їхні оселі.
JOSH|19|49|І скінчили вони посідати Край згідно з його границями. І дали Ізраїлеві сини спадок Ісусові, синові Навиновому, посеред себе.
JOSH|19|50|На Господній наказ дали йому те місто, яке він жадав: Тімнат-Серах на Єфремовій горі. І збудував він місто, та й осівся в ньому.
JOSH|19|51|Оце той спадок, що священик Елеазар і Ісус, син Навинів, та голови домів батьків давали племенам Ізраїлевих синів жеребком у Шіло перед Господнім лицем при вході до скинії заповіту. І покінчили вони ділити Край.
JOSH|20|1|І Господь промовляв до Ісуса, говорячи:
JOSH|20|2|Промовляй до Ізраїлевих синів, говорячи: Дайте собі міста на сховища, про які Я говорив вам через Мойсея,
JOSH|20|3|щоб утікав туди убійник, що заб'є кого ненароком невмисне, і вони будуть для вас на місце сховища від месника за кров.
JOSH|20|4|І втече він до одного з тих міст, і стане при вході міської брами, та й буде голосно говорити старшим того міста про свою справу. І вони візьмуть його до міста до себе, і дадуть йому місце, і він осяде з ними.
JOSH|20|5|А коли буде гнатися за ним месник, то не видадуть убійника в руку його, бо він невмисне забив свого ближнього, і не був йому ворогом ані вчора, ані позавчора.
JOSH|20|6|І буде він сидіти в тому місті, аж поки не стане перед громадою на суд, аж до смерти найвищого священика, що буде в тих днях. Тоді повернеться убійник, та й увійде до свого міста та до свого дому, до того міста, звідки він утік.
JOSH|20|7|І посвятили вони Кедеш в Ґалілі на Нефталимовій горі, і Сихем на Єфремовій горі та Кір'ят-Арбу, воно Ефрон, на горі Юдиній.
JOSH|20|8|А по той бік єрихонського Йордану на схід вони дали: Бецер на пустині, на рівнині, із Рувимового племени, і Рамот у Ґілеаді з Ґадового племени, і Ґалан у Башані з Манасіїного племени.
JOSH|20|9|Оце були міста призначення для всіх Ізраїлевих синів та для приходька, що мешкає чужинцем серед них, на сховище туди кожному, хто вб'є кого ненароком. І не помре він від руки месника за кров, аж поки не стане перед громадою.
JOSH|21|1|І підійшли голови домів батьків Левієвих до священика Елеазара й до Ісуса, сина Навинового, та до голів домів батьків племен Ізраїлевих синів,
JOSH|21|2|та й говорили до них у Шіло в ханаанському Краї, кажучи: Господь наказав був через Мойсея дати нам міста на сидіння, а їхні пасовиська для нашої худоби.
JOSH|21|3|І дали Ізраїлеві сини Левитам зо свого наділу на наказ Господній ті міста та їхні пасовиська.
JOSH|21|4|І вийшов жеребок для родів кегатеянина. І були синам священика Аарона з Левитів від племени Юдиного, і від племени Симеонового, і від племени Веніяминового тринадцять міст.
JOSH|21|5|А Кегатовим синам, що позосталися з родів племени Єфремового й з племени Данового та з половини племени Манасіїного жеребком дісталося десять міст.
JOSH|21|6|А для Ґершонових синів від родів Іссахарового племени, і від Асирового племени, і від Нефталимового племени, і від половини Манасіїного племени в Башані жеребком дісталося тринадцять міст.
JOSH|21|7|Мерарієвим синам за їхніми родами дісталося від племени Рувимового, і від племени Ґадового, і від племени Завулонового дванадцять міст.
JOSH|21|8|І дали Ізраїлеві сини Левитам ті міста та їхні пасовиська, як наказав був Господь через Мойсея, жеребком.
JOSH|21|9|І дали вони з племени синів Юдиних та з племени синів Симеонових ті міста, що будуть нижче названі йменням своїм.
JOSH|21|10|І було для Ааронових синів із родів кегатеянина, з Левієвих синів, бо їм був жеребок найперше.
JOSH|21|11|І дали їм місто Кір'ят, батька велетнів Арби, воно Хеврон, на Юдиних горах, та його пасовиська навколо нього.
JOSH|21|12|А мійське поле та оселі його дали Калеву, синові Єфуннеєвому, на власність його.
JOSH|21|13|А синам священика Аарона дали місто сховища вбійника: Хеврон та його пасовиська, і Лівну та її пасовиська,
JOSH|21|14|і Яттір та його пасовиська, і Ештемоа та її пасовиська,
JOSH|21|15|і Холон та його пасовиська, і Девір та його пасовиська,
JOSH|21|16|і Аїн та його пасовиська, і Ютту та її пасовиська, Бет-Шемеш та його пасовиська, дев'ять міст від двох тих племен.
JOSH|21|17|А від Веніяминового племени: Ґів'он та його пасовиська, Ґеву та її пасовиська,
JOSH|21|18|Анатоль та його пасовиська, і Алмон та його пасовиська, міст четверо.
JOSH|21|19|Усіх міст Ааронових синів, священиків, тринадцять міст та їхні пасовиська.
JOSH|21|20|А родам Кегатових синів, Левитам, що позостали від Кегатових синів, міста їхнього жеребка були від Єфремового племени.
JOSH|21|21|І дали їм місто сховища вбійника: Сихем та його пасовиська, на Єфремовій горі, і Ґезер та його пасовиська.
JOSH|21|22|І Ківцаїм та його пасовиська, і Бет-Хорон та його пасовиська, міст четверо.
JOSH|21|23|А від Данового племени: Елтеке та його пасовиська, Ґіббетон та його пасовиська,
JOSH|21|24|Айялон та його пасовиська, Ґат-Ріммон та його пасовиська, міст четверо.
JOSH|21|25|А від половини Манасіїного племени: Таанах та його пасовиська, і Ґат-Ріммон та його пасовиська, міст двоє.
JOSH|21|26|Усіх міст десять та їхні пасовиська для родів позосталих Кегатових синів.
JOSH|21|27|А для Ґершонових синів з Левієвих родів від половини Манасіїного племени місто сховища вбійника: Ґолан у Башані та його пасовиська, і Беештера та її пасовиська, міст двоє.
JOSH|21|28|А від Іссахарового племени: Кіш'йон та його пасовиська, Доврат та його пасовиська,
JOSH|21|29|Ярмут та його пасовиська, Ен-Ґаннім та його пасовиська, міст четверо.
JOSH|21|30|А від Асирового племени: Міш'ал та його пасовиська, Ардон та його пасовиська,
JOSH|21|31|Хелкат та його пасовиська, Рехов та його пасовиська, міст четверо.
JOSH|21|32|А від Нефталимового племени місто сховища вбійника: Кедеш у Ґаліл та його пасовиська, і Хаммот-Дор та його пасовиська, і Картан та його пасовиська, міст троє.
JOSH|21|33|Усіх міст Ґершонових за їхніми родами тринадцять міст та їхні пасовиська.
JOSH|21|34|А для родів Мерарієвих синів, Левитів, позосталих від племени Завулонового: Йокнеам та його пасовиська, Карта та її пасовиська.
JOSH|21|35|Дімна та її пасовиська, Нагалал та його пасовиська, міст четверо.
JOSH|21|36|А від Рувимового племени: Бецар та його пасовиська, і Ягца та її пасовиська,
JOSH|21|37|Кедемот та його пасовиська, і Мефаат та його пасовиська, міст четверо.
JOSH|21|38|А від Ґадового племени місто сховища вбійника: Рамот у Ґілеаді та його пасовиська, і Маханаїм та його пасовиська,
JOSH|21|39|Хешбон та його пасовиська, Язер та його пасовиська, усіх міст четверо.
JOSH|21|40|Усіх міст для Мерарієвих синів за їхніми родами, що позосталися з Левієвих родів, було за їхнім жеребком дванадцять міст.
JOSH|21|41|Усіх Левієвих міст серед власности Ізраїлевих синів сорок і вісім міст та їхні пасовиська.
JOSH|21|42|Будуть ті міста такі: кожне місто з пасовиськом його навколо нього, так для всіх тих міст.
JOSH|21|43|І дав Господь Ізраїлеві ввесь той Край, що присягнув був дати його їхнім батькам, і вони посіли його та й осілися в ньому.
JOSH|21|44|І Господь дав їм мир навколо, усе так, як присягнув був їхнім батькам. І ніхто зо всіх їхніх ворогів на встояв перед ними, усіх їхніх ворогів Господь дав у їхню руку.
JOSH|21|45|Нічого не було невиконаного з усього того доброго слова, що Господь говорив до Ізраїлевого дому, усе збулося.
JOSH|22|1|Тоді покликав Ісус племено Рувимове та Ґадове, та половину Манасіїного племени,
JOSH|22|2|та й сказав їм: Ви виконували все, що вам наказав був раб Господній Мойсей, і ви слухалися голосу мого про все, що я вам наказував.
JOSH|22|3|Ви оце не лишали братів своїх довгі дні аж до цього дня, і ви додержували виконання заповідей Господа, Бога вашого.
JOSH|22|4|А тепер Господь, Бог ваш, дав мир вашим братам, як вам говорив був. І тепер поверніться, та й ідіть собі до наметів своїх, до краю вашої власности, що вам дав Мойсей, раб Господній, на тім боці Йордану.
JOSH|22|5|Тільки дуже пильнуйте виконувати заповідь та Закона, що наказав був вам Мойсей, раб Господній: любити Господа, Бога вашого, і ходити всіма Його дорогами, і додержувати Його заповіді, і линути до Нього, і служити Йому всім вашим серцем та всією вашою душею.
JOSH|22|6|І поблагословив їх Ісус, та й послав їх, а вони пішли до наметів своїх.
JOSH|22|7|А половині Манасіїного племени Мойсей дав у Башані, а половині його дав Ісус з їхніми братами на цім боці Йордану на захід. І також, коли Ісус відпускав їх до їхніх наметів, то поблагословив їх,
JOSH|22|8|та й сказав до них, говорячи: Верніться до своїх наметів із великими маєтками та з дуже численною худобою, зо сріблом, і з золотом, і з міддю, і з залізом, і з дуже багатьома одежами. Поділіть здобич від ваших ворогів із вашими братами.
JOSH|22|9|І вернулися, і пішли сини Рувимові й сини Ґадові та половина Манасіїного племени від Ізраїлевих синів, із Шіло, що в ханаанському Краї, щоб піти до краю Ґілеад, до краю своєї власности, що посіли його на наказ Господній через Мойсея.
JOSH|22|10|І прийшли до йорданських могил, що в ханаанському Краї, і збудували там сини Рувимові й сини Ґадові та половина Манасіїного племени жертівника над Йорданом, жертівника великого на вид.
JOSH|22|11|І почули Ізраїлеві сини таке: Оце збудували сини Рувимові й сини Ґадові та половина Манасіїного племени жертівника навпроти ханаанського Краю, при йорданських могилах, на боці Ізраїлевих синів.
JOSH|22|12|І почули це Ізраїлеві сини, і була зібрана вся громада Ізраїлевих синів до Шіло, щоб піти на них війною.
JOSH|22|13|І послали Ізраїлеві сини до синів Рувимових і до синів Ґадових та до половини Манасіїного племени ґілеадського краю Пінхаса, сина священика Елеазара,
JOSH|22|14|та з ним десять начальників, по одному начальникові для батькового дому з усіх Ізраїлевих племен; а кожен із них голова дому їхніх батьків, вони для тисяч Ізраїлевих.
JOSH|22|15|І прийшли вони до синів Рувимових й до синів Ґадових та до половини Манасіїного племени до ґілеадського краю, та й говорили з ними, кажучи:
JOSH|22|16|Так сказала вся Господня громада: Що це за переступ, що ви спроневірилися ним проти Ізраїлевого Бога, щоб відвернутись сьогодні від Господа? Бо ви збудували собі жертівника, щоб сьогодні збунтуватися проти Господа.
JOSH|22|17|Чи нам мало Пеорового гріха, з якого ми не очистилися аж до цього дня, і була пораза в Господній громаді?
JOSH|22|18|А ви відвертаєтеся сьогодні від Господа. І станеться, ви збунутуєтеся сьогодні проти Господа, а Він узавтра розгнівається на всю Ізраїлеву громаду.
JOSH|22|19|І справді, якщо край вашої посілости нечистий, перейдіть собі до Краю Господньої посілости, що там пробуває Господня скинія, і візьміть посілість серед нас, а на Господа не бунтуйтеся, і не бунтуйтеся проти нас вашим збудуванням собі жертівника, окрім жертівника Господа, Бога нашого.
JOSH|22|20|Чи ж не Ахан, син Зерахів, спроневірився був переступом у заклятому, а гнів був на всю Ізраїлеву громаду? І він був єдиний чоловік, що не помер своєю смертю через свій гріх.
JOSH|22|21|І відповіли сини Рувимові, сини Ґадові та половина Манасіїного племени, і говорили з головами тисяч Ізраїлевих:
JOSH|22|22|Бог богів Господь, Бог богів Господь, Він знає, і Ізраїль він буде знати. Не пощади нас цього дня, якщо бунтом і якщо переступом проти Господа ми це зробили,
JOSH|22|23|якщо ми збудували собі жертівника на відвернення від Господа; а якщо ми будували на принесення цілопалення та жертви хлібної, і якщо на спорядження на ньому мирних жертов, то Господь Він відплатить,
JOSH|22|24|і якщо ми не зробили цього з обавою про таку річ, говорячи: Завтра скажуть ваші сини до наших синів, говорячи: Що вам до Господа, Бога Ізраїлевого?
JOSH|22|25|Бо Господь дав границю поміж нами та поміж вами, сини Рувимові та сини Ґадові, Йордан, нема вам наділу в Господі! І ваші сини відірвуть наших синів від боязні Господа.
JOSH|22|26|Тож сказали ми: Зробім собі, збудуймо жертівника не на цілопалення й не на жертву,
JOSH|22|27|але щоб він був свідком між нами та між вами, і між поколіннями нашими по нас, що ми служили служби Господні перед Його лицем нашими цілопаленнями, і нашими жертвами, і нашими жертвами мирними. І не скажуть ваші сини взавтра до наших синів: нема вам наділу в Господі!
JOSH|22|28|І сказали ми: І станеться, коли так скажуть до нас та до наших поколінь узавтра, то ми скажемо: Подивіться на вигляд жертівника, що зробили були наші батьки не на цілопалення й не на жертву, але щоб був він свідком між нами та між вами.
JOSH|22|29|Борони нас, Боже, бунтуватися нам проти Господа, і відвертатися сьогодні від Господа, щоб будувати жертівника на цілопалення, і на жертву хлібну, і на жертву, окрім жертівника Господа, Бога нашого, що перед скинією Його.
JOSH|22|30|І почув священик Пінхас та начальники громади й голови тисяч Ізраїлевих, що були з ним, ті слова, що казали сини Рувимові й сини Ґадові та сини Манасіїні, і було це добре в їхніх очах.
JOSH|22|31|І сказав Пінхас, син священика Елеазара, до синів Рувимових, і до синів Ґадових та до синів Манасіїних: Сьогодні ми пізнали, що Господь серед вас, що ви не спроневірилися Господеві тим переступом, тепер ви визволили Ізраїлевих синів від Господньої руки.
JOSH|22|32|І вернувся Пінхас, син священика Елеазара, та начальники від синів Рувимових, і від синів Ґадових з ґілеадського краю до Краю ханаанського до Ізраїлевих синів, і здали їм звіт.
JOSH|22|33|І була добра та річ в очах синів Ізраїлевих. І поблагословили Бога Ізраїлеві сини, і не сказали йти на них війною, щоб знищити край, що сини Рувимові та сини Ґадові сидять у ньому.
JOSH|22|34|І назвали сини Рувимові та сини Ґадові ім'я жертівникові: Ед, бо він свідок між нами, що Господь Він Бог.
JOSH|23|1|І сталося по багатьох днях по тому, як Господь дав мир Ізраїлеві від усіх їхніх ворогів навколо, а Ісус постарів, увійшов у літа,
JOSH|23|2|то покликав Ісус усього Ізраїля, його старших, і голів його, і суддів його, і урядників його, та й сказав до них: Я постарів, увійшов у літа.
JOSH|23|3|А ви бачили все, що зробив був Господь, Бог ваш, усім цим людям для вас, бо Господь, Бог ваш, Він Той воюючий для вас!
JOSH|23|4|Дивіться, ось я поділив вам жеребком цих позосталих людей на спадок для ваших племен від Йордану, і всі народи, що вигубив я, аж по море Велике, місце заходу сонця.
JOSH|23|5|А Господь, Бог ваш, Він пожене їх перед вами, і вижене їх перед вами, і ви посядете їхній Край, як говорив був Господь, Бог ваш, до вас.
JOSH|23|6|І ви будете дуже сильні, щоб виконувати й чинити все, написане в книзі Закону Мойсеєвого, щоб не відхилятися від нього ані праворуч, ані ліворуч,
JOSH|23|7|щоб ви не змішувалися з цими людьми, цими позосталими з вами, а ім'я їхніх богів ви не згадаєте, і не будете заприсягати ними, і не будете служити їм, і не будете вклонятися їм,
JOSH|23|8|бо ви будете горнутися тільки до Господа, Бога вашого, як робили ви аж до цього дня.
JOSH|23|9|І вигнав Господь перед вами народи великі та сильні, а ви не встояв ніхто перед вами аж до цього дня.
JOSH|23|10|Один чоловік із вас сам жене тисячу, бо Господь, Бог ваш Він той Вояк для вас, як говорив був Він вам.
JOSH|23|11|І будете ви дуже пильнувати про свої душі, щоб любити Господа, Бога вашого.
JOSH|23|12|Бо якщо справді будете ви відвертатися й приліпитеся до решти цих народів, цих позосталих із вами, і будете свататися з ними, і будете змішуватися з ними, а вони з вами,
JOSH|23|13|то дійсно будете ви знати, що Господь, Бог ваш, більш не гнатиме ці народи перед вами, і вони стануть для вас сіткою й пасткою, та батогом на ваші боки, та терням на ваші очі, аж поки ви не вигинете з-над цієї доброї землі, яку дав вам Господь, Бог ваш.
JOSH|23|14|А я оце сьогодні відходжу дорогою всієї землі. А ви будете знати всім своїм серцем та всією своєю душею, що не відпало ані одне слово зо всіх тих добрих слів, що про вас говорив був Господь, Бог ваш, усе збулося вам, не відпало з нього ані одне слово.
JOSH|23|15|І станеться, отак, як збулося вам усе те добре слово, що про вас говорив був Господь, Бог ваш, так наведе Господь на вас усе те слово зле, аж поки Він вигубить вас з-над цієї доброї землі, яку вам дав Господь, Бог ваш.
JOSH|23|16|Коли ви переступите заповіта Господа, Бога вашого, що Він наказав вам, і підете й будете служити іншим богам, і будете вклонятися їм, то запалиться гнів Господній на вас, і ви скоро погинете з того хорошого Краю, що його Він вам дав.
JOSH|24|1|І зібрав Ісус усі Ізраїлеві племена до Сихему, і покликав Ізраїлевих старших, і голів його, і суддів його, і урядників його, і поставали вони перед Божим лицем.
JOSH|24|2|І сказав Ісус до всього народу: Так сказав Господь, Бог Ізраїлів: По тім боці Річки сиділи були ваші батьки від віків: Терах, батько Авраамів та батько Нахорів, і служили іншим богам.
JOSH|24|3|І взяв Я вашого батька Авраама з того боку Річки, і водив його по всьому ханаанському Краї, і розмножив насіння його, і дав йому Ісака.
JOSH|24|4|І дав Я Ісакові Якова та Ісава, і дав Ісавові гору Сеїр, щоб її посів, а Яків та сини його зійшли до Єгипту.
JOSH|24|5|І послав Я Мойсея та Аарона, та й ударив Єгипет, як зробив Я серед нього, а потому Я вивів вас.
JOSH|24|6|І вивів Я ваших батьків із Єгипту, і ввійшли ви до моря, а Єгипет гнався за вашими батьками колесницями та верхівцями до Червоного моря.
JOSH|24|7|І кликали вони до Господа, і Він поклав темряву між вами та між Єгиптянином, і навів на нього море, і воно покрило його, і ваші очі бачили те, що зробив Я в Єгипті. І сиділи ви в пустині багато днів.
JOSH|24|8|І ввів я вас до краю амореян, що сидять по тім боці Йордану, і вони воювали з вами, а Я дав їх у вашу руку. І ви посіли їхній край, і Я вигубив їх перед вами.
JOSH|24|9|І встав був Балак, син Ціппорів, цар моавський, і воював з Ізраїлем. І він послав і покликав Валаама, Беорового сина, щоб проклясти вас.
JOSH|24|10|Та не хотів Я слухати Валаама, і він, благословляючи, поблагословив вас, і Я врятував вас від його руки.
JOSH|24|11|І перейшли ви Йордан, і прийшли до Єрихону. І воювали з вами господарі Єрихону: періззеянин, і ханаанеянин, і хіттеянин, і ґірґашеянин, і хіввеянин, і євусеянин, а Я дав їх у вашу руку.
JOSH|24|12|І послав Я перед вами шершня, і він вигнав їх перед вами, двох царів аморейських, не мечем твоїм і не луком твоїм.
JOSH|24|13|І дав Я вам Край, що над ним ти не трудився, і міста, що їх ви не будували, і ви осілися в них; виноградники та оливки, яких ви не садили, ви їли.
JOSH|24|14|А тепер бійтеся Господа й служіть Йому в невинності та в правді, і повідкидайте богів, яким служили ваші батьки на тому боці Річки та в Єгипті, та й служіть Господеві.
JOSH|24|15|А якщо зле в очах ваших служити Господеві, виберіть собі сьогодні, кому будете служити, чи богам, яким служили ваші батьки, що по тому боці Річки, та чи богам аморейським, що ви сидите в їхньому краї. А я та дім мій будемо служити Господеві.
JOSH|24|16|І відповів народ та й сказав: Борони, нас Боже, покинути Господа, щоб служити іншим богам!
JOSH|24|17|Бо Господь, Бог наш, Він Той, що вивів нас та наших батьків з єгипетського краю, з дому рабства, і що зробив на наших очах ті великі знамена, і стеріг нас на всій дорозі, що нею ми ходили, і по всіх народах, що ми перейшли серед них.
JOSH|24|18|І повиганяв Господь усі народи та амореянина, мешканця цього Краю, перед нами. І ми будемо служити Господеві, бо Він Бог наш.
JOSH|24|19|І сказав Ісус до народу: Ви не здолієте служити Господеві, бо Він Бог святий, Бог заздрісний Він. Не простить Він вашу провину та ваших гріхів.
JOSH|24|20|Коли ви покинете Господа, і будете служити чужим богам, то Він вернеться, і зробить вам зло, і вигубить вас по тому, як робив був добро вам.
JOSH|24|21|І сказав народ до Ісуса: Ні, таки Господеві будемо служити!
JOSH|24|22|І сказав Ісус до народу: Ви свідки на себе, що ви вибрали Господа служити Йому. І сказали вони: Свідки!
JOSH|24|23|А тепер покиньте чужих богів, що серед вас, і прихиліть своє серце до Господа, Бога Ізраїлевого.
JOSH|24|24|І сказав народ до Ісуса: Господеві, Богові нашому, ми будемо служити, а голосу Його будемо слухатися!
JOSH|24|25|І склав Ісус заповіта з народом того дня, і дав йому постанови та закони в Сихемі.
JOSH|24|26|І написав Ісус ті слова в книзі Божого Закону, і взяв великого каменя, та й поставив його там під тим дубом, що в Господній святині.
JOSH|24|27|І сказав Ісус до всього народу: Ось оцей камінь буде на нас на свідчення, бо він чув усі Господні слова, що Він говорив з нами. І він буде на вас за свідка, щоб ви не виреклися вашого Бога.
JOSH|24|28|І відпустив Ісус народ, кожного до спадку його.
JOSH|24|29|І сталося по тих випадках, і вмер Ісус, син Навинів, раб Господній, віку ста й десяти літ.
JOSH|24|30|І поховали його в границі спадку його, у Тімнат-Серахові, що в Єфремових горах, на північ від гори Ґааш.
JOSH|24|31|І служив Ізраїль Господеві по всі дні Ісуса та по всі дні старших, що продовжили дні свої по Ісусі, і що знали всякий чин Господній, що зробив Він Ізраїлеві.
JOSH|24|32|А Йосипові кості, які Ізраїлеві сини винесли були з Єгипту, поховали в Сихемі, на ділянці поля, що купив був Яків від синів Гамора, Сихемового батька, за сто кеситів.
JOSH|24|33|І Елеазар, син Ааронів, умер, і поховали його на верхів'ї Пінхаса, його сина, яке було йому дане на Єфремовій горі.
