GAL|1|1|Апостол Павло, поставлений ні від людей, ані від чоловіка, але від Ісуса Христа й Бога Отця, що з мертвих Його воскресив,
GAL|1|2|і присутня зо мною вся браття, до Церков галатійських:
GAL|1|3|благодать вам і мир від Бога, Отця нашого, і Господа Ісуса Христа,
GAL|1|4|що за наші гріхи дав Самого Себе, щоб від злого сучасного віку нас визволити, за волею Бога й Отця нашого,
GAL|1|5|Йому слава на віки вічні, амінь!
GAL|1|6|Дивуюся я, що ви так скоро відхилюєтесь від того, хто покликав Христовою благодаттю вас, на іншу Євангелію,
GAL|1|7|що не інша вона, але деякі є, що вас непокоять, і хочуть перевернути Христову Євангелію.
GAL|1|8|Але якби й ми або Ангол із неба зачав благовістити вам не те, що ми вам благовістили, нехай буде проклятий!
GAL|1|9|Як ми перше казали, і тепер знов кажу: коли хто вам не те благовістить, що ви прийняли, нехай буде проклятий!
GAL|1|10|Бо тепер чи я в людей шукаю признання чи в Бога? Чи людям дбаю я догоджати? Бо коли б догоджав я ще людям, я не був би рабом Христовим.
GAL|1|11|Звіщаю ж вам, браття, що Євангелія, яку я благовістив, вона не від людей.
GAL|1|12|Бо я не прийняв, ні навчився її від людини, але відкриттям Ісуса Христа.
GAL|1|13|Чули бо ви про моє поступовання перше в юдействі, що Божу Церкву жорстоко я переслідував та руйнував її.
GAL|1|14|І я перевищував в юдействі багатьох своїх ровесників роду мого, бувши запеклим прихильником моїх отцівських передань.
GAL|1|15|Коли ж Бог, що вибрав мене від утроби матері моєї і покликав благодаттю Своєю, уподобав
GAL|1|16|виявити мною Сина Свого, щоб благовістив я Його між поганами, я не радився зараз із тілом та кров'ю,
GAL|1|17|і не відправився в Єрусалим до апостолів, що передо мною були, а пішов я в Арабію, і знову вернувся в Дамаск.
GAL|1|18|По трьох роках потому пішов я в Єрусалим побачити Кифу, і в нього пробув днів із п'ятнадцять.
GAL|1|19|А іншого з апостолів я не бачив, крім Якова, брата Господнього.
GAL|1|20|А що вам пишу, ось кажу перед Богом, що я не обманюю!
GAL|1|21|Потому пішов я до сирських та кілікійських країн.
GAL|1|22|Церквам же Христовим в Юдеї я знаний не був особисто,
GAL|1|23|тільки чули вони, що той, що колись переслідував їх, благовістить тепер віру, що колись руйнував був її.
GAL|1|24|І славили Бога вони через мене!
GAL|2|1|Потому, по чотирнадцяти роках, я знову ходив в Єрусалим із Варнавою, взявши й Тита з собою.
GAL|2|2|А пішов я за відкриттям. І подав їм Євангелію, що її проповідую між поганами, особливо знатнішим, чи не дарма змагаюся я чи змагався.
GAL|2|3|Але й Тит, що зо мною, бувши греком, не був до обрізання змушений.
GAL|2|4|А щодо прибулих фальшивих братів, що прийшли підглядати нашу вільність, яку маємо в Христі Ісусі, щоб нас поневолити,
GAL|2|5|то ми їх не послухали ані на хвилю, і не піддалися були, щоб тривала в вас правда Євангелії.
GAL|2|6|Щождо тих, що за щось уважають себе, та якими колись вони були, то ні в чому різниці для мене нема, не дивиться Бог на особу людини! Бо ті, що за щось уважають себе, нічого мені не додали,
GAL|2|7|але навпаки, побачивши, що мені припоручена Євангелія для необрізаних, як Петрові для обрізаних,
GAL|2|8|бо Той, хто помагав Петрові в апостольстві між обрізаними, помагав і мені між поганами,
GAL|2|9|і, пізнавши ту благодать, що дана мені, Яків, і Кифа, і Іван, що стовпами вважаються, подали мені та Варнаві правиці спільноти, щоб ми для поган працювали, вони ж для обрізаних,
GAL|2|10|тільки щоб ми пам'ятали про вбогих, що я й пильнував був чинити таке.
GAL|2|11|Коли ж Кифа прийшов був до Антіохії, то відкрито я виступив супроти нього, заслуговував бо він на осуд.
GAL|2|12|Бо він перед тим, як прийшли були дехто від Якова, споживав із поганами. А коли прибули, став ховатися та відлучатися, боячися обрізаних.
GAL|2|13|А з ним лицемірили й інші юдеї, так що навіть Варнава пристав був до їхнього лицемірства.
GAL|2|14|А коли я побачив, що не йдуть вони рівно за євангельською правдою, то перед усіма сказав Кифі: Коли ти, бувши юдеєм, живеш по-поганському, а не по-юдейському, то нащо поган ти примушуєш жити по-юдейському?
GAL|2|15|Ми юдеї природою, а не грішники з поган...
GAL|2|16|А коли ми дізнались, що людина не може бути виправдана ділами Закону, але тільки вірою в Христа Ісуса, то ми ввірували в Христа Ісуса, щоб нам виправдатися вірою в Христа, а не ділами Закону. Бо жадна людина ділами Закону не буде виправдана!
GAL|2|17|Коли ж, шукаючи виправдання в Христі, ми й самі показалися грішниками, то хіба Христос слуга гріху? Зовсім ні!
GAL|2|18|Бо коли я будую знов те, що був зруйнував, то самого себе роблю злочинцем.
GAL|2|19|Бо Законом я вмер для Закону, щоб жити для Бога. Я розп'ятий з Христом.
GAL|2|20|І живу вже не я, а Христос проживає в мені. А що я живу в тілі тепер, живу вірою в Божого Сина, що мене полюбив, і видав за мене Самого Себе.
GAL|2|21|Божої благодаті я не відкидаю. Бо коли набувається правда Законом, то надармо Христос був умер!
GAL|3|1|О, ви нерозумні галати! Хто вас звів не коритися правді, вас, яким перед очима Ісус Христос переднакреслений був, як ніби між вами розп'ятий?
GAL|3|2|Це одне хочу знати від вас: чи ви прийняли Духа ділами Закону, чи із проповіді про віру?
GAL|3|3|Чи ж ви аж такі нерозумні? Духом почавши, кінчите тепер тілом?
GAL|3|4|Чи ви так багато терпіли надармо? Коли б тільки надармо!
GAL|3|5|Отже, Той, Хто вам Духа дає й чуда чинить між вами, чи чинить ділами Закону, чи із проповіді про віру?
GAL|3|6|Так як Авраам був увірував в Бога, і це залічено за праведність йому.
GAL|3|7|Тож знайте, що ті, хто від віри, то сини Авраамові.
GAL|3|8|І Писання, передбачивши, що вірою Бог виправдає поган, благовістило Авраамові: Благословляться в тобі всі народи!
GAL|3|9|Тому ті, хто від віри, будуть поблагословлені з вірним Авраамом.
GAL|3|10|А всі ті, хто на діла Закону покладається, вони під прокляттям. Бо написано: Проклятий усякий, хто не триває в усьому, що написано в книзі Закону, щоб чинити оте!
GAL|3|11|А що перед Богом Законом ніхто не виправдується, то це ясно, бо праведний житиме вірою.
GAL|3|12|А Закон не від віри, але хто чинитиме те, той житиме ним.
GAL|3|13|Христос відкупив нас від прокляття Закону, ставши прокляттям за нас, бо написано: Проклятий усякий, хто висить на дереві,
GAL|3|14|щоб Авраамове благословення в Ісусі Христі поширилося на поган, щоб обітницю Духа прийняти нам вірою.
GAL|3|15|Браття, кажу я по-людському: навіть людського затвердженого заповіту ніхто не відкидає та до нього не додає.
GAL|3|16|А обітниці дані були Авраамові й насінню його. Не говориться: і насінням, як про багатьох, але як про одного: і Насінню твоєму, яке є Христос.
GAL|3|17|А я кажу це, що заповіту, від Бога затвердженого, Закон, що прийшов по чотириста тридцяти роках, не відкидає, щоб обітницю він зруйнував.
GAL|3|18|Бо коли від Закону спадщина, то вже не з обітниці; Авраамові ж Бог дарував із обітниці.
GAL|3|19|Що ж Закон? Він був даний з причини переступів, аж поки прийде Насіння, якому обітниця дана була; він учинений був Анголами рукою посередника.
GAL|3|20|Але посередник не є для одного, Бог же один.
GAL|3|21|Отож, чи ж Закон проти Божих обітниць? Зовсім ні! Якби бо був даний Закон, щоб він міг оживляти, то праведність справді була б від Закону!
GAL|3|22|Та все зачинило Писання під гріх, щоб віруючим була дана обітниця з віри в Ісуса Христа.
GAL|3|23|Але поки прийшла віра, під Законом стережено нас, замкнених до приходу віри, що мала об'явитись.
GAL|3|24|Тому то Закон виховником був до Христа, щоб нам виправдатися вірою.
GAL|3|25|А як віра прийшла, то вже ми не під виховником.
GAL|3|26|Бо ви всі сини Божі через віру в Христа Ісуса!
GAL|3|27|Бо ви всі, що в Христа охристилися, у Христа зодягнулися!
GAL|3|28|Нема юдея, ні грека, нема раба, ані вільного, нема чоловічої статі, ані жіночої, бо всі ви один у Христі Ісусі!
GAL|3|29|А коли ви Христові, то ви Авраамове насіння й за обітницею спадкоємці.
GAL|4|1|Тож кажу я: поки спадкоємець дитина, він нічим від раба не різниться, хоч він пан над усім,
GAL|4|2|але під опікунами та керівниками знаходиться він аж до часу, що визначив батько.
GAL|4|3|Так і ми, поки дітьми були, то були поневолені стихіями світу.
GAL|4|4|Як настало ж виповнення часу, Бог послав Свого Сина, що родився від жони, та став під Законом,
GAL|4|5|щоб викупити підзаконних, щоб усиновлення ми прийняли.
GAL|4|6|А що ви сини, Бог послав у ваші серця Духа Сина Свого, що викликує: Авва, Отче!
GAL|4|7|Тому ти вже не раб, але син. А як син, то й спадкоємець Божий через Христа.
GAL|4|8|Та тоді, не знаючи Бога, служили ви тим, що з істоти богами вони не були.
GAL|4|9|А тепер, як пізнали ви Бога, чи краще як Бог вас пізнав, як вертаєтесь знов до слабих та вбогих стихій, яким хочете знов, як давніше, служити?
GAL|4|10|Ви вважаєте пильно на дні та на місяці, і на пори та роки.
GAL|4|11|Я боюся за вас, чи не дармо я працював коло вас?...
GAL|4|12|Прошу я вас, браття, будьте, як я, бо й я такий самий, як ви. Нічим ви мене не покривдили!
GAL|4|13|І знаєте ви, що в немочі тіла я перше звіщав вам Євангелію,
GAL|4|14|ви ж моєю спокусою в тілі моїм не погордували, і мене не відкинули, але, немов Ангола Божого, ви прийняли мене, як Христа Ісуса!
GAL|4|15|Тож де ваше тодішнє блаженство? Свідкую бо вам, що якби було можна, то ви вибрали б очі свої та мені віддали б!
GAL|4|16|Чи ж я став для вас ворогом, правду говорячи вам?
GAL|4|17|Недобре пильнують про вас, але вас відлучити хочуть, щоб ви пильнували про них.
GAL|4|18|То добре, пильнувати про добре постійно, а не тільки тоді, як приходжу до вас.
GAL|4|19|Дітки мої, я знову для вас терплю муки породу, поки образ Христа не відіб'ється в вас!
GAL|4|20|Я хотів би тепер бути в вас та змінити свій голос, бо маю я сумнів за вас.
GAL|4|21|Скажіть мені ви, що хочете бути під Законом: чи не слухаєтесь ви Закону?
GAL|4|22|Бо написано: Мав Авраам двох синів, одного від рабині, а другого від вільної.
GAL|4|23|Але той, хто був від рабині, народився за тілом, а хто був від вільної, за обітницею.
GAL|4|24|Розуміти це треба інакше, бо це два заповіти: один від гори Сінай, що в рабство народжує, а він то Аґар.
GAL|4|25|Бо Аґар то гора Сінай в Арабії, а відповідає сучасному Єрусалимові, який у рабстві з своїми дітьми.
GAL|4|26|А вишній Єрусалим вільний, він мати всім нам!
GAL|4|27|Бо написано: Звеселися, неплідна, ти, що не родиш! Гукай та викликуй ти, що в породі не мучилась, бо в полишеної значно більше дітей, ніж у тієї, що має вона чоловіка!
GAL|4|28|А ви, браття, діти обітниці за Ісаком!
GAL|4|29|Але як і тоді, хто родився за тілом, переслідував тих, хто родився за духом, так само й тепер.
GAL|4|30|Та що каже Писання? Прожени рабиню й сина її, бо не буде спадкувати син рабині разом із сином вільної.
GAL|4|31|Тому, браття, не сини ми рабині, але вільної!
GAL|5|1|Христос для волі нас визволив. Тож стійте в ній та не піддавайтеся знову в ярмо рабства!
GAL|5|2|Ось я, Павло, кажу вам, що коли ви обрізуєтесь, то нема вам тоді жадної користи від Христа.
GAL|5|3|І свідкую я знову всякому чоловікові, який обрізується, що повинен він виконати ввесь Закон.
GAL|5|4|Ви, що Законом виправдуєтесь, полишилися без Христа, відпали від благодаті!
GAL|5|5|Бо ми в дусі з віри чекаємо надії праведности.
GAL|5|6|Бо сили не має в Христі Ісусі ані обрізання, ані необрізання, але віра, що чинна любов'ю.
GAL|5|7|Бігли ви добре. Хто заборонив вам коритися правді?
GAL|5|8|Таке переконання не від Того, Хто вас покликав.
GAL|5|9|Трохи розчини квасить усе тісто!
GAL|5|10|Я в Господі маю надію на вас, що нічого іншого думати не будете ви. А хто вас непокоїть, осуджений буде, хоч би він хто був!
GAL|5|11|Чого ж, браття, мене ще переслідують, коли я обрізання ще проповідую? Тоді спокуса хреста в ніщо обертається!
GAL|5|12|О, коли б були навіть відсічені ті, хто підбурює вас!
GAL|5|13|Бо ви, браття, на волю покликані, але щоб ваша воля не стала приводом догоджати тілу, а любов'ю служити один одному!
GAL|5|14|Бо ввесь Закон в однім слові міститься: Люби свого ближнього, як самого себе!
GAL|5|15|Коли ж ви гризете та їсте один одного, то глядіть, щоб не знищили ви один одного!
GAL|5|16|І кажу: ходіть за духом, і не вчините пожадливости тіла,
GAL|5|17|бо тіло бажає противного духові, а дух противного тілу, і супротивні вони один одному, щоб ви чинили не те, чого хочете.
GAL|5|18|Коли ж дух вас провадить, то ви не під Законом.
GAL|5|19|Учинки тіла явні, то є: перелюб, нечистість, розпуста,
GAL|5|20|ідолослуження, чари, ворожнечі, сварка, заздрість, гнів, суперечки, незгоди, єресі,
GAL|5|21|завидки, п'янство, гулянки й подібне до цього. Я про це попереджую вас, як і попереджав був, що хто чинить таке, не вспадкують вони Царства Божого!
GAL|5|22|А плід духа: любов, радість, мир, довготерпіння, добрість, милосердя, віра,
GAL|5|23|лагідність, здержливість: Закону нема на таких!
GAL|5|24|А ті, що Христові Ісусові, розп'яли вони тіло з пожадливостями та з похотями.
GAL|5|25|Коли духом живемо, то й духом ходімо!
GAL|5|26|Не будьмо чванливі, не дражнімо один одного, не завидуймо один одному!
GAL|6|1|Браття, як людина й упаде в який прогріх, то ви, духовні, виправляйте такого духом лагідности, сам себе доглядаючи, щоб не спокусився й ти!
GAL|6|2|Носіть тягарі один одного, і так виконаєте закона Христового.
GAL|6|3|Коли бо хто думає, що він щось, бувши ніщо, сам себе той обманює.
GAL|6|4|Нехай кожен досліджує діло своє, і тоді матиме тільки в собі похвалу, а не в іншому!
GAL|6|5|Бо кожен нестиме свій власний тягар!
GAL|6|6|А хто слова навчається, нехай ділиться всяким добром із навчаючим.
GAL|6|7|Не обманюйтеся, Бог осміяний бути не може. Бо що тільки людина посіє, те саме й пожне!
GAL|6|8|Бо хто сіє для власного тіла свого, той від тіла тління пожне. А хто сіє для духа, той від духа пожне життя вічне.
GAL|6|9|А роблячи добре, не знуджуймося, бо часу свого пожнемо, коли не ослабнемо.
GAL|6|10|Тож тому, поки маємо час, усім робімо добро, а найбільш одновірним!
GAL|6|11|Погляньте, якими великими буквами я написав вам своєю рукою!
GAL|6|12|Усі ті, хто бажає хвалитися тілом, змушують вас обрізуватись, щоб тільки вони не були переслідувані за хреста Христового.
GAL|6|13|Бо навіть і ті, хто обрізується, самі не зберігають Закона, а хочуть, щоб ви обрізувались, щоб хвалитися їм вашим тілом.
GAL|6|14|А щодо мене, то нехай нічим не хвалюся, хіба тільки хрестом Господа нашого Ісуса Христа, що ним розп'ятий світ для мене, а я для світу.
GAL|6|15|Бо сили немає ані обрізання, ані необрізання, а створіння нове.
GAL|6|16|А всі ті, хто піде за цим правилом, мир та милість на них, і на Ізраїля Божого!
GAL|6|17|Зрештою, хай ніхто не турбує мене, бо ношу я Ісусові рани на тілі своїм!...
GAL|6|18|Благодать Господа нашого Ісуса Христа нехай буде з духом вашим, браття! Амінь.
