MATT|1|1|A record of the genealogy of Jesus Christ the son of David, the son of Abraham:
MATT|1|2|Abraham was the father of Isaac, Isaac the father of Jacob, Jacob the father of Judah and his brothers,
MATT|1|3|Judah the father of Perez and Zerah, whose mother was Tamar, Perez the father of Hezron, Hezron the father of Ram,
MATT|1|4|Ram the father of Amminadab, Amminadab the father of Nahshon, Nahshon the father of Salmon,
MATT|1|5|Salmon the father of Boaz, whose mother was Rahab, Boaz the father of Obed, whose mother was Ruth, Obed the father of Jesse,
MATT|1|6|and Jesse the father of King David. David was the father of Solomon, whose mother had been Uriah's wife,
MATT|1|7|Solomon the father of Rehoboam, Rehoboam the father of Abijah, Abijah the father of Asa,
MATT|1|8|Asa the father of Jehoshaphat, Jehoshaphat the father of Jehoram, Jehoram the father of Uzziah,
MATT|1|9|Uzziah the father of Jotham, Jotham the father of Ahaz, Ahaz the father of Hezekiah,
MATT|1|10|Hezekiah the father of Manasseh, Manasseh the father of Amon, Amon the father of Josiah,
MATT|1|11|and Josiah the father of Jeconiah and his brothers at the time of the exile to Babylon.
MATT|1|12|After the exile to Babylon: Jeconiah was the father of Shealtiel, Shealtiel the father of Zerubbabel,
MATT|1|13|Zerubbabel the father of Abiud, Abiud the father of Eliakim, Eliakim the father of Azor,
MATT|1|14|Azor the father of Zadok, Zadok the father of Akim, Akim the father of Eliud,
MATT|1|15|Eliud the father of Eleazar, Eleazar the father of Matthan, Matthan the father of Jacob,
MATT|1|16|and Jacob the father of Joseph, the husband of Mary, of whom was born Jesus, who is called Christ.
MATT|1|17|Thus there were fourteen generations in all from Abraham to David, fourteen from David to the exile to Babylon, and fourteen from the exile to the Christ.
MATT|1|18|This is how the birth of Jesus Christ came about: His mother Mary was pledged to be married to Joseph, but before they came together, she was found to be with child through the Holy Spirit.
MATT|1|19|Because Joseph her husband was a righteous man and did not want to expose her to public disgrace, he had in mind to divorce her quietly.
MATT|1|20|But after he had considered this, an angel of the Lord appeared to him in a dream and said, "Joseph son of David, do not be afraid to take Mary home as your wife, because what is conceived in her is from the Holy Spirit.
MATT|1|21|She will give birth to a son, and you are to give him the name Jesus, because he will save his people from their sins."
MATT|1|22|All this took place to fulfill what the Lord had said through the prophet:
MATT|1|23|"The virgin will be with child and will give birth to a son, and they will call him Immanuel"--which means, "God with us."
MATT|1|24|When Joseph woke up, he did what the angel of the Lord had commanded him and took Mary home as his wife.
MATT|1|25|But he had no union with her until she gave birth to a son. And he gave him the name Jesus.
MATT|2|1|After Jesus was born in Bethlehem in Judea, during the time of King Herod, Magi from the east came to Jerusalem
MATT|2|2|and asked, "Where is the one who has been born king of the Jews? We saw his star in the east and have come to worship him."
MATT|2|3|When King Herod heard this he was disturbed, and all Jerusalem with him.
MATT|2|4|When he had called together all the people's chief priests and teachers of the law, he asked them where the Christ was to be born.
MATT|2|5|"In Bethlehem in Judea," they replied, "for this is what the prophet has written:
MATT|2|6|"'But you, Bethlehem, in the land of Judah, are by no means least among the rulers of Judah; for out of you will come a ruler who will be the shepherd of my people Israel.'"
MATT|2|7|Then Herod called the Magi secretly and found out from them the exact time the star had appeared.
MATT|2|8|He sent them to Bethlehem and said, "Go and make a careful search for the child. As soon as you find him, report to me, so that I too may go and worship him."
MATT|2|9|After they had heard the king, they went on their way, and the star they had seen in the east went ahead of them until it stopped over the place where the child was.
MATT|2|10|When they saw the star, they were overjoyed.
MATT|2|11|On coming to the house, they saw the child with his mother Mary, and they bowed down and worshiped him. Then they opened their treasures and presented him with gifts of gold and of incense and of myrrh.
MATT|2|12|And having been warned in a dream not to go back to Herod, they returned to their country by another route.
MATT|2|13|When they had gone, an angel of the Lord appeared to Joseph in a dream. "Get up," he said, "take the child and his mother and escape to Egypt. Stay there until I tell you, for Herod is going to search for the child to kill him."
MATT|2|14|So he got up, took the child and his mother during the night and left for Egypt,
MATT|2|15|where he stayed until the death of Herod. And so was fulfilled what the Lord had said through the prophet: "Out of Egypt I called my son."
MATT|2|16|When Herod realized that he had been outwitted by the Magi, he was furious, and he gave orders to kill all the boys in Bethlehem and its vicinity who were two years old and under, in accordance with the time he had learned from the Magi.
MATT|2|17|Then what was said through the prophet Jeremiah was fulfilled:
MATT|2|18|"A voice is heard in Ramah, weeping and great mourning, Rachel weeping for her children and refusing to be comforted, because they are no more."
MATT|2|19|After Herod died, an angel of the Lord appeared in a dream to Joseph in Egypt
MATT|2|20|and said, "Get up, take the child and his mother and go to the land of Israel, for those who were trying to take the child's life are dead."
MATT|2|21|So he got up, took the child and his mother and went to the land of Israel.
MATT|2|22|But when he heard that Archelaus was reigning in Judea in place of his father Herod, he was afraid to go there. Having been warned in a dream, he withdrew to the district of Galilee,
MATT|2|23|and he went and lived in a town called Nazareth. So was fulfilled what was said through the prophets: "He will be called a Nazarene."
MATT|3|1|In those days John the Baptist came, preaching in the Desert of Judea
MATT|3|2|and saying, "Repent, for the kingdom of heaven is near."
MATT|3|3|This is he who was spoken of through the prophet Isaiah: "A voice of one calling in the desert, 'Prepare the way for the Lord, make straight paths for him.'"
MATT|3|4|John's clothes were made of camel's hair, and he had a leather belt around his waist. His food was locusts and wild honey.
MATT|3|5|People went out to him from Jerusalem and all Judea and the whole region of the Jordan.
MATT|3|6|Confessing their sins, they were baptized by him in the Jordan River.
MATT|3|7|But when he saw many of the Pharisees and Sadducees coming to where he was baptizing, he said to them: "You brood of vipers! Who warned you to flee from the coming wrath?
MATT|3|8|Produce fruit in keeping with repentance.
MATT|3|9|And do not think you can say to yourselves, 'We have Abraham as our father.' I tell you that out of these stones God can raise up children for Abraham.
MATT|3|10|The ax is already at the root of the trees, and every tree that does not produce good fruit will be cut down and thrown into the fire.
MATT|3|11|"I baptize you with water for repentance. But after me will come one who is more powerful than I, whose sandals I am not fit to carry. He will baptize you with the Holy Spirit and with fire.
MATT|3|12|His winnowing fork is in his hand, and he will clear his threshing floor, gathering his wheat into the barn and burning up the chaff with unquenchable fire."
MATT|3|13|Then Jesus came from Galilee to the Jordan to be baptized by John.
MATT|3|14|But John tried to deter him, saying, "I need to be baptized by you, and do you come to me?"
MATT|3|15|Jesus replied, "Let it be so now; it is proper for us to do this to fulfill all righteousness." Then John consented.
MATT|3|16|As soon as Jesus was baptized, he went up out of the water. At that moment heaven was opened, and he saw the Spirit of God descending like a dove and lighting on him.
MATT|3|17|And a voice from heaven said, "This is my Son, whom I love; with him I am well pleased."
MATT|4|1|Then Jesus was led by the Spirit into the desert to be tempted by the devil.
MATT|4|2|After fasting forty days and forty nights, he was hungry.
MATT|4|3|The tempter came to him and said, "If you are the Son of God, tell these stones to become bread."
MATT|4|4|Jesus answered, "It is written: 'Man does not live on bread alone, but on every word that comes from the mouth of God.'"
MATT|4|5|Then the devil took him to the holy city and had him stand on the highest point of the temple.
MATT|4|6|"If you are the Son of God," he said, "throw yourself down. For it is written: "'He will command his angels concerning you, and they will lift you up in their hands, so that you will not strike your foot against a stone.'"
MATT|4|7|Jesus answered him, "It is also written: 'Do not put the Lord your God to the test.'"
MATT|4|8|Again, the devil took him to a very high mountain and showed him all the kingdoms of the world and their splendor.
MATT|4|9|"All this I will give you," he said, "if you will bow down and worship me."
MATT|4|10|Jesus said to him, "Away from me, Satan! For it is written: 'Worship the Lord your God, and serve him only.'"
MATT|4|11|Then the devil left him, and angels came and attended him.
MATT|4|12|When Jesus heard that John had been put in prison, he returned to Galilee.
MATT|4|13|Leaving Nazareth, he went and lived in Capernaum, which was by the lake in the area of Zebulun and Naphtali--
MATT|4|14|to fulfill what was said through the prophet Isaiah:
MATT|4|15|"Land of Zebulun and land of Naphtali, the way to the sea, along the Jordan, Galilee of the Gentiles--
MATT|4|16|the people living in darkness have seen a great light; on those living in the land of the shadow of death a light has dawned."
MATT|4|17|From that time on Jesus began to preach, "Repent, for the kingdom of heaven is near."
MATT|4|18|As Jesus was walking beside the Sea of Galilee, he saw two brothers, Simon called Peter and his brother Andrew. They were casting a net into the lake, for they were fishermen.
MATT|4|19|"Come, follow me," Jesus said, "and I will make you fishers of men."
MATT|4|20|At once they left their nets and followed him.
MATT|4|21|Going on from there, he saw two other brothers, James son of Zebedee and his brother John. They were in a boat with their father Zebedee, preparing their nets. Jesus called them,
MATT|4|22|and immediately they left the boat and their father and followed him.
MATT|4|23|Jesus went throughout Galilee, teaching in their synagogues, preaching the good news of the kingdom, and healing every disease and sickness among the people.
MATT|4|24|News about him spread all over Syria, and people brought to him all who were ill with various diseases, those suffering severe pain, the demon-possessed, those having seizures, and the paralyzed, and he healed them.
MATT|4|25|Large crowds from Galilee, the Decapolis, Jerusalem, Judea and the region across the Jordan followed him.
MATT|5|1|Now when he saw the crowds, he went up on a mountainside and sat down. His disciples came to him,
MATT|5|2|and he began to teach them saying:
MATT|5|3|"Blessed are the poor in spirit, for theirs is the kingdom of heaven.
MATT|5|4|Blessed are those who mourn, for they will be comforted.
MATT|5|5|Blessed are the meek, for they will inherit the earth.
MATT|5|6|Blessed are those who hunger and thirst for righteousness, for they will be filled.
MATT|5|7|Blessed are the merciful, for they will be shown mercy.
MATT|5|8|Blessed are the pure in heart, for they will see God.
MATT|5|9|Blessed are the peacemakers, for they will be called sons of God.
MATT|5|10|Blessed are those who are persecuted because of righteousness, for theirs is the kingdom of heaven.
MATT|5|11|"Blessed are you when people insult you, persecute you and falsely say all kinds of evil against you because of me.
MATT|5|12|Rejoice and be glad, because great is your reward in heaven, for in the same way they persecuted the prophets who were before you.
MATT|5|13|"You are the salt of the earth. But if the salt loses its saltiness, how can it be made salty again? It is no longer good for anything, except to be thrown out and trampled by men.
MATT|5|14|"You are the light of the world. A city on a hill cannot be hidden.
MATT|5|15|Neither do people light a lamp and put it under a bowl. Instead they put it on its stand, and it gives light to everyone in the house.
MATT|5|16|In the same way, let your light shine before men, that they may see your good deeds and praise your Father in heaven.
MATT|5|17|"Do not think that I have come to abolish the Law or the Prophets; I have not come to abolish them but to fulfill them.
MATT|5|18|I tell you the truth, until heaven and earth disappear, not the smallest letter, not the least stroke of a pen, will by any means disappear from the Law until everything is accomplished.
MATT|5|19|Anyone who breaks one of the least of these commandments and teaches others to do the same will be called least in the kingdom of heaven, but whoever practices and teaches these commands will be called great in the kingdom of heaven.
MATT|5|20|For I tell you that unless your righteousness surpasses that of the Pharisees and the teachers of the law, you will certainly not enter the kingdom of heaven.
MATT|5|21|"You have heard that it was said to the people long ago, 'Do not murder, and anyone who murders will be subject to judgment.'
MATT|5|22|But I tell you that anyone who is angry with his brother will be subject to judgment. Again, anyone who says to his brother, 'Raca, 'is answerable to the Sanhedrin. But anyone who says, 'You fool!' will be in danger of the fire of hell.
MATT|5|23|"Therefore, if you are offering your gift at the altar and there remember that your brother has something against you,
MATT|5|24|leave your gift there in front of the altar. First go and be reconciled to your brother; then come and offer your gift.
MATT|5|25|"Settle matters quickly with your adversary who is taking you to court. Do it while you are still with him on the way, or he may hand you over to the judge, and the judge may hand you over to the officer, and you may be thrown into prison.
MATT|5|26|I tell you the truth, you will not get out until you have paid the last penny.
MATT|5|27|"You have heard that it was said, 'Do not commit adultery.'
MATT|5|28|But I tell you that anyone who looks at a woman lustfully has already committed adultery with her in his heart.
MATT|5|29|If your right eye causes you to sin, gouge it out and throw it away. It is better for you to lose one part of your body than for your whole body to be thrown into hell.
MATT|5|30|And if your right hand causes you to sin, cut it off and throw it away. It is better for you to lose one part of your body than for your whole body to go into hell.
MATT|5|31|"It has been said, 'Anyone who divorces his wife must give her a certificate of divorce.'
MATT|5|32|But I tell you that anyone who divorces his wife, except for marital unfaithfulness, causes her to become an adulteress, and anyone who marries the divorced woman commits adultery.
MATT|5|33|"Again, you have heard that it was said to the people long ago, 'Do not break your oath, but keep the oaths you have made to the Lord.'
MATT|5|34|But I tell you, Do not swear at all: either by heaven, for it is God's throne;
MATT|5|35|or by the earth, for it is his footstool; or by Jerusalem, for it is the city of the Great King.
MATT|5|36|And do not swear by your head, for you cannot make even one hair white or black.
MATT|5|37|Simply let your 'Yes' be 'Yes,' and your 'No,No'; anything beyond this comes from the evil one.
MATT|5|38|"You have heard that it was said, 'Eye for eye, and tooth for tooth.'
MATT|5|39|But I tell you, Do not resist an evil person. If someone strikes you on the right cheek, turn to him the other also.
MATT|5|40|And if someone wants to sue you and take your tunic, let him have your cloak as well.
MATT|5|41|If someone forces you to go one mile, go with him two miles.
MATT|5|42|Give to the one who asks you, and do not turn away from the one who wants to borrow from you.
MATT|5|43|"You have heard that it was said, 'Love your neighbor and hate your enemy.'
MATT|5|44|But I tell you: Love your enemies and pray for those who persecute you,
MATT|5|45|that you may be sons of your Father in heaven. He causes his sun to rise on the evil and the good, and sends rain on the righteous and the unrighteous.
MATT|5|46|If you love those who love you, what reward will you get? Are not even the tax collectors doing that?
MATT|5|47|And if you greet only your brothers, what are you doing more than others? Do not even pagans do that?
MATT|5|48|Be perfect, therefore, as your heavenly Father is perfect.
MATT|6|1|"Be careful not to do your 'acts of righteousness' before men, to be seen by them. If you do, you will have no reward from your Father in heaven.
MATT|6|2|"So when you give to the needy, do not announce it with trumpets, as the hypocrites do in the synagogues and on the streets, to be honored by men. I tell you the truth, they have received their reward in full.
MATT|6|3|But when you give to the needy, do not let your left hand know what your right hand is doing,
MATT|6|4|so that your giving may be in secret. Then your Father, who sees what is done in secret, will reward you.
MATT|6|5|"And when you pray, do not be like the hypocrites, for they love to pray standing in the synagogues and on the street corners to be seen by men. I tell you the truth, they have received their reward in full.
MATT|6|6|But when you pray, go into your room, close the door and pray to your Father, who is unseen. Then your Father, who sees what is done in secret, will reward you.
MATT|6|7|And when you pray, do not keep on babbling like pagans, for they think they will be heard because of their many words.
MATT|6|8|Do not be like them, for your Father knows what you need before you ask him.
MATT|6|9|"This, then, is how you should pray: "'Our Father in heaven, hallowed be your name,
MATT|6|10|your kingdom come, your will be done on earth as it is in heaven.
MATT|6|11|Give us today our daily bread.
MATT|6|12|Forgive us our debts, as we also have forgiven our debtors.
MATT|6|13|And lead us not into temptation, but deliver us from the evil one. '
MATT|6|14|For if you forgive men when they sin against you, your heavenly Father will also forgive you.
MATT|6|15|But if you do not forgive men their sins, your Father will not forgive your sins.
MATT|6|16|"When you fast, do not look somber as the hypocrites do, for they disfigure their faces to show men they are fasting. I tell you the truth, they have received their reward in full.
MATT|6|17|But when you fast, put oil on your head and wash your face,
MATT|6|18|so that it will not be obvious to men that you are fasting, but only to your Father, who is unseen; and your Father, who sees what is done in secret, will reward you.
MATT|6|19|"Do not store up for yourselves treasures on earth, where moth and rust destroy, and where thieves break in and steal.
MATT|6|20|But store up for yourselves treasures in heaven, where moth and rust do not destroy, and where thieves do not break in and steal.
MATT|6|21|For where your treasure is, there your heart will be also.
MATT|6|22|"The eye is the lamp of the body. If your eyes are good, your whole body will be full of light.
MATT|6|23|But if your eyes are bad, your whole body will be full of darkness. If then the light within you is darkness, how great is that darkness!
MATT|6|24|"No one can serve two masters. Either he will hate the one and love the other, or he will be devoted to the one and despise the other. You cannot serve both God and Money.
MATT|6|25|"Therefore I tell you, do not worry about your life, what you will eat or drink; or about your body, what you will wear. Is not life more important than food, and the body more important than clothes?
MATT|6|26|Look at the birds of the air; they do not sow or reap or store away in barns, and yet your heavenly Father feeds them. Are you not much more valuable than they?
MATT|6|27|Who of you by worrying can add a single hour to his life?
MATT|6|28|"And why do you worry about clothes? See how the lilies of the field grow. They do not labor or spin.
MATT|6|29|Yet I tell you that not even Solomon in all his splendor was dressed like one of these.
MATT|6|30|If that is how God clothes the grass of the field, which is here today and tomorrow is thrown into the fire, will he not much more clothe you, O you of little faith?
MATT|6|31|So do not worry, saying, 'What shall we eat?' or 'What shall we drink?' or 'What shall we wear?'
MATT|6|32|For the pagans run after all these things, and your heavenly Father knows that you need them.
MATT|6|33|But seek first his kingdom and his righteousness, and all these things will be given to you as well.
MATT|6|34|Therefore do not worry about tomorrow, for tomorrow will worry about itself. Each day has enough trouble of its own.
MATT|7|1|"Do not judge, or you too will be judged.
MATT|7|2|For in the same way you judge others, you will be judged, and with the measure you use, it will be measured to you.
MATT|7|3|"Why do you look at the speck of sawdust in your brother's eye and pay no attention to the plank in your own eye?
MATT|7|4|How can you say to your brother, 'Let me take the speck out of your eye,' when all the time there is a plank in your own eye?
MATT|7|5|You hypocrite, first take the plank out of your own eye, and then you will see clearly to remove the speck from your brother's eye.
MATT|7|6|"Do not give dogs what is sacred; do not throw your pearls to pigs. If you do, they may trample them under their feet, and then turn and tear you to pieces.
MATT|7|7|"Ask and it will be given to you; seek and you will find; knock and the door will be opened to you.
MATT|7|8|For everyone who asks receives; he who seeks finds; and to him who knocks, the door will be opened.
MATT|7|9|"Which of you, if his son asks for bread, will give him a stone?
MATT|7|10|Or if he asks for a fish, will give him a snake?
MATT|7|11|If you, then, though you are evil, know how to give good gifts to your children, how much more will your Father in heaven give good gifts to those who ask him!
MATT|7|12|So in everything, do to others what you would have them do to you, for this sums up the Law and the Prophets.
MATT|7|13|"Enter through the narrow gate. For wide is the gate and broad is the road that leads to destruction, and many enter through it.
MATT|7|14|But small is the gate and narrow the road that leads to life, and only a few find it.
MATT|7|15|"Watch out for false prophets. They come to you in sheep's clothing, but inwardly they are ferocious wolves.
MATT|7|16|By their fruit you will recognize them. Do people pick grapes from thornbushes, or figs from thistles?
MATT|7|17|Likewise every good tree bears good fruit, but a bad tree bears bad fruit.
MATT|7|18|A good tree cannot bear bad fruit, and a bad tree cannot bear good fruit.
MATT|7|19|Every tree that does not bear good fruit is cut down and thrown into the fire.
MATT|7|20|Thus, by their fruit you will recognize them.
MATT|7|21|"Not everyone who says to me, 'Lord, Lord,' will enter the kingdom of heaven, but only he who does the will of my Father who is in heaven.
MATT|7|22|Many will say to me on that day, 'Lord, Lord, did we not prophesy in your name, and in your name drive out demons and perform many miracles?'
MATT|7|23|Then I will tell them plainly, 'I never knew you. Away from me, you evildoers!'
MATT|7|24|"Therefore everyone who hears these words of mine and puts them into practice is like a wise man who built his house on the rock.
MATT|7|25|The rain came down, the streams rose, and the winds blew and beat against that house; yet it did not fall, because it had its foundation on the rock.
MATT|7|26|But everyone who hears these words of mine and does not put them into practice is like a foolish man who built his house on sand.
MATT|7|27|The rain came down, the streams rose, and the winds blew and beat against that house, and it fell with a great crash."
MATT|7|28|When Jesus had finished saying these things, the crowds were amazed at his teaching,
MATT|7|29|because he taught as one who had authority, and not as their teachers of the law.
MATT|8|1|When he came down from the mountainside, large crowds followed him.
MATT|8|2|A man with leprosy came and knelt before him and said, "Lord, if you are willing, you can make me clean."
MATT|8|3|Jesus reached out his hand and touched the man. "I am willing," he said. "Be clean!" Immediately he was cured of his leprosy.
MATT|8|4|Then Jesus said to him, "See that you don't tell anyone. But go, show yourself to the priest and offer the gift Moses commanded, as a testimony to them."
MATT|8|5|When Jesus had entered Capernaum, a centurion came to him, asking for help.
MATT|8|6|"Lord," he said, "my servant lies at home paralyzed and in terrible suffering."
MATT|8|7|Jesus said to him, "I will go and heal him."
MATT|8|8|The centurion replied, "Lord, I do not deserve to have you come under my roof. But just say the word, and my servant will be healed.
MATT|8|9|For I myself am a man under authority, with soldiers under me. I tell this one, 'Go,' and he goes; and that one, 'Come,' and he comes. I say to my servant, 'Do this,' and he does it."
MATT|8|10|When Jesus heard this, he was astonished and said to those following him, "I tell you the truth, I have not found anyone in Israel with such great faith.
MATT|8|11|I say to you that many will come from the east and the west, and will take their places at the feast with Abraham, Isaac and Jacob in the kingdom of heaven.
MATT|8|12|But the subjects of the kingdom will be thrown outside, into the darkness, where there will be weeping and gnashing of teeth."
MATT|8|13|Then Jesus said to the centurion, "Go! It will be done just as you believed it would." And his servant was healed at that very hour.
MATT|8|14|When Jesus came into Peter's house, he saw Peter's mother-in-law lying in bed with a fever.
MATT|8|15|He touched her hand and the fever left her, and she got up and began to wait on him.
MATT|8|16|When evening came, many who were demon-possessed were brought to him, and he drove out the spirits with a word and healed all the sick.
MATT|8|17|This was to fulfill what was spoken through the prophet Isaiah: "He took up our infirmities and carried our diseases."
MATT|8|18|When Jesus saw the crowd around him, he gave orders to cross to the other side of the lake.
MATT|8|19|Then a teacher of the law came to him and said, "Teacher, I will follow you wherever you go."
MATT|8|20|Jesus replied, "Foxes have holes and birds of the air have nests, but the Son of Man has no place to lay his head."
MATT|8|21|Another disciple said to him, "Lord, first let me go and bury my father."
MATT|8|22|But Jesus told him, "Follow me, and let the dead bury their own dead."
MATT|8|23|Then he got into the boat and his disciples followed him.
MATT|8|24|Without warning, a furious storm came up on the lake, so that the waves swept over the boat. But Jesus was sleeping.
MATT|8|25|The disciples went and woke him, saying, "Lord, save us! We're going to drown!"
MATT|8|26|He replied, "You of little faith, why are you so afraid?" Then he got up and rebuked the winds and the waves, and it was completely calm.
MATT|8|27|The men were amazed and asked, "What kind of man is this? Even the winds and the waves obey him!"
MATT|8|28|When he arrived at the other side in the region of the Gadarenes, two demon-possessed men coming from the tombs met him. They were so violent that no one could pass that way.
MATT|8|29|"What do you want with us, Son of God?" they shouted. "Have you come here to torture us before the appointed time?"
MATT|8|30|Some distance from them a large herd of pigs was feeding.
MATT|8|31|The demons begged Jesus, "If you drive us out, send us into the herd of pigs."
MATT|8|32|He said to them, "Go!" So they came out and went into the pigs, and the whole herd rushed down the steep bank into the lake and died in the water.
MATT|8|33|Those tending the pigs ran off, went into the town and reported all this, including what had happened to the demon-possessed men.
MATT|8|34|Then the whole town went out to meet Jesus. And when they saw him, they pleaded with him to leave their region.
MATT|9|1|Jesus stepped into a boat, crossed over and came to his own town.
MATT|9|2|Some men brought to him a paralytic, lying on a mat. When Jesus saw their faith, he said to the paralytic, "Take heart, son; your sins are forgiven."
MATT|9|3|At this, some of the teachers of the law said to themselves, "This fellow is blaspheming!"
MATT|9|4|Knowing their thoughts, Jesus said, "Why do you entertain evil thoughts in your hearts?
MATT|9|5|Which is easier: to say, 'Your sins are forgiven,' or to say, 'Get up and walk'?
MATT|9|6|But so that you may know that the Son of Man has authority on earth to forgive sins...." Then he said to the paralytic, "Get up, take your mat and go home."
MATT|9|7|And the man got up and went home.
MATT|9|8|When the crowd saw this, they were filled with awe; and they praised God, who had given such authority to men.
MATT|9|9|As Jesus went on from there, he saw a man named Matthew sitting at the tax collector's booth. "Follow me," he told him, and Matthew got up and followed him.
MATT|9|10|While Jesus was having dinner at Matthew's house, many tax collectors and "sinners" came and ate with him and his disciples.
MATT|9|11|When the Pharisees saw this, they asked his disciples, "Why does your teacher eat with tax collectors and 'sinners'?"
MATT|9|12|On hearing this, Jesus said, "It is not the healthy who need a doctor, but the sick.
MATT|9|13|But go and learn what this means: 'I desire mercy, not sacrifice.' For I have not come to call the righteous, but sinners."
MATT|9|14|Then John's disciples came and asked him, "How is it that we and the Pharisees fast, but your disciples do not fast?"
MATT|9|15|Jesus answered, "How can the guests of the bridegroom mourn while he is with them? The time will come when the bridegroom will be taken from them; then they will fast.
MATT|9|16|"No one sews a patch of unshrunk cloth on an old garment, for the patch will pull away from the garment, making the tear worse.
MATT|9|17|Neither do men pour new wine into old wineskins. If they do, the skins will burst, the wine will run out and the wineskins will be ruined. No, they pour new wine into new wineskins, and both are preserved."
MATT|9|18|While he was saying this, a ruler came and knelt before him and said, "My daughter has just died. But come and put your hand on her, and she will live."
MATT|9|19|Jesus got up and went with him, and so did his disciples.
MATT|9|20|Just then a woman who had been subject to bleeding for twelve years came up behind him and touched the edge of his cloak.
MATT|9|21|She said to herself, "If I only touch his cloak, I will be healed."
MATT|9|22|Jesus turned and saw her. "Take heart, daughter," he said, "your faith has healed you." And the woman was healed from that moment.
MATT|9|23|When Jesus entered the ruler's house and saw the flute players and the noisy crowd,
MATT|9|24|he said, "Go away. The girl is not dead but asleep." But they laughed at him.
MATT|9|25|After the crowd had been put outside, he went in and took the girl by the hand, and she got up.
MATT|9|26|News of this spread through all that region.
MATT|9|27|As Jesus went on from there, two blind men followed him, calling out, "Have mercy on us, Son of David!"
MATT|9|28|When he had gone indoors, the blind men came to him, and he asked them, "Do you believe that I am able to do this?Yes, Lord," they replied.
MATT|9|29|Then he touched their eyes and said, "According to your faith will it be done to you";
MATT|9|30|and their sight was restored. Jesus warned them sternly, "See that no one knows about this."
MATT|9|31|But they went out and spread the news about him all over that region.
MATT|9|32|While they were going out, a man who was demon-possessed and could not talk was brought to Jesus.
MATT|9|33|And when the demon was driven out, the man who had been mute spoke. The crowd was amazed and said, "Nothing like this has ever been seen in Israel."
MATT|9|34|But the Pharisees said, "It is by the prince of demons that he drives out demons."
MATT|9|35|Jesus went through all the towns and villages, teaching in their synagogues, preaching the good news of the kingdom and healing every disease and sickness.
MATT|9|36|When he saw the crowds, he had compassion on them, because they were harassed and helpless, like sheep without a shepherd.
MATT|9|37|Then he said to his disciples, "The harvest is plentiful but the workers are few.
MATT|9|38|Ask the Lord of the harvest, therefore, to send out workers into his harvest field."
MATT|10|1|He called his twelve disciples to him and gave them authority to drive out evil spirits and to heal every disease and sickness.
MATT|10|2|These are the names of the twelve apostles: first, Simon (who is called Peter) and his brother Andrew; James son of Zebedee, and his brother John;
MATT|10|3|Philip and Bartholomew; Thomas and Matthew the tax collector; James son of Alphaeus, and Thaddaeus;
MATT|10|4|Simon the Zealot and Judas Iscariot, who betrayed him.
MATT|10|5|These twelve Jesus sent out with the following instructions: "Do not go among the Gentiles or enter any town of the Samaritans.
MATT|10|6|Go rather to the lost sheep of Israel.
MATT|10|7|As you go, preach this message: 'The kingdom of heaven is near.'
MATT|10|8|Heal the sick, raise the dead, cleanse those who have leprosy, drive out demons. Freely you have received, freely give.
MATT|10|9|Do not take along any gold or silver or copper in your belts;
MATT|10|10|take no bag for the journey, or extra tunic, or sandals or a staff; for the worker is worth his keep.
MATT|10|11|"Whatever town or village you enter, search for some worthy person there and stay at his house until you leave.
MATT|10|12|As you enter the home, give it your greeting.
MATT|10|13|If the home is deserving, let your peace rest on it; if it is not, let your peace return to you.
MATT|10|14|If anyone will not welcome you or listen to your words, shake the dust off your feet when you leave that home or town.
MATT|10|15|I tell you the truth, it will be more bearable for Sodom and Gomorrah on the day of judgment than for that town.
MATT|10|16|I am sending you out like sheep among wolves. Therefore be as shrewd as snakes and as innocent as doves.
MATT|10|17|"Be on your guard against men; they will hand you over to the local councils and flog you in their synagogues.
MATT|10|18|On my account you will be brought before governors and kings as witnesses to them and to the Gentiles.
MATT|10|19|But when they arrest you, do not worry about what to say or how to say it. At that time you will be given what to say,
MATT|10|20|for it will not be you speaking, but the Spirit of your Father speaking through you.
MATT|10|21|"Brother will betray brother to death, and a father his child; children will rebel against their parents and have them put to death.
MATT|10|22|All men will hate you because of me, but he who stands firm to the end will be saved.
MATT|10|23|When you are persecuted in one place, flee to another. I tell you the truth, you will not finish going through the cities of Israel before the Son of Man comes.
MATT|10|24|"A student is not above his teacher, nor a servant above his master.
MATT|10|25|It is enough for the student to be like his teacher, and the servant like his master. If the head of the house has been called Beelzebub, how much more the members of his household!
MATT|10|26|"So do not be afraid of them. There is nothing concealed that will not be disclosed, or hidden that will not be made known.
MATT|10|27|What I tell you in the dark, speak in the daylight; what is whispered in your ear, proclaim from the roofs.
MATT|10|28|Do not be afraid of those who kill the body but cannot kill the soul. Rather, be afraid of the One who can destroy both soul and body in hell.
MATT|10|29|Are not two sparrows sold for a penny? Yet not one of them will fall to the ground apart from the will of your Father.
MATT|10|30|And even the very hairs of your head are all numbered.
MATT|10|31|So don't be afraid; you are worth more than many sparrows.
MATT|10|32|"Whoever acknowledges me before men, I will also acknowledge him before my Father in heaven.
MATT|10|33|But whoever disowns me before men, I will disown him before my Father in heaven.
MATT|10|34|"Do not suppose that I have come to bring peace to the earth. I did not come to bring peace, but a sword.
MATT|10|35|For I have come to turn "'a man against his father, a daughter against her mother, a daughter-in-law against her mother-in-law--
MATT|10|36|a man's enemies will be the members of his own household.'
MATT|10|37|"Anyone who loves his father or mother more than me is not worthy of me; anyone who loves his son or daughter more than me is not worthy of me;
MATT|10|38|and anyone who does not take his cross and follow me is not worthy of me.
MATT|10|39|Whoever finds his life will lose it, and whoever loses his life for my sake will find it.
MATT|10|40|"He who receives you receives me, and he who receives me receives the one who sent me.
MATT|10|41|Anyone who receives a prophet because he is a prophet will receive a prophet's reward, and anyone who receives a righteous man because he is a righteous man will receive a righteous man's reward.
MATT|10|42|And if anyone gives even a cup of cold water to one of these little ones because he is my disciple, I tell you the truth, he will certainly not lose his reward."
MATT|11|1|After Jesus had finished instructing his twelve disciples, he went on from there to teach and preach in the towns of Galilee.
MATT|11|2|When John heard in prison what Christ was doing, he sent his disciples
MATT|11|3|to ask him, "Are you the one who was to come, or should we expect someone else?"
MATT|11|4|Jesus replied, "Go back and report to John what you hear and see:
MATT|11|5|The blind receive sight, the lame walk, those who have leprosy are cured, the deaf hear, the dead are raised, and the good news is preached to the poor.
MATT|11|6|Blessed is the man who does not fall away on account of me."
MATT|11|7|As John's disciples were leaving, Jesus began to speak to the crowd about John: "What did you go out into the desert to see? A reed swayed by the wind?
MATT|11|8|If not, what did you go out to see? A man dressed in fine clothes? No, those who wear fine clothes are in kings' palaces.
MATT|11|9|Then what did you go out to see? A prophet? Yes, I tell you, and more than a prophet.
MATT|11|10|This is the one about whom it is written: "'I will send my messenger ahead of you, who will prepare your way before you.'
MATT|11|11|I tell you the truth: Among those born of women there has not risen anyone greater than John the Baptist; yet he who is least in the kingdom of heaven is greater than he.
MATT|11|12|From the days of John the Baptist until now, the kingdom of heaven has been forcefully advancing, and forceful men lay hold of it.
MATT|11|13|For all the Prophets and the Law prophesied until John.
MATT|11|14|And if you are willing to accept it, he is the Elijah who was to come.
MATT|11|15|He who has ears, let him hear.
MATT|11|16|"To what can I compare this generation? They are like children sitting in the marketplaces and calling out to others:
MATT|11|17|"'We played the flute for you, and you did not dance; we sang a dirge and you did not mourn.'
MATT|11|18|For John came neither eating nor drinking, and they say, 'He has a demon.'
MATT|11|19|The Son of Man came eating and drinking, and they say, 'Here is a glutton and a drunkard, a friend of tax collectors and "sinners."' But wisdom is proved right by her actions."
MATT|11|20|Then Jesus began to denounce the cities in which most of his miracles had been performed, because they did not repent.
MATT|11|21|"Woe to you, Korazin! Woe to you, Bethsaida! If the miracles that were performed in you had been performed in Tyre and Sidon, they would have repented long ago in sackcloth and ashes.
MATT|11|22|But I tell you, it will be more bearable for Tyre and Sidon on the day of judgment than for you.
MATT|11|23|And you, Capernaum, will you be lifted up to the skies? No, you will go down to the depths. If the miracles that were performed in you had been performed in Sodom, it would have remained to this day.
MATT|11|24|But I tell you that it will be more bearable for Sodom on the day of judgment than for you."
MATT|11|25|At that time Jesus said, "I praise you, Father, Lord of heaven and earth, because you have hidden these things from the wise and learned, and revealed them to little children.
MATT|11|26|Yes, Father, for this was your good pleasure.
MATT|11|27|"All things have been committed to me by my Father. No one knows the Son except the Father, and no one knows the Father except the Son and those to whom the Son chooses to reveal him.
MATT|11|28|"Come to me, all you who are weary and burdened, and I will give you rest.
MATT|11|29|Take my yoke upon you and learn from me, for I am gentle and humble in heart, and you will find rest for your souls.
MATT|11|30|For my yoke is easy and my burden is light."
MATT|12|1|At that time Jesus went through the grainfields on the Sabbath. His disciples were hungry and began to pick some heads of grain and eat them.
MATT|12|2|When the Pharisees saw this, they said to him, "Look! Your disciples are doing what is unlawful on the Sabbath."
MATT|12|3|He answered, "Haven't you read what David did when he and his companions were hungry?
MATT|12|4|He entered the house of God, and he and his companions ate the consecrated bread--which was not lawful for them to do, but only for the priests.
MATT|12|5|Or haven't you read in the Law that on the Sabbath the priests in the temple desecrate the day and yet are innocent?
MATT|12|6|I tell you that one greater than the temple is here.
MATT|12|7|If you had known what these words mean, 'I desire mercy, not sacrifice,' you would not have condemned the innocent.
MATT|12|8|For the Son of Man is Lord of the Sabbath."
MATT|12|9|Going on from that place, he went into their synagogue,
MATT|12|10|and a man with a shriveled hand was there. Looking for a reason to accuse Jesus, they asked him, "Is it lawful to heal on the Sabbath?"
MATT|12|11|He said to them, "If any of you has a sheep and it falls into a pit on the Sabbath, will you not take hold of it and lift it out?
MATT|12|12|How much more valuable is a man than a sheep! Therefore it is lawful to do good on the Sabbath."
MATT|12|13|Then he said to the man, "Stretch out your hand." So he stretched it out and it was completely restored, just as sound as the other.
MATT|12|14|But the Pharisees went out and plotted how they might kill Jesus.
MATT|12|15|Aware of this, Jesus withdrew from that place. Many followed him, and he healed all their sick,
MATT|12|16|warning them not to tell who he was.
MATT|12|17|This was to fulfill what was spoken through the prophet Isaiah:
MATT|12|18|"Here is my servant whom I have chosen, the one I love, in whom I delight; I will put my Spirit on him, and he will proclaim justice to the nations.
MATT|12|19|He will not quarrel or cry out; no one will hear his voice in the streets.
MATT|12|20|A bruised reed he will not break, and a smoldering wick he will not snuff out, till he leads justice to victory.
MATT|12|21|In his name the nations will put their hope."
MATT|12|22|Then they brought him a demon-possessed man who was blind and mute, and Jesus healed him, so that he could both talk and see.
MATT|12|23|All the people were astonished and said, "Could this be the Son of David?"
MATT|12|24|But when the Pharisees heard this, they said, "It is only by Beelzebub, the prince of demons, that this fellow drives out demons."
MATT|12|25|Jesus knew their thoughts and said to them, "Every kingdom divided against itself will be ruined, and every city or household divided against itself will not stand.
MATT|12|26|If Satan drives out Satan, he is divided against himself. How then can his kingdom stand?
MATT|12|27|And if I drive out demons by Beelzebub, by whom do your people drive them out? So then, they will be your judges.
MATT|12|28|But if I drive out demons by the Spirit of God, then the kingdom of God has come upon you.
MATT|12|29|"Or again, how can anyone enter a strong man's house and carry off his possessions unless he first ties up the strong man? Then he can rob his house.
MATT|12|30|"He who is not with me is against me, and he who does not gather with me scatters.
MATT|12|31|And so I tell you, every sin and blasphemy will be forgiven men, but the blasphemy against the Spirit will not be forgiven.
MATT|12|32|Anyone who speaks a word against the Son of Man will be forgiven, but anyone who speaks against the Holy Spirit will not be forgiven, either in this age or in the age to come.
MATT|12|33|"Make a tree good and its fruit will be good, or make a tree bad and its fruit will be bad, for a tree is recognized by its fruit.
MATT|12|34|You brood of vipers, how can you who are evil say anything good? For out of the overflow of the heart the mouth speaks.
MATT|12|35|The good man brings good things out of the good stored up in him, and the evil man brings evil things out of the evil stored up in him.
MATT|12|36|But I tell you that men will have to give account on the day of judgment for every careless word they have spoken.
MATT|12|37|For by your words you will be acquitted, and by your words you will be condemned."
MATT|12|38|Then some of the Pharisees and teachers of the law said to him, "Teacher, we want to see a miraculous sign from you."
MATT|12|39|He answered, "A wicked and adulterous generation asks for a miraculous sign! But none will be given it except the sign of the prophet Jonah.
MATT|12|40|For as Jonah was three days and three nights in the belly of a huge fish, so the Son of Man will be three days and three nights in the heart of the earth.
MATT|12|41|The men of Nineveh will stand up at the judgment with this generation and condemn it; for they repented at the preaching of Jonah, and now one greater than Jonah is here.
MATT|12|42|The Queen of the South will rise at the judgment with this generation and condemn it; for she came from the ends of the earth to listen to Solomon's wisdom, and now one greater than Solomon is here.
MATT|12|43|"When an evil spirit comes out of a man, it goes through arid places seeking rest and does not find it.
MATT|12|44|Then it says, 'I will return to the house I left.' When it arrives, it finds the house unoccupied, swept clean and put in order.
MATT|12|45|Then it goes and takes with it seven other spirits more wicked than itself, and they go in and live there. And the final condition of that man is worse than the first. That is how it will be with this wicked generation."
MATT|12|46|While Jesus was still talking to the crowd, his mother and brothers stood outside, wanting to speak to him.
MATT|12|47|Someone told him, "Your mother and brothers are standing outside, wanting to speak to you."
MATT|12|48|He replied to him, "Who is my mother, and who are my brothers?"
MATT|12|49|Pointing to his disciples, he said, "Here are my mother and my brothers.
MATT|12|50|For whoever does the will of my Father in heaven is my brother and sister and mother."
MATT|13|1|That same day Jesus went out of the house and sat by the lake.
MATT|13|2|Such large crowds gathered around him that he got into a boat and sat in it, while all the people stood on the shore.
MATT|13|3|Then he told them many things in parables, saying: "A farmer went out to sow his seed.
MATT|13|4|As he was scattering the seed, some fell along the path, and the birds came and ate it up.
MATT|13|5|Some fell on rocky places, where it did not have much soil. It sprang up quickly, because the soil was shallow.
MATT|13|6|But when the sun came up, the plants were scorched, and they withered because they had no root.
MATT|13|7|Other seed fell among thorns, which grew up and choked the plants.
MATT|13|8|Still other seed fell on good soil, where it produced a crop--a hundred, sixty or thirty times what was sown.
MATT|13|9|He who has ears, let him hear."
MATT|13|10|The disciples came to him and asked, "Why do you speak to the people in parables?"
MATT|13|11|He replied, "The knowledge of the secrets of the kingdom of heaven has been given to you, but not to them.
MATT|13|12|Whoever has will be given more, and he will have an abundance. Whoever does not have, even what he has will be taken from him.
MATT|13|13|This is why I speak to them in parables: "Though seeing, they do not see; though hearing, they do not hear or understand.
MATT|13|14|In them is fulfilled the prophecy of Isaiah: "'You will be ever hearing but never understanding; you will be ever seeing but never perceiving.
MATT|13|15|For this people's heart has become calloused; they hardly hear with their ears, and they have closed their eyes. Otherwise they might see with their eyes, hear with their ears, understand with their hearts and turn, and I would heal them.'
MATT|13|16|But blessed are your eyes because they see, and your ears because they hear.
MATT|13|17|For I tell you the truth, many prophets and righteous men longed to see what you see but did not see it, and to hear what you hear but did not hear it.
MATT|13|18|"Listen then to what the parable of the sower means:
MATT|13|19|When anyone hears the message about the kingdom and does not understand it, the evil one comes and snatches away what was sown in his heart. This is the seed sown along the path.
MATT|13|20|The one who received the seed that fell on rocky places is the man who hears the word and at once receives it with joy.
MATT|13|21|But since he has no root, he lasts only a short time. When trouble or persecution comes because of the word, he quickly falls away.
MATT|13|22|The one who received the seed that fell among the thorns is the man who hears the word, but the worries of this life and the deceitfulness of wealth choke it, making it unfruitful.
MATT|13|23|But the one who received the seed that fell on good soil is the man who hears the word and understands it. He produces a crop, yielding a hundred, sixty or thirty times what was sown."
MATT|13|24|Jesus told them another parable: "The kingdom of heaven is like a man who sowed good seed in his field.
MATT|13|25|But while everyone was sleeping, his enemy came and sowed weeds among the wheat, and went away.
MATT|13|26|When the wheat sprouted and formed heads, then the weeds also appeared.
MATT|13|27|"The owner's servants came to him and said, 'Sir, didn't you sow good seed in your field? Where then did the weeds come from?'
MATT|13|28|"'An enemy did this,' he replied. "The servants asked him, 'Do you want us to go and pull them up?'
MATT|13|29|"'No,' he answered, 'because while you are pulling the weeds, you may root up the wheat with them.
MATT|13|30|Let both grow together until the harvest. At that time I will tell the harvesters: First collect the weeds and tie them in bundles to be burned; then gather the wheat and bring it into my barn.'"
MATT|13|31|He told them another parable: "The kingdom of heaven is like a mustard seed, which a man took and planted in his field.
MATT|13|32|Though it is the smallest of all your seeds, yet when it grows, it is the largest of garden plants and becomes a tree, so that the birds of the air come and perch in its branches."
MATT|13|33|He told them still another parable: "The kingdom of heaven is like yeast that a woman took and mixed into a large amount of flour until it worked all through the dough."
MATT|13|34|Jesus spoke all these things to the crowd in parables; he did not say anything to them without using a parable.
MATT|13|35|So was fulfilled what was spoken through the prophet: "I will open my mouth in parables, I will utter things hidden since the creation of the world."
MATT|13|36|Then he left the crowd and went into the house. His disciples came to him and said, "Explain to us the parable of the weeds in the field."
MATT|13|37|He answered, "The one who sowed the good seed is the Son of Man.
MATT|13|38|The field is the world, and the good seed stands for the sons of the kingdom. The weeds are the sons of the evil one,
MATT|13|39|and the enemy who sows them is the devil. The harvest is the end of the age, and the harvesters are angels.
MATT|13|40|"As the weeds are pulled up and burned in the fire, so it will be at the end of the age.
MATT|13|41|The Son of Man will send out his angels, and they will weed out of his kingdom everything that causes sin and all who do evil.
MATT|13|42|They will throw them into the fiery furnace, where there will be weeping and gnashing of teeth.
MATT|13|43|Then the righteous will shine like the sun in the kingdom of their Father. He who has ears, let him hear.
MATT|13|44|"The kingdom of heaven is like treasure hidden in a field. When a man found it, he hid it again, and then in his joy went and sold all he had and bought that field.
MATT|13|45|"Again, the kingdom of heaven is like a merchant looking for fine pearls.
MATT|13|46|When he found one of great value, he went away and sold everything he had and bought it.
MATT|13|47|"Once again, the kingdom of heaven is like a net that was let down into the lake and caught all kinds of fish.
MATT|13|48|When it was full, the fishermen pulled it up on the shore. Then they sat down and collected the good fish in baskets, but threw the bad away.
MATT|13|49|This is how it will be at the end of the age. The angels will come and separate the wicked from the righteous
MATT|13|50|and throw them into the fiery furnace, where there will be weeping and gnashing of teeth.
MATT|13|51|"Have you understood all these things?" Jesus asked. "Yes," they replied.
MATT|13|52|He said to them, "Therefore every teacher of the law who has been instructed about the kingdom of heaven is like the owner of a house who brings out of his storeroom new treasures as well as old."
MATT|13|53|When Jesus had finished these parables, he moved on from there.
MATT|13|54|Coming to his hometown, he began teaching the people in their synagogue, and they were amazed. "Where did this man get this wisdom and these miraculous powers?" they asked.
MATT|13|55|"Isn't this the carpenter's son? Isn't his mother's name Mary, and aren't his brothers James, Joseph, Simon and Judas?
MATT|13|56|Aren't all his sisters with us? Where then did this man get all these things?"
MATT|13|57|And they took offense at him. But Jesus said to them, "Only in his hometown and in his own house is a prophet without honor."
MATT|13|58|And he did not do many miracles there because of their lack of faith.
MATT|14|1|At that time Herod the tetrarch heard the reports about Jesus,
MATT|14|2|and he said to his attendants, "This is John the Baptist; he has risen from the dead! That is why miraculous powers are at work in him."
MATT|14|3|Now Herod had arrested John and bound him and put him in prison because of Herodias, his brother Philip's wife,
MATT|14|4|for John had been saying to him: "It is not lawful for you to have her."
MATT|14|5|Herod wanted to kill John, but he was afraid of the people, because they considered him a prophet.
MATT|14|6|On Herod's birthday the daughter of Herodias danced for them and pleased Herod so much
MATT|14|7|that he promised with an oath to give her whatever she asked.
MATT|14|8|Prompted by her mother, she said, "Give me here on a platter the head of John the Baptist."
MATT|14|9|The king was distressed, but because of his oaths and his dinner guests, he ordered that her request be granted
MATT|14|10|and had John beheaded in the prison.
MATT|14|11|His head was brought in on a platter and given to the girl, who carried it to her mother.
MATT|14|12|John's disciples came and took his body and buried it. Then they went and told Jesus.
MATT|14|13|When Jesus heard what had happened, he withdrew by boat privately to a solitary place. Hearing of this, the crowds followed him on foot from the towns.
MATT|14|14|When Jesus landed and saw a large crowd, he had compassion on them and healed their sick.
MATT|14|15|As evening approached, the disciples came to him and said, "This is a remote place, and it's already getting late. Send the crowds away, so they can go to the villages and buy themselves some food."
MATT|14|16|Jesus replied, "They do not need to go away. You give them something to eat."
MATT|14|17|"We have here only five loaves of bread and two fish," they answered.
MATT|14|18|"Bring them here to me," he said.
MATT|14|19|And he directed the people to sit down on the grass. Taking the five loaves and the two fish and looking up to heaven, he gave thanks and broke the loaves. Then he gave them to the disciples, and the disciples gave them to the people.
MATT|14|20|They all ate and were satisfied, and the disciples picked up twelve basketfuls of broken pieces that were left over.
MATT|14|21|The number of those who ate was about five thousand men, besides women and children.
MATT|14|22|Immediately Jesus made the disciples get into the boat and go on ahead of him to the other side, while he dismissed the crowd.
MATT|14|23|After he had dismissed them, he went up on a mountainside by himself to pray. When evening came, he was there alone,
MATT|14|24|but the boat was already a considerable distance from land, buffeted by the waves because the wind was against it.
MATT|14|25|During the fourth watch of the night Jesus went out to them, walking on the lake.
MATT|14|26|When the disciples saw him walking on the lake, they were terrified. "It's a ghost," they said, and cried out in fear.
MATT|14|27|But Jesus immediately said to them: "Take courage! It is I. Don't be afraid."
MATT|14|28|"Lord, if it's you," Peter replied, "tell me to come to you on the water."
MATT|14|29|"Come," he said.
MATT|14|30|Then Peter got down out of the boat, walked on the water and came toward Jesus. But when he saw the wind, he was afraid and, beginning to sink, cried out, "Lord, save me!"
MATT|14|31|Immediately Jesus reached out his hand and caught him. "You of little faith," he said, "why did you doubt?"
MATT|14|32|And when they climbed into the boat, the wind died down.
MATT|14|33|Then those who were in the boat worshiped him, saying, "Truly you are the Son of God."
MATT|14|34|When they had crossed over, they landed at Gennesaret.
MATT|14|35|And when the men of that place recognized Jesus, they sent word to all the surrounding country. People brought all their sick to him
MATT|14|36|and begged him to let the sick just touch the edge of his cloak, and all who touched him were healed.
MATT|15|1|Then some Pharisees and teachers of the law came to Jesus from Jerusalem and asked,
MATT|15|2|"Why do your disciples break the tradition of the elders? They don't wash their hands before they eat!"
MATT|15|3|Jesus replied, "And why do you break the command of God for the sake of your tradition?
MATT|15|4|For God said, 'Honor your father and mother' and 'Anyone who curses his father or mother must be put to death.'
MATT|15|5|But you say that if a man says to his father or mother, 'Whatever help you might otherwise have received from me is a gift devoted to God,'
MATT|15|6|he is not to 'honor his father 'with it. Thus you nullify the word of God for the sake of your tradition.
MATT|15|7|You hypocrites! Isaiah was right when he prophesied about you:
MATT|15|8|"'These people honor me with their lips, but their hearts are far from me.
MATT|15|9|They worship me in vain; their teachings are but rules taught by men.'"
MATT|15|10|Jesus called the crowd to him and said, "Listen and understand.
MATT|15|11|What goes into a man's mouth does not make him 'unclean,' but what comes out of his mouth, that is what makes him 'unclean.'"
MATT|15|12|Then the disciples came to him and asked, "Do you know that the Pharisees were offended when they heard this?"
MATT|15|13|He replied, "Every plant that my heavenly Father has not planted will be pulled up by the roots.
MATT|15|14|Leave them; they are blind guides. If a blind man leads a blind man, both will fall into a pit."
MATT|15|15|Peter said, "Explain the parable to us."
MATT|15|16|"Are you still so dull?" Jesus asked them.
MATT|15|17|"Don't you see that whatever enters the mouth goes into the stomach and then out of the body?
MATT|15|18|But the things that come out of the mouth come from the heart, and these make a man 'unclean.'
MATT|15|19|For out of the heart come evil thoughts, murder, adultery, sexual immorality, theft, false testimony, slander.
MATT|15|20|These are what make a man 'unclean'; but eating with unwashed hands does not make him 'unclean.'"
MATT|15|21|Leaving that place, Jesus withdrew to the region of Tyre and Sidon.
MATT|15|22|A Canaanite woman from that vicinity came to him, crying out, "Lord, Son of David, have mercy on me! My daughter is suffering terribly from demon-possession."
MATT|15|23|Jesus did not answer a word. So his disciples came to him and urged him, "Send her away, for she keeps crying out after us."
MATT|15|24|He answered, "I was sent only to the lost sheep of Israel."
MATT|15|25|The woman came and knelt before him. "Lord, help me!" she said.
MATT|15|26|He replied, "It is not right to take the children's bread and toss it to their dogs."
MATT|15|27|"Yes, Lord," she said, "but even the dogs eat the crumbs that fall from their masters' table."
MATT|15|28|Then Jesus answered, "Woman, you have great faith! Your request is granted." And her daughter was healed from that very hour.
MATT|15|29|Jesus left there and went along the Sea of Galilee. Then he went up on a mountainside and sat down.
MATT|15|30|Great crowds came to him, bringing the lame, the blind, the crippled, the mute and many others, and laid them at his feet; and he healed them.
MATT|15|31|The people were amazed when they saw the mute speaking, the crippled made well, the lame walking and the blind seeing. And they praised the God of Israel.
MATT|15|32|Jesus called his disciples to him and said, "I have compassion for these people; they have already been with me three days and have nothing to eat. I do not want to send them away hungry, or they may collapse on the way."
MATT|15|33|His disciples answered, "Where could we get enough bread in this remote place to feed such a crowd?"
MATT|15|34|"How many loaves do you have?" Jesus asked. "Seven," they replied, "and a few small fish."
MATT|15|35|He told the crowd to sit down on the ground.
MATT|15|36|Then he took the seven loaves and the fish, and when he had given thanks, he broke them and gave them to the disciples, and they in turn to the people.
MATT|15|37|They all ate and were satisfied. Afterward the disciples picked up seven basketfuls of broken pieces that were left over.
MATT|15|38|The number of those who ate was four thousand, besides women and children.
MATT|15|39|After Jesus had sent the crowd away, he got into the boat and went to the vicinity of Magadan.
MATT|16|1|The Pharisees and Sadducees came to Jesus and tested him by asking him to show them a sign from heaven.
MATT|16|2|He replied, "When evening comes, you say, 'It will be fair weather, for the sky is red,'
MATT|16|3|and in the morning, 'Today it will be stormy, for the sky is red and overcast.' You know how to interpret the appearance of the sky, but you cannot interpret the signs of the times.
MATT|16|4|A wicked and adulterous generation looks for a miraculous sign, but none will be given it except the sign of Jonah." Jesus then left them and went away.
MATT|16|5|When they went across the lake, the disciples forgot to take bread.
MATT|16|6|"Be careful," Jesus said to them. "Be on your guard against the yeast of the Pharisees and Sadducees."
MATT|16|7|They discussed this among themselves and said, "It is because we didn't bring any bread."
MATT|16|8|Aware of their discussion, Jesus asked, "You of little faith, why are you talking among yourselves about having no bread?
MATT|16|9|Do you still not understand? Don't you remember the five loaves for the five thousand, and how many basketfuls you gathered?
MATT|16|10|Or the seven loaves for the four thousand, and how many basketfuls you gathered?
MATT|16|11|How is it you don't understand that I was not talking to you about bread? But be on your guard against the yeast of the Pharisees and Sadducees."
MATT|16|12|Then they understood that he was not telling them to guard against the yeast used in bread, but against the teaching of the Pharisees and Sadducees.
MATT|16|13|When Jesus came to the region of Caesarea Philippi, he asked his disciples, "Who do people say the Son of Man is?"
MATT|16|14|They replied, "Some say John the Baptist; others say Elijah; and still others, Jeremiah or one of the prophets."
MATT|16|15|"But what about you?" he asked. "Who do you say I am?"
MATT|16|16|Simon Peter answered, "You are the Christ, the Son of the living God."
MATT|16|17|Jesus replied, "Blessed are you, Simon son of Jonah, for this was not revealed to you by man, but by my Father in heaven.
MATT|16|18|And I tell you that you are Peter, and on this rock I will build my church, and the gates of Hades will not overcome it.
MATT|16|19|I will give you the keys of the kingdom of heaven; whatever you bind on earth will be bound in heaven, and whatever you loose on earth will be loosed in heaven."
MATT|16|20|Then he warned his disciples not to tell anyone that he was the Christ.
MATT|16|21|From that time on Jesus began to explain to his disciples that he must go to Jerusalem and suffer many things at the hands of the elders, chief priests and teachers of the law, and that he must be killed and on the third day be raised to life.
MATT|16|22|Peter took him aside and began to rebuke him. "Never, Lord!" he said. "This shall never happen to you!"
MATT|16|23|Jesus turned and said to Peter, "Get behind me, Satan! You are a stumbling block to me; you do not have in mind the things of God, but the things of men."
MATT|16|24|Then Jesus said to his disciples, "If anyone would come after me, he must deny himself and take up his cross and follow me.
MATT|16|25|For whoever wants to save his life will lose it, but whoever loses his life for me will find it.
MATT|16|26|What good will it be for a man if he gains the whole world, yet forfeits his soul? Or what can a man give in exchange for his soul?
MATT|16|27|For the Son of Man is going to come in his Father's glory with his angels, and then he will reward each person according to what he has done.
MATT|16|28|I tell you the truth, some who are standing here will not taste death before they see the Son of Man coming in his kingdom."
MATT|17|1|After six days Jesus took with him Peter, James and John the brother of James, and led them up a high mountain by themselves.
MATT|17|2|There he was transfigured before them. His face shone like the sun, and his clothes became as white as the light.
MATT|17|3|Just then there appeared before them Moses and Elijah, talking with Jesus.
MATT|17|4|Peter said to Jesus, "Lord, it is good for us to be here. If you wish, I will put up three shelters--one for you, one for Moses and one for Elijah."
MATT|17|5|While he was still speaking, a bright cloud enveloped them, and a voice from the cloud said, "This is my Son, whom I love; with him I am well pleased. Listen to him!"
MATT|17|6|When the disciples heard this, they fell facedown to the ground, terrified.
MATT|17|7|But Jesus came and touched them. "Get up," he said. "Don't be afraid."
MATT|17|8|When they looked up, they saw no one except Jesus.
MATT|17|9|As they were coming down the mountain, Jesus instructed them, "Don't tell anyone what you have seen, until the Son of Man has been raised from the dead."
MATT|17|10|The disciples asked him, "Why then do the teachers of the law say that Elijah must come first?"
MATT|17|11|Jesus replied, "To be sure, Elijah comes and will restore all things.
MATT|17|12|But I tell you, Elijah has already come, and they did not recognize him, but have done to him everything they wished. In the same way the Son of Man is going to suffer at their hands."
MATT|17|13|Then the disciples understood that he was talking to them about John the Baptist.
MATT|17|14|When they came to the crowd, a man approached Jesus and knelt before him.
MATT|17|15|"Lord, have mercy on my son," he said. "He has seizures and is suffering greatly. He often falls into the fire or into the water.
MATT|17|16|I brought him to your disciples, but they could not heal him."
MATT|17|17|"O unbelieving and perverse generation," Jesus replied, "how long shall I stay with you? How long shall I put up with you? Bring the boy here to me."
MATT|17|18|Jesus rebuked the demon, and it came out of the boy, and he was healed from that moment.
MATT|17|19|Then the disciples came to Jesus in private and asked, "Why couldn't we drive it out?"
MATT|17|20|He replied, "Because you have so little faith. I tell you the truth, if you have faith as small as a mustard seed, you can say to this mountain, 'Move from here to there' and it will move. Nothing will be impossible for you."
MATT|17|21|See Footnote
MATT|17|22|When they came together in Galilee, he said to them, "The Son of Man is going to be betrayed into the hands of men.
MATT|17|23|They will kill him, and on the third day he will be raised to life." And the disciples were filled with grief.
MATT|17|24|After Jesus and his disciples arrived in Capernaum, the collectors of the two-drachma tax came to Peter and asked, "Doesn't your teacher pay the temple tax?"
MATT|17|25|"Yes, he does," he replied. When Peter came into the house, Jesus was the first to speak. "What do you think, Simon?" he asked. "From whom do the kings of the earth collect duty and taxes--from their own sons or from others?"
MATT|17|26|"From others," Peter answered.
MATT|17|27|"Then the sons are exempt," Jesus said to him. "But so that we may not offend them, go to the lake and throw out your line. Take the first fish you catch; open its mouth and you will find a four-drachma coin. Take it and give it to them for my tax and yours."
MATT|18|1|At that time the disciples came to Jesus and asked, "Who is the greatest in the kingdom of heaven?"
MATT|18|2|He called a little child and had him stand among them.
MATT|18|3|And he said: "I tell you the truth, unless you change and become like little children, you will never enter the kingdom of heaven.
MATT|18|4|Therefore, whoever humbles himself like this child is the greatest in the kingdom of heaven.
MATT|18|5|"And whoever welcomes a little child like this in my name welcomes me.
MATT|18|6|But if anyone causes one of these little ones who believe in me to sin, it would be better for him to have a large millstone hung around his neck and to be drowned in the depths of the sea.
MATT|18|7|"Woe to the world because of the things that cause people to sin! Such things must come, but woe to the man through whom they come!
MATT|18|8|If your hand or your foot causes you to sin, cut it off and throw it away. It is better for you to enter life maimed or crippled than to have two hands or two feet and be thrown into eternal fire.
MATT|18|9|And if your eye causes you to sin, gouge it out and throw it away. It is better for you to enter life with one eye than to have two eyes and be thrown into the fire of hell.
MATT|18|10|"See that you do not look down on one of these little ones. For I tell you that their angels in heaven always see the face of my Father in heaven.
MATT|18|11|See Footnote
MATT|18|12|"What do you think? If a man owns a hundred sheep, and one of them wanders away, will he not leave the ninety-nine on the hills and go to look for the one that wandered off?
MATT|18|13|And if he finds it, I tell you the truth, he is happier about that one sheep than about the ninety-nine that did not wander off.
MATT|18|14|In the same way your Father in heaven is not willing that any of these little ones should be lost.
MATT|18|15|"If your brother sins against you, go and show him his fault, just between the two of you. If he listens to you, you have won your brother over.
MATT|18|16|But if he will not listen, take one or two others along, so that 'every matter may be established by the testimony of two or three witnesses.'
MATT|18|17|If he refuses to listen to them, tell it to the church; and if he refuses to listen even to the church, treat him as you would a pagan or a tax collector.
MATT|18|18|"I tell you the truth, whatever you bind on earth will be bound in heaven, and whatever you loose on earth will be loosed in heaven.
MATT|18|19|"Again, I tell you that if two of you on earth agree about anything you ask for, it will be done for you by my Father in heaven.
MATT|18|20|For where two or three come together in my name, there am I with them."
MATT|18|21|Then Peter came to Jesus and asked, "Lord, how many times shall I forgive my brother when he sins against me? Up to seven times?"
MATT|18|22|Jesus answered, "I tell you, not seven times, but seventy-seven times.
MATT|18|23|"Therefore, the kingdom of heaven is like a king who wanted to settle accounts with his servants.
MATT|18|24|As he began the settlement, a man who owed him ten thousand talents was brought to him.
MATT|18|25|Since he was not able to pay, the master ordered that he and his wife and his children and all that he had be sold to repay the debt.
MATT|18|26|"The servant fell on his knees before him. 'Be patient with me,' he begged, 'and I will pay back everything.'
MATT|18|27|The servant's master took pity on him, canceled the debt and let him go.
MATT|18|28|"But when that servant went out, he found one of his fellow servants who owed him a hundred denarii. He grabbed him and began to choke him. 'Pay back what you owe me!' he demanded.
MATT|18|29|"His fellow servant fell to his knees and begged him, 'Be patient with me, and I will pay you back.'
MATT|18|30|"But he refused. Instead, he went off and had the man thrown into prison until he could pay the debt.
MATT|18|31|When the other servants saw what had happened, they were greatly distressed and went and told their master everything that had happened.
MATT|18|32|"Then the master called the servant in. 'You wicked servant,' he said, 'I canceled all that debt of yours because you begged me to.
MATT|18|33|Shouldn't you have had mercy on your fellow servant just as I had on you?'
MATT|18|34|In anger his master turned him over to the jailers to be tortured, until he should pay back all he owed.
MATT|18|35|"This is how my heavenly Father will treat each of you unless you forgive your brother from your heart."
MATT|19|1|When Jesus had finished saying these things, he left Galilee and went into the region of Judea to the other side of the Jordan.
MATT|19|2|Large crowds followed him, and he healed them there.
MATT|19|3|Some Pharisees came to him to test him. They asked, "Is it lawful for a man to divorce his wife for any and every reason?"
MATT|19|4|"Haven't you read," he replied, "that at the beginning the Creator 'made them male and female,'
MATT|19|5|and said, 'For this reason a man will leave his father and mother and be united to his wife, and the two will become one flesh'?
MATT|19|6|So they are no longer two, but one. Therefore what God has joined together, let man not separate."
MATT|19|7|"Why then," they asked, "did Moses command that a man give his wife a certificate of divorce and send her away?"
MATT|19|8|Jesus replied, "Moses permitted you to divorce your wives because your hearts were hard. But it was not this way from the beginning.
MATT|19|9|I tell you that anyone who divorces his wife, except for marital unfaithfulness, and marries another woman commits adultery."
MATT|19|10|The disciples said to him, "If this is the situation between a husband and wife, it is better not to marry."
MATT|19|11|Jesus replied, "Not everyone can accept this word, but only those to whom it has been given.
MATT|19|12|For some are eunuchs because they were born that way; others were made that way by men; and others have renounced marriage because of the kingdom of heaven. The one who can accept this should accept it."
MATT|19|13|Then little children were brought to Jesus for him to place his hands on them and pray for them. But the disciples rebuked those who brought them.
MATT|19|14|Jesus said, "Let the little children come to me, and do not hinder them, for the kingdom of heaven belongs to such as these."
MATT|19|15|When he had placed his hands on them, he went on from there.
MATT|19|16|Now a man came up to Jesus and asked, "Teacher, what good thing must I do to get eternal life?"
MATT|19|17|"Why do you ask me about what is good?" Jesus replied. "There is only One who is good. If you want to enter life, obey the commandments."
MATT|19|18|"Which ones?" the man inquired.
MATT|19|19|Jesus replied, "'Do not murder, do not commit adultery, do not steal, do not give false testimony, honor your father and mother,' and 'love your neighbor as yourself.'"
MATT|19|20|"All these I have kept," the young man said. "What do I still lack?"
MATT|19|21|Jesus answered, "If you want to be perfect, go, sell your possessions and give to the poor, and you will have treasure in heaven. Then come, follow me."
MATT|19|22|When the young man heard this, he went away sad, because he had great wealth.
MATT|19|23|Then Jesus said to his disciples, "I tell you the truth, it is hard for a rich man to enter the kingdom of heaven.
MATT|19|24|Again I tell you, it is easier for a camel to go through the eye of a needle than for a rich man to enter the kingdom of God."
MATT|19|25|When the disciples heard this, they were greatly astonished and asked, "Who then can be saved?"
MATT|19|26|Jesus looked at them and said, "With man this is impossible, but with God all things are possible."
MATT|19|27|Peter answered him, "We have left everything to follow you! What then will there be for us?"
MATT|19|28|Jesus said to them, "I tell you the truth, at the renewal of all things, when the Son of Man sits on his glorious throne, you who have followed me will also sit on twelve thrones, judging the twelve tribes of Israel.
MATT|19|29|And everyone who has left houses or brothers or sisters or father or mother or children or fields for my sake will receive a hundred times as much and will inherit eternal life.
MATT|19|30|But many who are first will be last, and many who are last will be first.
MATT|20|1|"For the kingdom of heaven is like a landowner who went out early in the morning to hire men to work in his vineyard.
MATT|20|2|He agreed to pay them a denarius for the day and sent them into his vineyard.
MATT|20|3|"About the third hour he went out and saw others standing in the marketplace doing nothing.
MATT|20|4|He told them, 'You also go and work in my vineyard, and I will pay you whatever is right.'
MATT|20|5|So they went.
MATT|20|6|"He went out again about the sixth hour and the ninth hour and did the same thing. About the eleventh hour he went out and found still others standing around. He asked them, 'Why have you been standing here all day long doing nothing?'
MATT|20|7|"'Because no one has hired us,' they answered. "He said to them, 'You also go and work in my vineyard.'
MATT|20|8|"When evening came, the owner of the vineyard said to his foreman, 'Call the workers and pay them their wages, beginning with the last ones hired and going on to the first.'
MATT|20|9|"The workers who were hired about the eleventh hour came and each received a denarius.
MATT|20|10|So when those came who were hired first, they expected to receive more. But each one of them also received a denarius.
MATT|20|11|When they received it, they began to grumble against the landowner.
MATT|20|12|'These men who were hired last worked only one hour,' they said, 'and you have made them equal to us who have borne the burden of the work and the heat of the day.'
MATT|20|13|"But he answered one of them, 'Friend, I am not being unfair to you. Didn't you agree to work for a denarius?
MATT|20|14|Take your pay and go. I want to give the man who was hired last the same as I gave you.
MATT|20|15|Don't I have the right to do what I want with my own money? Or are you envious because I am generous?'
MATT|20|16|"So the last will be first, and the first will be last."
MATT|20|17|Now as Jesus was going up to Jerusalem, he took the twelve disciples aside and said to them,
MATT|20|18|"We are going up to Jerusalem, and the Son of Man will be betrayed to the chief priests and the teachers of the law. They will condemn him to death
MATT|20|19|and will turn him over to the Gentiles to be mocked and flogged and crucified. On the third day he will be raised to life!"
MATT|20|20|Then the mother of Zebedee's sons came to Jesus with her sons and, kneeling down, asked a favor of him.
MATT|20|21|"What is it you want?" he asked. She said, "Grant that one of these two sons of mine may sit at your right and the other at your left in your kingdom."
MATT|20|22|"You don't know what you are asking," Jesus said to them. "Can you drink the cup I am going to drink?We can," they answered.
MATT|20|23|Jesus said to them, "You will indeed drink from my cup, but to sit at my right or left is not for me to grant. These places belong to those for whom they have been prepared by my Father."
MATT|20|24|When the ten heard about this, they were indignant with the two brothers.
MATT|20|25|Jesus called them together and said, "You know that the rulers of the Gentiles lord it over them, and their high officials exercise authority over them.
MATT|20|26|Not so with you. Instead, whoever wants to become great among you must be your servant,
MATT|20|27|and whoever wants to be first must be your slave--
MATT|20|28|just as the Son of Man did not come to be served, but to serve, and to give his life as a ransom for many."
MATT|20|29|As Jesus and his disciples were leaving Jericho, a large crowd followed him.
MATT|20|30|Two blind men were sitting by the roadside, and when they heard that Jesus was going by, they shouted, "Lord, Son of David, have mercy on us!"
MATT|20|31|The crowd rebuked them and told them to be quiet, but they shouted all the louder, "Lord, Son of David, have mercy on us!"
MATT|20|32|Jesus stopped and called them. "What do you want me to do for you?" he asked.
MATT|20|33|"Lord," they answered, "we want our sight."
MATT|20|34|Jesus had compassion on them and touched their eyes. Immediately they received their sight and followed him.
MATT|21|1|As they approached Jerusalem and came to Bethphage on the Mount of Olives, Jesus sent two disciples,
MATT|21|2|saying to them, "Go to the village ahead of you, and at once you will find a donkey tied there, with her colt by her. Untie them and bring them to me.
MATT|21|3|If anyone says anything to you, tell him that the Lord needs them, and he will send them right away."
MATT|21|4|This took place to fulfill what was spoken through the prophet:
MATT|21|5|"Say to the Daughter of Zion, 'See, your king comes to you, gentle and riding on a donkey, on a colt, the foal of a donkey.'"
MATT|21|6|The disciples went and did as Jesus had instructed them.
MATT|21|7|They brought the donkey and the colt, placed their cloaks on them, and Jesus sat on them.
MATT|21|8|A very large crowd spread their cloaks on the road, while others cut branches from the trees and spread them on the road.
MATT|21|9|The crowds that went ahead of him and those that followed shouted, "Hosanna to the Son of David!Blessed is he who comes in the name of the Lord!Hosanna in the highest!"
MATT|21|10|When Jesus entered Jerusalem, the whole city was stirred and asked, "Who is this?"
MATT|21|11|The crowds answered, "This is Jesus, the prophet from Nazareth in Galilee."
MATT|21|12|Jesus entered the temple area and drove out all who were buying and selling there. He overturned the tables of the money changers and the benches of those selling doves.
MATT|21|13|"It is written," he said to them, "'My house will be called a house of prayer,' but you are making it a 'den of robbers.'"
MATT|21|14|The blind and the lame came to him at the temple, and he healed them.
MATT|21|15|But when the chief priests and the teachers of the law saw the wonderful things he did and the children shouting in the temple area, "Hosanna to the Son of David," they were indignant.
MATT|21|16|"Do you hear what these children are saying?" they asked him. "Yes," replied Jesus, "have you never read, "'From the lips of children and infants you have ordained praise'?"
MATT|21|17|And he left them and went out of the city to Bethany, where he spent the night.
MATT|21|18|Early in the morning, as he was on his way back to the city, he was hungry.
MATT|21|19|Seeing a fig tree by the road, he went up to it but found nothing on it except leaves. Then he said to it, "May you never bear fruit again!" Immediately the tree withered.
MATT|21|20|When the disciples saw this, they were amazed. "How did the fig tree wither so quickly?" they asked.
MATT|21|21|Jesus replied, "I tell you the truth, if you have faith and do not doubt, not only can you do what was done to the fig tree, but also you can say to this mountain, 'Go, throw yourself into the sea,' and it will be done.
MATT|21|22|If you believe, you will receive whatever you ask for in prayer."
MATT|21|23|Jesus entered the temple courts, and, while he was teaching, the chief priests and the elders of the people came to him. "By what authority are you doing these things?" they asked. "And who gave you this authority?"
MATT|21|24|Jesus replied, "I will also ask you one question. If you answer me, I will tell you by what authority I am doing these things.
MATT|21|25|John's baptism--where did it come from? Was it from heaven, or from men?"
MATT|21|26|They discussed it among themselves and said, "If we say, 'From heaven,' he will ask, 'Then why didn't you believe him?' But if we say, 'From men'--we are afraid of the people, for they all hold that John was a prophet."
MATT|21|27|So they answered Jesus, "We don't know." Then he said, "Neither will I tell you by what authority I am doing these things.
MATT|21|28|"What do you think? There was a man who had two sons. He went to the first and said, 'Son, go and work today in the vineyard.'
MATT|21|29|"'I will not,' he answered, but later he changed his mind and went.
MATT|21|30|"Then the father went to the other son and said the same thing. He answered, 'I will, sir,' but he did not go.
MATT|21|31|"Which of the two did what his father wanted?The first," they answered.
MATT|21|32|Jesus said to them, "I tell you the truth, the tax collectors and the prostitutes are entering the kingdom of God ahead of you. For John came to you to show you the way of righteousness, and you did not believe him, but the tax collectors and the prostitutes did. And even after you saw this, you did not repent and believe him.
MATT|21|33|"Listen to another parable: There was a landowner who planted a vineyard. He put a wall around it, dug a winepress in it and built a watchtower. Then he rented the vineyard to some farmers and went away on a journey.
MATT|21|34|When the harvest time approached, he sent his servants to the tenants to collect his fruit.
MATT|21|35|"The tenants seized his servants; they beat one, killed another, and stoned a third.
MATT|21|36|Then he sent other servants to them, more than the first time, and the tenants treated them the same way.
MATT|21|37|Last of all, he sent his son to them. 'They will respect my son,' he said.
MATT|21|38|"But when the tenants saw the son, they said to each other, 'This is the heir. Come, let's kill him and take his inheritance.'
MATT|21|39|So they took him and threw him out of the vineyard and killed him.
MATT|21|40|"Therefore, when the owner of the vineyard comes, what will he do to those tenants?"
MATT|21|41|"He will bring those wretches to a wretched end," they replied, "and he will rent the vineyard to other tenants, who will give him his share of the crop at harvest time."
MATT|21|42|Jesus said to them, "Have you never read in the Scriptures: "'The stone the builders rejected has become the capstone; the Lord has done this, and it is marvelous in our eyes'?
MATT|21|43|"Therefore I tell you that the kingdom of God will be taken away from you and given to a people who will produce its fruit.
MATT|21|44|He who falls on this stone will be broken to pieces, but he on whom it falls will be crushed."
MATT|21|45|When the chief priests and the Pharisees heard Jesus' parables, they knew he was talking about them.
MATT|21|46|They looked for a way to arrest him, but they were afraid of the crowd because the people held that he was a prophet.
MATT|22|1|Jesus spoke to them again in parables, saying:
MATT|22|2|"The kingdom of heaven is like a king who prepared a wedding banquet for his son.
MATT|22|3|He sent his servants to those who had been invited to the banquet to tell them to come, but they refused to come.
MATT|22|4|"Then he sent some more servants and said, 'Tell those who have been invited that I have prepared my dinner: My oxen and fattened cattle have been butchered, and everything is ready. Come to the wedding banquet.'
MATT|22|5|"But they paid no attention and went off--one to his field, another to his business.
MATT|22|6|The rest seized his servants, mistreated them and killed them.
MATT|22|7|The king was enraged. He sent his army and destroyed those murderers and burned their city.
MATT|22|8|"Then he said to his servants, 'The wedding banquet is ready, but those I invited did not deserve to come.
MATT|22|9|Go to the street corners and invite to the banquet anyone you find.'
MATT|22|10|So the servants went out into the streets and gathered all the people they could find, both good and bad, and the wedding hall was filled with guests.
MATT|22|11|"But when the king came in to see the guests, he noticed a man there who was not wearing wedding clothes.
MATT|22|12|'Friend,' he asked, 'how did you get in here without wedding clothes?' The man was speechless.
MATT|22|13|"Then the king told the attendants, 'Tie him hand and foot, and throw him outside, into the darkness, where there will be weeping and gnashing of teeth.'
MATT|22|14|"For many are invited, but few are chosen."
MATT|22|15|Then the Pharisees went out and laid plans to trap him in his words.
MATT|22|16|They sent their disciples to him along with the Herodians. "Teacher," they said, "we know you are a man of integrity and that you teach the way of God in accordance with the truth. You aren't swayed by men, because you pay no attention to who they are.
MATT|22|17|Tell us then, what is your opinion? Is it right to pay taxes to Caesar or not?"
MATT|22|18|But Jesus, knowing their evil intent, said, "You hypocrites, why are you trying to trap me?
MATT|22|19|Show me the coin used for paying the tax." They brought him a denarius,
MATT|22|20|and he asked them, "Whose portrait is this? And whose inscription?"
MATT|22|21|"Caesar's," they replied. Then he said to them, "Give to Caesar what is Caesar's, and to God what is God's."
MATT|22|22|When they heard this, they were amazed. So they left him and went away.
MATT|22|23|That same day the Sadducees, who say there is no resurrection, came to him with a question.
MATT|22|24|"Teacher," they said, "Moses told us that if a man dies without having children, his brother must marry the widow and have children for him.
MATT|22|25|Now there were seven brothers among us. The first one married and died, and since he had no children, he left his wife to his brother.
MATT|22|26|The same thing happened to the second and third brother, right on down to the seventh.
MATT|22|27|Finally, the woman died.
MATT|22|28|Now then, at the resurrection, whose wife will she be of the seven, since all of them were married to her?"
MATT|22|29|Jesus replied, "You are in error because you do not know the Scriptures or the power of God.
MATT|22|30|At the resurrection people will neither marry nor be given in marriage; they will be like the angels in heaven.
MATT|22|31|But about the resurrection of the dead--have you not read what God said to you,
MATT|22|32|'I am the God of Abraham, the God of Isaac, and the God of Jacob'? He is not the God of the dead but of the living."
MATT|22|33|When the crowds heard this, they were astonished at his teaching.
MATT|22|34|Hearing that Jesus had silenced the Sadducees, the Pharisees got together.
MATT|22|35|One of them, an expert in the law, tested him with this question:
MATT|22|36|"Teacher, which is the greatest commandment in the Law?"
MATT|22|37|Jesus replied: "'Love the Lord your God with all your heart and with all your soul and with all your mind.'
MATT|22|38|This is the first and greatest commandment.
MATT|22|39|And the second is like it: 'Love your neighbor as yourself.'
MATT|22|40|All the Law and the Prophets hang on these two commandments."
MATT|22|41|While the Pharisees were gathered together, Jesus asked them,
MATT|22|42|"What do you think about the Christ? Whose son is he?The son of David," they replied.
MATT|22|43|He said to them, "How is it then that David, speaking by the Spirit, calls him 'Lord'? For he says,
MATT|22|44|"'The Lord said to my Lord: "Sit at my right hand until I put your enemies under your feet."'
MATT|22|45|If then David calls him 'Lord,' how can he be his son?"
MATT|22|46|No one could say a word in reply, and from that day on no one dared to ask him any more questions.
MATT|23|1|Then Jesus said to the crowds and to his disciples:
MATT|23|2|"The teachers of the law and the Pharisees sit in Moses' seat.
MATT|23|3|So you must obey them and do everything they tell you. But do not do what they do, for they do not practice what they preach.
MATT|23|4|They tie up heavy loads and put them on men's shoulders, but they themselves are not willing to lift a finger to move them.
MATT|23|5|"Everything they do is done for men to see: They make their phylacteries wide and the tassels on their garments long;
MATT|23|6|they love the place of honor at banquets and the most important seats in the synagogues;
MATT|23|7|they love to be greeted in the marketplaces and to have men call them 'Rabbi.'
MATT|23|8|"But you are not to be called 'Rabbi,' for you have only one Master and you are all brothers.
MATT|23|9|And do not call anyone on earth 'father,' for you have one Father, and he is in heaven.
MATT|23|10|Nor are you to be called 'teacher,' for you have one Teacher, the Christ.
MATT|23|11|The greatest among you will be your servant.
MATT|23|12|For whoever exalts himself will be humbled, and whoever humbles himself will be exalted.
MATT|23|13|"Woe to you, teachers of the law and Pharisees, you hypocrites! You shut the kingdom of heaven in men's faces. You yourselves do not enter, nor will you let those enter who are trying to.
MATT|23|14|See Footnote
MATT|23|15|"Woe to you, teachers of the law and Pharisees, you hypocrites! You travel over land and sea to win a single convert, and when he becomes one, you make him twice as much a son of hell as you are.
MATT|23|16|"Woe to you, blind guides! You say, 'If anyone swears by the temple, it means nothing; but if anyone swears by the gold of the temple, he is bound by his oath.'
MATT|23|17|You blind fools! Which is greater: the gold, or the temple that makes the gold sacred?
MATT|23|18|You also say, 'If anyone swears by the altar, it means nothing; but if anyone swears by the gift on it, he is bound by his oath.'
MATT|23|19|You blind men! Which is greater: the gift, or the altar that makes the gift sacred?
MATT|23|20|Therefore, he who swears by the altar swears by it and by everything on it.
MATT|23|21|And he who swears by the temple swears by it and by the one who dwells in it.
MATT|23|22|And he who swears by heaven swears by God's throne and by the one who sits on it.
MATT|23|23|"Woe to you, teachers of the law and Pharisees, you hypocrites! You give a tenth of your spices--mint, dill and cummin. But you have neglected the more important matters of the law--justice, mercy and faithfulness. You should have practiced the latter, without neglecting the former.
MATT|23|24|You blind guides! You strain out a gnat but swallow a camel.
MATT|23|25|"Woe to you, teachers of the law and Pharisees, you hypocrites! You clean the outside of the cup and dish, but inside they are full of greed and self-indulgence.
MATT|23|26|Blind Pharisee! First clean the inside of the cup and dish, and then the outside also will be clean.
MATT|23|27|"Woe to you, teachers of the law and Pharisees, you hypocrites! You are like whitewashed tombs, which look beautiful on the outside but on the inside are full of dead men's bones and everything unclean.
MATT|23|28|In the same way, on the outside you appear to people as righteous but on the inside you are full of hypocrisy and wickedness.
MATT|23|29|"Woe to you, teachers of the law and Pharisees, you hypocrites! You build tombs for the prophets and decorate the graves of the righteous.
MATT|23|30|And you say, 'If we had lived in the days of our forefathers, we would not have taken part with them in shedding the blood of the prophets.'
MATT|23|31|So you testify against yourselves that you are the descendants of those who murdered the prophets.
MATT|23|32|Fill up, then, the measure of the sin of your forefathers!
MATT|23|33|"You snakes! You brood of vipers! How will you escape being condemned to hell?
MATT|23|34|Therefore I am sending you prophets and wise men and teachers. Some of them you will kill and crucify; others you will flog in your synagogues and pursue from town to town.
MATT|23|35|And so upon you will come all the righteous blood that has been shed on earth, from the blood of righteous Abel to the blood of Zechariah son of Berekiah, whom you murdered between the temple and the altar.
MATT|23|36|I tell you the truth, all this will come upon this generation.
MATT|23|37|"O Jerusalem, Jerusalem, you who kill the prophets and stone those sent to you, how often I have longed to gather your children together, as a hen gathers her chicks under her wings, but you were not willing.
MATT|23|38|Look, your house is left to you desolate.
MATT|23|39|For I tell you, you will not see me again until you say, 'Blessed is he who comes in the name of the Lord.'"
MATT|24|1|Jesus left the temple and was walking away when his disciples came up to him to call his attention to its buildings.
MATT|24|2|"Do you see all these things?" he asked. "I tell you the truth, not one stone here will be left on another; every one will be thrown down."
MATT|24|3|As Jesus was sitting on the Mount of Olives, the disciples came to him privately. "Tell us," they said, "when will this happen, and what will be the sign of your coming and of the end of the age?"
MATT|24|4|Jesus answered: "Watch out that no one deceives you.
MATT|24|5|For many will come in my name, claiming, 'I am the Christ, 'and will deceive many.
MATT|24|6|You will hear of wars and rumors of wars, but see to it that you are not alarmed. Such things must happen, but the end is still to come.
MATT|24|7|Nation will rise against nation, and kingdom against kingdom. There will be famines and earthquakes in various places.
MATT|24|8|All these are the beginning of birth pains.
MATT|24|9|"Then you will be handed over to be persecuted and put to death, and you will be hated by all nations because of me.
MATT|24|10|At that time many will turn away from the faith and will betray and hate each other,
MATT|24|11|and many false prophets will appear and deceive many people.
MATT|24|12|Because of the increase of wickedness, the love of most will grow cold,
MATT|24|13|but he who stands firm to the end will be saved.
MATT|24|14|And this gospel of the kingdom will be preached in the whole world as a testimony to all nations, and then the end will come.
MATT|24|15|"So when you see standing in the holy place 'the abomination that causes desolation,' spoken of through the prophet Daniel--let the reader understand--
MATT|24|16|then let those who are in Judea flee to the mountains.
MATT|24|17|Let no one on the roof of his house go down to take anything out of the house.
MATT|24|18|Let no one in the field go back to get his cloak.
MATT|24|19|How dreadful it will be in those days for pregnant women and nursing mothers!
MATT|24|20|Pray that your flight will not take place in winter or on the Sabbath.
MATT|24|21|For then there will be great distress, unequaled from the beginning of the world until now--and never to be equaled again.
MATT|24|22|If those days had not been cut short, no one would survive, but for the sake of the elect those days will be shortened.
MATT|24|23|At that time if anyone says to you, 'Look, here is the Christ!' or, 'There he is!' do not believe it.
MATT|24|24|For false Christs and false prophets will appear and perform great signs and miracles to deceive even the elect--if that were possible.
MATT|24|25|See, I have told you ahead of time.
MATT|24|26|"So if anyone tells you, 'There he is, out in the desert,' do not go out; or, 'Here he is, in the inner rooms,' do not believe it.
MATT|24|27|For as lightning that comes from the east is visible even in the west, so will be the coming of the Son of Man.
MATT|24|28|Wherever there is a carcass, there the vultures will gather.
MATT|24|29|"Immediately after the distress of those days "'the sun will be darkened, and the moon will not give its light; the stars will fall from the sky, and the heavenly bodies will be shaken.'
MATT|24|30|"At that time the sign of the Son of Man will appear in the sky, and all the nations of the earth will mourn. They will see the Son of Man coming on the clouds of the sky, with power and great glory.
MATT|24|31|And he will send his angels with a loud trumpet call, and they will gather his elect from the four winds, from one end of the heavens to the other.
MATT|24|32|"Now learn this lesson from the fig tree: As soon as its twigs get tender and its leaves come out, you know that summer is near.
MATT|24|33|Even so, when you see all these things, you know that it is near, right at the door.
MATT|24|34|I tell you the truth, this generation will certainly not pass away until all these things have happened.
MATT|24|35|Heaven and earth will pass away, but my words will never pass away.
MATT|24|36|"No one knows about that day or hour, not even the angels in heaven, nor the Son, but only the Father.
MATT|24|37|As it was in the days of Noah, so it will be at the coming of the Son of Man.
MATT|24|38|For in the days before the flood, people were eating and drinking, marrying and giving in marriage, up to the day Noah entered the ark;
MATT|24|39|and they knew nothing about what would happen until the flood came and took them all away. That is how it will be at the coming of the Son of Man.
MATT|24|40|Two men will be in the field; one will be taken and the other left.
MATT|24|41|Two women will be grinding with a hand mill; one will be taken and the other left.
MATT|24|42|"Therefore keep watch, because you do not know on what day your Lord will come.
MATT|24|43|But understand this: If the owner of the house had known at what time of night the thief was coming, he would have kept watch and would not have let his house be broken into.
MATT|24|44|So you also must be ready, because the Son of Man will come at an hour when you do not expect him.
MATT|24|45|"Who then is the faithful and wise servant, whom the master has put in charge of the servants in his household to give them their food at the proper time?
MATT|24|46|It will be good for that servant whose master finds him doing so when he returns.
MATT|24|47|I tell you the truth, he will put him in charge of all his possessions.
MATT|24|48|But suppose that servant is wicked and says to himself, 'My master is staying away a long time,'
MATT|24|49|and he then begins to beat his fellow servants and to eat and drink with drunkards.
MATT|24|50|The master of that servant will come on a day when he does not expect him and at an hour he is not aware of.
MATT|24|51|He will cut him to pieces and assign him a place with the hypocrites, where there will be weeping and gnashing of teeth.
MATT|25|1|"At that time the kingdom of heaven will be like ten virgins who took their lamps and went out to meet the bridegroom.
MATT|25|2|Five of them were foolish and five were wise.
MATT|25|3|The foolish ones took their lamps but did not take any oil with them.
MATT|25|4|The wise, however, took oil in jars along with their lamps.
MATT|25|5|The bridegroom was a long time in coming, and they all became drowsy and fell asleep.
MATT|25|6|"At midnight the cry rang out: 'Here's the bridegroom! Come out to meet him!'
MATT|25|7|"Then all the virgins woke up and trimmed their lamps.
MATT|25|8|The foolish ones said to the wise, 'Give us some of your oil; our lamps are going out.'
MATT|25|9|"'No,' they replied, 'there may not be enough for both us and you. Instead, go to those who sell oil and buy some for yourselves.'
MATT|25|10|"But while they were on their way to buy the oil, the bridegroom arrived. The virgins who were ready went in with him to the wedding banquet. And the door was shut.
MATT|25|11|"Later the others also came. 'Sir! Sir!' they said. 'Open the door for us!'
MATT|25|12|"But he replied, 'I tell you the truth, I don't know you.'
MATT|25|13|"Therefore keep watch, because you do not know the day or the hour.
MATT|25|14|"Again, it will be like a man going on a journey, who called his servants and entrusted his property to them.
MATT|25|15|To one he gave five talents of money, to another two talents, and to another one talent, each according to his ability. Then he went on his journey.
MATT|25|16|The man who had received the five talents went at once and put his money to work and gained five more.
MATT|25|17|So also, the one with the two talents gained two more.
MATT|25|18|But the man who had received the one talent went off, dug a hole in the ground and hid his master's money.
MATT|25|19|"After a long time the master of those servants returned and settled accounts with them.
MATT|25|20|The man who had received the five talents brought the other five. 'Master,' he said, 'you entrusted me with five talents. See, I have gained five more.'
MATT|25|21|"His master replied, 'Well done, good and faithful servant! You have been faithful with a few things; I will put you in charge of many things. Come and share your master's happiness!'
MATT|25|22|"The man with the two talents also came. 'Master,' he said, 'you entrusted me with two talents; see, I have gained two more.'
MATT|25|23|"His master replied, 'Well done, good and faithful servant! You have been faithful with a few things; I will put you in charge of many things. Come and share your master's happiness!'
MATT|25|24|"Then the man who had received the one talent came. 'Master,' he said, 'I knew that you are a hard man, harvesting where you have not sown and gathering where you have not scattered seed.
MATT|25|25|So I was afraid and went out and hid your talent in the ground. See, here is what belongs to you.'
MATT|25|26|"His master replied, 'You wicked, lazy servant! So you knew that I harvest where I have not sown and gather where I have not scattered seed?
MATT|25|27|Well then, you should have put my money on deposit with the bankers, so that when I returned I would have received it back with interest.
MATT|25|28|"'Take the talent from him and give it to the one who has the ten talents.
MATT|25|29|For everyone who has will be given more, and he will have an abundance. Whoever does not have, even what he has will be taken from him.
MATT|25|30|And throw that worthless servant outside, into the darkness, where there will be weeping and gnashing of teeth.'
MATT|25|31|"When the Son of Man comes in his glory, and all the angels with him, he will sit on his throne in heavenly glory.
MATT|25|32|All the nations will be gathered before him, and he will separate the people one from another as a shepherd separates the sheep from the goats.
MATT|25|33|He will put the sheep on his right and the goats on his left.
MATT|25|34|"Then the King will say to those on his right, 'Come, you who are blessed by my Father; take your inheritance, the kingdom prepared for you since the creation of the world.
MATT|25|35|For I was hungry and you gave me something to eat, I was thirsty and you gave me something to drink, I was a stranger and you invited me in,
MATT|25|36|I needed clothes and you clothed me, I was sick and you looked after me, I was in prison and you came to visit me.'
MATT|25|37|"Then the righteous will answer him, 'Lord, when did we see you hungry and feed you, or thirsty and give you something to drink?
MATT|25|38|When did we see you a stranger and invite you in, or needing clothes and clothe you?
MATT|25|39|When did we see you sick or in prison and go to visit you?'
MATT|25|40|"The King will reply, 'I tell you the truth, whatever you did for one of the least of these brothers of mine, you did for me.'
MATT|25|41|"Then he will say to those on his left, 'Depart from me, you who are cursed, into the eternal fire prepared for the devil and his angels.
MATT|25|42|For I was hungry and you gave me nothing to eat, I was thirsty and you gave me nothing to drink,
MATT|25|43|I was a stranger and you did not invite me in, I needed clothes and you did not clothe me, I was sick and in prison and you did not look after me.'
MATT|25|44|"They also will answer, 'Lord, when did we see you hungry or thirsty or a stranger or needing clothes or sick or in prison, and did not help you?'
MATT|25|45|"He will reply, 'I tell you the truth, whatever you did not do for one of the least of these, you did not do for me.'
MATT|25|46|"Then they will go away to eternal punishment, but the righteous to eternal life."
MATT|26|1|When Jesus had finished saying all these things, he said to his disciples,
MATT|26|2|"As you know, the Passover is two days away--and the Son of Man will be handed over to be crucified."
MATT|26|3|Then the chief priests and the elders of the people assembled in the palace of the high priest, whose name was Caiaphas,
MATT|26|4|and they plotted to arrest Jesus in some sly way and kill him.
MATT|26|5|"But not during the Feast," they said, "or there may be a riot among the people."
MATT|26|6|While Jesus was in Bethany in the home of a man known as Simon the Leper,
MATT|26|7|a woman came to him with an alabaster jar of very expensive perfume, which she poured on his head as he was reclining at the table.
MATT|26|8|When the disciples saw this, they were indignant. "Why this waste?" they asked.
MATT|26|9|"This perfume could have been sold at a high price and the money given to the poor."
MATT|26|10|Aware of this, Jesus said to them, "Why are you bothering this woman? She has done a beautiful thing to me.
MATT|26|11|The poor you will always have with you, but you will not always have me.
MATT|26|12|When she poured this perfume on my body, she did it to prepare me for burial.
MATT|26|13|I tell you the truth, wherever this gospel is preached throughout the world, what she has done will also be told, in memory of her."
MATT|26|14|Then one of the Twelve--the one called Judas Iscariot--went to the chief priests
MATT|26|15|and asked, "What are you willing to give me if I hand him over to you?" So they counted out for him thirty silver coins.
MATT|26|16|From then on Judas watched for an opportunity to hand him over.
MATT|26|17|On the first day of the Feast of Unleavened Bread, the disciples came to Jesus and asked, "Where do you want us to make preparations for you to eat the Passover?"
MATT|26|18|He replied, "Go into the city to a certain man and tell him, 'The Teacher says: My appointed time is near. I am going to celebrate the Passover with my disciples at your house.'"
MATT|26|19|So the disciples did as Jesus had directed them and prepared the Passover.
MATT|26|20|When evening came, Jesus was reclining at the table with the Twelve.
MATT|26|21|And while they were eating, he said, "I tell you the truth, one of you will betray me."
MATT|26|22|They were very sad and began to say to him one after the other, "Surely not I, Lord?"
MATT|26|23|Jesus replied, "The one who has dipped his hand into the bowl with me will betray me.
MATT|26|24|The Son of Man will go just as it is written about him. But woe to that man who betrays the Son of Man! It would be better for him if he had not been born."
MATT|26|25|Then Judas, the one who would betray him, said, "Surely not I, Rabbi?" Jesus answered, "Yes, it is you."
MATT|26|26|While they were eating, Jesus took bread, gave thanks and broke it, and gave it to his disciples, saying, "Take and eat; this is my body."
MATT|26|27|Then he took the cup, gave thanks and offered it to them, saying, "Drink from it, all of you.
MATT|26|28|This is my blood of the covenant, which is poured out for many for the forgiveness of sins.
MATT|26|29|I tell you, I will not drink of this fruit of the vine from now on until that day when I drink it anew with you in my Father's kingdom."
MATT|26|30|When they had sung a hymn, they went out to the Mount of Olives.
MATT|26|31|Then Jesus told them, "This very night you will all fall away on account of me, for it is written: "'I will strike the shepherd, and the sheep of the flock will be scattered.'
MATT|26|32|But after I have risen, I will go ahead of you into Galilee."
MATT|26|33|Peter replied, "Even if all fall away on account of you, I never will."
MATT|26|34|"I tell you the truth," Jesus answered, "this very night, before the rooster crows, you will disown me three times."
MATT|26|35|But Peter declared, "Even if I have to die with you, I will never disown you." And all the other disciples said the same.
MATT|26|36|Then Jesus went with his disciples to a place called Gethsemane, and he said to them, "Sit here while I go over there and pray."
MATT|26|37|He took Peter and the two sons of Zebedee along with him, and he began to be sorrowful and troubled.
MATT|26|38|Then he said to them, "My soul is overwhelmed with sorrow to the point of death. Stay here and keep watch with me."
MATT|26|39|Going a little farther, he fell with his face to the ground and prayed, "My Father, if it is possible, may this cup be taken from me. Yet not as I will, but as you will."
MATT|26|40|Then he returned to his disciples and found them sleeping. "Could you men not keep watch with me for one hour?" he asked Peter.
MATT|26|41|"Watch and pray so that you will not fall into temptation. The spirit is willing, but the body is weak."
MATT|26|42|He went away a second time and prayed, "My Father, if it is not possible for this cup to be taken away unless I drink it, may your will be done."
MATT|26|43|When he came back, he again found them sleeping, because their eyes were heavy.
MATT|26|44|So he left them and went away once more and prayed the third time, saying the same thing.
MATT|26|45|Then he returned to the disciples and said to them, "Are you still sleeping and resting? Look, the hour is near, and the Son of Man is betrayed into the hands of sinners.
MATT|26|46|Rise, let us go! Here comes my betrayer!"
MATT|26|47|While he was still speaking, Judas, one of the Twelve, arrived. With him was a large crowd armed with swords and clubs, sent from the chief priests and the elders of the people.
MATT|26|48|Now the betrayer had arranged a signal with them: "The one I kiss is the man; arrest him."
MATT|26|49|Going at once to Jesus, Judas said, "Greetings, Rabbi!" and kissed him.
MATT|26|50|Jesus replied, "Friend, do what you came for."
MATT|26|51|Then the men stepped forward, seized Jesus and arrested him. With that, one of Jesus' companions reached for his sword, drew it out and struck the servant of the high priest, cutting off his ear.
MATT|26|52|"Put your sword back in its place," Jesus said to him, "for all who draw the sword will die by the sword.
MATT|26|53|Do you think I cannot call on my Father, and he will at once put at my disposal more than twelve legions of angels?
MATT|26|54|But how then would the Scriptures be fulfilled that say it must happen in this way?"
MATT|26|55|At that time Jesus said to the crowd, "Am I leading a rebellion, that you have come out with swords and clubs to capture me? Every day I sat in the temple courts teaching, and you did not arrest me.
MATT|26|56|But this has all taken place that the writings of the prophets might be fulfilled." Then all the disciples deserted him and fled.
MATT|26|57|Those who had arrested Jesus took him to Caiaphas, the high priest, where the teachers of the law and the elders had assembled.
MATT|26|58|But Peter followed him at a distance, right up to the courtyard of the high priest. He entered and sat down with the guards to see the outcome.
MATT|26|59|The chief priests and the whole Sanhedrin were looking for false evidence against Jesus so that they could put him to death.
MATT|26|60|But they did not find any, though many false witnesses came forward.
MATT|26|61|Finally two came forward and declared, "This fellow said, 'I am able to destroy the temple of God and rebuild it in three days.'"
MATT|26|62|Then the high priest stood up and said to Jesus, "Are you not going to answer? What is this testimony that these men are bringing against you?"
MATT|26|63|But Jesus remained silent. The high priest said to him, "I charge you under oath by the living God: Tell us if you are the Christ, the Son of God."
MATT|26|64|"Yes, it is as you say," Jesus replied. "But I say to all of you: In the future you will see the Son of Man sitting at the right hand of the Mighty One and coming on the clouds of heaven."
MATT|26|65|Then the high priest tore his clothes and said, "He has spoken blasphemy! Why do we need any more witnesses? Look, now you have heard the blasphemy.
MATT|26|66|What do you think?He is worthy of death," they answered.
MATT|26|67|Then they spit in his face and struck him with their fists. Others slapped him
MATT|26|68|and said, "Prophesy to us, Christ. Who hit you?"
MATT|26|69|Now Peter was sitting out in the courtyard, and a servant girl came to him. "You also were with Jesus of Galilee," she said.
MATT|26|70|But he denied it before them all. "I don't know what you're talking about," he said.
MATT|26|71|Then he went out to the gateway, where another girl saw him and said to the people there, "This fellow was with Jesus of Nazareth."
MATT|26|72|He denied it again, with an oath: "I don't know the man!"
MATT|26|73|After a little while, those standing there went up to Peter and said, "Surely you are one of them, for your accent gives you away."
MATT|26|74|Then he began to call down curses on himself and he swore to them, "I don't know the man!"
MATT|26|75|Immediately a rooster crowed. Then Peter remembered the word Jesus had spoken: "Before the rooster crows, you will disown me three times." And he went outside and wept bitterly.
MATT|27|1|Early in the morning, all the chief priests and the elders of the people came to the decision to put Jesus to death.
MATT|27|2|They bound him, led him away and handed him over to Pilate, the governor.
MATT|27|3|When Judas, who had betrayed him, saw that Jesus was condemned, he was seized with remorse and returned the thirty silver coins to the chief priests and the elders.
MATT|27|4|"I have sinned," he said, "for I have betrayed innocent blood.What is that to us?" they replied. "That's your responsibility."
MATT|27|5|So Judas threw the money into the temple and left. Then he went away and hanged himself.
MATT|27|6|The chief priests picked up the coins and said, "It is against the law to put this into the treasury, since it is blood money."
MATT|27|7|So they decided to use the money to buy the potter's field as a burial place for foreigners.
MATT|27|8|That is why it has been called the Field of Blood to this day.
MATT|27|9|Then what was spoken by Jeremiah the prophet was fulfilled: "They took the thirty silver coins, the price set on him by the people of Israel,
MATT|27|10|and they used them to buy the potter's field, as the Lord commanded me."
MATT|27|11|Meanwhile Jesus stood before the governor, and the governor asked him, "Are you the king of the Jews?Yes, it is as you say," Jesus replied.
MATT|27|12|When he was accused by the chief priests and the elders, he gave no answer.
MATT|27|13|Then Pilate asked him, "Don't you hear the testimony they are bringing against you?"
MATT|27|14|But Jesus made no reply, not even to a single charge--to the great amazement of the governor.
MATT|27|15|Now it was the governor's custom at the Feast to release a prisoner chosen by the crowd.
MATT|27|16|At that time they had a notorious prisoner, called Barabbas.
MATT|27|17|So when the crowd had gathered, Pilate asked them, "Which one do you want me to release to you: Barabbas, or Jesus who is called Christ?"
MATT|27|18|For he knew it was out of envy that they had handed Jesus over to him.
MATT|27|19|While Pilate was sitting on the judge's seat, his wife sent him this message: "Don't have anything to do with that innocent man, for I have suffered a great deal today in a dream because of him."
MATT|27|20|But the chief priests and the elders persuaded the crowd to ask for Barabbas and to have Jesus executed.
MATT|27|21|"Which of the two do you want me to release to you?" asked the governor. "Barabbas," they answered.
MATT|27|22|"What shall I do, then, with Jesus who is called Christ?" Pilate asked. They all answered, "Crucify him!"
MATT|27|23|"Why? What crime has he committed?" asked Pilate. But they shouted all the louder, "Crucify him!"
MATT|27|24|When Pilate saw that he was getting nowhere, but that instead an uproar was starting, he took water and washed his hands in front of the crowd. "I am innocent of this man's blood," he said. "It is your responsibility!"
MATT|27|25|All the people answered, "Let his blood be on us and on our children!"
MATT|27|26|Then he released Barabbas to them. But he had Jesus flogged, and handed him over to be crucified.
MATT|27|27|Then the governor's soldiers took Jesus into the Praetorium and gathered the whole company of soldiers around him.
MATT|27|28|They stripped him and put a scarlet robe on him,
MATT|27|29|and then twisted together a crown of thorns and set it on his head. They put a staff in his right hand and knelt in front of him and mocked him. "Hail, king of the Jews!" they said.
MATT|27|30|They spit on him, and took the staff and struck him on the head again and again.
MATT|27|31|After they had mocked him, they took off the robe and put his own clothes on him. Then they led him away to crucify him.
MATT|27|32|As they were going out, they met a man from Cyrene, named Simon, and they forced him to carry the cross.
MATT|27|33|They came to a place called Golgotha (which means The Place of the Skull).
MATT|27|34|There they offered Jesus wine to drink, mixed with gall; but after tasting it, he refused to drink it.
MATT|27|35|When they had crucified him, they divided up his clothes by casting lots.
MATT|27|36|And sitting down, they kept watch over him there.
MATT|27|37|Above his head they placed the written charge against him: THIS IS JESUS, THE KING OF THE JEWS.
MATT|27|38|Two robbers were crucified with him, one on his right and one on his left.
MATT|27|39|Those who passed by hurled insults at him, shaking their heads
MATT|27|40|and saying, "You who are going to destroy the temple and build it in three days, save yourself! Come down from the cross, if you are the Son of God!"
MATT|27|41|In the same way the chief priests, the teachers of the law and the elders mocked him.
MATT|27|42|"He saved others," they said, "but he can't save himself! He's the King of Israel! Let him come down now from the cross, and we will believe in him.
MATT|27|43|He trusts in God. Let God rescue him now if he wants him, for he said, 'I am the Son of God.'"
MATT|27|44|In the same way the robbers who were crucified with him also heaped insults on him.
MATT|27|45|From the sixth hour until the ninth hour darkness came over all the land.
MATT|27|46|About the ninth hour Jesus cried out in a loud voice, "Eloi, Eloi, lama sabachthani?"--which means, "My God, my God, why have you forsaken me?"
MATT|27|47|When some of those standing there heard this, they said, "He's calling Elijah."
MATT|27|48|Immediately one of them ran and got a sponge. He filled it with wine vinegar, put it on a stick, and offered it to Jesus to drink.
MATT|27|49|The rest said, "Now leave him alone. Let's see if Elijah comes to save him."
MATT|27|50|And when Jesus had cried out again in a loud voice, he gave up his spirit.
MATT|27|51|At that moment the curtain of the temple was torn in two from top to bottom. The earth shook and the rocks split.
MATT|27|52|The tombs broke open and the bodies of many holy people who had died were raised to life.
MATT|27|53|They came out of the tombs, and after Jesus' resurrection they went into the holy city and appeared to many people.
MATT|27|54|When the centurion and those with him who were guarding Jesus saw the earthquake and all that had happened, they were terrified, and exclaimed, "Surely he was the Son of God!"
MATT|27|55|Many women were there, watching from a distance. They had followed Jesus from Galilee to care for his needs.
MATT|27|56|Among them were Mary Magdalene, Mary the mother of James and Joses, and the mother of Zebedee's sons.
MATT|27|57|As evening approached, there came a rich man from Arimathea, named Joseph, who had himself become a disciple of Jesus.
MATT|27|58|Going to Pilate, he asked for Jesus' body, and Pilate ordered that it be given to him.
MATT|27|59|Joseph took the body, wrapped it in a clean linen cloth,
MATT|27|60|and placed it in his own new tomb that he had cut out of the rock. He rolled a big stone in front of the entrance to the tomb and went away.
MATT|27|61|Mary Magdalene and the other Mary were sitting there opposite the tomb.
MATT|27|62|The next day, the one after Preparation Day, the chief priests and the Pharisees went to Pilate.
MATT|27|63|"Sir," they said, "we remember that while he was still alive that deceiver said, 'After three days I will rise again.'
MATT|27|64|So give the order for the tomb to be made secure until the third day. Otherwise, his disciples may come and steal the body and tell the people that he has been raised from the dead. This last deception will be worse than the first."
MATT|27|65|"Take a guard," Pilate answered. "Go, make the tomb as secure as you know how."
MATT|27|66|So they went and made the tomb secure by putting a seal on the stone and posting the guard.
MATT|28|1|After the Sabbath, at dawn on the first day of the week, Mary Magdalene and the other Mary went to look at the tomb.
MATT|28|2|There was a violent earthquake, for an angel of the Lord came down from heaven and, going to the tomb, rolled back the stone and sat on it.
MATT|28|3|His appearance was like lightning, and his clothes were white as snow.
MATT|28|4|The guards were so afraid of him that they shook and became like dead men.
MATT|28|5|The angel said to the women, "Do not be afraid, for I know that you are looking for Jesus, who was crucified.
MATT|28|6|He is not here; he has risen, just as he said. Come and see the place where he lay.
MATT|28|7|Then go quickly and tell his disciples: 'He has risen from the dead and is going ahead of you into Galilee. There you will see him.' Now I have told you."
MATT|28|8|So the women hurried away from the tomb, afraid yet filled with joy, and ran to tell his disciples.
MATT|28|9|Suddenly Jesus met them. "Greetings," he said. They came to him, clasped his feet and worshiped him.
MATT|28|10|Then Jesus said to them, "Do not be afraid. Go and tell my brothers to go to Galilee; there they will see me."
MATT|28|11|While the women were on their way, some of the guards went into the city and reported to the chief priests everything that had happened.
MATT|28|12|When the chief priests had met with the elders and devised a plan, they gave the soldiers a large sum of money,
MATT|28|13|telling them, "You are to say, 'His disciples came during the night and stole him away while we were asleep.'
MATT|28|14|If this report gets to the governor, we will satisfy him and keep you out of trouble."
MATT|28|15|So the soldiers took the money and did as they were instructed. And this story has been widely circulated among the Jews to this very day.
MATT|28|16|Then the eleven disciples went to Galilee, to the mountain where Jesus had told them to go.
MATT|28|17|When they saw him, they worshiped him; but some doubted.
MATT|28|18|Then Jesus came to them and said, "All authority in heaven and on earth has been given to me.
MATT|28|19|Therefore go and make disciples of all nations, baptizing them in the name of the Father and of the Son and of the Holy Spirit,
MATT|28|20|and teaching them to obey everything I have commanded you. And surely I am with you always, to the very end of the age."
