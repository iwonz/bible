JOEL|1|1|Verbum Domini, quod factum est ad loel filium Phatuel.
JOEL|1|2|Audite hoc, senes,et auribus percipite, omnes habitatores terrae,si factum est istud in diebus vestrisaut in diebus patrum vestrorum.
JOEL|1|3|Super hoc filiis vestris narrate,et filii vestri filiis suis,et filii eorum generationi alterae.
JOEL|1|4|Residuum erucae comedit locusta,et residuum locustae comedit bruchus,et residuum bruchi comedit gryllus.
JOEL|1|5|Expergiscimini, ebrii, et flete,et ululate, omnes, qui bibitis vinum,propter mustum,quoniam periit ab ore vestro.
JOEL|1|6|Gens enim ascendit super terram meamfortis et innumerabilis;dentes eius ut dentes leonis,et molares leaenae sunt ei.
JOEL|1|7|Posuit vineam meam in desertumet ficum meam in lignum confractum;nudans spoliavit eam et proiecit,albi facti sunt rami eius.
JOEL|1|8|Plange, quasi virgo accincta saccosuper virum pubertatis suae.
JOEL|1|9|Periit oblatio et libatiode domo Domini;luxerunt sacerdotesministri Domini.
JOEL|1|10|Depopulata est regio;luxit humus,quoniam devastatum est triticum,defecit mustum,elanguit oleum.
JOEL|1|11|Confundemini, agricolae,ululate, vinitores,super frumento et hordeo,quia periit messis agri.
JOEL|1|12|Vinea exaruit,et ficus elanguit,malogranatum et palma et malumet omnia ligna agri aruerunt,quia evanuit gaudiuma filiis hominum.
JOEL|1|13|Accingite vos et plangite, sacerdotes;ululate, ministri altaris.Ingredimini, cubate in sacco,ministri Dei mei,quoniam interiit de domo Dei vestrioblatio et libatio.
JOEL|1|14|Sanctificate ieiunium,vocate coetum,congregate senes,omnes habitatores terraein domum Dei vestri,et clamate ad Dominum:
JOEL|1|15|" Heu diei!Quia prope est dies Domini,et quasi vastitas a potente veniet.
JOEL|1|16|Numquid non coram oculis vestrisalimenta perierunt,de domo Dei nostrilaetitia et exsultatio?".
JOEL|1|17|Computruerunt seminasubtus glebas suas,demolita sunt horrea,dissipatae sunt apothecae,eo quod exaruit triticum.
JOEL|1|18|Quid ingemuit animal,perterrita sunt armenta boum,quia non est pascua eis?Sed et greges pecorum disperierunt.
JOEL|1|19|Ad te, Domine, clamo,quia ignis comeditpascua deserti,et flamma succenditomnia ligna agri.
JOEL|1|20|Sed et bestiae agrisuspirant ad te,quoniam exsiccati sunt fontes aquarum,et ignis devoravitpascua deserti.
JOEL|2|1|Canite tuba in Sion,ululate in monte sancto meo;conturbentur omnes habitatores terrae,quia venit dies Domini,quia prope est.
JOEL|2|2|Dies tenebrarum et caliginis,dies nubis et turbinis;quasi aurora expansa super montespopulus multus et fortis:similis ei non fuit a principio,et post eum non eritusque in annos generationis et generationis.
JOEL|2|3|Ante faciem eius ignis vorat,et post eum exurit flamma.Quasi hortus Eden terra coram eo,et post eum solitudo deserti;neque est quod effugiat eum.
JOEL|2|4|Quasi aspectus equorum aspectus eorum,et quasi equites sic current.
JOEL|2|5|Sicut sonitus quadrigarumsuper capita montium exsiliunt,sicut sonitus flammae ignisdevorantis stipulam,velut populus fortispraeparatus ad proelium.
JOEL|2|6|A facie eius cruciabuntur populi,omnes vultus candentes.
JOEL|2|7|Sicut fortes currunt,quasi viri bellatores ascendunt murum;unusquisque in viis suis graditur,et non declinant a semitis suis.
JOEL|2|8|Unusquisque fratrem suum non coarctat,singuli in calle suo ambulant,per media tela prorumpuntsine intermissione.
JOEL|2|9|Urbem ingrediuntur,in murum discurrunt,domos conscendunt,per fenestras intrant quasi fur.
JOEL|2|10|A facie eius contremuit terra,moti sunt caeli,sol et luna obtenebrati sunt,et stellae retraxerunt splendorem suum.
JOEL|2|11|Et Dominus dedit vocem suam ante faciem exercitus sui,quia multa sunt nimis castra eius,quia fortia et facientia verbum eius;magnus enim dies Dominiet terribilis valde, et quis sustinebit eum?
JOEL|2|12|" Nunc ergo,dicit Dominus,convertimini ad me in toto corde vestro,in ieiunio et in fletu et in planctu;
JOEL|2|13|et scindite corda vestra et non vestimenta vestra,et convertimini ad Dominum Deum vestrum,quia benignus et misericors est,patiens et multae misericordiaeet placabilis super malitia ".
JOEL|2|14|Quis scit, si convertatur et ignoscatet relinquat post se benedictionem,oblationem et libationemDomino Deo vestro?
JOEL|2|15|Canite tuba in Sion,sanctificate ieiunium, vocate coetum;congregate populum, sanctificate conventum,coadunate senes,
JOEL|2|16|congregate parvulos et sugentes ubera,egrediatur sponsus de cubili suo,et sponsa de thalamo suo.
JOEL|2|17|Inter vestibulum et altare plorentsacerdotes ministri Dominiet dicant: "Parce, Domine, populo tuoet ne des hereditatem tuam in opprobrium,ut dominentur eis nationes ".Quare dicent in populis: Ubi est Deus eorum "?
JOEL|2|18|Zelatus est Dominus terram suamet pepercit populo suo.
JOEL|2|19|Et respondit Dominus et dixit populo suo: Ecce ego mittam vobisfrumentum et vinum et oleum,et replebimini eis;et non dabo vos ultraopprobrium in gentibus.
JOEL|2|20|Et eum, qui ab aquilone est,procul faciam a vobiset expellam eum in terraminviam et desertam:facies eius contra mare orientale,et extremum eius ad mare occidentale;et ascendet foetor eius,et ascendet putredo eius,quia magna operatus est.
JOEL|2|21|Noli timere, terra;exsulta et laetare,quoniam magna Dominus operatus est.
JOEL|2|22|Nolite timere, animalia regionis,quia germinaverunt pascua deserti,quia lignum attulit fructum suum,ficus et vinea dederunt divitias suas.
JOEL|2|23|Et, filii Sion, exsultateet laetamini in Domino Deo vestro,quia dedit vobispluviam iustitiaeet descendere fecit ad vosimbrem matutinum et serotinum sicut prius.
JOEL|2|24|Et implebuntur areae frumento,et redundabunt torculariavino et oleo;
JOEL|2|25|et reddam vobis annos,quos comedit locusta, bruchuset gryllus et eruca,exercitus meus magnus,quem misi in vos.
JOEL|2|26|Et comedetis vescentes et saturabiminiet laudabitis nomen Domini Dei vestri,qui mirabilia fecit vobiscum;et non confundetur populus meus in sempiternum.
JOEL|2|27|Et scietis quia in medio Israel ego sum,et ego Dominus Deus vester,et non est amplius;et non confundetur populus meus in aeternum ".
JOEL|3|1|Et erit post haec:effundam spiritum meum super omnem carnem,et prophetabunt filii vestri et filiae vestrae,senes vestri somnia somniabunt,et iuvenes vestri visiones videbunt;
JOEL|3|2|sed et super servos meos et ancillasin diebus illis effundam spiritum meum.
JOEL|3|3|Et dabo prodigia in caelo et in terra,sanguinem et ignem et columnas fumi;
JOEL|3|4|sol convertetur in tenebras,et luna in sanguinem,antequam veniat dies Dominimagnus et horribilis.
JOEL|3|5|Et erit:omnis, qui invocaverit nomen Domini, salvus erit,quia in monte Sion et in Ierusalemerit salvatio, sicut dixit Dominus,et in residuis, quos Dominus vocaverit.
JOEL|4|1|Quia ecce in diebus illiset in tempore illo,cum convertero sortemIudae et Ierusalem,
JOEL|4|2|congregabo omnes genteset deducam eas in vallem Iosaphatet disceptabo cum eis ibisuper populo meo et hereditate mea Israel,quos disperserunt in nationibus,et terram meam diviserunt.
JOEL|4|3|Et super populum meum miserunt sortem;et dederunt puerum pro meretriceet puellam vendiderunt pro vino, ut biberent.
JOEL|4|4|Verum quid vobis et mihi, Tyrus et Sidon et omnes termini Philisthaeae? Numquid ultionem vos reddetis mihi? Et si ulciscimini vos contra me, cito velociter reddam ultionem vestram super caput vestrum.
JOEL|4|5|Argentum enim meum et aurum tulistis et pretiosa bona mea intulistis in delubra vestra.
JOEL|4|6|Et filios Iudae et filios Ierusalem vendidistis filiis Graecorum, ut longe faceretis eos de finibus suis.
JOEL|4|7|Ecce ego suscitabo eos de loco, in quo vendidistis eos, et reddam ultionem vestram in caput vestrum.
JOEL|4|8|Et vendam filios vestros et filias vestras in manibus filiorum Iudae; et venumdabunt eos Sabaeis, genti longinquae, quia Dominus locutus est.
JOEL|4|9|Clamate hoc in gentibus,sanctificate bellum,suscitate robustos;accedant, ascendantomnes viri bellatores.
JOEL|4|10|Concidite vomeres vestros in gladioset falces vestras in lanceas;infirmus dicat: Fortis ego sum ".
JOEL|4|11|Erumpite et venite,omnes gentes de circuitu,et congregamini ibi!Deduc, Domine, robustos tuos!
JOEL|4|12|Consurgant et ascendant gentesin vallem Iosaphat,quia ibi sedebo, ut iudicemomnes gentes in circuitu.
JOEL|4|13|Mittite falces,quoniam maturavit messis;venite et premite,quia plenum est torcular:exuberant torcularia,quia magna est malitia eorum.
JOEL|4|14|Populi, populiin valle Decisionis,quia iuxta est dies Dominiin valle Decisionis.
JOEL|4|15|Sol et luna obtenebrati sunt,et stellae retraxerunt splendorem suum.
JOEL|4|16|Et Dominus de Sion rugietet de Ierusalem dabit vocem suam;et movebuntur caeli et terra,et Dominus refugium populo suoet fortitudo filiis Israel.
JOEL|4|17|Et scietis quia ego Dominus Deus vesterhabitans in Sion monte sancto meo;et erit Ierusalem locus sanctus,et alieni non transibunt per eam amplius.
JOEL|4|18|Et erit in die illa:stillabunt montes mustum,et colles fluent lacte;et per omnes rivos Iudae ibunt aquae,et fons de domo Domini egredieturet irrigabit torrentem Settim.
JOEL|4|19|Aegyptus in desolationem erit,et Idumaea in desertum desolationis,pro eo quod inique egerint in filios Iudaeet effuderint sanguinem innocentem in terra eorum.
JOEL|4|20|Et Iuda in aeternum habitabitur,et Ierusalem in generationem et generationem;
JOEL|4|21|et vindicabo sanguinem eorum, quem non relinquam impunitum;et Dominus commoratur in Sion.
