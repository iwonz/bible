3JOHN|1|1|Старець улюбленому Гаєві, якого я направду люблю.
3JOHN|1|2|Улюблений, я молюся, щоб добре велося в усьому тобі, і щоб був ти здоровий, як добре ведеться душі твоїй.
3JOHN|1|3|Бо я дуже зрадів, як прийшли були браття, і засвідчили правду твою, як ти живеш у правді.
3JOHN|1|4|Я не маю більшої радости від цієї, щоб чути, що діти мої живуть у правді.
3JOHN|1|5|Улюблений, вірно ти чиниш, як що робиш для братті та для чужинців,
3JOHN|1|6|вони про любов твою свідчили Церкві; добре ти зробиш, як їх випровадиш, як достойно для Бога,
3JOHN|1|7|бо вийшли вони ради Ймення Його, нічого не взявши від поган.
3JOHN|1|8|Отож, ми повинні приймати таких, щоб бути співробітниками правді.
3JOHN|1|9|Я до Церкви писав був, але Діотреф, що любить бути першим у них, нас не приймає.
3JOHN|1|10|Тому то, коли я прийду, то згадаю про вчинки його, що їх робить, словами лихими обмовляючи нас. І він тим не задовольнюється, а й сам не приймає братів, і тим, що бажають приймати, боронить, і вигонить із Церкви.
3JOHN|1|11|Улюблений, не робися подібним до лихого, а до доброго: доброчинець від Бога, а злочинець Бога не бачив.
3JOHN|1|12|Про Димитрія свідчили всі й сама правда. І свідчимо й ми, а ви знаєте, що свідчення наше правдиве.
3JOHN|1|13|Багато хотів я писати, та не хочу писати до тебе чорнилом та очеретинкою,
3JOHN|1|14|але маю надію побачити тебе незабаром, і говорити устами до уст. (1-15) Мир тобі! Друзі вітають тебе. Привітай друзів пойменно! Амінь.
