2JOHN|1|1|Старець вибраній пані та дітям її, яких я поправді люблю, і не тільки я, але й усі, хто правду пізнав,
2JOHN|1|2|за правду, що в нас пробуває й повік буде з нами:
2JOHN|1|3|нехай буде з вами благодать, милість, мир від Бога Отця та Ісуса Христа, Сина Отцевого, у правді та в любові!
2JOHN|1|4|Я дуже зрадів, що між дітьми твоїми знайшов таких, що ходять у правді, як заповідь ми прийняли від Отця.
2JOHN|1|5|І тепер я благаю тебе, пані, не так, ніби пишу тобі нову заповідь, але ту, яку маємо від початку, щоб ми любили один одного!
2JOHN|1|6|А любов ця щоб ми жили згідно з Його заповідями. Це та заповідь, яку ви чули від початку, щоб ви згідно з нею жили.
2JOHN|1|7|Бо в світ увійшло багато обманців, які не визнають Ісуса Христа, що прийшов був у тілі. Такий то обманець та антихрист!
2JOHN|1|8|Пильнуйте себе, щоб ви не згубили того, над чим працювали, але щоб прийняли повну нагороду.
2JOHN|1|9|Кожен, хто робить переступ та не пробуває в науці Христовій, той Бога не має. А хто пробуває в науці Його, той має і Отця, і Сина.
2JOHN|1|10|Коли хто приходить до вас, але не приносить науки цієї, не приймайте до дому його, і не вітайте його!
2JOHN|1|11|Хто бо вітає його, той участь бере в лихих учинках його.
2JOHN|1|12|Багато я мав написати до вас, але не схотів на папері й чорнилом. Та маю надію прибути до вас, і говорити устами до уст, щоб повна була ваша радість!
2JOHN|1|13|Вітають тебе діти вибраної сестри твоєї. Амінь.
