HAG|1|1|In the second year of King Darius, on the first day of the sixth month, the word of the LORD came through the prophet Haggai to Zerubbabel son of Shealtiel, governor of Judah, and to Joshua son of Jehozadak, the high priest:
HAG|1|2|This is what the LORD Almighty says: "These people say, 'The time has not yet come for the LORD's house to be built.'"
HAG|1|3|Then the word of the LORD came through the prophet Haggai:
HAG|1|4|"Is it a time for you yourselves to be living in your paneled houses, while this house remains a ruin?"
HAG|1|5|Now this is what the LORD Almighty says: "Give careful thought to your ways.
HAG|1|6|You have planted much, but have harvested little. You eat, but never have enough. You drink, but never have your fill. You put on clothes, but are not warm. You earn wages, only to put them in a purse with holes in it."
HAG|1|7|This is what the LORD Almighty says: "Give careful thought to your ways.
HAG|1|8|Go up into the mountains and bring down timber and build the house, so that I may take pleasure in it and be honored," says the LORD.
HAG|1|9|"You expected much, but see, it turned out to be little. What you brought home, I blew away. Why?" declares the LORD Almighty. "Because of my house, which remains a ruin, while each of you is busy with his own house.
HAG|1|10|Therefore, because of you the heavens have withheld their dew and the earth its crops.
HAG|1|11|I called for a drought on the fields and the mountains, on the grain, the new wine, the oil and whatever the ground produces, on men and cattle, and on the labor of your hands."
HAG|1|12|Then Zerubbabel son of Shealtiel, Joshua son of Jehozadak, the high priest, and the whole remnant of the people obeyed the voice of the LORD their God and the message of the prophet Haggai, because the LORD their God had sent him. And the people feared the LORD.
HAG|1|13|Then Haggai, the LORD's messenger, gave this message of the LORD to the people: "I am with you," declares the LORD.
HAG|1|14|So the LORD stirred up the spirit of Zerubbabel son of Shealtiel, governor of Judah, and the spirit of Joshua son of Jehozadak, the high priest, and the spirit of the whole remnant of the people. They came and began to work on the house of the LORD Almighty, their God,
HAG|1|15|on the twenty-fourth day of the sixth month in the second year of King Darius.
HAG|2|1|On the twenty-first day of the seventh month, the word of the LORD came through the prophet Haggai:
HAG|2|2|"Speak to Zerubbabel son of Shealtiel, governor of Judah, to Joshua son of Jehozadak, the high priest, and to the remnant of the people. Ask them,
HAG|2|3|'Who of you is left who saw this house in its former glory? How does it look to you now? Does it not seem to you like nothing?
HAG|2|4|But now be strong, O Zerubbabel,' declares the LORD. 'Be strong, O Joshua son of Jehozadak, the high priest. Be strong, all you people of the land,' declares the LORD, 'and work. For I am with you,' declares the LORD Almighty.
HAG|2|5|'This is what I covenanted with you when you came out of Egypt. And my Spirit remains among you. Do not fear.'
HAG|2|6|"This is what the LORD Almighty says: 'In a little while I will once more shake the heavens and the earth, the sea and the dry land.
HAG|2|7|I will shake all nations, and the desired of all nations will come, and I will fill this house with glory,' says the LORD Almighty.
HAG|2|8|'The silver is mine and the gold is mine,' declares the LORD Almighty.
HAG|2|9|'The glory of this present house will be greater than the glory of the former house,' says the LORD Almighty. 'And in this place I will grant peace,' declares the LORD Almighty."
HAG|2|10|On the twenty-fourth day of the ninth month, in the second year of Darius, the word of the LORD came to the prophet Haggai:
HAG|2|11|"This is what the LORD Almighty says: 'Ask the priests what the law says:
HAG|2|12|If a person carries consecrated meat in the fold of his garment, and that fold touches some bread or stew, some wine, oil or other food, does it become consecrated?'" The priests answered, "No."
HAG|2|13|Then Haggai said, "If a person defiled by contact with a dead body touches one of these things, does it become defiled?Yes," the priests replied, "it becomes defiled."
HAG|2|14|Then Haggai said, "'So it is with this people and this nation in my sight,' declares the LORD. 'Whatever they do and whatever they offer there is defiled.
HAG|2|15|"'Now give careful thought to this from this day on -consider how things were before one stone was laid on another in the LORD's temple.
HAG|2|16|When anyone came to a heap of twenty measures, there were only ten. When anyone went to a wine vat to draw fifty measures, there were only twenty.
HAG|2|17|I struck all the work of your hands with blight, mildew and hail, yet you did not turn to me,' declares the LORD.
HAG|2|18|'From this day on, from this twenty-fourth day of the ninth month, give careful thought to the day when the foundation of the LORD's temple was laid. Give careful thought:
HAG|2|19|Is there yet any seed left in the barn? Until now, the vine and the fig tree, the pomegranate and the olive tree have not borne fruit. "'From this day on I will bless you.'"
HAG|2|20|The word of the LORD came to Haggai a second time on the twenty-fourth day of the month:
HAG|2|21|"Tell Zerubbabel governor of Judah that I will shake the heavens and the earth.
HAG|2|22|I will overturn royal thrones and shatter the power of the foreign kingdoms. I will overthrow chariots and their drivers; horses and their riders will fall, each by the sword of his brother.
HAG|2|23|"'On that day,' declares the LORD Almighty, 'I will take you, my servant Zerubbabel son of Shealtiel,' declares the LORD, 'and I will make you like my signet ring, for I have chosen you,' declares the LORD Almighty."
