1JOHN|1|1|That which was from the beginning, which we have heard, which we have seen with our eyes, which we looked upon and have touched with our hands, concerning the word of life-
1JOHN|1|2|the life was made manifest, and we have seen it, and testify to it and proclaim to you the eternal life, which was with the Father and was made manifest to us-
1JOHN|1|3|that which we have seen and heard we proclaim also to you, so that you too may have fellowship with us; and indeed our fellowship is with the Father and with his Son Jesus Christ.
1JOHN|1|4|And we are writing these things so that our joy may be complete.
1JOHN|1|5|This is the message we have heard from him and proclaim to you, that God is light, and in him is no darkness at all.
1JOHN|1|6|If we say we have fellowship with him while we walk in darkness, we lie and do not practice the truth.
1JOHN|1|7|But if we walk in the light, as he is in the light, we have fellowship with one another, and the blood of Jesus his Son cleanses us from all sin.
1JOHN|1|8|If we say we have no sin, we deceive ourselves, and the truth is not in us.
1JOHN|1|9|If we confess our sins, he is faithful and just to forgive us our sins and to cleanse us from all unrighteousness.
1JOHN|1|10|If we say we have not sinned, we make him a liar, and his word is not in us.
1JOHN|2|1|My little children, I am writing these things to you so that you may not sin. But if anyone does sin, we have an advocate with the Father, Jesus Christ the righteous.
1JOHN|2|2|He is the propitiation for our sins, and not for ours only but also for the sins of the whole world.
1JOHN|2|3|And by this we know that we have come to know him, if we keep his commandments.
1JOHN|2|4|Whoever says "I know him" but does not keep his commandments is a liar, and the truth is not in him,
1JOHN|2|5|but whoever keeps his word, in him truly the love of God is perfected. By this we may be sure that we are in him:
1JOHN|2|6|whoever says he abides in him ought to walk in the same way in which he walked.
1JOHN|2|7|Beloved, I am writing you no new commandment, but an old commandment that you had from the beginning. The old commandment is the word that you have heard.
1JOHN|2|8|At the same time, it is a new commandment that I am writing to you, which is true in him and in you, because the darkness is passing away and the true light is already shining.
1JOHN|2|9|Whoever says he is in the light and hates his brother is still in darkness.
1JOHN|2|10|Whoever loves his brother abides in the light, and in him there is no cause for stumbling.
1JOHN|2|11|But whoever hates his brother is in the darkness and walks in the darkness, and does not know where he is going, because the darkness has blinded his eyes.
1JOHN|2|12|I am writing to you, little children, because your sins are forgiven for his name's sake.
1JOHN|2|13|I am writing to you, fathers, because you know him who is from the beginning. I am writing to you, young men, because you have overcome the evil one. I write to you, children, because you know the Father.
1JOHN|2|14|I write to you, fathers, because you know him who is from the beginning. I write to you, young men, because you are strong, and the word of God abides in you, and you have overcome the evil one.
1JOHN|2|15|Do not love the world or the things in the world. If anyone loves the world, the love of the Father is not in him.
1JOHN|2|16|For all that is in the world- the desires of the flesh and the desires of the eyes and pride in possessions- is not from the Father but is from the world.
1JOHN|2|17|And the world is passing away along with its desires, but whoever does the will of God abides forever.
1JOHN|2|18|Children, it is the last hour, and as you have heard that antichrist is coming, so now many antichrists have come. Therefore we know that it is the last hour.
1JOHN|2|19|They went out from us, but they were not of us; for if they had been of us, they would have continued with us. But they went out, that it might become plain that they all are not of us.
1JOHN|2|20|But you have been anointed by the Holy One, and you all have knowledge.
1JOHN|2|21|I write to you, not because you do not know the truth, but because you know it, and because no lie is of the truth.
1JOHN|2|22|Who is the liar but he who denies that Jesus is the Christ? This is the antichrist, he who denies the Father and the Son.
1JOHN|2|23|No one who denies the Son has the Father. Whoever confesses the Son has the Father also.
1JOHN|2|24|Let what you heard from the beginning abide in you. If what you heard from the beginning abides in you, then you too will abide in the Son and in the Father.
1JOHN|2|25|And this is the promise that he made to us- eternal life.
1JOHN|2|26|I write these things to you about those who are trying to deceive you.
1JOHN|2|27|But the anointing that you received from him abides in you, and you have no need that anyone should teach you. But as his anointing teaches you about everything- and is true and is no lie, just as it has taught you- abide in him.
1JOHN|2|28|And now, little children, abide in him, so that when he appears we may have confidence and not shrink from him in shame at his coming.
1JOHN|2|29|If you know that he is righteous, you may be sure that everyone who practices righteousness has been born of him.
1JOHN|3|1|See what kind of love the Father has given to us, that we should be called children of God; and so we are. The reason why the world does not know us is that it did not know him.
1JOHN|3|2|Beloved, we are God's children now, and what we will be has not yet appeared; but we know that when he appears we will be like him, because we shall see him as he is.
1JOHN|3|3|And everyone who thus hopes in him purifies himself as he is pure.
1JOHN|3|4|Everyone who makes a practice of sinning also practices lawlessness; sin is lawlessness.
1JOHN|3|5|You know that he appeared to take away sins, and in him there is no sin.
1JOHN|3|6|No one who abides in him keeps on sinning; no one who keeps on sinning has either seen him or known him.
1JOHN|3|7|Little children, let no one deceive you. Whoever practices righteousness is righteous, as he is righteous.
1JOHN|3|8|Whoever makes a practice of sinning is of the devil, for the devil has been sinning from the beginning. The reason the Son of God appeared was to destroy the works of the devil.
1JOHN|3|9|No one born of God makes a practice of sinning, for God's seed abides in him, and he cannot keep on sinning because he has been born of God.
1JOHN|3|10|By this it is evident who are the children of God, and who are the children of the devil: whoever does not practice righteousness is not of God, nor is the one who does not love his brother.
1JOHN|3|11|For this is the message that you have heard from the beginning, that we should love one another.
1JOHN|3|12|We should not be like Cain, who was of the evil one and murdered his brother. And why did he murder him? Because his own deeds were evil and his brother's righteous.
1JOHN|3|13|Do not be surprised, brothers, that the world hates you.
1JOHN|3|14|We know that we have passed out of death into life, because we love the brothers. Whoever does not love abides in death.
1JOHN|3|15|Everyone who hates his brother is a murderer, and you know that no murderer has eternal life abiding in him.
1JOHN|3|16|By this we know love, that he laid down his life for us, and we ought to lay down our lives for the brothers.
1JOHN|3|17|But if anyone has the world's goods and sees his brother in need, yet closes his heart against him, how does God's love abide in him?
1JOHN|3|18|Little children, let us not love in word or talk but in deed and in truth.
1JOHN|3|19|By this we shall know that we are of the truth and reassure our heart before him;
1JOHN|3|20|for whenever our heart condemns us, God is greater than our heart, and he knows everything.
1JOHN|3|21|Beloved, if our heart does not condemn us, we have confidence before God;
1JOHN|3|22|and whatever we ask we receive from him, because we keep his commandments and do what pleases him.
1JOHN|3|23|And this is his commandment, that we believe in the name of his Son Jesus Christ and love one another, just as he has commanded us.
1JOHN|3|24|Whoever keeps his commandments abides in him, and he in them. And by this we know that he abides in us, by the Spirit whom he has given us.
1JOHN|4|1|Beloved, do not believe every spirit, but test the spirits to see whether they are from God, for many false prophets have gone out into the world.
1JOHN|4|2|By this you know the Spirit of God: every spirit that confesses that Jesus Christ has come in the flesh is from God,
1JOHN|4|3|and every spirit that does not confess Jesus is not from God. This is the spirit of the antichrist, which you heard was coming and now is in the world already.
1JOHN|4|4|Little children, you are from God and have overcome them, for he who is in you is greater than he who is in the world.
1JOHN|4|5|They are from the world; therefore they speak from the world, and the world listens to them.
1JOHN|4|6|We are from God. Whoever knows God listens to us; whoever is not from God does not listen to us. By this we know the Spirit of truth and the spirit of error.
1JOHN|4|7|Beloved, let us love one another, for love is from God, and whoever loves has been born of God and knows God.
1JOHN|4|8|Anyone who does not love does not know God, because God is love.
1JOHN|4|9|In this the love of God was made manifest among us, that God sent his only Son into the world, so that we might live through him.
1JOHN|4|10|In this is love, not that we have loved God but that he loved us and sent his Son to be the propitiation for our sins.
1JOHN|4|11|Beloved, if God so loved us, we also ought to love one another.
1JOHN|4|12|No one has ever seen God; if we love one another, God abides in us and his love is perfected in us.
1JOHN|4|13|By this we know that we abide in him and he in us, because he has given us of his Spirit.
1JOHN|4|14|And we have seen and testify that the Father has sent his Son to be the Savior of the world.
1JOHN|4|15|Whoever confesses that Jesus is the Son of God, God abides in him, and he in God.
1JOHN|4|16|So we have come to know and to believe the love that God has for us. God is love, and whoever abides in love abides in God, and God abides in him.
1JOHN|4|17|By this is love perfected with us, so that we may have confidence for the day of judgment, because as he is so also are we in this world.
1JOHN|4|18|There is no fear in love, but perfect love casts out fear. For fear has to do with punishment, and whoever fears has not been perfected in love.
1JOHN|4|19|We love because he first loved us.
1JOHN|4|20|If anyone says, "I love God," and hates his brother, he is a liar; for he who does not love his brother whom he has seen cannot love God whom he has not seen.
1JOHN|4|21|And this commandment we have from him: whoever loves God must also love his brother.
1JOHN|5|1|Everyone who believes that Jesus is the Christ has been born of God, and everyone who loves the Father loves whomever has been born of him.
1JOHN|5|2|By this we know that we love the children of God, when we love God and obey his commandments.
1JOHN|5|3|For this is the love of God, that we keep his commandments. And his commandments are not burdensome.
1JOHN|5|4|For everyone who has been born of God overcomes the world. And this is the victory that has overcome the world- our faith.
1JOHN|5|5|Who is it that overcomes the world except the one who believes that Jesus is the Son of God?
1JOHN|5|6|This is he who came by water and blood- Jesus Christ; not by the water only but by the water and the blood. And the Spirit is the one who testifies, because the Spirit is the truth.
1JOHN|5|7|For there are three that testify:
1JOHN|5|8|the Spirit and the water and the blood; and these three agree.
1JOHN|5|9|If we receive the testimony of men, the testimony of God is greater, for this is the testimony of God that he has borne concerning his Son.
1JOHN|5|10|Whoever believes in the Son of God has the testimony in himself. Whoever does not believe God has made him a liar, because he has not believed in the testimony that God has borne concerning his Son.
1JOHN|5|11|And this is the testimony, that God gave us eternal life, and this life is in his Son.
1JOHN|5|12|Whoever has the Son has life; whoever does not have the Son of God does not have life.
1JOHN|5|13|I write these things to you who believe in the name of the Son of God that you may know that you have eternal life.
1JOHN|5|14|And this is the confidence that we have toward him, that if we ask anything according to his will he hears us.
1JOHN|5|15|And if we know that he hears us in whatever we ask, we know that we have the requests that we have asked of him.
1JOHN|5|16|If anyone sees his brother committing a sin not leading to death, he shall ask, and God will give him life- to those who commit sins that do not lead to death. There is sin that leads to death; I do not say that one should pray for that.
1JOHN|5|17|All wrongdoing is sin, but there is sin that does not lead to death.
1JOHN|5|18|We know that everyone who has been born of God does not keep on sinning, but he who was born of God protects him, and the evil one does not touch him.
1JOHN|5|19|We know that we are from God, and the whole world lies in the power of the evil one.
1JOHN|5|20|And we know that the Son of God has come and has given us understanding, so that we may know him who is true; and we are in him who is true, in his Son Jesus Christ. He is the true God and eternal life.
1JOHN|5|21|Little children, keep yourselves from idols.
