ESTH|1|1|І сталося за днів Ахашвероша, це той Ахашверош, що царював від Індії аж до Етіопії, сто й двадцять і сім округ,
ESTH|1|2|за тих днів, коли цар Ахашверош засів на троні свого царства, на замку Сузи.
ESTH|1|3|Третього року свого царювання справив він гостину для всіх своїх князів та для своїх слуг війська перського та мідійського, старших та правителів округ,
ESTH|1|4|показуючи багатство слави царства свого й пишну славу своєї величности довгі дні, сто й вісімдесят день.
ESTH|1|5|А по скінченні цих днів справив цар для всього народу, що знаходився в замку Сузи, від великого й аж до малого, гостину на сім день на садковому подвір'ї царського палацу.
ESTH|1|6|Біла, зелена та блакитна тканина, тримана віссоновими та пурпуровими шнурами, висіла на срібних стовпцях та мармурових колонах. Золоті та срібні ложа стояли на підлозі з плиток з зеленого, білого, жовтого й чорного мармуру.
ESTH|1|7|А напої подавали в золотому посуді, в посуді все різному, і царського вина було вельми щедро, за великою спроможністю царя.
ESTH|1|8|А пиття було за встановленим порядком, ніхто не примушував, бо цар так установив усім значним свого дому, щоб чинили за вподобою кожного.
ESTH|1|9|Також цариця Вашті справила гостину для жінок в царському домі царя Ахашвероша.
ESTH|1|10|Сьомого дня, коли цареві стало весело на серці від вина, він сказав Мегуманові, Біззеті, Харвоні, Біґті, і Аваґті, Зетарові та Каркасові, сімом евнухам, які служили перед обличчям царя Ахашвероша,
ESTH|1|11|привести царицю Вашті перед цареве обличчя в короні царській, щоб показати народам та зверхникам її красу, бо була вона вродливого вигляду.
ESTH|1|12|Та цариця Вашті відмовилася прийти за царським словом, що було передане їй через евнухів. І сильно загнівався цар, і в ньому горіла його лютість!
ESTH|1|13|І сказав цар до мудреців, що знають часи бо так царська справа йшла перед усіма, що знали закона та право,
ESTH|1|14|а близькими до нього були: Каршена, Шетар, Адмата, Паршіш, Мерес, Марсена, Мемухан, сім князів перських та мідійських, які бачать цареве обличчя й сидять перші в царстві:
ESTH|1|15|Як велить закон, щоб зробити з царицею Вашті за те, що не виконала слова царя Ахашвероша, переданого їй через евнухів?
ESTH|1|16|І сказав Мемухан перед царем та князями: Не перед самим царем провинилася цариця Вашті, але й перед усіма князями та перед усіма народами, що по всіх округах царя Ахашвероша.
ESTH|1|17|Бо царицин учинок дійде до всіх жінок, і спричиниться до погордження їхніх чоловіків в їхніх очах, бо будуть говорити: Цар Ахашверош сказав був привести царицю перед обличчя своє, та вона не прийшла!
ESTH|1|18|І цього дня казатимуть те саме княгині перські та мідійські, що почують про царицин учинок, до всіх царських князів, і буде багато погорди та гніву!
ESTH|1|19|Якщо цареві це добре, нехай вийде царський наказ від нього й нехай буде записане в законах Персії та Мідії, і нехай не поминеться, щоб Вашті більш не приходила перед обличчя царя Ахашвероша, а її царювання цар дасть іншій, ліпшій від неї.
ESTH|1|20|А коли почується царський наказ, який цар зробить відомим у всім своїм царстві, хоч яке велике воно, то всі жінки віддадуть честь своїм чоловікам, від великого й аж до малого.
ESTH|1|21|І була приємна ця рада в очах царя та князів, і цар зробив за Мемухановим словом.
ESTH|1|22|І порозсилав він листи до всіх царських округ, до кожної округи письмом її, і до кожного народу мовою його, щоб кожен чоловік був паном у домі своєму, і говорив про це мовою свого народу.
ESTH|2|1|По цих подіях, коли затихла лютість царя Ахашвероша, згадав він про Вашті, і що вона зробила, і що було заряджене про неї.
ESTH|2|2|І сказали царські отроки, його слуги: Нехай пошукають для царя дівчат, уродливих на вигляд паннів,
ESTH|2|3|і нехай цар призначить урядників по всіх округах свого царства, і нехай вони зберуть усіх дівчат, паннів уродливого вигляду, до замку Сузи, до дому жінок під руку Геґая, царського євнуха, сторожа жінок, і дати їм потрібне для їхнього причепурення.
ESTH|2|4|А та дівчина, що буде найкраща в царських очах, буде царювати замість Вашті. І була приємна ця рада у царевих очах, і він зробив так.
ESTH|2|5|А в замку Сузи був один юдеянин, а ім'я йому Мордехай, син Яіра, сина Шім'ї, сина Кішового, муж Веніяминівець,
ESTH|2|6|що був узятий з Єрусалиму з тим полоном, який був узятий разом з Єхонією, царем Юдиним, якого взяв був Навуходоносор, цар вавилонський.
ESTH|2|7|І він виховував Гадассу, вона ж Естер, дочку свого дядька, бо не мала вона ні батька, ні матері. А ця дівчина була хорошої постави та вродливого вигляду, а коли помер її батько та мати її, Мордехай узяв її собі за дочку.
ESTH|2|8|І сталося, коли був оголошений царський наказ та закон його, і коли збирали багато дівчат до замку Сузи під руку Геґая, то взята була й Естер до царського дому під руку Геґая, сторожа жінок.
ESTH|2|9|І була та дівчина хороша в його очах, і мала ласку перед ним, і він приспішив видати їй потрібне для її причепурення й її частки, та дати їй сімох відповідних дівчат із царського дому. І він перемістив її та дівчат її до найкращого місця в домі жінок.
ESTH|2|10|Естер не виявила ні про народ свій, ні про місце свого народження, бо Мордехай наказав їй, щоб цього вона не виявляла.
ESTH|2|11|А кожного дня Мордехай ходив до подвір'я дому жінок, щоб довідатись, як мається Естер та що вона робить.
ESTH|2|12|А коли приходила черга для кожної дівчини входити до царя Ахашвероша, коли кінчалися дванадцять місяців установленого порядку для жінок, бо так виповнялися дні їхнього причепурювання: шість місяців мирровою оливою, а шість місяців пахощами та іншим потрібним для причепурювання жінок,
ESTH|2|13|то з тим дівчина приходила до царя: давалося їй усе, що вона скаже, щоб воно йшло з нею з дому жінок до дому царського.
ESTH|2|14|Ввечорі вона приходила, а ранком вона верталася до другого дому жінок під руку Шаазґаза, царського евнуха, сторожа наложниць. Вона вже не входила до царя, хіба б що цар пожадав її, і вона була покликана за ім'ям.
ESTH|2|15|А коли настала черга для Естери, дочки Авіхая, Мордехаєвого дядька, що взяв її собі за дочку, щоб іти до царя, вона нічого не жадала, як тільки того, що казав Геґай, царський евнух, сторож жінок. І Естер мала ласку в очах усіх, хто її бачив!
ESTH|2|16|І була взята Естер до царя Ахашвероша, до царського дому його, десятого місяця, він місяць тевет, сьомого року царювання його.
ESTH|2|17|І цар покохав Естер понад усіх жінок, і вона мала прихильність та ласку перед його обличчям понад усіх дівчат, і він поклав царську корону на її голову, і зробив її царицею замість Вашті.
ESTH|2|18|І справив цар велику гостину для всіх своїх князів та своїх слуг, гостину для Естери, і зробив полегшення для округ, і дав дарунка за царською спроможністю.
ESTH|2|19|А коли збирали дівчат другий раз, то Мордехай сидів при царській брамі.
ESTH|2|20|Естер же не виявляла місця свого народження та народу свого, як наказав був їй Мордехай, бо Естер виконувала Мордехаєве слово так, як коли була в нього на вихованні.
ESTH|2|21|Тими днями, коли Мордехай сидів у царській брамі, розгнівалися Біґтан та Тереш, два царські евнухи зо сторожів порогів, і задумували простягнути руку на царя Ахашвероша.
ESTH|2|22|І стала відома ця річ Мордехаєві, і він доніс про це цариці Естер, а Естер переказала цареві в імені Мордехая.
ESTH|2|23|І була розвідана ця справа, і знайдено так, і ті обоє були повішені на шибениці. І було записане це в хроніці перед обличчям царським.
ESTH|3|1|По цих подіях цар Ахашверош звеличив Гамана, сина Гаммедатового, аґаґ'янина, і повищив його, і поставив його крісло понад усіх князів, що були з ним.
ESTH|3|2|А всі цареві раби, що були в царській брамі, падали на коліна та вклонялися Гаманові, бо так про нього наказав цар. А Мордехай не падав на коліна й не вклонявся.
ESTH|3|3|І сказали царські раби, що були в царській брамі, до Мордехая: Чого ти переступаєш царевого наказа?
ESTH|3|4|І сталося, як вони говорили до нього день-у-день, а він не слухався їх, то вони донесли Гаманові, щоб побачити, чи втримається Мордехай у своїм слові, бо він виявив їм, що він юдеянин.
ESTH|3|5|І побачив Гаман, що Мордехай не падає на коліна й не вклоняється йому, і Гаман переповнився лютістю...
ESTH|3|6|І погорджував він у своїх очах простягнути руку свою не тільки на Мордехая, самого його, бо донесли йому про Мордехаїв народ, і Гаман шукав випадку вигубити всіх юдеян, що були в усьому Ахашверошевому царстві, народ Мордехаїв.
ESTH|3|7|Першого місяця, він місяць нісан, дванадцятого року царя Ахашвероша, кидано пура, цебто жеребка, перед Гаманом із дня на день та з місяця на місяць, і жереб упав на дванадцятий місяць, він місяць адар.
ESTH|3|8|І сказав Гаман до царя Ахашвероша: Є один народ, розпорошений та поділений між народами в усіх округах твого царства, а закони їх різняться від законів усіх народів і законів царських вони не виконують, і цареві не варто позоставляти їх.
ESTH|3|9|Якщо це цареві вгодне, нехай буде написано вигубити їх, а я відважу десять тисяч талантів срібла на руки робітників, щоб унесли до царських скарбниць!
ESTH|3|10|І зняв цар персня свого зо своєї руки, і дав його Гаманові, синові Гаммедатовому, аґаґ'янинові, ненависникові юдеїв.
ESTH|3|11|І сказав цар до Гамана: Це срібло віддаю тобі, і дається тобі й той народ, щоб робити з ним, як угодно в очах твоїх!
ESTH|3|12|І були покликані царські писарі першого місяця тринадцятого дня в ньому, і було написано все так, як наказав Гаман до царських сатрапів та до намісників, що були над кожною скругою, і до князів кожного народу, до кожної округи письмом його, і до кожного народу мовою його; в імені царя Ахашвероша було написано, і припечатано було царським перснем.
ESTH|3|13|І були послані листи через гінців до всіх царських округ, щоб були повигублювані, побиті та понищені всі юдеї від хлопця й аж до старого, діти та жінки одного тринадцятого дня місяця дванадцятого, він місяць адар, а здобич по них пограбувати.
ESTH|3|14|Відпис із цього листа щоб був виданий як закон, у кожній окрузі, і оголошений для всіх народів, щоб були готові на цей день.
ESTH|3|15|Гінці вийшли, пігнані царевим словом. А закон був виданий в замку Сузи. А цар та Гаман сіли до пиття, а місто Сузи було в замішанні.
ESTH|4|1|А Мордехай довідався про все, що було зроблено. І роздер Мордехай одежу свою, і зодягнув веретище та посипався попелом, і вийшов на середину міста, та й кричав криком сильним та гірким!
ESTH|4|2|І прийшов він аж під царську браму, бо не можна було входити в царську браму в веретищному убранні.
ESTH|4|3|А в кожній окрузі та місці, куди доходило слово царя та його закон, були для юдеїв велика жалоба, і піст, і плач, і голосіння, а веретище та попел були ложем для багатьох...
ESTH|4|4|І прийшли дівчата Естерині й евнухи її, та й донесли їй про це. І дуже затремтіла цариця, і послала одежу зодягнути Мордехая та зняти з нього його веретище, та він не прийняв.
ESTH|4|5|І покликала Естер Гатаха, одного з евнухів царя, якого він приставив до неї, і наказала йому довідатися про Мордехая, що то з ним, і чого то жалоба?
ESTH|4|6|І вийшов Гатах на міську площу, що перед царською брамою.
ESTH|4|7|І виявив йому Мордехай усе, що спіткало його, і про суму срібла, яку Гаман сказав відважити до царської скарбниці за юдеїв, щоб вигубити їх.
ESTH|4|8|І він дав йому відписа листа закону, що був виданий у Сузах на вигублення їх, щоб показав Естері, та щоб доніс їй, і щоб наказав їй піти до царя благати його та просити перед його обличчям за її народ.
ESTH|4|9|І прийшов Гатах, і доніс Естері Мордехаєві слова.
ESTH|4|10|І сказала Естер до Гатаха, і наказала йому переказати Мордехаєві:
ESTH|4|11|Усі царські раби та народ царських округ знають, що кожен чоловік та жінка, що прийде до царя до внутрішнього подвір'я непокликаний, один йому закон, убити його, окрім того, кому цар простягне золоте берло, і буде він жити. А мене не кличуть входити до царя от уже тридцять день...
ESTH|4|12|І переказали Мордехаєві Естерині слова.
ESTH|4|13|І сказав Мордехай відповісти Естері: Не думай в душі своїй, що втечеш до царського дому одна з усіх юдеїв...
ESTH|4|14|Бо якщо справді будеш ти мовчати цього часу, то полегшення та врятування прийде для юдеїв з іншого місця, а ти та дім твого батька погинете. А хто знає, чи не на час, як оцей, досягла ти царства!...
ESTH|4|15|І сказала Естер відповісти Мордехаєві:
ESTH|4|16|Іди, збери всіх юдеїв, що знаходяться в Сузах, і постіть за мене, і не їжте й не пийте три дні, ніч та день. Також я та дівчата мої будемо постити так, і так прийду до царя, хоч це не буде за законом. А якщо я загину, то загину...
ESTH|4|17|І пішов Мордехай, і зробив усе, як звеліла йому Естер.
ESTH|5|1|І сталося третього дня, і вбрала Естер царські шати, та й стала на внутрішньому подвір'ї царського дому, навпроти царського дому. А цар сидів на троні свого царства в царському домі навпроти входу до дому.
ESTH|5|2|І сталося, як цар побачив царицю Естер, що стоїть у брамі, то знайшла вона ласку в очах його. І цар простягнув Естері золоте берло, що в руці його, а Естер підійшла й доторкнулася до кінця берла.
ESTH|5|3|І сказав до неї цар: Що тобі, царице Естер? І яке прохання твоє? Якщо побажаєш аж до половини царства, то буде дане тобі!
ESTH|5|4|А Естер відказала: Якщо це цареві вгодне, нехай прийде цар та Гаман сьогодні на гостину, яку я вчиню йому!
ESTH|5|5|І сказав цар: Скоріше покличте Гамана, щоб виконати Естерині слова! І прийшов цар та Гаман у гостину, що вчинила Естер.
ESTH|5|6|І сказав цар до Естери при питті вина: Яке жадання твоє? І буде тобі дане. І яке прохання твоє? Якщо побажаєш аж до половини царства, то буде зроблене!
ESTH|5|7|І відповіла Естер та й сказала: Моє жадання та моє прохання таке:
ESTH|5|8|Якщо знайшла я ласку в царевих очах, і якщо це цареві вгодне, щоб вволити жадання моє й щоб виконати прохання моє, нехай прийде цар та Гаман на гостину, що зроблю їм, і взавтра я зроблю за царевим словом.
ESTH|5|9|І вийшов Гаман того дня радісний та добросердий. Та коли Гаман побачив Мордехая в царській брамі, і він не встав і не затремтів перед ним, то Гаман переповнився лютістю на Мордехая.
ESTH|5|10|Та стримався Гаман, і прийшов до свого дому. І послав він покликати своїх приятелів та жінку свою Зереш.
ESTH|5|11|І розповів їм Гаман про славу свого багатства, та про численність синів своїх, та про все, як звеличив його цар, і як підняв його понад князів та слуг царевих.
ESTH|5|12|І сказав Гаман: А цариця Естер не привела з царем на гостину, яку зробила, нікого, крім мене. І також назавтра я покликаний до неї з царем!
ESTH|5|13|Та все це нічого не варте мені цього часу, доки я бачу того юдея Мордехая, що сидить у царській брамі!...
ESTH|5|14|І сказала до нього жінка його Зереш та всі його приятелі: Нехай приготують шибеницю, високу на п'ятдесят ліктів, а ранком скажи цареві, і нехай повісять на ній Мордехая, і підеш з царем радісний на гостину! І була приємна та рада для Гамана, і зробив він ту шибеницю.
ESTH|6|1|Тієї ночі втік був сон від царя, і він сказав принести Книгу пам'яток, Хроніки, і вони читалися перед обличчям царським.
ESTH|6|2|І знайдене було написане, що Мордехай доніс на Біґдана та Тереша, двох царських евнухів, зо сторожів порога, що задумували були простягнути руку на царя Ахашвероша.
ESTH|6|3|І сказав цар: Яка честь та гідність зроблена Мордехаєві за це? І сказали цареві отроки, що прислуговували йому: Нічого йому не зроблено...
ESTH|6|4|І спитав цар: Хто на подвір'ї? А Гаман прийшов на зовнішнє подвір'я царського дому, щоб сказати цареві повісити Мордехая на тій шибениці, яку приготовив для нього.
ESTH|6|5|І сказали отроки царя до нього: Ось Гаман стоїть на подвір'ї. І сказав цар: Нехай увійде!
ESTH|6|6|І Гаман увійшов, а цар йому сказав: Що зробити з чоловіком, якому цар хоче чести? І подумав Гаман у серці своїм: Кому ж цар зажадає вчинити честь більше, як мені?
ESTH|6|7|І відповів Гаман цареві: Тому чоловікові, якому цар жадає чести,
ESTH|6|8|нехай принесуть цареву одежу, яку цар зодягав, та коня, що цар їздив на ньому, і щоб була дана царська корона на його голову.
ESTH|6|9|І дати цю одежу та цього коня на руку котрогось із старших князів царевих. І нехай зодягнуть того чоловіка, якому цар жадає чести, і нехай возять його на коні на міській площі, і нехай кличуть перед ним: Так робиться мужеві, якому цар жадає чести!
ESTH|6|10|І сказав цар до Гамана: Поспіши, візьми одежу та коня, як казав ти, і зроби так юдеєві Мордехаєві, що сидить у царській брамі. Не пропусти нічого зо всього, що ти говорив!
ESTH|6|11|І взяв Гаман одежу та коня, і зодягнув Мордехая, і возив його на міській площі, і кричав перед ним: Так робиться мужеві, якому цар жадає чести!
ESTH|6|12|І вернувся Мордехай до царської брами, а Гаман поспішив до дому свого сумний та закривши голову...
ESTH|6|13|І розповів Гаман жінці своїй Зереші та всім приятелям своїм усе, що спіткало його. І сказали йому мудреці його та жінка його Зереш: Якщо з юдейського насіння Мордехай, перед яким зачав ти падати, то не переможеш його, бо дійсно впадеш перед ним!...
ESTH|6|14|Ще вони говорили з ним, а евнухи царські прибули й поспішили відвести Гамана на гостину, яку зробила Естер.
ESTH|7|1|І прийшов цар та Гаман на гостину цариці Естер.
ESTH|7|2|І сказав цар до Естери також другого дня при питті вина: Яке жадання твоє? І буде тобі дане. І яке прохання твоє? Якщо побажаєш аж до половини царства, то буде зроблено!
ESTH|7|3|І відповіла цариця Естер та й сказала: Якщо знайшла я ласку в очах твоїх, о царю, і якщо це цареві вгодне, нехай буде дане мені життя моє на жадання моє, а народ мій на прохання моє!
ESTH|7|4|Бо продані ми, я та народ мій, на вигублення, на забій та на погибіль... Та коли б ми були продані на рабів та на невільниць, мовчала б я, бо цей утиск був би не вартий царевого занепокоєння...
ESTH|7|5|Тоді сказав цар Ахашверош, і повів до цариці Естери: Хто то він, і де той, що його серце наповнило його відвагою чинити так?
ESTH|7|6|І сказала Естер: Ненависник та ворог це злий Гаман! І Гаман перелякався перед обличчям царя та цариці...
ESTH|7|7|А цар у своїй лютості устав від гостини, і вийшов до палацового саду. А Гаман став просити царицю Естер за життя своє, бо побачив, що загрожує йому лихо від царя...
ESTH|7|8|І цар вернувся з палацового саду до дому пиття вина, а Гаман припав до ліжка, що на ньому була Естер. І цар сказав: Чи хочеш також збезчестити царицю в мене в домі? Як тільки це слово вийшло з царевих уст, то закрили Гаманове обличчя...
ESTH|7|9|І сказав Харвона, один з евнухів перед царевим обличчям: Та ось шибениця, яку зробив Гаман для Мордехая, що говорив добре на царя, яка стоїть у Гамановому домі, висока на п'ятдесят ліктів. І сказав цар: Повісьте його на ній!
ESTH|7|10|І повісили Гамана на шибениці, яку він приготовив був для Мордехая, а лютість царева втихла...
ESTH|8|1|Того дня цар Ахашверош віддав цариці Естері дім Гамана, ненависника юдеїв, а Мордехай став перед цареве обличчя, бо Естер виявила, хто він для неї.
ESTH|8|2|І зняв цар свого персня, що забрав від Гамана, та й дав його Мордехаєві, а Естер настановила Мордехая над Гамановим домом.
ESTH|8|3|І Естер далі говорила перед обличчям царя. І впала вона перед його ногами, і плакала та благала його відвернути лихо аґаґ'янина Гамана та задуми його, які задумував був на юдеїв...
ESTH|8|4|І простягнув цар до Естери золоте берло, а Естер устала й стала перед царевим обличчям,
ESTH|8|5|та й сказала: Якщо це цареві вгодне, й якщо знайшла я ласку перед обличчям його, і вгодна ця річ перед царевим обличчям та вгодна я в очах його, нехай буде написано, щоб були повернені ті листи задумів аґаґ'янина Гамана, Гаммедатового сина, що написав був повигублювати юдеїв, які є в царевих округах.
ESTH|8|6|Бо як я могла б дивитися на лихо, що спіткає народ мій, і як я могла б дивитися на загибіль роду свого?
ESTH|8|7|І сказав цар Ахашверош до цариці Естери та до юдеянина Мордехая: Ось я дав Естері дім Гамана, а його повісили на шибениці за те, що простяг був руку свою на юдеїв.
ESTH|8|8|А ви пишіть до юдеїв, як добре в ваших очах, в імені царя, і припечатайте царським перснем, бо листа, що був написаний в імені царя та був припечатаний царським перснем, не можна відмінити.
ESTH|8|9|І були покликані царські писарі того часу, місяця третього, він місяць сіван, двадцять і третього дня в ньому, і було написане все, як наказав був Мордехай, до юдеїв, і до сатрапів, і намісників, і зверхників округ, що від Году й аж до Кушу, сто й двадцять і сім округ, і до кожної округи письмом її, і до кожного народу мовою його, та до юдеїв їхнім письмом та їхньою мовою.
ESTH|8|10|І понаписував він листи в імені царя Ахашвероша, і поприпечатував перснем царським, і послав через гінців на конях, які їздять на державних конях, конях баских,
ESTH|8|11|що цар дав право юдеям, які живуть у кожному місті, зібратися й стати за своє життя, вигубити, забити та погубити всяке військо народу та округи, що ненавидять їх, дітей та жінок, а здобич по них розграбувати,
ESTH|8|12|одного дня по всіх округах царя Ахашвероша, тринадцятого дня дванадцятого місяця, він місяць адар.
ESTH|8|13|Відпис цього листа щоб був виданий, як закон, у кожній окрузі, посланий був відкритий для всіх народів, і щоб юдеї були готові на той день помститися на своїх ворогах.
ESTH|8|14|Гінці, що поїхали верхи на швидких конях, вийшли, приспішені та пігнані царським словом. А цей наказ був даний у замку Сузи.
ESTH|8|15|А Мордехай вийшов з-перед царевого обличчя в царській одежі, блакитній та білій, а на ньому велика золота корона та віссонний і пурпуровий завій. І місто Сузи раділо та тішилося!
ESTH|8|16|Юдеям було тоді світло, і радість, і веселість, і честь!
ESTH|8|17|І в кожній окрузі та в кожному місті, куди досягає слово царя та закон його, була юдеям радість та веселість, бенкет та свято! І багато-хто з народів краю стали юдеями, бо на них напав страх перед юдеям.
ESTH|9|1|А дванадцятого місяця, він місяць адар, тринадцятого дня в ньому, коли наказ царя та закон його мали бути виконані, дня, коли вороги юдеїв сподівалися запанувати над ними, повернулося те так, що вони, юдеї, запанували над ненависниками своїми,
ESTH|9|2|зібралися юдеї в своїх містах по всіх округах царя Ахашвероша, щоб простягнути руку на тих, що задумували їм лихо, та ніхто не став перед ними, бо страх перед ними напав на всі народи.
ESTH|9|3|А всі зверхники округ, і сатрапи, і намісники, і виконавці царської праці підтримували юдеїв, бо напав на них страх перед Мордехаєм.
ESTH|9|4|Бо Мордехай став великим у царському домі, а вістка про нього покотилась по всіх округах, бо той чоловік, Мордехай, усе ріс.
ESTH|9|5|І били юдеї всіх своїх ворогів, побиваючи мечем, і забиваючи та вигублюючи їх, і робили з своїми ворогами за своєю волею.
ESTH|9|6|А в замку Сузи юдеї позабивали та повигублювали п'ять сотень чоловіка,
ESTH|9|7|і Паршандату, і Далфона, і Аспату,
ESTH|9|8|і Пората, і Адалію, і Арідата,
ESTH|9|9|і Пармашту, і Арісая, і Арідая, і Вайзата,
ESTH|9|10|десятьох синів Гамана, Гаммедатового сина, ненависника юдеїв, забили, а на грабунок не простягли своєї руки.
ESTH|9|11|Того дня число забитих у замку Сузи прийшло перед цареве обличчя.
ESTH|9|12|І сказав цар до цариці Естери: У замку Сузи юдеї позабивали та повигублювали п'ять сотень чоловіка та десятьох Гаманових синів. Що вони зробили в решті царевих округ? І яке жадання твоє? І буде тобі вволене. І яке ще прохання твоє? І буде зроблене.
ESTH|9|13|І відповіла Естер: Якщо це цареві вгодне, нехай буде дане юдеям, що в Сузах, також узавтра вчинити за законом цього дня, а десятьох Гаманових синів нехай повісять на шибениці.
ESTH|9|14|І сказав цар, щоб було зроблено так, і був даний закон у Сузах, а десятьох Гаманових синів повісили.
ESTH|9|15|І зібралися юдеї, що в Сузах, також чотирнадцятого дня місяця адар, і вибили в Сузах три сотні чоловіка, а на грабунок не простягли своєї руки.
ESTH|9|16|А решта юдеїв, що жили по царських округах, зібралися та й стали до бою за своє життя, і відпочили від ворогів своїх. І позабивали вони між своїми ненависниками сімдесят і п'ять тисяч, а на грабунок не простягли своєї руки.
ESTH|9|17|Це було тринадцятого дня місяця адара, а чотирнадцятого в ньому настав мир, і зробили його днем гостини та радости.
ESTH|9|18|А юдеї, що в Сузах, збиралися тринадцятого дня в ньому та чотирнадцятого в ньому, а мир мали п'ятнадцятого дня в ньому, і зробили його днем гостини та радости.
ESTH|9|19|Тому то юдеї неогороджених селищ, що сидять по неогороджених містах, роблять чотирнадцятий день місяця адара днем радости й гостини та свята, та днем посилання дарунків один одному.
ESTH|9|20|А Мордехай описав ці події, і порозсилав листи до всіх юдеїв, що по всіх округах царя Ахашвероша, до близьких та далеких,
ESTH|9|21|щоб вони постановили святкувати чотирнадцятий день місяця адара та п'ятнадцятий день у ньому кожного року,
ESTH|9|22|які ті дні, коли юдеї відпочили від ворогів своїх, і як той місяць, коли їм сум обернувся на радість, жалоба на свято, щоб зробити їх днями гостини та радости, і посилання дарунків один одному та дарунків убогим.
ESTH|9|23|І прийняли юдеї це, що зачали робити, і про що написав їм Мордехай,
ESTH|9|24|що аґаґ'янин Гаман, син Гаммедатів, ненависник усіх юдеїв, замишляв був на юдеїв, щоб вигубити їх, і кидав пура, цебто жеребка, на збентеження їх та на згубу їхню.
ESTH|9|25|Та коли прийшла вона, Естер, перед обличчя, царя він наказав листом: Нехай обернеться його злий задум, якого він задумав був на юдеїв, на його голову! І повісили його та синів його на шибениці.
ESTH|9|26|Тому то й назвали ці дні: Пурім, від імени пур. Тому то згідно зо всіма словами цього листа, і що вони бачили про це й що трапилося з ними,
ESTH|9|27|юдеї постановили й прийняли на себе й на нащадків своїх, та на всіх, хто поєднається з ними, і не відступлять, але щоб святкувати два ті дні кожного року згідно з написаним про них та згідно з їхнім часом.
ESTH|9|28|А дні ці мають споминатися та святкуватися в кожному поколінні, у кожному роді, у кожній окрузі, у кожному місті. А ці дні, Пурім, не минуться між юдеями, а пам'ять про них не скінчиться з їхнього насіння.
ESTH|9|29|І написала цариця Естер, дочка Авіхаїлова, та юдеянин Мордехай з сильним домаганням другий раз про те, щоб виконувати цього листа про Пурім.
ESTH|9|30|І порозсилав він листи до всіх юдеїв, до ста й двадцяти й семи округ Ахашверошового царства, зо словами миру та правди,
ESTH|9|31|щоб вони виконували ті дні Пурім у їх означених часах, як постановив про них юдеянин Мордехай та цариця Естер, і як вони самі постановили на себе та на нащадків своїх приписи постів та їхнього голосіння.
ESTH|9|32|А Естерин наказ ствердив ці приписи про Пурім, і було це записане в книгу.
ESTH|10|1|І наклав цар Ахашверош данину на землю та на морські острови.
ESTH|10|2|А ввесь чин його сили та його лицарських діл, і виразний опис величности Мордехая, що звеличив його цар, ось вони описані в Книзі Хронік царів мідійських та перських.
ESTH|10|3|Бо юдеянин Мордехай був другий по царі Ахашвероші, і великий для юдеїв, і милий для багатьох братів своїх, який шукав добра для народу свого й говорив мир! для всіх нащадків своїх.
