2KGS|1|1|亚哈 死后， 摩押 背叛 以色列 。
2KGS|1|2|亚哈谢 在 撒玛利亚 ，一日从楼上的栏杆跌下来，就病了。于是他派使者，对他们说：“你们去问 以革伦 的神明 巴力．西卜 ，我这病是否能痊愈。”
2KGS|1|3|但耶和华的使者对 提斯比 人 以利亚 说：“你起来，上去迎见 撒玛利亚 王的使者，对他们说：‘你们去问 以革伦 的神明 巴力．西卜 ，是因为 以色列 中没有上帝吗？’
2KGS|1|4|所以耶和华如此说：‘你必不能下你所上的床，因为你一定会死！’” 以利亚 就去了。
2KGS|1|5|使者回到王那里，王对他们说：“你们为什么回来了呢？”
2KGS|1|6|他们对王说：“有一个人上来迎见我们，对我们说：‘去，回到差你们来的王那里，对他说：耶和华如此说，你派人去问 以革伦 的神明 巴力．西卜 ，是因为 以色列 中没有上帝吗？所以你必不能下所上的床，你一定会死。’”
2KGS|1|7|王对他们说：“上来迎见你们，告诉你们这些话的人是什么样子呢？”
2KGS|1|8|他们对王说：“这人身穿毛衣 ，腰束皮带。”王说：“他一定是 提斯比 人 以利亚 。”
2KGS|1|9|于是，王派了一个五十夫长，带领五十人到 以利亚 那里。他上来，看哪， 以利亚 正坐在山顶上。五十夫长对他说：“神人哪，王吩咐你下来！”
2KGS|1|10|以利亚 回答五十夫长说：“我若是神人，愿火从天上降下来，吞灭你和你的五十个人！”于是有火从天上降下来，吞灭五十夫长和他的五十个人。
2KGS|1|11|王又派另一个五十夫长，带领五十人到 以利亚 那里。五十夫长对他说：“神人哪，王这样吩咐，快快下来！”
2KGS|1|12|以利亚 回答他们说：“我若是神人，愿火从天上降下来，吞灭你和你的五十个人！”于是上帝的火 从天上降下来，吞灭五十夫长和他的五十个人。
2KGS|1|13|王第三次又派一个五十夫长，带领五十人去。第三个五十夫长上去，双膝跪在 以利亚 面前，哀求他说：“神人哪，愿我的性命和你这五十个仆人的性命在你眼中看为宝贵！
2KGS|1|14|看哪，已经有火从天上降下来，吞灭前两次来的五十夫长和他们的五十个人，现在愿我的性命在你眼中看为宝贵！”
2KGS|1|15|耶和华的使者对 以利亚 说：“你跟他下去，不要怕他！” 以利亚 就起来，跟他下到王那里去。
2KGS|1|16|他对王说：“耶和华如此说：‘你派人去问 以革伦 的神明 巴力．西卜 ，是因为 以色列 中没有上帝可以让你求问他的话吗？所以你必不能下所上的床，你一定会死！’”
2KGS|1|17|亚哈谢 死了，正如耶和华藉 以利亚 所说的话。 犹大 王 约沙法 的儿子 约兰 第二年， 亚哈谢 的兄弟 约兰 接续他作王，因 亚哈谢 没有儿子。
2KGS|1|18|亚哈谢 其余所做的事，不都写在《以色列诸王记》上吗？
2KGS|2|1|耶和华要用旋风接 以利亚 升天的时候， 以利亚 与 以利沙 从 吉甲 往前行。
2KGS|2|2|以利亚 对 以利沙 说：“耶和华差遣我往 伯特利 去，你可以留在这里。” 以利沙 说：“我指着永生的耶和华，又指着你的性命起誓，我必不离开你。”于是二人下到 伯特利 。
2KGS|2|3|在 伯特利 的先知的门徒出来，到 以利沙 那里，对他说：“耶和华今日要接你的师父离开你 ，你知不知道？”他说：“我知道，你们不要作声。”
2KGS|2|4|以利亚 对 以利沙 说：“耶和华差遣我往 耶利哥 去，你可以留在这里。” 以利沙 说：“我指着永生的耶和华，又指着你的性命起誓，我必不离开你。”于是二人到了 耶利哥 。
2KGS|2|5|在 耶利哥 的先知的门徒来靠近 以利沙 ，对他说：“耶和华今日要接你的师父离开你，你知不知道？”他说：“我知道，你们不要作声。”
2KGS|2|6|以利亚 对 以利沙 说：“耶和华差遣我往 约旦河 去，你可以留在这里。” 以利沙 说：“我指着永生的耶和华，又指着你的性命起誓，我必不离开你。”于是二人一同往前行。
2KGS|2|7|有五十个先知的门徒同去，远远地站在他们对面；他们二人在 约旦河 边站住。
2KGS|2|8|以利亚 卷起自己的外衣，用来打水，水就左右分开，二人走干地过去。
2KGS|2|9|过去之后， 以利亚 对 以利沙 说：“我未被接去离开你以前，你要我为你做什么，只管求。” 以利沙 说：“愿感动你的灵双倍感动我。”
2KGS|2|10|以利亚 说：“你求的是一件难事。我被接去离开你的时候，你若看见我，就必得着；若不然，就得不着了。”
2KGS|2|11|他们边走边说话的时候，看哪，有火马和火焰车出现，把二人隔开， 以利亚 就乘旋风升天去了。
2KGS|2|12|以利沙 看见，就呼叫说：“我父啊！我父啊！ 以色列 的战车骑兵啊！” 以利沙 不再看见他的时候，就把自己的衣服撕为两片。
2KGS|2|13|他拾起 以利亚 身上掉下来的外衣，回去站在 约旦河 边。
2KGS|2|14|他用 以利亚 身上掉下来的外衣打水，说：“耶和华－ 以利亚 的上帝在哪里呢？”打水之后，水也左右分开， 以利沙 就过去了。
2KGS|2|15|在 耶利哥 的先知的门徒从对面看见他，说：“感动 以利亚 的灵临到 以利沙 身上了。”他们就来迎接他，俯伏于地，向他下拜，
2KGS|2|16|对他说：“看哪，仆人这里有五十个壮士，请你让他们去寻找你师父，或者耶和华的灵将他提起来，投在某山某谷。” 以利沙 说：“你们不必派人去。”
2KGS|2|17|他们再三催促，直到他不好意思，就说：“你们派人去吧！”他们就派了五十个人去，寻找了三天，也没有找着他。
2KGS|2|18|以利沙 仍然留在 耶利哥 ，他们回到他那里，他对他们说：“我不是告诉你们不必去吗？”
2KGS|2|19|耶利哥城 的人对 以利沙 说：“看哪，这城的地势美好，正如我主所看见的，只是水质恶劣，地也没有生产。”
2KGS|2|20|以利沙 说：“你们拿一个新的瓶子来，里面装盐。”他们就拿给他。
2KGS|2|21|他出去到了水源，把盐倒在那里，说：“耶和华如此说：‘我治好了这水，从那里不会再有死亡和不生产的事了。’”
2KGS|2|22|于是那水治好了，直到今日，正如 以利沙 所说的话。
2KGS|2|23|以利沙 从那里上 伯特利 去。正上路的时候，有些孩童从城里出来，讥笑他，对他说：“秃头的，上去吧！秃头的，上去吧！”
2KGS|2|24|他转过身来瞪着他们，奉耶和华的名诅咒他们。于是有两只母熊从林中出来，撕裂他们当中的四十二个孩童。
2KGS|2|25|以利沙 从 伯特利 上 迦密山 ，又从那里回到 撒玛利亚 。
2KGS|3|1|犹大 王 约沙法 第十八年， 亚哈 的儿子 约兰 在 撒玛利亚 登基，作 以色列 王十二年。
2KGS|3|2|他行耶和华眼中看为恶的事，但不致像他父母所行的，因为他除掉他父所造 巴力 的柱像。
2KGS|3|3|然而，他依恋 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪，总不离开。
2KGS|3|4|摩押 王 米沙 牧养许多羊，曾向 以色列 王进贡十万羔羊和十万公绵羊的毛。
2KGS|3|5|亚哈 死后， 摩押 王背叛 以色列 王。
2KGS|3|6|那时 约兰 王出 撒玛利亚 ，数点 以色列 众人。
2KGS|3|7|他向前行，派人到 犹大 王 约沙法 那里，说：“ 摩押 王背叛我，你肯同我去攻打 摩押 吗？” 约沙法 说：“我肯上去，你我不分彼此，我的军队就是你的军队，我的马就是你的马。”
2KGS|3|8|然后 约沙法 说：“我们从哪条路上去呢？” 约兰 说：“从 以东 旷野的路上去。”
2KGS|3|9|于是， 以色列 王和 犹大 王，以及 以东 王，都一同去。他们绕行了七日的路程，军队和所带的牲畜都没有水喝。
2KGS|3|10|以色列 王说：“哀哉！耶和华召集我们这三王，是要交在 摩押 人的手里。”
2KGS|3|11|约沙法 说：“这里不是有耶和华的先知吗？我们可以托他求问耶和华。” 以色列 王的一个大臣回答说：“这里有 沙法 的儿子 以利沙 ，就是从前服事 以利亚 的 。”
2KGS|3|12|约沙法 说：“他必有耶和华的话。”于是 以色列 王、 约沙法 和 以东 王都下去见他。
2KGS|3|13|以利沙 对 以色列 王说：“我跟你有什么关系呢？去问你父亲的先知和你母亲的先知吧！” 以色列 王对他说：“不，因为耶和华召集我们这三王，是要交在 摩押 人的手里。”
2KGS|3|14|以利沙 说：“我指着所事奉永生的万军之耶和华起誓，我若不看 犹大 王 约沙法 的情面，必不理你，不睬你。
2KGS|3|15|现在你们给我找一个弹琴的人来。”弹琴的人弹奏的时候，耶和华的手就按在 以利沙 身上。
2KGS|3|16|他就说：“耶和华如此说：‘你们要在这谷中到处挖沟。’
2KGS|3|17|因为耶和华如此说：‘你们虽不见风，也不见雨，这谷却必满了水，使你们和你们的牛羊牲畜都有水喝。’
2KGS|3|18|在耶和华眼中这还算是小事，他也必将 摩押 人交在你们手中。
2KGS|3|19|你们必攻破一切堡垒和美好的城镇，砍伐各种好树，塞住一切水泉，用石头毁坏一切良田。”
2KGS|3|20|到了早晨，约在献祭的时候，看哪，有水从 以东 而来，遍地就满了水。
2KGS|3|21|摩押 众人听见这三王上来要与他们打仗，凡能束上腰带的，无论老少，都被召集站在边界上。
2KGS|3|22|摩押 人清早起来，日光照在水上，他们看见对面水红如血，
2KGS|3|23|就说：“这是血啊！必是三王互相击杀，全都灭亡了。 摩押 人哪，我们现在去抢夺财物吧！”
2KGS|3|24|摩押 人到了 以色列 营， 以色列 人起来攻打他们，他们就在 以色列 人面前逃跑。 以色列 人追杀 摩押 人，直杀入 摩押 境内 。
2KGS|3|25|他们拆毁 摩押 的城镇，各人抛石头填满一切良田，塞住一切水泉，砍伐各种好树，只剩下 吉珥．哈列设 的石墙，但甩石的兵仍然包围攻打那城。
2KGS|3|26|摩押 王见战事激烈，对他不利，就率领七百个拿刀的兵，想突围逃到 以东 王那里，却没有成功。
2KGS|3|27|于是他在城墙上，把那应当接续他作王的长子献为燔祭。 有极大的愤怒临到 以色列 ，于是三王离开 摩押 王，各自回本地去了。
2KGS|4|1|有个先知门徒的妻子哀求 以利沙 说：“你的仆人，我丈夫死了，他敬畏耶和华是你所知道的。现在有债主来，要带走我的两个孩子给他作奴隶。”
2KGS|4|2|以利沙 对她说：“我可以为你做什么呢？告诉我，你家里有什么？”她说：“婢女家中除了一瓶油之外，什么也没有。”
2KGS|4|3|以利沙 说：“你到外面去向所有的邻舍借器皿，要空的器皿，不要少借。
2KGS|4|4|然后你回家，关上门，你和你儿子在里面把油倒在所有的器皿里，倒满了就放在一边。”
2KGS|4|5|于是妇人离开 以利沙 去了。她关上门，把自己和儿子关在家里。他们把器皿拿给她，她就倒油。
2KGS|4|6|器皿都满了，她对儿子说：“再给我拿器皿来。”儿子对她说：“没有器皿了。”油就止住了。
2KGS|4|7|妇人去告诉神人，神人说：“你去卖了油还债，你和你两个儿子可以靠着所剩的过活。”
2KGS|4|8|一日， 以利沙 经过 书念 ，在那里有一个富有的妇人强留他吃饭。此后， 以利沙 每次经过就转到那里去吃饭。
2KGS|4|9|妇人对丈夫说：“看哪，我知道那常从我们这里经过的是神圣的神人。
2KGS|4|10|我们可以为他盖一间有墙的小阁楼，里面安放床榻、桌子、椅子、灯台。每当他来到我们这里，就可以住在那里。”
2KGS|4|11|一日， 以利沙 来到那里，转进那阁楼，躺卧在那里。
2KGS|4|12|以利沙 吩咐仆人 基哈西 说：“你叫这 书念 妇人来。”他把妇人叫了来，妇人就站在 以利沙 面前。
2KGS|4|13|以利沙 吩咐仆人说：“你对她说：‘看哪，你为我们费了许多心思，我可以为你做什么呢？我可以为你向王或元帅求什么呢？’”她说：“我已住在自己百姓之中。”
2KGS|4|14|以利沙 说：“究竟可以为她做什么呢？” 基哈西 说：“她真的没有儿子，她丈夫也老了。”
2KGS|4|15|以利沙 说：“叫她回来。”于是他叫了她来，她就站在门口。
2KGS|4|16|以利沙 说：“明年这时候 ，你必抱一个儿子。”她说：“神人，我主啊，不要这样欺哄婢女。”
2KGS|4|17|妇人果然怀孕，到了明年那时候，生了一个儿子，正如 以利沙 向她所说的。
2KGS|4|18|孩子长大，一日出去到他父亲和收割的人那里。
2KGS|4|19|他对父亲说：“我的头啊，我的头啊！”他父亲对仆人说：“把他抱到他母亲那里。”
2KGS|4|20|仆人抱去，交给他母亲。孩子坐在母亲的膝上，到中午就死了。
2KGS|4|21|他母亲上去，把他放在神人的床上，关了门出来，
2KGS|4|22|呼叫她丈夫说：“你叫一个仆人给我牵一匹驴来，我要赶去见神人，然后回来。”
2KGS|4|23|丈夫说：“今日不是初一，也不是安息日，你为何要到他那里去呢？”妇人说：“平安无事。”
2KGS|4|24|于是她备上驴，对仆人说：“走，赶紧走，除非我吩咐你，不要为了我而慢下来。”
2KGS|4|25|妇人往 迦密山 去，到了神人那里。 神人远远看见她，对仆人 基哈西 说：“看哪， 书念 的妇人来了！
2KGS|4|26|现在你跑去迎接她，对她说，你平安吗？你丈夫平安吗？孩子平安吗？”她说：“平安。”
2KGS|4|27|妇人上了山，到神人那里，就抱住神人的脚。 基哈西 前来要推开她，神人说：“由她吧！因为她心里愁苦。但耶和华向我隐瞒这事，没有告诉我。”
2KGS|4|28|妇人说：“我何尝向我主求过儿子呢？我岂不是说过，不要欺哄我吗？”
2KGS|4|29|以利沙 吩咐 基哈西 说：“你束上腰，手拿我的杖前去。若遇见人，不要向他问安，人若向你问安，也不要回答。要把我的杖放在孩子脸上。”
2KGS|4|30|孩子的母亲说：“我指着永生的耶和华，又指着你的性命起誓，我必不离开你。”于是 以利沙 起身，随着她去了。
2KGS|4|31|基哈西 在他们以先去了，把杖放在孩子脸上，却没有声音，也没有动静。 基哈西 回去，迎见 以利沙 ，告诉他说：“孩子还没有醒过来。”
2KGS|4|32|以利沙 进了屋子，看哪，孩子死了，放在自己的床上。
2KGS|4|33|他进去，关上门，只有他们两个人，他就向耶和华祈祷。
2KGS|4|34|他上去伏在孩子身上，口对口，眼对眼，手对手。他伏在孩子身上，孩子的身体就渐渐暖和了。
2KGS|4|35|然后他下来，在屋里来回走了一趟，又上去伏在孩子身上。孩子打了七个喷嚏，眼睛就睁开了。
2KGS|4|36|以利沙 叫 基哈西 说：“你叫这 书念 妇人来。”于是他叫了她来。妇人来到 以利沙 那里， 以利沙 说：“把你儿子抱起来。”
2KGS|4|37|妇人就进来，在 以利沙 脚前俯伏于地，向他下拜，然后抱起她儿子出去了。
2KGS|4|38|以利沙 回到 吉甲 ，那地正有饥荒。先知的门徒坐在他面前，他吩咐仆人说：“你把大锅放在火上，给先知的门徒熬汤。”
2KGS|4|39|有一个人去到田野摘菜，发现一棵野瓜藤，就摘了满满一兜的野瓜回来，切了放进熬汤的锅中，并不知道那是什么。
2KGS|4|40|他们把汤倒出来给大家吃。他们吃汤里东西的时候，喊叫说：“神人哪，锅子里的东西会死人！”所以他们不能吃了。
2KGS|4|41|以利沙 说：“拿点面来。”他把面撒在锅中，说：“倒出来，给大家吃吧！”锅中就没有毒了。
2KGS|4|42|有一个人从 巴力．沙利沙 来，带着初熟果子的食物、二十个大麦做的饼和新麦穗，装在袋子里送给神人。神人说：“把这些给大家吃。”
2KGS|4|43|仆人说：“这些岂可摆在一百人面前呢？” 以利沙 说：“你只管给大家吃吧！因为耶和华如此说，他们必吃了，还有剩下的。”
2KGS|4|44|仆人就摆在他们面前，他们吃了，还有剩下，正如耶和华所说的。
2KGS|5|1|亚兰 王的元帅 乃缦 在他主人面前是一个伟大的人，得王的喜悦，因为耶和华曾藉他使 亚兰 人得胜。他虽然是大能的勇士，却染上了痲疯 。
2KGS|5|2|亚兰 人成群出征的时候，从 以色列 地掳了一个小女孩，她就服事 乃缦 的妻子。
2KGS|5|3|她对女主人说：“我希望主人去见 撒玛利亚 的先知，他必能治好主人的痲疯。”
2KGS|5|4|乃缦 去告诉他主人说，从 以色列 地来的女孩如此如此说。
2KGS|5|5|亚兰 王说：“你可以去，我也会送信给 以色列 王。”于是 乃缦 手里带十他连得银子、六千舍客勒金子和十套衣裳去了。
2KGS|5|6|他带着这信给 以色列 王，说：“现在你接到这信，看哪，我派臣仆 乃缦 到你这里来，你要治好他的痲疯。”
2KGS|5|7|以色列 王读了信就撕裂衣服，说：“我岂是上帝，能使人死使人活呢？这人竟派人来，叫我治好一个人的痲疯。你们要知道，看，这人是找机会来跟我吵架的。”
2KGS|5|8|神人 以利沙 听见 以色列 王撕裂衣服，就派人到王那里，说：“你为什么撕裂衣服呢？让那人到我这里来，他会知道 以色列 中有先知。”
2KGS|5|9|于是 乃缦 带着车马到了 以利沙 的家，站在门前。
2KGS|5|10|以利沙 派一个使者，对 乃缦 说：“去，在 约旦河 中沐浴七次，你的肉就必复原，你会得洁净。”
2KGS|5|11|乃缦 却发怒走了。他说：“看哪，我以为他必定会出来，到我这里，站着求告耶和华－他上帝的名，在患处上摇手，治好这痲疯。
2KGS|5|12|大马士革 的 亚玛拿河 和 法珥法河 岂不比 以色列 的一切水更好吗？我难道不可以在那里沐浴而得洁净吗？”于是他生气，转身走了。
2KGS|5|13|他的仆人近前来，对他说：“我父啊，先知若吩咐你做一件大事，你岂不做吗？何况是吩咐你去沐浴，得洁净呢？”
2KGS|5|14|于是 乃缦 下去，照着神人的话，在 约旦河 里浸了七次。他的肉复原，好像小孩的肉，他就洁净了。
2KGS|5|15|乃缦 带着所有跟随他的人，回到神人那里，站在他面前，说：“看哪，我知道，除了 以色列 ，全地没有上帝。现在请你收下仆人的礼物。”
2KGS|5|16|以利沙 说：“我指着所事奉永生的耶和华起誓，我必不接受。” 乃缦 再三请他收下，他却不肯。
2KGS|5|17|乃缦 说：“你若不肯，请把两匹骡子能驮的土赐给仆人，仆人必不再把燔祭或祭物献给别神，只献给耶和华。
2KGS|5|18|惟有一件事，愿耶和华饶恕你仆人：我主人进 临门 庙在那里叩拜的时候，他总是扶着我的手，所以我也在 临门 庙叩拜。我在 临门 庙叩拜的这事，愿耶和华饶恕你仆人。”
2KGS|5|19|以利沙 对他说：“你平安地回去吧！” 乃缦 离开他去了。走了一小段路，
2KGS|5|20|神人 以利沙 的仆人 基哈西 说：“看哪，我主人不愿从这 亚兰 人 乃缦 手里接受他带来的礼物，我指着永生的耶和华起誓，我必跑去追上他，向他拿些东西。”
2KGS|5|21|于是 基哈西 去追 乃缦 。 乃缦 看见有人追来，就下车迎着他，说：“都平安吗？”
2KGS|5|22|他说：“都平安！我主人派我来说：‘看哪，现在有两个年轻人，是先知的门徒，从 以法莲 山区来到我这里，请你给他们一他连得银子，两套衣裳。’”
2KGS|5|23|乃缦 说：“好啊，请收下二他连得。”他再三请求，就把二他连得银子装在两个袋子里，连同两套衣裳交给两个仆人；他们就在 基哈西 前头抬着走。
2KGS|5|24|到了山冈， 基哈西 从他们手中接过来，放在屋里，打发这些人走了。
2KGS|5|25|基哈西 进去，站在主人面前。 以利沙 对他说：“ 基哈西 ，你从哪里来？”他说：“仆人哪里也没去。”
2KGS|5|26|以利沙 对他说：“那人下车转过来迎着你的时候，我的心岂没有去呢？这岂是接受银子，接受衣裳、橄榄园、葡萄园、牛羊、仆婢的时候呢？
2KGS|5|27|因此， 乃缦 的痲疯必紧随你和你的后裔，直到永远。” 基哈西 从 以利沙 面前出去，就长了痲疯，像雪一样。
2KGS|6|1|先知的门徒对 以利沙 说：“看哪，我们在你面前居住的地方，那里对我们太窄小了。
2KGS|6|2|让我们往 约旦河 去，各人从那里取一根木料，在那里为自己建造居住的地方。”他说：“你们去吧！”
2KGS|6|3|有一人说：“请你与仆人同去。”他说：“我可以去。”
2KGS|6|4|于是 以利沙 与他们同去。到了 约旦河 ，他们砍伐树木。
2KGS|6|5|有一人砍树的时候，斧子的头掉在水里，他就喊着说：“不好了！我主啊，斧子是借来的。”
2KGS|6|6|神人说：“掉在哪里了？”他把那地方指给 以利沙 看。 以利沙 砍了一块木头，抛在水里，就使斧子的头浮上来了。
2KGS|6|7|以利沙 说：“拿起来吧！”那人就伸手拿起来了。
2KGS|6|8|亚兰 王与 以色列 作战，他和臣仆商议说：“我要在某处某处安营 。”
2KGS|6|9|神人派人到 以色列 王那里，说：“你要小心，不要从某处经过，因为 亚兰 人下到那里去了。”
2KGS|6|10|以色列 王派人到神人告诉他的地方去。神人警告他，他就在那里有所防备，不止一两次。
2KGS|6|11|亚兰 王因这事心里气愤，召了臣仆来，对他们说：“我们当中有谁帮助 以色列 王，你们不告诉我吗？”
2KGS|6|12|有一个臣仆说：“不，我主，我王！只有 以色列 中的先知 以利沙 ，把王在卧房所说的话告诉 以色列 王。”
2KGS|6|13|王说：“你们去查看他在哪里，我好派人去捉拿他。”有人告诉王说：“看哪，他在 多坍 。”
2KGS|6|14|王就派遣车马和大军往那里去，夜间他们到了，围困那城。
2KGS|6|15|神人的仆人清早起来出去，看哪，车马军兵围困了城。仆人对神人说：“不好了！我主啊，我们该怎么办呢？”
2KGS|6|16|神人说：“不要惧怕！因与我们同在的比与他们同在的更多。”
2KGS|6|17|以利沙 祷告说：“耶和华啊，求你开他的眼目，使他能看见。”耶和华开了这年轻人的眼目，他就看见了，看哪，满山有火马和火焰车围绕 以利沙 。
2KGS|6|18|亚兰 人下到 以利沙 那里， 以利沙 向耶和华祷告说：“求你击打这国，使他们眼目失明。”耶和华就照 以利沙 的话，击打他们，使他们眼目失明。
2KGS|6|19|以利沙 对他们说：“这不是那条路，也不是那座城。你们跟我走，我必领你们到你们要寻找的人那里。”于是他领他们到了 撒玛利亚 。
2KGS|6|20|他们进了 撒玛利亚 ， 以利沙 说：“耶和华啊，求你开这些人的眼目，使他们能看见。”耶和华开了他们的眼目，他们就看见了，看哪，是在 撒玛利亚城 中。
2KGS|6|21|以色列 王看见他们，就对 以利沙 说：“我父啊，我真的可以击杀他们吗？”
2KGS|6|22|他说：“不可击杀！这些人岂是你用刀用弓掳来给你击杀的呢？当在他们面前摆设饮食给他们吃喝，让他们回到他们主人那里。”
2KGS|6|23|王为他们预备了盛大的宴席。他们吃喝完了，王就送他们回到他们主人那里。此后， 亚兰 的军队不再侵犯 以色列 地了。
2KGS|6|24|此后， 亚兰 王 便．哈达 召集他的全军，上来围困 撒玛利亚 。
2KGS|6|25|看哪，被围困的时候， 撒玛利亚 有大饥荒，甚至一个驴头值八十舍客勒，四分之一卡布 的鸽子粪值五舍客勒。
2KGS|6|26|一日， 以色列 王在城墙上经过，有一个妇人向他呼叫说：“我主，我王啊！求你帮助。”
2KGS|6|27|王说：“耶和华不帮助你，我从哪里帮助你呢？是从禾场，或从压酒池吗？”
2KGS|6|28|王对妇人说：“你有什么事？”她说：“这妇人对我说：‘把你的儿子交出来，我们今日可以吃他，明日可以吃我的儿子。’
2KGS|6|29|我们就煮了我的儿子吃了。次日我对她说：‘要把你的儿子交出来，我们可以吃。’她却把她的儿子藏起来。”
2KGS|6|30|王听见妇人的话，就撕裂衣服；那时，王在城墙上经过，百姓看见了，看哪，王贴身穿着麻布。
2KGS|6|31|王说：“我今日若容许 沙法 的儿子 以利沙 的头还留在他身上，愿上帝重重惩罚我！”
2KGS|6|32|那时， 以利沙 正坐在家中，有长老与他同坐。王派一个人先去，使者还没有到， 以利沙 对长老说：“你们看，这凶手之子派人来斩我的头。你们注意，当使者来到，你们就关上门，把他关在门外。在他后头不就是他主人的脚步声吗？”
2KGS|6|33|正与他们说话的时候，看哪，使者 下到他那里，说：“看哪，这灾祸是从耶和华来的，我何必再仰望耶和华呢？”
2KGS|7|1|以利沙 说：“你们要听耶和华的话，耶和华如此说：明日约这时候，在 撒玛利亚 城门口，一细亚细面只卖一舍客勒，二细亚大麦也卖一舍客勒。”
2KGS|7|2|有一个搀扶王的军官回答神人说：“看哪，即使耶和华打开天上的窗户，也不可能有这事。” 以利沙 说：“看哪，你必亲眼看见，在那里却吃不到什么。”
2KGS|7|3|在城门口有四个长痲疯的人，他们彼此说：“我们为何坐在这里等死呢？
2KGS|7|4|我们若说要进城去，城里有饥荒，我们必死在那里。若我们在这里坐着不动，也必死。现在，来吧，我们去向 亚兰 人的军队投降。若他们饶我们的命，我们就活着；若杀我们，我们就死吧！”
2KGS|7|5|黄昏的时候，他们起来往 亚兰 人的军营去；到了营边，看哪，没有一人在那里。
2KGS|7|6|因为主使 亚兰 人的军队听见战车战马的声音，大军的声音，他们就彼此说：“看哪，这必是 以色列 王雇用 赫 人诸王和 埃及 诸王来攻击我们。”
2KGS|7|7|所以，在黄昏的时候他们起来逃跑，撇下帐棚、马、驴，把军营留在原处，只顾逃命。
2KGS|7|8|那些长痲疯的人到了营边，进了一座帐棚，吃了喝了，从当中拿走金银和衣服，收藏起来。他们又回来，进了另一座帐棚，从当中拿走财物去收藏。
2KGS|7|9|那时，他们彼此说：“我们所做的不对了！这一天是有好消息的日子，我们竟不作声！若等到天亮，我们就有罪了。现在，来，我们去向王室报信吧！”
2KGS|7|10|他们就去叫守城门的人，告诉他们说：“我们到了 亚兰 人的军营，看哪，没有一人在那里，也无人声，只有拴着的马和驴，帐棚都留在原处。”
2KGS|7|11|守城门的人就呼叫，他们向城内的王室报信。
2KGS|7|12|王夜间起来，对臣仆说：“我告诉你们 亚兰 人向我们做的事。他们知道我们饥饿，所以离营，埋伏在田野，说：‘ 以色列 人出城的时候，我们活捉他们，我们就可以进到城里去。’”
2KGS|7|13|王的一个臣仆回答说：“不如叫人从城里剩下的马中取五匹，看哪，这些马像 以色列 大众一样 ，快要灭亡了；我们派人去窥探吧！”
2KGS|7|14|于是他们取了两辆车和马，王派人去跟踪 亚兰 人的军队，说：“你们去窥探吧。”
2KGS|7|15|他们去跟踪 亚兰 人，直到 约旦河 。看哪，整条路上都是 亚兰 人匆忙逃跑时所丢弃的衣服和器具，使者就回来向王报告。
2KGS|7|16|百姓就出去，掳掠 亚兰 人的军营。于是一细亚细面只卖一舍客勒，二细亚大麦也卖一舍客勒，正如耶和华所说的。
2KGS|7|17|王派搀扶他的那军官在城门指挥，百姓在城门把他踩死了，正如神人在王下到他那里的时候所说的。
2KGS|7|18|神人曾对王说：“明日约这时候，在 撒玛利亚 城门口，二细亚大麦只卖一舍客勒，一细亚细面也卖一舍客勒。”
2KGS|7|19|那军官回答神人说：“看哪，即使耶和华打开天上的窗户，也不可能有这事。”神人说：“看哪，你必亲眼看见，在那里却吃不到什么。”
2KGS|7|20|这话果然应验在他身上，因为百姓在城门把他踩死了。
2KGS|8|1|以利沙 曾对他救活的孩子的母亲说：“你和你的全家要起身，往你可住的地方去住，因为耶和华已令饥荒降在这地七年。”
2KGS|8|2|妇人就起身，照神人的话去做，带着全家往 非利士 人的地去，寄居了七年。
2KGS|8|3|过了七年，那妇人从 非利士 人的地回来，就出去为自己的房屋田地哀求王。
2KGS|8|4|那时王正与神人的仆人 基哈西 谈话，说：“你把 以利沙 所做的一切大事告诉我。”
2KGS|8|5|基哈西 告诉王 以利沙 如何使死人复活，看哪， 以利沙 所救活的孩子的母亲正为自己的房屋田地来哀求王。 基哈西 说：“我主我王，这就是那妇人，这是她的儿子，就是 以利沙 所救活的。”
2KGS|8|6|王问那妇人，她就把事情告诉王。于是王为她派一个官员，说：“凡属这妇人的都还给她，自从她离开本地直到今日，她田地的出产也都还给她。”
2KGS|8|7|以利沙 来到 大马士革 ， 亚兰 王 便．哈达 正患病。有人告诉王说：“神人来到这里了。”
2KGS|8|8|王就吩咐 哈薛 说：“你带着礼物去见神人，托他求问耶和华，我这病能不能好？”
2KGS|8|9|于是 哈薛 用四十匹骆驼，驮着 大马士革 的各样美物为礼物，去迎见 以利沙 。 哈薛 到了那里，站在他面前，说：“你儿子 亚兰 王 便．哈达 派我到你这里，问说：‘我这病会不会好？’”
2KGS|8|10|以利沙 对 哈薛 说：“你回去告诉他说：‘你一定会好。’但耶和华指示我，他必定会死。”
2KGS|8|11|神人定睛看着 哈薛 ，直到他感到羞愧。神人就哭了。
2KGS|8|12|哈薛 说：“我主为什么哭？”他说：“因为我知道你必虐待 以色列 人，用火焚烧他们的堡垒，用刀杀死他们的壮丁，摔死他们的婴孩，剖开他们的孕妇。”
2KGS|8|13|哈薛 说：“仆人算什么，不过是一条狗，怎么能行这大事呢？” 以利沙 说：“耶和华指示我，你必作 亚兰 王。”
2KGS|8|14|哈薛 离开 以利沙 ，回到他主人那里。主人对他说：“ 以利沙 对你说了什么？”他说：“他告诉我你必能好。”
2KGS|8|15|次日， 哈薛 拿被子浸在水中，蒙住王的脸，王就死了。于是 哈薛 篡了他的位。
2KGS|8|16|亚哈 的儿子 以色列 王 约兰 第五年－ 约沙法 曾作 犹大 王 － 犹大 王 约沙法 的儿子 约兰 登基作了 犹大 王。
2KGS|8|17|约兰 登基的时候年三十二岁，在 耶路撒冷 作王八年。
2KGS|8|18|他行 以色列 诸王的道，正如 亚哈 家所行的，因他娶了 亚哈 的女儿为妻，行耶和华眼中看为恶的事。
2KGS|8|19|耶和华却因他仆人 大卫 的缘故，不肯灭绝 犹大 ，要照他所应许的，永远赐灯光给 大卫 和他的子孙。
2KGS|8|20|约兰 在位期间， 以东 背叛，自己立王治理他们，脱离 犹大 的权势。
2KGS|8|21|约兰 率领他所有的战车过到 撒益 去。他夜间起来，攻打围困他的 以东 人和战车长； 犹大 军兵逃跑，各回自己的帐棚去了；
2KGS|8|22|这样， 以东 背叛，脱离 犹大 的管辖，直到今日。那时 立拿 也背叛了。
2KGS|8|23|约兰 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|8|24|约兰 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 亚哈谢 接续他作王。
2KGS|8|25|亚哈 的儿子 以色列 王 约兰 第十二年， 犹大 王 约兰 的儿子 亚哈谢 登基。
2KGS|8|26|他登基的时候年二十二岁，在 耶路撒冷 作王一年。他母亲名叫 亚她利雅 ，是 以色列 王 暗利 的孙女。
2KGS|8|27|亚哈谢 行 亚哈 家的道，行耶和华眼中看为恶的事，与 亚哈 家一样，因为他是 亚哈 家的女婿。
2KGS|8|28|他与 亚哈 的儿子 约兰 同往 基列 的 拉末 去，与 亚兰 王 哈薛 交战。 亚兰 人打伤了 约兰 ，
2KGS|8|29|约兰 王回到 耶斯列 ，医治在 拉末 与 亚兰 王 哈薛 打仗时，被 亚兰 人击打所受的伤。 约兰 的儿子 犹大 王 亚哈谢 因为 亚哈 的儿子 约兰 病了，就下到 耶斯列 看望他。
2KGS|9|1|以利沙 先知叫了一个先知的门徒来，吩咐他：“你束上腰，手拿这瓶膏油往 基列 的 拉末 去。
2KGS|9|2|你到了那里，要在那里寻找 宁示 的孙子， 约沙法 的儿子 耶户 。你去，使他从弟兄中起来，带他进最里面的内室，
2KGS|9|3|把瓶里的膏油倒在他头上，说：‘耶和华如此说：我膏你作 以色列 王。’然后你就开门逃跑，不要等候。”
2KGS|9|4|于是那青年，那年轻的先知往 基列 的 拉末 去了。
2KGS|9|5|他到了那里，看哪，众军官都坐着，就说：“长官，我有话对你说。” 耶户 说：“你要对我们哪一个说呢？”他说：“长官，我要对你说。”
2KGS|9|6|耶户 就起来，进了内室，那青年把膏油倒在他头上，对他说：“耶和华－ 以色列 的上帝如此说：‘我膏你作耶和华百姓 以色列 的王。
2KGS|9|7|你要击杀你主人 亚哈 的全家，我好在 耶洗别 身上，为我仆人众先知和耶和华所有仆人的血伸冤。
2KGS|9|8|亚哈 全家都必灭亡，凡属 亚哈 的男丁，无论是奴役的、自由的，我必从 以色列 中剪除。
2KGS|9|9|我必使 亚哈 的家像 尼八 儿子 耶罗波安 的家，又像 亚希雅 儿子 巴沙 的家。
2KGS|9|10|至于 耶洗别 ，狗必在 耶斯列 田里吃她，无人埋葬。’”于是那青年就开门逃跑了。
2KGS|9|11|耶户 出来，回到他主人的臣仆那里，有一人问他说：“平安吗？这疯狂的人为什么到你这里来呢？”他对他们说：“你们认得那人，也知道他在胡说。”
2KGS|9|12|他们说：“说谎！告诉我们吧。”他说：“他如此如此对我说：‘耶和华如此说：我膏你作 以色列 的王。’”
2KGS|9|13|他们各人就急忙把自己的衣服铺在台阶的上层，在 耶户 的下面；他们吹角，说：“ 耶户 作王了！”
2KGS|9|14|这样， 宁示 的孙子， 约沙法 的儿子 耶户 背叛了 约兰 。先前 约兰 和 以色列 众人因为 亚兰 王 哈薛 的缘故，把守 基列 的 拉末 。
2KGS|9|15|后来 约兰 王回到 耶斯列 ，医治他与 亚兰 王 哈薛 打仗时，被 亚兰 人击打所受的伤。 耶户 说：“若你们有这样的意思，就不要让人溜出城，到 耶斯列 去报信。”
2KGS|9|16|于是 耶户 驾战车往 耶斯列 去，因为 约兰 卧病在那里。 犹大 王 亚哈谢 已经下去看望他。
2KGS|9|17|有一个守望的人站在 耶斯列 的城楼上，看见 耶户 带着一队人来，就说：“我看见一队人。” 约兰 说：“派一个骑兵去迎接他们，问说：‘平安吗？’”
2KGS|9|18|骑兵就去迎接 耶户 ，说：“王如此说：‘平安吗？’”耶户说：“平安不平安跟你有什么关系呢？转身跟在我后面吧！”守望的人说：“使者到了他们那里，却不回来。”
2KGS|9|19|王又派第二个骑兵去。这人到了他们那里，说：“王如此说：‘平安吗？’” 耶户 说：“平安不平安跟你有什么关系呢？转身跟在我后面吧！”
2KGS|9|20|守望的人又说：“他到了他们那里，也不回来。车驾得很凶猛，好像 宁示 的孙子 耶户 在驾车。”
2KGS|9|21|约兰 吩咐说：“套车！”人就给他套车。 以色列 王 约兰 和 犹大 王 亚哈谢 各坐自己的车出去迎接 耶户 ，在 耶斯列 人 拿伯 的田那里遇见他。
2KGS|9|22|约兰 见 耶户 就说：“ 耶户 ，平安吗？” 耶户 说：“你母亲 耶洗别 的淫行邪术这样多，怎么能平安呢？”
2KGS|9|23|约兰 用手转过车来逃跑，对 亚哈谢 说：“ 亚哈谢 啊，反了！”
2KGS|9|24|耶户 全力拉弓，射中 约兰 两臂中间，箭从心窝穿出， 约兰 就仆倒在车上。
2KGS|9|25|耶户 对他的军官 毕甲 说：“把他抛在 耶斯列 人 拿伯 的田里。你当记得，你我一同驾车跟随他父亲 亚哈 的时候，耶和华对 亚哈 说了预言，
2KGS|9|26|耶和华说：‘我昨日看见 拿伯 的血和他众子的血，我发誓我必在这块田上报应你。’这是耶和华说的。现在你要照着耶和华的话，把他抛在这田里。”
2KGS|9|27|犹大 王 亚哈谢 看见了，就沿着 伯．哈干 的路逃跑。 耶户 追赶他，说：“把这人也击杀在车上，在靠近 以伯莲 的 姑珥 坡上 。”他逃到 米吉多 ，就死在那里。
2KGS|9|28|他的臣仆用车把他的尸体运回 耶路撒冷 ，与他祖先同葬在 大卫城 ，他自己的坟墓里。
2KGS|9|29|亚哈 的儿子 约兰 第十一年， 亚哈谢 登基作了 犹大 王。
2KGS|9|30|耶户 到了 耶斯列 。 耶洗别 听见了，就画眼影、梳头，从窗户往外观看。
2KGS|9|31|耶户 进了城门， 耶洗别 说：“杀主人的 心利 啊，平安吗？”
2KGS|9|32|耶户 向窗户抬头，说：“有谁顺从我？谁？”有两三个太监向外看他。
2KGS|9|33|耶户 说：“把她抛下来！”他们就把她抛下来。她的血溅在墙上和马上， 耶户 践踏在她身上。
2KGS|9|34|耶户 进去，吃了喝了，说：“你们去处理这被诅咒的妇人，埋了她，因为她是王的女儿。”
2KGS|9|35|他们去了，要埋葬她，却只找到她的头骨和脚，以及手掌。
2KGS|9|36|他们回来报告 耶户 ， 耶户 说：“这正应验耶和华藉他仆人 提斯比 人 以利亚 所说的话，说：‘在 耶斯列 田里，狗必吃 耶洗别 的肉，
2KGS|9|37|耶洗别 的尸体必在 耶斯列 田里的地面上如同粪土，甚至没有人可说：这是 耶洗别 。’”
2KGS|10|1|亚哈 有七十个儿子在 撒玛利亚 。 耶户 写信送到 撒玛利亚 ，给 耶斯列 的领袖和长老 ，以及教养 亚哈 众儿子的人，说：
2KGS|10|2|“你们主人的众儿子既然在你们那里，你们又有战车、马匹、兵器、坚固城，现在你们接了这信，
2KGS|10|3|可以在你们主人的众儿子中选一个贤能正直的，使他坐他父亲的王位，你们也可以为你们主人的家作战。”
2KGS|10|4|他们却非常惧怕，说：“看哪，两个王在他面前尚且站立不住，我们怎能站立得住呢？”
2KGS|10|5|王宫总管、市长和长老，并教养众儿子的人，派人到 耶户 那里，说：“我们是你的仆人，凡你所吩咐的，我们都必遵行。我们不立谁作王，你看怎样好就怎样做吧。”
2KGS|10|6|耶户 写第二封信给他们，说：“你们若归顺我，听从我的话，明日这时候，要带着你们主人众儿子的首级，来到 耶斯列 我这里。”那时王的儿子七十人都住在城中教养他们的那些尊贵人家里。
2KGS|10|7|信一到他们那里，他们就把王的七十个儿子杀了，将首级装在筐里，送到 耶斯列 ， 耶户 那里。
2KGS|10|8|有使者来告诉 耶户 说：“他们把王众儿子的首级送来了。” 耶户 说：“把首级分成两堆，放在城门口，直到早晨。”
2KGS|10|9|次日早晨， 耶户 出来，站着对众百姓说：“你们都是公义的！看哪，我背叛了我的主人，把他杀了，但这所有的人又是谁杀的呢？
2KGS|10|10|由此可知，耶和华指着 亚哈 家所说的话一句也没有落空，因为耶和华实现了他藉他仆人 以利亚 所说的话。”
2KGS|10|11|凡 亚哈 家在 耶斯列 所剩下的，他的大臣、密友、祭司， 耶户 全都杀了，没有留下一个幸存者。
2KGS|10|12|耶户 起身往 撒玛利亚 去。路途中，在牧人聚集的 伯．艾克特 ，
2KGS|10|13|耶户 遇见 犹大 王 亚哈谢 的兄弟，说：“你们是谁？”他们说：“我们是 亚哈谢 的兄弟，现在下去要向王和太后的众儿子问安。”
2KGS|10|14|耶户 说：“活捉他们！”人就活捉了他们，把他们杀在 伯．艾克特 的坑边，共四十二人，一个也没有留下。
2KGS|10|15|耶户 从那里往前行，遇见 利甲 的儿子 约拿达 来迎接他， 耶户 向他问安，对他说：“你的心 ，像我的心待你的心那样正直吗？” 约拿达 说：“是。” 耶户 说：“若是这样，请你伸出手来。”他伸出手， 耶户 就拉他上车。
2KGS|10|16|耶户 说：“你和我同去，看我为耶和华怎样热心。”于是他们请他坐在车上。
2KGS|10|17|到了 撒玛利亚 ， 耶户 把 亚哈 家在 撒玛利亚 剩下的人全都杀了，直到灭尽，正如耶和华对 以利亚 所说的话。
2KGS|10|18|耶户 召集众百姓，对他们说：“ 亚哈 事奉 巴力 还不够热心， 耶户 更要热心。
2KGS|10|19|现在你们召集 巴力 的众先知和所有拜 巴力 的人，以及 巴力 的众祭司，都到我这里来，一个也不可缺少，因为我要给 巴力 献大祭；凡不来的必不得活。” 耶户 行诡诈，为要消灭拜 巴力 的人。
2KGS|10|20|耶户 说：“要为 巴力 召集严肃会！”于是他们宣告了。
2KGS|10|21|耶户 派人走遍 以色列 ；凡拜 巴力 的人都来齐了，没有留下一个不来的。他们进了 巴力 庙， 巴力 庙中前后都挤满了人。
2KGS|10|22|耶户 对掌管服装的人说：“拿出袍子来，给所有拜 巴力 的人穿。”他就拿出礼服来给了他们。
2KGS|10|23|耶户 和 利甲 的儿子 约拿达 进了 巴力 庙，对拜 巴力 的人说：“你们要搜查察看，不可以有耶和华的仆人在你们这里，只可以有拜 巴力 的人。”
2KGS|10|24|他们进去，献上祭物和燔祭． 耶户 先安排八十人在庙外，说：“我把这些人交在你们手中，谁放走其中一人，谁就要以命偿命！”
2KGS|10|25|耶户 献完了燔祭，就对护卫兵和众军官说：“进去杀他们，不要让一人逃脱！”护卫兵和军官用刀杀了他们，将尸体抛出去，然后进入 巴力 庙的堡垒，
2KGS|10|26|将 巴力 庙中的柱像都 拿出来焚烧。
2KGS|10|27|他们毁坏 巴力 的柱像，拆毁了 巴力 庙当厕所，直到今日。
2KGS|10|28|这样， 耶户 在 以色列 中消灭了 巴力 。
2KGS|10|29|只是 耶户 不离开 尼八 的儿子 耶罗波安 使 以色列 人陷入罪里的那罪，就是拜 伯特利 和 但 的金牛犊。
2KGS|10|30|耶和华对 耶户 说：“因你办好我眼中看为正的事，照我的心意待 亚哈 家，你的子孙必接续你坐 以色列 的王位，直到第四代。”
2KGS|10|31|只是 耶户 不尽心遵守耶和华－ 以色列 上帝的律法，不离开 耶罗波安 使 以色列 人陷入罪里的那罪。
2KGS|10|32|在那些日子，耶和华开始削弱 以色列 。 哈薛 在 以色列 各边界攻击他们，
2KGS|10|33|就是 约旦河 东 基列 全地，从靠近 亚嫩谷 边的 亚罗珥 起，包括 基列 和 巴珊 ，就是 迦得 人、 吕便 人、 玛拿西 人的地。
2KGS|10|34|耶户 其余的事，凡他所做的和他英勇的事迹，不都写在《以色列诸王记》上吗？
2KGS|10|35|耶户 与他祖先同睡，葬在 撒玛利亚 ，他儿子 约哈斯 接续他作王。
2KGS|10|36|耶户 在 撒玛利亚 作 以色列 王二十八年。
2KGS|11|1|亚哈谢 的母亲 亚她利雅 见她儿子死了，就起来剿灭王室所有的后裔。
2KGS|11|2|但 约兰 王的女儿， 亚哈谢 的妹妹 约示巴 ，将 亚哈谢 的儿子 约阿施 从被杀的王子中偷出来，把他和他的奶妈藏在卧房里，躲避了 亚她利雅 ，没有被杀。
2KGS|11|3|亚她利雅 治理这地的时候， 约阿施 和他的奶妈在耶和华的殿里藏了六年。
2KGS|11|4|第七年， 耶何耶大 派人叫 迦利 人和护卫兵的众百夫长来，领他们进耶和华的殿，与他们立约，使他们在耶和华殿里起誓，又把王的儿子指给他们看，
2KGS|11|5|吩咐他们说：“你们要这样做：你们当中在安息日值班的，三分之一要把守王宫，
2KGS|11|6|三分之一要在 苏珥门 ，三分之一要在护卫兵院的后门；你们要这样轮流把守王宫。
2KGS|11|7|你们安息日所有不值班的两队人员要在耶和华的殿里护卫王；
2KGS|11|8|各人手拿兵器，四围保护王。凡擅自闯入你们行列的，要被处死。王出入的时候，你们当跟随他。”
2KGS|11|9|众百夫长就照着 耶何耶大 祭司一切所吩咐的去做，各带自己的人，无论安息日值班或不值班的，都到 耶何耶大 祭司那里。
2KGS|11|10|祭司就把耶和华殿里所藏 大卫 王的枪和盾牌交给百夫长。
2KGS|11|11|护卫兵手中各拿兵器，在祭坛和殿那里，从殿南到殿北，站在王的四围。
2KGS|11|12|耶何耶大 领 约阿施 出来，给他戴上冠冕，把律法书交给他，膏他作王；众人都鼓掌说：“愿王万岁！”
2KGS|11|13|亚她利雅 听见护卫兵和百姓的声音，就进耶和华的殿，到百姓那里。
2KGS|11|14|她观看，看哪，王照仪式站在柱旁，百夫长和号手在王旁边，国中的众百姓欢乐吹号。 亚她利雅 就撕裂衣服，喊着说：“反了！反了！”
2KGS|11|15|耶何耶大 祭司吩咐管军兵的百夫长，对他们说：“把她从行列之间赶出去，凡跟随她的必用刀杀死！”因为祭司说：“不可在耶和华殿里杀她。”
2KGS|11|16|他们就下手拿住她；她进入通往王宫的 马门 ，就在那里被杀。
2KGS|11|17|耶何耶大 使王和百姓与耶和华立约，作耶和华的子民，又使王与百姓立约。
2KGS|11|18|于是国中的众百姓都到 巴力 庙去，拆毁了庙，彻底打碎祭坛和偶像，又在坛前把 巴力 的祭司 玛坦 杀了。 耶何耶大 祭司派官员看守耶和华的殿，
2KGS|11|19|又率领百夫长， 迦利 人和护卫兵，以及国中的众百姓，请王从耶和华的殿下来，由护卫兵的门进入王宫，他就坐上王位。
2KGS|11|20|国中的众百姓都欢乐，合城也都平静。他们已将 亚她利雅 在王宫那里用刀杀了。
2KGS|11|21|约阿施 登基的时候年方七岁。
2KGS|12|1|耶户 第七年， 约阿施 登基，在 耶路撒冷 作王四十年。他母亲名叫 西比亚 ，是 别是巴 人。
2KGS|12|2|约阿施 在 耶何耶大 祭司教导他的一切日子，行耶和华眼中看为正的事。
2KGS|12|3|只是丘坛还没有废去，百姓仍在丘坛献祭烧香。
2KGS|12|4|约阿施 对众祭司说：“凡献到耶和华殿分别为圣的银子，无论是人的赎价，各人生命的赎价， 或自愿献给耶和华殿的银子，
2KGS|12|5|祭司可以各自从认识的人收取，用来修理殿的破坏之处，就是在那里发现的一切破坏之处。”
2KGS|12|6|然而，到了 约阿施 王第二十三年，祭司仍未修理殿的破坏之处。
2KGS|12|7|所以 约阿施 王召了 耶何耶大 祭司和众祭司来，对他们说：“你们怎么不修理殿的破坏之处呢？现在，不要再从认识的人收银子了，但要为了殿的破坏之处，把银子交出来。”
2KGS|12|8|众祭司答应不再收百姓的银子，也不再修理殿的破坏之处。
2KGS|12|9|耶何耶大 祭司取了一个柜子，在柜盖上钻了一个洞，放在祭坛旁，在进耶和华殿的右边；守门的祭司将献到耶和华殿的一切银子投在柜里。
2KGS|12|10|他们见柜里的银子多了，就叫王的书记和大祭司上来，将耶和华殿里所得的银子数点了，包起来。
2KGS|12|11|他们把秤好了的银子交在管理耶和华殿督工的手里，督工就支付给木匠和建造耶和华殿的工人，
2KGS|12|12|瓦匠和石匠，又买木料和凿成的石头，用来修理耶和华殿的破坏之处，以及其他修理殿的各项费用。
2KGS|12|13|但这些献到耶和华殿的银子，并没有用来造耶和华殿里的银杯、钳子、盘子、号筒和其他的金银器皿。
2KGS|12|14|他们把这银子交给工人，用来整修耶和华的殿。
2KGS|12|15|他们不用跟这些经手接受银子去支付工人的人算账，因为这些人办事诚实。
2KGS|12|16|赎愆祭和赎罪祭的银子没有献到耶和华的殿里，都归给祭司。
2KGS|12|17|那时， 亚兰 王 哈薛 上来攻打 迦特 ，攻取了它。 哈薛 就定意上来攻打 耶路撒冷 。
2KGS|12|18|犹大 王 约阿施 将他祖先 犹大 王 约沙法 、 约兰 、 亚哈谢 所分别为圣的物和自己所分别为圣的物，以及耶和华殿与王宫府库里所有的金子都送给 亚兰 王 哈薛 ； 哈薛 就不上 耶路撒冷 来了。
2KGS|12|19|约阿施 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|12|20|约阿施 的臣仆起来背叛，在下到 悉拉 路上的 米罗 宫那里把他杀了。
2KGS|12|21|杀他的臣仆就是 示米押 的儿子 约撒拔 和 朔默 的儿子 约萨拔 。他与祖先同葬在 大卫城 ，他儿子 亚玛谢 接续他作王。
2KGS|13|1|亚哈谢 的儿子 犹大 王 约阿施 第二十三年， 耶户 的儿子 约哈斯 在 撒玛利亚 登基作 以色列 王十七年。
2KGS|13|2|约哈斯 行耶和华眼中看为恶的事，效法 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪，总不离开。
2KGS|13|3|于是，耶和华的怒气向 以色列 发作，将他们屡次交在 亚兰 王 哈薛 和他儿子 便．哈达 的手里。
2KGS|13|4|约哈斯 恳求耶和华，耶和华就应允他，因为耶和华看见 以色列 所受的欺压，因 亚兰 王欺压他们。
2KGS|13|5|耶和华赐给 以色列 一位拯救者，使他们脱离 亚兰 人的手，于是 以色列 人仍旧安居在自己的帐棚里。
2KGS|13|6|然而他们不离开 耶罗波安 家使 以色列 陷入罪里的那罪，仍行在罪中，并且在 撒玛利亚 留下 亚舍拉 。
2KGS|13|7|亚兰 王灭绝 约哈斯 的军队，践踏他们如禾场上的尘沙，只给 约哈斯 留下五十骑兵，十辆战车，一万步兵。
2KGS|13|8|约哈斯 其余的事，凡他所做的和他英勇的事迹，不都写在《以色列诸王记》上吗？
2KGS|13|9|约哈斯 与他祖先同睡，葬在 撒玛利亚 ，他儿子 约阿施 接续他作王。
2KGS|13|10|犹大 王 约阿施 第三十七年， 约哈斯 的儿子 约阿施 在 撒玛利亚 登基作 以色列 王十六年。
2KGS|13|11|他行耶和华眼中看为恶的事，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的一切罪，仍行在罪中。
2KGS|13|12|约阿施 其余的事，凡他所做的和他与 犹大 王 亚玛谢 交战的英勇事迹，不都写在《以色列诸王记》上吗？
2KGS|13|13|约阿施 与他祖先同睡， 耶罗波安 坐上他的王位。 约阿施 与 以色列 诸王一同葬在 撒玛利亚 。
2KGS|13|14|以利沙 得了致命的病， 以色列 王 约阿施 下来看他，伏在他脸上哭泣，说：“我父啊！我父啊！ 以色列 的战车和骑兵啊！”
2KGS|13|15|以利沙 对他说：“把弓箭拿来。”王就拿了弓箭来。
2KGS|13|16|以利沙 对 以色列 王说：“你用手开弓。”王就用手开弓。 以利沙 按手在王的手上，
2KGS|13|17|说：“打开朝东的窗户。”他就打开。 以利沙 说：“射箭！”他就射箭。 以利沙 说：“这是耶和华得胜的箭，是战胜 亚兰 人的箭，因为你必在 亚弗 攻打 亚兰 人，直到灭尽他们。”
2KGS|13|18|以利沙 又说：“拿几枝箭来。”他就拿了来。 以利沙 对 以色列 王说：“打地吧！”他打了三次，就停止了。
2KGS|13|19|神人向他发怒，说：“你应当击打五六次，就能攻打 亚兰 人直到灭尽；现在你只能打败 亚兰 人三次。”
2KGS|13|20|以利沙 死了，人把他埋葬了。新的一年， 摩押 人成群结队入侵境内。
2KGS|13|21|有人正在埋葬死人，看哪，他们看见一群人来，就把死人抛在 以利沙 的坟墓里，逃跑了。死人一碰到 以利沙 的骸骨，就活过来，用脚站了起来。
2KGS|13|22|约哈斯 在位年间， 亚兰 王 哈薛 屡次欺压 以色列 。
2KGS|13|23|耶和华却因与 亚伯拉罕 、 以撒 、 雅各 所立的约，仍施恩给 以色列 人，怜悯他们，眷顾他们，不肯灭尽他们，直到现在 仍不赶逐他们离开自己面前。
2KGS|13|24|亚兰 王 哈薛 死了，他儿子 便．哈达 接续他作王。
2KGS|13|25|从前 哈薛 和 约阿施 的父亲 约哈斯 交战，攻取了些城镇，现在 约哈斯 的儿子 约阿施 三次打败 哈薛 的儿子 便．哈达 ，从他手中收回了 以色列 的城镇。
2KGS|14|1|约哈斯 的儿子 以色列 王 约阿施 第二年， 犹大 王 约阿施 的儿子 亚玛谢 登基。
2KGS|14|2|他登基的时候年二十五岁，在 耶路撒冷 作王二十九年。他母亲名叫 约耶但 ，是 耶路撒冷 人。
2KGS|14|3|亚玛谢 行耶和华眼中看为正的事，但不如他祖先 大卫 。他效法他父亲 约阿施 一切所行的。
2KGS|14|4|只是丘坛还没有废去，百姓仍在丘坛献祭烧香。
2KGS|14|5|王国在他手里巩固的时候，他就把杀他父王的臣仆杀了，
2KGS|14|6|却没有处死杀王凶手的儿子，正如 摩西 律法书上耶和华所吩咐的说：“不可因子杀父，也不可因父杀子，各人要为自己的罪而死。”
2KGS|14|7|亚玛谢 在 盐谷 杀了一万 以东 人，又在战役中攻取了 西拉 ，称它为 约帖 ，直到今日。
2KGS|14|8|那时， 亚玛谢 派使者到 耶户 的孙子， 约哈斯 的儿子 以色列 王 约阿施 那里，说：“来，让我们面对面较量吧！”
2KGS|14|9|以色列 王 约阿施 派人去见 犹大 王 亚玛谢 ，说：“ 黎巴嫩 的蒺藜派人去见 黎巴嫩 的香柏树，说：‘将你的女儿嫁给我的儿子。’但有一只野兽经过 黎巴嫩 ，把蒺藜践踏了。
2KGS|14|10|你果然打败了 以东 ，就心高气傲。你以此为荣，就待在自己家里算了吧，为何要惹祸，使自己和 犹大 一同败亡呢？”
2KGS|14|11|亚玛谢 却不肯听从。于是 以色列 王 约阿施 上来，在 犹大 的 伯．示麦 与 犹大 王 亚玛谢 面对面较量。
2KGS|14|12|犹大 败在 以色列 面前，他们逃跑，各人逃回自己的帐棚去了。
2KGS|14|13|以色列 王 约阿施 在 伯．示麦 擒住 亚哈谢 的孙子， 约阿施 的儿子 犹大 王 亚玛谢 ，就来到 耶路撒冷 ，拆毁 耶路撒冷 的城墙，从 以法莲门 直到 角门 共四百肘。
2KGS|14|14|他又拿了耶和华殿里与王宫府库里所有的金银和器皿，并带着人质，回 撒玛利亚 去了。
2KGS|14|15|约阿施 其余所做的事和他英勇的事迹，以及他与 犹大 王 亚玛谢 交战的事，不都写在《以色列诸王记》上吗？
2KGS|14|16|约阿施 与他祖先同睡，与 以色列 诸王一同葬在 撒玛利亚 ，他儿子 耶罗波安 接续他作王。
2KGS|14|17|约哈斯 的儿子 以色列 王 约阿施 死后， 犹大 王 约阿施 的儿子 亚玛谢 又活了十五年。
2KGS|14|18|亚玛谢 其余的事，不都写在《犹大列王记》上吗？
2KGS|14|19|耶路撒冷 有人背叛 亚玛谢 ， 亚玛谢 逃往 拉吉 ；他们却派人追到 拉吉 ，在那里杀了他。
2KGS|14|20|有人用马将他驮回，葬在 耶路撒冷 ，与他祖先一同葬在 大卫城 。
2KGS|14|21|犹大 众百姓立 亚撒利雅 接续他父亲 亚玛谢 作王，那时他年十六岁。
2KGS|14|22|亚玛谢 王与他祖先同睡之后， 亚撒利雅 收复 以拉他 回归 犹大 ，又重新整修。
2KGS|14|23|约阿施 的儿子 犹大 王 亚玛谢 第十五年， 以色列 王 约阿施 的儿子 耶罗波安 在 撒玛利亚 登基，作王四十一年。
2KGS|14|24|他行耶和华眼中看为恶的事，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的一切罪。
2KGS|14|25|他收回 以色列 边界之地，从 哈马口 直到 亚拉巴海 ，正如耶和华－ 以色列 的上帝藉他仆人 迦特．希弗 人 亚米太 的儿子 约拿 先知所说的。
2KGS|14|26|因耶和华看见 以色列 非常艰苦的困境；没有奴役的，没有自由的，也没有人来帮助 以色列 。
2KGS|14|27|耶和华并没有说要将 以色列 的名从天下涂抹，却要藉 约阿施 的儿子 耶罗波安 拯救他们。
2KGS|14|28|耶罗波安 其余的事，凡他所做的和他英勇的事迹，他怎样作战，怎样收复 大马士革 和先前属 犹大 的 哈马 回归 以色列 ，不都写在《以色列诸王记》上吗？
2KGS|14|29|耶罗波安 与他祖先 以色列 诸王同睡，他儿子 撒迦利雅 接续他作王。
2KGS|15|1|以色列 王 耶罗波安 第二十七年， 犹大 王 亚玛谢 的儿子 亚撒利雅 登基。
2KGS|15|2|他登基的时候年十六岁，在 耶路撒冷 作王五十二年。他母亲名叫 耶可利雅 ，是 耶路撒冷 人。
2KGS|15|3|亚撒利雅 行耶和华眼中看为正的事，效法他父亲 亚玛谢 一切所行的。
2KGS|15|4|只是丘坛还没有废去，百姓仍在丘坛献祭烧香。
2KGS|15|5|耶和华降灾于王，使他长了痲疯，直到死的那日。他住在隔离的行宫里，他儿子 约坦 管理王的家，治理这地的百姓。
2KGS|15|6|亚撒利雅 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|15|7|亚撒利雅 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 约坦 接续他作王。
2KGS|15|8|犹大 王 亚撒利雅 第三十八年， 耶罗波安 的儿子 撒迦利雅 登基，在 撒玛利亚 作 以色列 王六个月。
2KGS|15|9|他行耶和华眼中看为恶的事，效法他祖先所行的，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪。
2KGS|15|10|雅比 的儿子 沙龙 背叛他，在百姓面前 击杀他，篡了他的位。
2KGS|15|11|撒迦利雅 其余的事，看哪，都写在《以色列诸王记》上。
2KGS|15|12|这就是耶和华应许 耶户 的话：“你的子孙必坐 以色列 的王位，直到第四代。”这事果然发生了。
2KGS|15|13|犹大 王 乌西雅 第三十九年， 雅比 的儿子 沙龙 登基，在 撒玛利亚 作王一个月。
2KGS|15|14|迦底 的儿子 米拿现 从 得撒 上 撒玛利亚 ，杀了 雅比 的儿子 沙龙 ，篡了他的位。
2KGS|15|15|沙龙 其余的事和他阴谋背叛的事，看哪，都写在《以色列诸王记》上。
2KGS|15|16|那时， 米拿现 从 得撒 起击杀 提斐萨 和城中所有的人，以及它周围的地区，因为他们没有给他开城门。他击杀他们，剖开其中所有的孕妇。
2KGS|15|17|犹大 王 亚撒利雅 第三十九年， 迦底 的儿子 米拿现 登基，在 撒玛利亚 作 以色列 王十年。
2KGS|15|18|他行耶和华眼中看为恶的事，终生不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪。
2KGS|15|19|亚述 王 普勒 来攻击这地， 米拿现 给他一千他连得银子，为了请 普勒 帮助他巩固他所掌握的国度。
2KGS|15|20|米拿现 向 以色列 所有的富豪索取银子，要他们各出五十舍客勒，交给 亚述 王。于是 亚述 王回去了，不在境内停留。
2KGS|15|21|米拿现 其余的事，凡他所做的，不都写在《以色列诸王记》上吗？
2KGS|15|22|米拿现 与他祖先同睡，他儿子 比加辖 接续他作王。
2KGS|15|23|犹大 王 亚撒利雅 第五十年， 米拿现 的儿子 比加辖 登基，在 撒玛利亚 作 以色列 王二年。
2KGS|15|24|他行耶和华眼中看为恶的事，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪。
2KGS|15|25|比加辖 的将军， 利玛利 的儿子 比加 背叛他，在 撒玛利亚 王宫的堡垒杀了他。 亚珥歌伯 和 亚利耶 并 基列 的五十人帮助 比加 ； 比加 击杀他，篡了他的位。
2KGS|15|26|比加辖 其余的事，凡他所做的，看哪，都写在《以色列诸王记》上。
2KGS|15|27|犹大 王 亚撒利雅 第五十二年， 利玛利 的儿子 比加 登基，在 撒玛利亚 作 以色列 王二十年。
2KGS|15|28|他行耶和华眼中看为恶的事，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪。
2KGS|15|29|在 以色列 王 比加 的日子， 亚述 王 提革拉．毗列色 来夺取 以云 、 亚伯．伯．玛迦 、 亚挪 、 基低斯 、 夏琐 、 基列 、 加利利 和 拿弗他利 全地，把这些地方的居民都掳到 亚述 去了。
2KGS|15|30|乌西雅 的儿子 约坦 第二十年， 以拉 的儿子 何细亚 背叛 利玛利 的儿子 比加 ，击杀他，篡了他的位。
2KGS|15|31|比加 其余的事，凡他所做的，看哪，都写在《以色列诸王记》上。
2KGS|15|32|利玛利 的儿子 以色列 王 比加 第二年， 犹大 王 乌西雅 的儿子 约坦 登基。
2KGS|15|33|他登基的时候年二十五岁，在 耶路撒冷 作王十六年。他母亲名叫 耶路沙 ，是 撒督 的女儿。
2KGS|15|34|约坦 行耶和华眼中看为正的事，效法他父亲 乌西雅 一切所行的。
2KGS|15|35|只是丘坛还没有废去，百姓仍在丘坛献祭烧香。 约坦 建了耶和华殿的 上门 。
2KGS|15|36|约坦 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|15|37|在那些日子，耶和华开始差 亚兰 王 利汛 和 利玛利 的儿子 比加 去攻击 犹大 。
2KGS|15|38|约坦 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 亚哈斯 接续他作王。
2KGS|16|1|利玛利 的儿子 比加 第十七年， 犹大 王 约坦 的儿子 亚哈斯 登基。
2KGS|16|2|他登基的时候年二十岁，在 耶路撒冷 作王十六年。他不像他祖先 大卫 行耶和华－他上帝眼中看为正的事，
2KGS|16|3|却行 以色列 诸王的道，又照着耶和华从 以色列 人面前赶出的外邦人所行可憎的事，使他的儿子经火，
2KGS|16|4|并在丘坛上、山冈上、各青翠树下献祭烧香。
2KGS|16|5|那时， 亚兰 王 利汛 和 利玛利 的儿子 以色列 王 比加 上来攻打 耶路撒冷 ，围困 亚哈斯 ，却不能打胜。
2KGS|16|6|当时 亚兰 王 利汛 收复 以拉他 回归 亚兰 ，把 犹大 人从 以拉他 赶出去。 以东 人来到 以拉他 ，住在那里，直到今日。
2KGS|16|7|亚哈斯 派使者到 亚述 王 提革拉．毗列色 那里，说：“我是你的仆人，你的儿子。现在 亚兰 王和 以色列 王攻击我，求你上来，救我脱离他们的手。”
2KGS|16|8|亚哈斯 将耶和华殿里和王宫府库里所有的金银都送给 亚述 王为礼物。
2KGS|16|9|亚述 王答应了他，上去攻打 大马士革 ，攻下了城，杀了 利汛 ，把居民掳到 吉珥 。
2KGS|16|10|亚哈斯 王到 大马士革 迎接 亚述 王 提革拉．毗列色 ，在 大马士革 看见一座坛。 亚哈斯 王把坛的规模和样式，以及作法的细节，送到 乌利亚 祭司那里。
2KGS|16|11|乌利亚 祭司照着 亚哈斯 王从 大马士革 所送来的一切，在 亚哈斯 王还未从 大马士革 回来之前，筑了一座坛。
2KGS|16|12|王从 大马士革 回来，看见坛，走近坛前，在坛上献祭。
2KGS|16|13|他烧燔祭和素祭，献浇酒祭，将平安祭牲的血洒在坛上。
2KGS|16|14|他移动耶和华面前的铜坛，从殿的前面，新坛和耶和华殿的中间，搬到新坛的北边。
2KGS|16|15|亚哈斯 王吩咐 乌利亚 祭司说：“早晨的燔祭、晚上的素祭，王的燔祭、素祭，国内众百姓的燔祭、素祭、浇酒祭都要烧在大坛上。燔祭牲和其他祭牲的血全都要洒在这坛上。至于铜坛，我要作求问之用。”
2KGS|16|16|乌利亚 祭司就照着 亚哈斯 王所吩咐的一切做了。
2KGS|16|17|亚哈斯 王把盆座四面的嵌边拆下来，把盆从座上挪下来，又将铜海从驮铜海的铜牛上搬下来，放在石板铺的地上。
2KGS|16|18|他为了 亚述 王的缘故，在耶和华的殿里移动 殿里为安息日所盖的遮棚 和王从外面进来的入口。
2KGS|16|19|亚哈斯 其余所做的事，不都写在《犹大列王记》上吗？
2KGS|16|20|亚哈斯 与他祖先同睡， 与他祖先同葬在 大卫城 ，他儿子 希西家 接续他作王。
2KGS|17|1|犹大 王 亚哈斯 第十二年， 以拉 的儿子 何细亚 在 撒玛利亚 登基作 以色列 王九年。
2KGS|17|2|他行耶和华眼中看为恶的事，只是不像在他以前的 以色列 诸王。
2KGS|17|3|亚述 王 撒缦以色 上来攻击 何细亚 ， 何细亚 就服事他，向他进贡。
2KGS|17|4|何细亚 背叛，派使者到 埃及 王 梭 那里 ，不照往年所行的向 亚述 王进贡。 亚述 王知道了，就逮捕他，把他囚在监里。
2KGS|17|5|亚述 王上来攻击 以色列 全地，上到 撒玛利亚 ，围困这城三年。
2KGS|17|6|何细亚 第九年， 亚述 王攻取了 撒玛利亚 ，把 以色列 人掳到 亚述 ，安置在 哈腊 与 歌散 的 哈博河 边，以及 玛代 人的城镇。
2KGS|17|7|这是因为 以色列 人得罪了那领他们出 埃及 地、脱离 埃及 王法老之手的耶和华－他们的上帝，去敬畏别神，
2KGS|17|8|随从耶和华在 以色列 人面前所赶出外邦人的风俗和 以色列 诸王所立的规条。
2KGS|17|9|以色列 人暗中行不正的事，违背耶和华－他们的上帝，在他们所有的城镇，从了望楼直到坚固城，建筑丘坛；
2KGS|17|10|在各高冈上、各青翠树下立柱像和 亚舍拉 ；
2KGS|17|11|在各丘坛上烧香，效法耶和华在他们面前赶出的外邦人所行的，又行恶事，惹耶和华发怒。
2KGS|17|12|他们事奉偶像，耶和华对他们说：“你们不可做这事。”
2KGS|17|13|耶和华藉众先知、先见劝戒 以色列 和 犹大 说：“当离开你们的恶行，谨守我的诫命律例，遵行我吩咐你们祖先、藉我仆人众先知所传给你们的一切律法。”
2KGS|17|14|他们却不听从，竟硬着颈项，像他们祖先一样，不信服耶和华－他们的上帝。
2KGS|17|15|他们厌弃他的律例，和他与他们列祖所立的约，以及他劝戒他们的话，去随从虚无的神明 ，自己成为虚妄，效法周围的列国，就是耶和华嘱咐他们不可效法的。
2KGS|17|16|他们离弃耶和华－他们上帝的一切诫命，为自己铸造了两个牛犊的像，立了 亚舍拉 ，敬拜天上的万象，事奉 巴力 ，
2KGS|17|17|使他们的儿女经火，占卜，行法术，出卖自己，行耶和华眼中看为恶的事，惹他发怒。
2KGS|17|18|所以耶和华向 以色列 大大发怒，从自己面前赶出他们，只剩下 犹大 一个支派。
2KGS|17|19|但是， 犹大 也不遵守耶和华－他们上帝的诫命，效法 以色列 所立的规条。
2KGS|17|20|耶和华就厌弃 以色列 所有的后裔，使他们受苦，把他们交在抢夺他们的人手中，直到他把他们从自己面前赶出去。
2KGS|17|21|当他使 以色列 从 大卫 家分离出来的时候，他们立 尼八 的儿子 耶罗波安 作王。 耶罗波安 引诱 以色列 不随从耶和华，陷入大罪中。
2KGS|17|22|以色列 人行 耶罗波安 所犯的一切罪，总不离开，
2KGS|17|23|以致耶和华把他们从自己面前赶出去，正如他藉他仆人众先知所说的。这样， 以色列 人从自己的土地被掳到 亚述 ，直到今日。
2KGS|17|24|亚述 王从 巴比伦 、 古他 、 亚瓦 、 哈马 和 西法瓦音 迁移人来，安置在 撒玛利亚 的城镇，代替 以色列 人；他们就占据了 撒玛利亚 ，住在城中。
2KGS|17|25|他们开始住在那里的时候，不敬畏耶和华，所以耶和华叫狮子进入他们中间，咬死了一些人。
2KGS|17|26|有人对 亚述 王说：“你所迁移安置在 撒玛利亚 城镇的各国的人，他们不知道那地之上帝的规矩，所以他叫狮子进入他们中间。看哪，狮子咬死了他们，因为他们不知道那地之上帝的规矩。”
2KGS|17|27|亚述 王吩咐说：“当派一个从那里掳来的祭司回去，叫他住在那里，将那地之上帝的规矩指导他们。”
2KGS|17|28|于是有一个从 撒玛利亚 掳去的祭司回来，住在 伯特利 ，教导他们怎样敬畏耶和华。
2KGS|17|29|然而，各国的人在所住的城里为自己制造神像，安置在 撒玛利亚 人所建有丘坛的庙中。
2KGS|17|30|巴比伦 人造 疏割．比讷 像； 古他 人造 匿甲 像； 哈马 人造 亚示玛 像；
2KGS|17|31|亚瓦 人造 匿哈 和 他珥他 像； 西法瓦音 人用火焚烧儿女，献给 西法瓦音 的神明 亚得米勒 和 亚拿米勒 。
2KGS|17|32|他们惧怕耶和华，却从他们中间立丘坛的祭司，在丘坛的庙中为他们献祭。
2KGS|17|33|他们惧怕耶和华，但又事奉自己的神明，从何邦迁来，就随从那里的风俗，
2KGS|17|34|直到如今仍照先前的风俗去行。 他们不敬畏耶和华，不遵守耶和华吩咐 雅各 后裔的律例、典章、律法、诫命； 雅各 就是从前耶和华起名叫 以色列 的。
2KGS|17|35|耶和华曾与他们立约，吩咐他们说：“不可敬畏别神，不可跪拜事奉它们，也不可向它们献祭。
2KGS|17|36|惟有那用大能和伸出来的膀臂领你们出 埃及 地的耶和华，你们当敬畏他，向他跪拜，向他献祭。
2KGS|17|37|他给你们写的律例、典章、律法、诫命，你们应当永远谨守遵行。你们不可敬畏别神。
2KGS|17|38|你们不可忘记我与你们所立的约，也不可敬畏别神。
2KGS|17|39|只要敬畏耶和华－你们的上帝，他必救你们脱离一切仇敌的手。”
2KGS|17|40|他们却不听从，仍照先前的风俗去行。
2KGS|17|41|这样，这些国家又惧怕耶和华，又事奉他们的偶像。他们子子孙孙也都照样行，效法他们的祖宗，直到今日。
2KGS|18|1|以拉 的儿子 以色列 王 何细亚 第三年， 犹大 王 亚哈斯 的儿子 希西家 登基。
2KGS|18|2|他登基的时候年二十五岁，在 耶路撒冷 作王二十九年。他母亲名叫 亚比 ，是 撒迦利雅 的女儿。
2KGS|18|3|希西家 行耶和华眼中看为正的事，效法他祖先 大卫 一切所行的。
2KGS|18|4|他废去丘坛，毁坏柱像，砍下 亚舍拉 ，打碎 摩西 所造的铜蛇，因为到那时 以色列 人仍向铜蛇烧香。人叫铜蛇为 尼忽士但 。
2KGS|18|5|希西家 倚靠耶和华－ 以色列 的上帝，在他之前和在他之后的 犹大 列王中没有一个像他一样的。
2KGS|18|6|因为他紧紧跟随耶和华，谨守耶和华所吩咐 摩西 的诫命，总不离开。
2KGS|18|7|耶和华与他同在，他无论往何处去尽都亨通。他背叛 亚述 王，不服事他。
2KGS|18|8|希西家 攻击 非利士 人，直到 迦萨 ，以及所属的领土，从了望楼到坚固城。
2KGS|18|9|希西家 王第四年，也就是 以拉 的儿子 以色列 王 何细亚 第七年， 亚述 王 撒缦以色 上来围困 撒玛利亚 。
2KGS|18|10|过了三年，他们攻取了城。 希西家 第六年， 以色列 王 何细亚 第九年， 撒玛利亚 被攻取了。
2KGS|18|11|亚述 王把 以色列 人掳到 亚述 ，安置在 哈腊 与 歌散 的 哈博河 边，以及 玛代 人的城镇。
2KGS|18|12|这是因为他们不听从耶和华－他们的上帝的话，违背了他的约；他们既不听从，也不遵行耶和华仆人 摩西 一切所吩咐的。
2KGS|18|13|希西家 王十四年， 亚述 王 西拿基立 上来攻击 犹大 的一切坚固的城，将城攻取。
2KGS|18|14|犹大 王 希西家 派人到 拉吉 ， 亚述 王那里，说：“我错了，求你撤退离开我；凡你罚我的，我必承当。”于是 亚述 王罚 犹大 王 希西家 三百他连得银子，三十他连得金子。
2KGS|18|15|希西家 把耶和华殿里和王宫府库里所有的银子都给了他。
2KGS|18|16|那时， 犹大 王 希西家 将耶和华殿门上的金子和他自己包在柱子上的金子都刮下来，给了 亚述 王。
2KGS|18|17|亚述 王从 拉吉 差遣元帅 、太监长 和将军 率领大军前往 耶路撒冷 ，到 希西家 王那里去。他们上来，到 耶路撒冷 。他们上来之后，站在 上池 的水沟旁，在往漂布地的大路上。
2KGS|18|18|他们呼叫王， 希勒家 的儿子 以利亚敬 宫廷总管， 舍伯那 书记和 亚萨 的儿子 约亚 史官就出来见他们。
2KGS|18|19|将军对他们说：“你们去告诉 希西家 ，大王 亚述 王如此说：‘你倚靠什么，让你如此自信满满？
2KGS|18|20|你说，你有打仗的计谋和能力，我看不过是空话。你到底倚靠谁，竟敢背叛我呢？
2KGS|18|21|现在，看哪，你自己所倚靠的 埃及 是那断裂的苇杖，人若倚靠这杖，它就刺进他的手，穿透它。 埃及 王法老向所有倚靠他的人都是这样。
2KGS|18|22|你们若对我说：我们倚靠耶和华－我们的上帝， 希西家 岂不是将上帝的丘坛和祭坛废去，并且吩咐 犹大 和 耶路撒冷 的人说：你们当在 耶路撒冷 这坛前敬拜吗？
2KGS|18|23|现在你与我主 亚述 王打赌，我给你两千匹马，看你能否派得出骑士来骑它们。
2KGS|18|24|若不然，怎能使我主臣仆中最小的一个军官转脸而逃呢？你难道要倚靠 埃及 的战车和骑兵吗？
2KGS|18|25|现在我上来攻击毁灭这地方，岂不是出于耶和华吗？耶和华吩咐我说，你上去攻击这地，毁灭它吧！’”
2KGS|18|26|希勒家 的儿子 以利亚敬 ， 舍伯那 和 约亚 对将军说：“求你用 亚兰 话对仆人说，因为我们听得懂；不要用 犹大 话对我们说，免得传到城墙上百姓的耳中。”
2KGS|18|27|将军对他们说：“我主差遣我来，岂是单对你和你的主人说这些话吗？不也是对这些坐在城墙上、要与你们一同吃自己粪、喝自己尿的人说的吗？”
2KGS|18|28|于是 亚述 将军站着，用 犹大 话大声喊着说：“你们当听大王 亚述 王的话，
2KGS|18|29|王如此说：‘你们不要被 希西家 欺哄了，因他不能救你们脱离我的手。
2KGS|18|30|不要听凭 希西家 说服你们倚靠耶和华，他说，耶和华必要拯救我们，这城必不交在 亚述 王的手中。’
2KGS|18|31|你们不要听 希西家 的话！因 亚述 王如此说：‘你们要与我讲和，出来投降我，各人就可以吃自己葡萄树和无花果树的果子，喝自己井里的水，
2KGS|18|32|等我来领你们到一个地方，与你们本地一样，就是有五谷和新酒之地，有粮食和葡萄园之地，有橄榄树和蜂蜜之地，好使你们存活，不至于死。不要听 希西家 的话，因为他误导你们说：耶和华必拯救我们。
2KGS|18|33|列国的神明有哪一个曾救它本国脱离 亚述 王的手呢？
2KGS|18|34|哈马 、 亚珥拔 的神明在哪里呢？ 西法瓦音 、 希拿 、 以瓦 的神明在哪里呢？ 它们曾救 撒玛利亚 脱离我的手吗？
2KGS|18|35|这些国的神明有谁曾救自己的国脱离我的手呢？难道耶和华能救 耶路撒冷 脱离我的手吗？’”
2KGS|18|36|百姓静默不言，一句不答，因为 希西家 王曾吩咐说：“不要回答他。”
2KGS|18|37|当下， 希勒家 的儿子 以利亚敬 宫廷总管、 舍伯那 书记和 亚萨 的儿子 约亚 史官，都撕裂衣服，来到 希西家 那里，将 亚述 将军的话告诉他。
2KGS|19|1|希西家 王听见了，就撕裂衣服，披上麻布，进了耶和华的殿。
2KGS|19|2|他差遣 以利亚敬 宫廷总管和 舍伯那 书记，并祭司中年长的，都披上麻布，到 亚摩斯 的儿子 以赛亚 先知那里去。
2KGS|19|3|他们对他说：“ 希西家 如此说：‘今日是急难、惩罚、凌辱的日子，就如婴孩快要出生，却没有力气生产。
2KGS|19|4|或许耶和华－你的上帝听见 亚述 将军一切的话，就是他主人 亚述 王差他来辱骂永生上帝的话，耶和华－你的上帝就斥责所听见的这些话。求你为幸存的余民扬声祷告。’”
2KGS|19|5|希西家 王的臣仆来到 以赛亚 那里的时候，
2KGS|19|6|以赛亚 对他们说：“要对你们的主人这样说，耶和华如此说：‘你听见 亚述 王的仆人亵渎我的话，不要惧怕。
2KGS|19|7|看哪，我必惊动他的心 ，他要听见风声就归回本地，在那里我必使他倒在刀下。’”
2KGS|19|8|亚述 将军听见 亚述 王已拔营离开 拉吉 ，就启程返回，正遇见 亚述 王去攻打 立拿 。
2KGS|19|9|亚述 王听见有人谈论 古实 王 特哈加 说：“看哪，他出来要与你争战。”于是 亚述 王又差使者去见 希西家 ，说：
2KGS|19|10|“你们要对 犹大 王 希西家 如此说：‘不要听你所倚靠的上帝欺哄你说： 耶路撒冷 必不交在 亚述 王的手中。
2KGS|19|11|看哪，你总听说 亚述 诸王向列国所行的是尽行灭绝，难道你能幸免吗？
2KGS|19|12|我祖先所毁灭的，就是 歌散 、 哈兰 、 利色 和 提．拉撒 的 伊甸 人；这些国的神明何曾拯救他们呢？
2KGS|19|13|哈马 的王， 亚珥拔 的王， 西法瓦音城 的王， 希拿 和 以瓦 的王，都在哪里呢？’”
2KGS|19|14|希西家 从使者手里接过书信，读完了，就上耶和华的殿，在耶和华面前展开书信。
2KGS|19|15|希西家 向耶和华祷告说：“坐在基路伯之上耶和华－ 以色列 的上帝啊，你，惟有你是地上万国的上帝，你创造了天和地。
2KGS|19|16|耶和华啊，求你侧耳而听；耶和华啊，求你睁眼而看，听 西拿基立 差遣使者辱骂永生上帝的话。
2KGS|19|17|耶和华啊， 亚述 诸王果然使列国和列国之地变为荒芜，
2KGS|19|18|将列国的神像扔在火里，因为它们不是上帝，是人手所造的，是木头、石头，所以被灭绝了。
2KGS|19|19|耶和华－我们的上帝啊，现在求你救我们脱离 亚述 王的手，使地上万国都知道惟独你－耶和华是上帝！”
2KGS|19|20|亚摩斯 的儿子 以赛亚 差人去见 希西家 ，说：“耶和华－ 以色列 的上帝如此说：你因 亚述 王 西拿基立 的事向我祈求，我已听见了。
2KGS|19|21|耶和华论他这样说： ‘少女 锡安 藐视你，嘲笑你； 耶路撒冷 向你摇头。
2KGS|19|22|‘你辱骂谁，亵渎谁， 扬起声来，高举眼目攻击谁呢？ 你攻击的是 以色列 的圣者。
2KGS|19|23|你藉你的使者辱骂主说： 我率领许多战车登上高山， 到 黎巴嫩 的顶端； 我要砍伐其中高大的香柏树 和上好的松树； 我必进到极遥远的住所， 进入最茂盛的森林里。
2KGS|19|24|我已经在外邦挖井喝水； 我必用脚掌踏干 埃及 一切的河流。
2KGS|19|25|‘你岂没有听见 我早先所定、古时所立、现今实现的事吗？ 就是让你去毁坏坚固的城镇，使它们变为废墟；
2KGS|19|26|城里的居民力量微小， 他们惊惶羞愧； 像野草，像青菜， 如房顶上的草， 又如未长成而枯干的禾稼。
2KGS|19|27|‘你坐下，你出去，你进来， 你向我发烈怒，我都知道。
2KGS|19|28|因你向我发烈怒， 你的狂傲上达我耳中， 我要用钩子钩住你的鼻子， 将嚼环放在你口里， 使你从原路转回去。’
2KGS|19|29|“这是给你的预兆：你们今年要吃野生的，明年也要吃自长的；后年，你们就要耕种收割，栽葡萄园，吃其中的果子。
2KGS|19|30|犹大 家所逃脱剩余的，仍要往下扎根，向上结果。
2KGS|19|31|必有剩余的民从 耶路撒冷 而出，有逃脱的人从 锡安山 而来。万军之耶和华的热心必成就这事。
2KGS|19|32|“所以耶和华论 亚述 王如此说：他必不得来到这城，也不在这里射箭，不得拿盾牌到城前，也不建土堆攻城。
2KGS|19|33|他从哪条路来，必从那条路回去，必不得来到这城。这是耶和华说的。
2KGS|19|34|因我为自己的缘故，又为我仆人 大卫 的缘故，必保护拯救这城。”
2KGS|19|35|当夜，耶和华的使者出去，在 亚述 营中杀了十八万五千人。清早有人起来，看哪，都是死尸。
2KGS|19|36|亚述 王 西拿基立 就拔营回去，住在 尼尼微 。
2KGS|19|37|一日，他在他的神明 尼斯洛 庙里叩拜，他儿子 亚得米勒 和 沙利色 用刀杀了他，然后逃到 亚拉腊 地；他儿子 以撒．哈顿 接续他作王。
2KGS|20|1|那些日子， 希西家 病得要死， 亚摩斯 的儿子 以赛亚 先知来见他，对他说：“耶和华如此说：‘你当留遗嘱给你的家，因为你必死，不能活了。’”
2KGS|20|2|希西家 转脸朝墙，向耶和华祷告说：
2KGS|20|3|“耶和华啊，求你记念我在你面前怎样存完全的心，按诚实行事，又做你眼中看为善的事。” 希西家 就痛哭。
2KGS|20|4|以赛亚 出来，还没有离开中院，耶和华的话就临到他，说：
2KGS|20|5|“你回去告诉我百姓的君王 希西家 说：耶和华－你祖先 大卫 的上帝如此说：‘我听见了你的祷告，看见了你的眼泪。看哪，我必医治你；到第三日，你必上到耶和华的殿。
2KGS|20|6|我必加添你十五年的寿数，并且我要救你和这城脱离 亚述 王的手。我为自己和我仆人 大卫 的缘故，必保护这城。’”
2KGS|20|7|以赛亚 说：“取一块无花果饼来。”人就取了来，贴在疮上，王就痊愈了。
2KGS|20|8|希西家 对 以赛亚 说：“耶和华必医治我，到第三日我能上耶和华的殿，有什么预兆呢？”
2KGS|20|9|以赛亚 说：“耶和华必成就他所说的这话。这是耶和华给你的预兆：你要日影向前进十度呢？或是要往后退十度呢？”
2KGS|20|10|希西家 说：“日影向前进十度容易；不，让日影往后退十度吧。”
2KGS|20|11|以赛亚 先知求告耶和华，耶和华就使 亚哈斯 日晷上照下来的日影，往后退了十度。
2KGS|20|12|那时， 巴拉但 的儿子， 巴比伦 王 米罗达．巴拉但 听见 希西家 生病了，就送书信和礼物给他。
2KGS|20|13|希西家 听使者的话 ，就将自己一切宝库里的金子、银子、香料、贵重的膏油和他军械库里的兵器，以及他所有的财宝，都给他们看；在他家中和全国之内， 希西家 没有一样东西不给他们看的。
2KGS|20|14|于是 以赛亚 先知到 希西家 王那里去，对他说：“这些人说了些什么？他们从哪里来见你？” 希西家 说：“他们从远方的 巴比伦 来。”
2KGS|20|15|以赛亚 说：“他们在你家里看见了什么？” 希西家 说：“凡我家中所有的，他们都看见了；我财宝中没有一样东西不给他们看的。”
2KGS|20|16|以赛亚 对 希西家 说：“你要听耶和华的话：
2KGS|20|17|耶和华说：‘看哪，日子将到，凡你家里所有的，并你祖先积蓄到如今的一切，都要被掳到 巴比伦 去，不留下一样；
2KGS|20|18|从你本身所生的孩子，其中必有被掳到 巴比伦 王宫当太监的。’”
2KGS|20|19|希西家 对 以赛亚 说：“你所说耶和华的话甚好。”因为他想：“在我有生之年岂不是有太平和安稳吗？”
2KGS|20|20|希西家 其余的事和他一切英勇的事迹，他怎样造池、挖沟、引水入城，不都写在《犹大列王记》上吗？
2KGS|20|21|希西家 与他祖先同睡，他儿子 玛拿西 接续他作王。
2KGS|21|1|玛拿西 登基的时候年十二岁，在 耶路撒冷 作王五十五年。他母亲名叫 协西巴 。
2KGS|21|2|玛拿西 行耶和华眼中看为恶的事，效法耶和华在 以色列 人面前赶出的列国那些可憎的事。
2KGS|21|3|他重新建筑他父亲 希西家 所毁坏的丘坛，又为 巴力 筑坛，造 亚舍拉 ，效法 以色列 王 亚哈 所行的，敬拜天上的万象，事奉它们。
2KGS|21|4|他在耶和华殿中筑坛，耶和华曾指着这殿说：“我必立我的名在 耶路撒冷 。”
2KGS|21|5|他在耶和华殿的两个院子为天上的万象筑坛，
2KGS|21|6|并使他的儿子经火，又观星象，行法术，求问招魂的和行巫术的，多行耶和华眼中看为恶的事，惹他发怒。
2KGS|21|7|他又把自己所造的 亚舍拉 雕像立在殿内，耶和华曾对 大卫 和他儿子 所罗门 说：“我在 以色列 众支派中所选择的 耶路撒冷 和这殿，必立我的名，直到永远。
2KGS|21|8|只要 以色列 人谨守遵行我一切所吩咐的和我仆人 摩西 所吩咐的一切律法，我就不再使他们的脚挪移，离开我所赐给他们列祖之土地。”
2KGS|21|9|他们却不听从，并且 玛拿西 引诱他们行恶，比耶和华在 以色列 人面前所灭的列国更严重。
2KGS|21|10|耶和华藉他仆人众先知说：
2KGS|21|11|“因 犹大 王 玛拿西 行这些可憎的恶事，比先前 亚摩利 人所行的一切更坏，使 犹大 人拜偶像，陷入罪里，
2KGS|21|12|所以耶和华－ 以色列 的上帝如此说：看哪，我必降祸于 耶路撒冷 和 犹大 ，凡听见的人都必双耳齐鸣。
2KGS|21|13|我必用量 撒玛利亚 的准绳和 亚哈 家的铅垂线拉在 耶路撒冷 之上；我必擦拭 耶路撒冷 ，如人擦盘子，把盘子翻过来。
2KGS|21|14|我必撇弃我产业中的余民，把他们交在仇敌手中，使他们成为所有仇敌的掳物和掠物，
2KGS|21|15|因为自从他们的祖先出 埃及 的那日直到今日，他们常行我眼中看为恶的事，惹我发怒。”
2KGS|21|16|玛拿西 行耶和华眼中看为恶的事，使 犹大 陷入罪里，又流许多无辜人的血，直到这血充满了 耶路撒冷 ，从这边到那边。
2KGS|21|17|玛拿西 其余的事，凡他所做的和他所犯的罪，不都写在《犹大列王记》上吗？
2KGS|21|18|玛拿西 与他祖先同睡，葬在自己王宫的园子， 乌撒 园里，他儿子 亚们 接续他作王。
2KGS|21|19|亚们 登基的时候年二十二岁，在 耶路撒冷 作王二年。他母亲名叫 米舒利密 ，是 约提巴 人 哈鲁斯 的女儿。
2KGS|21|20|亚们 行耶和华眼中看为恶的事，效法他父亲 玛拿西 所行的。
2KGS|21|21|他行他父亲一切所行的道，事奉他父亲所事奉的偶像，敬拜它们，
2KGS|21|22|离弃耶和华－他列祖的上帝，不遵行耶和华的道。
2KGS|21|23|亚们 的臣仆背叛他，在宫里杀了王。
2KGS|21|24|但这地的百姓杀了所有背叛 亚们 王的人；这地的百姓立他儿子 约西亚 接续他作王。
2KGS|21|25|亚们 其余所做的事，不都写在《犹大列王记》上吗？
2KGS|21|26|亚们 葬在 乌撒 园内自己的坟墓里，他儿子 约西亚 接续他作王。
2KGS|22|1|约西亚 登基的时候年八岁，在 耶路撒冷 作王三十一年。他母亲名叫 耶底大 ，是 波斯加 人 亚大雅 的女儿。
2KGS|22|2|约西亚 行耶和华眼中看为正的事，行他祖先 大卫 一切所行的道，不偏左右。
2KGS|22|3|约西亚 王十八年，王派 米书兰 的孙子， 亚萨利雅 的儿子 沙番 书记上耶和华殿去，说：
2KGS|22|4|“你上到 希勒家 大祭司那里，请他把奉献到耶和华殿的银子，就是门口的守卫从百姓中收来的银子，结算清楚，
2KGS|22|5|交在管理耶和华殿督工的手里，由他们支付给在耶和华殿里做工的人，好修理殿的破坏之处，
2KGS|22|6|就是木匠、工人和瓦匠，又买木料和凿成的石头，来整修殿宇。
2KGS|22|7|但他们不用跟这些经手接受银子的人算帐，因为这些人办事诚实。”
2KGS|22|8|希勒家 大祭司对 沙番 书记说：“我在耶和华殿里发现了律法书。” 希勒家 把书递给 沙番 ， 沙番 就读了。
2KGS|22|9|沙番 书记到王那里，把这事回覆王说：“你的仆人已把殿里所发现的银子倒出来，交在管理耶和华殿督工的手里了。”
2KGS|22|10|沙番 书记又向王报告说：“ 希勒家 祭司递给我一卷书。” 沙番 就在王面前朗读那书。
2KGS|22|11|王听见律法书上的话，就撕裂衣服。
2KGS|22|12|王吩咐 希勒家 祭司与 沙番 的儿子 亚希甘 、 米该亚 的儿子 亚革波 、 沙番 书记和王的臣仆 亚撒雅 ，说：
2KGS|22|13|“你们去，以所发现这书上的话，为我、为百姓、为全 犹大 求问耶和华；因为我们祖先没有听从这书上的话，没有遵照一切所写有关我们的 去行，耶和华就向我们大发烈怒。”
2KGS|22|14|于是， 希勒家 祭司和 亚希甘 、 亚革波 、 沙番 、 亚撒雅 都去见 户勒大 女先知，她是掌管礼服的 沙龙 的妻子； 沙龙 是 哈珥哈斯 的孙子， 特瓦 的儿子。 户勒大 住在 耶路撒冷 第二区。他们向她请教。
2KGS|22|15|她对他们说：“耶和华－ 以色列 的上帝如此说：‘你们可以回覆那派你们来见我的人说，
2KGS|22|16|耶和华如此说：看哪，我必照着 犹大 王所读那书上的一切话，降祸于这地方和其上的居民。
2KGS|22|17|因为他们离弃我，向别神烧香，用他们手所做的一切惹我发怒，所以我的愤怒必向这地方发作，总不止息。’
2KGS|22|18|然而，派你们来求问耶和华的 犹大 王，你们要这样回覆他：‘耶和华－ 以色列 的上帝如此说：至于你所听见的话，
2KGS|22|19|就是听见我指着这地方和其上的居民说，要使这地方变为荒芜、百姓受诅咒的话，你的心就软化，在耶和华面前谦卑下来，撕裂衣服，向我哭泣，因此我应允你。这是耶和华说的。
2KGS|22|20|因此，看哪，我必使你归到你祖先那里，平安地进入坟墓；我要降于这地方的一切灾祸，你不会亲眼看见。’”他们就去把这话回覆王。
2KGS|23|1|王派人召集 犹大 和 耶路撒冷 的众长老来。
2KGS|23|2|王和 犹大 众人、 耶路撒冷 的居民、祭司、先知，以及所有的百姓，无论大小，都一同上到耶和华的殿去；王把耶和华殿里所发现的约书上一切的话读给他们听。
2KGS|23|3|王站在柱子旁边，在耶和华面前立约，要尽心尽性跟从耶和华，遵守他的诫命、法度、律例，实行这书上所写这约的话。全体百姓都愿遵守所立的约。
2KGS|23|4|王吩咐 希勒家 大祭司和副祭司，以及把守殿门的，把那些为 巴力 和 亚舍拉 ，以及天上万象所造的器皿，都从耶和华殿里搬出来，在 耶路撒冷 外 汲沦 的田间烧了，把灰拿到 伯特利 去。
2KGS|23|5|从前 犹大 列王所立拜偶像的祭司，在 犹大 城镇的丘坛和 耶路撒冷 周围烧香，现在王都废去，他们是向 巴力 和日、月、行星，以及天上万象烧香的人。
2KGS|23|6|他把 亚舍拉 从耶和华殿里搬到 耶路撒冷 外的 汲沦溪 ，在 汲沦溪 边焚烧，打碎成灰，把灰撒在平民的坟上。
2KGS|23|7|他又拆毁耶和华殿里男的庙妓的屋子，就是妇女在那里为 亚舍拉 编织衣服的屋子。
2KGS|23|8|他从 犹大 的城镇将众祭司带来，从 迦巴 直到 别是巴 ，玷污祭司烧香的丘坛。他又拆毁城门旁的丘坛，这丘坛是在 约书亚 市长的城门前，在人进城门的左边。
2KGS|23|9|只是丘坛的祭司不登 耶路撒冷 耶和华的坛，仅在他们弟兄中间吃无酵饼。
2KGS|23|10|他又玷污 欣嫩子谷 的 陀斐特 ，不许人在那里使儿女经火献给 摩洛 。
2KGS|23|11|他把在耶和华殿门旁、靠近 拿单．米勒 官员走廊的屋子， 犹大 列王献给太阳的马废去，且用火焚烧献给太阳的战车。
2KGS|23|12|犹大 列王在 亚哈斯 楼房顶上所筑的坛和 玛拿西 在耶和华殿两院中所筑的坛，王都拆毁，从那里移走 ，把灰倒在 汲沦溪 中。
2KGS|23|13|从前 以色列 王 所罗门 在 耶路撒冷 东边、 邪僻山 南边为 西顿 人可憎的 亚斯她录 、 摩押 人可憎的 基抹 、 亚扪 人可憎的 米勒公 所筑的丘坛，王都玷污了，
2KGS|23|14|又打碎柱像，砍下 亚舍拉 ，用人的骨头填满那地方。
2KGS|23|15|此外，在 伯特利 丘坛的坛，就是 尼八 的儿子 耶罗波安 所筑、使 以色列 人陷入罪里的，他也把这坛和丘坛都拆毁了，又焚烧丘坛 ，打碎成灰，并焚烧了 亚舍拉 。
2KGS|23|16|约西亚 转头，看见山上的坟墓，就派人取出坟墓里的骸骨，烧在坛上，玷污了坛，正如从前 耶罗波安 在节期中站在坛旁时，耶和华藉神人所宣告的话。 约西亚 转头看见了宣告这些话的神人的坟墓。
2KGS|23|17|他说：“我看见的这碑是什么呢？”那城里的人对他说：“这是神人的坟墓，他从 犹大 来，宣告了王向 伯特利 的坛所做的这些事。”
2KGS|23|18|约西亚 说：“让他安息吧！不要挪移他的骸骨。”他们就保存了他的骸骨和从 撒玛利亚 来的那先知的骸骨。
2KGS|23|19|从前 以色列 诸王在 撒玛利亚 的城镇所建一切惹动怒气的丘坛的庙， 约西亚 也都废去了，正如他在 伯特利 所做的。
2KGS|23|20|他又把在那里所有丘坛的祭司都杀在坛上，并在坛上烧人的骨头。于是他回 耶路撒冷 去了。
2KGS|23|21|王吩咐众百姓说：“你们当照这约书上所写的，向耶和华－你们的上帝守逾越节。”
2KGS|23|22|自从士师治理 以色列 ，到 以色列 诸王、 犹大 列王在位的一切日子，从来没有守过这样的逾越节，
2KGS|23|23|只有在 约西亚 王十八年，才在 耶路撒冷 向耶和华守这逾越节。
2KGS|23|24|此外，在 犹大 地和 耶路撒冷 所见那些招魂的、行巫术的，家中的神像和偶像，以及一切可憎之物， 约西亚 尽都除掉，实行了 希勒家 祭司在耶和华殿里所发现的律法书上所写的话。
2KGS|23|25|在 约西亚 以前，没有王像他尽心、尽性、尽力地归向耶和华，遵行 摩西 的一切律法；在他以后，也没有兴起一个王像他。
2KGS|23|26|然而，耶和华向 犹大 所发猛烈的怒气仍不止息，因为 玛拿西 种种的恶事激怒了他。
2KGS|23|27|耶和华说：“我也必将 犹大 从我面前赶出，如同赶出 以色列 一样。我必撇弃我从前所选择的这城 耶路撒冷 和我所说我的名必留在那里的殿。”
2KGS|23|28|约西亚 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|23|29|约西亚 的日子， 埃及 王法老 尼哥 上到 幼发拉底河 ，到 亚述 王那里； 约西亚 王去迎击他。 埃及 王在 米吉多 看见 约西亚 ，就杀了他。
2KGS|23|30|他的臣仆用车把他的尸体从 米吉多 送到 耶路撒冷 ，葬在他自己的坟墓里。这地的百姓选 约西亚 的儿子 约哈斯 ，膏立他，接续他父亲作王。
2KGS|23|31|约哈斯 登基的时候年二十三岁，在 耶路撒冷 作王三个月。他母亲名叫 哈慕她 ，是 立拿 人 耶利米 的女儿。
2KGS|23|32|约哈斯 行耶和华眼中看为恶的事，效法他祖先一切所行的。
2KGS|23|33|法老 尼哥 把 约哈斯 监禁在 哈马 地的 利比拉 ，不许他在 耶路撒冷 作王 ，又罚这地一百他连得银子，一他连得金子。
2KGS|23|34|法老 尼哥 立 约西亚 的儿子 以利亚敬 接续他父亲 约西亚 作王，给他改名叫 约雅敬 ，却把 约哈斯 带到 埃及 ，他就死在那里。
2KGS|23|35|约雅敬 进贡金银给法老，照着法老的指示在这地征收银子，向这地的百姓按各人的能力索取金银，要送给法老 尼哥 。
2KGS|23|36|约雅敬 登基的时候年二十五岁，在 耶路撒冷 作王十一年。他母亲名叫 西布大 ，是 鲁玛 人 毗大雅 的女儿。
2KGS|23|37|约雅敬 行耶和华眼中看为恶的事，效法他祖先一切所行的。
2KGS|24|1|约雅敬 的日子， 巴比伦 王 尼布甲尼撒 上来； 约雅敬 服事他三年，以后又背叛他。
2KGS|24|2|耶和华派 迦勒底 、 亚兰 、 摩押 和 亚扪 人的军队来攻击 约雅敬 ；耶和华派他们来攻击 犹大 ，要毁灭它，正如耶和华藉他仆人众先知所说的话。
2KGS|24|3|这事临到 犹大 ，诚然是出于耶和华的命令 ，要把 犹大 从自己面前赶出去，是因 玛拿西 所犯的一切罪，
2KGS|24|4|又因他流无辜人的血，使无辜人的血充满 耶路撒冷 ；耶和华不愿赦免。
2KGS|24|5|约雅敬 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|24|6|约雅敬 与他祖先同睡，他儿子 约雅斤 接续他作王。
2KGS|24|7|埃及 王不再从他的国出征，因为 巴比伦 王把 埃及 王所管之地，从 埃及 溪谷直到 幼发拉底河 都夺去了。
2KGS|24|8|约雅斤 登基的时候年十八岁，在 耶路撒冷 作王三个月。他母亲名叫 尼护施她 ，是 耶路撒冷 人 以利拿单 的女儿。
2KGS|24|9|约雅斤 行耶和华眼中看为恶的事，效法他父亲一切所行的。
2KGS|24|10|那时， 巴比伦 王 尼布甲尼撒 的军兵上到 耶路撒冷 ，城被围困。
2KGS|24|11|当他的军兵围困城的时候， 巴比伦 王 尼布甲尼撒 亲自来到 耶路撒冷 。
2KGS|24|12|犹大 王 约雅斤 和他母亲、臣仆、王子、官员一同出来，向 巴比伦 王投降。 巴比伦 王俘掳了他，那时是 巴比伦 王第八年。
2KGS|24|13|巴比伦 王把耶和华殿里和王宫里一切的宝物从那里拿走，又把 以色列 王 所罗门 所造耶和华殿里一切的金器都毁坏了，正如耶和华所说的。
2KGS|24|14|他把全 耶路撒冷 众领袖和所有大能的勇士，共一万人，连同所有的木匠和铁匠都掳了去，只留下这地最贫穷的百姓。
2KGS|24|15|他把 约雅斤 和他的母亲、后妃、官员，以及这地的贵族，都从 耶路撒冷 掳到 巴比伦 去了，
2KGS|24|16|又把所有的勇士七千人，木匠和铁匠一千人，全是能上阵的勇士，都掳到 巴比伦 去了。
2KGS|24|17|巴比伦 王立 约雅斤 的叔父 玛探雅 取代他作王，给 玛探雅 改名叫 西底家 。
2KGS|24|18|西底家 登基的时候年二十一岁，在 耶路撒冷 作王十一年。他母亲名叫 哈慕她 ，是 立拿 人 耶利米 的女儿。
2KGS|24|19|西底家 行耶和华眼中看为恶的事，正如 约雅敬 一切所行的。
2KGS|24|20|因此，耶和华向 耶路撒冷 和 犹大 发怒，以致把他们从自己面前赶出去。 西底家 背叛 巴比伦 王。
2KGS|25|1|西底家 作王第九年十月初十， 巴比伦 王 尼布甲尼撒 率领全军前来攻击 耶路撒冷 ，对城安营，四围筑堡垒攻城。
2KGS|25|2|城被围困，直到 西底家 王十一年。
2KGS|25|3|四月初九，城里的饥荒非常严重，当地的百姓都没有粮食。
2KGS|25|4|城被攻破，士兵全都在夜间从靠近王的花园、两城墙中间的门逃跑。 迦勒底 人正在四围攻城，王就往 亚拉巴 逃去。
2KGS|25|5|迦勒底 的军队追赶王，在 耶利哥 的平原追上他；他的全军都离开他溃散了。
2KGS|25|6|迦勒底 人就拿住王，带他到 利比拉 的 巴比伦 王那里；他们就判他的罪。
2KGS|25|7|他们在 西底家 眼前杀了他的儿女，挖了 西底家 的眼睛，用铜链锁着他，带到 巴比伦 去。
2KGS|25|8|巴比伦 王 尼布甲尼撒 十九年五月初七， 巴比伦 王的臣仆 尼布撒拉旦 护卫长进入 耶路撒冷 ，
2KGS|25|9|他焚烧了耶和华的殿、王宫和 耶路撒冷 一切的房屋；用火焚烧所有大户人家的房屋。
2KGS|25|10|跟从护卫长的 迦勒底 全军拆毁了 耶路撒冷 四围的城墙。
2KGS|25|11|那时 尼布撒拉旦 护卫长将城里剩下的百姓和那些投降 巴比伦 王的人，以及其余的众人，都掳去了。
2KGS|25|12|但护卫长留下一些当地最穷的人，叫他们修整葡萄园，耕种田地。
2KGS|25|13|耶和华殿的铜柱并殿内的盆座和铜海， 迦勒底 人都打碎了，把那些铜运到 巴比伦 去。
2KGS|25|14|他们又带走锅、铲子、钳子、勺子和供奉用的一切铜器；
2KGS|25|15|火盆和碗，无论金的银的，护卫长都带走了；
2KGS|25|16|还有 所罗门 为耶和华殿所造的两根柱子、一个铜海和盆座，这一切器皿的铜多得无法可秤。
2KGS|25|17|这一根柱子高十八肘，柱上有铜顶，铜顶高三肘；铜顶的周围有网子和石榴，也都是铜的。第二根柱子与此相同，也有网子。
2KGS|25|18|护卫长拿住 西莱雅 大祭司、 西番亚 副祭司和门口的三个守卫，
2KGS|25|19|又从城中拿住一个管理士兵的官 ，并在城里所找到王面前的五个亲信，和召募当地百姓之将军的书记官，以及在城中找到的六十个当地百姓。
2KGS|25|20|尼布撒拉旦 护卫长把这些人带到 利比拉 的 巴比伦 王那里。
2KGS|25|21|巴比伦 王击杀他们，在 哈马 地的 利比拉 把他们处死。这样， 犹大 人就被掳去离开本地。
2KGS|25|22|至于 犹大 地剩下的百姓，就是 巴比伦 王 尼布甲尼撒 所留下的， 巴比伦 王立了 沙番 的孙子， 亚希甘 的儿子 基大利 作他们的省长。
2KGS|25|23|所有的军官和属他们的人听见 巴比伦 王立了 基大利 作省长， 尼探雅 的儿子 以实玛利 、 加利亚 的儿子 约哈难 、 尼陀法 人 单户蔑 的儿子 西莱雅 、 玛迦 人的儿子 雅撒尼亚 ，和属他们的人，都来到 米斯巴 的 基大利 那里。
2KGS|25|24|基大利 向他们和属他们的人起誓说：“你们不必惧怕 迦勒底 臣仆，只管住在这地，服事 巴比伦 王，就可以得福。”
2KGS|25|25|七月中，王室后裔 以利沙玛 的孙子， 尼探雅 的儿子 以实玛利 带着十个人来，击杀了 基大利 和同他在 米斯巴 的 犹大 人与 迦勒底 人，把他们杀死。
2KGS|25|26|于是众人，无论大小，连同军官，因为惧怕 迦勒底 人，都起身逃到 埃及 去了。
2KGS|25|27|巴比伦 王 以未．米罗达 作王的元年，就是 犹大 王 约雅斤 被掳后三十七年，十二月二十七日，他使 犹大 王 约雅斤 抬起头来，提他出监，
2KGS|25|28|对他说好话，使他的位高过与他一同被掳在 巴比伦 众王的位；
2KGS|25|29|又给他脱了囚服，使他终身常在 巴比伦 王面前吃饭。
2KGS|25|30|王赐给他日常需用的食物，每日一份，终身都是这样。
