NUM|1|1|І Господь промовляв до Мойсея в Сінайській пустині в скинії заповіту першого дня другого місяця, другого року від виходу їх з єгипетського краю, говорячи:
NUM|1|2|Перелічіть усю громаду Ізраїлевих синів за родами їхніми, за домами їхніх батьків числом усіх чоловічої статі за їх головами,
NUM|1|3|від віку двадцяти літ і вище, кожного, хто здатний до війська в Ізраїлі, за військовими відділами їхніми перелічіть їх ти та Аарон.
NUM|1|4|А з вами будуть по одному мужеві для племени; той муж голова дому батьків своїх він.
NUM|1|5|А оце ймення тих мужів, що стануть із вами: для Рувима Еліцур, син Шедеурів;
NUM|1|6|для Симеона Шелуміїл, син Цурішаддаїв;
NUM|1|7|для Юди Нахшон, син Аммінадавів;
NUM|1|8|для Іссахара Натанаїл, син Цуарів;
NUM|1|9|для Завулона Елів, син Хелонів;
NUM|1|10|для Йосипових синів, від Єфрема Елішама, син Аммігудів; від Манасії Гамаліїл, син Педацурів;
NUM|1|11|для Веніямина Авідан, син Ґід'оніїв;
NUM|1|12|для Дана Ахіезер, син Аммішаддаїв;
NUM|1|13|для Асира Паґ'іїл, син Охранів;
NUM|1|14|для Ґада Ел'ясаф, син Деуїлів;
NUM|1|15|для Нефталима Ахіра, син Енанів.
NUM|1|16|Оце покликані громади, начальники племен їхніх батьків. Вони голови тисяч Ізраїлевих.
NUM|1|17|І взяв Мойсей та Аарон тих мужів, що були названі пойменно,
NUM|1|18|і вони зібрали всю ту громаду першого дня другого місяця. І вони виявили родоводи свої за домами їхніх батьків числом імен від віку двадцяти літ і вище, за головами їх,
NUM|1|19|як Господь наказав був Мойсеєві. І він перелічив їх у Сінайській пустині.
NUM|1|20|І було синів Рувима, перворідного Ізраїлевого, їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен за головами їх, усіх чоловічої статі від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|21|перелічені їхні від Рувимового племені сорок і шість тисяч і п'ятсот.
NUM|1|22|У Симеонових синів їхніх нащадків за їхніми родами, за домами їхніх батьків перелік їх числом імен за головами їхніми, усі чоловічої статі від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|23|перелічені їхні від Симеонового племени п'ятдесят і дев'ять тисяч і триста.
NUM|1|24|У Ґадових синів їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|25|перелічені їхні від Ґадового племени сорок і п'ять тисяч і шістсот і п'ятдесят.
NUM|1|26|У Юдових синів їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|27|перелічені їхні від Юдового племени сімдесят і чотири тисячі й шістсот.
NUM|1|28|У Іссахарових синів їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|29|перелічені їхні від Іссахарового племени п'ятдесят і чотири тисячі й чотириста.
NUM|1|30|У Завулонових синів їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|31|перелічені їхні від Завулонового племени п'ятдесят і сім тисяч і чотириста.
NUM|1|32|У Йосипових синів: у Єфремових синів їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|33|перелічені їхні від Єфремового племени сорок тисяч і п'ятсот.
NUM|1|34|У синів Манасії їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|35|перелічені їхні від племени Манасіїного тридцять і дві тисячі й двісті.
NUM|1|36|У Веніяминових синів їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|37|перелічені їхні від Веніяминового племени тридцять і п'ять тисяч і чотириста.
NUM|1|38|У Данових синів їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|39|перелічені їхні від Данового племени шістдесят і дві тисячі й сімсот.
NUM|1|40|У Асирових синів їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|41|перелічені їхні від Асирового племени, сорок і одна тисяча й п'ятсот.
NUM|1|42|У синів Нефталимових їхніх нащадків за їхніми родами, за домами їхніх батьків числом імен від віку двадцяти літ і вище, кожен, хто здатний до війська,
NUM|1|43|перелічені їхні від племени Нефталимового п'ятдесят і три тисячі й чотириста.
NUM|1|44|Оце ті перелічені, кого перелічив Мойсей й Аарон та Ізраїлеві начальники, дванадцятеро мужа, вони були по одному мужеві для дому батьків своїх.
NUM|1|45|І були всі перелічені з Ізраїлевих синів за домами батьків своїх від віку двадцяти літ і вище, кожен, хто здатний до війська, в Ізраїлі,
NUM|1|46|і були всі перелічені шістсот тисяч і три тисячі й п'ятсот і п'ятдесят.
NUM|1|47|А Левити не були перелічені серед них за племенем батьків своїх.
NUM|1|48|І Господь промовляв до Мойсея, говорячи:
NUM|1|49|Тільки Левієвого племени не переглянеш і не перелічиш їх серед Ізраїлевих синів.
NUM|1|50|А ти постав Левитів наглядачами над скинією свідоцтва, і над усіма речами її та над усім, що її. Вони будуть носити скинію та всі її речі, і вони будуть обслуговувати її, і отаборяться навколо скинії.
NUM|1|51|А коли скинія буде рушати, Левити розберуть її, а коли буде спинятися скинія, Левити поставлять її. А якщо наблизиться чужий, він нехай буде забитий.
NUM|1|52|І отаборяться Ізраїлеві сини кожен у таборі своїм, і кожен при своїм прапорі за своїми військовими відділами.
NUM|1|53|А Левити отаборяться навколо скинії свідоцтва, щоб не було гніву на громаду Ізраїлевих синів. І будуть Левити виконувати сторожу скинії свідоцтва.
NUM|1|54|І зробили Ізраїлеві сини, згідно зо всім, як наказав був Господь Мойсеєві, так зробили вони.
NUM|2|1|І Господь промовляв до Мойсея та до Аарона, говорячи:
NUM|2|2|Отаборяться Ізраїлеві сини кожен при прапорі своїм за ознаками домів своїх батьків, навпроти скинії заповіту навколо отаборяться.
NUM|2|3|Напереді на схід отаборяться: прапор Юдиного табору за своїми військовими відділами, а начальник Юдиних синів Нахшон, син Аммінадавів;
NUM|2|4|а його військо та його перелік сімдесят і чотири тисячі й шістсот.
NUM|2|5|А при ньому отабориться Іссахарове плем'я, а начальник Іссахарових синів Натанаїл, син Цуарів;
NUM|2|6|а його військо та його перелік п'ятдесят і чотири тисячі й чотириста.
NUM|2|7|Плем'я Завулонове, а начальник Завулонових синів Еліяв, син Хелонів;
NUM|2|8|а його військо та його перелік п'ятдесят і сім тисяч і чотириста.
NUM|2|9|Усіх перелічених Юдиного табору сто тисяч і вісімдесят тисяч і шість тисяч і чотириста за своїми військовими відділами. Вони рушать найперше.
NUM|2|10|Прапор Рувимового табору на південь, за військовими відділами своїми, а начальник Рувимових синів Еліцур, син Шедеурів;
NUM|2|11|а його військо та його перелік сорок і шість тисяч і п'ятсот.
NUM|2|12|А при ньому отабориться Симеонове плем'я, а начальник Симеонових синів Шелуміїл, син Цурішаддаїв;
NUM|2|13|а його військо та його перелік п'ятдесят і дев'ять тисяч і триста.
NUM|2|14|І Ґадове плем'я, а начальник Ґадових синів Ел'ясаф, син Реуїлів;
NUM|2|15|а його військо та його перелік сорок і п'ять тисяч і шістсот і п'ятдесят.
NUM|2|16|Усіх перелічених Рувимового табору сто тисяч і п'ятдесят і одна тисяча й чотириста й п'ятдесят за своїми військовими відділами. Вони рушать другі.
NUM|2|17|І як рушить скинія заповіту, то табір Левитів буде серед таборів. Як вони отаборяться, так вирушать, кожен на своїм місці за своїми прапорами.
NUM|2|18|Прапор Єфремового табору за військовими відділами своїми на захід, а начальник Єфремових синів Елішама, син Аммігудів;
NUM|2|19|а його військо та їхній перелік сорок тисяч і п'ятсот.
NUM|2|20|А при ньому плем'я Манасіїне, а начальник синів Манасіїних Гамаліїл, син Педацурів;
NUM|2|21|а його військо та їхній перелік тридцять і дві тисячі й двісті.
NUM|2|22|І Веніяминове плем'я, а начальник Веніяминових синів Авідан, син Ґід'оніїв;
NUM|2|23|а його військо та їхній перелік тридцять і п'ять тисяч і чотириста.
NUM|2|24|Усіх перелічених Єфремового табору сто тисяч і вісім тисяч і сто за своїми військовими відділами. Вони рушать треті.
NUM|2|25|Прапор Данового табору північ, за своїми військовими відділами, а начальник Данових синів Ахіезер, син Аммішаддаїв;
NUM|2|26|а його військо та їхній перелік шістдесят і дві тисячі й сімсот.
NUM|2|27|А при ньому отабориться Асирове плем'я, а начальник Асирових синів Паґ'іїл, син Охранів;
NUM|2|28|а його військо та їхній перелік сорок і одна тисяча й п'ятсот.
NUM|2|29|І плем'я Нефталимове, а начальник синів Нефталимових Ахіра, син Енанів;
NUM|2|30|а його військо та їхній перелік п'ятдесят і три тисячі й чотириста.
NUM|2|31|Усіх перелічених Данового табору сто тисяч і п'ятдесят і сім тисяч і шістсот. Вони рушать наостанку за прапорами своїми.
NUM|2|32|Оце перелічені Ізраїлевих синів за домами батьків своїх, усіх перелічених тих таборів за своїми військовими відділами шістсот тисяч і три тисячі й п'ятсот і п'ятдесят.
NUM|2|33|А Левити не перелічені серед Ізраїлевих синів, як Господь наказав був Мойсеєві.
NUM|2|34|І Ізраїлеві сини зробили все, що Господь наказав був Мойсеєві, так вони таборували за прапорами своїми, і так рушали кожен за своїми родами при домі своїх батьків.
NUM|3|1|А оце нащадки Ааронові та Мойсеєві в дні, коли Господь промовляв до Мойсея на Сінайській горі.
NUM|3|2|І оце імена Ааронових синів: перворідний Надав, і Авігу, Елеазар та Ітамар.
NUM|3|3|Оце імена Ааронових синів, помазаних священиків, що він посвятив їх бути священиками.
NUM|3|4|Та помер Надав та Авігу перед Господнім лицем, коли вони принесли були чужий огонь перед Господнім лицем у Сінайській пустині, а синів у них не було. І були священиками Елеазар та Ітамар за життя батька свого Аарона.
NUM|3|5|І Господь промовляв до Мойсея, говорячи:
NUM|3|6|Приведи Левієве плем'я, і постав його перед священиком Аароном, і вони будуть услуговувати йому.
NUM|3|7|І будуть вони виконувати сторожу його та всієї громади перед скинією заповіту, щоб виконувати службу скинійну.
NUM|3|8|І будуть вони стерегти всі речі скинії заповіту та сторожу Ізраїлевих синів, щоб виконувати службу скинійну.
NUM|3|9|І даси Левитів Ааронові та синам його, власне йому вони дані від Ізраїлевих синів.
NUM|3|10|А Аарона та синів його постав, щоб вони пильнували свого священства, а чужий, хто наблизиться, буде забитий.
NUM|3|11|І Господь промовляв до Мойсея, говорячи:
NUM|3|12|А Я оце взяв Левитів з-посеред Ізраїлевих синів замість кожного перворідного, що розкривають утробу, з Ізраїлевих синів. І будуть Левити Мої,
NUM|3|13|бо Мій кожен перворідний. Того дня, коли Я був ударив кожного перворідного в єгипетськім краї, Я посвятив Собі кожного перворідного в Ізраїлі від людини аж до скотини, Мої вони будуть. Я Господь!
NUM|3|14|І Господь промовляв до Мойсея в Сінайській пустині, говорячи:
NUM|3|15|Перелічи Левієвих синів за домами їхніх батьків, за родами їхніми, кожного чоловічої статі від місячного віку й вище перелічиш їх.
NUM|3|16|І Мойсей перелічив їх за Господнім словом, як йому наказано.
NUM|3|17|І були за йменнями своїми оці Левієві сини: Ґершон, і Кегат, і Мерарі.
NUM|3|18|А оце імена Ґершонових синів за їхніми родами: Лівні та Шім'ї.
NUM|3|19|А сини Кегатові за їхніми родами: Амрам і Їцгар, Хеврон і Уззіїл.
NUM|3|20|А сини Мерарі за їхніми родами: Махлі та Муші. Оце вони, роди Левієві, за домами своїх батьків.
NUM|3|21|Від Ґершона: рід Лівнієвих та рід Шім'їєвих. Оце вони, роди Ґершонових.
NUM|3|22|Перелічені їхні числом кожного чоловічої статі від місячного віку й вище, перелічені їхні сім тисяч і п'ятсот.
NUM|3|23|Роди Ґершонових будуть таборувати за наметом на захід.
NUM|3|24|А начальник батьківського дому Ґершонових Ел'ясаф, син Лаїлів.
NUM|3|25|А догляд Ґершонових синів у скинії заповіту: скинія внутрішня і намет зовнішній, і покриття його, і завіса входу скинії заповіту,
NUM|3|26|і запони подвір'я, і заслона входу подвір'я, що на скинії та на жертівнику навколо, і шнури її до всієї служби його.
NUM|3|27|А від Кегата: рід Амрамових, і рід Іцхарових, і рід Хевронових, і рід Оззіїлових, оце вони, роди Кегатових.
NUM|3|28|Числом кожного чоловічої статі від місячного віку й вище, вісім тисяч і шістсот, що пильнували сторожу святині.
NUM|3|29|Роди Кегатових синів отаборяться на подовжньому боці скинії на південь.
NUM|3|30|А начальник батькового дому родів Кегатових Еліцафан, син Уззіїлів.
NUM|3|31|А їхній догляд: ковчег, і стіл, і свічник, і жертівники, і святі речі, що служать ними, і завіса, і вся служба при тому.
NUM|3|32|А начальник Левієвих начальників Елеазар, син священика Аарона, що мав догляд над тими, хто пильнує сторожу святині.
NUM|3|33|Від Мерарі: рід Махлієвих, і рід Мушієвих, оце вони, роди Мерарієві.
NUM|3|34|А перелічені їхні числом кожного чоловічої статі від місячного віку й вище, шість тисяч і двісті.
NUM|3|35|А начальник батьківського дому Мерарієвих родів Цуріїл, син Авіхаїлів. Вони отаборяться на подовжнім боці скинії на північ.
NUM|3|36|А догляд сторожі Мерарієвих синів: дошки скинії, і засови її, і стовпи її, і підстави її, і всі речі її, і вся служба її,
NUM|3|37|і стовпи подвір'я навколо, і їхні підстави, і кілки їхні, і їхні шнури.
NUM|3|38|А ті, що таборують спереду перед скинією, перед скинією заповіту на схід, Мойсей й Аарон та сини його, вони виконують сторожу святині, сторожу за Ізраїлевих синів. А чужий, хто наблизиться, буде забитий.
NUM|3|39|Усі перелічені Левитів, що перелічив Мойсей та Аарон на Господній наказ за їхніми родами, кожен чоловічої статі від місячного віку й вище, двадцять і дві тисячі.
NUM|3|40|І сказав Господь до Мойсея: Перелічи всіх перворідних чоловічої статі Ізраїлевих синів від місячного віку й вище, і перелічи число імен їх.
NUM|3|41|І візьми для мене Левитів Я Господь! замість кожного перворідного Ізраїлевих синів, а худобу Левитів замість кожного перворідного серед худоби Ізраїлевих синів.
NUM|3|42|І перелічив Мойсей, як Господь наказав був йому, усіх перворідних серед Ізраїлевих синів.
NUM|3|43|І було всіх перворідних чоловічої статі числом імен від місячного віку й вище, за їхніми переліченими двадцять і дві тисячі двісті і сімдесят і три.
NUM|3|44|І Господь промовляв до Мойсея, говорячи:
NUM|3|45|Візьми Левитів замість кожного перворідного серед Ізраїлевих синів, а худобу Левитів замість їхньої худоби, і будуть Левити Мої. Я Господь!
NUM|3|46|А на окуп тих двохсот і семидесяти і трьох, що позостали понад Левитами з перворідного Ізраїлевих синів,
NUM|3|47|то візьми по п'яти шеклів на голову, на міру шеклем святині візьмеш, двадцять ґер шекель,
NUM|3|48|і даси ті гроші Ааронові та синам його, як окуп за позосталих серед них.
NUM|3|49|І взяв Мойсей гроші окупу від позосталих понад викуплених Левитами,
NUM|3|50|від перворідного Ізраїлевих синів узяв він ті гроші, тисячу і триста і шістдесят і п'ять на міру шеклем святині.
NUM|3|51|І дав Мойсей гроші окупу Ааронові та синами його за Господнім наказом, як Господь наказав був Мойсеєві.
NUM|4|1|І Господь промовляв до Мойсея й до Аарона, говорячи:
NUM|4|2|Перелічи Кегатових синів серед синів Левієвих за їхніми родами, за домами їхніх батьків
NUM|4|3|від віку тридцяти літ і вище й аж до віку п'ятидесяти літ, кожного, хто здатний до війська, щоб виконувати працю в наметі скинії заповіту.
NUM|4|4|Оце служба Кегатових синів у скинії заповіту: носити Святеє Святих.
NUM|4|5|Коли табір рушатиме, то ввійде Аарон та сини його, та й здіймуть завісу заслони, і покриють нею ковчега свідоцтва.
NUM|4|6|І дадуть на нього шкуряне тахашеве накриття, і розкладуть згори покривало, усе з блакиті, і накладуть держаки його.
NUM|4|7|А на столі показних хлібів розкладуть блакитну шату, і дадуть на нього миски, і ложки, і чаші, і кухлі на лиття, і хліб повсякчасний буде на ньому.
NUM|4|8|І розкладуть на них шату з червені, і покриють її шкуряним тахашевим покриттям, і накладуть держаки його.
NUM|4|9|І візьмуть блакитну шату, і покриють свічника освітлення, і лямпадки його, і щипці його, і його лопатки на вугіль, і всі посудини для оливи його, якими служать при ньому,
NUM|4|10|і покриють його і ввесь посуд його шкуряним тахашевим покриттям, і покладуть на держаки.
NUM|4|11|А на золотий жертівник розкладуть блакитну шату, і покриють його шкуряним тахашевим покриттям, і вкладуть його держаки.
NUM|4|12|І візьмуть увесь посуд служення, що ним служать у святині, і дадуть до блакитної шати, і покриють їх шкуряним тахашевим покриттям, і покладуть на держаки.
NUM|4|13|І заберуть попіл із жертівника, і розкладуть на ньому шату пурпурову,
NUM|4|14|і покладуть на нього ввесь посуд його, що ним служать на ньому: лопатки на вугіль, видельця, і шуфлі, і кропильниці, ввесь посуд жертівника; і розкладуть на ньому шкуряне тахашеве покриття, і вкладуть держаки його.
NUM|4|15|І скінчить Аарон та сини покривати святиню та ввесь святий посуд, коли табір рушає, а потім увійдуть Кегатові сини, щоб нести але не доторкнуться до святого, щоб не повмирати.
NUM|4|16|А догляд Елеазара, сина священика Аарона, олива освітлення, і кадило пахощів, і повсякчасна хлібна жертва, і олива помазання, догляд усієї скинії та всього, що в ній, у святині та в речах її.
NUM|4|17|І Господь промовляв до Мойсея й до Аарона, говорячи:
NUM|4|18|Не винищуйте племени Кегатових родів з-посеред Левитів.
NUM|4|19|І оце зробіть їм, і будуть жити й не повмирають, коли вони підходять до Святого Святих: увійдуть Аарон та сини його, і розмістять їх одного по одному на службі його та на ношенні його.
NUM|4|20|А самі вони не ввійдуть, щоб ані на хвилю не бачити святині, і щоб не повмирати.
NUM|4|21|І Господь промовляв до Мойсея, говорячи:
NUM|4|22|Перелічи також Ґершонових синів, вони за домами свої батьків, за родами своїми,
NUM|4|23|від віку тридцяти літ і вище аж до віку п'ятидесяти літ перелічиш їх усіх, хто здатний для праці, щоб служити в скинії заповіту.
NUM|4|24|Оце служба Ґершонових родів, на службу й на ношення:
NUM|4|25|вони будуть носити покривала скинії, і скинію заповіту, покриття її й покриття тахашеве, що на ній згори, і завісу входу скинії заповіту,
NUM|4|26|і запони подвір'я, і заслону входу брами подвір'я, що при скинії та при жертівнику навколо, і шнури їхні, і ввесь посуд служби їх, і все, що буде зроблене для них, і будуть служити вони.
NUM|4|27|На наказ Аарона та синів його буде вся служба Ґершонових синів щодо всього ношення їхнього та щодо всієї служби їхньої. І доручите їм пильнувати про все, що вони будуть носити.
NUM|4|28|Оце служба родів Ґершонових синів у скинії заповіту, а їхня сторожа у руці Ітамара, сина священика Ааронового.
NUM|4|29|Синів Мерарієвих за родами їхніми, за домами їхніх батьків перелічиш їх
NUM|4|30|від віку тридцяти літ і вище, й аж до віку п'ятидесяти літ, перелічиш їх кожного, хто здатний для праці, щоб служити в скинії заповіту.
NUM|4|31|А оце те, що вони повинні носити під час їхньої служби в скинії заповіту: дошки скинії, і засуви її, і стовпи її, і підстави її,
NUM|4|32|і стовпи подвір'я навколо, і їхні підстави, і їхні кілки, і їхні шнури, зо всіма їхніми речами, і зо всією службою їхньою, і пойменно перелічиш речі, що вони дбають про їхнє ношення.
NUM|4|33|Оце служба родин синів Мерарієвих щодо всієї їхньої служби в скинії заповіту під рукою Ітамара, сина священика Аарона.
NUM|4|34|І перелічив Мойсей та Аарон, та начальники громади Кегатових синів за їхніми родами й за домами їхніх батьків
NUM|4|35|від віку тридцяти літ і вище, і аж до віку п'ятидесяти літ, кожного, хто входить до відділу на службу в скинії заповіту.
NUM|4|36|І було їхніх перелічених за їхніми родами дві тисячі сімсот і п'ятдесят.
NUM|4|37|Оце перелічені Кегатових родів, кожен, хто працює в скинії заповіту, що перелічив Мойсей та Аарон за Господнім наказом через Мойсея.
NUM|4|38|А перелічені Ґершонових синів за своїми родами та за домами своїх батьків
NUM|4|39|від віку тридцяти літ і вище, і аж до віку п'ятидесяти літ, кожен, хто входить до відділу на службу в скинії заповіту,
NUM|4|40|і було їхніх перелічених за родами їхніми, за домами своїх батьків дві тисячі й шістсот і тридцять.
NUM|4|41|Оце перелічені родів Ґершонових синів, кожен, хто працює в скинії заповіту, що перелічив Мойсей та Аарон за Господнім наказом.
NUM|4|42|А перелічені родів синів Мерарієвих за їхніми родами, за домами своїх батьків
NUM|4|43|від віку тридцяти літ і вище, і аж до віку п'ятидесяти літ, кожен, хто входить до відділу на службу в скинії заповіту,
NUM|4|44|і було їхніх перелічених за родами їхніми три тисячі й двісті.
NUM|4|45|Оце перелічені родів синів Мерарієвих, що перелічив Мойсей та Аарон за Господнім наказом через Мойсея.
NUM|4|46|Усі перелічені Левити, кого перелічив Мойсей й Аарон та Ізраїлеві начальники, за родами своїми, за домами своїх батьків
NUM|4|47|від віку тридцяти літ і вище, і аж до віку п'ятидесяти літ, кожен, хто входить, щоб виконувати працю служби й працю ношення в скинії заповіту,
NUM|4|48|і було їхніх перелічених вісім тисяч і п'ятсот і вісімдесят.
NUM|4|49|За Господнім наказом перелічено їх через Мойсея кожного на службі його та на ношенні його. І були перелічені, як Господь наказав був Мойсеєві.
NUM|5|1|І Господь промовляв до Мойсея, говорячи:
NUM|5|2|Накажи Ізраїлевим синам, і нехай повисилають з табору кожного прокаженого, і кожного течивого, і кожного нечистого через доторкнення до мертвого тіла.
NUM|5|3|І чоловіка й жінку будете висилати, поза табір будете висилати їх, і вони не занечистять таборів своїх, що Я серед них пробуваю.
NUM|5|4|І зробили так Ізраїлеві сини, і повисилали їх поза табір, як Господь промовляв був Мойсеєві, так зробили Ізраїлеві сини.
NUM|5|5|І Господь промовляв до Мойсея, говорячи:
NUM|5|6|Промовляй до Ізраїлевих синів: Чоловік або жінка, коли зробить який людський гріх, чинячи тим спроневірення проти Господа, і завинить душа та,
NUM|5|7|то вони визнають свій гріх, що зробили, і кожен зверне найперше ціну провини своєї, і додасть до неї п'ятину її, та й дасть тому, кому завинив він.
NUM|5|8|А якщо в того чоловіка нема викупника, щоб йому звернути ту ціну провини, то провина та буде звернена Господеві, і буде це священикові, опріч барана очищення, що ним очистить його.
NUM|5|9|А кожне приношення зо всяких святощів Ізраїлевих синів, що принесуть священикові, буде йому.
NUM|5|10|І що хто посвятить, буде йому. Що хто дасть священикові, буде йому.
NUM|5|11|І Господь промовляв до Мойсея, говорячи:
NUM|5|12|Промовляй до Ізраїлевих синів і скажи їм: Кожен чоловік, коли жінка його зрадить і спроневірить його,
NUM|5|13|і буде хто злягатися з нею і буде затаєне від очей її чоловіка, і буде заховане, і вона занечиститься, а свідка проти неї нема, і вона не буде схоплена,
NUM|5|14|та на ньому перейде дух ревнощів, і він буде ревнивий за свою жінку, що вона занечищена; або перейде на ньому дух ревнощів, і він буде ревнивий за свою жінку, а вона не була занечищена,
NUM|5|15|то приведе той чоловік свою жінку до священика, і принесе за неї жертву її, десяту частину ефи ячної муки, оливи на неї виллє, і не дасть на неї ладану, бо це хлібна жертва ревнощів, жертва пригадувальна, що пригадує провину.
NUM|5|16|І священик приведе її, і поставить перед Господнім лицем.
NUM|5|17|І візьме священик святої води в глиняну посудину, і пороху, що буде на долівці скинії, візьме священик, та й дасть до води.
NUM|5|18|І поставить священик ту жінку перед лицем Господнім, і відкриє голову тієї жінки, і дасть на руки її хлібну жертву пригадувальну, це хлібна жертва ревнощів. А в руці священика буде гірка вода, що наводить прокляття.
NUM|5|19|І закляне її священик та й скаже до жінки: Якщо ніхто не лежав із тобою, і якщо ти не зрадила нечистим гріхом, живши з чоловіком своїм, очисться від гіркої води, що наводить прокляття!
NUM|5|20|А коли ж ти зрадила, живши з чоловіком своїм, і коли ти занечистилась, і хтось злігся з тобою, крім твого чоловіка,
NUM|5|21|і закляне священик ту жінку клятвою прокляття, і скаже священик тій жінці: Нехай дасть тебе Господь на прокляття та клятву серед народу твого тим, що Господь зробить стегно твоє опалим, а живіт твій напухлим,
NUM|5|22|і ввійде ця вода, що наводить прокляття, до нутра твого, щоб зробити живіт напухлим, і щоб зробити стегно опалим. А жінка та скаже: Амінь, амінь!
NUM|5|23|І напише священик ті прокляття на звої, й обмиє гіркою водою,
NUM|5|24|і напоїть ту жінку гіркою водою, що наводить прокляття; і ввійде в неї та вода, що наводить прокляття, і дає гіркий біль.
NUM|5|25|І візьме священик із руки тієї жінки ту хлібну жертву ревнощів, і буде колихати ту хлібну жертву перед Господнім лицем, та й принесе її до жертівника.
NUM|5|26|І візьме священик жменю з хлібної жертви, як пригадувальну частину, та й спалить на жертівнику. А потім напоїть ту жінку водою.
NUM|5|27|І напоїть водою, і станеться, якщо була вона занечищена й спроневірила своєму чоловікові, то ввійде в неї та вода, що наводить прокляття, і дасть гіркий біль, і опухне живіт її, і западе стегно її, і стане та жінка прокляттям серед народу свого.
NUM|5|28|А якщо та жінка не була занечищена, і чиста вона, то буде очищена, і буде здатна родити дітей.
NUM|5|29|Оце закон про ревнощі, коли зрадить жінка чоловікові своєму, і занечиститься,
NUM|5|30|або коли на чоловіка найде дух ревнощів, і він буде ревнивий за жінку свою, то поставить ту жінку перед Господнім лицем, а священик виконає над нею ввесь цей закон.
NUM|5|31|І буде очищений той чоловік від гріха, а жінка та понесе свій гріх.
NUM|6|1|І Господь промовляв до Мойсея, говорячи:
NUM|6|2|Промовляй до Ізраїлевих синів, і скажи їм: Чоловік або жінка, коли вирішиться скласти обітницю назіра, щоб посвятити себе Господеві,
NUM|6|3|то він стримається від вина та п'янкого напою, не буде пити оцту винного та оцту з п'янкого напою, і жодного виноградного соку не питиме, і не їстиме ані свіжого, ані сухого винограду.
NUM|6|4|Усі дні посвячення свого не буде він їсти нічого, що зроблене з винограду, від зернят аж до лушпиння.
NUM|6|5|Усі дні його посвячення на назіра бритва не торкнеться голови його; аж до виповнення днів, що посвятить Господеві, він буде святий, мусить запустити волосся голови своєї!
NUM|6|6|Усі дні посвячення його Господеві не підійде він до мертвого тіла,
NUM|6|7|навіть через батька свого та через матір свою, через брата свого та через сестру свою не занечиститься ними, коли б вони померли, бо на голові його посвячення Богу його.
NUM|6|8|Усі дні посвячення його святий він для Господа.
NUM|6|9|А коли хто помре при ньому несподівано нагло, і він занечистить цим голову свого посвячення, то оголить голову свою в день очищення свого, сьомого дня оголить її.
NUM|6|10|А восьмого дня він принесе дві горлиці або двоє голубенят до священика до входу скинії заповіту.
NUM|6|11|І священик принесе одне на жертву за гріх, а одне на цілопалення, і очистить його з того, що занечистився він мертвим тілом, і посвятить його голову того дня.
NUM|6|12|І почне він знову дні посвячення свого Господеві, і принесе однорічне ягня на жертву за провину. А перші дні його будуть надаремні, бо занечистилося його посвячення.
NUM|6|13|І оце закон про назіра: того дня, коли виповнюються дні його посвячення, священик приведе його до входу скинії заповіту.
NUM|6|14|І принесе він Господеві жертву свою, одне безвадне однорічне ягня на цілопалення, і одну безвадну однорічну вівцю на жертву за гріх, і одного безвадного барана на жертву мирну,
NUM|6|15|і кіш опрісноків із пшеничної муки, калачі, мішані в оливі, і прісні коржі, помазані оливою, і хлібну їхню жертву, і їхні литі жертви.
NUM|6|16|І принесе священик перед Господнє лице, і принесе його жертву за гріх та його цілопалення.
NUM|6|17|А барана принесе мирною жертвою для Господа на коші опрісноків, і священик принесе його хлібну жертву та його жертву литу.
NUM|6|18|І оголить той назір голову свого посвячення у входа скинії заповіту, і візьме волосся голови свого посвячення та й покладе на огонь, що під мирною жертвою.
NUM|6|19|І візьме священик варену лопатку з барана, і одного прісного калача з коша, і одного прісного коржика, та й дасть на долоні назіра, як він оголить голову свого посвячення.
NUM|6|20|І священик буде колихати їх, як колихання перед Господнім лицем. Це святощ для священика, понад грудину колихання й понад стегно приношення. А по цьому той назір може пити вино.
NUM|6|21|Оце закон про назіра, що обіцяє свою жертву Господеві за своє посвячення, крім того, на що спроможна рука його. За обітницею своєю, що обіцює, так він зробить за законом про посвячення його.
NUM|6|22|І Господь промовляв до Мойсея, говорячи:
NUM|6|23|Промовляй до Аарона та до синів його, говорячи: Так благословляйте Ізраїлевих синів, говорячи їм:
NUM|6|24|Нехай Господь поблагословить тебе, і нехай Він тебе стереже!
NUM|6|25|Нехай Господь засяє на тебе лицем Своїм, і нехай буде милостивий до тебе!
NUM|6|26|Нехай Господь зверне на тебе лице Своє, і хай дасть тобі мир!
NUM|6|27|Вони будуть кликати Ймення Моє на Ізраїлевих синів, а Я благословлятиму їх!
NUM|7|1|І сталося того дня, коли Мойсей закінчив ставити скинію, і помазав її, і посвятив її та всі речі її, і жертівника та всі речі його, і помазав їх та посвятив їх,
NUM|7|2|то поприносили Ізраїлеві начальники, голови домів своїх батьків, вони начальники племен, вони ті, що стояли над переліком,
NUM|7|3|і принесли свою жертву перед Господнє лице: шість критих возів, і дванадцять волів, віз на двох начальників, а віл на одного, і поставили їх перед скинію.
NUM|7|4|І промовив Господь до Мойсея, говорячи:
NUM|7|5|Візьми від них, і будуть вони, щоб виконувати службу скинії заповіту, і даси їх Левитам, кожному за службою його.
NUM|7|6|І взяв Мойсей вози та воли, та й дав їх Левитам:
NUM|7|7|два вози та чотири воли дав Ґершоновим синам, за їхньою службою,
NUM|7|8|а чотири вози та вісім волів дав синам Мерарієвим за їхньою службою під рукою Ітамара, сина священика Аарона.
NUM|7|9|А Кегатовим синам не дав, бо на них лежить служба святині, на плечах повинні носити.
NUM|7|10|І поприносили начальники жертву на понову жертівника в день його помазання, і поприносили начальники свою жертву перед жертівника.
NUM|7|11|А Господь промовляв до Мойсея: По одному начальнику на день нехай приносять своє приношення на понову жертівника.
NUM|7|12|І був той, хто першого дня приніс своє приношення, Нахшон, син Аммінадавів, Юдиного племени.
NUM|7|13|А жертва його: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|14|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|15|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|16|один козел на жертву за гріх,
NUM|7|17|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце приношення Нахшона, Аммінадавого сина.
NUM|7|18|Другого дня приніс Натанаїл, син Цуарів, начальник Іссахарів.
NUM|7|19|Приніс він своє приношення: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|20|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|21|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|22|один козел на жертву за гріх,
NUM|7|23|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Натанаїла, Цуарового сина.
NUM|7|24|Третього дня начальник Завулонових синів Еліяв, син Хелонів.
NUM|7|25|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|26|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|27|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|28|один козел на жертву за гріх,
NUM|7|29|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Еліява, Хелонового сина.
NUM|7|30|Четвертого дня начальник Рувимових синів Еліцур, син Шедеурів.
NUM|7|31|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|32|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|33|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|34|один козел на жертву за гріх,
NUM|7|35|на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Еліцура, Шедеурового сина.
NUM|7|36|П'ятого дня начальник Симеонових синів Шелуміїл, син Цурішаддаїв.
NUM|7|37|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|38|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|39|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|40|один козел на жертву за гріх,
NUM|7|41|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Шелуміїла, Цурішаддаєвого сина.
NUM|7|42|Шостого дня начальник Ґадових синів Ел'ясаф, син Деуїлів.
NUM|7|43|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|44|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|45|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|46|один козел на жертву за гріх,
NUM|7|47|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Ел'ясафа, Деуїлового сина.
NUM|7|48|Сьомого дня начальник Єфремових синів Елішама, син Аммігудів.
NUM|7|49|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|50|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|51|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|52|один козел на жертву за гріх,
NUM|7|53|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Елішами, Аммігудового сина.
NUM|7|54|Восьмого дня начальник синів Манасії, Гамаліїл, син Педоцурів.
NUM|7|55|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|56|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|57|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|58|один козел на жертву за гріх,
NUM|7|59|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Гамаліїла, Педоцурового сина.
NUM|7|60|Дев'ятого дня начальник Веніяминових синів Авідан, син Ґід'оніїв.
NUM|7|61|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|62|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|63|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|64|один козел на жертву за гріх,
NUM|7|65|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Авідана, Ґід'онієвого сина.
NUM|7|66|Десятого дня начальник Данових синів Ахіезер, син Аммішаддаїв.
NUM|7|67|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на хлібну жертву,
NUM|7|68|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|69|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|70|один козел на жертву за гріх,
NUM|7|71|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Ахіезера, Аммішаддаєвого сина.
NUM|7|72|Одинадцятого дня начальник Асирових синів Паґ'іїл, син Охранів.
NUM|7|73|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на мучну жертву,
NUM|7|74|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|75|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|76|один козел на жертву за гріх,
NUM|7|77|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Паґ'іїла, Охранового сина.
NUM|7|78|Дванадцятого дня начальник Нефталимових синів Ахіра, син Енанів.
NUM|7|79|Його жертва: одна срібна миска, сто й тридцять шеклів вага її, одна срібна кропильниця, сімдесят шеклів на міру шеклем святині, обидві повні пшеничної муки, мішаної в оливі, на мучну жертву,
NUM|7|80|одна кадильниця, десять шеклів золота, повна кадила,
NUM|7|81|одне теля, один баран, одне однорічне ягня на цілопалення,
NUM|7|82|один козел на жертву за гріх,
NUM|7|83|а на мирну жертву два воли, п'ять баранів, п'ять козлів, п'ять ягнят однорічних, оце жертва Ахіри, Енанового сина.
NUM|7|84|Оце обряд освячення жертівника в дні його помазання, від Ізраїлевих начальників: срібних мисок дванадцять, срібних кропильниць дванадцять, золотих кадильниць дванадцять,
NUM|7|85|сто й тридцять шеклів одна срібна миска, і сімдесят одна кропильниця. Усе срібло посудин дві тисячі й чотириста шеклів на міру шеклем святині.
NUM|7|86|Кадильниць золотих дванадцять, повні кадила, по десяти шеклів кадильниця на міру шеклем святині; усе золото кадильниць сто й двадцять шеклів.
NUM|7|87|Уся велика худоба на цілопалення: дванадцять телят, баранів дванадцять, ягнят однорічних дванадцять, та жертва хлібна їх, і козлів дванадцять на жертву за гріх.
NUM|7|88|А вся худоба мирної жертви: двадцять і чотири теляті, баранів шістдесят, козлів шістдесят, ягнят однорічних шістдесят. Оце обряд освячення жертівника по помазанні його.
NUM|7|89|А коли Мойсей входив до скинії заповіту, щоб говорити з Ним, то він чув голос, що говорив до нього з-понад віка, яке на ковчезі свідоцтва, з-поміж обох херувимів говорив Він до нього.
NUM|8|1|І Господь промовляв до Мойсея, говорячи:
NUM|8|2|Промовляй до Аарона та й скажи йому: Коли ти світитимеш лямпадки, то з переду свічника будуть світити сім лямпадок.
NUM|8|3|І Аарон зробив так, з переду свічника засвітив його лямпадки, як Господь наказав був Мойсеєві.
NUM|8|4|А оце робота свічника: він куття золоте аж до підстави його, аж до квіток його куття він. За взірцем, що Господь показав був Мойсеєві, так він зробив свічника.
NUM|8|5|І Господь промовляв до Мойсея, говорячи:
NUM|8|6|Візьми Левитів з-посеред Ізраїлевих синів, та й очисть їх.
NUM|8|7|І так зробиш їм, щоб очистити їх: покропи на них водою жертви за гріх, і нехай обголять бритвою все тіло своє, і нехай виперуть одежу свою, і стануть чисті.
NUM|8|8|І вони візьмуть теля, а його хлібна жертва пшенична мука, мішана в оливі, і друге теля візьмеш на жертву за гріх.
NUM|8|9|І приведеш Левитів до скинії заповіту, і збереш усю громаду Ізраїлевих синів.
NUM|8|10|І приведеш Левитів перед Господнє лице, а Ізраїлеві сини покладуть свої руки на Левитів.
NUM|8|11|І буде Аарон посвячувати Левитів, як посвячення перед Господнім лицем від Ізраїлевих синів, і будуть вони на роботу Господньої служби.
NUM|8|12|А Левити покладуть свої руки на голову телят, і зроби одного жертвою за гріх, а одного цілопаленням для Господа, щоб очистити Левитів.
NUM|8|13|І поставиш Левитів перед Аароном та перед синами його, і будеш посвячувати їх, як посвячення для Господа.
NUM|8|14|І відділиш Левитів з-поміж Ізраїлевих синів, і будуть Левити Мої.
NUM|8|15|А по цьому Левити ввійдуть, щоб служити в скинії заповіту, і ти їх очистиш, і віддаси їх, як жертву посвячення,
NUM|8|16|бо вони дані, Мені вони дані з-поміж Ізраїлевих синів; замість перворідного кожного з Ізраїлевих синів, що розкриває кожну утробу, узяв Я їх Собі,
NUM|8|17|бо Мій кожен перворідний серед Ізраїлевих синів, серед людини й серед худоби; того дня, коли Я побивав кожного перворідного в єгипетськім краї, Я посвятив їх Собі.
NUM|8|18|І взяв Я Левитів замість кожного перворідного серед Ізраїлевих синів.
NUM|8|19|І дав Я Левитів, як дар Ааронові та синам його з-поміж Ізраїлевих синів, щоб вони чинили службу Ізраїлевих синів в скинії заповіту, щоб очищали Ізраїлевих синів, щоб не було поразки серед Ізраїлевих синів, щоб Ізраїлеві сини підходили до святині.
NUM|8|20|І зробив Мойсей й Аарон та вся громада Ізраїлевих синів для Левитів усе, як Господь наказав був Мойсеєві про Левитів, так зробили їм Ізраїлеві сини.
NUM|8|21|І очистилися Левити, і випрали одяг свій, а Аарон посвятив їх перед Господнім лицем, і очистив їх Аарон, щоб стали чистими.
NUM|8|22|А по тому ввійшли Левити, щоб виконувати свою службу в скинії заповіту перед Аароном та перед синами його. Як Господь наказав був Мойсеєві про Левитів, так їм зробили вони.
NUM|8|23|І Господь промовляв до Мойсея, говорячи:
NUM|8|24|Оце щодо Левитів: від віку двадцяти й п'яти літ і вище ввійдуть вони до праці на службу скинії заповіту.
NUM|8|25|А від віку п'ятидесяти літ відійдуть від служби, і не будуть уже служити.
NUM|8|26|І будуть вони обслуговувати братів своїх у скинії заповіту, щоб виконувати сторожу, а служби не будуть робити. Так зробиш Левитам у їхній службі.
NUM|9|1|І Господь промовляв до Мойсея в Сінайській пустині другого року по виході з єгипетського краю, першого місця, говорячи:
NUM|9|2|І нехай справлять Ізраїлеві сини Пасху в означений час.
NUM|9|3|Чотирнадцятого дня цього місяця надвечір справите її означеного часу його, за всіма постановами її та за всіма уставами її спорядите її.
NUM|9|4|І Мойсей промовляв до Ізраїлевих синів, щоб справили Пасху.
NUM|9|5|І справили вони Пасху першого місяця, чотирнадцятого дня місяця надвечір у Сінайській пустині, усе, як Господь наказав був Мойсеєві, так зробили Ізраїлеві сини.
NUM|9|6|Та були люди, що були нечисті від дотику до тіла померлої людини, і не могли справити Пасху того дня. І прийшли вони того дня до Мойсея й до Аарона,
NUM|9|7|та й сказали ті люди до нього: Ми нечисті через дотик до тіла померлої людини. Чому ми будемо позбавлені ласки принести жертву Господню означеного часу серед Ізраїлевих синів?
NUM|9|8|І сказав до них Мойсей: Постійте, а я послухаю, що Господь накаже про вас.
NUM|9|9|І Господь промовляв до Мойсея, говорячи:
NUM|9|10|Промовляй до Ізраїлевих синів, говорячи: Кожен чоловік із вас, або з ваших нащадків, коли буде нечистий через дотик до мертвого тіла, або буде в далекій дорозі, то й він справить Пасху для Господа.
NUM|9|11|Місяця другого, чотирнадцятого дня надвечір спорядять вони її, з опрісноками та з гірким зіллям будуть їсти її.
NUM|9|12|Не позоставлять із неї до ранку, а костей не зламають у ній, за повною постановою Пасхи справлять її.
NUM|9|13|А чоловік, який чистий, а в дорозі не є, і стримається споряджати Пасху, то буде винищена душа та з народу її, бо Господньої жервти він не приніс означеного часу її. Гріх свій понесе той чоловік!
NUM|9|14|А коли перебуватиме з вами приходько, то справить він Пасху для Господа, за постановою про Пасху та за уставом про неї, так зробить. Постанова одна буде для вас, і для приходька, і для тубільця землі.
NUM|9|15|А того дня, коли поставлено скинію, хмара покрила скинію над ковчегом свідоцтва. А ввечорі було над скинією, як подоба огню, аж до ранку.
NUM|9|16|Так завжди бувало: удень покривала його та хмара, а вночі подоба огню.
NUM|9|17|І коли підіймалася хмара з-над скинії, то потому рушали Ізраїлеві сини, а на тому місці, на якому хмара ставала, там таборували Ізраїлеві сини.
NUM|9|18|На Господній наказ рушали Ізраїлеві сини, і на Господній наказ таборували. Усі ті дні, коли хмара перебувала над скинією, вони таборували.
NUM|9|19|А коли хмара багато днів позоставалася над скинією, то Ізраїлеві сини виконували Господню сторожу, і не рушали.
NUM|9|20|І бувало, що хмара була над скинією полічені дні, то вони на Господній наказ таборували, і на Господній наказ рушали.
NUM|9|21|І бувало, що хмара була від вечора аж до ранку, а підіймалася хмара вранці, то рушали вони. Або день і ніч була, і підіймалася хмара, то рушали вони.
NUM|9|22|Або два дні, або місяць, або рік хмара була над нею, над скинією, Ізраїлеві сини таборували, і не рушали, а коли вона підіймалась, рушали вони.
NUM|9|23|На Господній наказ таборували вони, і на Господній наказ рушали вони. Вони виконували Господню сторожу на Господній наказ через Мойсея.
NUM|10|1|Господь промовляв до Мойсея, говорячи:
NUM|10|2|Зроби собі дві срібні сурмі, куттям зробиш їх; і будуть вони тобі на скликання громади та на рушання таборів.
NUM|10|3|І засурмлять у них, і збереться до тебе громада при вході скинії зборів.
NUM|10|4|А якщо засурмлять в одну, то зберуться до тебе начальники, голови Ізраїлевих тисяч.
NUM|10|5|А засурмлять на сполох, то рушать табори, що таборують на сході.
NUM|10|6|А засурмите на сполох удруге, то рушать табори, що таборують на півдні, будуть сурмити на сполох, щоб рушали вони.
NUM|10|7|А на скликання зборів засурмите, але без сполоху.
NUM|10|8|А сурмити в сурми будуть Ааронові сини, священики. І ці сурмлення будуть для вас на вічну постанову для ваших поколінь.
NUM|10|9|А коли підете війною в вашому Краю на ворога, що гнобить вас, і засурмите на сполох, то ви будете згадані перед лицем Господа, Бога вашого, і будете спасені від ваших ворогів.
NUM|10|10|А в день вашої радости, і в ваші свята та першого дня ваших місяців засурмите в ті сурми на ваших цілопаленнях та на мирних жертвах ваших, і вони будуть вам на пригад перед лицем вашого Бога. Я Господь, Бог ваш!
NUM|10|11|І сталося, другого року, другого місяця, дванадцятого дня місяця піднялася хмара з-над скинії свідоцтва.
NUM|10|12|І рушили Ізраїлеві сини з Сінайської пустині на походи свої, і хмара спинилася в пустині Паран.
NUM|10|13|І рушили вони вперше за Господнім наказом через Мойсея.
NUM|10|14|І найперш рушив прапор табору синів Юдиних за своїми військовими відділами, а над військом його Нахшон, син Аммінадавів.
NUM|10|15|А над військом племени синів Іссахара Натанаїл, син Цуарів.
NUM|10|16|А над військом племени Завулонових синів Еліяв, син Хелонів.
NUM|10|17|І була розібрана скинія, і рушили Ґершонові сини та сини Мерарієві, носії скинії.
NUM|10|18|І рушив прапор табору Рувима за своїми військовими відділами, а над військом його Еліцур, син Шедеурів.
NUM|10|19|А над військом племени Симеонових синів Шелуміїл, син Цурішаддаїв.
NUM|10|20|А над військом племени Ґадових синів Ел'ясаф, син Деуїлів.
NUM|10|21|І рушили сини Кегатові, носії святині, та й поставили скинію до приходу їх, усіх інших.
NUM|10|22|І рушив прапор табору синів Єфремових за своїми військовими відділами, а над військом його Елішама, син Аммігудів.
NUM|10|23|А над військом племени синів Манасіїних Гамаліїл, син Педацурів.
NUM|10|24|А над військом племени Веніяминових синів Авідан, син Ґідеонів.
NUM|10|25|І рушив прапор табору синів Данових як задня сторожа для всіх таборів за своїми військовими відділами, а над військом його Ахіезер, син Аммішаддаїв.
NUM|10|26|А над військом племени Асирових синів Паґ'іїл, син Охрана.
NUM|10|27|А над військом племени синів Нефталимових Ахіра, син Енанів.
NUM|10|28|Оце походи Ізраїлевих синів за їхніми військовими відділами. І рушили вони.
NUM|10|29|І сказав Мойсей до Ховава, сина мідіянітянина Реуїла, Мойсеєвого тестя: Ми рушаємо до того місця, що про нього Господь був сказав: Його дам вам. Ходи ж із нами, і ми зробимо тобі добро, бо Господь промовляв був добро про Ізраїля.
NUM|10|30|Та той відказав йому: Не піду, але піду до краю свого та до місця своєї батьківщини.
NUM|10|31|А Мойсей відказав: Не покидай нас, бо через те, що ти знаєш наше таборування в пустині, то будеш нам очима.
NUM|10|32|І станеться, коли підеш із нами, то те добро, що Господь учинить нам, ми його вчинимо тобі.
NUM|10|33|І рушили вони від Господньої гори триденною дорогою. А ковчег заповіту Господнього рушав перед ними триденною дорогою, щоб вивідати для них місце спинитися.
NUM|10|34|А хмара Господня була над ними вдень, коли вони рушали з табору.
NUM|10|35|І бувало, коли ковчег вирушав, то Мойсей промовляв: Устань же, о Господи, і хай розпорошаться Твої вороги, і хай повтікають Твої ненависники з-перед Твойого лиця.
NUM|10|36|А коли він ставав, то говорив: Вернися, о Господи, до десятьтисячок тисяч Ізраїля!
NUM|11|1|І став народ голосно нарікати до Господніх ушей. І почув Господь, і запалав Його гнів, і загорівся між ними Господній огонь, та й пожер їх у кінці табору.
NUM|11|2|І народ став кричати до Мойсея. А Мойсей помолився до Господа, і погас той огонь.
NUM|11|3|І він назвав ім'я того місця: Тав'ера, бо між ними горів був Господній огонь.
NUM|11|4|А збиранина, що була серед нього, стала вередувати, і також Ізраїлеві сини стали плакати з ними та говорити: Хто нагодує нас м'ясом?
NUM|11|5|Ми згадуємо рибу, що їли в Єгипті даремно, огірки й дині, і пір, і цибулю, і часник.
NUM|11|6|А тепер душа наша в'яне, немає нічого, тільки манна нам перед очима.
NUM|11|7|А манна як коріяндрове насіння вона, а вигляд її, як вигляд кришталу.
NUM|11|8|Люди розходилися, і збирали її та мололи жорнами або товкли в ступі, і варили в горшку та й робили з неї калачі. А смак її був, як смак олійного коржа.
NUM|11|9|А коли роса спадала на табір, спадала й та манна на нього.
NUM|11|10|І почув Мойсей, що народ плаче в родинах своїх, кожен при вході намету свого. І сильно запалав гнів Господній, і в очах Мойсеєвих то було зле.
NUM|11|11|І сказав Мойсей до Господа: Нащо вчинив Ти зло своєму рабові, і чому я не знайшов милости в очах Твоїх, що Ти поклав тягара всього народу на мене?
NUM|11|12|Чи я був вагітний усім тим народом, чи я його породив, що Ти кажеш мені: Неси його на лоні своїм, як мамка носить ссунця, до землі, яку Ти присягнув батькам його?
NUM|11|13|Звідки мені взяти м'яса, щоб дати всьому цьому народові? Бо вони плачуть передо мною, говорячи: Дай же нам м'яса, і ми будемо їсти!
NUM|11|14|Не подолаю я сам носити всього цього народа, бо він тяжчий за мене!
NUM|11|15|А якщо Ти таке мені робиш, то краще забий мене, якщо я знайшов милість в очах Твоїх, щоб я не побачив нещастя свого!
NUM|11|16|І сказав Господь до Мойсея: Збери ж мені сімдесятеро люда зо старших Ізраїлевих, яких знаєш, що вони старші народу та його наглядачі, і візьми їх до скинії заповіту, і стануть вони там із тобою.
NUM|11|17|І Я зійду, і буду розмовляти там із тобою, і візьму від Духа, що на тобі, і покладу на них, і вони носитимуть із тобою тягара того народу, і не будеш носити ти сам.
NUM|11|18|А до народу скажи: Освятіться назавтра, і будете їсти м'ясо, бо ви плакали до Господніх ушей, говорячи: Хто дасть нам їсти м'яса, бо добре було нам в Єгипті? І дасть Господь вам м'яса, і ви будете їсти.
NUM|11|19|Не один день будете ви їсти, і не два дні, і не п'ять день, і не десять день, і не двадцять день,
NUM|11|20|але цілий місяць, аж поки не вийде воно з ваших ніздрів, і стане вам на огиду, бо ви знехтували собі Господа, що серед вас, і плакали перед лицем Його, говорячи: Чого це ми вийшли з Єгипту?
NUM|11|21|І сказав Мойсей: Шістсот тисяч піхоти той народ, що я серед нього, а Ти сказав: Я дам їм м'яса, і вони будуть їсти місяць часу.
NUM|11|22|Чи худоба дрібна та худоба велика заріжеться для них, і вистачить їм? Чи також збереться для них уся морська риба, і вистачить їм?
NUM|11|23|А Господь сказав до Мойсея: Чи Господня рука буває коротка? Тепер ти побачиш, чи сповниться тобі Моє слово, чи ні.
NUM|11|24|І вийшов Мойсей, і промовляв до того народу Господні слова. І зібрав він сімдесятеро чоловіка зо старших народу, і поставив їх навколо скинії.
NUM|11|25|І зійшов Господь у хмарі, та й промовляв до нього, і взяв від Духа, що на ньому, і дав на сімдесят чоловіка старших. І сталося, як спочив на них Дух той, то вони стали пророкувати, та потім перестали.
NUM|11|26|І зосталося двоє людей в таборі, ім'я одному Елдад, а ймення другому Медад. І спочив на них Дух; а вони були серед записаних, та не вийшли до скинії, і пророкували в таборі.
NUM|11|27|І побіг юнак, і промовив до Мойсея й сказав: Елдад і Медад пророкують у таборі!
NUM|11|28|І відповів Ісус, син Навинів, Мойсеїв слуга від своєї молодости, та й сказав: Пане мій Мойсею, заборони їм!
NUM|11|29|І сказав йому Мойсей: Чи ти заздрісний за мене? О, якби то ввесь Господній народ став пророками, коли б дав Господь Духа Свого і на них!
NUM|11|30|І вернувся Мойсей до табору, він та старші Ізраїлеві.
NUM|11|31|І знявся вітер від Господа, і навіяв перепелиці від моря, і опустив їх над табором, як денна дорога туди й як денна дорога сюди навколо табору, і коло двох ліктів на поверхні землі.
NUM|11|32|І встав народ, і цілий той день і цілу ту ніч, і цілий день назавтра збирали перепелицю. Хто збирав мало, той зібрав десять хомерів, і порозкладали їх собі скрізь навколо табору.
NUM|11|33|Те м'ясо було ще між їхніми зубами, поки було пожуване, а гнів Господній запалився на народ! І вдарив Господь дуже великою поразкою в народ...
NUM|11|34|І названо ймення того місця: Ківрот-Гаттаава, бо там поховали народ пожадливий.
NUM|11|35|З Ківрот-Гаттаави рушили люди до Гацероту, і були в Гацероті.
NUM|12|1|І нарікали Маріям та Аарон на Мойсея за жінку кушитянку, що взяв, бо він узяв був жінку кушитянку.
NUM|12|2|І казали вони: Чи тільки з Мойсеєм Господь говорив? Чи ж не говорив Він також із нами? І почув це Господь.
NUM|12|3|А той муж, Мойсей, був найлагідніший за всяку людину, що на поверхні землі.
NUM|12|4|І нагло сказав Господь до Мойсея й до Аарона та до Маріям: Вийдіть ви троє до скинії заповіту. І вони троє вийшли.
NUM|12|5|І зійшов Господь у стовпі хмари, і став при вході скинії, та й покликав Аарона й Маріям. І вийшли обоє вони.
NUM|12|6|І сказав Він: Послухайте ж ви Моїх слів: Якщо буде між вами пророк, то Я, Господь, дамся пізнати в видінні йому, у сні говорити з ним буду.
NUM|12|7|Не так раб мій Мойсей: у всім домі Моїм він довірений!
NUM|12|8|Говорю Я з ним уста до уст, а не видінням і не загадками, і Образ Господа він оглядає. І чому не боялися ви нарікать на Мойсея, Мойого раба?
NUM|12|9|І запалав гнів Господній на них, і Він пішов,
NUM|12|10|а хмара відступила з-над скинії. А ось Маріям прокажена, збілівши, як сніг! І обернувся Аарон до Маріям, аж ось вона прокажена!
NUM|12|11|І сказав Аарон до Мойсея: Будь ласкав, мій пане, не поклади ж на нас гріха, що були ми нерозумні та що прогрішились!
NUM|12|12|Нехай же не буде вона, як та мертва дитина, що, як виходить з утроби матері своєї, то зітліла половина тіла її.
NUM|12|13|І Мойсей кликав до Господа, говорячи: Боже, вилікуй же її!
NUM|12|14|І сказав Господь до Мойсея: А коли б її батько справді плюнув на обличчя її, чи не буде вона сім день засоромлена? Вона буде замкнена сім день поза табором, а потім повернеться.
NUM|12|15|І була замкнена Маріям поза табором сім день, а народ не рушив аж до повернення Маріям.
NUM|12|16|А потім рушив народ із Гацероту, і таборував у пустині Паран.
NUM|13|1|І промовляв Господь до Мойсея, говорячи:
NUM|13|2|Пошли людей, і вони розвідають ханаанський Край, що Я даю Ізраїлевим синам; пошлете по одному чоловікові від племени своїх батьків, кожного начальника в них.
NUM|13|3|І послав їх Мойсей з пустині Паран за Господнім наказом. Усі вони мужі достойні, вони голови Ізраїлевих синів.
NUM|13|4|А оце ймення їх: для Рувимового племени Шаммуа, син Заккурів;
NUM|13|5|для Симеонового племени Шафат, син Хоріїв;
NUM|13|6|для Юдиного племени Калев, син Єфуннеїв;
NUM|13|7|для Іссахарового племени Їґ'ал, син Йосипів;
NUM|13|8|для Єфремового племени Осія, син Навинів;
NUM|13|9|для Веніяминового племени Палті, син Рафуїв;
NUM|13|10|для Завулонового племени Ґаддіїл, син Содіїв;
NUM|13|11|для Йосипового племени, для племени Манасіїного Ґадді, син Сусіїв;
NUM|13|12|для Данового племени Амміїл, син Ґемалліїв;
NUM|13|13|для Асирового племени Сетур, син Михаїлів;
NUM|13|14|для Нефталимового племени Нахбі, син Вофсіїв;
NUM|13|15|для Ґадового племени Ґеуїл, син Махіїв.
NUM|13|16|Оце ймення тих людей, що Мойсей послав був розвідати той Край. І назвав Мойсей Осію, Навинового сина: Ісус.
NUM|13|17|І послав їх Мойсей розвідати Край ханаанський, та й промовив до них: Підіть тут на південь, і ввійдете на гору,
NUM|13|18|та й побачите той Край який він, і народ, що сидить у ньому, чи сильний він, чи слабий, чи малий він, чи численний?
NUM|13|19|І який той Край, що він сидить у ньому, чи він добрий чи злий? І які ті міста, що він сидить у них, чи в таборах, чи в твердинях?
NUM|13|20|І яка та земля, чи масна вона, чи пісна? Чи є на ній дерево, чи ні? І будьте відважні, і візьміть з плоду землі; а дні ці дні виноградного первоплоду.
NUM|13|21|І знялися вони, і розвідали той Край від пустині Цін аж до Рехова, у напрямі до Хамоту.
NUM|13|22|І пішли вони на південь, і прибули аж до Хеврону, а там були Ахіман, Шешай та Талмай, нащадки велетня. А Хеврон був збудований за сім літ перед Цоаном єгипетським.
NUM|13|23|І прибули вони аж до долини Ешколу, і витяли там галузку з одним гроном винограду, і вдвох понесли його на жердині; також узяли із гранатів та з фіґ.
NUM|13|24|Те місце назвали: Нахал-Ешкол, через те гроно, що Ізраїлеві сини витяли були там.
NUM|13|25|І вернулися вони з розвідки того Краю по сорока днях.
NUM|13|26|І пішли, і прийшли вони до Мойсея й до Аарона та до всієї громади Ізраїлевих синів, до пустині Паран, до Кадешу, і здали справу їм та всій тій громаді, і показали плід того Краю.
NUM|13|27|І вони розповіли йому та й сказали: Прибули ми до Краю, куди ти послав був нас, а він тече молоком та медом, а оце плід його!
NUM|13|28|Та народ той, що сидить у тім Краї, міцний, а міста укріплені, дуже великі. А також бачили ми там нащадків велетня...
NUM|13|29|Амалик сидить у краї південнім, а хіттеянин, і євусеянин, і амореянин сидять на горі, а ханаанеянин сидить над морем та при Йордані.
NUM|13|30|А Калев утихомирював народ перед Мойсеєм та й сказав: Конче ввійдемо ми й заволодіємо ним, бо ми справді переможем його!
NUM|13|31|Та люди, що ходили з ним, сказали: Ми не зможемо ввійти до того народу, бо він сильніший за нас...
NUM|13|32|І пустили вони між Ізраїлевими синами злу вістку про той Край, що розвідали його, говорячи: Той Край, що ми перейшли по ньому, щоб розвідати його, це край, який поїдає своїх мешканців. А ввесь той народ, що ми бачили в ньому, люди високі на зріст.
NUM|13|33|І там ми бачили велетнів, синів Енака, з роду велетнів, і були ми в своїх очах немов та сарана, і такими були ми і в їхніх очах.
NUM|14|1|І зняла зойк уся та громада, та й заголосила. І плакав народ той тієї ночі.
NUM|14|2|І нарікали на Мойсея та на Аарона всі Ізраїлеві сини. І сказала до них вся громада: О, якби ми померли були в єгипетськім краї, або щоб ми померли були в цій пустині!
NUM|14|3|І нащо Господь провадить нас до того Краю, щоб нам попадати від меча? Жінки наші та діти наші стануть здобиччю... Чи не краще нам вернутися до Єгипту?
NUM|14|4|І сказали вони один до одного: Оберімо собі голову, та й вертаймось до Єгипту!
NUM|14|5|І впали Мойсей та Аарон на обличчя свої перед усім збором громади Ізраїлевих синів.
NUM|14|6|А Ісус, син Навинів, та Калев, син Єфуннеїв, із тих, що розвідували той Край, пороздирали одежу свою,
NUM|14|7|та й сказали до всієї громади Ізраїлевих синів, говорячи: Той Край, що перейшли ми по ньому, щоб розвідати його, Край той дуже-дуже хороший!
NUM|14|8|Якщо Господь уподобає Собі нас, то впровадить нас до того Краю, і дасть його нам, Край, який тече молоком та медом.
NUM|14|9|Тільки не бунтуйтесь проти Господа, і не бійтеся народу того Краю, бо вони хліб для нас! Їхня тінь відійшла від них, а з нами Господь, не бійтеся їх!
NUM|14|10|І сказала була вся громада, щоб камінням закидати їх, та слава Господня появилася в скинії заповіту всім Ізраїлевим синам...
NUM|14|11|І промовив Господь до Мойсея: Аж доки буде цей народ зневажати Мене, і аж доки не будуть вони вірувати в Мене, у всі ті ознаки, що Я учинив був серед нього?
NUM|14|12|Ударю його поразою, і позбавлю його насліддя, а тебе зроблю народом більшим і сильнішим від нього.
NUM|14|13|І сказав Мойсей до Господа: І почує Єгипет, що Ти з-посеред нього вивів Своєю силою народ цей,
NUM|14|14|та й скаже до мешканців цього Краю, які чули, що Ти Господь серед цього народу, що око-в-око являєшся Ти, Господи, а хмара Твоя стоїть над ними, і що Ти ходиш перед ними в стовпі хмари вдень, а в стовпі огню вночі,
NUM|14|15|якщо заб'єш Ти цей народ, як одну людину, то скажуть ті люди, що чули слух про Тебе, говорячи:
NUM|14|16|Через неспроможність Господа впровадити той народ до Краю, якого Він заприсяг був їм, вигубив їх у пустині...
NUM|14|17|А тепер нехай же звеличиться сила Господня, як Ти наказав був, говорячи:
NUM|14|18|Господь довготерпеливий, і багатомилостивий, Він прощає провину та переступ, і не очистить винного, а карає провину батьків на третіх і на четвертих поколіннях.
NUM|14|19|Прости ж провину цього народу через велику милість Свою, як прощав Ти цьому народові від Єгипту й аж сюди!
NUM|14|20|А Господь сказав: Я простив за словом твоїм.
NUM|14|21|Але, як Я живий, слава Господня наповнить увесь оцей Край.
NUM|14|22|Тому всі ті люди, що бачили славу Мою та ознаки Мої, що чинив Я в Єгипті та в пустині, але випробовували Мене оце десять раз та не слухалися голосу Мого,
NUM|14|23|поправді кажу, не побачать вони того Краю, що Я заприсяг був їхнім батькам. І всі, хто зневажає Мене, не побачать його!
NUM|14|24|Але раб Мій Калев за те, що з ним був дух інший, і він виконував накази Мої, то Я введу його до того Краю, куди він увійшов був, і потомство його оволодіє ним.
NUM|14|25|А амаликитянин та ханаанеянин сидить у долині. Узавтра оберніться, та й рушайте на пустиню дорогою Червоного моря!
NUM|14|26|І Господь промовляв до Мойсея й до Аарона, говорячи:
NUM|14|27|Аж доки цій злій громаді нарікати на Мене? Нарікання Ізраїлевих синів, що вони нарікають на Мене, Я чув.
NUM|14|28|Скажи їм: Живий Я! Мова Господня: Поправді кажу, як ви говорили до ушей Моїх, так Я зроблю вам.
NUM|14|29|У цій пустині попадають ваші трупи, та всі перелічені ваші всім вашим числом від віку двадцяти літ і вище, що нарікали на Мене.
NUM|14|30|Поправді кажу, ви не ввійдете до того Краю, що Я підносив був на присягу руку Свою, що будете перебувати в нім, окрім Калева, сина Єфуннеєвого, та Ісуса, сина Навинового.
NUM|14|31|А діти ваші, що про них казали ви: станете здобиччю ворогові, то впроваджу Я їх, і пізнають вони цей Край, яким ви обридили.
NUM|14|32|І ваші власні трупи попадають у цій пустині!
NUM|14|33|А ваші сини будуть блукати на пустині сорок літ, і відповідатимуть за зраду вашу, аж поки вигинуть ваші трупи на пустині.
NUM|14|34|Числом тих днів, що розвідували ви той Край, сорок день, будете ви нести ваші гріхи по року за день сорок літ, і пізнаєте, що значить бути покинутими Мною!
NUM|14|35|Я, Господь, говорив: Поправді кажу, оце зроблю всій цій злій громаді, що змовляється проти Мене: у цій пустині вигинуть, і тут повмирають.
NUM|14|36|А ті люди, яких Мойсей послав був розвідати той Край, коли вернулися, то зробили, що вся громада нарікала на нього, і пустили злу вістку на той Край,
NUM|14|37|то ті люди, що пустили були злу вістку на той Край, повмирали від порази перед Господнім лицем.
NUM|14|38|А Ісус, син Навинів, та Калев, син Єфуннеїв, жили з тих людей, що ходили розвідати той Край.
NUM|14|39|І говорив Мойсей ці слова до всіх Ізраїлевих синів, і народ був у тяжкій жалобі!
NUM|14|40|І повставали вони рано вранці, та й повиходили на верхів'я гори, говорячи: Ось ми, і ми підемо до місця, що Господь був сказав, бо ми прогрішили.
NUM|14|41|А Мойсей сказав: Чому ж ви переступаєте наказ Господній? Таж це не вдасться!
NUM|14|42|Не виходьте, бо Господь не серед вас, а то будете побиті своїми ворогами.
NUM|14|43|Бо там перед вами амаликитянин і ханаанеянин, і ви попадаєте від меча, бо ви відвернулися від Господа, і не буде Господь із вами.
NUM|14|44|Але вони осмілилися вийти на верхів'я гори, а ковчег свідоцтва Господнього та Мойсей не рушилися з-посеред табору.
NUM|14|45|І зійшов амаликитянин та ханаанеянин, що сидить на тій горі, та й побили їх, і били їх аж до Хорми.
NUM|15|1|І Господь промовляв до Мойсея, говорячи:
NUM|15|2|Промовляй до Ізраїлевих синів і скажеш їм: Коли ви ввійдете до Краю ваших осель, що Я даю вам,
NUM|15|3|і принесете огняну жертву для Господа, цілопалення, або криваву жертву на сповнення обітниці, або в дарі, або в означених часах при спорядженні любих пахощів для Господа з худоби великої або з худоби дрібної,
NUM|15|4|то той, хто приносить, принесе свою жертву для Господа, хлібну жертву, десяту частину ефи пшеничної муки, мішаної в чверті гіна оливи,
NUM|15|5|і вина для литої жертви принесеш чверть гіна на цілопалення або для жертви для кожного ягняти.
NUM|15|6|Або для барана принесеш хлібну жертву, дві десятих частини ефи пшеничної муки, мішаної в оливі третьої частини гіна.
NUM|15|7|І вина для литої жертви третю частину гіна, принесеш пахощі любі для Господа.
NUM|15|8|А коли принесеш молодого бичка як цілопалення, або як жертву на сповнення обітниці, або як мирну жертву для Господа,
NUM|15|9|то принесеш молодого бичка і хлібну жертву, три десяті частини ефи пшеничної муки, мішаної в оливі половини гіна.
NUM|15|10|І принесеш на литу жертву пів гіна вина, жертва огняна, пахощі любі для Господа.
NUM|15|11|Так буде робитися для одного вола, або для одного барана, або для ягняти з-поміж овець, або з-поміж кіз.
NUM|15|12|За числом жертов, що принесете, так зробите для кожної, за числом їх.
NUM|15|13|Кожен тубілець так принесе це, щоб принести огняну жертву, пахощі любі для Господа.
NUM|15|14|А коли з вами буде тимчасово мешкати приходько, або той, що серед вас, постанова для ваших поколінь, то він принесе огняну жертву, пахощі любі для Господа, як принесете ви, так принесе й він.
NUM|15|15|Збори, постанова одна для вас та для приходька, що мешкає тимчасово, постанова вічна для ваших поколінь: як ви, так і приходько буде перед Господнім лицем!
NUM|15|16|Один закон і одна постанова буде вам і приходькові, що мешкає тимчасово з вами.
NUM|15|17|І Господь промовляв до Мойсея, говорячи:
NUM|15|18|Промовляй до синів Ізраїлевих, та й скажи їм: Як ви ввійдете до Краю, що Я впроваджую вас туди,
NUM|15|19|то станеться, коли ви їстимете хліб того Краю, ви принесете приношення для Господа.
NUM|15|20|Як початок діж ваших, калача принесете на приношення, як приношення току, принесете його.
NUM|15|21|Від початку діж ваших дасте Господеві приношення, постанова для ваших поколінь!
NUM|15|22|А коли ви помилитеся, і не виконаєте всіх тих заповідей, що Господь говорив до Мойсея,
NUM|15|23|усього, що наказав вам Господь через Мойсея, від дня, коли Господь наказав був і далі для ваших поколінь,
NUM|15|24|то станеться, коли зроблено помилку через недогляд громади, нехай вся громада принесе одного бичка, молоде з великої худоби, на цілопалення, на пахощі любі для Господа, а хлібна його жертва та лита жертва його за постановою, і козла на жертву за гріх.
NUM|15|25|І очистить священик всю громаду синів Ізраїлевих, і буде прощено їм, бо то помилка, а вони принесли жертву свою, жертву огняну для Господа та жертву свою за гріх перед лице Господнє за свою помилку.
NUM|15|26|І буде прощено всій громаді Ізраїлевих синів та приходькові, що мешкає тимчасово серед них, бо то помилковий гріх усього народу.
NUM|15|27|А якщо згрішить помилково одна душа, то вона принесе однорічну козу на жертву за гріх.
NUM|15|28|І очистить священик ту душу, що помилилась, що згрішила помилково перед Господнім лицем, на очищення її, і буде прощено їй.
NUM|15|29|Тубільцеві серед Ізраїлевих синів та приходькові, що мешкає тимчасово серед них, закон один буде вам для того, хто зробить гріх помилково.
NUM|15|30|А та душа, що зробить зухвалою рукою, чи з тубільця, чи з приходька, він Господа зневажає, і буде винищена душа та з-посеред народу її.
NUM|15|31|Бо він знехтував слово Господа, і зламав Його заповідь, конче буде винищена душа та, гріх її на ній.
NUM|15|32|І були Ізраїлеві сини в пустині, та й знайшли чоловіка, що збирає дрова суботнього дня.
NUM|15|33|І привели його ті, хто знайшов його, як збирав дрова, до Мойсея й до Аарона та до всієї громади.
NUM|15|34|І взяли його під сторожу, бо не було вирішене, що зробити йому.
NUM|15|35|І сказав Господь до Мойсея: Конче буде забитий цей чоловік, закидати його камінням усій громаді поза табором!
NUM|15|36|І випровадила його вся громада поза табір, та й закидала його камінням, і він помер, як Господь наказав був Мойсеєві.
NUM|15|37|І сказав Господь до Мойсея, говорячи:
NUM|15|38|Промовляй до Ізраїлевих синів, та й скажи їм: Нехай вони зроблять собі кутаси на краях своїх одеж, вони й їхні покоління, і дадуть на кутаса поли блакитну нитку.
NUM|15|39|І буде вона вам за кутаса, і будете бачити його, і пам'ятатимете всі Господні заповіді, і виконаєте їх, і не будете оглядатися за серцем своїм та за очима своїми, за якими йдучи, ви зраджуєте,
NUM|15|40|щоб згадували ви та виконували всі Мої заповіді, і будьте святі для вашого Бога!
NUM|15|41|Я Господь, Бог ваш, що вивів вас з єгипетського краю, щоб бути вашим Богом. Я Господь, Бог ваш!
NUM|16|1|І взяли Корей, син Їцгара, сина Кегата, сина Левієвого, і Датан, і Авірон, сини Еліявові, та Он, син Пелета, сини Рувимові,
NUM|16|2|та й повстали проти Мойсея, а з ними двісті й п'ятдесят мужа Ізраїлевих синів, начальники громади, закликувані на збори, люди вельможні.
NUM|16|3|І зібралися вони на Мойсея та на Аарона, та й сказали до них: Досить вам, бо вся громада усі вони святі, а серед них Господь! І чому ви несетеся понад зборами Господніми?
NUM|16|4|І почув це Мойсей, та й упав на обличчя своє.
NUM|16|5|І промовив він до Корея та до всієї громади його, говорячи: Уранці Господь дасть знати, хто Його та хто святий, щоб наблизити його до Себе; а кого вибере, того Він і наблизить до Себе.
NUM|16|6|Зробіть ви оце: візьміть собі кадильниці, Корею та вся громадо твоя,
NUM|16|7|і дайте в них огню та покладіть на них кадила перед Господнє лице взавтра. І станеться, той чоловік, що Господь його вибере, він святий. Досить вам, Левієві сини!
NUM|16|8|І сказав Мойсей до Корея: Слухайте ж, Левієві сини,
NUM|16|9|чи вам мало, що Бог Ізраїлів відділив вас від Ізраїлевої громади, щоб наблизити вас до Себе, і щоб ви виконували службу Господньої скинії, і стояли перед громадою, щоб служити їй?
NUM|16|10|І Він наблизив тебе та всіх братів твоїх, Левієвих синів, із тобою; а ти будеш домагатися ще й священства?.
NUM|16|11|Тому ти та вся громада твоя змовилися проти Господа. А Аарон, що він, що ви ремствуєте проти нього?
NUM|16|12|І послав Мойсей та Аарон закликати Датана й Авірона, синів Еліявових, та сказали вони: Не вийдемо!
NUM|16|13|Чи мало того, що ти вивів нас із краю, який тече молоком та медом, щоб повбивати нас у пустині? Хочеш ще панувати над нами, щоб бути також вельможею?
NUM|16|14|Ти не впровадив нас ані до Краю, що тече молоком та медом, ані не дав нам на власність поля та виноградники. Чи ти вибереш очі цим людям? Не вийдемо!
NUM|16|15|А Мойсей сильно запалився, та й сказав до Господа: Не обернися до їхнього приношення! Я не взяв від них жодного осла, і зла не вчинив жодному з них!
NUM|16|16|І сказав Мойсей до Корея: Ти та вся громада твоя будьте перед Господнім лицем, ти й вони та Аарон узавтра.
NUM|16|17|І візьміть кожен свою кадильницю, і покладіть на неї кадила та й принесете перед Господнє лице кожен кадильницю свою, двісті й п'ятдесят кадильниць, і ти та Аарон, кожен кадильницю свою.
NUM|16|18|І взяли кожен кадильницю свою, і поклали на них огню, і поклали на неї кадила, та й стали при вході скинії заповіту, а також Мойсей та Аарон.
NUM|16|19|І Корей зібрав на них усю громаду до входу скинії заповіту. І показалася слава Господня всій громаді!
NUM|16|20|І промовив Господь до Мойсея та до Аарона, говорячи:
NUM|16|21|Відділіться від цієї громади, Я винищу їх умить!
NUM|16|22|А вони попадали на обличчя свої та й сказали: Боже, Боже духів і кожного тіла! Як згрішить один чоловік, чи Ти будеш гніватися на всю громаду?
NUM|16|23|І Господь промовляв до Мойсея, говорячи:
NUM|16|24|Скажи до громади, говорячи: Відступіться зо всіх боків від місця мешкання Корея, Датана й Авірона!
NUM|16|25|І встав Мойсей, і пішов до Датана та Авірона, і пішли за ним старші Ізраїлеві.
NUM|16|26|І він промовляв до громади, говорячи: Відступіть від наметів тих несправедливих людей, і не доторкніться до всього, що їхнє, щоб і ви не загинули за всі їхні гріхи!
NUM|16|27|І вони відступилися від місця мешкання Корея, Датана й Авірона зо всіх боків; а Датан та Авірон вийшли, і стояли при вході наметів своїх, і жінки їх, і сини їх, та діти їхні.
NUM|16|28|І сказав Мойсей: Оцим пізнаєте, що Господь послав мене зробити всі діла ці, що вони не з моєї вигадки.
NUM|16|29|Якщо вони повмирають, як умирає кожна людина, і їх спіткає доля кожної людини, то не Господь послав мене!
NUM|16|30|А коли Господь створить щось нове, і земля відкриє уста свої та й поглине їх та все, що їхнє, і вони зійдуть живі до шеолу, то пізнаєте, що люди образили Господа.
NUM|16|31|І сталося, як скінчив він говорити всі ці слова, то розступилася та земля, що під ними!
NUM|16|32|А земля відкрила свої уста, та й поглинула їх, і доми їхні, і кожну людину, що Кореєва, та ввесь їх маєток.
NUM|16|33|І зійшли вони та все, що їхнє, живі до шеолу, і накрила їх земля, і вони погинули з-посеред збору!
NUM|16|34|А ввесь Ізраїль, що був навколо них, повтікав на їхній крик, бо казали: Щоб земля не поглинула й нас!
NUM|16|35|І вийшов огонь від Господа, та й поїв тих двісті й п'ятдесят чоловіка, що приносили кадило!
NUM|16|36|(17-1) І Господь промовляв до Мойсея, говорячи:
NUM|16|37|(17-2) Скажи до Елеазара, сина священика Аарона, і нехай він позбирає ті кадильниці з-посеред погорілища, а огонь повикидає геть, бо вони освятилися,
NUM|16|38|(17-3) кадильниці тих грішників, їхньою смертю. І нехай і вони зроблять із них биті бляхи на покриття для жертівника, бо приносили їх перед Господнє лице, і вони освятилися. І будуть вони знаком для Ізраїлевих синів.
NUM|16|39|(17-4) І взяв священик Елеазар мідяні кадильниці, що приносили їх ті, що спалені, і перекували їх на покриття для жертівника,
NUM|16|40|(17-5) пам'ятка для Ізраїлевих синів, щоб чужий чоловік, хто не з Ааронового насіння, не наближався кадити кадило перед Господнім лицем, щоб не сталося з ними, як із Кореєм та з громадою його, як Господь говорив йому через Мойсея.
NUM|16|41|(17-6) А назавтра вся громада Ізраїлевих синів нарікали на Мойсея та на Аарона, говорячи: Ви повбивали Господній народ!
NUM|16|42|(17-7) І сталося, коли громада збиралася на Мойсея та на Аарона, то обернулися вони до скинії заповіту, аж ось покрила її хмара, і показалася слава Господня!
NUM|16|43|(17-8) І ввійшли Мойсей та Аарон до переду скинії заповіту.
NUM|16|44|(17-9) І Господь промовляв до Мойсея, говорячи:
NUM|16|45|(17-10) Вийдіть з-посеред цієї громади, а Я винищу їх умить! І вони попадали на обличчя свої.
NUM|16|46|(17-11) І сказав Мойсей до Аарона: Візьми кадильницю, і поклади на неї огню від жертівника, і поклади кадила, та й понеси швидко до громади, та й очисть її, бо вийшов гнів від Господнього лиця, і розпочалася поразка.
NUM|16|47|(17-12) І взяв Аарон, як говорив Мойсей, і побіг до середини зборів, аж ось розпочалася поразка народу! І він поклав кадила, і очистив народ.
NUM|16|48|(17-13) І став він поміж умерлими та поміж живими, і затрималась та поразка.
NUM|16|49|(17-14) І було померлих поразкою чотирнадцять тисяч і сімсот, окрім померлих у справі Корея.
NUM|16|50|(17-15) І вернувся Аарон до Мойсея до входу скинії заповіту, а поразка припинилася.
NUM|17|1|(17-16) І Господь промовляв до Мойсея, говорячи:
NUM|17|2|(17-17) Промовляй до Ізраїлевих синів, і візьми від них по одній палиці для батьківського дому, від усіх їхніх начальників для дому їхніх батьків, дванадцять палиць; і напиши ймення кожного на палиці його.
NUM|17|3|(17-18) А Ааронове ймення напишеш на Левієвій палиці, бо одна палиця для голови дому батьків їх.
NUM|17|4|(17-19) І покладеш їх у скинії заповіту перед ковчегом свідоцтва, де Я, за умовою, буду являтися вам.
NUM|17|5|(17-20) І станеться, той чоловік, що Я виберу його, його палиця зацвіте. І Я відхилю від Себе нарікання Ізраїлевих синів, що вони нарікають на вас.
NUM|17|6|(17-21) І Мойсей промовляв до Ізраїлевих синів, і дали йому всі їхні начальники по палиці від кожного начальника для дому їхніх батьків, дванадцять палиць. А палиця Ааронова серед їхніх палиць.
NUM|17|7|(17-22) І поклав Мойсей ті палиці перед Господнім лицем у скинії заповіту.
NUM|17|8|(17-23) І сталося назавтра, і ввійшов Мойсей до скинії заповіту, аж ось зацвіла Ааронова палиця для Левієвого дому, і пустила пуп'янки, і зацвіла квіткою, і випустила дозрілі мигдалі!
NUM|17|9|(17-24) І виніс Мойсей усі ті палиці з-перед Господнього лиця до всіх Ізраїлевих синів, і вони побачили, і взяли кожен свою палицю.
NUM|17|10|(17-25) І сказав Господь до Мойсея: Верни Ааронову палицю до ковчегу свідоцтва, щоб берегти на ознаку для неслухняних синів, і спиниш їхні нарікання проти Мене, щоб не повмирали вони.
NUM|17|11|(17-26) І зробив так Мойсей, як Господь наказав був йому, так він і зробив.
NUM|17|12|(17-27) І сказали Ізраїлеві сини до Мойсея, говорячи: Тож ми повмираємо, погинемо, усі ми погинемо!
NUM|17|13|(17-28) Кожен, хто наблизиться до Господньої скинії, помре. Чи ж ми дорешти вимремо?
NUM|18|1|І сказав Господь до Аарона: Ти й сини твої та дім батька твого з тобою понесете на собі гріх щодо святині; і ти, і сини твої з тобою понесете на собі гріх щодо вашого священства.
NUM|18|2|А також ти наблизиш до себе братів своїх, плем'я Левіїне, плем'я батька свого, і вони злучаться з тобою, і будуть прислужувати тобі, а ти й сини твої з тобою будете перед скинією свідоцтва.
NUM|18|3|І будуть вони виконувати твою сторожу та строжу всієї скинії, тільки до речей святині та до жертівника не приступлять, щоб не повмирали як вони, так і ви.
NUM|18|4|І злучаться вони з тобою, і будуть виконувати сторожу скинії заповіту, для всякої служби в скинії, а чужий не приступить до вас.
NUM|18|5|І будете ви виконувати сторожу святині та сторожу жертівника, щоб не було вже гніву на Ізраїлевих синів.
NUM|18|6|А Я оце взяв ваших братів Левитів з-посеред Ізраїлевих синів для вас, як дар вони дані Господеві, щоб виконувати службу скинії заповіту.
NUM|18|7|А ти та сини твої з тобою будете допильновувати ваше священство для всякої речі жертівника та для того, що поза завісою, і будете робити. Як службу дару даю Я священство вам, а чужий, хто приступить, буде забитий.
NUM|18|8|І Господь промовляв до Аарона: Я оце доручив тобі пильнувати за приношеннями Моїми. Від усього посвяченого синами Ізраїлевими Я дав частку тобі та для синів твоїх на вічну постанову.
NUM|18|9|Оце буде тобі з найсвятіших жертов, без огню: кожна їхня хлібна жертва, і кожна їхня жертва за гріх, і кожна їхня жертва за провину, що звернуть Мені як найсвятіше, тобі це та для твоїх синів!
NUM|18|10|На найсвятішому місці будеш ти їсти оце. Кожен чоловічої статі буде їсти, це буде святість для тебе.
NUM|18|11|А це тобі приношення їхнього дару всіх колихань Ізраїлевих синів, Я дав їх тобі, і синам твоїм та дочкам твоїм з тобою на вічну постанову, кожен чистий у твоїм домі буде це їсти.
NUM|18|12|Усе найкраще зо свіжої оливи, і все найкраще з молодого вина та збіжжя, їхні первоплоди, що вони дадуть Господеві, Я віддав їх тобі.
NUM|18|13|Первоплоди усього, що в їхньому Краю, що вони принесуть Господеві, будуть для тебе, кожен чистий у твоїм домі буде те їсти.
NUM|18|14|Усе закляте між Ізраїлем буде тобі.
NUM|18|15|Усе, що розкриває утробу кожного тіла, що принесуть Господеві з-поміж людей та з-поміж скотини, буде для тебе. Тільки конче викупиш перворідного людини, і перворідне з нечистої худобини викупиш.
NUM|18|16|А викуп його: від місячного віку викупиш за твоєю оцінкою, п'ять шеклів срібла на міру шеклем святині, двадцять ґер він.
NUM|18|17|Тільки перворідного з волів, або перворідного з овечок, або перворідного з кіз не викупиш, вони святість: їхньою кров'ю окропиш жертівника, а їхній лій спалиш, як огняну жертву на любі пахощі для Господа.
NUM|18|18|А їхнє м'ясо буде для тебе, як грудина колихання, і як стегно правиці буде для тебе.
NUM|18|19|Усі святощі приношення, що Ізраїлеві сини принесуть для Господа, Я віддав тобі, і синам твоїм та дочкам твоїм із тобою, вічною постановою. Це міцний заповіт, він вічний перед Господнім лицем для тебе та для насіння твого з тобою.
NUM|18|20|І сказав Господь до Аарона: У їхньому Краю ти не будеш мати власности, і не буде тобі частки між ними, Я частка твоя та власність твоя поміж Ізраїлевими синами!
NUM|18|21|А Левієвим синам Я дав ось кожну десятину в Ізраїлі на спадщину, взамін за їхню службу, бо вони виконують службу скинії заповіту.
NUM|18|22|І Ізраїлеві сини не приступлять уже до скинії заповіту, щоб не понести гріха, і не вмерти.
NUM|18|23|І буде Левит сам виконувати службу скинії заповіту, і сам понесе вину свою. Це вічна постанова для ваших поколінь, а між Ізраїлевими синами не будуть вони дідичити спадщину,
NUM|18|24|бо десятину Ізраїлевих синів, що вони принесуть як приношення для Господа, Я дав Левитам за спадщину. Тому Я сказав до них: Між Ізраїлевими синами не будуть вони дідичити спадщину.
NUM|18|25|І Господь промовляв до Мойсея, говорячи:
NUM|18|26|А до Левитів будеш ти промовляти та й скажеш їм: Коли візьмете від Ізраїлевих синів ту десятину, що Я дав вам від них на ваше спадщину, то ви принесете з неї Господнє приношення, десятину з десятини.
NUM|18|27|І буде пораховане ваше приношення як збіжжя з току, і як повня з кадки чавила.
NUM|18|28|Так принесете й ви Господнє приношення зо всіх ваших десятин, що візьмете від Ізраїлевих синів, і дасте з того Господнє приношення священикові Ааронові.
NUM|18|29|Зо всіх ваших дарів принесе кожен Господнє приношення, зо всього найкращого посвячення з нього.
NUM|18|30|І скажи їм: коли ви будете приносити найкраще з нього, то це порахується Левитам, як урожай току, і як урожай кадки чавила.
NUM|18|31|І будете їсти це на кожному місці ви та дім ваш, бо це нагорода для вас взамін за вашу службу в скинії заповіту.
NUM|18|32|І ви не понесете через це гріха, коли будете приносити найкраще з нього, а святощів Ізраїлевих синів не збезчестите, і не повмираєте.
NUM|19|1|І Господь промовляв до Мойсея та до Аарона, говорячи:
NUM|19|2|Промовляй до Ізраїлевих синів, і нехай вони візьмуть для тебе безвадну руду ялівку, що в ній нема вади, що на неї не накладали ярма.
NUM|19|3|І дасте її до священика Елеазара, а він виведе її поза табір. І заріжуть її перед ним.
NUM|19|4|І візьме Елеазар пальцем своїм її крови, та й покропить кров'ю її перед скинії заповіту сім раз.
NUM|19|5|І спалиться та ялівка на його очах, шкура її, і м'ясо її, і кров її з її нечистостями спалиться.
NUM|19|6|І візьме священик кедрове дерево, і ісоп та червень, та й кине до середини погорілища тієї ялівки.
NUM|19|7|І випере той священик шати свої та обмиє тіло своє в воді, а потім увійде до табору. І буде той священик нечистий аж до вечора.
NUM|19|8|А той, хто палить її, випере одежу свою в воді й обмиє тіло своє в воді, та й буде нечистий аж до вечора.
NUM|19|9|І збере чистий чоловік попіл тієї ялівки, і покладе поза табором в чистому місці, і буде це для громади Ізраїлевих синів на сховок для очищальної води, це жертва за гріх.
NUM|19|10|А той, хто збирає попіл тієї ялівки, випере одежу свою, і буде нечистий аж до вечора. І це буде на вічну постанову для Ізраїлевих синів та для приходька, що мешкає серед них тимчасово.
NUM|19|11|А той, хто доторкається до всякого мертвого тіла людини, то буде нечистий сім день.
NUM|19|12|Він очиститься тим попелом дня третього та дня сьомого, і буде чистий. А якщо він не очиститься дня третього та дня сьомого, не буде чистий.
NUM|19|13|Кожен, хто доторкується до померлого, до тіла людини, що померла, і не очиститься, він занечистив Господню скинію, і буде винищена душа та з Ізраїля, бо очищальна вода не була покроплена на нього, нечистий він буде, нечистість його в ньому.
NUM|19|14|Оце той закон: коли в наметі помре людина, то кожен, хто входить до того намету, та все, що в наметі, буде нечисте сім день.
NUM|19|15|І кожна відкрита посудина, що на ній нема міцно прив'язаного накриття, нечиста вона.
NUM|19|16|А кожен, хто доторкнеться на поверхні поля до трупа від меча, або до померлого, або до костей людини, або до гробу, буде нечистий сім день.
NUM|19|17|І візьмуть для того нечистого пороху з погорілища жертви за гріх, і наллють на нього живої води до посуду.
NUM|19|18|А чистий чоловік візьме ісопу, і вмочить у ту воду, та й покропить на того намета, і на всі посудини, і на душі ті, що були там, та на того, хто доторкується до тієї кістки, або до трупа, або до померлого, або до гробу.
NUM|19|19|І покропить той чистий на нечистого дня третього та дня сьомого, та й очистить його сьомого дня. І випере він одежу свою й обмиє в воді, і стане чистий увечері.
NUM|19|20|А чоловік, що стане нечистим і не очиститься, то буде знищена душа та з-посеред збору, бо він занечистив Господню святиню, очищальна вода не була кроплена на нього, нечистий він.
NUM|19|21|І буде це для них на вічну постанову, а той, хто кропить очищальну воду, випере одежу свою, а хто доторкається до очищальної води, буде нечистий аж до вечора.
NUM|19|22|А кожен, до кого доторкнеться нечистий, буде нечистий, а особа, що доторкується, буде нечиста аж до вечора.
NUM|20|1|І ввійшли Ізраїлеві сини, уся громада, до пустині Цін першого місяця, та й засів народ у Кадеші. І померла там Маріям, і була там похована.
NUM|20|2|І не було води для громади, і вони зібралися проти Мойсея та проти Аарона.
NUM|20|3|І сварився той народ із Мойсеєм, та й сказали, говорячи: О, якби ми повмирали були, коли наші брати вмирали перед Господнім лицем!
NUM|20|4|І нащо ви привели Господню громаду на цю пустиню, щоб повмирали тут ми та худоба наша?
NUM|20|5|І нащо ви вивели нас із Єгипту, щоб привести нас на це зле місце? Тут не родить збіжжя, ані фіґи, ані виноград, ані гранатове яблуко, і навіть немає напитись води!
NUM|20|6|І ввійшли Мойсей та Аарон від громади до входу скинії заповіту, та й попадали на обличчя свої. І слава Господня появилася їм!
NUM|20|7|І Господь промовляв до Мойсея, говорячи:
NUM|20|8|Візьми жезло, та збери громаду ти та брат твій Аарон, і скажете до тієї скелі на їхніх очах, і вона дасть свою воду. І виведеш для них воду з тієї скелі, та й напоїш ту громаду та їхню худобу.
NUM|20|9|І взяв Мойсей те жезло з-перед Господнього лиця, як Він наказав був йому.
NUM|20|10|І зібрали Мойсей та Аарон громаду перед тією скелею. І сказав він до них: Послухайте ж, неслухняні, чи з цієї скелі ми виведемо для вас воду?
NUM|20|11|І підніс Мойсей руку свою, та й ударив ту скелю своїм жезлом два рази, і вийшло багато води! І пила громада та їхня худоба!...
NUM|20|12|І сказав Господь до Мойсея та до Аарона: За те, що ви не ввірували в Мене, щоб явилася святість Моя на очах Ізраїлевих синів, ви не введете цієї громади до Краю, що Я дав їм.
NUM|20|13|Це вода Меріви, де сварилися Ізраїлеві сини з Господом, і святість Його явилася їм.
NUM|20|14|І послав Мойсей послів із Кадешу до царя едомського сказати: Так каже брат твій Ізраїль: Ти знаєш усю тяготу, що впала на нас.
NUM|20|15|І зійшли були наші батьки до Єгипту, і сиділи ми в Єгипті багато часу, а Єгипет чинив зло нам та батькам нашим.
NUM|20|16|І голосили ми до Господа, і Він почув наш голос, та й послав Ангола, і вивів нас із Єгипту, а оце ми в Кадеші, що при самім кінці твоєї границі.
NUM|20|17|Нехай же ми перейдемо через твій край! Ми не підемо полем та виноградником, і не будемо пити води з криниці, ми підемо дорогою царською, не збочимо ні праворуч, ні ліворуч, аж поки не перейдемо границі твоєї.
NUM|20|18|І сказав до нього Едом: Ти не перейдеш у мене, бо інакше я з мечем вийду проти тебе!
NUM|20|19|І сказали йому Ізраїлеві сини: Ми підемо битою дорогою, а якщо будемо пити воду твою я та худоба моя, то я дам заплату за неї. Нічого більше, тільки нехай перейду я своїми ногами!
NUM|20|20|А той відказав: Не перейдеш! І вийшов Едом навпроти нього з численним народом та з сильною рукою.
NUM|20|21|І відмовив Едом дати Ізраїлеві перейти його границі, і Ізраїль збочив від нього.
NUM|20|22|І рушили з Кадешу, і вийшли Ізраїлеві сини, уся громада, до Гор-гори.
NUM|20|23|І сказав Господь до Мойсея та до Аарона на Гор-горі, на границі едомського краю, говорячи:
NUM|20|24|Нехай прилучиться Аарон до своєї рідні, бо він не ввійде до того Краю, що Я дав Ізраїлевим синам, через те, що ви були неслухняні наказу Моєму при воді Меріви.
NUM|20|25|Візьми Аарона та сина його Елеазара, та й виведи їх на Гор-гору.
NUM|20|26|І нехай Аарон здійме шати свої, і зодягне в них сина свого Елеазара, і Аарон буде забраний, та й помре там.
NUM|20|27|І зробив Мойсей, як Господь наказав був, і вийшли вони на Гор-гору на очах усієї громади.
NUM|20|28|І зняв Мойсей з Аарона шати його, і зодягнув у них сина його Елеазара, і Аарон помер там на верхів'ї гори. І зійшов Мойсей та Елеазар із гори.
NUM|20|29|І бачила вся громада, що помер Аарон, і оплакував Аарона ввесь Ізраїлів дім тридцять день.
NUM|21|1|І почув ханаанеянин, цар Араду, що сидів на полудні, що Ізраїль увійшов дорогою Атарім, і він став воювати з Ізраїлем, і взяв у нього до неволі полонених.
NUM|21|2|І склав Ізраїль обітницю Господеві й сказав: Якщо справді даси Ти народ той у мою руку, то я вчиню їхні міста закляттям.
NUM|21|3|І вислухав Господь голос Ізраїлів, і дав йому ханаанеянина, і він учинив закляттям їх та їхні міста, і назвав ім'я тому міста: Хорма.
NUM|21|4|І рушили вони з Гор-гори дорогою Червоного моря, щоб обійти едомський край. І підупала душа того народу в тій дорозі.
NUM|21|5|І промовляв той народ проти Бога та проти Мойсея: Нащо ви вивели нас із Єгипту, щоб ми повмирали в пустині? Бож нема тут хліба й нема води, а душі нашій обридла ця непридатна їжа.
NUM|21|6|І послав Господь на той народ зміїв сарафів, і вони кусали народ. І померло багато народу з Ізраїля.
NUM|21|7|І прийшов народ до Мойсея та й сказав: Згрішили ми, бо говорили проти Господа та проти тебе. Молися до Господа, і нехай Він забере від нас цих зміїв. І молився Мойсей за народ.
NUM|21|8|І сказав Господь до Мойсея: Зроби собі сарафа, і вистав його на жердині. І станеться, кожен покусаний, як погляне на нього, то буде жити.
NUM|21|9|І зробив Мойсей мідяного змія, і виставив його на жердині. І сталося, якщо змій покусав кого, то той дивився на мідяного змія і жив!
NUM|21|10|І рушили Ізраїлеві сини, і таборували в Овоті.
NUM|21|11|І рушили вони з Овоту, і таборували в Ійє-Гааварімі, на пустині, що перед Моавом, від сходу сонця.
NUM|21|12|Звідти вони рушили, і таборували в долині Зереду.
NUM|21|13|Звідти рушили й таборували на тім боці Арнону в пустині, що виходить із аморейської границі, бо Арнон границя Моаву між Моавом та амореянином.
NUM|21|14|Тому розповідається в Книжці воєн Господніх: Вагев у Суфі, і потоки Арнону,
NUM|21|15|і спад потоків, що збочив на місце Ару, і на моавську границю опертий.
NUM|21|16|А звідти до Бееру. Це той Беер, що про нього сказав Господь до Мойсея: Збери народ, і нехай Я дам їм воду.
NUM|21|17|Тоді заспівав був Ізраїль цю пісню: Піднесися, кринице, співайте про неї!
NUM|21|18|Криниця, вельможі копали її, її викопали народні достойники берлом, жезлами своїми. А з Мідбару до Маттани,
NUM|21|19|а з Маттани до Нахаліїлу, а з Нахаліїлу до Бамоту,
NUM|21|20|а з Бамоту до долини, що на моавському полі, у верхівки Пісґі, що звернена до пустині.
NUM|21|21|І послав Ізраїль послів до Сигона аморейського царя, говорячи:
NUM|21|22|Нехай я перейду в твоїм краї! Ми не збочимо ні на поле, ні на виноградник, не будемо пити води з криниці, ми підемо царською дорогою, аж поки перейдемо землю твою.
NUM|21|23|І не дав Сигон Ізраїлеві перейти в границі його. І зібрав Сигон увесь свій народ, та й вийшов навпроти Ізраїля на пустині, і прибув до Йогці, і воював з Ізраїлем.
NUM|21|24|І вдарив його Ізраїль вістрям меча, і посів край його від Арнону аж до Яббоку, аж до синів Аммону, бо Аз границя синів Аммону.
NUM|21|25|І позабирав Ізраїль усі ті міста. І осів Ізраїль у всіх аморейських містах: у Хешбоні й по всіх залежних містах його.
NUM|21|26|Бо Хешбон місто Сигона, царя аморейського він; і він воював з першим моавським царем, і забрав увесь його край з його руки аж до Арнону.
NUM|21|27|Тому й розповідають кобзарі: Підіть до Хешбону, нехай він збудується, і хай міцно поставиться місто Сигонове.
NUM|21|28|Бо вийшов огонь із Хешбону, а полум'я з міста Сигонового, він місто моавське пожер, володарів арнонських висот.
NUM|21|29|Горе тобі, о Моаве, ти згинув, народе Кемошів! Він зробив був синів своїх утікачами, а дочок своїх дав у неволю Сигону, царю аморейському.
NUM|21|30|І розбили ми їх, згинув Хешбон до Дівону, і ми попустошили аж до Нофаху, що аж до Медви.
NUM|21|31|І Ізраїль осів в аморейському краї.
NUM|21|32|І послав Мойсей розвідати про Язера, і вони здобули його залежні міста, і заволоділи амореянином, що жив там.
NUM|21|33|І повернулись вони, і пішли дорогою Башану. І вийшов Оґ, цар башанський, насупроти них, він та ввесь його народ, на війну до Едреї.
NUM|21|34|І сказав Господь до Мойсея: Не бійся його, бо в руку твою дав Я його й увесь народ його та край його, і зробиш йому, як зробив ти Сигону, цареві аморейському, що сидів у Хешбоні.
NUM|21|35|І вони побили його й синів його та ввесь народ його, так що нікого не зосталося. І вони заволоділи краєм його.
NUM|22|1|І рушили Ізраїлеві сини, та й таборували в моавських степах по тім боці приєрихонського Йордану.
NUM|22|2|І побачив Балак, син Ціппорів, усе, що зробив Ізраїль амореянинові.
NUM|22|3|І дуже злякався Моав того народу, бо він був великий. І настрашився Моав Ізраїлевих синів.
NUM|22|4|І сказав Моав до мідіянських старших: Тепер повискубує оця громада всі наші околиці, як вискубує віл польову зеленину. А Балак, син Ціппорів, був того часу моавським царем.
NUM|22|5|І послав він послів до Валаама, Беорового сина, до Петору, що над Річкою, до краю синів народу його, щоб покликати його, говорячи: Ось вийшов народ із Єгипту, ось покрив він поверхню землі, і сидить навпроти мене.
NUM|22|6|А тепер ходи ж, прокляни мені цей народ, бо він міцніший за мене. Може я потраплю вдарити його, і вижену його з краю, бо знаю, що кого ти поблагословиш, той благословенний, а кого проклянеш, проклятий.
NUM|22|7|І пішли моавські старші та старші Мідіяну, а дарунки за чари в руці їх, і прийшли до Валаама, та й промовляли до нього Балакові слова.
NUM|22|8|А він їм сказав: Ночуйте тут цієї ночі, і я перекажу вам слово, як Господь промовлятиме до мене. І зостались моавські вельможі в Валаама.
NUM|22|9|І прийшов Бог до Валаама та й сказав: Хто ці люди з тобою?
NUM|22|10|І сказав Валаам до Бога: Балак, син Ціппорів, цар моавський, послав до мене сказати:
NUM|22|11|Ось народ виходить з Єгипту, і закрив поверхню землі; тепер іди ж, прокляни мені його, може я потраплю воювати з ним, і вижену його.
NUM|22|12|І сказав Бог до Валаама: Не підеш ти з ними, не проклянеш того народу, бо благословенний він!
NUM|22|13|І встав Валаам уранці та й сказав до Балакових вельмож: Вертайтесь до свого краю, бо відмовив Господь позволити мені піти з вами.
NUM|22|14|І встали моавські вельможі, і прийшли до Балака та й сказали: Відмовив Валаам піти з нами.
NUM|22|15|А Балак знову послав вельмож, більше й поважніших від тих.
NUM|22|16|І прибули вони до Валаама та й сказали йому: Так сказав Балак, син Ціппорів: Не стримуйся прийти до мене,
NUM|22|17|бо справді дуже вшаную тебе, і все, що скажеш мені, зроблю. І ходи ж, прокляни мені народ той!
NUM|22|18|І відповів Валаам, і сказав Балаковим рабам: Якщо Балак дасть мені повний свій дім срібла та золота, то й тоді я не зможу переступити наказу Господа, Бога мого, щоб зробити річ малу чи річ велику.
NUM|22|19|А тепер посидьте й ви тут цієї ночі, а я пізнаю, що ще Господь буде говорити мені.
NUM|22|20|І прийшов Бог уночі до Валаама та й сказав йому: Якщо ці люди прийшли покликати тебе, устань, іди з ними. Але тільки те, що Я промовлятиму до тебе, те ти зробиш.
NUM|22|21|І встав Валаам уранці, і осідлав свою ослицю, та й пішов із моавськими вельможами.
NUM|22|22|І запалився гнів Божий, що він іде. І став Ангол Господній на дорозі за перешкоду йому, а він їде на своїй ослиці, і двоє слуг його з ним.
NUM|22|23|І побачила та ослиця Господнього Ангола, що стоїть на дорозі, а витягнений меч його в руці його. І збочила ослиця з дороги, і пішла полем, а Валаам ударив ослицю, щоб збочила на дорогу.
NUM|22|24|І став Ангол Господній на стежці виноградників, стіна з цієї сторони, і стіна з тієї.
NUM|22|25|І побачила та ослиця Господнього Ангола, і притиснулася до стіни, та й притиснула до стіни Валаамову ногу. І він далі її бив.
NUM|22|26|І Ангол Господній знов перейшов, і став у тісному місці, де нема дороги збочити ні праворуч, ні ліворуч.
NUM|22|27|І побачила та ослиця Господнього Ангола і лягла під Валаамом. І запалився гнів Валаамів, і він ударив ослицю києм.
NUM|22|28|І відкрив Господь уста ослиці, і сказала вона до Валаама: Що я зробила тобі, що ти оце тричі вдарив мене?
NUM|22|29|І сказав Валаам до ослиці: Бо ти виставила мене на сміх. Коли б меч був у руці моїй, то тепер я забив би тебе!
NUM|22|30|І сказала ослиця до Валаама: Чи ж я не ослиця твоя, що ти їздив на мені, скільки живеш, аж до цього дня? Чи ж справді звикла я робити тобі так? І він відказав: Ні!
NUM|22|31|І відкрив Господь очі Валаамові, і побачив він Господнього Ангола, що стоїть на дорозі, а його витягнений меч у руці його. І схилився він, і впав на обличчя своє.
NUM|22|32|І сказав до нього Ангол Господній: Нащо ти вдарив ослицю свою оце тричі? Ось я вийшов за перешкоду, бо ця дорога погибельна передо мною.
NUM|22|33|І побачила мене ця ослиця, і збочила перед лицем моїм ось власне тричі. І коли б вона не збочила була перед лицем моїм, то тепер я й забив би тебе, а її позоставив би живою.
NUM|22|34|І сказав Валаам до Господнього Ангола: Я згрішив, бо не знав, що ти стоїш на дорозі навпроти мене. А тепер, якщо це зле в очах твоїх, то я вернуся собі.
NUM|22|35|І сказав Ангол Господній до Валаама: Іди з цими людьми, і те слово, що скажу тобі, його тільки будеш говорити. І пішов Валаам з Балаковими вельможами.
NUM|22|36|І почув Балак, що прийшов Валаам, і вийшов навпроти нього до Їр-Моаву, що на границі Арнону, що на краю границі.
NUM|22|37|І сказав Балак до Валаама: Чи ж справді не послав я до тебе, щоб покликати тебе, чому ж не пішов ти до мене? Чи справді я не потраплю вшанувати тебе?
NUM|22|38|І сказав Валаам до Балака: Ось я прибув до тебе тепер. Чи потраплю я сказати щось? Те слово, що Бог вкладе в уста мої, його тільки я буду промовляти.
NUM|22|39|І пішов Валаам із Балаком, і прибули вони до Кір'ят-Хуцоту.
NUM|22|40|І приніс Балак на жертву худобу велику та худобу дрібну, і послав Валаамові та вельможам, що з ним.
NUM|22|41|І сталося вранці, і взяв Балак Валаама, та й вивів його на Бамот-Баал, щоб побачив ізвідти тільки частину того народу.
NUM|23|1|І сказав Валаам до Балака: Збудуй мені тут сім жертівників, і приготуй мені тут сім бичків та сім баранів.
NUM|23|2|І зробив Балак, як Валаам говорив. І приніс Балак та Валаам бичка та барана на кожному жертівнику.
NUM|23|3|І сказав Валаам до Балака: Стань над своїм цілопаленням, а я піду, може стріну Господа навпроти себе, і що Він об'явить мені, я перекажу тобі. І він пішов на лису гору.
NUM|23|4|І стрівся Валаамові Бог, і сказав він Йому: Сім жертівників склав я, і приніс бичка та барана на кожному жертівнику.
NUM|23|5|І вклав Господь слово до Валаамових уст та й сказав: Вернись до Балака, і будеш так промовляти.
NUM|23|6|І вернувсь він до нього, аж ось він стоїть над своїм цілопаленням, він та всі вельможі моавські.
NUM|23|7|І він виголосив свою приповістку пророчу й сказав: Із Араму мене припровадив Балак, цар моавський, з гір сходу: Іди ж, прокляни мені Якова, а йди ж, скажи зло на Ізраїля!
NUM|23|8|Що ж я буду того проклинати, що Бог не прокляв був його? І що ж буду казать зло на того, що гніву на нього не має Господь?
NUM|23|9|Бо я бачу його з вершка скель, і з пагірків його оглядаю, тож народ пробуває самітно, а серед людей не рахується.
NUM|23|10|Хто ж перелічив порох Яковів, і хто зрахував пил Ізраїлів? Хай душа моя вмре смертю праведних, і кінець мій хай буде такий, як його!
NUM|23|11|І сказав Балак до Валаама: Що ти зробив мені? Я взяв тебе, щоб ти прокляв моїх ворогів, а оце ти справді поблагословив їх!
NUM|23|12|А той відповів та й сказав: Чи ж не те, що Господь вкладе в мої уста, я буду пильнувати, щоб те говорити?
NUM|23|13|І сказав до нього Балак: Ходи ж зо мною до іншого місця, звідки побачиш його. Тільки частину його будеш бачити, а всього його не побачиш. І прокляни мені його, мого ворога, звідти!
NUM|23|14|І він узяв його на Седе-Цофім, на верхів'я Пісґі, і збудував сім жертівників, і приніс бичка та барана на кожнім жертівнику.
NUM|23|15|І сказав він до Балака: Стань тут над своїм цілопаленням, а я стріну там Господа.
NUM|23|16|І стрів Господь Валаама, і вклав слово до уст його та й сказав: Вернися до Балака, і будеш так промовляти.
NUM|23|17|І прийшов він до нього, аж ось він стоїть над своїм цілопаленням, а з ним вельможі моавські. І сказав йому Балак: Що ж говорив Господь?
NUM|23|18|І він виголосив свою приповістку пророчу й сказав: Устань же, Балаку, та й слухай, нахили своє ухо до мене, о сину Ціппорів!
NUM|23|19|Бог не чоловік, щоб неправду казати, і Він не син людський, щоб Йому жалкувати. Чи ж Він був сказав і не зробить, чи ж Він говорив та й не виконає?
NUM|23|20|Оце я одержав наказа поблагословити, і поблагословив Він, і я того не відверну!
NUM|23|21|Не видно страждання між Яковом, і не запримітно нещастя в Ізраїлі, з ним Господь, його Бог, а між ним голосний крик на славу Царя!
NUM|23|22|Бог, що вивів був їх із Єгипту, Він для нього, як міць однорожця!
NUM|23|23|Бо нема ворожби поміж Яковом, і чарів нема між Ізраїлем, тепер буде сказане Якову та Ізраїлеві, що Бог учинив.
NUM|23|24|Тож устане народ, як левиця, і підійметься він, немов лев! Він не ляже, аж поки не буде він жерти здобичу, і аж поки не буде він пить кров забитих!
NUM|23|25|І сказав Балак до Валаама: Ні проклинати не проклинай його, ні благословити не благословляй його!
NUM|23|26|І сказав Валаам, і відповів до Балака: Чи ж не казав я тобі, говорячи: Усе, що буде промовляти Господь, те зроблю?
NUM|23|27|І сказав Балак до Валаама: Ходи ж, візьму тебе ще до іншого місця, може сподобається в Божих очах, і ти звідти проклянеш мені його.
NUM|23|28|І взяв Балак Валаама на верхів'я Пеору, що звернений до пустині.
NUM|23|29|І сказав Валаам до Балака: Збудуй мені тут сім жертівників, і приготуй мені тут сім бичків та сім баранів.
NUM|23|30|І зробив Балак, як сказав був Валаам, і приніс бичка та барана на кожному жертівнику.
NUM|24|1|І побачив Валаам, що Господеві вгодно поблагословити Ізраїля, і не пішов, як кожного разу, на ворожбу, і звернув лице своє до пустині.
NUM|24|2|І звів Валаам очі свої, та й побачив Ізраїля, що пробував за своїми племенами. І на ньому був Дух Божий!
NUM|24|3|І він виголосив свою приповістку пророчу й сказав: Мова Валаама, сина Беорового, і мова мужа з очима відкритими,
NUM|24|4|це мова того, хто слухається Божих слів, хто бачить видіння Всемогутнього, що падає він, але очі відкриті йому.
NUM|24|5|Які, Якове, гарні намети твої, місця перебування твойого, Ізраїлю!
NUM|24|6|Вони розтяглися, немов ті долини, немов ті садки понад річкою, вони як дерева алойні, що Господь насадив, як кедри над водами!
NUM|24|7|Вода потече з його відер, а насіння його над великими водами. Його цар стане вищий за Аґаґа, і царство його піднесеться.
NUM|24|8|Із Єгипту Бог вивів його, Він для нього як міць однорожця! Поїсть він людей, що ворожі йому, і їхні кості потрощить, а стріли його поламає.
NUM|24|9|Нахилився він, ліг, немов лев, і як левиця, хто підійме його? Хто благословляє тебе той благословенний, а хто проклинає тебе той проклятий!
NUM|24|10|І запалав гнів Балаків на Валаама, і сплеснув він у долоні свої! І сказав Балак до Валаама: Я покликав тебе проклясти ворогів моїх, а ти ось, благословляючи, поблагословив їх оце тричі!
NUM|24|11|А тепер утікай собі до свого місця! Я сказав був: конче пошаную тебе, та ось стримав тебе Господь від пошани.
NUM|24|12|І сказав Валаам до Балака: Чи ж не казав я також до посланців твоїх, яких послав ти до мене, говорячи:
NUM|24|13|Якщо Балак дасть мені повний свій дім срібла та золота, то й тоді я не зможу переступити наказу Господнього, щоб зробити добре чи зле з власної волі, що казатиме Господь, те я буду говорити!
NUM|24|14|А тепер я оце йду до народу свого. Ходи ж, я звіщу тобі, що зробить той народ твоєму народові на кінці днів.
NUM|24|15|І він виголосив свою приповістку пророчу й сказав: Мова Валаама, сина Беорового, і мова мужа з очима відкритими,
NUM|24|16|мова того, хто слухається Божих слів, і знає думку Всевишнього, хто бачить видіння Всемогутнього, що падає він, але очі відкриті йому.
NUM|24|17|Я бачу його, та не тепер, дивлюся на нього, та він не близький! Сходить зоря он від Якова, і підіймається берло з Ізраїля, ламає він скроні Моава та черепа всіх синів Сифа!
NUM|24|18|І стане Едом за спадщину, і стане Сеїр за посілість своїх ворогів, а Ізраїль робитиме справи великі!
NUM|24|19|І той запанує, хто з Якова, і вигубить рештки із міста.
NUM|24|20|І побачив він Амалика, і виголосив свою приповістку пророчу й сказав: Початок народів Амалик, та загине наприкінці й він!
NUM|24|21|І побачив він кенеянина, і виголосив свою приповістку пророчу й сказав: Міцна ця оселя твоя, і поклав ти на скелі гніздо своє!
NUM|24|22|Але вигублений буде Каїн, незабаром Ашшур поневолить тебе!
NUM|24|23|І він виголосив свою приповістку пророчу й сказав: О, хто ж буде жити, як зачне Бог робити оце?
NUM|24|24|І кораблі припливуть від кіттеїв, і Ашшура впокорять, і Евера впокорять. Та загине наприкінці й він!
NUM|24|25|І встав Валаам і пішов, та й вернувся до місця свого. А Балак також пішов на дорогу свою.
NUM|25|1|І осівся Ізраїль у Шіттімі, і народ зачав ходити на розпусту до моавських дочок,
NUM|25|2|а вони закликали народ до жертов їхнім богам, і народ їв та вклонявся богам їхнім.
NUM|25|3|І Ізраїль приліпився був до пеорського Ваала. І запалав гнів Господній на Ізраїля.
NUM|25|4|І сказав Господь до Мойсея: Візьми всіх голів народу, та й повішай їх для Господа навпроти сонця. І відвернеться палючий Господній гнів від Ізраїля.
NUM|25|5|І сказав Мойсей до Ізраїлевих суддів: Позабивайте кожен мужів своїх, приліплених до пеорського Ваала.
NUM|25|6|Аж ось прийшов один із Ізраїлевих синів, та й привів до братів своїх мідіянітянку на очах Мойсея й на очах усієї громади Ізраїлевих синів, а вони плакали при вході скинії заповіту.
NUM|25|7|І побачив це Пінхас, син Елеазара, сина священика Аарона. І встав він з-посеред громади, і взяв списа в свою руку.
NUM|25|8|І ввійшов він за Ізраїлевим мужем до середини мешкання, та й пробив їх обох ізраїльтянина та ту жінку, аж через її черево. І була стримана поразка Ізраїлевих синів.
NUM|25|9|І померло в поразці двадцять і чотири тисячі.
NUM|25|10|І промовив Господь до Мойсея, говорячи:
NUM|25|11|Пінхас, син Елеазара, сина священика Аарона, відвернув Мою лють від Ізраїлевих синів, коли він запалився горливістю Моєю серед них. І Я не вигубив Ізраїлевих синів у Своїй горливості.
NUM|25|12|Тому скажи: ось Я даю йому свого заповіта: мир.
NUM|25|13|І буде йому та насінню його по нім заповіт вічного священства за те, що він запалився для Бога свого, і очистив Ізраїлевих синів.
NUM|25|14|А ймення забитого Ізраїлевого мужа, що був забитий з тією мідіянітянкою, Зімрі, син Салу, начальник батькового дому Симеона.
NUM|25|15|І ім'я тієї забитої мідіянітської жінки Козбі, дочка Цура, що був головою племен батькового дому в Мідіяні.
NUM|25|16|І Господь промовляв до Мойсея, говорячи:
NUM|25|17|Ненавидіти мідіянітів, і будете їх забивати!
NUM|25|18|Бож вони ненавидять вас у своїх підступах, що зводили вас через Пеора, і через Козбі, дочку мідіянітського начальника, сестру їх, забиту дня поразки за Пеора.
NUM|26|1|І сталося по поразці, і сказав Господь до Мойсея й до Елеазара, сина священика Аарона, говорячи:
NUM|26|2|Перелічіть усю громаду Ізраїлевих синів від віку двадцяти літ і вище за домами їхніх батьків, кожного, хто здатний до війська в Ізраїлі.
NUM|26|3|І говорив до них Мойсей та священик Елеазар у моавських степах над приєрихонським Йорданом, говорячи:
NUM|26|4|Перелічіть від віку двадцяти літ і вище, як наказав був Господь Мойсеєві і Ізраїлевим синам, що виходили з єгипетського краю.
NUM|26|5|Рувим, перворідний Ізраїлів. Рувимові сини: Ханох рід Ханохів, від Паллу рід Паллуїв,
NUM|26|6|від Хецрона рід Хецронів, від Кармі рід Карміїв.
NUM|26|7|Оце Рувимові роди. І були їхні перелічені: сорок і три тисячі й сімсот і тридцять.
NUM|26|8|А сини Паллуєві: Еліяв.
NUM|26|9|А сини Еліявові: Немуїл, і Датан, і Авірон. Це той Датан та Авірон, покликані громади, що підбурювали проти Мойсея та проти Аарона в Кореєвій громаді, коли вони підбурювали на Господа.
NUM|26|10|І відкрила земля свої уста, та й поглинула їх та Корея при смерті тієї громади, коли огонь пожер був двісті і п'ятдесят люда, і стали вони за ознаку.
NUM|26|11|А Кореєві сини не померли.
NUM|26|12|Сини Симеонові за їхніми родами: від Немуїла рід Немуїлів, від Яміна рід Ямінів, від Яхіна рід Яхінів,
NUM|26|13|від Зераха рід Зерахів, від Саула рід Саулів.
NUM|26|14|Оце Симеонові роди, двадцять і дві тисячі й двісті.
NUM|26|15|Сини Ґадові за їхніми родами: від Цефона рід Цефонів, від Хаґґі рід Хаґґіїв, від Шуні рід Шуніїв,
NUM|26|16|від Озні рід Озніїв, від Ері рід Еріїв,
NUM|26|17|від Арода рід Ародів, від Ар'елі рід Ар'еліїв.
NUM|26|18|Оце роди Ґадових синів, за їхнім переліченням: сорок тисяч і п'ятсот.
NUM|26|19|Сини Юдині: Ер та Онан; і помер Ер та Онан у ханаанськім Краї.
NUM|26|20|І були Юдині сини за їхніми родами: від Шели рід Шелин, від Переца рід Переців, від Зераха рід Зерахів.
NUM|26|21|А Перецеві сини були: від Хецрона рід Хецронів, від Хамула рід Хамулів.
NUM|26|22|Оце Юдини роди за їхнім переліченням: сімдесят і шість тисяч і п'ятсот.
NUM|26|23|Сини Іссахарові за їхніми родами: Тола рід Толин, від Цувви рід Цуввин,
NUM|26|24|від Яшува рід Яшувів, від Шімрона рід Шімронів.
NUM|26|25|Оце Іссахарові роди за їхнім переліченням: шістдесят і чотири тисячі й триста.
NUM|26|26|Сини Завулонові за їхніми родами: від Середа рід Середів, від Елона рід Елонів, від Яхлеїла рід Яхлеїлів.
NUM|26|27|Оце Завулонові роди за їхнім переліченням: шістдесят тисяч і п'ятсот.
NUM|26|28|Сини Йосипа за їхніми родами: Манасія та Єфрем.
NUM|26|29|Сини Манасіїні: від Махіра рід Махірів, а Махір породив Ґілеада, від Ґілеада рід Ґілеадів.
NUM|26|30|Оце Ґілеадові сини: Єзер рід Єзерів, від Хелека рід Хелеків,
NUM|26|31|і Асріїл рід Асріїлів, і Шехем рід Шехемів,
NUM|26|32|і Шеміда рід Шемідин, і Хефер рід Хеферів.
NUM|26|33|А Целофхад, син Хеферів, не мав синів, а тільки дочок. А ймення дочок: Махла й Ноа, Хоґла, Мілка й Тірца.
NUM|26|34|Оце роди Манасіїні, а їхні перелічені: п'ятдесят і дві тисячі й сімсот.
NUM|26|35|Оце Єфремові сини за їхніми родами: від Шутелаха рід Шутелахів, від Бехера рід Бехерів, від Тахана рід Таханів.
NUM|26|36|А оце Шутелахові сини: від Ерана рід Еранів.
NUM|26|37|Оце роди Єфремових синів за їхнім переліченням: тридцять і дві тисячі і п'ятсот. Оце Йосипові сини за їхніми родами.
NUM|26|38|Сини Веніяминові за їхніми родами: від Бели рід Белин, від Ашбела рід Ашбелів, від Ахірама рід Ахірамів,
NUM|26|39|від Шефуфама рід Шефуфамів, від Хуфама рід Хуфамів.
NUM|26|40|А сини Белині були: Ард, і Нааман, від Арда рід Ардів, від Наамана рід Нааманів.
NUM|26|41|Оце Веніяминові сини за їхніми родами, а перелічені їхні: сорок і п'ять тисяч і шістсот.
NUM|26|42|Оце Данові сини за їхніми родами: від Шухама рід Шухамів. Оце Данові роди за їхніми родами.
NUM|26|43|Всі Шухамові роди за їхнім переліченням: шістдесят і чотири тисячі і чотириста.
NUM|26|44|Асирові сини за їхніми родами: від Їмни рід Їмнин, від Їшві рід Їшвіїв, від Берії рід Беріїв.
NUM|26|45|Сини Берії: від Хевера рід Хеверів, від Малкіїла рід Малкіїлів,
NUM|26|46|а ймення Асирової дочки Сарах.
NUM|26|47|Оце роди Асирових синів за їхнім переліченням: п'ятдесят і три тисячі й чотириста.
NUM|26|48|Сини Нефталимові за їхніми родами: від Яхцеїла рід Яхцеїлів, від Ґуні рід Ґуніїв,
NUM|26|49|від Єцера рід Єцерів, від Шіллема рід Шіллемів.
NUM|26|50|Оце роди Нефталимові за їхніми родами й за їхнім переліченням: сорок і п'ять тисяч і чотириста.
NUM|26|51|Оце перелічені Ізраїлевих синів: шістсот тисяч і тисяча й сімсот і тридцять.
NUM|26|52|І промовив Господь до Мойсея, говорячи:
NUM|26|53|Для цих буде поділений Край у спадок за числом імен.
NUM|26|54|Численному примножиш спадщину його, а малому зменшиш спадок його, кожному за переліченням його буде дана спадщина його.
NUM|26|55|Тільки жеребком поділиться землю, вони будуть володіти за іменами племен їхніх батьків.
NUM|26|56|За жеребком буде поділена спадщина його поміж численним та малим.
NUM|26|57|А оце перелічені Левити за їхніми родами: від Ґершона рід Ґершонів, від Кегата рід Кегатів, від Мерарі рід Мераріїв.
NUM|26|58|Оце роди Левієві: рід Левіїв, рід Хевроніїв, рід Махліїв, рід Мушіїв, рід Кореїв, а Кегат породив Амрама.
NUM|26|59|А ймення Амрамової жінки Йохевед, дочка Левієва, що вродила її Левієві жінка його в Єгипті, а вона вродила Амрамові Аарона, і Мойсея, і сестру їх Маріям.
NUM|26|60|І вродилися Ааронові Надав, й Авігу, й Елеазар, й Ітамар.
NUM|26|61|А Надав та Авігу померли, коли вони приносили чужий огонь перед Господнє лице.
NUM|26|62|І були їхні перелічені двадцять і три тисячі, кожен чоловічої статі від місячного віку й вище; бо вони не були перелічені серед Ізраїлевих синів, не дана бо їм спадщина серед Ізраїлевих синів.
NUM|26|63|Оце перелічені Мойсея та священика Елеазара, що перелічували Ізраїлевих синів у моавських степах над приєрихонським Йорданом.
NUM|26|64|А серед тих не було вже нікого з перелічених Мойсея та священика Аарона, що перелічували Ізраїлевих синів на Сінайській пустині,
NUM|26|65|бо Господь був сказав їм: Конче повмираєте ви на пустині. І не позостався з них ніхто, крім Калева, сина Єфуннеєвого, та Ісуса, сина Навинового.
NUM|27|1|І прийшли дочки Целофхада, сина Хеферового, сина Ґілеадового, сина Махірового, сина Манасіїного, з родів Манасії, сина Йосипового, а оце ймення дочок його: Махла, Ноа, і Хоґла, і Мілка, і Тірца.
NUM|27|2|І стали вони перед Мойсеєм і перед священиком Елеазаром та перед начальниками, і всією громадою при вході скинії заповіту, говорячи:
NUM|27|3|Наш батько помер у пустині, і він не був серед громади змовників на Господа в Кореєвій громаді, бо він помер за свій гріх, а синів він не мав.
NUM|27|4|Чому ймення нашого батька буде відняте з-посеред його роду, що немає в нього сина? Дай же нам володіння серед братів нашого батька!
NUM|27|5|І приніс Мойсей їхню справу перед Господнє лице.
NUM|27|6|І сказав Господь до Мойсея, говорячи:
NUM|27|7|Целофхадові дочки слушно говорять. Конче даси їм володіння спадкове серед братів їхнього батька, і зробиш, щоб перейшла їм спадщина їхнього батька.
NUM|27|8|А до Ізраїлевих синів будеш промовляти, говорячи: Коли хто помре, а сина в нього нема, то зробите, щоб спадок його перейшов дочці його.
NUM|27|9|А якщо в нього немає дочки, то дасте спадщину його братам його.
NUM|27|10|А якщо в нього немає братів, то дасте спадок його братам батька його.
NUM|27|11|А якщо в його батька немає братів, то дасте спадщину його родичеві, близькому йому з його роду, і він посяде його. А це стане для Ізраїлевих синів на правну постанову, як Господь наказав був Мойсеєві.
NUM|27|12|І сказав Господь до Мойсея: Вийди на цю гору Аварім, і побач той Край, що Я дав Ізраїлевим синам.
NUM|27|13|І побачиш його, і будеш прилучений до своєї рідні і ти, як був прилучений твій брат Аарон,
NUM|27|14|бо ви були неслухняні наказам Моїм у пустині Цін при сварці громади, щоб явилася святість Моя через воду на їхніх очах. Це вода Меріви Кадеської в пустині Цін.
NUM|27|15|І промовив Господь до Мойсея, говорячи:
NUM|27|16|Нехай призначить Господь, Бог духів і кожного тіла, чоловіка над громадою,
NUM|27|17|що вийде перед ними, і що ввійде перед ними, і що випровадить їх, і що впровадить їх, і не буде Господня громада, як отара, що не має пастуха.
NUM|27|18|І сказав Господь до Мойсея: Візьми собі Ісуса, Навинового сина, мужа, що в ньому Дух, і покладеш свою руку на нього.
NUM|27|19|І поставиш його перед священиком Елеазаром та перед усією громадою, і накажеш йому на їхніх очах.
NUM|27|20|І даси на нього з влади своєї, щоб чула вся громада Ізраїлевих синів.
NUM|27|21|І стане він перед священиком Елеазаром, і він запитає для нього вироку уріму перед Господнім лицем. І за наказом його вийдуть, і за наказом його ввійдуть він та всі Ізраїлеві сини з ним і вся громада.
NUM|27|22|І зробив Мойсей, як Господь наказав був йому. І взяв він Ісуса, і поставив його перед Елеазаром та перед усією громадою.
NUM|27|23|І поклав він руки свої на нього, і заповів йому, як Господь промовляв через Мойсея.
NUM|28|1|І Господь промовляв до Мойсея, говорячи:
NUM|28|2|Накажи Ізраїлевим синам, і скажи їм: Ви будете пильнувати жертву Мою, хліб Мій для огняних Моїх жертов, пахощі любі Мої, щоб приносити Мені означеного часу.
NUM|28|3|І скажи їм: Оце огняна жертва, що принесете Господеві: безвадні однорічні ягнята, двоє на день, цілопалення завжди.
NUM|28|4|Одне ягня принесеш уранці, а ягня друге принесеш надвечір.
NUM|28|5|І десяту частину ефи пшеничної муки на хлібну жертву, мішану в товченій оливі чверть гіна.
NUM|28|6|Це стале цілопалення, принесене на Сінайській горі на пахощі любі, огняна жертва для Господа.
NUM|28|7|А лита жертва його чверть гіна для одного ягняти. У святині принесеш литу жертву вина для Господа.
NUM|28|8|А друге ягня принесеш надвечір, принесеш як хлібну жертву ранку й як жертву литу його, це огняна жертва, любі пахощі для Господа.
NUM|28|9|А суботнього дня двоє однорічних безвадних ягнят, і дві десяті пшеничної муки, жертва хлібна, мішана в оливі, і жертва лита його.
NUM|28|10|Це суботнє цілопалення щосуботи його, окрім цілопалення сталого та його литої жертви.
NUM|28|11|А першого дня ваших місяців принесете цілопалення для Господа: бички, молоде з великої худоби два, і одного барана, однорічні ягнята сім безвадних,
NUM|28|12|і три десяті ефи пшеничної муки, жертву хлібну, мішану в оливі, для одного бичка, і дві десяті пшеничної муки, жертву хлібну, мішану в оливі, для одного барана,
NUM|28|13|і по десятій частині ефи пшеничної муки, жертву хлібну, мішану в оливі, для одного ягняти. Це цілопалення, пахощі любі, огняна жертва для Господа.
NUM|28|14|А їхні литі жертви: пів гіна вина буде для бика, а третина гіна для барана, а четвертина гіна для ягняти. Це новомісячне цілопалення кожного молодика, для всіх молодиків року.
NUM|28|15|І буде принесений один козел на жертву за гріх для Господа, крім сталого цілопалення, і лита жертва його.
NUM|28|16|А першого місяця, чотирнадцятого дня місяця Пасха для Господа.
NUM|28|17|А п'ятнадцятого дня того місяця свято, сім день опрісноки їсти.
NUM|28|18|Першого дня святі збори, жодного робочого зайняття не будете робити.
NUM|28|19|І принесете огняну жертву, цілопалення для Господа: бички, молоде з великої худоби два, і одного барана, і сім однорічних ягнят, безвадні вони будуть у вас.
NUM|28|20|А їхня хлібна жертва пшенична мука, мішана в оливі, принесете три десяті ефи для бичка й дві десяті для барана.
NUM|28|21|По десятій частині ефи принесеш для одного ягняти, так для семи ягнят.
NUM|28|22|І одного козла жертви за гріх на очищення вас,
NUM|28|23|окрім цілопалення ранку, що належить до сталого цілопалення, принесете оце.
NUM|28|24|Як оце, будете приносити щоденно сім день хліб огняної жертви, любі пахощі для Господа; окрім сталого цілопалення буде це принесене, і лита жертва його.
NUM|28|25|А сьомого дня будуть для вас святі збори, жодного робочого зайняття не будете робити.
NUM|28|26|А дня первоплодів, коли приносите нову хлібну жертву для Господа в ваших тижнях, будуть для вас святі збори, жодного робочого зайняття не будете робити.
NUM|28|27|І принесете цілопалення на любі пахощі для Господа: бички, молоде з великої худоби два, барана одного, сім ягнят однорічних.
NUM|28|28|А їхня хлібна жертва: пшенична мука, мішана в оливі, три десяті ефи для одного бичка, дві десяті для одного барана,
NUM|28|29|по десятій частині ефи для одного ягняти, так для семи ягнят.
NUM|28|30|Козел один, на очищення вас,
NUM|28|31|окрім сталого цілопалення та хлібної його жертви це принесете, вони будуть безвадні у вас, і їхні литі жертви.
NUM|29|1|А сьомого місяця, першого дня місяця святі збори будуть для вас, жодного робочого зайняття не будете робити, це буде для вас день сурмлення.
NUM|29|2|І спорядите цілопалення на пахощі любі для Господа: бичка, молоде з великої худоби, одного, барана одного, однорічні ягнята, семеро безвадних.
NUM|29|3|А їхня хлібна жертва: пшенична мука, мішана в оливі, три десяті ефи для бичка, дві десяті для барана,
NUM|29|4|і одна десята для одного ягняти, так для семи ягнят,
NUM|29|5|і один козел, жертва за гріх, на очищення вас,
NUM|29|6|окрім новомісячного цілопалення й хлібної його жертви та цілопалення сталого, і хлібної його жертви та їхніх литих жертов за їхньою постановою, на любі пахощі, огняна жертва для Господа.
NUM|29|7|А десятого дня того сьомого місяця будуть для вас святі збори, і будете впокоряти свої душі, жодного зайняття не будете робити.
NUM|29|8|І принесете цілопалення для Господа, любі пахощі: бичка, молоде з великої худоби, одного, барана одного, однорічних ягнят семеро, безвадні будуть у вас.
NUM|29|9|А їхня хлібна жертва: пшенична мука, мішана в оливі, три десяті ефи для бичка, дві десяті для одного барана,
NUM|29|10|по десятій для одного ягняти, так для семи ягнят.
NUM|29|11|Козел один, жертва за гріх, окрім жертви за гріх очищення й сталого цілопалення, і його жертви хлібної та їхніх литих жертов.
NUM|29|12|А п'ятнадцятого дня сьомого місяця будуть для вас святі збори, жодного робочого заняття не будете робити, і будете святкувати сім день для Господа.
NUM|29|13|І принесете цілопалення, огняну жертву, пахощі любі для Господа: бички, молоде з великої худоби, тринадцятеро, барани два, однорічних ягнят чотирнадцятеро, безвадні будуть вони.
NUM|29|14|А хлібна їхня жертва: пшенична мука, мішана в оливі, три десяті ефи для кожного з тринадцяти бичків, дві десяті для одного барана, для двох баранів,
NUM|29|15|і по десятій для кожного з чотирнадцяти ягнят,
NUM|29|16|і один козел, жертва за гріх, окрім сталого цілопалення, його хлібної жертви та його жертви литої.
NUM|29|17|А другого дня: бички, молоде з великої худоби, дванадцятеро, барани два, однорічні ягнята чотирнадцятеро, безвадні.
NUM|29|18|А хлібна їхня жертва та їхні литі жертви для бичків, для баранів і для ягнят за числом їх, за постановою.
NUM|29|19|І козел один, жертва за гріх, окрім сталого цілопалення й хлібної його жертви та їхніх литих жертов.
NUM|29|20|А третього дня: бички одинадцятеро, барани два, однорічні ягнята чотирнадцятеро, безвадні.
NUM|29|21|А хлібна їхня жертва та їхні литі жертви для бичків, для баранів і для ягнят за числом їх, за постановою.
NUM|29|22|І козел жертви за гріх один, окрім сталого цілопалення й його хлібної жертви та його литої жертви.
NUM|29|23|А четвертого дня: бички десятеро, барани два, однорічні ягнята чотирнадцятеро, безвадні.
NUM|29|24|Хлібна їхня жертва та їхні литі жертви для бичків, для баранів і для ягнят за числом їх, за постановою.
NUM|29|25|І козел один, жертва за гріх, окрім сталого цілопалення їхньої хлібної жертви та їхньої литої жертви.
NUM|29|26|А п'ятого дня: бички дев'ятеро, барани два, однорічні ягнята чотирнадцятеро, безвадні.
NUM|29|27|А хлібна їхня жертва та їхні литі жертви для бичків, для баранів і для ягнят за числом їх, за постановою.
NUM|29|28|І козел жертви за гріх один, окрім сталого цілопалення та його хлібної жертви та його литої жертви.
NUM|29|29|А шостого дня: бички восьмеро, барани двоє, однорічні ягнята чотирнадцятеро, безвадні.
NUM|29|30|А хлібна їхня жертва та їхні литі жертви для бичків, для баранів і для ягнят за числом їх за постановою.
NUM|29|31|І козел жертви за гріх один, окрім сталого цілопалення його хлібної жертви та його литих жертов.
NUM|29|32|А сьомого дня: бички семеро, барани двоє, однорічні ягнята чотирнадцятеро, безвадні.
NUM|29|33|А хлібна їхня жертва та їхні литі жертви для бичків, для баранів і для ягнят за числом їх, за постановою.
NUM|29|34|І козел жертви за гріх один, окрім сталого цілопалення його хлібної жертви та його литої жертви.
NUM|29|35|А восьмого дня буде для вас віддання свята, жодного робочого зайняття не будете робити.
NUM|29|36|І принесете цілопалення, огняну жертву, пахощі любі для Господа: бичка одного, барана одного, однорічних ягнят семеро, безвадні.
NUM|29|37|Хлібна їхня жертва та їхні литі жертви для бичка, для барана й для ягнят за числом їх, за постановою.
NUM|29|38|І козел жертви за гріх один, окрім сталого цілопалення та його хлібної жертви та його литої жертви.
NUM|29|39|це принесете для Господа в ваші свята, окрім ваших обітниць та ваших дарів, для ваших цілопалень, і для ваших хлібних жертов, і для ваших литих жертов, і для ваших жертов мирних.
NUM|29|40|(30-1) І Мойсей сказав Ізраїлевим синам усе так, як Господь наказав Мойсеєві.
NUM|30|1|(30-2) І Промовляв Мойсей до голів племен Ізраїлевих синів, говорячи: Оце та річ, що Господь наказав:
NUM|30|2|(30-3) Коли хто складає обітницю для Господа або присягне присягу заректи зарока на душу свою, хай той не порушить свого слова, нехай зробить усе, як вийшло було з його уст.
NUM|30|3|(30-4) А жінка, коли складає обітницю для Господа, і зарече зарока в домі свого батька в своїй молодості,
NUM|30|4|(30-5) і почує її батько обітницю її та зарока, що зарекла на свою душу, та буде мовчати їй батько її, то будуть важні всі обітниці її, і буде важний кожен зарік її, що вона зарекла на душу свою.
NUM|30|5|(30-6) А якщо батько її заборонить їй того дня, коли був почув, усі обітниці її та зароки її, що зарекла на свою душу, то не будуть вони важні, а Господь пробачить їй, бо її батько заборонив їй.
NUM|30|6|(30-7) А якщо буде вона заміжня, а обітниці її на ній або мова уст її, що зарекла на душу свою,
NUM|30|7|(30-8) і почує її чоловік, і буде мовчати їй того дня, коли почує, то будуть важні обітниці її, і зароки її, що зарекла на свою душу, будуть важні.
NUM|30|8|(30-9) А якщо того дня, коли чоловік її почув, він заборонить їй і уневажнить обітниці її, що на ній, і мову уст її, що зарекла на свою душу, то Господь пробачить їй.
NUM|30|9|(30-10) А обітниця вдови та розведеної, усе, що зарекла на свою душу, буде важне на ній.
NUM|30|10|(30-11) А якщо вона обітувала в домі свого чоловіка, або зарекла зарока на свою душу присягою,
NUM|30|11|(30-12) а чоловік її чув та змовчав їй, не заборонив їй, то будуть важні всі обітниці її, і кожен зарік, що зарекла на свою душу, буде важний.
NUM|30|12|(30-13) А якщо справді уневажнить їх чоловік її того дня, коли він почує, то все, що вийшло з її уст для її обітниць та для зароків душі її, не буде важне, її чоловік уневажнив їх, і Господь простить їй.
NUM|30|13|(30-14) Кожна обітниця й кожна присяга зароку впокоряти свою душу, чоловік її зробить важною, або чоловік її уневажнить її.
NUM|30|14|(30-15) А якщо чоловік її, замовчуючи, буде мовчати їй з дня на день, то зробить важними всі її обітниці, або всі її зароки, що на ній; зробив їх важними, бо він мовчав їй того дня, коли був почув.
NUM|30|15|(30-16) А якщо справді уневажнить він їх по тому, як був почув, то понесе він гріх її.
NUM|30|16|(30-17) Оце постанови, що Господь наказав був Мойсеєві, у цій справі між чоловіком та його жінкою, між батьком та його дочкою в її молодості в домі батька свого.
NUM|31|1|І Господь промовляв до Мойсея, говорячи:
NUM|31|2|Пімсти мідіянітам за кривду Ізраїлевих синів, потім будеш прилучений до своєї рідні.
NUM|31|3|І промовив Мойсей до народу, говорячи: Озбройте з-поміж себе людей для війська, і будуть вони на мідіян, щоб дати Господню пімсту на мідіян.
NUM|31|4|По тисячі з племені зо всіх Ізраїлевих племен пошлете до війська.
NUM|31|5|І були призначені з Ізраїлевих тисяч тисяча з племені дванадцять тисяч узброєних для війська.
NUM|31|6|І послав їх Мойсей тисячу з кожного племени до їх війська, і Пінхаса, сина священика Елеазара, на війну, і святий посуд, і сурми для сурмлення в його руці.
NUM|31|7|І рушили війною на Мідіяна, як наказав був Господь Мойсеєві, і позабивали кожного чоловічої статі.
NUM|31|8|І крім тих забитих, позабивали мідіянських царів: Евія, і Рекема, і Цура, і Хура, і Реву, п'ять мідіянських царів, і Валаама, Беорового сина, забили мечем.
NUM|31|9|І полонили Ізраїлеві сини мідіянських жінок і їхніх дітей, і всю їхню худобу, і всі їхні стада та ввесь їх маєток пограбували.
NUM|31|10|А всі їхні міста по їхніх осадах та всі їхні оселі попалили огнем.
NUM|31|11|І позабирали вони все захоплене й усю здобич, людей та худобу.
NUM|31|12|І вони привели до Мойсея й до священика Елеазара та до громади Ізраїлевих синів полонених і здобич, і захоплене до табору, до моавських степів, що над приєрихонським Йорданом.
NUM|31|13|І вийшли Мойсей і священик Елеазар та всі начальники громади назустріч їм поза табір.
NUM|31|14|І розгнівався Мойсей на військових провідників, тисячників та сотників, що верталися з війська тієї війни.
NUM|31|15|І сказав до них Мойсей: Чи ви позоставили живими всіх жінок?
NUM|31|16|Тож вони були для Ізраїлевих синів за радою Валаама причиною на відступлення від Господа через Пеора! І була поразка в Господній громаді.
NUM|31|17|А тепер позабивайте кожного хлопця між дітьми, і кожну жінку, що познала чоловіка на мужеськім ложі, повбивайте.
NUM|31|18|А всіх молодих жінок, що не познали мужеського ложа, зоставте живими для себе.
NUM|31|19|А ви пробудьте поза табором сім день. Кожен, хто забив кого, і кожен, хто доторкався трупа, очистьтеся дня третього й дня сьомого ви та ваші бранці.
NUM|31|20|І ви очистите кожну одежу, і кожну шкуряну річ, і все зроблене з козиної вовни, і кожну дерев'яну річ.
NUM|31|21|І сказав священик Елеазар воїнам, що ходили на війну: Оце постанова закону, що Господь наказав був Мойсеєві:
NUM|31|22|Тільки золото й срібло, мідь, залізо, цину та олово,
NUM|31|23|кожну річ, що видержить в огні, перепровадите через огонь, і стане чиста, тільки перше очищальною водою очиститься; а все, що не видержує огню, перепровадите через воду.
NUM|31|24|І виперете одежу свою сьомого дня, і станете чисті, а потому ввійдете до табору.
NUM|31|25|І Господь промовляв до Мойсея, говорячи:
NUM|31|26|Перелічи здобич бранців між людьми й між худобою ти й священик Елеазар та голови батьківських домів громади.
NUM|31|27|І поділиш ту здобич пополовині між учасниками війни, що входять до війська, і між усією громадою.
NUM|31|28|І принесеш данину для Господа від військових, що входять до війська, одну душу від п'яти сотень від людини й від великої худоби, і від ослів, і від худоби дрібної.
NUM|31|29|З їхньої половини візьми, і даси священикові Елеазарові як Господнє приношення.
NUM|31|30|А з половини Ізраїлевих синів візьмеш одного вийнятого з п'ятидесяти з людини, з худоби великої, з ослів та з худоби дрібної, з кожної скотини, та й даси їх Левитам, що виконують сторожу Господньої скинії.
NUM|31|31|І зробив Мойсей та священик Елеазар, як Господь наказав був Мойсеєві.
NUM|31|32|І була здобич, позостале грабунку, що захопили були військові: дрібної худоби шістсот тисяч і сімдесят тисяч і п'ять тисяч.
NUM|31|33|А худоба велика сімдесят і дві тисячі.
NUM|31|34|І осли шістдесят і одна тисяча.
NUM|31|35|А душ людських із жінок, що не пізнали мужеського ложа, усіх душ тридцять і дві тисячі.
NUM|31|36|І була половина, частка тих, що входили до війська, число худоби дрібної триста тисяч і тридцять тисяч і сім тисяч і п'ять сотень.
NUM|31|37|І була данина для Господа з худоби дрібної, шість сотень сімдесят і п'ять.
NUM|31|38|А худоба велика: тридцять і шість тисяч, а їхня данина для Господа сімдесят і двоє.
NUM|31|39|А осли: тридцять тисяч і п'ять сотень, а їхня данина для Господа шістдесят і один.
NUM|31|40|А душ людських: шістнадцять тисяч, а їхня данина для Господа тридцять і дві душі.
NUM|31|41|І дав Мойсей данину Господнього приношення священикові Елеазарові, як Господь наказав був Мойсеєві.
NUM|31|42|І з половини Ізраїлевих синів, що Мойсей відділив, від людей, що вирушали на війну,
NUM|31|43|і була громадська половина з дрібної худоби триста тисяч і тридцять тисяч і сім тисяч і п'ять сотень.
NUM|31|44|А худоба велика тридцять і шість тисяч.
NUM|31|45|А осли тридцять тисяч і п'ять сотень.
NUM|31|46|А людських душ шістнадцять тисяч,
NUM|31|47|і взяв Мойсей з половини Ізраїлевих синів вийнятого одного з п'ятидесяти з людини та зо скотини, та й дав їх Левитам, що виконують сторожу Господньої скинії, як Господь наказав був Мойсеєві.
NUM|31|48|І прийшли до Мойсея старшини над тисячами війська, тисячники та сотники,
NUM|31|49|та й сказали Мойсеєві: Твої раби перелічили військових, що під нашою рукою, і нікого з нас не бракувало.
NUM|31|50|І ми принесли Господню жертву, кожен, хто знайшов що з золота, ланцюжок на ноги, і нараменник, перстень, сережки та нашийника на очищення наших душ перед Господнім лицем.
NUM|31|51|І взяв Мойсей та священик Елеазар від них те золото, кожну зроблену річ.
NUM|31|52|І було всього золота приношення, що принесли для Господа, шістнадцять тисяч сімсот і п'ятдесят шеклів від тисячників і від сотників.
NUM|31|53|Військові грабували кожен для себе.
NUM|31|54|І взяв Мойсей та священик Елеазар те золото від тисячників та сотників, і внесли його до скинії заповіту, пам'ятка для Ізраїлевих синів перед Господнім лицем.
NUM|32|1|А в Рувимових синів та в синів Ґадових були великі стада, дуже численні. І побачили вони край Язерський та край Ґілеадський, а ото це місце місце добре для худоби.
NUM|32|2|І прийшли Ґадові сини та сини Рувимові, та й сказали до Мойсея й до священика Елеазара та до громадських начальників, говорячи:
NUM|32|3|Аторот, і Дівон, і Язер, і Німра, і Хешбон, і Ел'але і Севам, і Нево, і Беон,
NUM|32|4|та земля, що Господь побив був перед Ізраїлевою громадою, вона земля добра для худоби, а в твоїх рабів є худоба.
NUM|32|5|І сказали вони: Якщо ми знайшли ласку в очах твоїх, то нехай дано буде ту землю твоїм рабам на володіння. Не перепроваджуй нас через Йордан!
NUM|32|6|І сказав Мойсей до Ґадових синів та до синів Рувимових: Чи брати ваші підуть на війну, а ви будете тут сидіти?
NUM|32|7|І для чого ви стримуєте серце Ізраїлевих синів від переходу до того Краю, що дав їм Господь?
NUM|32|8|Так зробили були ваші батьки, коли я посилав їх із Кадеш-Барнеа побачити той Край.
NUM|32|9|І ввійшли вони в Ешкольську долину, і побачили були той Край, і стримали серце Ізраїлевих синів, щоб не входити до того Краю, що дав їм Господь.
NUM|32|10|І запалився Господній гнів того дня, і присягнув Він, говорячи:
NUM|32|11|Поправді кажу, не побачать ці люди, що виходять з Єгипту, від віку двадцяти літ і вище, тієї землі, що Я присягнув був Авраамові, Ісакові та Якову, бо вони не виконували наказів Моїх,
NUM|32|12|окрім Калева, Єфуннеєвого сина, кеніззеянина, та Ісуса, сина Навинового, бо вони виконували накази за Господом.
NUM|32|13|І запалився був гнів Господній на Ізраїля, і Він зробив, що вони ходили по пустині сорок літ, аж поки не скінчилося все те покоління, що робило зло в Господніх очах.
NUM|32|14|А оце стали ви замість ваших батьків, як нащадки грішних людей, щоб збільшити ще палючий гнів Господній на Ізраїля.
NUM|32|15|Бо як ви відвернетесь від Нього, то Він ще далі триматиме його в пустині, і ви спричините згубу всьому цьому народові.
NUM|32|16|А вони підійшли до нього та й сказали: Ми побудуємо тут кошари для нашої худоби та міста для наших дітей,
NUM|32|17|а ми самі узброїмося, готові до бою перед Ізраїлевими синами, аж поки не введемо їх до їхнього місця. А діти наші осядуть по твердинних містах, охороняючи себе перед мешканцями цієї землі.
NUM|32|18|Ми не вернемось до наших домів, аж поки Ізраїлеві сини не заволодіють кожен спадком своїм.
NUM|32|19|Бо ми не будемо володіти з ними по той бік Йордану й далі, бо прийшла нам наша спадщина з цього боку Йордану на схід.
NUM|32|20|І сказав їм Мойсей: Якщо ви зробите цю річ, якщо ви узброїтесь на війну перед Господнім лицем,
NUM|32|21|і перейде кожен ваш узброєний Йордан перед Господнім лицем, аж поки Він не вижене ворогів Своїх перед Собою,
NUM|32|22|то буде здобутий той Край перед Господнім лицем, і ви потому вернетеся, і будете невинні перед Господом та перед Ізраїлем. І буде вам цей Край на володіння перед Господнім лицем.
NUM|32|23|А якщо не зробите так, то ви згрішили Господеві, і знайте, що ваш гріх знайде вас!
NUM|32|24|Побудуйте собі міста для ваших дітей, та кошари для ваших отар. А що вийшло з ваших уст, те зробіть.
NUM|32|25|І сказали Ґадові сини та сини Рувимові до Мойсея, говорячи: Раби твої зроблять, як пан наш приказує.
NUM|32|26|Діти наші, жінки наші, стадо наше та вся наша худоба будуть там, у ґілеадських містах.
NUM|32|27|А раби твої перейдуть, кожен військовий озброєний, перед Господнім лицем на війну, як пан наш наказує.
NUM|32|28|І Мойсей наказав про них священикові Елеазарові й Ісусові, синові Навиновому, та головам батьківських домів племен Ізраїлевих синів.
NUM|32|29|І сказав Мойсей до них: Якщо Ґадові сини та сини Рувимові перейдуть із вами Йордан, кожен озброєний на війну перед лицем Господнім, і буде здобутий Край перед вами, то дасте їм ґілеадський край на володіння.
NUM|32|30|А якщо вони не перейдуть з вами озброєні, то отримають володіння серед вас в ханаанському Краї.
NUM|32|31|І відповіли Ґадові сини та сини Рувимові, говорячи: Що говорив Господь до твоїх рабів, так зробимо.
NUM|32|32|Ми перейдемо озброєні перед Господнім лицем до ханаанського Краю, а з нами буде наше володіння по цей бік Йордану.
NUM|32|33|І Мойсей дав їм, Ґадовим синам і синам Рувимовим та половині племені Манасії, Йосипового сина, царство Сігона, царя аморейського, і царство Оґа, царя башанського, той Край по містах його, у границях міст того Краю навколо.
NUM|32|34|І збудували Ґадові сини Дівон, і Атарот, і Ароер,
NUM|32|35|і Атарот Шофан, і Язер, і Йоґбегу,
NUM|32|36|і Бет-Німру, і Бет-Гаран, твердинні міста та кошари для отари.
NUM|32|37|У Рувимові сини збудували: Хешбон, і Ел'але, і Кір'ятаїм,
NUM|32|38|і Нево, і Баал-Меон, зміненоіменні, і Сивму, і назвали йменнями міста, що вони збудували.
NUM|32|39|І пішли сини Махіра, сина Манасії, до Ґілеаду, та й здобули його, і позбавили спадщини амореянина, що в ньому.
NUM|32|40|І дав Мойсей Ґілеад Махірові, синові Манасії, і той осів у ньому.
NUM|32|41|А Яір, син Манасіїн, пішов і здобув їхні села, та й назвав їх: Яірові села.
NUM|32|42|А Новах пішов та й здобув Кенат та залежні від нього міста, і назвав його своїм ім'ям: Новах.
NUM|33|1|Оце походи Ізраїлевих синів, що вийшли з єгипетського краю за своїми військовими відділами під рукою Мойсея та Аарона.
NUM|33|2|А Мойсей написав їхні виходи з їхніми походами за Господнім наказом, і оце їхні походи за їхніми виходами.
NUM|33|3|І рушили вони з Рамесесу першого місяця, п'ятнадцятого дня першого місяця, другого дня по Пасці вийшли Ізраїлеві сини сильною рукою на очах усього Єгипту.
NUM|33|4|А Єгипет ховав, кого побив Господь серед них, кожного перворідного, а над їхніми богами зробив Господь суди.
NUM|33|5|І рушили Ізраїлеві сини з Рамесесу, і таборували в Суккоті.
NUM|33|6|І рушили з Суккоту й таборували в Етамі, що на краю пустині.
NUM|33|7|І рушили з Етаму, а вернулися до Пі-Хіроту, що перед Баал-Цефоном, і таборували перед Міґдолом.
NUM|33|8|І рушили з-перед Хіроту, і перейшли серед моря до пустині, і йшли триденною дорогою в Етамській пустині, і таборували в Марі.
NUM|33|9|І рушили з Мари й увійшли до Еліму, а в Елімі дванадцять джерел води та сімдесят пальм, і таборували там.
NUM|33|10|І рушили з Еліму й таборували над Червоним морем.
NUM|33|11|І рушили з-над Червоного моря й таборували в пустині Сін.
NUM|33|12|І рушили з пустині Сін і таборували в Дофці.
NUM|33|13|І рушили з Дофки й таборували в Алуші.
NUM|33|14|І рушили з Алушу й таборували в Ріфідімі, і не було там води на пиття для народу.
NUM|33|15|І рушили з Ріфідіму й таборували в пустині Сінай.
NUM|33|16|І рушили з пустині Сінай і таборували в Ківрот-Гаттааві.
NUM|33|17|І рушили з Ківрот-Гаттаави й таборували в Хацероті.
NUM|33|18|І рушили з Хацероту й таборували в Рітмі.
NUM|33|19|І рушили з Рітми й таборували в Ріммоні Переца.
NUM|33|20|І рушили з Ріммону Переца й таборували в Лівні.
NUM|33|21|І рушили з Лівни й таборували в Ріссі.
NUM|33|22|І рушили з Рісси й таборували в Кегелаті.
NUM|33|23|І рушили з Кегелати й таборували на горі Шефер.
NUM|33|24|І рушили з гори Шефер і таборували в Хараді.
NUM|33|25|І рушили з Харади й таборували в Макгелоті.
NUM|33|26|І рушили з Макгелоту й таборували в Тахаті.
NUM|33|27|І рушили з Тахату й таборували в Тераху.
NUM|33|28|І рушили з Тераху й таборували в Мітці.
NUM|33|29|І рушили з Мітки й таборували в Хашмоні.
NUM|33|30|І рушили з Хашмони й таборували в Мосероті.
NUM|33|31|І рушили з Мосероту й таборували в Бене-Яакані.
NUM|33|32|І рушили з Бене-Яакану й таборували в Хорі Ґідґаду.
NUM|33|33|І рушили з Хору Ґідґаду й таборували в Йотваті.
NUM|33|34|І рушили з Йотвати й таборували в Авроні.
NUM|33|35|І рушили з Аврони й таборували в Ецйон-Ґевері.
NUM|33|36|І рушили з Ецйон-Ґеверу й таборували в пустині Цін, це Кадеш.
NUM|33|37|І рушили з Кадешу й таборували на Гор-горі, на краю едомської землі.
NUM|33|38|І зійшов священик Аарон на Гор-гору з Господнього наказу, та й помер там сорокового року виходу Ізраїлевих синів з єгипетського краю, п'ятого місяця, першого дня місяця.
NUM|33|39|А Аарон був віку ста й двадцяти й трьох літ, коли помер він на Гор-горі.
NUM|33|40|І почув ханаанеянин, цар Араду, а він сидів на півдні в Краї ханаанськім, що йдуть Ізраїлеві сини.
NUM|33|41|І рушили від Гор-гори й таборували в Цалмоні.
NUM|33|42|І рушили з Цалмони й таборували в Пуноні.
NUM|33|43|І рушили з Пунону й таборували в Овоті.
NUM|33|44|І рушили з Овоту й таборували в Ійє-Гааварімі, на моавській границі.
NUM|33|45|І рушили з Ійїму й таборували в Дівоні Ґаду.
NUM|33|46|І рушили з Дівону Ґаду й таборували в Алмон-Дівлатаймі.
NUM|33|47|І рушили з Алмон-Дівлатайми й таборували в горах Аварім перед Нево.
NUM|33|48|І рушили з гір Аварім, і таборували в моавських степах.
NUM|33|49|І таборували вони над Йорданом від Бет-Єшмоту аж до Авел-Шіттіму в моавських степах.
NUM|33|50|І Господь промовляв до Мойсея в моавських степах над приєрихонським Йорданом, говорячи:
NUM|33|51|Промовляй до Ізраїлевих синів та й скажеш до них: Коли ви перейдете Йордан до ханаанського Краю,
NUM|33|52|то проженете всіх мешканців того Краю перед собою, і понищите всі їхні зображення, і всіх литих ідолів їхніх понищите, і всі їхні висоти поруйнуєте.
NUM|33|53|І ви заволодієте тим Краєм, і осядете в ньому, бо Я дав вам той Край на власність.
NUM|33|54|І ви заволодієте тим Краєм жеребком за вашими родами: численному збільшите власність його, а малому зменшите власність його, де вийде йому жеребок, туди йому буде, за племенами ваших батьків будете володіти собі.
NUM|33|55|А якщо ви не виженете мешканців того Краю від себе, то будуть ті, кого позоставите з них, колючками в ваших очах та тернями в ваших боках. І будуть вас утискати на тій землі, що на ній ви сидітимете.
NUM|33|56|І станеться, як Я думав був учинити їм, учиню те вам.
NUM|34|1|І Господь промовляв до Мойсея, говорячи:
NUM|34|2|Накажи Ізраїлевим синам та й скажи їм: Коли ви ввійдете до ханаанського Краю, це буде той Край, що припаде вам у спадщині, ханаанський Край по границях його.
NUM|34|3|І буде вам південна сторона від пустині Цін при Едомі, і буде вам південна границя від кінця Солоного моря на схід.
NUM|34|4|І скерується вам та границя з полудня до Маале-Акраббіму, і перейде до Ціну, і будуть виходи її з полудня до Кадеш-Барнеа. І вийде вона до Хацар-Аддару й перейде до Ацмону.
NUM|34|5|І скерується границя з Ацмону до єгипетського потоку, і будуть її виходи до моря.
NUM|34|6|А границя західня, буде для вас море Велике, це буде для вас західня границя.
NUM|34|7|А оце буде для вас північна границя: від Великого моря визначите собі за границю Гор-гору.
NUM|34|8|Від Гор-гори визначите в напрямі до Гамату, і будуть виходи границі до Цедаду.
NUM|34|9|І вийде границя до Зіфрону, і будуть її виходи до Гацар-Енану. Це буде вам північна границя.
NUM|34|10|І визначите собі за границю на схід від Гацар-Енану до Шефаму.
NUM|34|11|І зійде границя від Шефаму до Рівли, на схід Аіну. І зійде границя, і дійде на беріг Кінеретського моря на схід.
NUM|34|12|І зійде границя до Йордану, і будуть її виходи море Солоне. Це буде для вас Край по його границях навколо.
NUM|34|13|І Мойсей наказав Ізраїлевим синам, говорячи: Оце та земля, що ви поділите собі її жеребком, що Господь наказав дати дев'яти племенам і половині племені.
NUM|34|14|Бо взяли плем'я Рувимових синів за домами батьків своїх, і плем'я Ґадових синів за домами батьків своїх, і половина племени Манасіїного взяли спадщину свою,
NUM|34|15|два племені й половина племени взяли вже свою спадщину з того боку приєрихонського Йордану на схід та на південь.
NUM|34|16|І Господь промовляв до Мойсея, говорячи:
NUM|34|17|Оце імена тих мужів, що поділять для вас той Край на спадок: священик Елеазар та Ісус, син Навинів,
NUM|34|18|та візьмете по одному князеві з племени, щоб поділити той Край на власність.
NUM|34|19|А оце ймення тих мужів: для Юдиного племени Калев, син Єфуннеїв;
NUM|34|20|а для племени Симеонових синів Шемуїл, син Аммігудів;
NUM|34|21|а для племени Веніяминового Елідад, син Кіслонів;
NUM|34|22|для племени Данових синів князь Буккі, син Йоґліїв;
NUM|34|23|для Йосипових синів, для племени синів Манасіїних князь Ханніїл, син Ефодів;
NUM|34|24|а для племени Єфремових синів князь Кемуїл, син Шіфтанів;
NUM|34|25|а для племени Завулонових синів князь Еліцафан, син Парнахів;
NUM|34|26|а для племени Іссахарових синів князь Палтіїл, син Аззана;
NUM|34|27|а для племени Асирових синів князь Ахігуд, син Шеломіїв;
NUM|34|28|а для племени синів Нефталимових князь Педаїл, син Аммігудів.
NUM|34|29|Оце ті, кому наказав Господь поділити ханаанський Край на спадщину для Ізраїлевих синів.
NUM|35|1|І Господь промовляв до Мойсея на моавських степах над приєрихонським Йорданом, говорячи:
NUM|35|2|Накажи Ізраїлевим синам, і нехай вони дадуть Левитам зо спадку свого володіння міста на сидіння; і пасовисько для міст навколо них дасте ви Левитам.
NUM|35|3|І будуть ті міста їм на сидіння, а їхні пасовиська будуть для їхньої скотини, і для їхньої худоби та для всієї їхньої звірини.
NUM|35|4|А пасовиська тих міст, що дасте Левитам, будуть тягнутись від міської стіни й назовні тисяча локтів навколо.
NUM|35|5|І відміряєте поза містом на східню сторону дві тисячі ліктів, і на південну сторону дві тисячі ліктів, і на західню сторону дві тисячі ліктів, і на північну сторону дві тисячі ліктів, а місто усередині. Це будуть для вас міські пасовиська.
NUM|35|6|А з міст, що дасте Левитам, буде шість міст на сховища, що дасте, щоб утікати туди убійникові. А окрім них дасте сорок і два міста.
NUM|35|7|Усі ті міста, що дасте Левитам, сорок і вісім їхніх міст та їхні пасовиська.
NUM|35|8|А ті міста, що дасте з володіння Ізраїлевих синів, від більшого дасте більше, а від меншого менше, кожен за спадком своїм, яким володітиме, дасть із своїх міст Левитам.
NUM|35|9|І Господь промовляв до Мойсея, говорячи:
NUM|35|10|Промовляй до Ізраїлевих синів та й скажи їм: Коли ви перейдете Йордан до ханаанського Краю,
NUM|35|11|то виберіть собі міста, вони будуть на сховища для вас, і втече туди убійник, що заб'є душу невмисне.
NUM|35|12|І будуть для вас ті міста на сховища перед месником, і не помре убійник, поки не стане на суд перед громадою.
NUM|35|13|А ті міста, що дасте, шість міст на сховища буде для вас.
NUM|35|14|Три місті дасте по той бік Йордану, а три місті дасте в ханаанському Краї, вони будуть міста на сховища.
NUM|35|15|Ці шість міст будуть на сховища для Ізраїлевих синів, і для приходька та для осілого серед них, щоб утік туди кожен, хто заб'є кого невмисне.
NUM|35|16|А коли б хто вдарив кого залізним знаряддям, а той помер, він убійник, буде конче забитий той убійник.
NUM|35|17|А якщо вдарив його каменем, що був у руці, що від нього можна померти, і той помер, він убійник, буде конче забитий той убійник.
NUM|35|18|Або вдарив його дерев'яним знаряддям, що було в руці, що від нього можна померти, і той помер, він убійник, буде конче забитий той убійник.
NUM|35|19|Месник за кров він заб'є убійника; як спіткає його, він заб'є його.
NUM|35|20|А якщо пхне його з ненависти, або кине на нього чим навмисне, а той помре,
NUM|35|21|або з ворогування вдарив його своєю рукою, а той помер, буде конче забитий той, хто вдарив, він убійник; месник за кров заб'є убійника, як спіткає його.
NUM|35|22|А як хто випадково, без ненависти пхнув кого або кинув на нього невмисне якимбудь знаряддям,
NUM|35|23|або якимбудь каменем, що від нього можна померти, кинув на нього не бачачи, і той помер, а він не був ворог йому й не шукав йому зла,
NUM|35|24|то розсудить громада між убійником та між месником за кров за цими постановами.
NUM|35|25|І громада визволить убійника з руки месника за кров, і громада верне його до міста сховища його, що втік був туди. І осяде він у ньому аж до смерти найвищого священика, помазаного святою оливою.
NUM|35|26|А якщо убійник, виходячи, вийде з границі міста сховища його, куди втік був,
NUM|35|27|і знайде його месник за кров поза границями міста сховища його, і замордує месник за кров убійника, нема йому вини крови!
NUM|35|28|Бо він повинен сидіти в місті сховища свого аж до смерти найвищого священика. А по смерті найвищого священика вернеться убійник до землі володіння свого.
NUM|35|29|І буде це для вас на правну постанову для ваших поколінь по всіх ваших оселях.
NUM|35|30|Коли хто заб'є кого, то месник за словами свідків заб'є убійника. А одного свідка не досить проти кого, щоб осудити на смерть.
NUM|35|31|І не візьмете окупу для душі убійника, що він повинен умерти, бо буде він конче забитий.
NUM|35|32|І не візьмете окупу від змушеного втікати до міста сховища його, щоб вернувся сидіти в Краю до смерти священика.
NUM|35|33|І не збезчестите того Краю, що ви в ньому, бо та кров вона безчестить Край, а Краєві не прощається за кров, що пролита в ньому, як тільки кров'ю того, хто її пролив.
NUM|35|34|І не занечистиш того Краю, що ви сидите в ньому, що Я пробуваю серед нього. Бо Я Господь, що пробуваю посеред синів Ізраїлевих!
NUM|36|1|І поприходили голови батьківських домів родів синів Ґілеада, сина Махіра, сина Манасіїного з родів Йосипових синів, і промовили перед Мойсеєм та перед князями, головами батьківських домів Ізраїлевих синів,
NUM|36|2|і сказали: Господь наказав моєму панові дати жеребком цей Край Ізраїлевим синам, і пан мій отримав Господнього наказа дати спадок нашого брата Целофхада його дочкам.
NUM|36|3|І якщо вони будуть за жінок кому з синів інших племен Ізраїлевих синів, то буде віднята їхня спадщина зо спадку наших батьків, і буде додане над спадок тому племені, що вони стануть їм за жінок, а з жеребка нашого спадку буде відняте.
NUM|36|4|А якщо Ізраїлевим синам буде ювілей, то буде їхня спадщина додана до спадку племени, що стануть їм за жінок, і їхня спадщина буде віднята від спадку племени наших батьків.
NUM|36|5|І наказав Мойсей Ізраїлевим синам за Господнім наказом, говорячи: Слушно говорить плем'я Йосипових синів.
NUM|36|6|Оце та річ, що Господь заповів про Целофхадових дочок, говорячи: Вони стануть за жінок тим, хто їм подобається, тільки родові племени їхнього батька вони стануть за жінок.
NUM|36|7|І не буде переходити спадщина Ізраїлевих синів від племени до племени, бо кожен із Ізраїлевих синів буде держатися спадщини племени своїх батьків.
NUM|36|8|А кожна дочка, що посяде спадщину від племени Ізраїлевих синів, стане за жінку одному з роду племени батька свого, щоб Ізраїлеві сини володіли кожен спадком батьків своїх.
NUM|36|9|І не буде переходити спадок від племени до іншого племени, бо кожен із племен Ізраїлевих синів буде держатися спадку свого.
NUM|36|10|Як Господь наказав був Мойсеєві, так учинили Целофхадові дочки.
NUM|36|11|І стали Целофхадові дочки: Махла, Тірца, і Хоґла, і Мілка, і Ноа за жінок для синів дядьків своїх.
NUM|36|12|Тим, що з родів синів Манасіїних, сина Йосипового, стали вони за жінок, а їхня спадщина залишилася за племенем роду їхнього батька.
NUM|36|13|Оце заповіді та постанови, що Господь наказав був через Мойсея Ізраїлевим синам у моавських степах над приєрихонським Йорданом.
