PHIL|1|1|Paul and Timothy, servants of Christ Jesus, To all the saints in Christ Jesus at Philippi, together with the overseers and deacons:
PHIL|1|2|Grace and peace to you from God our Father and the Lord Jesus Christ.
PHIL|1|3|I thank my God every time I remember you.
PHIL|1|4|In all my prayers for all of you, I always pray with joy
PHIL|1|5|because of your partnership in the gospel from the first day until now,
PHIL|1|6|being confident of this, that he who began a good work in you will carry it on to completion until the day of Christ Jesus.
PHIL|1|7|It is right for me to feel this way about all of you, since I have you in my heart; for whether I am in chains or defending and confirming the gospel, all of you share in God's grace with me.
PHIL|1|8|God can testify how I long for all of you with the affection of Christ Jesus.
PHIL|1|9|And this is my prayer: that your love may abound more and more in knowledge and depth of insight,
PHIL|1|10|so that you may be able to discern what is best and may be pure and blameless until the day of Christ,
PHIL|1|11|filled with the fruit of righteousness that comes through Jesus Christ--to the glory and praise of God.
PHIL|1|12|Now I want you to know, brothers, that what has happened to me has really served to advance the gospel.
PHIL|1|13|As a result, it has become clear throughout the whole palace guard and to everyone else that I am in chains for Christ.
PHIL|1|14|Because of my chains, most of the brothers in the Lord have been encouraged to speak the word of God more courageously and fearlessly.
PHIL|1|15|It is true that some preach Christ out of envy and rivalry, but others out of goodwill.
PHIL|1|16|The latter do so in love, knowing that I am put here for the defense of the gospel.
PHIL|1|17|The former preach Christ out of selfish ambition, not sincerely, supposing that they can stir up trouble for me while I am in chains.
PHIL|1|18|But what does it matter? The important thing is that in every way, whether from false motives or true, Christ is preached. And because of this I rejoice.
PHIL|1|19|Yes, and I will continue to rejoice, for I know that through your prayers and the help given by the Spirit of Jesus Christ, what has happened to me will turn out for my deliverance.
PHIL|1|20|I eagerly expect and hope that I will in no way be ashamed, but will have sufficient courage so that now as always Christ will be exalted in my body, whether by life or by death.
PHIL|1|21|For to me, to live is Christ and to die is gain.
PHIL|1|22|If I am to go on living in the body, this will mean fruitful labor for me. Yet what shall I choose? I do not know!
PHIL|1|23|I am torn between the two: I desire to depart and be with Christ, which is better by far;
PHIL|1|24|but it is more necessary for you that I remain in the body.
PHIL|1|25|Convinced of this, I know that I will remain, and I will continue with all of you for your progress and joy in the faith,
PHIL|1|26|so that through my being with you again your joy in Christ Jesus will overflow on account of me.
PHIL|1|27|Whatever happens, conduct yourselves in a manner worthy of the gospel of Christ. Then, whether I come and see you or only hear about you in my absence, I will know that you stand firm in one spirit, contending as one man for the faith of the gospel
PHIL|1|28|without being frightened in any way by those who oppose you. This is a sign to them that they will be destroyed, but that you will be saved--and that by God.
PHIL|1|29|For it has been granted to you on behalf of Christ not only to believe on him, but also to suffer for him,
PHIL|1|30|since you are going through the same struggle you saw I had, and now hear that I still have.
PHIL|2|1|If you have any encouragement from being united with Christ, if any comfort from his love, if any fellowship with the Spirit, if any tenderness and compassion,
PHIL|2|2|then make my joy complete by being like-minded, having the same love, being one in spirit and purpose.
PHIL|2|3|Do nothing out of selfish ambition or vain conceit, but in humility consider others better than yourselves.
PHIL|2|4|Each of you should look not only to your own interests, but also to the interests of others.
PHIL|2|5|Your attitude should be the same as that of Christ Jesus:
PHIL|2|6|Who, being in very nature God, did not consider equality with God something to be grasped,
PHIL|2|7|but made himself nothing, taking the very nature of a servant, being made in human likeness.
PHIL|2|8|And being found in appearance as a man, he humbled himself and became obedient to death--even death on a cross!
PHIL|2|9|Therefore God exalted him to the highest place and gave him the name that is above every name,
PHIL|2|10|that at the name of Jesus every knee should bow, in heaven and on earth and under the earth,
PHIL|2|11|and every tongue confess that Jesus Christ is Lord, to the glory of God the Father.
PHIL|2|12|Therefore, my dear friends, as you have always obeyed--not only in my presence, but now much more in my absence--continue to work out your salvation with fear and trembling,
PHIL|2|13|for it is God who works in you to will and to act according to his good purpose.
PHIL|2|14|Do everything without complaining or arguing,
PHIL|2|15|so that you may become blameless and pure, children of God without fault in a crooked and depraved generation, in which you shine like stars in the universe
PHIL|2|16|as you hold out the word of life--in order that I may boast on the day of Christ that I did not run or labor for nothing.
PHIL|2|17|But even if I am being poured out like a drink offering on the sacrifice and service coming from your faith, I am glad and rejoice with all of you.
PHIL|2|18|So you too should be glad and rejoice with me.
PHIL|2|19|I hope in the Lord Jesus to send Timothy to you soon, that I also may be cheered when I receive news about you.
PHIL|2|20|I have no one else like him, who takes a genuine interest in your welfare.
PHIL|2|21|For everyone looks out for his own interests, not those of Jesus Christ.
PHIL|2|22|But you know that Timothy has proved himself, because as a son with his father he has served with me in the work of the gospel.
PHIL|2|23|I hope, therefore, to send him as soon as I see how things go with me.
PHIL|2|24|And I am confident in the Lord that I myself will come soon.
PHIL|2|25|But I think it is necessary to send back to you Epaphroditus, my brother, fellow worker and fellow soldier, who is also your messenger, whom you sent to take care of my needs.
PHIL|2|26|For he longs for all of you and is distressed because you heard he was ill.
PHIL|2|27|Indeed he was ill, and almost died. But God had mercy on him, and not on him only but also on me, to spare me sorrow upon sorrow.
PHIL|2|28|Therefore I am all the more eager to send him, so that when you see him again you may be glad and I may have less anxiety.
PHIL|2|29|Welcome him in the Lord with great joy, and honor men like him,
PHIL|2|30|because he almost died for the work of Christ, risking his life to make up for the help you could not give me.
PHIL|3|1|Finally, my brothers, rejoice in the Lord! It is no trouble for me to write the same things to you again, and it is a safeguard for you.
PHIL|3|2|Watch out for those dogs, those men who do evil, those mutilators of the flesh.
PHIL|3|3|For it is we who are the circumcision, we who worship by the Spirit of God, who glory in Christ Jesus, and who put no confidence in the flesh--
PHIL|3|4|though I myself have reasons for such confidence. If anyone else thinks he has reasons to put confidence in the flesh, I have more:
PHIL|3|5|circumcised on the eighth day, of the people of Israel, of the tribe of Benjamin, a Hebrew of Hebrews; in regard to the law, a Pharisee;
PHIL|3|6|as for zeal, persecuting the church; as for legalistic righteousness, faultless.
PHIL|3|7|But whatever was to my profit I now consider loss for the sake of Christ.
PHIL|3|8|What is more, I consider everything a loss compared to the surpassing greatness of knowing Christ Jesus my Lord, for whose sake I have lost all things. I consider them rubbish, that I may gain Christ
PHIL|3|9|and be found in him, not having a righteousness of my own that comes from the law, but that which is through faith in Christ--the righteousness that comes from God and is by faith.
PHIL|3|10|I want to know Christ and the power of his resurrection and the fellowship of sharing in his sufferings, becoming like him in his death,
PHIL|3|11|and so, somehow, to attain to the resurrection from the dead.
PHIL|3|12|Not that I have already obtained all this, or have already been made perfect, but I press on to take hold of that for which Christ Jesus took hold of me.
PHIL|3|13|Brothers, I do not consider myself yet to have taken hold of it. But one thing I do: Forgetting what is behind and straining toward what is ahead,
PHIL|3|14|I press on toward the goal to win the prize for which God has called me heavenward in Christ Jesus.
PHIL|3|15|All of us who are mature should take such a view of things. And if on some point you think differently, that too God will make clear to you.
PHIL|3|16|Only let us live up to what we have already attained.
PHIL|3|17|Join with others in following my example, brothers, and take note of those who live according to the pattern we gave you.
PHIL|3|18|For, as I have often told you before and now say again even with tears, many live as enemies of the cross of Christ.
PHIL|3|19|Their destiny is destruction, their god is their stomach, and their glory is in their shame. Their mind is on earthly things.
PHIL|3|20|But our citizenship is in heaven. And we eagerly await a Savior from there, the Lord Jesus Christ,
PHIL|3|21|who, by the power that enables him to bring everything under his control, will transform our lowly bodies so that they will be like his glorious body.
PHIL|4|1|Therefore, my brothers, you whom I love and long for, my joy and crown, that is how you should stand firm in the Lord, dear friends!
PHIL|4|2|I plead with Euodia and I plead with Syntyche to agree with each other in the Lord.
PHIL|4|3|Yes, and I ask you, loyal yokefellow, help these women who have contended at my side in the cause of the gospel, along with Clement and the rest of my fellow workers, whose names are in the book of life.
PHIL|4|4|Rejoice in the Lord always. I will say it again: Rejoice!
PHIL|4|5|Let your gentleness be evident to all. The Lord is near.
PHIL|4|6|Do not be anxious about anything, but in everything, by prayer and petition, with thanksgiving, present your requests to God.
PHIL|4|7|And the peace of God, which transcends all understanding, will guard your hearts and your minds in Christ Jesus.
PHIL|4|8|Finally, brothers, whatever is true, whatever is noble, whatever is right, whatever is pure, whatever is lovely, whatever is admirable--if anything is excellent or praiseworthy--think about such things.
PHIL|4|9|Whatever you have learned or received or heard from me, or seen in me--put it into practice. And the God of peace will be with you.
PHIL|4|10|I rejoice greatly in the Lord that at last you have renewed your concern for me. Indeed, you have been concerned, but you had no opportunity to show it.
PHIL|4|11|I am not saying this because I am in need, for I have learned to be content whatever the circumstances.
PHIL|4|12|I know what it is to be in need, and I know what it is to have plenty. I have learned the secret of being content in any and every situation, whether well fed or hungry, whether living in plenty or in want.
PHIL|4|13|I can do everything through him who gives me strength.
PHIL|4|14|Yet it was good of you to share in my troubles.
PHIL|4|15|Moreover, as you Philippians know, in the early days of your acquaintance with the gospel, when I set out from Macedonia, not one church shared with me in the matter of giving and receiving, except you only;
PHIL|4|16|for even when I was in Thessalonica, you sent me aid again and again when I was in need.
PHIL|4|17|Not that I am looking for a gift, but I am looking for what may be credited to your account.
PHIL|4|18|I have received full payment and even more; I am amply supplied, now that I have received from Epaphroditus the gifts you sent. They are a fragrant offering, an acceptable sacrifice, pleasing to God.
PHIL|4|19|And my God will meet all your needs according to his glorious riches in Christ Jesus.
PHIL|4|20|To our God and Father be glory for ever and ever. Amen.
PHIL|4|21|Greet all the saints in Christ Jesus. The brothers who are with me send greetings.
PHIL|4|22|All the saints send you greetings, especially those who belong to Caesar's household.
PHIL|4|23|The grace of the Lord Jesus Christ be with your spirit. Amen.
