ACTS|1|1|提阿非羅 啊，我在第一本書中已論到耶穌從開頭所做和所教導的一切事，
ACTS|1|2|直到他藉著聖靈吩咐所揀選的使徒後，被接上升的日子為止。
ACTS|1|3|他受害以後，用許多確據向使徒顯明自己是活著的，在四十天之中向他們顯現，並講說上帝國的事。
ACTS|1|4|耶穌和他們聚集的時候，囑咐他們說：「不要離開 耶路撒冷 ，但要等候父的應許，就是你們聽見我說過的。
ACTS|1|5|約翰 是用水施洗，但過了不多幾天，你們要在聖靈裏受洗。」
ACTS|1|6|他們聚集的時候，問耶穌：「主啊，你就要在這時候復興 以色列 國嗎？」
ACTS|1|7|耶穌對他們說：「父憑著自己的權柄所定的時候和日期，不是你們可以知道的。
ACTS|1|8|但聖靈降臨在你們身上，你們就必得著能力，並要在 耶路撒冷 、 猶太 全地和 撒瑪利亞 ，直到地極，作我的見證。」
ACTS|1|9|說了這些話，他們正看的時候，他被接上升，有一朵雲彩從他們眼前把他接去。
ACTS|1|10|他升上去的時候，他們定睛望天，看哪，有兩個人身穿白衣站在他們旁邊，
ACTS|1|11|說：「 加利利 人哪，你們為甚麼站著望天呢？這離開你們被接升天的耶穌，你們見他怎樣升上天去，他也要怎樣來臨。」
ACTS|1|12|有一座山，名叫 橄欖山 ，離 耶路撒冷 不遠，有安息日可行走的路程 。那時，門徒從那裏回 耶路撒冷 去，
ACTS|1|13|他們一進城，就上了所住的樓房；在那裏有 彼得 、 約翰 、 雅各 、 安得烈 、 腓力 、 多馬 、 巴多羅買 、 馬太 、 亞勒腓 的兒子 雅各 、激進黨的 西門 ，和 雅各 的兒子 猶大 。
ACTS|1|14|這些人和幾個婦人，包括耶穌的母親 馬利亞 ，和耶穌的兄弟，都同心合意地恆切禱告。
ACTS|1|15|那時，有許多人聚會，約有一百二十名， 彼得 在弟兄中間站起來，說：
ACTS|1|16|「諸位弟兄，聖經的話必須應驗。聖經中，聖靈曾藉 大衛 的口預先說到那領人來拿耶穌的 猶大 ；
ACTS|1|17|他本來算是我們中的一個，並且得了這一份使徒的職任。
ACTS|1|18|這人用他不義的代價買了一塊田，以後身子仆倒，肚腹崩裂，腸子都流出來。
ACTS|1|19|住在 耶路撒冷 的人都知道這事，所以按著他們當地的話把那塊田叫 亞革大馬 ，就是「血田」的意思。
ACTS|1|20|因為《詩篇》上寫著： 「願他的住處變為廢墟， 無人在內居住。」 又說： 「願別人得他的職分。」
ACTS|1|21|所以，主耶穌在我們中間出入的整段時間，就是從 約翰 施洗起，直到主離開我們被接上升的日子為止，必須從那常與我們一起的人中，立一位與我們同作耶穌復活的見證。」
ACTS|1|22|
ACTS|1|23|於是他們推舉兩個人，就是那叫 巴撒巴 ，又稱為 猶士都 的 約瑟 ，和 馬提亞 。
ACTS|1|24|眾人禱告說：「主啊，你知道萬人的心，求你從這兩個人中指明你所揀選的是哪一位，
ACTS|1|25|去得這使徒的職任；這職位 猶大 已經丟棄，往自己的地方去了。」
ACTS|1|26|於是眾人為他們搖籤，搖出 馬提亞 來；他就和十一個使徒同列。
ACTS|2|1|五旬節那日到了，他們全都聚集在一起。
ACTS|2|2|忽然，有響聲從天上下來，好像一陣大風吹過，充滿了他們所坐的整座屋子；
ACTS|2|3|又有舌頭如火焰向他們顯現，分開落在他們每個人身上。
ACTS|2|4|他們都被聖靈充滿，就按著聖靈所賜的口才說起別國的話來。
ACTS|2|5|那時，有從天下各國來的虔誠的 猶太 人，住在 耶路撒冷 。
ACTS|2|6|這聲音一響，許多人都來聚集，各人因為聽見門徒用他們各自的鄉談說話，就甚納悶，
ACTS|2|7|都詫異驚奇說：「看哪，這些說話的不都是 加利利 人嗎？
ACTS|2|8|我們每個人怎麼聽見他們說我們生來所用的鄉談呢？
ACTS|2|9|我們 帕提亞 人、 瑪代 人、 以攔 人，和住在 美索不達米亞 、 猶太 、 加帕多家 、 本都 、 亞細亞 、
ACTS|2|10|弗呂家 、 旁非利亞 、 埃及 的人，並靠近 古利奈 的 利比亞 一帶地方的人，僑居的 羅馬 人，
ACTS|2|11|包括 猶太 人和皈依 猶太 教的人， 克里特 人和 阿拉伯 人，都聽見他們用我們的鄉談講論上帝的大作為。」
ACTS|2|12|眾人就都驚奇困惑，彼此說：「這是甚麼意思呢？」
ACTS|2|13|還有人譏誚，說：「他們是灌滿了新酒吧！」
ACTS|2|14|彼得 和十一個使徒站起來，他就高聲向眾人說：「 猶太 人和所有住在 耶路撒冷 的人哪，這件事你們要知道，要側耳聽我的話。
ACTS|2|15|這些人並不像你們所想的喝醉了，因為現在才早晨九點鐘。
ACTS|2|16|這正是藉著先知 約珥 所說的：
ACTS|2|17|『上帝說： 在末後的日子， 我要將我的靈澆灌凡血肉之軀的。 你們的兒女要說預言； 你們的少年要見異象； 你們的老人要做異夢。
ACTS|2|18|在那些日子，我要把我的靈澆灌， 甚至給我的僕人和婢女， 他們要說預言。
ACTS|2|19|在天上，我要顯出奇事， 在地下，我要顯出神蹟， 有血，有火，有煙霧。
ACTS|2|20|太陽要變為黑暗， 月亮要變為血， 這都在主大而光榮的日子未到以前。
ACTS|2|21|那時，凡求告主名的都必得救。』
ACTS|2|22|「 以色列 人哪，你們要聽我這些話： 拿撒勒 人耶穌就是上帝以異能、奇事、神蹟向你們證明出來的人，這些事是上帝藉著他在你們中間施行，正如你們自己知道的。
ACTS|2|23|他既按著上帝確定的旨意和預知被交與人，你們就藉著不法之人的手把他釘在十字架上，殺了。
ACTS|2|24|上帝卻將死的痛苦解除，使他復活了，因為他原不能被死拘禁。
ACTS|2|25|大衛 指著他說： 『我看見 主常在我眼前， 他在我右邊，使我不至於動搖。
ACTS|2|26|所以我心裏歡喜，我的舌頭快樂， 而且我的肉身要安居在指望中。
ACTS|2|27|因你必不將我的靈魂撇在陰間， 也不讓你的聖者見朽壞。
ACTS|2|28|你已將生命的道路指示我， 必使我在你面前充滿快樂。』
ACTS|2|29|「諸位弟兄，先祖 大衛 的事，我可以坦然地對你們說：他死了，也埋葬了，而且他的墳墓直到今日還在我們這裏。
ACTS|2|30|既然 大衛 是先知，他知道上帝曾向他起誓，要從他的後裔中立一位坐在他的寶座上。
ACTS|2|31|他預先看見了，就講論基督的復活，說： 『他不被撇在陰間； 他的肉身也不見朽壞。』
ACTS|2|32|這耶穌，上帝已經使他復活了，我們都是這事的見證人。
ACTS|2|33|他既被高舉在上帝的右邊，又從父受了所應許的聖靈，就把你們所看見所聽見的，澆灌下來。
ACTS|2|34|大衛 並沒有升到天上，但他自己說： 『主對我主說： 你坐在我的右邊，
ACTS|2|35|等我使你的仇敵作你的腳凳。』
ACTS|2|36|故此， 以色列 全家當確實知道，你們釘在十字架上的這位耶穌，上帝已經立他為主，為基督了。」
ACTS|2|37|眾人聽見這話，覺得扎心，就對 彼得 和其餘的使徒說：「諸位弟兄，我們該怎樣做呢？」
ACTS|2|38|彼得 對他們說：「你們各人要悔改，奉耶穌基督的名受洗，使你們的罪得赦免，就會領受所賜的聖靈。
ACTS|2|39|因為這應許是給你們和你們的兒女，並一切在遠方的人，就是給所有主—我們的上帝所召來的人。」
ACTS|2|40|彼得 還用更多別的話作見證，勸勉他們說：「你們當救自己脫離這彎曲的世代。」
ACTS|2|41|於是領受他話的人，都受了洗；那一天，門徒約添了三千人。
ACTS|2|42|他們都專注於使徒的教導和彼此的團契，擘餅和祈禱。
ACTS|2|43|眾人都心存敬畏；使徒們 又行了許多奇事神蹟。
ACTS|2|44|信的人都聚在一處，凡物公用，
ACTS|2|45|又賣了田產和家業，照每一個人所需要的分給他們。
ACTS|2|46|他們天天同心合意恆切地在聖殿裏敬拜，且在家中 擘餅，存著歡喜坦誠的心用飯，
ACTS|2|47|讚美上帝，得全體百姓的喜愛。主將得救的人天天加給他們。
ACTS|3|1|下午三點鐘禱告的時候， 彼得 和 約翰 上聖殿去。
ACTS|3|2|一個從母腹裏就是瘸腿的人正被人抬來，他們天天把他放在聖殿的一個叫 美門 的門口，求進聖殿的人施捨。
ACTS|3|3|他看見 彼得 、 約翰 將要進聖殿，就求他們施捨。
ACTS|3|4|彼得 和 約翰 定睛看他， 彼得 說：「看著我們！」
ACTS|3|5|那人就注目看他們，指望從他們得著甚麼。
ACTS|3|6|彼得 卻說：「金銀我都沒有，但我把我有的給你：奉 拿撒勒 人耶穌基督的名起來 行走！」
ACTS|3|7|於是 彼得 拉著他的右手，扶他起來；他的腳和踝骨立刻健壯了，
ACTS|3|8|就跳起來，站著，又開始行走。他跟他們進了聖殿，邊走邊跳，讚美上帝。
ACTS|3|9|百姓都看見他又行走，又讚美上帝，
ACTS|3|10|認得他是那素常坐在聖殿的 美門 口求人施捨的，就因他所遇到的事滿心驚訝詫異。
ACTS|3|11|那人正在稱為 所羅門 的廊下，拉住 彼得 和 約翰 ，大家都覺得很驚訝，一齊跑到他們那裏。
ACTS|3|12|彼得 看見，就對百姓說：「 以色列 人哪，為甚麼因這事而驚訝呢？為甚麼定睛看我們，以為我們憑自己的能力和虔誠使這人行走呢？
ACTS|3|13|亞伯拉罕 的上帝、 以撒 的上帝、 雅各 的上帝，就是我們列祖的上帝，已經榮耀了他的僕人耶穌，這耶穌就是你們交付官府的那位， 彼拉多 決定要釋放他時，你們卻在 彼拉多 面前棄絕了他。
ACTS|3|14|你們棄絕了那聖潔公義者，反而要求釋放一個兇手給你們。
ACTS|3|15|你們殺了那生命的創始者，上帝卻叫他從死人中復活；我們都是這事的見證人。
ACTS|3|16|因信他的名，他的名使你們所看見所認識的這人健壯了；正是他所賜的信心使這人在你們眾人面前完全好了。
ACTS|3|17|「如今，弟兄們，我知道你們做這事是出於無知，你們的官長也是如此。
ACTS|3|18|但上帝藉著眾先知的口預先宣告過基督將要受害的事，就這樣應驗了。
ACTS|3|19|所以，你們當悔改歸正，使你們的罪得以塗去，
ACTS|3|20|這樣，那安舒的日子就必從主面前來到；主也必差遣所預定給你們的基督耶穌來臨。
ACTS|3|21|他必須留在天上，直到萬物復興的時候，就是上帝自古藉著聖先知的口所說的。
ACTS|3|22|摩西 曾說：『主—你們 的上帝要從你們弟兄中給你們興起一位先知像我，凡他向你們所說的一切，你們都要聽從。
ACTS|3|23|凡不聽從那先知的，必將從民中滅絕。』
ACTS|3|24|從 撒母耳 以來和後繼的眾先知，凡說預言的，也都曾宣告這些日子。
ACTS|3|25|你們是先知的子孫，也是上帝與你們 祖宗所立之約的子孫，就是對 亞伯拉罕 說：『地上萬族都將因你的後裔得福。』
ACTS|3|26|上帝既興起他的僕人，就先差他到你們這裏來，賜福給你們，使各人回轉，離開你們的邪惡。」
ACTS|4|1|彼得 和 約翰 正向百姓說話的時候，祭司們、守殿官和撒都該人來了，
ACTS|4|2|就很煩惱，因為使徒們教導百姓，傳揚在耶穌的事上證明有死人復活，
ACTS|4|3|於是下手拿住他們；因為天已經晚了，就把他們押在拘留所到第二天。
ACTS|4|4|但聽道的人有許多信了，男人的數目約有五千。
ACTS|4|5|第二天，官長、長老和文士在 耶路撒冷 聚集，
ACTS|4|6|又有 亞那 大祭司、 該亞法 、 約翰 、 亞歷山大 ，和大祭司的親族都在那裏。
ACTS|4|7|他們叫使徒站在中間，問他們：「你們憑甚麼能力，奉誰的名做這事呢？」
ACTS|4|8|那時， 彼得 被聖靈充滿，對他們說：「民間的官長和長老啊，
ACTS|4|9|倘若今日我們被查問是因為在殘障的人身上所行的善事，就是這人怎麼得了痊癒，
ACTS|4|10|那麼，你們大家和 以色列 全民都當知道，站在你們面前的這人得痊癒，是因你們所釘在十字架、上帝使他從死人中復活的 拿撒勒 人耶穌基督的名。
ACTS|4|11|這位耶穌是： 『你們匠人所丟棄的石頭， 已成了房角的頭塊石頭。』
ACTS|4|12|除他以外，別無拯救，因為在天下人間，沒有賜下別的名，我們可以靠著得救。」
ACTS|4|13|他們見 彼得 、 約翰 的膽量，又看出他們原是沒有學問的平民，就很驚訝，認出他們曾是跟耶穌一起的；
ACTS|4|14|又看見那治好了的人和他們一同站著，就無話可駁。
ACTS|4|15|於是他們吩咐他們兩人從議會退出，就彼此商議，
ACTS|4|16|說：「我們當怎樣辦這兩個人呢？因為他們誠然行了一件明顯的神蹟，凡住在 耶路撒冷 的人都知道，我們也不能否認。
ACTS|4|17|但為避免這事越發在民間傳揚，我們必須威嚇他們，叫他們不可再奉這名對任何人講論。」
ACTS|4|18|於是他們叫了兩人來，禁止他們，再不可奉耶穌的名講論或教導人。
ACTS|4|19|彼得 和 約翰 回答他們說：「聽從你們，不聽從上帝，在上帝面前合理不合理，你們自己判斷吧！
ACTS|4|20|我們所看見所聽見的，我們不能不說。」
ACTS|4|21|官長為百姓的緣故，想不出任何法子懲罰他們，只好威嚇一番就把他們釋放了；這是因眾人為了所行的奇事都歸榮耀與上帝。
ACTS|4|22|原來經歷這神蹟醫好的人有四十多歲了。
ACTS|4|23|二人既被釋放，就到自己的人那裏去，把祭司長和長老所說的話都告訴他們。
ACTS|4|24|他們聽見了，就同心合意地高聲向上帝說：「主宰啊！你是那創造天、地、海和其中萬物的；
ACTS|4|25|你曾藉著聖靈託你僕人—我們祖宗 大衛 的口說： 『外邦為甚麼擾動？ 萬民為甚麼謀算虛妄的事？
ACTS|4|26|地上的君王都站穩， 臣宰也聚集一處， 要對抗主，對抗主的受膏者 』。
ACTS|4|27|希律 和 本丟．彼拉多 ，同外邦人和 以色列 民，果然在這城裏聚集，要攻打你所膏的聖僕耶穌，
ACTS|4|28|做了你手和你旨意所預定必成就的事。
ACTS|4|29|主啊，現在求你鑒察，他們的威嚇，使你僕人放膽講你的道，
ACTS|4|30|伸出你的手來，讓醫治、神蹟、奇事藉著你聖僕耶穌的名行出來。」
ACTS|4|31|他們禱告完了，聚會的地方震動；他們都被聖靈充滿，放膽傳講上帝的道。
ACTS|4|32|許多信徒都一心一意，沒有一人說他的任何東西是自己的，都是大家公用。
ACTS|4|33|使徒以大能見證主耶穌 復活；眾人也都蒙了大恩。
ACTS|4|34|他們當中沒有一個缺乏的，因為凡有田產房屋的都賣了，把所賣的錢拿來，
ACTS|4|35|放在使徒腳前，照每人所需要的，分給每人。
ACTS|4|36|有一個 利未 人，名叫 約瑟 ，使徒稱他為 巴拿巴 （ 巴拿巴 翻出來就是安慰之子），生在 塞浦路斯 。
ACTS|4|37|他有田地，也賣了，把錢拿來，放在使徒腳前。
ACTS|5|1|有一個人，名叫 亞拿尼亞 ，同他的妻子 撒非喇 ，賣了田產，
ACTS|5|2|把錢私自留下一部分，他的妻子也知道，其餘的部分拿來放在使徒腳前。
ACTS|5|3|彼得 說：「 亞拿尼亞 ！為甚麼撒但充滿了你的心，使你欺騙聖靈，把賣田地的錢私自留下一部分呢？
ACTS|5|4|田地還沒有賣，不是你自己的嗎？既賣了，錢不是你作主嗎？你怎麼心裏會想這樣做呢？你不是欺騙人，是欺騙上帝！」
ACTS|5|5|亞拿尼亞 一聽見這些話，就仆倒，斷了氣；所有聽見的人都非常懼怕。
ACTS|5|6|有些年輕人起來，把他裹好，抬出去埋葬了。
ACTS|5|7|約過了三小時，他的妻子進來，還不知道所發生的事。
ACTS|5|8|彼得 對她說：「你告訴我，你們賣田地的錢就是這些嗎？」她說：「就是這些。」
ACTS|5|9|彼得 對她說：「你們為甚麼同謀來試探主的靈呢？你看，埋葬你丈夫之人的腳已到門口，他們也要把你抬出去。」
ACTS|5|10|她立刻仆倒在 彼得 腳前，斷了氣。那些年輕人進來，見她已經死了，就把她抬出去，埋在她丈夫旁邊。
ACTS|5|11|全教會和所有聽見這些事的人都非常懼怕。
ACTS|5|12|主藉使徒的手在民間行了許多神蹟奇事；他們都同心合意地聚集在 所羅門 的廊下。
ACTS|5|13|其餘的人沒有一個敢接近他們，百姓卻尊重他們。
ACTS|5|14|信主的人越發增添，連男帶女都很多，
ACTS|5|15|甚至有人將病人抬到街上，放在床上或褥子上，好讓 彼得 走過來的時候，或者影子投在一些人身上。
ACTS|5|16|還有許多人帶著病人和被污靈纏磨的，從 耶路撒冷 四圍的城鎮來，他們全都得了醫治。
ACTS|5|17|於是，大祭司採取行動，他和他所有一起的人，就是撒都該派的人，滿心忌恨，
ACTS|5|18|就下手拿住使徒，把他們押在公共拘留所內。
ACTS|5|19|但在夜間主的使者開了監門，領他們出來，說：
ACTS|5|20|「你們去，站在聖殿裏，把這生命的一切話講給百姓聽。」
ACTS|5|21|使徒聽了這話，天將亮的時候就進聖殿裏去教導人。大祭司和他一起的人來了，叫齊議會的人和 以色列 人的眾長老，然後派人到監牢裏去把使徒提出來。
ACTS|5|22|但差役到了，不見他們在監裏，就回來稟報，
ACTS|5|23|說：「我們看見監牢關得很緊，警衛也站在門外，但打開門來，裏面一個人都不見。」
ACTS|5|24|守殿官和祭司長聽了這些話，心裏困惑，不知這事將來如何。
ACTS|5|25|有一個人來稟報說：「你們押在監裏的人，現在站在聖殿裏教導百姓。」
ACTS|5|26|於是守殿官和差役去帶使徒來，並沒有用暴力，因為怕百姓用石頭打他們。
ACTS|5|27|他們把使徒帶來了，就叫他們站在議會前。大祭司問他們，
ACTS|5|28|說：「我們不是嚴嚴地禁止你們，不可奉這名教導人嗎？ 看，你們倒把你們的道理充滿了 耶路撒冷 ，想要叫這人的血歸到我們身上！」
ACTS|5|29|彼得 和眾使徒回答：「我們必須順從上帝，勝於順從人。
ACTS|5|30|你們掛在木頭上殺害的耶穌，我們祖宗的上帝已經使他復活了。
ACTS|5|31|上帝把他高舉在自己的右邊，使他作元帥，作救主，使 以色列 人得以悔改，並且罪得赦免。
ACTS|5|32|我們是這些事的見證人；上帝賜給順從的人的聖靈也為這些事作見證。」
ACTS|5|33|議會的人聽了極其惱怒，想要殺他們。
ACTS|5|34|但有一個法利賽人，名叫 迦瑪列 ，是眾百姓所敬重的律法教師，他在議會中站起來，吩咐人把使徒暫且帶到外面去，
ACTS|5|35|然後對眾人說：「 以色列 人哪，對於這些人，你們應當小心怎樣處理。
ACTS|5|36|從前 杜達 出現，自命不凡，附從他的人數約有四百；他被殺後，附從他的人全都散了，歸於無有。
ACTS|5|37|此後，登記戶籍的時候，又有 加利利 的 猶大 出現，引誘百姓跟從他，他也滅亡，附從他的人也都四散了。
ACTS|5|38|現在，我勸你們不要管這些人，任憑他們吧！他們所謀所為若是出於人，必要敗壞；
ACTS|5|39|若是出於上帝，你們就不能敗壞他們，恐怕你們倒是攻擊上帝了。」 議會的人被他說服了，
ACTS|5|40|就叫使徒來，把他們打了，又吩咐他們不可奉耶穌的名講道，然後把他們釋放了。
ACTS|5|41|他們歡歡喜喜地離開議會，因他們算配為這名受辱。
ACTS|5|42|他們就每日在聖殿裏，在家裏 ，不住地教導人，傳耶穌是基督的福音。
ACTS|6|1|那些日子，門徒增多，有說希臘話的 猶太 人向 希伯來 人發怨言，因為在日常的供給上忽略了他們的寡婦。
ACTS|6|2|十二使徒叫眾門徒來，說：「我們撇下上帝的道去管理飯食，是不合宜的。
ACTS|6|3|所以弟兄們，當從你們中間選出七個有好名聲、滿有聖靈和智慧，我們派他們管理這事。
ACTS|6|4|至於我們，我們要專注於祈禱和傳道的事奉。」
ACTS|6|5|這話使全會眾都喜悅，就揀選了 司提反 —他是一個滿有信心和聖靈的人；他們又揀選了 腓利 、 伯羅哥羅 、 尼迦挪 、 提門 、 巴米拿 ，並皈依 猶太 教的 安提阿 人 尼哥拉 ，
ACTS|6|6|叫他們站在使徒面前，使徒禱告後，就為他們按手。
ACTS|6|7|上帝的道興旺起來；在 耶路撒冷 門徒數目增加得很多，也有許多祭司聽從了這信仰。
ACTS|6|8|司提反 滿有恩惠和能力，在民間行了大奇事和神蹟。
ACTS|6|9|當時有從稱為「自由人」會堂，並 古利奈 、 亞歷山大 會堂來的人，還有些從 基利家 、 亞細亞 來的人，起來和 司提反 辯論。
ACTS|6|10|司提反 是以智慧和聖靈說話，眾人抵擋不住，
ACTS|6|11|就收買人來說：「我們聽見他說褻瀆 摩西 和上帝的話。」
ACTS|6|12|他們又煽動百姓、長老和文士，就突然來捉拿他，把他帶到議會去，
ACTS|6|13|設下假見證，說：「這個人不斷地說話，侮辱神聖的地方和律法。
ACTS|6|14|我們曾聽見他說，這 拿撒勒 人耶穌要毀壞這地方，也要改變 摩西 所交給我們的規矩。」
ACTS|6|15|在議會裏坐著的人都定睛看他，見他的面貌好像天使的面貌。
ACTS|7|1|大祭司說：「果真有這些事嗎？」
ACTS|7|2|司提反 說：「諸位父老弟兄請聽！從前我們的祖宗 亞伯拉罕 在 美索不達米亞 ，還沒有住在 哈蘭 的時候，榮耀的上帝向他顯現，
ACTS|7|3|對他說：『你要離開本地和親族，往我所要指示你的地去。』
ACTS|7|4|他就離開 迦勒底 人的地方，住在 哈蘭 。他父親死了以後，上帝使他從那裏搬到你們現在所住的地方。
ACTS|7|5|在這裏上帝並沒有給他產業，連立足的地方都沒有，但應許要將這地賜給他和他的後裔為業，雖然那時他還沒有兒子。
ACTS|7|6|上帝這樣說：『他的後裔必寄居外邦，那裏的人要使他們作奴隸，苦待他們四百年。』
ACTS|7|7|上帝又說：『但我要懲罰使他們作奴隸的那國。以後他們要出來，在這地方事奉我。』
ACTS|7|8|上帝又賜他割禮的約。於是 亞伯拉罕 生了 以撒 ，在第八日給他行了割禮；後來 以撒 生 雅各 ， 雅各 生十二位先祖。
ACTS|7|9|「先祖嫉妒 約瑟 ，把他賣到 埃及 去，上帝卻與他同在，
ACTS|7|10|救他脫離一切苦難，又使他在 埃及 王法老面前蒙恩，又有智慧。法老派他作 埃及 國的宰相兼管法老的全家。
ACTS|7|11|後來全 埃及 和 迦南 遭遇饑荒和大災難，我們的祖宗絕了糧。
ACTS|7|12|雅各 聽見在 埃及 有糧，就打發我們的祖宗初次往那裏去。
ACTS|7|13|第二次 約瑟 與兄弟們相認，法老才認識他的家族。
ACTS|7|14|約瑟 就打發人，請父親 雅各 和全族七十五個人都來。
ACTS|7|15|於是 雅各 下了 埃及 ，後來他和我們的祖宗都死在那裏；
ACTS|7|16|他們又被遷到 示劍 ，葬於 亞伯拉罕 在 示劍 用銀子從 哈抹 子孫 買來的墳墓裏。
ACTS|7|17|「當上帝應許 亞伯拉罕 的日期將到的時候， 以色列 人在 埃及 人丁興旺，
ACTS|7|18|直到另一位不認識 約瑟 的王興起統治 埃及 。
ACTS|7|19|他用詭計待我們的宗族，苦待我們的祖宗，強迫他們丟棄嬰孩，使嬰孩不能存活。
ACTS|7|20|就在那時， 摩西 生了下來，上帝看為俊美，在父親家裏被撫養了三個月。
ACTS|7|21|他被丟棄的時候，法老的女兒拾了去，當自己的兒子撫養。
ACTS|7|22|摩西 學了 埃及 人一切的學問，說話辦事都有才能。
ACTS|7|23|「他到了四十歲，心中起意去看望他的弟兄 以色列 人。
ACTS|7|24|他見他們中的一個人受冤屈，就庇護他，為那被壓迫的人報仇，打死了那 埃及 人。
ACTS|7|25|他以為他的弟兄們必明白上帝是藉他的手搭救他們，他們卻不明白。
ACTS|7|26|第二天，他遇見有人在打架，就想勸他們和好，說：『二位，你們是弟兄，為甚麼彼此欺負呢？』
ACTS|7|27|那欺負鄰舍的人把他推開，說：『誰立你作我們的領袖和審判官呢？
ACTS|7|28|難道你要殺我像昨天殺那 埃及 人一樣嗎？』
ACTS|7|29|摩西 聽見這話就逃走了，寄居於 米甸 地，在那裏生了兩個兒子。
ACTS|7|30|「過了四十年，在 西奈山 的曠野，有一位天使在荊棘的火焰中向 摩西 顯現。
ACTS|7|31|摩西 見了那異象，覺得很驚訝，正往前觀看的時候，有主的聲音說：
ACTS|7|32|『我是你列祖的上帝，就是 亞伯拉罕 、 以撒 、 雅各 的上帝。』 摩西 戰戰兢兢，不敢觀看。
ACTS|7|33|主對他說：『把你腳上的鞋脫下來，因為你所站的地方是聖地。
ACTS|7|34|我的百姓在 埃及 所受的困苦，我確實看見了；他們悲嘆的聲音，我也聽見了。我下來要救他們。現在，你來，我要差你往 埃及 去。』
ACTS|7|35|「這 摩西 就是有人曾棄絕他說『誰立你作我們的領袖和審判官』的，上帝卻藉那在荊棘中顯現的天使的手差派他作領袖，作解救者。
ACTS|7|36|這人領 以色列 人出來，在 埃及 地，在 紅海 ，在曠野的四十年間行了奇事神蹟。
ACTS|7|37|這人是 摩西 ，就是那曾對 以色列 人說『上帝要從你們弟兄中給你們興起一位先知像我』的。
ACTS|7|38|這人是那曾在曠野的會眾中和 西奈山 上，與那對他說話的天使同在，又與我們祖宗同在的，他領受了活潑的聖言傳給我們。
ACTS|7|39|我們的祖宗不肯聽從，反棄絕他，他們的心轉向 埃及 ，
ACTS|7|40|對 亞倫 說：『你為我們造神明，在我們前面引路，因為領我們出 埃及 地的這個 摩西 ，我們不知道他遭遇了甚麼事。』
ACTS|7|41|那時，他們造了一個牛犢，又拿祭物獻給那像，為自己手所做的工作歡躍。
ACTS|7|42|但是上帝轉臉不顧，任憑他們祭拜天上的日月星辰，正如先知書上所寫的： 『 以色列 家啊，你們四十年間在曠野， 何曾將犧牲和祭物獻給我？
ACTS|7|43|你們抬著 摩洛 的帳幕 和 理番 ──你們神明的星， 就是你們所造為要敬拜的像。 因此，我要把你們遷到 巴比倫 外去。』
ACTS|7|44|「我們的祖宗在曠野，有作證的會幕，是上帝吩咐 摩西 照著他所看見的樣式做的。
ACTS|7|45|這帳幕，我們的祖宗同 約書亞 相繼承受了，當上帝在他們面前趕走外邦人的時候，他們把這帳幕搬進承受為業之地，直存到 大衛 的日子。
ACTS|7|46|大衛 在上帝面前蒙恩，祈求為 雅各 的家 預備居所。
ACTS|7|47|但卻是 所羅門 為上帝造成殿宇。
ACTS|7|48|其實，至高者並不住人手所造的，就如先知所言：
ACTS|7|49|『主說：天是我的寶座， 地是我的腳凳。 你們要為我造怎樣的殿宇？ 哪裏是我安歇的地方呢？
ACTS|7|50|這一切不都是我手所造的嗎？』
ACTS|7|51|「你們這硬著頸項，心與耳未受割禮的人哪，時常抗拒聖靈！你們的祖宗怎樣，你們也怎樣。
ACTS|7|52|先知中有哪一個不是受你們祖宗的迫害呢？他們把預先宣告那義者要來的人殺了。如今你們成了那義者的出賣者和兇手了。
ACTS|7|53|你們領受了天使所傳佈的律法，竟不遵守。」
ACTS|7|54|眾人聽見這些話，心中極其惱怒，向 司提反 咬牙切齒。
ACTS|7|55|但 司提反 滿有聖靈，定睛望天，看見上帝的榮耀，又看見耶穌站在上帝的右邊，
ACTS|7|56|就說：「我看見天開了，人子站在上帝的右邊。」
ACTS|7|57|眾人大聲喊叫，摀著耳朵，齊心衝向他，
ACTS|7|58|把他推到城外，用石頭打他。作見證的人把他們的衣裳放在一個名叫 掃羅 的青年腳前。
ACTS|7|59|他們正用石頭打 司提反 的時候，他呼求說：「主耶穌啊，求你接納我的靈魂！」
ACTS|7|60|然後他跪下來，大聲喊著：「主啊，不要將這罪歸於他們！」說了這話，就長眠了。
ACTS|8|1|掃羅 也贊同處死他。從那一天開始， 耶路撒冷 的教會遭受到大迫害，除了使徒以外，眾門徒都分散在 猶太 和 撒瑪利亞 各處。
ACTS|8|2|有些虔誠的人把 司提反 埋葬了，為他大大哀哭。
ACTS|8|3|掃羅 卻殘害教會，挨家挨戶地進去，拉著男女關在監裏。
ACTS|8|4|那些分散的人往各地去傳福音的道。
ACTS|8|5|腓利 下 撒瑪利亞城 去 ，向當地人宣講基督。
ACTS|8|6|眾人都聚精會神，同心合意地聽 腓利 所說的話，一邊聽他的話，一邊看他所行的神蹟。
ACTS|8|7|因為有許多人被污靈附著，那些污靈大聲呼叫，從他們身上出來；還有許多癱瘓的、瘸腿的都得了醫治。
ACTS|8|8|那城裏，有極大的喜樂。
ACTS|8|9|有一個人名叫 西門 ，向來在那城裏行邪術，自命為大人物，使 撒瑪利亞 的居民驚奇。
ACTS|8|10|所有的人，從小到大都聽從他，說：「這個人就是上帝的能力，那稱為大能者的。」
ACTS|8|11|他們聽從他，因他很久以來用邪術使他們驚奇。
ACTS|8|12|當他們信了 腓利 所傳上帝國的福音和耶穌基督的名，連男帶女都受了洗。
ACTS|8|13|西門 自己也信了；既受了洗，就常與 腓利 在一處，看見他所行的神蹟和大異能，就覺得很驚奇。
ACTS|8|14|在 耶路撒冷 的使徒聽見 撒瑪利亞 人領受了上帝的道，就打發 彼得 和 約翰 到他們那裏去。
ACTS|8|15|兩個人下去，就為他們禱告，要讓他們領受聖靈，
ACTS|8|16|因為聖靈還沒有降在他們任何一個人身上，他們只奉主耶穌的名受了洗。
ACTS|8|17|於是使徒按手在他們頭上，他們就領受了聖靈。
ACTS|8|18|西門 看見使徒一按手，就有聖靈賜下，就拿錢給使徒，
ACTS|8|19|說：「請把這權柄也給我，使我手按著誰，誰就可以領受聖靈。」
ACTS|8|20|彼得 對他說：「你的銀子和你一同滅亡吧！因為你想上帝的恩賜是可以用錢買的。
ACTS|8|21|你在這道上無份無關；因為你在上帝面前心懷不正。
ACTS|8|22|你要為你這樣的惡而悔改，祈求主，或者你心裏的意念可得赦免。
ACTS|8|23|我看出你正在苦膽之中，被不義捆綁著。」
ACTS|8|24|西門 回答說：「請你們為我求主，使你們所說的，沒有一樣臨到我身上。」
ACTS|8|25|使徒既作了見證，並且宣講了主的道，就回 耶路撒冷 去，一路在 撒瑪利亞 好些村莊傳揚福音。
ACTS|8|26|有主的一個使者對 腓利 說：「起來！向南走，往那從 耶路撒冷 下 迦薩 的路上去。」那路是曠野。
ACTS|8|27|腓利 就起身去了。不料，有一個 埃塞俄比亞 人，是個有大權的太監，在 埃塞俄比亞 女王 甘大基 的手下總管銀庫，他上 耶路撒冷 去禮拜。
ACTS|8|28|回程中，他坐在車上，正念著 以賽亞 先知的書，
ACTS|8|29|聖靈對 腓利 說：「你去！靠近那車走。」
ACTS|8|30|腓利 就跑到太監那裏，聽見他正在念 以賽亞 先知的書，就說：「你明白你所念的嗎？」
ACTS|8|31|他說：「沒有人指教我，怎能明白呢？」於是他請 腓利 上車，與他同坐。
ACTS|8|32|他所念的那段經文是這樣： 「他像羊被牽去宰殺， 又像羔羊在剪毛的人手下無聲， 他也是這樣不開口。
ACTS|8|33|他卑微的時候，得不到公義的審判， 誰能述說他的身世？ 因為他的生命從地上被奪去。」
ACTS|8|34|太監回答 腓利 說：「請問，先知說這話是指誰，是指自己，還是指別人呢？」
ACTS|8|35|腓利 就開口，從這段經文開始，對他傳講耶穌的福音。
ACTS|8|36|二人正沿路往前走，到了有水的地方，太監說：「看哪！這裏有水，有甚麼能阻止我受洗呢？」
ACTS|8|37|
ACTS|8|38|於是他吩咐把車停下來， 腓利 和太監二人一同下到水裏， 腓利 就給他施洗。
ACTS|8|39|他們從水裏上來，主的靈把 腓利 提了去，太監再也看不見他了，就歡歡喜喜地上路。
ACTS|8|40|後來有人在 亞鎖都 遇見 腓利 ；他走遍那地方，在各城宣揚福音，一直到 凱撒利亞 。
ACTS|9|1|掃羅 不斷用威嚇兇悍的口氣向主的門徒說話。他去見大祭司，
ACTS|9|2|要求發信給 大馬士革 的各會堂，若是找著信奉這道的人，無論男女，都准他捆綁帶到 耶路撒冷 。
ACTS|9|3|掃羅 在途中，將到 大馬士革 的時候，忽然有一道光從天上下來，四面照射著他，
ACTS|9|4|他就仆倒在地，聽見有聲音對他說：「 掃羅 ！ 掃羅 ！你為甚麼迫害我？」
ACTS|9|5|他說：「主啊！你是誰？」主說：「我就是你所迫害的耶穌。
ACTS|9|6|起來！進城去，你應該做的事，必有人告訴你。」
ACTS|9|7|同行的人站在那裏，說不出話來，因為他們聽見聲音，卻看不見人。
ACTS|9|8|掃羅 從地上起來，睜開眼睛，竟不能看見甚麼。有人拉他的手，領他進了 大馬士革 。
ACTS|9|9|他三天甚麼都看不見，也不吃也不喝。
ACTS|9|10|那時，在 大馬士革 有一個門徒，名叫 亞拿尼亞 。主在異象中對他說：「 亞拿尼亞 ！」他說：「主啊，我在這裏。」
ACTS|9|11|主對他說：「起來！往那叫 直街 的路去，在 猶大 的家裏，去找一個 大數 人，名叫 掃羅 ；他正在禱告，
ACTS|9|12|在異象中 看見了一個人，名叫 亞拿尼亞 ，進來為他按手，讓他能再看得見。」
ACTS|9|13|亞拿尼亞 回答：「主啊，我聽見許多人講到這個人，說他怎樣在 耶路撒冷 多多苦待你的聖徒，
ACTS|9|14|並且他在這裏有從祭司長得來的權柄，要捆綁一切求告你名的人。」
ACTS|9|15|主對他說：「你只管去。他是我所揀選的器皿，要在外邦人、君王和 以色列 人面前宣揚我的名。
ACTS|9|16|我也要指示他，為我的名必須受許多的苦難。」
ACTS|9|17|亞拿尼亞 就去了，進入那家，把手按在 掃羅 身上，說：「 掃羅 弟兄，在你來的路上向你顯現的主，就是耶穌，打發我來，叫你能再看得見，又被聖靈充滿。」
ACTS|9|18|掃羅 的眼睛上立刻好像有鱗一般的東西掉下來，他就能再看得見，於是他起來，受了洗，
ACTS|9|19|吃過飯體力就恢復了。 掃羅 和 大馬士革 的門徒一起住了些日子，
ACTS|9|20|立刻在各會堂裏傳揚耶穌，說他是上帝的兒子。
ACTS|9|21|凡聽見的人都很驚奇，說：「在 耶路撒冷 殘害求告這名的不就是這個人嗎？他不是到這裏來要捆綁他們，帶到祭司長那裏去嗎？」
ACTS|9|22|但 掃羅 越發有能力，駁倒住在 大馬士革 的 猶太 人，證明耶穌是基督。
ACTS|9|23|過了好些日子， 猶太 人商議要殺 掃羅 ，
ACTS|9|24|但他們的計謀被 掃羅 知道了。他們晝夜在城門守候著要殺他。
ACTS|9|25|他的門徒就在夜間用筐子把他從城牆上縋了下去。
ACTS|9|26|掃羅 到了 耶路撒冷 ，想與門徒結交，大家卻都怕他，不信他是門徒。
ACTS|9|27|只有 巴拿巴 接待他，領他去見使徒，把他在路上怎麼看見主，主怎麼向他說話，他在 大馬士革 怎麼奉耶穌的名放膽傳道，都述說出來。
ACTS|9|28|於是 掃羅 在 耶路撒冷 同門徒出入來往，奉主的名放膽傳道，
ACTS|9|29|並和說 希臘 話的 猶太 人講論辯駁，他們卻想法子要殺他。
ACTS|9|30|弟兄們知道了，就帶他下 凱撒利亞 ，送他往 大數 去。
ACTS|9|31|那時， 猶太 、 加利利 、 撒瑪利亞 各處的教會都得平安，建立起來，凡事敬畏主，蒙聖靈的安慰，人數逐漸增多。
ACTS|9|32|彼得 在眾信徒中到處奔波的時候，也到了住在 呂大 的聖徒那裏。
ACTS|9|33|他在那裏遇見一個人，名叫 以尼雅 ，得了癱瘓，在褥子上躺了八年。
ACTS|9|34|彼得 對他說：「 以尼雅 ，耶穌基督醫好你了，起來！整理你的褥子吧。」他立刻就起來了。
ACTS|9|35|凡住 呂大 和 沙崙 的人都看見了他，就歸向主。
ACTS|9|36|在 約帕 有一個女門徒，名叫 大比大 ，翻出來的意思是 多加 ；她廣行善事，多施賙濟。
ACTS|9|37|當時，她患病死了，有人把她清洗後，停在樓上。
ACTS|9|38|呂大 原與 約帕 相近；門徒聽見 彼得 在那裏，就派兩個人去見他，央求他說：「請快到我們那裏去，不要耽延。」
ACTS|9|39|彼得 就起身和他們同去。他到了，就有人領他上樓。眾寡婦都站在 彼得 旁邊哭，拿 多加 與她們同在時所做的內衣外衣給他看。
ACTS|9|40|彼得 叫她們都出去，然後跪下禱告，轉身對著屍體說：「 大比大 ，起來！」她就睜開眼睛，看見 彼得 ，就坐了起來。
ACTS|9|41|彼得 伸手扶她起來，叫那些聖徒和寡婦都進來，把 多加 活活地交給他們。
ACTS|9|42|這事傳遍了 約帕 ，就有許多人信了主。
ACTS|9|43|此後， 彼得 在 約帕 一個皮革匠 西門 的家裏住了好些日子。
ACTS|10|1|在 凱撒利亞 有一個人名叫 哥尼流 ，是 意大利 營的百夫長。
ACTS|10|2|他是個虔誠人，他和全家都敬畏上帝。他多多賙濟百姓，常常向上帝禱告。
ACTS|10|3|有一天，約在下午三點鐘，他在異象中清楚看見上帝的一個使者進來，到他那裏，對他說：「 哥尼流 。」
ACTS|10|4|哥尼流 定睛看他，驚惶地說：「主啊，甚麼事？」天使對他說：「你的禱告和你的賙濟已達到上帝面前，蒙記念了。
ACTS|10|5|現在你要派人往 約帕 去，請一位稱為 彼得 的 西門 來。
ACTS|10|6|他住在一個皮革匠 西門 的家裏，房子就在海邊。」
ACTS|10|7|向他說話的天使離開後， 哥尼流 叫了兩個僕人和常伺候他的一個虔誠的兵來，
ACTS|10|8|把一切的事都講給他們聽，然後就派他們往 約帕 去。
ACTS|10|9|第二天，他們走路將近那城，約在正午， 彼得 上房頂去禱告。
ACTS|10|10|他覺得餓了，想要吃。那家的人正預備飯的時候， 彼得 魂遊象外，
ACTS|10|11|看見天開了，有一塊好像大布的東西降下，四角 吊著縋在地上，
ACTS|10|12|裏面有地上各樣四腳的走獸、爬蟲和天上的飛鳥。
ACTS|10|13|又有聲音對他說：「 彼得 ，起來！宰了吃。」
ACTS|10|14|彼得 卻說：「主啊，絕對不可！凡污俗和不潔淨的東西，我從來沒有吃過。」
ACTS|10|15|第二次有聲音再對他說：「上帝所潔淨的，你不可當作污俗的。」
ACTS|10|16|這樣一連三次，那東西隨即收回天上去了。
ACTS|10|17|正當 彼得 心裏困惑，不知所看見的異象是甚麼意思時， 哥尼流 所差來的人已經找到了 西門 的家，站在門外，
ACTS|10|18|喊著問有沒有一位稱為 彼得 的 西門 住在這裏。
ACTS|10|19|彼得 還在思考那異象的時候，聖靈對他說：「有三個人來找你。
ACTS|10|20|起來，下去，跟他們同去，不要疑惑，因為是我差他們來的。」
ACTS|10|21|於是 彼得 下去見那些人，說：「我就是你們要找的人，你們是為了甚麼緣故在這裏？」
ACTS|10|22|他們說：「百夫長 哥尼流 是個義人，敬畏上帝，為 猶太 全民族所稱讚。他蒙一位聖天使指示，叫他請你到他家裏去，要聽你講話。」
ACTS|10|23|彼得 就請他們進去住宿。 次日，他起身和他們同去，還有 約帕 的幾個弟兄跟他一起去。
ACTS|10|24|又次日，他 進入 凱撒利亞 ， 哥尼流 已經請了他的親朋好友在等候他們。
ACTS|10|25|彼得 一進去， 哥尼流 就迎接他，俯伏在他腳前拜他。
ACTS|10|26|但是 彼得 拉他起來，說：「你起來，我自己也不過是人。」
ACTS|10|27|彼得 和他一邊說話一邊進去，見有好些人聚集，
ACTS|10|28|就對他們說：「你們知道， 猶太 人和別國的人結交來往本是不合規矩的，但上帝已經指示我，無論甚麼人都不可看作污俗或不潔淨的。
ACTS|10|29|所以，我一被邀請，沒有推辭就來了。現在請問，你們為甚麼叫我來呢？」
ACTS|10|30|哥尼流 說：「四天前，這個時候，我在家中守著下午三點鐘的禱告，忽然有一個人穿著明亮的衣裳站在我面前，
ACTS|10|31|說：『 哥尼流 ，你的禱告已蒙垂聽，你的賙濟在上帝面前已蒙記念了。
ACTS|10|32|你要派人往 約帕 去，請那稱為 彼得 的 西門 來，他住在海邊一個皮革匠 西門 的家裏。』
ACTS|10|33|所以我立刻派人去請你。你來了真好。現在我們都在上帝面前，要聽主 吩咐你的一切話。」
ACTS|10|34|彼得 開口說：「我真的看出上帝是不偏待人的。
ACTS|10|35|不但如此，在各國中那敬畏他而行義的人都為他所悅納。
ACTS|10|36|上帝藉著耶穌基督—他是萬有的主—傳和平的福音，把這道傳給 以色列 人。
ACTS|10|37|這話在 約翰 傳揚洗禮以後，從 加利利 起，傳遍了 猶太 。上帝怎樣以聖靈和能力膏了 拿撒勒 人耶穌，這都是你們知道的。他到處奔波，行善事，醫好凡被魔鬼壓制的人，因為上帝與他同在。
ACTS|10|38|
ACTS|10|39|他在 猶太 人之地和 耶路撒冷 所行的一切事，有我們作見證人。他們竟把他掛在木頭上殺了。
ACTS|10|40|第三天，上帝使他復活，使他顯現出來；
ACTS|10|41|不是顯現給所有的人看，而是顯現給上帝預先所揀選為他作見證的人看，就是我們這些在他從死人中復活以後和他同吃同喝的人。
ACTS|10|42|他吩咐我們傳道給眾人，證明他是上帝所立定，要作審判活人、死人的審判者。
ACTS|10|43|眾先知也為這人作見證：凡信他的人，必藉著他的名得蒙赦罪。」
ACTS|10|44|彼得 還在說這些話的時候，聖靈降在一切聽道的人身上。
ACTS|10|45|那些奉割禮的信徒和 彼得 同來，見聖靈的恩賜也澆在外邦人身上，就都驚奇；
ACTS|10|46|因聽見他們說方言 ，稱讚上帝為大。於是 彼得 回答：
ACTS|10|47|「這些人既受了聖靈，跟我們一樣，誰能阻止用水給他們施洗呢？」
ACTS|10|48|他就吩咐奉耶穌基督的名給他們施洗。於是他們請 彼得 住了幾天。
ACTS|11|1|使徒和在 猶太 的眾弟兄聽到外邦人也領受了上帝的道。
ACTS|11|2|等到 彼得 上了 耶路撒冷 ，那些奉割禮的信徒和他爭辯，
ACTS|11|3|說：「你竟進入未受割禮之人當中，和他們一同吃飯！」
ACTS|11|4|彼得 就開始把這事逐一向他們解釋，說：
ACTS|11|5|「我在 約帕城 裏禱告的時候，魂遊象外，看見異象，有一塊好像大布的東西降下，四角吊著從天縋下，直來到我跟前。
ACTS|11|6|我定睛觀看，見內中有地上四腳的牲畜、野獸、爬蟲和天上的飛鳥。
ACTS|11|7|我還聽見有聲音對我說：『 彼得 ，起來！宰了吃。』
ACTS|11|8|我說：『主啊，絕對不可！凡污俗或不潔淨的東西從來沒有進過我的口。』
ACTS|11|9|第二次，有聲音從天上回答：『上帝所潔淨的，你不可當作污俗的。』
ACTS|11|10|這樣一連三次，然後一切就都收回天上去了。
ACTS|11|11|正當那時，有三個從 凱撒利亞 差來見我的人，站在我們 所住的屋子門前。
ACTS|11|12|聖靈吩咐我和他們同去，不要疑惑，還有這六位弟兄也跟我一起去，我們進了那人的家。
ACTS|11|13|那人就告訴我們，他如何看見一位天使站在他家裏，說：『你派人往 約帕 去，請那稱為 彼得 的 西門 來，
ACTS|11|14|他有話要告訴你，因這些話你和你的全家都可以得救。』
ACTS|11|15|我一開始講話，聖靈就降在他們身上，正像當初降在我們身上一樣。
ACTS|11|16|我就想起主的話如何說：『 約翰 用水施洗，但你們要在聖靈裏受洗。』
ACTS|11|17|既然上帝給他們恩賜，像在我們信主耶穌基督的時候給了我們一樣，我是誰，能攔阻上帝嗎？」
ACTS|11|18|眾人聽見這些話，就不說話了，只歸榮耀給上帝，說：「這樣看來，上帝也賜恩給外邦人，使他們悔改得生命了。」
ACTS|11|19|那些因 司提反 的事遭患難而四處分散的門徒，直走到 腓尼基 、 塞浦路斯 和 安提阿 。他們不向別人講道，只向 猶太 人講。
ACTS|11|20|但內中有 塞浦路斯 和 古利奈 人，他們到了 安提阿 也向 希臘 人傳講主耶穌的福音 。
ACTS|11|21|主的手與他們同在，信而歸主的人數很多。
ACTS|11|22|這風聲傳到 耶路撒冷 教會的人耳中，他們就打發 巴拿巴 到 安提阿 去。
ACTS|11|23|他到了那裏，看見上帝所賜的恩就歡喜，勸勉眾人要立定心志，恆久靠主。
ACTS|11|24|這 巴拿巴 原是個好人，滿有聖靈和信心，於是有許多人歸服了主。
ACTS|11|25|他又往 大數 去找 掃羅 ，
ACTS|11|26|找著了，就帶他到 安提阿 去。他們足有一年和教會一同聚集，教導了許多人。門徒稱為「基督徒」是從 安提阿 開始的。
ACTS|11|27|當那些日子，有幾位先知從 耶路撒冷 下到 安提阿 。
ACTS|11|28|內中有一位，名叫 亞迦布 ，站起來，藉著聖靈指示普天下將有大饑荒；這事在 克勞第 年間果然實現了。
ACTS|11|29|於是門徒決定，照各人的力量捐錢，送去供給住在 猶太 的弟兄。
ACTS|11|30|他們就這樣做了，託 巴拿巴 和 掃羅 的手送到眾長老那裏。
ACTS|12|1|約在那時候， 希律 王下手苦待教會中的一些人，
ACTS|12|2|用刀殺了 約翰 的哥哥 雅各 。
ACTS|12|3|他見 猶太 人喜歡這事，也去拿住 彼得 。那時候正是除酵節期間。
ACTS|12|4|希律 捉了 彼得 ，押在監裏，交給四班士兵看守，每班四個人，企圖要在逾越節後把他提出來，當著百姓辦他。
ACTS|12|5|於是 彼得 被囚在監裏，教會卻為他切切禱告上帝。
ACTS|12|6|希律 將要提他出來的前一夜， 彼得 被兩條鐵鏈鎖著，睡在兩個士兵當中；門前還有警衛看守。
ACTS|12|7|忽然，有主的一個使者顯現，牢房裏有光照耀；天使拍 彼得 的肋旁，叫醒了他，說：「快起來！」鐵鏈就從他手上脫落下來。
ACTS|12|8|天使對他說：「束上腰帶，穿上鞋子。」他就照著做了。天使又對他說：「披上外衣，跟我來。」
ACTS|12|9|彼得 就出來跟著他走，不知道天使所做是真的，以為見了異象。
ACTS|12|10|他們經過了第一層和第二層監牢，就來到往城內的鐵門，那門就自動給他們開了。他們出來，走過一條街，忽然天使離開他去了。
ACTS|12|11|彼得 清醒過來，說：「現在我真知道主差遣他的使者，救我脫離 希律 的手，和 猶太 人所期待的一切。」
ACTS|12|12|他明白了，就到那稱為 馬可 的 約翰 的母親 馬利亞 家去，在那裏已有好些人聚集禱告。
ACTS|12|13|彼得 敲外門時，有一個使女，名叫 羅大 ，出來應門，
ACTS|12|14|認出是 彼得 的聲音，歡喜得顧不了開門，就跑進去報信，說 彼得 站在門外。
ACTS|12|15|他們對她說：「你瘋了！」使女堅持真有其事。他們說：「那是他的天使。」
ACTS|12|16|彼得 不停地敲門；他們開了門，一見是他，就很驚奇。
ACTS|12|17|彼得 做個手勢，要他們不作聲，就告訴他們主怎樣領他出監；又說：「你們要把這些事告訴 雅各 和眾弟兄。」然後，他離開往別處去了。
ACTS|12|18|到了天亮，士兵中起了不少騷動，不知道 彼得 到哪裏去了。
ACTS|12|19|希律 找他，找不著，就審問警衛，下令帶走他們處死。後來 希律 離開 猶太 ，下 凱撒利亞 去，住在那裏。
ACTS|12|20|希律 向 推羅 和 西頓 的人發怒。他們那一帶地方是從王的土地供應糧食的，因此就託了王的內侍大臣 伯拉斯都 的情，一心來求和。
ACTS|12|21|希律 在所定的日子，穿上朝服，坐在位上，對他們演講。
ACTS|12|22|民眾一直喊著：「這是神明的聲音，不是人的聲音。」
ACTS|12|23|希律 不歸榮耀給上帝，所以主的使者立刻擊打他，他被蟲咬，就斷了氣。
ACTS|12|24|上帝的道日見興旺，越發廣傳。
ACTS|12|25|巴拿巴 和 掃羅 完成了供給的事，就回到 耶路撒冷 ，帶著稱為 馬可 的 約翰 同去。
ACTS|13|1|在 安提阿 的教會中，有幾位先知和教師，就是 巴拿巴 和稱為 尼結 的 西面 、 古利奈 人 路求 ，與 希律 分封王一起長大的 馬念 ，和 掃羅 。
ACTS|13|2|他們在事奉主和禁食的時候，聖靈說：「要為我分派 巴拿巴 和 掃羅 去做我召他們做的工作。」
ACTS|13|3|於是他們禁食禱告後，給 巴拿巴 和 掃羅 按手，然後派遣他們走了。
ACTS|13|4|他們既蒙聖靈差遣，就下到 西流基 ，從那裏坐船往 塞浦路斯 去，
ACTS|13|5|到了 撒拉米 ，就在 猶太 人各會堂裏宣講上帝的道，也有 約翰 作他們的幫手。
ACTS|13|6|他們走遍全島，直到 帕弗 ，在那裏遇見一個術士— 猶太 人的假先知，名叫 巴耶穌 。
ACTS|13|7|這人常和 士求．保羅 省長在一起。 士求．保羅 是個通達人，他請 巴拿巴 和 掃羅 來，要聽上帝的道。
ACTS|13|8|只是術士 以呂馬 (他的名字翻出來就是行法術的意思)敵對使徒，設法使省長遠離這信仰。
ACTS|13|9|掃羅 ，又名 保羅 ，被聖靈充滿，定睛看他，
ACTS|13|10|說：「你這充滿各樣詭詐奸惡，魔鬼的兒子，一切正義的仇敵，你還不停止扭曲主的正道嗎？
ACTS|13|11|現在你看，主的手臨到你身上，你會瞎眼，暫時看不見日光。」立刻迷濛和黑暗籠罩著他，他到處摸索，求人拉著手領他。
ACTS|13|12|省長看見所發生的事就信了，因對主的教導感到驚奇。
ACTS|13|13|保羅 和他的同伴從 帕弗 開船，來到 旁非利亞 的 別加 ， 約翰 卻離開他們，回 耶路撒冷 去了。
ACTS|13|14|他們從 別加 往前行，來到 彼西底 的 安提阿 。在安息日，他們進了會堂就坐下。
ACTS|13|15|在讀完了律法和先知的書，會堂主管們叫人過去，對他們說：「二位弟兄，你們若有甚麼勸勉眾人的話，請說。」
ACTS|13|16|保羅 就站起來，做個手勢，說：「諸位 以色列 人和一切敬畏上帝的人，請聽。
ACTS|13|17|這 以色列 民的上帝揀選了我們的祖宗，當百姓寄居 埃及 的時候抬舉他們，用大能的手領他們從那地出來。
ACTS|13|18|他在曠野容忍 他們，約有四十年。
ACTS|13|19|他消滅了 迦南 地七族的人後，把那地分給他們為業，
ACTS|13|20|約有四百五十年。此後 ，他給他們設立士師，直到 撒母耳 先知的時候。
ACTS|13|21|從那時起，他們要求立一個王，上帝就將 便雅憫 支派中 基士 的兒子 掃羅 給他們作王，共四十年。
ACTS|13|22|他廢了 掃羅 之後，就興起 大衛 作他們的王，又為他作見證說：『我尋得 耶西 的兒子 大衛 ，他是合我心意的人，他要遵行我一切的旨意。』
ACTS|13|23|從這人的後裔中，上帝已經照著所應許的為 以色列 人興起一位救主，就是耶穌。
ACTS|13|24|在他沒有出來以前， 約翰 已向 以色列 全民宣講悔改的洗禮。
ACTS|13|25|約翰 快走完他的人生路程時，說：『你們以為我是誰？我不是 ；但是有一位在我以後來的，我就是解他腳上的鞋帶也不配。』
ACTS|13|26|「諸位弟兄— 亞伯拉罕 的子孫和你們中間敬畏上帝的人哪，這救世的道是傳給我們的。
ACTS|13|27|耶路撒冷 的居民和他們的官長，因為不認識這基督，也不明白每安息日所讀的先知的書，把他定了死罪，正應驗了先知的預言。
ACTS|13|28|雖然他們查不出他有該死的罪狀，還是要求 彼拉多 把他殺了。
ACTS|13|29|他們既實現了經上指著他所記的一切話，就從木頭上把他取下來，放在墳墓裏。
ACTS|13|30|上帝卻使他從死人中復活。
ACTS|13|31|有許多日子，他向那些從 加利利 同他上 耶路撒冷 的人顯現，這些人如今在民間成為他的見證人。
ACTS|13|32|我們報好信息給你們，就是那應許祖宗的話，
ACTS|13|33|上帝已經向我們這些作他們兒女的 應驗，使耶穌復活了。正如《詩篇》第二篇上記著： 『你是我的兒子， 我今日生了你。』
ACTS|13|34|論到上帝使他從死人中復活，不再歸於朽壞，他曾這樣說： 『我必將所應許 大衛 那聖潔、 可靠的恩典賜給你們。』
ACTS|13|35|所以他也在另一篇說： 『你必不讓你的聖者見朽壞。』
ACTS|13|36|大衛 在世的時候，遵行了上帝的旨意就長眠了 ，歸到他祖宗那裏，已見朽壞；
ACTS|13|37|惟獨上帝使他復活的那一位，他並未見朽壞。
ACTS|13|38|所以弟兄們，你們當知道：赦罪的道是由這人傳給你們的，
ACTS|13|39|你們靠 摩西 的律法在不得稱義的一切事上，每一個信靠這位耶穌的都得稱義了。
ACTS|13|40|所以，你們要小心，免得先知書上所說的臨到你們：
ACTS|13|41|『要觀看，你們這些藐視的人， 要驚訝，要滅亡， 因為在你們的日子，我行一件事， 雖有人告訴你們，你們總是不信。』」
ACTS|13|42|他們走出會堂的時候，眾人請他們在下一個安息日再講這些話給他們聽。
ACTS|13|43|散會以後，有許多 猶太 人和敬虔的皈依 猶太 教的人跟從了 保羅 和 巴拿巴 。二人對他們講話，勸他們務要恆久倚靠上帝的恩典。
ACTS|13|44|到下一個安息日，全城的人幾乎都聚集起來，要聽主的道 。
ACTS|13|45|但 猶太 人看見這麼多的人，就滿心嫉妒，辯駁 保羅 所說的話，並且毀謗他。
ACTS|13|46|於是 保羅 和 巴拿巴 放膽說：「上帝的道本應先傳給你們；只因你們棄絕這道，斷定自己不配得永生，我們就轉向外邦人。
ACTS|13|47|因為主曾這樣吩咐我們： 『我已經立你作萬邦之光， 使你施行我的救恩，直到地極。』」
ACTS|13|48|外邦人聽見這話很歡喜，讚美主的道，凡被指定得永生的人都信了。
ACTS|13|49|於是主的道傳遍了那一帶地方。
ACTS|13|50|但 猶太 人挑唆虔敬尊貴的婦女和城內有名望的人，迫害 保羅 和 巴拿巴 ，把他們趕出境外。
ACTS|13|51|二人對著眾人跺掉腳上的塵土，然後往 以哥念 去了。
ACTS|13|52|門徒滿心喜樂，又被聖靈充滿。
ACTS|14|1|同樣的事也發生在 以哥念 。 保羅 和 巴拿巴 進了 猶太 人的會堂，在那裏講道，所以有很多 猶太 人和 希臘 人都信了。
ACTS|14|2|但那不順從的 猶太 人煽動外邦人，使他們心裏仇恨弟兄。
ACTS|14|3|二人在那裏住了好些日子，倚靠主放膽講道，主藉他們的手施行神蹟奇事，證明他恩惠的道。
ACTS|14|4|城裏的眾人卻分裂了：有依附 猶太 人的，有依附使徒的。
ACTS|14|5|那時，外邦人、 猶太 人和他們的官長，一齊擁上來，要凌辱使徒，用石頭打他們。
ACTS|14|6|使徒知道了，就逃到 呂高尼 的 路司得 和 特庇 兩個城，以及周圍地方去，
ACTS|14|7|在那裏繼續傳福音。
ACTS|14|8|路司得城 裏有一個兩腳無力的人，他從母腹裏就是瘸腿的，老是坐著，從來沒有走過。
ACTS|14|9|他聽 保羅 講道； 保羅 定睛看他，見他有信心，可得痊癒，
ACTS|14|10|就大聲說：「起來！兩腳站直。」那人就跳起來，開始行走。
ACTS|14|11|眾人看見 保羅 所做的事，就用 呂高尼 話大聲說：「有神明藉著人形降臨在我們中間了。」
ACTS|14|12|於是他們稱 巴拿巴 為 宙斯 ，稱 保羅 為 希耳米 ，因為他總是帶頭說話。
ACTS|14|13|城外有 宙斯 廟的祭司牽著牛，拿著花環，來到門前，要同眾人一起獻祭。
ACTS|14|14|巴拿巴 和 保羅 二位使徒聽見，就撕開衣裳，跳進眾人中間，喊著：
ACTS|14|15|「諸位，為甚麼做這些事呢？我們也是人，性情和你們一樣。我們傳福音給你們，是要你們離棄這些虛妄的事，歸向那創造天、地、海和其中萬物的永生的上帝。
ACTS|14|16|他在從前的世代，任憑萬國各行其道；
ACTS|14|17|然而他未嘗不為自己留下證據來，就如常行善事，從天降雨，賞賜豐年，使你們飲食飽足，滿心喜樂。」
ACTS|14|18|二人說了這些話，總算攔住眾人不獻祭給他們。
ACTS|14|19|但有些 猶太 人，從 安提阿 和 以哥念 來，挑唆眾人，並且用石頭打 保羅 ，以為他死了，就把他拖到城外。
ACTS|14|20|當門徒圍著他的時候，他站了起來，走進城去。第二天， 保羅 同 巴拿巴 往 特庇 去。
ACTS|14|21|保羅 和 巴拿巴 對那城裏的人傳了福音，使好些人成為門徒後，又回 路司得 、 以哥念 、 安提阿 去，
ACTS|14|22|堅固門徒的心，勸他們持守他們的信仰，說：「我們進入上帝的國，必須經歷許多艱難。」
ACTS|14|23|二人在各教會中選立了長老，禁食禱告後，把他們交託給他們所信的主。
ACTS|14|24|二人經過 彼西底 來到 旁非利亞 ，
ACTS|14|25|在 別加 講了道，就下 亞大利 去，
ACTS|14|26|從那裏坐船回 安提阿 去。當初，眾人就在這地方，把他們交託在上帝的恩典中，要完成現在所做的工。
ACTS|14|27|他們一到那裏，就聚集了會眾，述說上帝藉他們所行的一切事，並且上帝怎樣為外邦人開了信道的門。
ACTS|14|28|二人在那裏同門徒住了一段日子。
ACTS|15|1|有幾個人從 猶太 下來，教導弟兄們說：「你們若不按照 摩西 的規矩受割禮，不能得救。」
ACTS|15|2|保羅 和 巴拿巴 跟他們發生了激烈的爭執和辯論；大家就決定指派 保羅 、 巴拿巴 和本會的幾個人，為所辯論的事上 耶路撒冷 去見使徒和長老。
ACTS|15|3|於是教會為他們送行。他們經過 腓尼基 、 撒瑪利亞 ，沿途敘說外邦人歸主的事，使眾弟兄都非常歡喜。
ACTS|15|4|他們到了 耶路撒冷 ，教會、使徒和長老都接待他們，他們就述說上帝同他們所做的一切事。
ACTS|15|5|惟有幾個法利賽派的信徒起來，說：「必須給外邦人行割禮，吩咐他們遵守 摩西 的律法。」
ACTS|15|6|使徒和長老聚集商議這事。
ACTS|15|7|辯論了許久後， 彼得 站起來，對他們說：「諸位弟兄，你們知道上帝早已在你們中間揀選了我，讓外邦人從我口中得聽福音之道，而且相信。
ACTS|15|8|知道人心的上帝也為他們作了見證，賜聖靈給他們，正如給我們一樣；
ACTS|15|9|又藉著信潔淨了他們的心，他們和我們之間並沒有甚麼分別。
ACTS|15|10|現在你們為甚麼試探上帝，要把我們祖宗和我們所不能負的軛放在門徒的頸項上呢？
ACTS|15|11|相反地，我們相信，我們得救是因主耶穌的恩典，和他們一樣。」
ACTS|15|12|眾人都默默無聲，聽 巴拿巴 和 保羅 述說上帝藉著他們在外邦人中所行的神蹟和奇事。
ACTS|15|13|他們講完了， 雅各 回答說：「諸位弟兄，請聽我說。
ACTS|15|14|剛才 西門 述說上帝當初怎樣眷顧外邦人，從他們中間選取人民歸於自己的名下；
ACTS|15|15|眾先知的話也與這意思相符合。
ACTS|15|16|正如經上所寫的： 『此後，我要回來， 重新修造 大衛 倒塌了的帳幕， 從廢墟中重新修造， 把它建立起來，
ACTS|15|17|使剩餘的人， 就是凡稱我名的外邦人， 都尋求主。 這話是自古以來顯明這些事的主說的。』
ACTS|15|18|
ACTS|15|19|所以，我的意見是不可難為那歸向上帝的外邦人；
ACTS|15|20|但是要寫信吩咐他們禁戒偶像所玷污的東西、血和勒死的牲畜 ，禁戒淫亂。
ACTS|15|21|因為歷代以來， 摩西 的書在各城都有人宣講，每逢安息日，也在會堂裏誦讀。」
ACTS|15|22|那時，使徒、長老和全教會認為應從他們中間揀選人，差他們和 保羅 、 巴拿巴 一同到 安提阿 去，所揀選的就是稱為 巴撒巴 的 猶大 和 西拉 。這二人在弟兄中是領袖。
ACTS|15|23|他們帶去的信說：「使徒和作長老的弟兄們向 安提阿 、 敘利亞 、 基利家 外邦眾弟兄問安。
ACTS|15|24|我們聽說，有幾個人從我們這裏出去 ，用一些話騷擾你們，使你們的心困惑， 其實我們並沒有吩咐他們。
ACTS|15|25|我們認為，既然我們同心定意，就揀選幾個人，派他們同我們所親愛的 巴拿巴 和 保羅 到你們那裏去。
ACTS|15|26|這二人曾為我主耶穌基督的名不顧自己的性命。
ACTS|15|27|所以我們派 猶大 和 西拉 去，他們也會親口述說這些事。
ACTS|15|28|因為聖靈和我們決定除了這幾件重要的事，不將別的重擔放在你們身上，
ACTS|15|29|就是禁戒偶像所玷污的東西、血和勒死的牲畜，禁戒淫亂。這幾件你們若能自己禁戒就好了。祝你們安康！」
ACTS|15|30|他們既奉了差遣就下 安提阿 去，聚集會眾，把書信交給他們。
ACTS|15|31|眾人念了，因為信上鼓勵的話而感到欣慰。
ACTS|15|32|猶大 和 西拉 自己也是先知，就用許多話勸勉弟兄，堅固他們。
ACTS|15|33|二人住了些日子，弟兄們打發他們平平安安地回到差遣他們的人那裏去。
ACTS|15|34|
ACTS|15|35|但 保羅 和 巴拿巴 仍留在 安提阿 ，和許多別的人一同教導，並傳揚主的道。
ACTS|15|36|過了些日子， 保羅 對 巴拿巴 說：「讓我們回到從前宣揚主道的各城，看看弟兄們的情況如何。」
ACTS|15|37|巴拿巴 有意要帶稱為 馬可 的 約翰 同去；
ACTS|15|38|但 保羅 認為不宜帶他去，因為 馬可 從前在 旁非利亞 離開他們，不和他們一起工作。
ACTS|15|39|於是二人起了爭執，甚至彼此分手。 巴拿巴 帶著 馬可 ，坐船往 塞浦路斯 去；
ACTS|15|40|保羅 則揀選了 西拉 ，也出發了，蒙弟兄們把他交於主的恩典中。
ACTS|15|41|他就走遍了 敘利亞 、 基利家 ，堅固眾教會。
ACTS|16|1|後來， 保羅 來到 特庇 ，又到 路司得 。在那裏有一個門徒，名叫 提摩太 ，是信主的 猶太 婦人的兒子，他父親卻是 希臘 人。
ACTS|16|2|路司得 和 以哥念 的弟兄都稱讚他。
ACTS|16|3|保羅 要帶他同去，只因那些地方的 猶太 人都知道他父親是 希臘 人，就給他行了割禮。
ACTS|16|4|他們經過各城，把 耶路撒冷 使徒和長老所決定的規條交給門徒遵守。
ACTS|16|5|於是眾教會信心越發堅固，人數天天增加。
ACTS|16|6|因為聖靈禁止他們在 亞細亞 講道，他們就經過 弗呂家 、 加拉太 一帶地方。
ACTS|16|7|到了 每西亞 的邊界，他們想要往 庇推尼 去，耶穌的靈卻不許。
ACTS|16|8|他們就越過 每西亞 ，下 特羅亞 去。
ACTS|16|9|夜間，有異象向 保羅 顯現。有一個 馬其頓 人站著求他說：「請你過來，到 馬其頓 來幫助我們！」
ACTS|16|10|保羅 既看見這異象，我們就立即設法往 馬其頓 去，認為上帝呼召我們傳福音給那裏的人。
ACTS|16|11|我們從 特羅亞 開船，直行駛到 撒摩特喇 ，第二天到了 尼亞坡里 ；
ACTS|16|12|從那裏來到 腓立比 ，就是 馬其頓 這一帶的一個重要城市 ，也是 羅馬 的駐防城。我們在這城裏住了幾天。
ACTS|16|13|在安息日，我們出城門，到了河邊，知道那裏有一個禱告的地方 ，我們就坐下來對那些聚會的婦女講道。
ACTS|16|14|有一個賣紫色布的婦人，名叫 呂底亞 ，是 推雅推喇城 的人，素來敬拜上帝。她在聽著，主就開導她的心，使她留心聽 保羅 所講的話。
ACTS|16|15|她和她一家都領了洗，就求我們說：「你們若以為我是真心信主的 ，請到我家裏來住。」於是她堅決請我們留下。
ACTS|16|16|後來，我們往那禱告的地方去時，有一個被占卜的靈附身的使女迎面走來，她使用法術使她的主人們發了大財。
ACTS|16|17|她跟隨 保羅 和我們，喊著說：「這些人是至高上帝的僕人，對你們傳講救人的道路。」
ACTS|16|18|她一連好幾天這樣喊叫， 保羅 就心中厭煩，轉身對那靈說：「我奉耶穌基督的名吩咐你從她身上出來！」那靈立刻出來了。
ACTS|16|19|使女的主人們見發財的指望沒有了，就揪住 保羅 和 西拉 ，拉他們到市上去見官；
ACTS|16|20|又帶他們到行政官長們面前，說：「這些騷擾我們城的，他們是 猶太 人，
ACTS|16|21|竟傳佈我們 羅馬 人所不可接受、不可遵守的規矩。」
ACTS|16|22|群眾就一齊起來攻擊他們。官長們吩咐撕開他們的衣裳，用棍子打；
ACTS|16|23|打了許多棍，就把他們下在監裏，囑咐獄警嚴緊看守。
ACTS|16|24|獄警領了這樣的命令，就把他們下在內監，兩腳拴在木架上。
ACTS|16|25|約在半夜， 保羅 和 西拉 正在禱告，唱詩讚美上帝，眾囚犯也側耳聽著的時候，
ACTS|16|26|忽然，地大震動，甚至監牢的地基都搖動了，監門立刻全開，眾囚犯的鎖鏈也都解開了。
ACTS|16|27|獄警一醒，看見監門全開，以為囚犯已經逃走，就拔刀要自殺。
ACTS|16|28|保羅 大聲呼叫：「不要傷害自己！我們都在這裏。」
ACTS|16|29|獄警叫人拿燈來，就衝進去，戰戰兢兢地俯伏在 保羅 和 西拉 面前。
ACTS|16|30|然後獄警領他們出來，說：「二位先生，我必須做甚麼才可以得救？」
ACTS|16|31|他們說：「當信主耶穌，你和你一家都必得救 。」
ACTS|16|32|他們就把主的道講給他和他全家的人聽。
ACTS|16|33|當夜，就在那時候，獄警把他們帶去，洗他們的傷；他和他所有的家人立刻都受了洗。
ACTS|16|34|於是獄警領他們上自己的家裏去，給他們擺上飯。他和全家的人，因為信了上帝，都滿心喜樂。
ACTS|16|35|到了天亮，官長們打發差役來，說：「釋放那兩個人吧。」
ACTS|16|36|獄警就把這些話告訴 保羅 ：「官長們打發人來，要釋放你們，現在可以出監，平平安安去吧。」
ACTS|16|37|保羅 卻說：「我們是 羅馬 人，並沒有定罪，他們竟在公眾面前打了我們，又把我們下在監裏；現在要私下趕我們出去嗎？這不行！叫他們自己來領我們出去吧！」
ACTS|16|38|差役把這些話回稟官長們；官長們聽見他們是 羅馬 人，就害怕了，
ACTS|16|39|於是來勸他們，領他們出來，請他們離開那城。
ACTS|16|40|二人出了監牢，往 呂底亞 家裏去，見了弟兄們，勸慰他們一番，就離開了。
ACTS|17|1|保羅 和 西拉 經過 暗妃坡里 、 亞波羅尼亞 ，來到 帖撒羅尼迦 ，在那裏有 猶太 人的會堂。
ACTS|17|2|保羅 照他素常的規矩進去，一連三個安息日，根據聖經與他們辯論，
ACTS|17|3|講解和說明基督必須受害，從死人中復活；又說：「我所傳給你們的這位耶穌就是基督。」
ACTS|17|4|他們中間有些人聽了勸，就跟從 保羅 和 西拉 ，還有許多虔敬的 希臘 人，尊貴的婦女也不少。
ACTS|17|5|但不信的 猶太 人心裏嫉妒，聚集了些市井流氓，搭夥成群，煽動全城的人闖進 耶孫 的家，要把 保羅 和 西拉 帶到民眾那裏。
ACTS|17|6|那些人找不著他們，就把 耶孫 和幾個弟兄拉到地方官那裏，喊叫著：「這些攪亂天下的人也到這裏來了，
ACTS|17|7|耶孫 竟收留他們。這些人都違背凱撒的命令，說另有一個王耶穌。」
ACTS|17|8|眾人和地方官聽見這些話，就惶恐了，
ACTS|17|9|於是收了 耶孫 和其餘的人的保證金後，釋放了他們。
ACTS|17|10|當夜，弟兄們立刻送 保羅 和 西拉 往 庇哩亞 去；二人到了，就進入 猶太 人的會堂。
ACTS|17|11|這地方的 猶太 人比 帖撒羅尼迦 的人開明，熱心領受這道，天天查考聖經，要知道這道是否真實。
ACTS|17|12|所以，他們中間有許多信了，又有 希臘 的尊貴婦人，男人也不少。
ACTS|17|13|但 帖撒羅尼迦 的 猶太 人知道 保羅 又在 庇哩亞 傳上帝的道，就往那裏去，煽動挑撥群眾。
ACTS|17|14|於是，弟兄們立刻送 保羅 到海邊去， 西拉 和 提摩太 卻仍留在 庇哩亞 。
ACTS|17|15|護送 保羅 的人帶他到了 雅典 ，他們領了 保羅 的命令，叫 西拉 和 提摩太 趕快到他那裏來，然後回去了。
ACTS|17|16|保羅 在 雅典 等候他們的時候，看見滿城都是偶像，就心裏非常難過。
ACTS|17|17|於是他在會堂裏與 猶太 人和虔敬的人，以及每日在市場上所遇見的人辯論。
ACTS|17|18|還有 伊壁鳩魯 和 斯多亞 兩派的哲學家也與他爭辯。有的說：「這胡言亂語的要說甚麼？」有的說：「他似乎是宣傳外邦鬼神的。」這是因 保羅 傳講耶穌與復活的福音。
ACTS|17|19|他們就把他帶到 亞略巴古 ，說：「你所講的這新學說，我們也可以知道嗎？
ACTS|17|20|因為你有些奇怪的事傳到我們耳中，我們想知道這些事是甚麼意思。」
ACTS|17|21|原來所有的 雅典 人和居住在那裏的外國人都無暇管別的事，只是談談或聽聽新聞。
ACTS|17|22|保羅 站在 亞略巴古 當中，說：「諸位 雅典 人！我看你們凡事很敬畏鬼神。
ACTS|17|23|我到處走走的時候，仔細觀察你們所敬拜的，發現一座壇，上面寫著『獻給未識之神明』。你們所不認識而敬拜的，我現在向你們宣告：
ACTS|17|24|他是創造宇宙和其中萬物的上帝；他既是天地的主，就不住在人手所造的殿宇裏，
ACTS|17|25|也不用人手去服侍，好像缺少甚麼似的；自己倒將生命、氣息、萬物賜給萬人。
ACTS|17|26|他從一人 造出萬族，居住在全地面上，並且預先定準他們的年限和所住的疆界，
ACTS|17|27|為要使他們尋求上帝，或者可以揣摩而找到他，其實他離我們各人不遠。
ACTS|17|28|我們生活、行動、存在都在於他。就如你們的詩人也有人說：『我們也是他所生的。』
ACTS|17|29|既然我們是上帝所生的，就不應該以為上帝的神性像人用手藝和心思所雕刻的金、銀、石像一般。
ACTS|17|30|世人蒙昧無知的時候，上帝並不追究，如今卻吩咐各處的人都要悔改。
ACTS|17|31|因為他已經定了日子，要藉著他所設立的人按公義審判天下，並且使他從死人中復活，給萬人作可信的憑據。」
ACTS|17|32|眾人聽見死人復活的話，就有人譏誚他；又有人說：「我們會再聽你講這事。」
ACTS|17|33|於是 保羅 從他們當中出去了。
ACTS|17|34|但有幾個人依附他，信了主，其中有 亞略巴古 的議員 丟尼修 ，和一個名叫 大馬哩 的婦人，還有幾個與他們一起的人。
ACTS|18|1|這些事以後， 保羅 離開 雅典 ，來到 哥林多 。
ACTS|18|2|他遇見一個生在 本都 的 猶太 人，名叫 亞居拉 。不久前，他帶著妻子 百基拉 從 意大利 來，因為 克勞第 命令所有的 猶太 人都離開 羅馬 。 保羅 去投靠他們。
ACTS|18|3|他們本是製造帳棚為業。 保羅 因與他們同業，就和他們同住，一同做工。
ACTS|18|4|每逢安息日， 保羅 在會堂裏辯論，勸導 猶太 人和 希臘 人。
ACTS|18|5|西拉 和 提摩太 從 馬其頓 來的時候， 保羅 正專心傳道，向 猶太 人證明耶穌是基督。
ACTS|18|6|當他們抗拒他、毀謗他的時候，他就抖掉衣裳的灰塵，對他們說：「你們的罪歸到你們自己的頭上，與我無干。從今以後，我要往外邦人那裏去。」
ACTS|18|7|於是他離開那裏，到了一個人的家裏，他名叫 提多．猶士都 ，是敬拜上帝的人，他的家靠近會堂。
ACTS|18|8|會堂的主管 基利司布 和全家都信了主，還有許多 哥林多 人聽了就信，而且受了洗。
ACTS|18|9|夜間，主在異象中對 保羅 說：「不要怕，只管講，不要沉默，
ACTS|18|10|有我與你同在，沒有人會下手害你，因為在這城裏有許多屬我的人。」
ACTS|18|11|保羅 在那裏住了一年六個月，將上帝的道教導他們。
ACTS|18|12|到 迦流 作 亞該亞 省長的時候， 猶太 人齊心起來攻擊 保羅 ，拉他到法庭，
ACTS|18|13|說：「這個人教唆人不按著律法敬拜上帝。」
ACTS|18|14|保羅 剛要開口， 迦流 對 猶太 人說：「你們這些 猶太 人哪！如果是為冤枉或奸惡的事，我理當耐性聽你們。
ACTS|18|15|既然你們所爭論的是關乎用字、名目和你們的律法，你們自己去辦吧！這樣的事我不願意審問。」
ACTS|18|16|於是，他把他們逐出法庭。
ACTS|18|17|眾人就揪住會堂的主管 所提尼 ，在法庭前打他。這些事 迦流 都不管。
ACTS|18|18|保羅 又住了好些日子，就辭別了弟兄，坐船到 敘利亞 去。 百基拉 、 亞居拉 和他同去。他因為許過願，就在 堅革哩 剃了頭髮。
ACTS|18|19|到了 以弗所 ， 保羅 就把他們留在那裏，自己進了會堂，和 猶太 人辯論。
ACTS|18|20|眾人請他多住些日子，他沒有答應，
ACTS|18|21|就辭別他們，說：「上帝若許可，我還要回到你們這裏來。」於是他上船離開 以弗所 。
ACTS|18|22|他在 凱撒利亞 下了船，上 耶路撒冷 去問候教會，隨後下 安提阿 去。
ACTS|18|23|他在那裏住了些日子，又離開了那裏，逐一經過 加拉太 和 弗呂家 各地方，堅固眾門徒。
ACTS|18|24|有一個生在 亞歷山大 的 猶太 人，名叫 亞波羅 ，來到 以弗所 ，他很有口才，很會講解聖經。
ACTS|18|25|這人已經在主的道路上受了訓練，心裏火熱，精確地講論和教導耶穌的事；可是他只知道 約翰 的洗禮。
ACTS|18|26|他開始在會堂裏放膽講道； 百基拉 、 亞居拉 聽見，就接他來，將上帝的道路 給他更精確地講解。
ACTS|18|27|他想要往 亞該亞 去，弟兄們就勉勵他，並寫信請門徒們接待他，他到了那裏，多多幫助那些蒙恩信主的人，
ACTS|18|28|因為他在公眾面前極力駁倒 猶太 人，引聖經證明耶穌是基督。
ACTS|19|1|亞波羅 在 哥林多 的時候， 保羅 經過了內陸地區，來到 以弗所 ，在那裏他遇見幾個門徒，
ACTS|19|2|問他們：「你們信的時候領受了聖靈沒有？」他們說：「沒有，我們連甚麼是聖靈都沒有聽過。」
ACTS|19|3|保羅 說：「這樣，你們受的是甚麼洗呢？」他們說：「是受了 約翰 的洗。」
ACTS|19|4|保羅 說：「 約翰 所施的是悔改的洗禮，他告訴百姓當信那在他以後要來的那位，就是耶穌。」
ACTS|19|5|他們聽見這話以後，就奉主耶穌的名受洗。
ACTS|19|6|保羅 給他們按手，聖靈就降在他們身上，他們開始說方言 和說預言。
ACTS|19|7|他們約有十二個人。
ACTS|19|8|保羅 進會堂，一連三個月放膽講道，辯論上帝國的事，勸導眾人。
ACTS|19|9|後來，有些人心裏剛硬不信，在眾人面前毀謗這道； 保羅 就離開他們，也叫門徒與他們分開，就在 推喇奴 的講堂天天辯論。
ACTS|19|10|這樣有兩年之久，使一切住在 亞細亞 的，無論是 猶太 人是 希臘 人，都聽見主的道。
ACTS|19|11|上帝藉 保羅 的手行了些奇異的神蹟，
ACTS|19|12|甚至有人從 保羅 身上拿走手巾或圍裙放在病人身上，病就消除了，邪靈也出去了。
ACTS|19|13|那時，有幾個巡迴各處念咒趕鬼的 猶太 人，擅自利用主耶穌的名，向那些被邪靈所附的人說：「我奉 保羅 所傳的耶穌命令你們出來！」
ACTS|19|14|做這事的是 猶太 祭司長 士基瓦 的七個兒子。
ACTS|19|15|但邪靈回答他們：「耶穌我知道， 保羅 我也認識，你們卻是誰呢？」
ACTS|19|16|被邪靈所附的人就撲到他們身上，制伏他們，勝過他們，使他們赤著身子，受了傷，從那房子裏逃出去了。
ACTS|19|17|凡住在 以弗所 的，無論是 猶太 人是 希臘 人，都知道這件事，也都懼怕；主耶穌的名從此就更被尊為大了。
ACTS|19|18|許多已經信的人來承認並公開自己所行的事。
ACTS|19|19|又有許多平素行邪術的人把他們的書都拿來，堆積在眾人面前焚燒。他們計算書價，得知共值五萬塊銀錢。
ACTS|19|20|這樣，主的道大大興旺，而且普遍傳開了。
ACTS|19|21|這些事過後， 保羅 心裏決定要經過 馬其頓 、 亞該亞 ，就往 耶路撒冷 去。他說：「我到了那裏以後，也必須到 羅馬 去看看。」
ACTS|19|22|於是他差遣兩個助手 提摩太 和 以拉都 往 馬其頓 去，自己暫時留在 亞細亞 。
ACTS|19|23|那時，因這道路而起的騷動不小。
ACTS|19|24|有一個銀匠，名叫 底米丟 ，是製造 亞底米 神銀龕的，他使從事這手藝的人生意發達。
ACTS|19|25|他聚集他們和同行的工人，說：「諸位，你們知道我們是倚靠這生意發財的。
ACTS|19|26|你們看到，也聽見這 保羅 不但在 以弗所 ，也幾乎在 亞細亞 全地，引誘迷惑了許多人，說：『人手所做的不是神明。』
ACTS|19|27|這樣，不僅我們這行業陷入被藐視的危險，就是大女神 亞底米 的廟也要被人輕看，連 亞細亞 全地和普天下所敬拜的女神的威望也受損害了。」
ACTS|19|28|眾人聽見，就怒氣沖沖，喊著說：「大哉， 以弗所 人的 亞底米 ！」
ACTS|19|29|於是滿城都騷動起來。眾人抓住與 保羅 同行的 馬其頓 人 該猶 和 亞里達古 ，齊心衝進劇場。
ACTS|19|30|保羅 想要進到民眾那裏，門徒卻不許他去。
ACTS|19|31|連 亞細亞 的幾位官員，是 保羅 的朋友，也打發人來勸他不要冒險到劇場裏去。
ACTS|19|32|聚集的人亂成一團，有的喊這個，有的喊那個，大半不知道為了甚麼聚集。
ACTS|19|33|猶太 人把 亞歷山大 推出去，人群中有人慫恿他，他就做手勢，要向民眾申訴。
ACTS|19|34|但他們一認出他是 猶太 人，大家就異口同聲喊著：「大哉， 以弗所 人的 亞底米 ！」約喊了兩小時。
ACTS|19|35|城裏的書記官安撫了群眾後，說：「 以弗所 人哪，誰不知道 以弗所 人的城是看守大 亞底米 的廟和從 宙斯 那裏落下來的像的守護者呢？
ACTS|19|36|既然這些事是駁不倒的，你們就要安靜下來，不可妄動。
ACTS|19|37|你們把這些人帶來，他們並沒有偷竊廟中之物，也沒有褻瀆我們的女神。
ACTS|19|38|如果 底米丟 和他同行的手藝人有控告的事，自有公堂，也有省長，他們可以彼此控告。
ACTS|19|39|你們若有別的事請求，可以在合法的集會裏解決。
ACTS|19|40|今日的擾亂本是無緣無故的，有被控告的危險。這次的騷動，我們也說不出理由來。」
ACTS|19|41|他說完這些話，就叫眾人散會。
ACTS|20|1|騷亂平定以後， 保羅 請門徒來，勸勉了他們，就辭別他們，往 馬其頓 去。
ACTS|20|2|他走遍那一帶地方，用許多話勸勉門徒，然後來到 希臘 ，
ACTS|20|3|在那裏住了三個月。他快要坐船往 敘利亞 去的時候， 猶太 人設計害他，他就決定從 馬其頓 回去。
ACTS|20|4|同他到 亞細亞 去的，有 庇哩亞 人 畢羅斯 的兒子 所巴特 ， 帖撒羅尼迦 人 亞里達古 和 西公都 ，還有 特庇 人 該猶 和 提摩太 ，又有 亞細亞 人 推基古 和 特羅非摩 。
ACTS|20|5|這些人先走，在 特羅亞 等候我們。
ACTS|20|6|過了除酵節的日子，我們從 腓立比 開船，五天以後到了 特羅亞 ，和他們相會，在那裏住了七天。
ACTS|20|7|七日的第一日，我們聚會擘餅的時候， 保羅 因次日要起行，就為他們講道，直講到半夜。
ACTS|20|8|我們聚會的那座樓上有好些燈火。
ACTS|20|9|有一個少年，名叫 猶推古 ，坐在窗口上，沉沉入睡。 保羅 講了多時，少年睡熟了，從三層樓上掉下去，扶起來時已經死了。
ACTS|20|10|保羅 下去，伏在他身上，抱著他，說：「你們不要慌亂，他還有氣呢！」
ACTS|20|11|保羅 又上樓去，擘餅，吃了，再講了許久，直到天亮才離開。
ACTS|20|12|他們把那活過來的孩子帶走，大家得到很大的安慰。
ACTS|20|13|我們先上船，起航往 亞朔 去，想要在那裏接 保羅 ；因為他是這樣安排的，他自己本來打算要走陸路。
ACTS|20|14|他既在 亞朔 與我們相會，我們就接他上船，來到 米推利尼 。
ACTS|20|15|我們從那裏開船，第二天到了 基阿 的對岸；再下一天，在 撒摩 靠岸，又過了一天，到了 米利都 。
ACTS|20|16|因為 保羅 早已決定要越過 以弗所 ，免得在 亞細亞 耽延，他急忙前行，假如可能的話，在五旬節前能趕到 耶路撒冷 。
ACTS|20|17|保羅 從 米利都 打發人往 以弗所 去，請教會的長老來。
ACTS|20|18|他們來了， 保羅 對他們說：「你們自己知道，自從我到 亞細亞 的第一天，我怎樣跟你們相處，
ACTS|20|19|怎樣凡事謙卑，以眼淚服侍主，又因 猶太 人的謀害經歷試煉。
ACTS|20|20|你們也知道，凡對你們有益的，我沒有一樣隱瞞不說的，或在公眾面前，或在每一個人的家裏，我都教導你們，
ACTS|20|21|不論 猶太 人和 希臘 人，我都已證明他們當在上帝面前悔改，信靠我們的主耶穌。
ACTS|20|22|現在我被聖靈催迫 要往 耶路撒冷 去，雖然不知道在那裏會遭遇甚麼事，
ACTS|20|23|但知道聖靈在各城裏向我指證，說有捆鎖與患難等著我。
ACTS|20|24|我卻不以性命為念，只要走完我的路程，完成我從主耶穌所領受的職分，為上帝恩典的福音作見證。
ACTS|20|25|「我素常在你們中間到處傳講上帝的國；現在我知道，你們眾人以後不會再見到我的面了。
ACTS|20|26|所以我今日向你們作證，你們中間無論何人死亡，罪不在我。
ACTS|20|27|因為上帝一切的旨意，我並沒有退縮不傳給你們的。
ACTS|20|28|聖靈立你們作全群的監督，你們就當為自己謹慎，也為全群謹慎，牧養上帝 的教會，就是他用自己血所買來的 。
ACTS|20|29|我知道，在我離開以後必有兇暴的豺狼進入你們中間，不顧惜羊群。
ACTS|20|30|就是你們中間也必有人起來，說悖謬的話，要引誘門徒跟從他們。
ACTS|20|31|所以你們要警醒，記念我三年之久，晝夜不斷地流淚勸戒你們各人。
ACTS|20|32|現在我把你們交託給上帝和他恩惠的道；這道能建立你們，使你們和一切成聖的人同得基業。
ACTS|20|33|我未曾貪圖一個人的金、銀或衣服。
ACTS|20|34|你們自己知道，我靠兩隻手工作來供給我和同工的需用。
ACTS|20|35|我凡事給你們作榜樣，叫你們知道應當這樣勞苦，扶助軟弱的人，又當記念主耶穌的話，說：『施比受更為有福。』」
ACTS|20|36|保羅 說完了這些話，就和大家跪下來禱告。
ACTS|20|37|眾人痛哭，抱著 保羅 的頸項跟他親吻。
ACTS|20|38|叫他們最傷心的，就是他說「以後不會再見到我的面」那句話。於是他們送他上船去了。
ACTS|21|1|我們離別了眾人，就開船直航到 哥士 ，第二天到了 羅底 ，又從那裏到 帕大喇 。
ACTS|21|2|我們遇見一隻船要往 腓尼基 去，就上船起航。
ACTS|21|3|我們望見 塞浦路斯 ，就從南邊行過，往 敘利亞 去，在 推羅 上岸，因為船要在那裏卸貨。
ACTS|21|4|我們在那裏找到了一些門徒，就住了七天。他們藉著聖靈的感動，告訴 保羅 不要上 耶路撒冷 去。
ACTS|21|5|幾天之後，我們又出發前行。他們眾人同妻子兒女都送我們到城外，我們都跪在灘上禱告，彼此辭別。
ACTS|21|6|我們上了船，他們就回家去了。
ACTS|21|7|我們從 推羅 行完航程，來到了 多利買 ，問候那裏的弟兄，和他們同住了一天。
ACTS|21|8|第二天，我們離開那裏，來到 凱撒利亞 ，就進了傳福音的 腓利 家裏，和他同住；他是那七個執事裏的一個。
ACTS|21|9|他有四個女兒，都是未出嫁的，都會說預言。
ACTS|21|10|我們在那裏多住了好幾天，有一個先知，名叫 亞迦布 ，從 猶太 下來。
ACTS|21|11|他到了我們這裏，就拿 保羅 的腰帶，捆上自己的手腳，說：「聖靈這樣說：『 猶太 人在 耶路撒冷 要如此捆綁這腰帶的主人，把他交在外邦人手裏。』」
ACTS|21|12|我們聽見這些話，就跟當地的人苦勸 保羅 不要上 耶路撒冷 去。
ACTS|21|13|於是 保羅 回答：「你們為甚麼這樣痛哭，使我心碎呢？我為主耶穌的名，不但被人捆綁，就是死在 耶路撒冷 也是願意的。」
ACTS|21|14|既然 保羅 不聽勸，我們就住了口，只說：「願主的旨意成就。」
ACTS|21|15|過了這幾天，我們收拾行李上 耶路撒冷 去。
ACTS|21|16|有 凱撒利亞 的幾個門徒和我們同去，帶我們到一個早期的門徒 塞浦路斯 人 拿孫 的家裏，請我們與他同住。
ACTS|21|17|我們到了 耶路撒冷 ，弟兄們歡歡喜喜地接待我們。
ACTS|21|18|第二天， 保羅 同我們去見 雅各 ；所有的長老也都在場。
ACTS|21|19|保羅 向他們問安，然後將上帝用他在外邦人中所做的事奉，一一述說了。
ACTS|21|20|他們聽見了，就歸榮耀給上帝，對 保羅 說：「弟兄，你看 猶太 人中有數以萬計的信徒，而他們都是熱心於律法的人。
ACTS|21|21|他們曾聽見人說，你教導所有在外邦的 猶太 人離棄 摩西 ，對他們說，不要給孩子行割禮，也不要遵守規矩。
ACTS|21|22|眾人必聽見你來了，這可怎麼辦呢？
ACTS|21|23|你就照著我們的話做吧！我們這裏有四個人，都有願在身。
ACTS|21|24|你帶他們去，與他們一同行潔淨的禮，替他們繳納規費，讓他們得以剃頭。這樣，眾人就會知道，先前所聽見關於你的事都是假的；而且也知道，你自己為人循規蹈矩，遵行律法。
ACTS|21|25|至於信主的外邦人， 我們已經根據我們的決議寫信，叫他們要禁戒偶像所玷污的東西、血和勒死的牲畜，禁戒淫亂。」
ACTS|21|26|於是 保羅 帶著那四個人，第二天與他們一同行了潔淨禮，進了聖殿，報告潔淨期滿的日子，等候祭司為他們各人獻上祭物。
ACTS|21|27|那七日將完，從 亞細亞 來的 猶太 人看見 保羅 在聖殿裏，就煽動所有的群眾，下手拿住他，
ACTS|21|28|喊著：「 以色列 人哪，來幫忙！這就是在各處教導眾人糟蹋我們百姓、律法和這地方的人。不但如此，他還帶了 希臘 人進聖殿，污穢了這聖地。」
ACTS|21|29|這話是因他們曾看見 以弗所 人 特羅非摩 跟 保羅 一起在城裏，以為 保羅 帶他進了聖殿。
ACTS|21|30|於是全城都騷動，百姓一齊跑來，拿住 保羅 ，拉他出聖殿，殿門立刻都關了。
ACTS|21|31|他們正想要殺他，有人報信給營裏的千夫長，說 耶路撒冷 全城都亂了。
ACTS|21|32|千夫長立刻帶著士兵和幾個百夫長，跑下去到他們那裏。他們見了千夫長和士兵，就停下來不打 保羅 。
ACTS|21|33|於是千夫長上前拿住他，吩咐用兩條鐵鏈捆鎖，又問他是甚麼人，做了甚麼事。
ACTS|21|34|群眾中有的喊這個，有的喊那個；因為這樣亂嚷，千夫長無法知道實情，就下令將 保羅 帶進營樓去。
ACTS|21|35|保羅 一走上臺階，群眾擠得兇猛，士兵只得將 保羅 抬起來。
ACTS|21|36|一群人跟在後面，喊著：「除掉他！」
ACTS|21|37|保羅 快要被帶進營樓時，對千夫長說：「我可以對你說句話嗎？」千夫長說：「你懂得 希臘 話嗎？
ACTS|21|38|那你就不是從前作亂、帶領四千兇徒往曠野去的那 埃及 人了。」
ACTS|21|39|保羅 說：「我本是 猶太 人，生在 基利家 的 大數 ，並不是無名小城的公民。求你准我對百姓說話。」
ACTS|21|40|千夫長准了。 保羅 就站在臺階上，向百姓做了個手勢，要他們靜下來， 保羅 就用 希伯來 話對他們說：
ACTS|22|1|「諸位父老弟兄，請聽我現在對你們的申辯。」
ACTS|22|2|他們聽 保羅 說的是 希伯來 話，就更加安靜了。
ACTS|22|3|保羅 說：「我原是 猶太 人，生在 基利家 的 大數 ，但在這城裏長大，在 迦瑪列 門下按著我們祖宗嚴緊的律法受教，熱心事奉上帝，就如你們大家今日一樣。
ACTS|22|4|我也曾迫害信奉這道路的人，置他們於死地，無論男女都捆綁，關在監裏。
ACTS|22|5|這是大祭司和議會的眾長老都可以給我作證的。我又從他們那裏領了致弟兄們的書信，往 大馬士革 去，要把在那裏的信徒綁起來，帶到 耶路撒冷 受刑。」
ACTS|22|6|「當我走近 大馬士革 的時候，約在中午，忽然有一道大光從天上下來，照射在我周圍。
ACTS|22|7|我就仆倒在地，聽見有聲音對我說：『 掃羅 ！ 掃羅 ！你為甚麼迫害我？』
ACTS|22|8|我回答：『主啊！你是誰？』他對我說：『我就是你所迫害的 拿撒勒 人耶穌。』
ACTS|22|9|跟我一起的人看見了那光，卻沒有聽見那位對我說話的聲音。
ACTS|22|10|我說：『主啊，我該做甚麼？』主說：『起來，進 大馬士革 去，在那裏有人會把指派你做的一切事告訴你。』
ACTS|22|11|我因那光的閃耀不能看見，跟我一起的人就拉著我的手進了 大馬士革 。
ACTS|22|12|「那裏有一個人，名叫 亞拿尼亞 ，按著律法是虔誠人，為所有住在那裏的 猶太 人所稱讚。
ACTS|22|13|他來見我，站在旁邊，對我說：『 掃羅 弟兄，你看見吧！』就在那時，我恢復視覺，看見了他。
ACTS|22|14|他又說：『我們祖宗的上帝揀選了你，讓你明白他的旨意，又看見那義者，聽見他口中所出的聲音。
ACTS|22|15|因為你要將所看見的、所聽見的，對著萬人作他的見證人。
ACTS|22|16|現在你為甚麼耽延呢？起來，受洗，求告他的名，洗去你的罪。』」
ACTS|22|17|「後來，我回到 耶路撒冷 ，在聖殿裏禱告的時候，魂遊象外，
ACTS|22|18|看見主對我說：『你趕緊離開 耶路撒冷 ，越快越好，因為這裏的人不接受你為我作的見證。』
ACTS|22|19|我就說：『主啊，他們都知道，我從前在各會堂裏把信你的人監禁，又鞭打他們。
ACTS|22|20|當你的見證人 司提反 被害流血的時候，我也站在一旁贊同；又為打死他的人看守衣裳。』
ACTS|22|21|主對我說：『你去吧！我要差你到遠方外邦人那裏去。』」
ACTS|22|22|眾人聽他說到這句話，就高聲說：「這樣的人，從地上除掉他吧！他是該死的。」
ACTS|22|23|大家一邊喧嚷一邊摔衣裳，向空中撒灰塵。
ACTS|22|24|千夫長下令把 保羅 帶進營樓，叫人用鞭子拷問他，要知道他們向他這樣喧嚷是甚麼緣故。
ACTS|22|25|他們剛用皮條把他捆上的時候， 保羅 對站在旁邊的百夫長說：「一個 羅馬 人，又未被定罪，你們就鞭打他是合法的嗎？」
ACTS|22|26|百夫長聽見這話，就去見千夫長，報告說：「你要怎麼辦呢？這個人是 羅馬 人。」
ACTS|22|27|千夫長就來問 保羅 ：「你告訴我，你是 羅馬 人嗎？」 保羅 說：「是。」
ACTS|22|28|千夫長回答：「我用了許多銀子才得到 羅馬 公民的身份。」 保羅 說：「我生來就是。」
ACTS|22|29|於是那些要拷問 保羅 的人立刻離開他走了。千夫長一知道他是 羅馬 人，又因為曾捆綁了他，也害怕起來。
ACTS|22|30|第二天，千夫長為要知道 猶太 人控告 保羅 的實情，就解開他，下令祭司長們和全議會的人都聚集，然後將 保羅 帶下來，叫他站在他們面前。
ACTS|23|1|保羅 定睛看著議會的人，說：「諸位弟兄，我在上帝面前，行事為人都是憑著清白的良心，直到今日。」
ACTS|23|2|亞拿尼亞 大祭司就吩咐旁邊站著的人打他的嘴。
ACTS|23|3|這時， 保羅 對他說：「你這粉飾的牆，上帝要打你！你坐堂是要按律法審問我，你竟違背律法，命令人打我嗎？」
ACTS|23|4|站在旁邊的人說：「你竟敢辱罵上帝的大祭司嗎？」
ACTS|23|5|保羅 說：「弟兄們，我不知道他是大祭司；因為經上記著：『不可毀謗你百姓的官長。』」
ACTS|23|6|保羅 看出他們一部分是撒都該人，一部分是法利賽人，就在議會中喊著：「諸位弟兄，我是法利賽人，也是法利賽人的子孫。我現在受審問是為有關死人復活的盼望。」
ACTS|23|7|說了這話，法利賽人和撒都該人爭論起來，會眾分為兩派。
ACTS|23|8|因為撒都該人一方面說沒有復活，另一方面沒有天使和鬼魂；法利賽人卻承認兩方面都有。
ACTS|23|9|於是大大地爭吵起來；有幾個法利賽派的文士站起來爭辯說：「我們看不出這人有甚麼錯處；說不定有鬼魂或者天使對他說過話呢！」
ACTS|23|10|那時爭辯越來越大，千夫長恐怕 保羅 被他們扯碎了，就命令士兵下去，把他從眾人當中搶出來，帶進營樓去。
ACTS|23|11|當夜，主站在 保羅 旁邊，說：「放心吧！你怎樣在 耶路撒冷 為我作見證，也必怎樣在 羅馬 為我作見證。」
ACTS|23|12|到了天亮， 猶太 人同謀起誓，說「若不先殺 保羅 就不吃不喝」。
ACTS|23|13|參與這陰謀的有四十多人。
ACTS|23|14|他們來見祭司長和長老，說：「我們已經發了重誓，若不先殺 保羅 就甚麼也不吃。
ACTS|23|15|現在你們和議會要通知千夫長，叫他把 保羅 帶到你們這裏來，假裝要詳細調查他的事；我們已經預備好，在他來到這裏以前就殺掉他。」
ACTS|23|16|保羅 的外甥聽見他們設下埋伏，就來到營樓裏告訴 保羅 。
ACTS|23|17|保羅 請一個百夫長來，說：「你領這青年去見千夫長，他有事告訴他。」
ACTS|23|18|於是百夫長把他領去見千夫長，說：「被囚的 保羅 請我到他那裏，求我領這青年來見你；他有事告訴你。」
ACTS|23|19|千夫長就拉著他的手，走到一旁，私下問他：「你有甚麼事告訴我呢？」
ACTS|23|20|他說：「 猶太 人已經約定，要求你明天把 保羅 帶到議會去，假裝要詳細查問他的事。
ACTS|23|21|你切不要隨從他們，因為他們有四十多人埋伏，已經起誓，若不先殺掉 保羅 就不吃不喝。現在都預備好了，只等你的允准。」
ACTS|23|22|於是千夫長打發那青年走，囑咐他：「不要告訴人，你已將這些事報告我了。」
ACTS|23|23|於是，千夫長叫了兩個百夫長來，說：「預備步兵二百、騎兵七十、長槍手二百，今夜九點往 凱撒利亞 去；
ACTS|23|24|也要預備牲口讓 保羅 騎上，護送到 腓力斯 總督那裏去。」
ACTS|23|25|千夫長又寫了公文，大略說：
ACTS|23|26|「 克勞第．呂西亞 向 腓力斯 總督大人請安。
ACTS|23|27|這個人被 猶太 人拿住，快被殺害時，我得知他是 羅馬 人，就帶士兵下去，把他救了出來。
ACTS|23|28|因為我要知道他們告他的罪狀，就帶他下到他們的議會去。
ACTS|23|29|我查知他被告發是因他們律法上的爭論，並沒有甚麼該死或該監禁的罪名。
ACTS|23|30|後來有人把要害他的計謀告訴我，我立刻把他解到你那裏去，又命令告他的人在你面前告他。 」
ACTS|23|31|於是士兵照所命令他們的，連夜把 保羅 帶到 安提帕底 。
ACTS|23|32|第二天，由騎兵護送 保羅 ，他們就回營樓去。
ACTS|23|33|騎兵來到 凱撒利亞 ，把公文呈給總督，就叫 保羅 站在他面前。
ACTS|23|34|總督讀了公文，問 保羅 是哪一省的人；一知道他是 基利家 人，
ACTS|23|35|就說：「等告你的人來到，我才詳細聽你。」於是他命令把 保羅 拘留在 希律 的衙門裏。
ACTS|24|1|過了五天， 亞拿尼亞 大祭司、幾個長老和一個叫 帖土羅 的律師下來，向總督控告 保羅 。
ACTS|24|2|保羅 一被傳來， 帖土羅 就開始控告他，說：「 腓力斯 大人，我們因你得以享受國泰民安，並且這一國的弊病，因著你的遠見得以改革。
ACTS|24|3|我們隨時隨地都滿心感激不盡。
ACTS|24|4|為了不敢耽擱你太久，我只求你寬容一下，聽我們說幾句話。
ACTS|24|5|我們看這個人如同瘟疫一般，是鼓動普天下所有的 猶太 人作亂的人，又是 拿撒勒 教派裏的一個頭目。
ACTS|24|6|他甚至連聖殿也要污穢，我們就把他捉拿了。
ACTS|24|7|
ACTS|24|8|你自己審問他，就可以知道我們所控告他的一切事了。」
ACTS|24|9|眾 猶太 人也隨著控告他，說：「這些事情確是這樣。」
ACTS|24|10|總督示意叫 保羅 說話， 保羅 就回答：「我知道你在本國作法官多年，所以我樂意為自己申辯。
ACTS|24|11|你查問就可以知道，從我上 耶路撒冷 去禮拜到今日不過十二天。
ACTS|24|12|他們並沒有看見我在聖殿裏跟人辯論，或在會堂裏、在城裏煽動群眾。
ACTS|24|13|也不能對你證實他們現在所控告我的事。
ACTS|24|14|但有一件事我向你承認，就是我正按著他們所稱為異端的道事奉我祖宗的上帝，又信合乎律法和先知書上所記載的一切。
ACTS|24|15|我對上帝存著這些人自己也接受的盼望，就是義人和不義的人都要復活。
ACTS|24|16|因此，我勉勵自己，對上帝對人，時常存著無虧的良心。
ACTS|24|17|過了幾年，我帶著賙濟本國的捐項和供物上去。
ACTS|24|18|正獻的時候，他們看見我在聖殿裏已經潔淨了，並沒有聚眾，也沒有吵嚷，
ACTS|24|19|惟有幾個從 亞細亞 來的 猶太 人—他們若有控告我的事，應當到你面前來告我。
ACTS|24|20|不然，讓這些人自己說，他們看出我站在議會前的時間，有甚麼不對的地方。
ACTS|24|21|縱然有，也不過是為了一句話，就是我站在他們中間喊說：『我今日在你們面前受審，是為了死人復活。』」
ACTS|24|22|腓力斯 本是詳細認識這道，就拖延他們，說：「且等 呂西亞 千夫長下來，我再審判你們的案。」
ACTS|24|23|於是他下令百夫長看守 保羅 ，要從寬待他，不可攔阻他的親友來供給他。
ACTS|24|24|過了幾天， 腓力斯 和他夫人 猶太 女子 土西拉 一同來到，就叫 保羅 來，聽他講論信基督耶穌的事。
ACTS|24|25|保羅 講論公義、節制和將來的審判， 腓力斯 害怕起來，就回答：「你暫且去吧！等我有機會時再來叫你。」
ACTS|24|26|腓力斯 又指望 保羅 送他銀錢，所以屢次叫他來，和他談論。
ACTS|24|27|過了兩年， 波求．非斯都 接了 腓力斯 的任； 腓力斯 要討 猶太 人的喜歡，就把 保羅 留在監裏。
ACTS|25|1|非斯都 到省裏上任，過了三天，就從 凱撒利亞 上 耶路撒冷 去。
ACTS|25|2|祭司長和 猶太 人的領袖向他控告 保羅 ；又央求他，
ACTS|25|3|向他求情要對付 保羅 ，把他提到 耶路撒冷 來，他們要在路上埋伏殺害他。
ACTS|25|4|非斯都 就回答：「 保羅 押在 凱撒利亞 ，我自己快要往那裏去。」
ACTS|25|5|他又說：「所以，你們中間有權的人與我一同下去，那人若有甚麼不是，就讓他們控告他。」
ACTS|25|6|非斯都 在他們那裏住了不超過八天或十天，就下 凱撒利亞 去；第二天開庭，下令把 保羅 提上來。
ACTS|25|7|保羅 來了，那些從 耶路撒冷 下來的 猶太 人周圍站著，提出許多嚴重而不能證實的事控告他。
ACTS|25|8|保羅 申辯說：「無論 猶太 人的律法，或是聖殿，或是凱撒，我都沒有干犯。」
ACTS|25|9|但 非斯都 要討 猶太 人的喜歡，就回答 保羅 說：「你願意上 耶路撒冷 去，在那裏為這些事受我的審判嗎？」
ACTS|25|10|保羅 說：「我現在站在凱撒的審判臺前，這就是我應當受審的地方。我並沒有對 猶太 人做過甚麼不對的事，這也是你明明知道的。
ACTS|25|11|我若做了不對的事，犯了甚麼該死的罪，就是死我也不辭。他們所控告我的事若都不實，就沒有人能把我交給他們。我要向凱撒上訴。」
ACTS|25|12|非斯都 和議會商量了，就回答：「既然你要向凱撒上訴，你就到凱撒那裏去吧。」
ACTS|25|13|過了些日子， 亞基帕 王和 百妮基 來到 凱撒利亞 ，拜訪 非斯都 。
ACTS|25|14|他們在那裏住了好些日子， 非斯都 將 保羅 的案件向王陳述，說：「這裏有一個人，是 腓力斯 留在監裏的。
ACTS|25|15|我在 耶路撒冷 的時候，祭司長和 猶太 的長老把他的事稟報了，要求定他的罪。
ACTS|25|16|我回覆他們，無論甚麼人，被告還沒有和原告當面對質，沒有機會為所控告的事申辯，就先定他罪的，這不是 羅馬 人的規矩。
ACTS|25|17|及至他們都來到這裏，我沒有耽誤，第二天就開庭，下令把那人提上來。
ACTS|25|18|控告他的人站起來告他，所控告的並沒有任何我所預料的那等惡 事。
ACTS|25|19|不過，有幾樣辯論是有關他們自己敬鬼神的事，以及一個名叫耶穌的人，他已經死了， 保羅 卻說他是活著的。
ACTS|25|20|我對這些事不知該怎樣處理，所以問他是否願意上 耶路撒冷 去，在那裏為這些事接受審判。
ACTS|25|21|但 保羅 要求我留下他，要聽皇上判斷，我就下令把他留下，等我解他到凱撒那裏去。」
ACTS|25|22|亞基帕 對 非斯都 說：「我也願意親自聽聽這個人。」 非斯都 說：「明天你就可以聽他。」
ACTS|25|23|第二天， 亞基帕 和 百妮基 大張旗鼓而來，與眾千夫長和城裏的顯要進了大廳。 非斯都 一聲令下，就有人將 保羅 帶進來。
ACTS|25|24|非斯都 說：「 亞基帕 王和在這裏的諸位，你們看這個人，他就是所有在 耶路撒冷 和這裏的 猶太 人曾向我懇求呼叫，說不可容他再活著的。
ACTS|25|25|但我查明他並沒有犯甚麼該死的罪，並且他自己也已向皇帝上訴了，所以我決定把他解去。
ACTS|25|26|論到這個人，我沒有確實的事可以奏明主上。因此，我帶他到你們面前，尤其到你 亞基帕 王面前，為要在查問之後有所呈奏。
ACTS|25|27|因為據我看，解送囚犯而不指明他的罪狀是不合理的。」
ACTS|26|1|亞基帕 對 保羅 說：「准你為自己申訴。」於是 保羅 伸手辯護說：
ACTS|26|2|「 亞基帕 王啊， 猶太 人所控告我的一切事，今日得以在你面前辯護，實為萬幸。
ACTS|26|3|更慶幸的是你熟悉 猶太 人的規矩和他們的爭論；所以，求你耐心聽我。
ACTS|26|4|「我自幼為人如何，從起初在本國的同胞中，以及在 耶路撒冷 ，所有的 猶太 人都知道。
ACTS|26|5|他們若肯作見證，就知道我從起初是按著我們教中最嚴緊的教門作了法利賽人。
ACTS|26|6|現在我站在這裏受審，是為了對上帝向我們祖宗的應許存著盼望。
ACTS|26|7|這應許，我們十二個支派，晝夜切切地事奉上帝，都指望得著。王啊，我正是因這指望被 猶太 人控告。
ACTS|26|8|上帝使死人復活，你們為甚麼判斷為不可信呢？
ACTS|26|9|「從前我自己認為必須竭力反對 拿撒勒 人耶穌的名，
ACTS|26|10|我在 耶路撒冷 也曾這樣做過；我不但從祭司長得了權柄，把許多聖徒收在監裏，而且他們被殺，我也表示 贊成。
ACTS|26|11|在各會堂，我屢次用刑強迫他們說褻瀆的話，我非常厭惡他們，甚至追逼他們，直到外邦的城鎮。」
ACTS|26|12|「那時，我帶著祭司長的權柄和命令往 大馬士革 去。
ACTS|26|13|王啊！我在路上，中午的時候，看見從天上有一道光，比太陽還亮，四面照射著我和跟我同行的人。
ACTS|26|14|我們都仆倒在地，我就聽見有聲音用 希伯來 話對我說：『 掃羅 ！ 掃羅 ！你為甚麼迫害我？你用腳踢刺棒是自找苦吃的！』
ACTS|26|15|我說：『主啊，你是誰？』主說：『我就是你所迫害的耶穌。
ACTS|26|16|起來，站著，我向你顯現的目的是要派你作僕役，為你所看見我 的事，和我將要指示你的事作見證人。
ACTS|26|17|我也要救你脫離百姓和外邦人的手。我差你到他們那裏去，
ACTS|26|18|要開他們的眼睛，使他們從黑暗中轉向光明，從撒但權下歸向上帝；使他們因信我而得蒙赦罪，和一切成聖的人同得基業。』」
ACTS|26|19|「因此， 亞基帕 王啊！我沒有違背那從天上來的異象；
ACTS|26|20|我先在 大馬士革 ，後在 耶路撒冷 和 猶太 全地，以及外邦，勸勉他們應當悔改歸向上帝，行事與悔改的心相稱。
ACTS|26|21|為這緣故， 猶太 人在聖殿裏拿住我，想要殺我。
ACTS|26|22|然而，我蒙上帝的幫助，直到今日還站立得穩，向尊貴的和卑微的作見證。我所講的，並不外乎眾先知和 摩西 所說將來必成的事，
ACTS|26|23|就是基督必須受害，並且首先從死人中復活，把亮光傳給 猶太 人和外邦人。」
ACTS|26|24|保羅 這樣申訴時， 非斯都 大聲說：「 保羅 ，你瘋了！你的學問太大，反使你瘋了！」
ACTS|26|25|保羅 說：「 非斯都 大人，我不是瘋了，我說的乃是真實和清醒的話。
ACTS|26|26|王也知道這些事，所以對王大膽直言，我深信這些事沒有一件能向王隱瞞的，因為都不是在背地裏做的。
ACTS|26|27|亞基帕 王啊，你信先知嗎？我知道你是信的。」
ACTS|26|28|亞基帕 對 保羅 說：「你想稍微勸一勸就能說服我作基督徒了嗎？」
ACTS|26|29|保羅 說：「無論少勸還是多勸，我向上帝所求的，不但你一個人，就是今天所有聽我說話的人都要像我一樣，只是不要有這些鎖鏈。」
ACTS|26|30|於是，王和總督以及 百妮基 跟同坐的人都站起來，
ACTS|26|31|退到裏面，彼此談論說：「這個人並沒有犯甚麼該死該監禁的罪。」
ACTS|26|32|亞基帕 對 非斯都 說：「這人若沒有向凱撒上訴，早就被釋放了。」
ACTS|27|1|既然 非斯都 決定要我們坐船往 意大利 去，就將 保羅 和別的囚犯交給御營裏的一個名叫 猶流 的百夫長。
ACTS|27|2|有一隻 亞大米田 的船要開往 亞細亞 沿海一帶地方去，我們上了那船，就起航了；有 馬其頓 的 帖撒羅尼迦 人 亞里達古 和我們同去。
ACTS|27|3|第二天，我們到了 西頓 。 猶流 寬待 保羅 ，准他往朋友那裏去，受他們的照應。
ACTS|27|4|我們又從那裏開船，因為遇到逆風，就貼著 塞浦路斯 的背風岸航行，
ACTS|27|5|渡過了 基利家 、 旁非利亞 一帶的海面，就到了 呂家 的 每拉 。
ACTS|27|6|在那裏，百夫長找到一隻 亞歷山大 的船要往 意大利 去，就叫我們上了那船。
ACTS|27|7|一連多日，船行得很慢，我們好不容易才來到 革尼土 的對面；又因被風攔阻，我們就貼著 克里特 島背風岸，從 撒摩尼 對面航行。
ACTS|27|8|我們沿岸前進，十分艱難，來到一個名叫 佳澳 的地方，離那裏不遠有 拉西亞城 。
ACTS|27|9|航行的日子久了，已經過了禁食的節期，行船又危險， 保羅 就建議，
ACTS|27|10|對眾人說：「諸位，我看這次航行，不但貨物和船要受損傷，大遭破壞，連我們的性命也難保。」
ACTS|27|11|但百夫長信從船長和船主，不信 保羅 所說的。
ACTS|27|12|且因在這港口不適宜過冬，船上大多數的人都主張開船離開這地方，或者能到 非尼基 去過冬。 非尼基 是 克里特 的一個港口，一面朝西南，一面朝西北。
ACTS|27|13|當南風微微吹起時，他們以為對目的地已有了把握，就起錨，貼近 克里特 開去。
ACTS|27|14|過了不久，有一股叫「友拉革羅」的東北巨風從島上撲來，
ACTS|27|15|船被風抓住，無法頂風航行，我們只好任它漂流。
ACTS|27|16|我們貼著一個叫 高大 的小島的背風岸急航，好不容易才保住了救生艇。
ACTS|27|17|既然把救生艇拉上來，他們就用纜索捆綁船底，又恐怕在 賽耳底 淺灘上擱淺，就落了篷，任船漂流。
ACTS|27|18|我們被風浪逼得很急，第二天眾人就把貨物拋在海裏。
ACTS|27|19|第三天，他們又親手把船上的器具拋棄了。
ACTS|27|20|許多天都沒有看到太陽和星辰，又有狂風大浪催逼，我們獲救的指望都放棄了。
ACTS|27|21|眾人已有好幾天沒有吃東西， 保羅 就出來站在他們中間，說：「諸位，你們本該聽我的話不離開 克里特 島，就不致遭到這樣的損失和破壞。
ACTS|27|22|現在我勸你們放心，除了損失這條船，你們中間沒有一人會喪失性命。
ACTS|27|23|因為昨夜，我所屬所事奉的上帝的使者站在我旁邊，
ACTS|27|24|說：『 保羅 ，不要害怕，你必定站在凱撒面前；並且上帝已把安全賜給與你同船的人了。』
ACTS|27|25|所以，諸位可以放心，我信上帝怎樣對我說，事情也要怎樣成就；
ACTS|27|26|只是我們必須在一個島上擱淺。」
ACTS|27|27|到了第十四天夜間，船在 亞得里亞海 漂來漂去。約在半夜，水手以為漸近旱地，
ACTS|27|28|就去探測深淺，探得有十二丈 ；稍往前行，又探深淺，探得有九丈。
ACTS|27|29|恐怕我們撞到礁石，他們就從船尾拋下四個錨，盼望天亮。
ACTS|27|30|水手想棄船逃走，把救生艇縋下海裏，假裝要從船頭拋錨的樣子。
ACTS|27|31|保羅 對百夫長和士兵說：「這些人若不留在船上，你們就不能獲救。」
ACTS|27|32|於是士兵砍斷救生艇的繩子，由它漂去。
ACTS|27|33|天快亮的時候， 保羅 勸眾人都用餐，說：「你們一直捱餓等候，不吃甚麼，已經十四天了。
ACTS|27|34|所以我勸你們吃點東西，這是關乎你們獲救的，因為你們各人連一根頭髮也不至於掉落。」
ACTS|27|35|保羅 說了這話，就拿起餅來，在眾人面前祝謝了上帝，然後擘開來吃。
ACTS|27|36|於是他們都放心，就吃了。
ACTS|27|37|我們在船上的共有二百七十六個人。
ACTS|27|38|他們吃飽了，為要使船輕一點，就把船上的麥子拋到海裏。
ACTS|27|39|天亮的時候，他們不認得那地方，只見一個有岸可登的海灣，就想法子看能不能把船靠岸。
ACTS|27|40|於是他們砍斷纜索，把錨丟到海裏，同時也鬆開舵繩，拉起頭篷，順風向著岸行去。
ACTS|27|41|但碰到兩水夾流的地方，就擱了淺，船頭膠住不動，船尾被浪的猛力衝壞了 。
ACTS|27|42|士兵的意思要把囚犯都殺了，免得有游水脫逃的。
ACTS|27|43|但百夫長要救 保羅 ，不准他們任意而行，就吩咐會游水的，跳下水去，先上岸；
ACTS|27|44|其餘的人則用板子或船的碎片上岸。這樣，眾人都獲救，上了岸。
ACTS|28|1|我們既已獲救，才知道那島名叫 馬耳他 。
ACTS|28|2|當地人非常友善地接待我們；因為正在下雨，天氣又冷，他們就生了火歡迎我們眾人。
ACTS|28|3|那時， 保羅 拾起一捆柴，放在火中，有一條毒蛇，因為熱的緣故鑽了出來，纏住他的手。
ACTS|28|4|當地的人看見那毒蛇懸在他手上，就彼此說：「這人必是個兇手，雖然他從海裏獲救，天理仍不容他活著。」
ACTS|28|5|保羅 竟把那毒蛇甩在火裏，並沒有受傷。
ACTS|28|6|當地的人想他快要腫起來，或是忽然倒下死了，但等了好久，見他沒有甚麼異樣，就轉念說他是個神明。
ACTS|28|7|離那地方不遠有一些田產，是島長 部百流 的。他接納我們，盡情款待了我們三日。
ACTS|28|8|當時， 部百流 的父親臥病不起，患了熱病和痢疾。 保羅 進去見他，為他禱告按手，治好了他。
ACTS|28|9|從此，島上其餘的病人也都來，得了醫治。
ACTS|28|10|他們又多方面尊敬我們，到了開船的時候，又把我們所需用的東西送到船上。
ACTS|28|11|過了三個月，我們上了 亞歷山大 的船起航。這船以「 宙斯 雙子」為記，是在那海島過冬的。
ACTS|28|12|我們到了 敘拉古 ，停泊了三日；
ACTS|28|13|又從那裏起錨開船， 來到 利基翁 。過了一天，起了南風，第二天就來到 部丟利 。
ACTS|28|14|我們在那裏遇見一些弟兄，他們請我們同住了七天。就這樣，我們來到 羅馬 。
ACTS|28|15|那裏的弟兄們一聽見我們的消息，就到 亞比烏 市和 三館 來迎接我們。 保羅 見了他們，就感謝上帝，越發壯膽。
ACTS|28|16|我們進了 羅馬城 ， 保羅 蒙准和那個看守他的兵另住在一處。
ACTS|28|17|過了三天， 保羅 請當地 猶太 人的領袖來。他們來了， 保羅 對他們說：「諸位弟兄，雖然我沒有做甚麼事干犯本國的百姓和我們祖宗的規矩，卻在 耶路撒冷 被囚禁，交在 羅馬 人的手裏。
ACTS|28|18|他們審問了我，有意要釋放我，因為在我身上並沒有該死的罪狀。
ACTS|28|19|但 猶太 人反對，我不得已只好上訴於凱撒，並不是有甚麼事要控告我本國的百姓。
ACTS|28|20|為這緣故，我請你們來見我當面談話，我原是為 以色列 人所指望的那位才被這鐵鏈捆綁的。」
ACTS|28|21|他們對他說：「我們並沒有接到從 猶太 寄來有關於你的信，也沒有弟兄到這裏來向我們報告，或說你有甚麼不好的地方。
ACTS|28|22|但我們願意聽聽你的意見，因為我們知道這教門是到處遭人反對的。」
ACTS|28|23|他們和 保羅 約定了日子，就有許多人到他的住處來。 保羅 從早到晚向他們講解這事，為上帝的國作證，並引 摩西 的律法和先知的書勸導他們信從耶穌。
ACTS|28|24|他所說的話，有的信，有的不信。
ACTS|28|25|他們間彼此不合，就分散了；未散以先， 保羅 說了一句話：「聖靈藉 以賽亞 先知向你們祖宗所說的話是對的。
ACTS|28|26|他說： 『你去對這百姓說： 你們聽了又聽，卻不明白； 看了又看，卻看不清。
ACTS|28|27|因為這百姓的心麻木， 耳朵塞著， 眼睛閉著， 免得眼睛看見， 耳朵聽見， 心裏明白，回轉過來， 我會醫治他們。』
ACTS|28|28|所以，你們當知道，上帝這救恩已經傳給外邦人；他們會聽的。」
ACTS|28|29|
ACTS|28|30|保羅 在自己所租的房子裏住了足足兩年。凡來見他的人，他都接待，
ACTS|28|31|放膽傳講上帝的國，並教導主耶穌基督的事，沒有人禁止。
