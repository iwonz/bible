1TIM|1|1|奉我們的救主上帝，和我們的盼望基督耶穌的命令，作基督耶穌使徒的 保羅 ，
1TIM|1|2|寫信給那因信主作我真兒子的 提摩太 。願恩惠、憐憫、平安 從父上帝和我們主基督耶穌歸給你！
1TIM|1|3|我往 馬其頓 去的時候，曾勸你留在 以弗所 ，好囑咐某些人不可傳別的教義，
1TIM|1|4|也不要聽從無稽的傳說和冗長的家譜；這樣的事只會引起爭論，無助於上帝的計劃，這計劃是憑著信才能了解的。
1TIM|1|5|但命令的目的就是愛；這愛是出於清潔的心、無愧的良心和無偽的信心。
1TIM|1|6|有人偏離了這些而轉向空談，
1TIM|1|7|想要作律法教師，卻不明白自己所講的是甚麼，也不知道所主張的是甚麼。
1TIM|1|8|我們知道，只要人善用律法，律法是好的；
1TIM|1|9|因為知道律法不是為義人訂立的，而是為不法和叛逆的，不虔誠和犯罪的，不聖潔和戀世俗的，弒父母和殺人的，
1TIM|1|10|犯淫亂和親男色的，拐賣人口和說謊話的，並起假誓的，或是為任何違背健全教義的事訂立的。
1TIM|1|11|這是按照可稱頌、榮耀之上帝交託我的福音說的。
1TIM|1|12|我感謝那賜給我力量的我們的主基督耶穌，因為他認為我可信任，派我服事他。
1TIM|1|13|我從前是褻瀆、迫害、侮慢上帝的人；然而我還蒙了憐憫，因為我是在不信、不明白的時候做的。
1TIM|1|14|而且我們的主的恩典格外豐盛，使我在基督耶穌裏有信心和愛心。
1TIM|1|15|這話可信，值得完全接受：「基督耶穌到世上來是要拯救罪人」，而在罪人中我是個罪魁。
1TIM|1|16|然而，我蒙了憐憫，好讓基督耶穌在我這罪魁身上顯明他完全的忍耐，給後來信他得永生的人作榜樣。
1TIM|1|17|願尊貴、榮耀歸給永世的君王，那不朽壞、看不見、獨一的上帝，直到永永遠遠。阿們！
1TIM|1|18|我兒 提摩太 啊，我照從前指著你的預言把這命令交託你，使你能藉著這些預言打那美好的仗，
1TIM|1|19|常存信心和無愧的良心。有些人丟棄良心，在信仰上觸了礁；
1TIM|1|20|其中有 許米乃 和 亞歷山大 ，我已經把他們交給撒但，讓他們學會不再褻瀆。
1TIM|2|1|所以，我勸你，首先要為人人祈求、禱告、代求、感謝；
1TIM|2|2|為君王和一切在位的，也要如此，使我們能夠敬虔端正地過平穩寧靜的生活。
1TIM|2|3|這是好的，在我們的救主上帝面前可蒙悅納。
1TIM|2|4|他願意人人得救，並得以認識真理。
1TIM|2|5|因為只有一位上帝， 在上帝和人之間也只有一位中保， 是成為人的基督耶穌。
1TIM|2|6|他獻上自己作人人的贖價； 在適當的時候這事已經證實了。
1TIM|2|7|我為此奉派作傳道，作使徒，在信仰和真理上作外邦人的教師。我說的是真話，不是說謊。
1TIM|2|8|我希望男人舉起聖潔的手隨處禱告，不發怒，不爭論。
1TIM|2|9|我也希望女人以端正、克制和合乎體統的服裝打扮自己，不以編髮、金飾、珍珠和名貴衣裳來打扮。
1TIM|2|10|要有善行，這才與自稱為敬畏上帝的女人相稱。
1TIM|2|11|女人要事事順服地安靜學習。
1TIM|2|12|我不許女人教導，也不許她管轄男人，只要安靜。
1TIM|2|13|因為 亞當 先被造，然後才是 夏娃 ；
1TIM|2|14|亞當 並沒有受騙，而是女人受騙，陷在過犯裏。
1TIM|2|15|然而，女人若持守信心、愛心，又聖潔克制，就必藉著生產而得救。
1TIM|3|1|「若有人想望監督的職分，他是在羨慕一件好事」，這話是可信的。
1TIM|3|2|監督必須無可指責，只作一個婦人的丈夫，有節制、克己、端正，樂意接待外人，善於教導，
1TIM|3|3|不酗酒，不打人；要溫和，不好鬥，不貪財。
1TIM|3|4|要好好管理自己的家，使兒女順服，凡事莊重。
1TIM|3|5|人若不知道管理自己的家，怎能照管上帝的教會呢？
1TIM|3|6|剛信主的，不可作監督，恐怕他自高自大，落在魔鬼所受的懲罰裏。
1TIM|3|7|監督也必須在教外有好名聲，免得被人毀謗，落在魔鬼的羅網裏。
1TIM|3|8|同樣，執事也必須莊重，不一口兩舌，不好酒，不貪不義之財；
1TIM|3|9|要存清白的良心固守信仰的奧祕。
1TIM|3|10|這些人也要先受考驗，若沒有可責之處，才讓他們作執事。
1TIM|3|11|同樣，女執事 也必須莊重，不說閒話，有節制，凡事忠心。
1TIM|3|12|執事只作一個婦人的丈夫，要好好管兒女和自己的家。
1TIM|3|13|因為善於作執事的，為自己得到美好的地位，並且無懼地堅信在基督耶穌裏的信仰。
1TIM|3|14|我希望盡快到你那裏去，所以先把這些事寫給你；
1TIM|3|15|倘若我延誤了，你也可以知道在上帝的家中該怎樣做。這家就是永生上帝的教會，真理的柱石和根基。
1TIM|3|16|敬虔的奧祕是公認為偉大的： 上帝在肉身顯現， 被聖靈稱義， 被天使看見， 被傳於外邦， 被世人信服， 被接在榮耀裏。
1TIM|4|1|聖靈明說，在末後的時期必有人離棄信仰，去聽信那誘惑人的邪靈和鬼魔的教訓。
1TIM|4|2|這是出於撒謊者的假冒；這些人的良心如同被熱鐵烙了一般。
1TIM|4|3|他們禁止嫁娶，又禁戒食物—就是上帝所造、讓那信而明白真理的人存感謝的心領受的。
1TIM|4|4|上帝所造之物樣樣都是好的，若存感謝的心領受，沒有一樣是不可吃的，
1TIM|4|5|都因上帝的話和人的祈禱而成為聖潔了。
1TIM|4|6|你若把這些事提醒弟兄們，就是基督耶穌的好執事，在信仰的話語和你向來所服從的正確教義上得到了栽培。
1TIM|4|7|要棄絕那世俗的言語和老婦的無稽傳說。要在敬虔上操練自己：
1TIM|4|8|因操練身體有些益處；但敬虔在各方面都有益，它有現今和未來的生命的應許。
1TIM|4|9|這話可信，值得完全接受。
1TIM|4|10|我們勞苦，努力 正是為此，因為我們的指望在乎永生的上帝。他是人人的救主，更是信徒的救主。
1TIM|4|11|你要囑咐和教導這些事。
1TIM|4|12|不可叫人小看你年輕，總要在言語、行為、愛心、信心、清潔上，都作信徒的榜樣。
1TIM|4|13|要以宣讀聖經，勸勉，教導為念，直等到我來。
1TIM|4|14|不要忽略你所得的恩賜，就是從前藉著預言、在眾長老按手的時候賜給你的。
1TIM|4|15|這些事你要殷勤去做，並要在這些事上專心，讓眾人看出你的長進來。
1TIM|4|16|要謹慎自己和自己的教導，要在這些事上恆心，因為這樣做，既能救自己，又能救聽你的人。
1TIM|5|1|不可嚴責老年人，要勸他如同父親。要待年輕人如同弟兄，
1TIM|5|2|年老婦女如同母親。要清清潔潔地待年輕婦女如同姊妹。
1TIM|5|3|要尊敬真正守寡的婦人。
1TIM|5|4|寡婦若有兒女，或有孫兒女，要讓兒孫先在自己家中學習行孝，報答親恩，因為這在上帝面前是可蒙悅納的。
1TIM|5|5|獨居無靠的真寡婦只仰賴上帝，晝夜不住地祈求禱告。
1TIM|5|6|但好宴樂的寡婦活著也算是死了。
1TIM|5|7|這些事，你要囑咐她們，讓她們無可指責。
1TIM|5|8|若有人不照顧親屬，尤其是自己家裏的人，就是背棄信仰，還不如不信的人。
1TIM|5|9|寡婦登記，年齡必須在六十歲以上，只作一個丈夫的妻子，
1TIM|5|10|又有行善的名聲，就如養育兒女，收留外人，洗聖徒的腳，救濟遭難的人，竭力行各樣善事。
1TIM|5|11|至於年輕的寡婦，你要拒絕登記，因為她們情慾衝動、背棄基督的時候，就想嫁人，
1TIM|5|12|她們因廢棄了當初所許的願而被定罪。
1TIM|5|13|同時，她們又學了懶惰，習慣於挨家閒逛；不但懶惰，而且說長道短，好管閒事，說些不該說的話。
1TIM|5|14|所以，我希望年輕的寡婦嫁人，生養兒女，治理家務，不讓敵人有辱罵的把柄，
1TIM|5|15|因為已經有一些人轉去隨從撒但了。
1TIM|5|16|信主的婦女若有親戚是寡婦，要救濟她們，不可拖累教會，好使教會能救濟真正無助的寡婦。
1TIM|5|17|善於督導教會的長老，尤其是勤勞講道教導人的，應該得到加倍的敬奉。
1TIM|5|18|因為經上說：「牛在踹穀的時候，不可籠住牠的嘴」；又說：「工人得工資是應當的。」
1TIM|5|19|有控告長老的案件，非有兩三個證人就不要受理。
1TIM|5|20|繼續犯罪的人，要在眾人面前責備他，使其餘的人也有所懼怕。
1TIM|5|21|我在上帝、基督耶穌和蒙揀選的天使面前囑咐你要遵守這些話，不可存成見，做事也不可偏心。
1TIM|5|22|不可急於給人行按手禮；也不可在別人的罪上有份，要保守自己純潔。
1TIM|5|23|為了你的胃，又常患病，不要只喝水，要稍微喝點酒。
1TIM|5|24|有些人的罪是明顯的，已先受審判了；有些人的罪是隨後跟著來。
1TIM|5|25|同樣，善行也有明顯的，就是那不明顯的也不能隱藏。
1TIM|6|1|凡負軛作奴隸的，要認為自己的主人配受各樣的尊敬，免得上帝的名和教導被人褻瀆。
1TIM|6|2|奴隸若有信主的主人，不可因他是主內弟兄就輕看他們，更要越發服侍他們，因為得到服侍的益處的正是信徒，是蒙愛的人。 你要教導人和勸勉這些事。
1TIM|6|3|若有人傳別的教義，不符合我們主耶穌基督純正的話語與合乎敬虔的教導，
1TIM|6|4|他是自高自大，一無所知，專好爭辯，擅於舌戰，因而生出嫉妒、紛爭、毀謗、惡意猜疑，
1TIM|6|5|和心術不正與喪失真理的人不停地爭吵，以敬虔為得利的門路。
1TIM|6|6|其實，敬虔加上知足就是大利。
1TIM|6|7|因為我們沒有帶甚麼到世上來， 也不能帶甚麼去；
1TIM|6|8|只要有衣有食， 我們就該知足。
1TIM|6|9|但那些想要發財的人就陷在誘惑、羅網和許多無知有害的慾望中，使人沉淪，以致敗壞和滅亡。
1TIM|6|10|貪財是萬惡之根。有人因貪戀錢財而背離信仰，用許多愁苦把自己刺透了。
1TIM|6|11|但你這屬上帝的人哪，要逃避這些事；要追求公義、敬虔、信心、愛心、忍耐、溫柔。
1TIM|6|12|你要為信仰打那美好的仗；要持定永生，你為此被召，也已經在許多見證人面前作了那美好的見證。
1TIM|6|13|我在那賜生命給萬物的上帝面前，並在向 本丟．彼拉多 作過那美好見證的基督耶穌面前囑咐你 ：
1TIM|6|14|要守這命令，毫不玷污，無可指責，直到我們的主耶穌基督顯現。
1TIM|6|15|到了適當的時候都要顯明出來： 他是那可稱頌、獨一的權能者， 萬王之王， 萬主之主，
1TIM|6|16|就是那獨一不死、 住在人不能靠近的光裏， 是人未曾看見，也是不能看見的。 願尊貴和永遠的權能都歸給他。阿們！
1TIM|6|17|至於那些今世富足的人，你要囑咐他們不要自高，也不要倚賴靠不住的錢財；要倚靠那厚賜萬物給我們享受的上帝。
1TIM|6|18|又要囑咐他們行善，在好事上富足，甘心施捨，樂意分享，
1TIM|6|19|為自己積存財富，而為將來打美好的根基，好使他們能把握那真正的生命。
1TIM|6|20|提摩太 啊，要持守所給你的託付。要躲避世俗的空談和那假冒知識的矛盾言論。
1TIM|6|21|有人自稱有這知識而偏離了信仰。 願恩惠與你們同在！
