DAN|1|1|Anno tertio regni Ioachim regis Iudae venit Nabuchodonosor rex Babylonis Ierusalem et obsedit eam;
DAN|1|2|et tradidit Dominus in manu eius Ioachim regem Iudae et partem vasorum domus Dei, et asportavit ea in terram Sennaar in domum deorum suorum et vasa intulit in domum thesauri deorum suorum.
DAN|1|3|Et ait rex Asfanaz praeposito eunuchorum suorum, ut introduceret de filiis Israel et de semine regio et tyrannorum
DAN|1|4|pueros, in quibus nulla esset macula, decoros forma et eruditos omni sapientia, cautos scientia et doctos disciplina, et qui possent stare in palatio regis, et ut docerent eos litteras et linguam Chaldaeorum.
DAN|1|5|Et constituit eis rex annonam per singulos dies de cibis suis et de vino, unde bibebat ipse, ut enutriti tribus annis postea starent in conspectu regis.
DAN|1|6|Fuerunt ergo inter eos de filiis Iudae Daniel, Ananias, Misael et Azarias.
DAN|1|7|Et imposuit eis praepositus eunuchorum nomina: Danieli Baltassar et Ananiae Sedrac, Misaeli Misac et Azariae Abdenago.
DAN|1|8|Proposuit autem Daniel in corde suo, ne pollueretur de mensa regis neque de vino potus eius, et rogavit eunuchorum praepositum, ne contaminaretur.
DAN|1|9|Dedit autem Deus Danieli gratiam et misericordiam in conspectu principis eunuchorum;
DAN|1|10|et ait princeps eunuchorum ad Daniel: " Timeo ego dominum meum regem, qui constituit vobis cibum et potum; qui si viderit vultus vestros macilentiores prae ceteris adulescentibus coaevis vestris, condemnabitis caput meum regi ".
DAN|1|11|Et dixit Daniel ad custodem, quem constituerat princeps eunuchorum super Daniel, Ananiam, Misael et Azariam:
DAN|1|12|" Tenta nos, obsecro, servos tuos diebus decem, et dentur nobis legumina ad vescendum et aqua ad bibendum;
DAN|1|13|et videantur in conspectu tuo vultus nostri et vultus puerorum, qui vescuntur cibo regio, et, sicut videris, facies cum servis tuis ".
DAN|1|14|Qui, audito sermone huiuscemodi, tentavit eos diebus decem.
DAN|1|15|Post dies autem decem apparuerunt vultus eorum meliores et corpulentiores prae omnibus pueris, qui vescebantur cibo regio.
DAN|1|16|Porro custos tollebat cibaria et vinum potus eorum dabatque eis legumina.
DAN|1|17|Quattuor autem pueris his dedit Deus scientiam et disciplinam in omni scriptura et sapientia, Danieli autem intellegentiam omnium visionum et somniorum.
DAN|1|18|Completis itaque diebus, post quos dixerat rex, ut introducerentur, introduxit eos praepositus eunuchorum in conspectu Nabuchodonosor.
DAN|1|19|Cumque locutus eis fuisset rex, non sunt inventi de universis tales ut Daniel, Ananias, Misael et Azarias; et steterunt in conspectu regis.
DAN|1|20|Et omne verbum sapientiae et intellectus, quod sciscitatus est ab eis, rex invenit in eis decuplum super cunctos hariolos et magos, qui erant in universo regno eius.
DAN|1|21|Fuit autem Daniel usque ad annum primum Cyri regis.
DAN|2|1|In anno secundo regni Nabu chodonosor vidit Nabuchodo nosor somnium, et conterritus est spiritus eius, et somnus eius fugit ab eo.
DAN|2|2|Praecepit autem rex, ut convocarentur harioli et magi et malefici et Chaldaei et indicarent regi somnia sua; qui cum venissent, steterunt coram rege.
DAN|2|3|Et dixit ad eos rex: " Vidi somnium, et spiritus meus conterritus est, ut intellegat somnium ".
DAN|2|4|Responderuntque Chaldaei regi Aramaice: " Rex, in sempiternum vive! Dic somnium servis tuis, et interpretationem eius indicabimus ".
DAN|2|5|Et respondens rex ait Chaldaeis: " Sermo recessit a me. Nisi indicaveritis mihi somnium et coniecturam eius, in frusta concidemini, et domus vestrae in sterquilinium ponentur;
DAN|2|6|si autem somnium et coniecturam eius narraveritis, praemia et dona et honorem multum accipietis a me. Somnium igitur et interpretationem eius indicate mihi ".
DAN|2|7|Responderunt secundo atque dixerunt: " Rex somnium dicat servis suis, et interpretationem illius indicabimus ".
DAN|2|8|Respondit rex et ait: " Certe novi quia tempus redimitis, scientes quod recesserit a me sermo.
DAN|2|9|Si ergo somnium non indicaveritis mihi, una est de vobis sententia. Et verbum fallax et deceptione plenum composuistis, ut loquamini mihi, donec tempus pertranseat; somnium itaque dicite mihi, ut sciam quod interpretationem eius loquamini mihi ".
DAN|2|10|Respondentes ergo Chaldaei coram rege dixerunt: " Non est homo super terram qui sermonem regis possit indicare; quapropter neque regum quisquam magnus et potens verbum huiuscemodi sciscitatur ab omni hariolo et mago et Chaldaeo.
DAN|2|11|Sermo enim, quem tu quaeris, rex, gravis est, nec reperietur quisquam qui indicet illum in conspectu regis, exceptis diis, quorum non est cum hominibus conversatio ".
DAN|2|12|Quo audito, rex in furore et in ira magna praecepit, ut perirent omnes sapientes Babylonis.
DAN|2|13|Et egressa sententia, ut sapientes interficerentur, quaerebantur Daniel et socii eius, ut perirent.
DAN|2|14|Tunc Daniel interrogavit cum consilio et prudentia Arioch, principem militiae regis, qui egressus fuerat ad interficiendos sapientes Babylonis;
DAN|2|15|respondens dixit ad Arioch, qui a rege potestatem acceperat, quam ob causam tam crudelis sententia a facie esset regis egressa. Cum ergo rem indicasset Arioch Danieli,
DAN|2|16|Daniel ingressus rogavit regem, ut tempus daret sibi ad solutionem indicandam regi;
DAN|2|17|et ingressus est domum suam Ananiaeque, Misaeli et Azariae sociis suis indicavit negotium,
DAN|2|18|ut quaererent misericordiam a facie Dei caeli super sacramento isto et non perirent Daniel et socii eius cum ceteris sapientibus Babylonis.
DAN|2|19|Tunc Danieli per visionem nocte mysterium revelatum est, et benedixit Daniel Deo caeli
DAN|2|20|et locutus Daniel ait: Sit nomen Dei benedictuma saeculo et usque in saeculum,quia sapientia et fortitudo eius sunt;
DAN|2|21|et ipse mutat tempora et aetates,transfert atque constituit reges,dat sapientiam sapientibuset scientiam intellegentibus disciplinam:
DAN|2|22|ipse revelat profunda et absconditaet novit in tenebris constituta,et lux cum eo inhabitat,
DAN|2|23|Tibi, Deus patrum meorum, confiteor teque laudo,quia sapientiam et fortitudinem dedisti mihiet nunc ostendisti mihi, quae rogavimus te,quia sermonem regis aperuisti nobis ".
DAN|2|24|Propterea Daniel, ingressus ad Arioch, quem constituerat rex, ut perderet sapientes Babylonis, sic ei locutus est: " Sapientes Babylonis ne perdas; introduc me in conspectu regis et solutionem regi enarrabo ".
DAN|2|25|Tunc Arioch festinus introduxit Danielem ad regem et dixit ei: " Inveni hominem de filiis transmigrationis Iudae, qui solutionem regi annuntiet ".
DAN|2|26|Respondit rex et dixit Danieli, cuius nomen erat Baltassar: " Putasne vere potes mihi indicare somnium, quod vidi, et interpretationem eius?".
DAN|2|27|Et respondens Daniel coram rege ait: " Mysterium, quod rex interrogat, sapientes, magi et harioli et haruspices non queunt indicare regi;
DAN|2|28|sed est Deus in caelo revelans mysteria, qui indicavit tibi, rex Nabuchodonosor, quae ventura sunt in novissimis temporibus. Somnium tuum et visiones capitis tui in cubili tuo huiuscemodi sunt:
DAN|2|29|Tu, rex, cogitare coepisti in strato tuo quid esset futurum post haec; et, qui revelat mysteria, ostendit tibi, quae ventura sunt.
DAN|2|30|Mihi quoque non in sapientia, quae est in me plus quam in cunctis viventibus, sacramentum hoc revelatum est, sed ut interpretatio regi manifesta fieret, et cogitationes mentis tuae scires.
DAN|2|31|Tu, rex, videbas, et ecce statua una grandis: statua illa magna et statura sublimis stabat contra te, et intuitus eius erat terribilis.
DAN|2|32|Huius statuae caput ex auro optimo erat, pectus autem et brachia de argento, porro venter et femora ex aere,
DAN|2|33|tibiae autem ferreae, pedum quaedam pars erat ferrea, quaedam autem fictilis.
DAN|2|34|Videbas ita, donec abscissus est lapis sine manibus et percussit statuam in pedibus eius ferreis et fictilibus et comminuit eos;
DAN|2|35|tunc contrita sunt pariter ferrum, testa, aes, argentum et aurum, et fuerunt quasi folliculus ex areis aestivis, et rapuit ea ventus, nullusque locus inventus est eis; lapis autem, qui percusserat statuam, factus est mons magnus et implevit universam terram.
DAN|2|36|Hoc est somnium; interpretationem quoque eius dicemus coram te, rex.
DAN|2|37|Tu rex regum es, et Deus caeli regnum et fortitudinem et imperium et gloriam dedit tibi;
DAN|2|38|et omnia, in quibus habitant filii hominum et bestiae agri volucresque caeli, dedit in manu tua et te dominum universorum constituit: tu es caput aureum.
DAN|2|39|Et post te consurget regnum aliud minus te et regnum tertium aliud aereum, quod imperabit universae terrae.
DAN|2|40|Et regnum quartum erit robustum velut ferrum; quomodo ferrum comminuit et domat omnia, et sicut ferrum comminuens conteret et comminuet omnia haec.
DAN|2|41|Porro quia vidisti pedum et digitorum partem testae figuli et partem ferream, regnum divisum erit; et robur ferri erit ei, secundum quod vidisti ferrum mixtum testae ex luto.
DAN|2|42|Et digitos pedum ex parte ferreos et ex parte fictiles, ex parte regnum erit solidum et ex parte contritum.
DAN|2|43|Quod autem vidisti ferrum mixtum testae ex luto, commiscebuntur quidem humano semine, sed non adhaerebunt sibi, sicuti ferrum misceri non potest testae.
DAN|2|44|In diebus autem regnorum illorum suscitabit Deus caeli regnum, quod in aeternum non dissipabitur, et regnum populo alteri non tradetur: comminuet et consumet universa regna haec, et ipsum stabit in aeternum.
DAN|2|45|Secundum quod vidisti quod de monte abscisus est lapis sine manibus et comminuit testam et ferrum et aes et argentum et aurum, Deus magnus ostendit regi, quae ventura sunt postea; et verum est somnium et fidelis interpretatio eius ".
DAN|2|46|Tunc rex Nabuchodonosor cecidit in faciem suam et Danielem adoravit et hostias et incensum praecepit, ut sacrificarent ei.
DAN|2|47|Loquens ergo rex ait Danieli: " Vere Deus vester Deus deorum est et Dominus regum et revelans mysteria, quoniam potuisti aperire sacramentum hoc ".
DAN|2|48|Tunc rex Danielem in sublime extulit et munera multa et magna dedit ei et constituit eum principem super omnes provincias Babylonis et principem praefectorum super cunctos sapientes Babylonis.
DAN|2|49|Daniel autem postulavit a rege et constituit super opera provinciae Babylonis Sedrac, Misac et Abdenago; ipse autem Daniel erat in foribus regis.
DAN|3|1|Nabuchodonosor rex fecit sta tuam auream altitudine cubito rum sexaginta, latitudine cubitorum sex; et statuit eam in campo Dura in provincia Babylonis.
DAN|3|2|Itaque Nabuchodonosor rex misit ad congregandos satrapas, magistratus et iudices, duces et tyrannos et praefectos omnesque principes provinciarum, ut convenirent ad dedicationem statuae, quam erexerat Nabuchodonosor rex.
DAN|3|3|Tunc congregati sunt satrapae, magistratus et iudices, duces et tyranni et optimates, qui erant in potestatibus constituti, et universi principes provinciarum ad dedicationem statuae, quam erexerat Nabuchodonosor rex. Stabant autem in conspectu statuae, quam posuerat Nabuchodonosor,
DAN|3|4|et praeco clamabat valenter: " Vobis dicitur, populi, tribus et linguae:
DAN|3|5|in hora, qua audieritis sonitum tubae et fistulae et citharae, sambucae et psalterii et symphoniae et universi generis musicorum, cadentes adorate statuam auream, quam constituit Nabuchodonosor rex.
DAN|3|6|Si quis autem non prostratus adoraverit, eadem hora mittetur in fornacem ignis ardentis ".
DAN|3|7|Post haec igitur, statim ut audierunt omnes populi sonitum tubae, fistulae et citharae, sambucae et psalterii et symphoniae et omnis generis musicorum, cadentes omnes populi tribus et linguae adoraverunt statuam auream, quam constituerat Nabuchodonosor rex.
DAN|3|8|Statimque et in ipso tempore accedentes viri Chaldaei accusaverunt Iudaeos
DAN|3|9|dixeruntque Nabuchodonosor regi: " Rex, in aeternum vive!
DAN|3|10|Tu, rex, posuisti decretum, ut omnis homo, qui audierit sonitum tubae, fistulae et citharae, sambucae et psalterii et symphoniae et universi generis musicorum, prosternat se et adoret statuam auream;
DAN|3|11|si quis autem non procidens adoraverit, mittetur in fornacem ignis ardentis.
DAN|3|12|Sunt ergo viri Iudaei, quos constituisti super opera provinciae Babylonis, Sedrac, Misac et Abdenago; viri isti te, rex, non honorant: deos tuos non colunt et statuam auream, quam erexisti, non adorant ".
DAN|3|13|Tunc Nabuchodonosor in furore et in ira praecepit, ut adducerentur Sedrac, Misac et Abdenago; tunc viri illi adducti sunt in conspectu regis.
DAN|3|14|Pronuntiansque Nabuchodonosor rex ait eis: " Verene, Sedrac, Misac et Abdenago, deos meos non colitis et statuam auream, quam constitui, non adoratis?
DAN|3|15|Numquid estis nunc parati, quacumque hora audieritis sonitum tubae, fistulae, citharae, sambucae, psalterii et symphoniae omnisque generis musicorum, prosternere vos et adorare statuam, quam feci? Quod si non adoraveritis, eadem hora mittemini in fornacem ignis ardentis; et quis est deus, qui eripiat vos de manu mea? ".
DAN|3|16|Respondentes Sedrac, Misac et Abdenago dixerunt regi Nabuchodonosor: " Non oportet nos de hac re respondere tibi:
DAN|3|17|Si enim Deus noster, quem colimus, potest eripere nos de camino ignis ardentis, et de manu tua, rex, liberabit.
DAN|3|18|Quod si noluerit, notum sit tibi, rex, quia deos tuos non colimus et statuam auream, quam erexisti, non adoramus ".
DAN|3|19|Tunc Nabuchodonosor repletus est furore, et aspectus faciei illius immutatus est super Sedrac, Misac et Abdenago; et respondens praecepit, ut succenderetur fornax septuplum quam succendi consueverat;
DAN|3|20|et viris fortissimis de exercitu suo iussit, ut ligarent Sedrac, Misac et Abdenago et mitterent eos in fornacem ignis ardentis;
DAN|3|21|et confestim viri illi vincti, cum bracis suis et tiaris et calceamentis et vestibus missi sunt in medium fornacis ignis ardentis;
DAN|3|22|itaque, quia iussio regis urgebat, et fornax succensa erat nimis, viros illos, qui miserant Sedrac, Misac et Abdenago, interfecit flamma ignis.
DAN|3|23|Viri autem tres, Sedrac, Misac et Abdenago, ceciderunt in medio camino ignis ardentis colligati.Quae sequuntur in Hebraeis voluminibus non repperi).
DAN|3|24|Et ambulabant in medio flammae laudantes Deum et benedicentes Domino.
DAN|3|25|Stans autem Azarias oravit sic aperiensque os suum in medio ignis ait:
DAN|3|26|" Benedictus es, Domine, Deus patrum nostrorum,et laudabilis et gloriosum nomen tuum in saecula,
DAN|3|27|quia iustus es in omnibus, quae fecisti nobis,et universa opera tua vera, et viae tuae rectae,et omnia iudicia tua veritas.
DAN|3|28|Iudicia enim vera fecistiiuxta omnia, quae induxisti super noset super civitatem sanctam patrum nostrorum Ierusalem,quia in veritate et in iudicio induxisti omnia haecpropter peccata nostra.
DAN|3|29|Peccavimus enim et inique egimus recedentes a teet deliquimus in omnibus;
DAN|3|30|et praecepta tua non audivimusnec observavimusnec fecimus, sicut praeceperas nobis,ut bene nobis esset.
DAN|3|31|Omnia ergo, quae induxisti super nos,et universa, quae fecisti nobis,vero iudicio fecisti;
DAN|3|32|et tradidisti nos in manibus inimicorum nostroruminiquorum et pessimorum praevaricatorumqueet regi iniusto et pessimo ultra omnem terram.
DAN|3|33|Et nunc non possumus aperire os;confusio et opprobrium facta suntservis tuis et his, qui colunt te.
DAN|3|34|Ne, quaesumus, tradas nos in perpetuumpropter nomen tuumet ne dissipes testamentum tuum
DAN|3|35|neque auferas misericordiam tuam a nobispropter Abraham dilectum tuumet Isaac servum tuumet Israel sanctum tuum,
DAN|3|36|quibus dixistiquod multiplicares semen eorum sicut stellas caeliet sicut arenam, quae est in litore maris;
DAN|3|37|quia, Domine,imminuti sumus plus quam omnes gentessumusque humiles in universa terrahodie propter peccata nostra;
DAN|3|38|et non est in tempore hocprinceps et propheta et duxneque holocaustum neque sacrificiumneque oblatio neque incensumneque locus primitiarum coram te,ut possimus invenire misericordiam;
DAN|3|39|sed in anima contrita et spiritu humilitatis suscipiamursicut in holocausto arietum et taurorum
DAN|3|40|et sicut in milibus agnorum pinguium;sic fiat sacrificium nostrum in conspectu tuo hodie,et perfice subsequentes te,quoniam non est confusio confidentibus in te.
DAN|3|41|Et nunc sequimur te in toto cordeet timemus te et quaerimus faciem tuam;
DAN|3|42|ne confundas nos,sed fac nobiscum iuxta mansuetudinem tuamet secundum multitudinem misericordiae tuae
DAN|3|43|et erue nos in mirabilibus tuiset da gloriam nomini tuo, Domine.
DAN|3|44|Et confundantur omnes, qui ostendunt servis tuis mala;confundantur absque ulla potentia,et robur eorum conteratur.
DAN|3|45|Sciant quia tu es Dominus,Deus solus et gloriosus super orbem terrarum ".
DAN|3|46|Et non cessabant, qui immiserant eos, ministri regis succendere fornacem naphta et stuppa et pice et malleolis,
DAN|3|47|et effundebatur flamma super fornacem cubitis quadraginta novem
DAN|3|48|et erupit et incendit, quos repperit iuxta fornacem de Chaldaeis.
DAN|3|49|Angelus autem Domini descendit cum Azaria et sociis eius in fornacem et excussit flammam ignis de fornace
DAN|3|50|et fecit medium fornacis quasi ventum roris flantem; et non tetigit eos omnino ignis neque contristavit nec quidquam molestiae intulit.
DAN|3|51|Tunc hi tres, quasi ex uno ore, laudabant et glorificabant et benedicebant Deo in fornace dicentes:
DAN|3|52|" Benedictus es, Domine, Deus patrum nostrorum,et laudabilis et superexaltatus in saecula;et benedictum nomen gloriae tuae sanctumet superlaudabile et superexaltatum in saecula.
DAN|3|53|Benedictus es in templo sanctae gloriae tuaeet superlaudabilis et supergloriosus in saecula.
DAN|3|54|Benedictus es in throno regni tuiet superlaudabilis et superexaltatus in saecula.
DAN|3|55|Benedictus es, qui intueris abyssos sedens super cherubim,et laudabilis et superexaltatus in saecula.
DAN|3|56|Benedictus es in firmamento caeliet laudabilis et gloriosus in saecula.
DAN|3|57|Benedicite, omnia opera Domini, Domino,laudate et superexaltate eum in saecula.
DAN|3|58|Benedicite, caeli, Domino,laudate et superexaltate eum in saecula.
DAN|3|59|Benedicite, angeli Domini, Domino,laudate et superexaltate eum in saecula.
DAN|3|60|Benedicite, aquae omnes, quae super caelos sunt, Domino,laudate et superexaltate eum in saecula.
DAN|3|61|Benedicat omnis virtus Domino,laudate et superexaltate eum in saecula.
DAN|3|62|Benedicite, sol et luna, Domino,laudate et superexaltate eum in saecula.
DAN|3|63|Benedicite, stellae caeli, Domino,laudate et superexaltate eum in saecula.
DAN|3|64|Benedicite, omnis imber et ros, Domino,laudate et superexaltate eum in saecula.
DAN|3|65|Benedicite, omnes venti, Domino,laudate et superexaltate eum in saecula.
DAN|3|66|Benedicite, ignis et aestus, Domino,laudate et superexaltate eum in saecula.
DAN|3|67|Benedicite, frigus et aestus, Domino,laudate et superexaltate eum in saecula.
DAN|3|68|Benedicite, rores et pruina, Domino,laudate et superexaltate eum in saecula.
DAN|3|69|Benedicite, gelu et frigus, Domino,laudate et superexaltate eum in saecula.
DAN|3|70|Benedicite, glacies et nives, Domino,laudate et superexaltate eum in saecula.
DAN|3|71|Benedicite, noctes et dies, Domino,laudate et superexaltate eum in saecula.
DAN|3|72|Benedicite, lux et tenebrae, Domino,laudate et superexaltate eum in saecula.
DAN|3|73|Benedicite, fulgura et nubes, Domino,laudate et superexaltate eum in saecula.
DAN|3|74|Benedicat terra Dominum,laudet et superexaltet eum in saecula.
DAN|3|75|Benedicite, montes et colles, Domino,laudate et superexaltate eum in saecula.
DAN|3|76|Benedicite, universa germinantia in terra, Domino,laudate et superexaltate eum in saecula.
DAN|3|77|Benedicite, maria et flumina, Domino,laudate et superexaltate eum in saecula.
DAN|3|78|Benedicite, fontes, Domino,laudate et superexaltate eum in saecula.
DAN|3|79|Benedicite, cete et omnia quae moventur in aquis, Domino,laudate et superexaltate eum in saecula.
DAN|3|80|Benedicite, omnes volucres caeli, Domino,laudate et superexaltate eum in saecula.
DAN|3|81|Benedicite, omnes bestiae et pecora, Domino,laudate et superexaltate eum in saecula.
DAN|3|82|Benedicite, filii hominum, Domino,laudate et superexaltate eum in saecula.
DAN|3|83|Benedic, Israel, Domino,laudate et superexaltate eum in saecula.
DAN|3|84|Benedicite, sacerdotes Domini, Domino,laudate et superexaltate eum in saecula.
DAN|3|85|Benedicite, servi Domini, Domino,laudate et superexaltate eum in saecula.
DAN|3|86|Benedicite, spiritus et animae iustorum, Domino,laudate et superexaltate eum in saecula.
DAN|3|87|Benedicite, sancti et humiles corde, Domino,laudate et superexaltate eum in saecula.
DAN|3|88|Benedicite, Anania, Azaria, Misael, Domino,laudate et superexaltate eum in saecula;quia eruit nos de inferno et salvos fecit de manu mortiset liberavit nos de medio fornacis ardentis flammaeet de medio ignis eruit nos.
DAN|3|89|Confitemini Domino, quoniam bonus,quoniam in saeculum misericordia eius.
DAN|3|90|Benedicite, omnes, qui timetis Dominum, Deo deorum;laudate et confitemini ei, quia in saecula misericordia eius ".Hucusque non habetur in Hebraeo et, quae posuimus, de Theodotionis editione translata sunt).
DAN|3|91|24 Tunc Nabuchodonosor rex obstupuit et surrexit propere; respondens ait optimatibus suis: " Nonne tres viros misimus in medium ignis compeditos?". Qui respondentes dixerunt regi: " Vere, rex ".
DAN|3|92|25 Respondit et ait: " Ecce ego video viros quattuor solutos et ambulantes in medio ignis, et nihil corruptionis in eis est, et species quarti similis filio deorum ".
DAN|3|93|26 Tunc accessit Nabuchodonosor ad ostium fornacis ignis ardentis et ait: " Sedrac, Misac et Abdenago, servi Dei excelsi, egredimini et venite. Statimque egressi sunt Sedrac, Misac et Abdenago de medio ignis.
DAN|3|94|27 Et congregati satrapae, magistratus et iudices et potentes regis contemplabantur viros illos, quoniam nihil potestatis habuisset ignis in corporibus eorum, et capillus capitis eorum non esset adustus, et sarabara eorum non fuissent immutata, et odor ignis non transisset per eos.
DAN|3|95|28 Et erumpens Nabuchodonosor ait: " Benedictus Deus eorum, Sedrac, Misac et Abdenago, qui misit angelum suum et eruit servos suos, qui crediderunt in eo, et verbum regis immutaverunt et tradiderunt corpora sua, ne servirent et ne adorarent omnem deum, excepto Deo suo.
DAN|3|96|29 A me ergo positum est decretum, ut omnis populus, tribus et lingua quaecumque locuta fuerit blasphemiam contra Deum Sedrac, Misac et Abdenago, in frusta concidatur, et domus eius in sterquilinium fiat, eo quod non est Deus alius, qui possit ita salvare ".
DAN|3|97|30 Tunc rex promovit Sedrac, Misac et Abdenago in provincia Babylonis.
DAN|3|98|31 Nabuchodonosor rex omnibus populis, gentibus et linguis, quae habitant in universa terra: " Pax vobis multiplicetur.
DAN|3|99|32 Signa et mirabilia, quae fecit apud me Deus excelsus, placuit mihi praedicare:
DAN|3|100|33 Signa eius quam magna sunt,et mirabilia eius quam fortia!Et regnum eius regnum sempiternum,et potestas eius in generationem et generationem ".
DAN|4|1|Ego Nabuchodonosor quietus eram in domo mea et florens in palatio meo;
DAN|4|2|somnium vidi, quod perterruit me, et cogitationes in stratu meo et visiones capitis mei conturbaverunt me.
DAN|4|3|Et per me propositum est decretum, ut introducerentur in conspectu meo cuncti sapientes Babylonis, ut solutionem somnii indicarent mihi.
DAN|4|4|Tunc ingrediebantur harioli, magi, Chaldaei et haruspices; et somnium narravi in conspectu eorum, et solutionem eius non indicaverunt mihi;
DAN|4|5|donec denique ingressus est in conspectu meo Daniel, cui nomen Baltassar secundum nomen dei mei et qui habet spiritum deorum sanctorum in semetipso. Et somnium coram ipso locutus sum:
DAN|4|6|Baltassar, princeps hariolorum, quem ego scio quod spiritum deorum sanctorum habeas in te, et omne sacramentum non est impossibile tibi, visiones somnii mei, quas vidi, et solutionem eius narra.
DAN|4|7|Visio capitis mei in cubili meo:Videbam, et ecce arbor in medio terrae,et altitudo eius nimia.
DAN|4|8|Magna arbor et fortis,et proceritas eius contingens caelum;aspectus illius erat usque ad terminos universae terrae.
DAN|4|9|Folia eius pulcherrima,et fructus eius nimius,et esca universorum in ea.Subter eam habitabant bestiae agri,et in ramis eius conversabantur volucres caeli,et ex ea vescebatur omnis caro.
DAN|4|10|Videbam in visione capitis mei super stratum meum,et ecce vigil et sanctus de caelo descendit.
DAN|4|11|Clamavit fortiter et sic ait:Succidite arborem et praecidite ramos eius,excutite folia eius et dispergite fructus eius.Fugiant bestiae de sub ea,et volucres de ramis eius.
DAN|4|12|Verumtamen germen radicum eius in terra siniteet in vinculo ferreo et aereo in herbis agri,et rore caeli tingatur,et cum feris pars eius in herba terrae.
DAN|4|13|Cor eius ab humano commutetur,et cor ferae detur ei,et septem tempora mutentur super eum.
DAN|4|14|In sententia vigilum decretum est,et sermo sanctorum petitio,ut cognoscant viventesquoniam dominatur Excelsus in regno hominumet, cuicumque voluerit, dabit illudet humillimum hominem constituet super eo".
DAN|4|15|Hoc somnium vidi ego rex Nabuchodonosor. Tu ergo, Baltassar, interpretationem narra, quia omnes sapientes regni mei non queunt solutionem edicere mihi; tu autem potes, quia spiritus deorum sanctorum in te est ".
DAN|4|16|Tunc Daniel, cuius nomen Baltassar, obstupuit quasi una hora, et cogitationes eius conturbabant eum. Respondens autem rex ait: " Baltassar, somnium et interpretatio eius non conturbent te ". Respondit Baltassar et dixit: " Domine mi, somnium his, qui te oderunt, et interpretatio eius hostibus tuis sit.
DAN|4|17|Arborem, quam vidisti sublimem atque robustam, cuius altitudo pertingit ad caelum, et aspectus illius in omnem terram,
DAN|4|18|et rami eius pulcherrimi, et fructus eius nimius, et esca omnium in ea, subter eam habitantes bestiae agri, et in ramis eius commorantes aves caeli,
DAN|4|19|tu es, rex, qui magnificatus es et invaluisti, et magnitudo tua crevit et pervenit usque ad caelum, et potestas tua in terminos terrae.
DAN|4|20|Quod autem vidit rex vigilem et sanctum descendere de caelo et dicere: Succidite arborem et dissipate illam; attamen germen radicum eius in terra dimittite, et vinculo ferreo et aereo in herbis agri, et rore caeli conspergatur, et cum feris sit pars eius, donec septem tempora mutentur super eum",
DAN|4|21|haec est interpretatio, rex, et sententia Altissimi, quae pervenit super dominum meum regem:
DAN|4|22|et eicient te ab hominibus, et cum bestiis feris erit habitatio tua, et fenum ut boves comedes et rore caeli infunderis; septem quoque tempora mutabuntur super te, donec scias quod dominetur Excelsus super regnum hominum et, cuicumque voluerit, det illud.
DAN|4|23|Quod autem praeceperunt, ut relinqueretur germen radicum eius, id est arboris, regnum tuum tibi manebit, postquam cognoveris potestatem caeli.
DAN|4|24|Quam ob rem, rex, consilium meum placeat tibi, et peccata tua eleemosynis redime et iniquitates tuas misericordiis pauperum; sic longitudo erit prosperitati tuae ".
DAN|4|25|Omnia haec venerunt super Nabuchodonosor regem.
DAN|4|26|Post finem mensium duodecim in palatio regni Babylonis deambulabat;
DAN|4|27|responditque rex et ait: " Nonne haec est Babylon magna, quam ego aedificavi in domum regni, in robore fortitudinis meae et in gloria decoris mei? ".
DAN|4|28|Cum adhuc sermo esset in ore regis, vox de caelo ruit: " Tibi dicitur, Nabuchodonosor rex: Regnum tuum transiit a te,
DAN|4|29|et ab hominibus te eicient, et cum bestiis feris erit habitatio tua: fenum quasi boves comedes; et septem tempora mutabuntur super te, donec scias quod dominetur Excelsus in regno hominum et, cuicumque voluerit, det illud ".
DAN|4|30|Eadem hora sermo completus est super Nabuchodonosor, et ex hominibus abiectus est et fenum ut boves comedit, et rore caeli corpus eius infectum est, donec capilli eius in similitudinem aquilarum crescerent, et ungues eius quasi avium.
DAN|4|31|" Igitur post finem dierum ego Nabuchodonosor oculos meos ad caelum levavi, et sensus meus redditus est mihi, et Altissimo benedixi et Viventem in sempiternum laudavi et glorificavi,quia potestas eius potestas sempiterna,et regnum eius in generationem et generationem;
DAN|4|32|et omnes habitatores terrae apud eum in nihilum reputati sunt:iuxta voluntatem enim suam facittam in virtutibus caeli quam in habitatoribus terrae,et non est qui resistat manui eiuset dicat ei: "Quid facis?".
DAN|4|33|In ipso tempore sensus meus reversus est ad me, et ad honorem regni mei maiestas mea et splendor meus reversa sunt ad me; et optimates mei et magistratus mei requisierunt me, et in regno meo constitutus sum, et magnificentia amplior addita est mihi.
DAN|4|34|Nunc igitur ego Nabuchodonosor laudo et magnifico et glorifico Regem caeli, quia omnia opera eius veritas, et viae eius iudicium, et gradientes in superbia potest humiliare ".
DAN|5|1|Balthasar rex fecit grande con vivium optimatibus suis mille et coram his milibus vinum bibebat.
DAN|5|2|Balthasar ergo praecepit iam temulentus, ut afferrentur vasa aurea et argentea, quae asportaverat Nabuchodonosor pater eius de templo, quod fuit in Ierusalem, ut biberent in eis rex et optimates eius uxoresque eius et concubinae.
DAN|5|3|Tunc allata sunt vasa aurea, quae asportaverat de templo, quod fuerat in Ierusalem; et biberunt in eis rex et optimates eius, uxores et concubinae illius:
DAN|5|4|bibebant vinum et laudabant deos suos aureos et argenteos, aereos, ferreos ligneosque et lapideos.
DAN|5|5|In eadem hora apparuerunt digiti manus hominis et scripserunt contra candelabrum in superficie parietis palatii regis; et rex aspiciebat articulos manus scribentis.
DAN|5|6|Tunc regis facies commutata est, et cogitationes eius conturbabant eum, et compages renum eius solvebantur, et genua eius ad se invicem collidebantur.
DAN|5|7|Exclamavit itaque rex fortiter, ut introducerent magos, Chaldaeos et haruspices; et proloquens rex ait sapientibus Babylonis: " Quicumque legerit scripturam hanc et interpretationem eius manifestam mihi fecerit, purpura vestietur et torquem auream habebit in collo et tertius in regno meo dominabitur ".
DAN|5|8|Tunc ingressi sunt omnes sapientes regis et non potuerunt nec scripturam legere nec interpretationem indicare regi;
DAN|5|9|unde rex Balthasar satis conturbatus est, et vultus illius immutatus est super eum, sed et optimates eius turbabantur.
DAN|5|10|Regina autem, sermonum regis optimatiumque eius causa, domum convivii ingressa est; et regina proloquens ait: " Rex, in aeternum vive! Non te conturbent cogitationes tuae, neque facies tua immutetur.
DAN|5|11|Est vir in regno tuo, qui spiritum deorum sanctorum habet in se, et in diebus patris tui scientia et intellegentia et sapientia quasi sapientia deorum inventae sunt in eo; nam et rex Nabuchodonosor pater tuus principem magorum, incantatorum, Chaldaeorum et haruspicum constituit eum; pater tuus, o rex,
DAN|5|12|quia spiritus amplior et prudentia intellegentiaque et interpretatio somniorum et ostensio secretorum ac solutio ligatorum inventae sunt in eo, in Daniele, cui rex posuit nomen Baltassar. Nunc itaque Daniel vocetur et interpretationem narrabit ".
DAN|5|13|Igitur introductus est Daniel coram rege; ad quem praefatus rex ait: " Tu es Daniel de filiis captivitatis Iudae, quem adduxit rex pater meus de Iuda?
DAN|5|14|Audivi de te quoniam spiritum deorum habeas, et scientia intellegentiaque ac sapientia ampliores inventae sint in te.
DAN|5|15|Et nunc introgressi sunt in conspectu meo sapientes, magi, ut scripturam hanc legerent et interpretationem eius indicarent mihi et nequiverunt sensum huius sermonis edicere.
DAN|5|16|Porro ego audivi de te quod possis obscura interpretari et ligata dissolvere; si ergo vales scripturam legere et interpretationem eius indicare mihi, purpura vestieris et torquem auream circa collum tuum habebis et tertius in regno meo princeps eris ".
DAN|5|17|Tunc respondens Daniel ait coram rege: " Munera tua sint tibi, et dona tua alteri da; scripturam autem legam tibi, rex, et interpretationem eius ostendam tibi.
DAN|5|18|O rex, Deus altissimus regnum et magnificentiam et gloriam et honorem dedit Nabuchodonosor patri tuo.
DAN|5|19|Et propter magnificentiam, quam dederat ei, universi populi, tribus et linguae tremebant et metuebant eum; quos volebat, interficiebat et, quos volebat, percutiebat et, quos volebat, exaltabat et, quos volebat, humiliabat.
DAN|5|20|Quando autem elevatum est cor eius, et spiritus illius obfirmatus est ad superbiam, depositus est de solio regni sui, et gloria eius ablata est ab eo;
DAN|5|21|et a filiis hominum eiectus est, sed et cor eius cum bestiis positum est, et cum onagris erat habitatio eius, fenum quoque ut boves comedebat, et rore caeli corpus eius infectum est, donec cognosceret quod potestatem haberet Deus altissimus in regno hominum et, quemcumque voluerit, suscitabit super illud.
DAN|5|22|Tu quoque filius eius, Balthasar, non humiliasti cor tuum, cum scires haec omnia,
DAN|5|23|sed adversum Dominum caeli elevatus es, et vasa domus eius allata sunt coram te, et tu et optimates tui et uxores tuae et concubinae tuae vinum bibistis in eis; deos quoque argenteos et aureos et aereos, ferreos ligneosque et lapideos, qui non vident neque audiunt neque sentiunt, laudasti, porro Deum, qui habet flatum tuum in manu sua et omnes vias tuas, non glorificasti.
DAN|5|24|Idcirco ab eo missi sunt articuli manus, et scriptura haec exarata est.
DAN|5|25|Haec est autem scriptura, quae digesta est: mane, thecel, upharsin.
DAN|5|26|Et haec est interpretatio sermonis: mane, numeravit Deus regnum tuum et complevit illud;
DAN|5|27|thecel, appensus es in statera et inventus es minus habens;
DAN|5|28|phares, divisum est regnum tuum et datum est Medis et Persis ".
DAN|5|29|Tunc, iubente Balthasar, indutus est Daniel purpura, et circumdata est torques aurea collo eius, et praedicatum est de eo quod haberet potestatem tertius in regno suo.
DAN|5|30|Eadem nocte interfectus est Balthasar rex Chaldaeorum.
DAN|6|1|Et Darius Medus successit in regnum annos natus sexaginta duos.
DAN|6|2|Placuit Dario et constituit super regnum satrapas centum viginti, ut essent in toto regno suo,
DAN|6|3|et super eos principes tres, ex quibus Daniel unus erat, ut satrapae illis redderent rationem, et rex non sustineret molestiam.
DAN|6|4|Igitur ille Daniel superabat omnes principes et satrapas, quia spiritus Dei amplior erat in eo. Porro rex cogitabat constituere eum super omne regnum;
DAN|6|5|unde principes et satrapae quaerebant, ut invenirent occasionem Danieli ex latere regni, nullamque causam et suspicionem reperire potuerunt, eo quod fidelis esset, et omnis culpa et suspicio non inveniretur in eo.
DAN|6|6|Dixerunt ergo viri illi: " Non inveniemus Danieli huic aliquam occasionem, nisi forte inveniamus adversus eum in lege Dei sui ".
DAN|6|7|Tunc principes et satrapae illi concurrerunt ad regem et sic locuti sunt ei: " Darie rex, in aeternum vive!
DAN|6|8|Consilium inierunt cuncti principes regni, magistratus et satrapae, optimates et iudices, ut decretum regis promulget et edictum confirmet, ut omnis, qui petierit aliquam petitionem a quocumque deo et homine usque ad dies triginta, nisi a te, rex, mittatur in lacum leonum.
DAN|6|9|Nunc itaque, rex, confirma sententiam et signa decretum, ut non immutetur iuxta legem Medorum et Persarum, quam praevaricari non licet ".
DAN|6|10|Porro rex Darius signavit edictum et decretum.
DAN|6|11|Daniel autem, cum comperisset decretum signatum esse, ingressus est domum suam et, fenestris apertis in cenaculo suo contra Ierusalem, tribus temporibus in die flectebat genua sua et adorabat confitebaturque coram Deo suo, sicut et ante facere consueverat.
DAN|6|12|Viri ergo illi accesserunt et invenerunt Danielem orantem et obsecrantem Deum suum.
DAN|6|13|Tunc accesserunt et locuti sunt coram rege super edicto: " Rex, numquid non signasti decretum, ut omnis homo, qui rogaret quemquam de diis et hominibus usque ad dies triginta, nisi a te, rex, mitteretur in lacum leonum? ". Respondens rex ait: " Verus est sermo iuxta decretum Medorum atque Persarum, quod praevaricari non licet ".
DAN|6|14|Tunc respondentes dixerunt coram rege: " Daniel de filiis captivitatis Iudae non curavit de te, rex, et de edicto, quod constituisti, sed tribus temporibus per diem orat obsecratione sua".
DAN|6|15|Quod verbum cum audisset, rex satis contristatus est; et pro Daniele posuit cor, ut liberaret eum, et usque ad occasum solis laborabat, ut erueret illum.
DAN|6|16|Viri autem illi accesserunt ad regem et dixerunt ei: " Scito, rex, quia lex Medorum est atque Persarum, ut omne decretum et edictum, quod constituit rex, non liceat immutari ".
DAN|6|17|Tunc rex praecepit, et adduxerunt Danielem et miserunt eum in lacum leonum. Dixitque rex Danieli: " Deus tuus, quem colis semper, ipse liberet te ".
DAN|6|18|Allatusque est lapis unus et positus est super os laci; quem obsignavit rex anulo suo et anulo optimatum suorum, ne quid fieret contra Danielem.
DAN|6|19|Et abiit rex in domum suam et dormivit incenatus, cibique non sunt illati coram eo; insuper et somnus recessit ab eo.
DAN|6|20|Tunc rex primo diluculo consurgens festinus ad lacum leonum perrexit;
DAN|6|21|appropinquansque lacui Danielem voce lacrimabili inclamavit et affatus est Danielem: " Daniel, serve Dei viventis, Deus tuus, cui tu servis semper, putasne valuit liberare te a leonibus?".
DAN|6|22|Et Daniel regi respondens ait: " Rex, in aeternum vive!
DAN|6|23|Deus meus misit angelum suum et conclusit ora leonum, et non nocuerunt mihi, quia coram eo iustitia inventa est in me; sed et coram te, rex, delictum non feci ".
DAN|6|24|Tunc rex vehementer gavisus est super eo et Danielem praecepit educi de lacu; eductusque est Daniel de lacu, et nulla laesio inventa est in eo, quia credidit Deo suo.
DAN|6|25|Dixit autem rex, et adducti sunt viri illi, qui accusaverant Danielem, et in lacum leonum missi sunt, ipsi et filii eorum et uxores eorum, et non pervenerunt usque ad pavimentum laci, donec potirentur eis leones, et omnia ossa eorum comminuerunt.
DAN|6|26|Tunc Darius rex scripsit universis populis, tribubus et linguis, habitantibus in universa terra: "Pax vobis multiplicetur!
DAN|6|27|A me constitutum est decretum, ut in universo imperio regni mei tremescant et paveant Deum Danielis:ipse est enim Deus vivenset permanens in saecula,et regnum eius non dissipabitur,et potestas eius usque in aeternum;
DAN|6|28|ipse liberator atque salvatoret faciens signa et mirabiliain caelo et in terra.Liberavit autem Danielemde manu leonum ".
DAN|6|29|Porro Daniel prosperatus est in regno Darii et in regno Cyri Persae.
DAN|7|1|Anno primo Balthasar regis Babylonis Daniel somnium vidit et visionem capitis eius in cubili suo; tunc et somnium scripsit. Caput verborum, quae locutus est.
DAN|7|2|Respondit Daniel et dixit: " Videbam in visione mea nocte: et ecce quattuor venti caeli conturbabant mare Magnum,
DAN|7|3|et quattuor bestiae grandes ascendebant de mari diversae inter se.
DAN|7|4|Prima quasi leaena et alas habebat aquilae; aspiciebam, donec evulsae sunt alae eius; et sublata est de terra et super pedes quasi homo stetit, et cor hominis datum est ei.
DAN|7|5|Et ecce bestia alia, secunda, similis urso in parte stetit, et tres costae erant in ore eius et in dentibus eius; et sic dicebant ei: "Surge, comede carnes plurimas".
DAN|7|6|Post hoc aspiciebam, et ecce alia quasi pardus et alas habebat avis quattuor super se, et quattuor capita erant in bestia; et potestas data est ei.
DAN|7|7|Post hoc aspiciebam in visione noctis, et ecce bestia quarta terribilis atque mirabilis et fortis nimis; dentes ferreos habebat magnos, comedens atque comminuens et reliqua pedibus suis conculcans; dissimilis autem erat ceteris bestiis, quas videram ante eam, et habebat cornua decem.
DAN|7|8|Considerabam cornua, et ecce cornu aliud parvulum ortum est de medio eorum, et tria de cornibus primis evulsa sunt a facie eius; et ecce oculi quasi oculi hominis erant in cornu isto, et os loquens ingentia.
DAN|7|9|Aspiciebam,donec throni positi sunt,et Antiquus dierum sedit.Vestimentum eius quasi nix candidum,et capilli capitis eius quasi lana munda;thronus eius flammae ignis,rotae eius ignis accensus.
DAN|7|10|Fluvius igneus effluebatet egrediebatur a facie eius;milia milium ministrabant ei,et decies milies centena milia assistebant ei:iudicium sedit,et libri aperti sunt.
DAN|7|11|Aspiciebam tunc propter vocem sermonum grandium, quos cornu illud loquebatur; et vidi quoniam interfecta esset bestia, et perisset corpus eius, et tradita esset ad comburendum igni;
DAN|7|12|aliarum quoque bestiarum ablata esset potestas, et tempora vitae constituta essent eis usque ad tempus et tempus.
DAN|7|13|Aspiciebam ergo in visione noctis:et ecce cum nubibus caeliquasi Filius hominis veniebatet usque ad Antiquum dierum pervenit,et in conspectu eius obtulerunt eum;
DAN|7|14|et data sunt ei potestas et honor et regnum;et omnes populi, tribus et linguaeipsi servierunt:potestas eius potestas aeterna,quae non auferetur,et regnum eius, quod non corrumpetur.
DAN|7|15|Horruit spiritus meus: ego Daniel territus sum in his, et visiones capitis mei conturbaverunt me.
DAN|7|16|Accessi ad unum de assistentibus et veritatem quaerebam ab eo de omnibus his; qui dixit mihi et interpretationem sermonum edocuit me:
DAN|7|17|"Hae bestiae magnae quattuor, quattuor regna consurgent de terra;
DAN|7|18|suscipient autem regnum sancti Dei altissimi et obtinebunt regnum usque in saeculum et saeculum saeculorum".
DAN|7|19|Post hoc volui diligenter discere de bestia quarta, quae erat dissimilis valde ab omnibus his et terribilis nimis, dentes ferrei et ungues eius aerei, comedens et comminuens et reliquias pedibus suis conculcans,
DAN|7|20|et de cornibus decem, quae habebat in capite, et de alio, quod ortum fuerat ante, et ceciderant tria cornua, de cornu illo, quod habebat oculos et os loquens grandia et maius erat ceteris.
DAN|7|21|Aspiciebam, et ecce cornu illud faciebat bellum adversus sanctos et praevalebat eis,
DAN|7|22|donec venit Antiquus dierum et iudicium dedit sanctis Excelsi, et tempus advenit, et regnum obtinuerunt sancti.
DAN|7|23|Et sic ait: "Bestia quarta regnum quartum erit in terra, quod maius erit omnibus regnis et devorabit universam terram et conculcabit et comminuet eam.
DAN|7|24|Porro cornua decem regni decem reges erunt; et alius consurget post eos et ipse potentior erit prioribus et tres reges humiliabit
DAN|7|25|et sermones contra Excelsum loquetur et sanctos Altissimi conteret et putabit quod possit mutare tempora et legem, et tradentur in manu eius usque ad tempus et tempora et dimidium temporis;
DAN|7|26|et iudicium sedebit, et potentiam eius auferent, ut conteratur et dispereat usque in finem;
DAN|7|27|regnum autem et potestas et magnitudo regnorum, quae sunt subter omne caelum, detur populo sanctorum Altissimi, cuius regnum regnum sempiternum est, et omnes reges servient ei et oboedient" ".
DAN|7|28|Hucusque finis verbi. Ego Daniel multum cogitationibus meis conturbabar, et facies mea mutata est in me; verbum autem in corde meo conservavi.
DAN|8|1|Anno tertio regni Balthasar regis visio apparuit mihi, ego Daniel, post id quod mihi apparuerat in principio.
DAN|8|2|Vidi in visione, et factum est, dum viderem, eram in Susis castro, quod est in Elam provincia; vidi autem in visione esse me super rivum Ulai.
DAN|8|3|Et levavi oculos meos et vidi: et ecce aries unus stabat ante rivum habens cornua et cornua excelsa et unum excelsius altero, et excelsius crescebat in postero.
DAN|8|4|Vidi arietem cornibus ventilantem contra occidentem et contra aquilonem et contra meridiem, et omnes bestiae non poterant resistere ei neque liberari de manu eius; fecitque secundum voluntatem suam et magnificatus est.
DAN|8|5|Et ego intellegebam: ecce autem hircus caprarum veniebat ab occidente super faciem totius terrae et non tangebat terram; porro hircus habebat cornu insigne inter oculos suos.
DAN|8|6|Et venit usque ad arietem illum cornutum, quem videram stantem ante rivum, et cucurrit ad eum in impetu fortitudinis suae.
DAN|8|7|Vidi eum appropinquantem prope arietem, et efferatus est in eum et percussit arietem et comminuit duo cornua eius, et non poterat aries resistere ei; cumque eum misisset in terram, conculcavit, et nemo quibat liberare arietem de manu eius.
DAN|8|8|Hircus autem caprarum magnus factus est nimis; cumque crevisset, fractum est cornu magnum, et orta sunt quattuor cornua loco illius per quattuor ventos caeli.
DAN|8|9|De uno autem ex eis egressum est cornu unum modicum et factum est grande contra meridiem et contra orientem et contra fortitudinem
DAN|8|10|et magnificatum est usque ad fortitudinem caeli et deiecit de fortitudine et de stellis et conculcavit eas;
DAN|8|11|et usque ad principem fortitudinis magnificatum est et ab eo tulit iuge sacrificium et deiecit locum sanctificationis eius.
DAN|8|12|Militia autem data est contra iuge sacrificium propter peccata, et prostrata est veritas in terra; cornu autem fecit et prosperatum est.
DAN|8|13|Et audivi unum de sanctis loquentem, et dixit unus sanctus alteri, nescio cui, loquenti: " Usquequo visio et iuge sacrificium et peccatum desolationis, quae facta est, et sanctuarium et fortitudo conculcabitur?.
DAN|8|14|Et dixit ei: " Usque ad vesperam et mane, dies duo milia trecenti; et mundabitur sanctuarium ".
DAN|8|15|Factum est autem cum viderem ego Daniel visionem et quaererem intellegentiam, ecce stetit in conspectu meo quasi species viri;
DAN|8|16|et audivi vocem viri inter Ulai, et clamavit et ait: " Gabriel, fac intellegere istum visionem ".
DAN|8|17|Et venit et stetit iuxta, ubi ego stabam; cumque venisset, pavens corrui in faciem meam, et ait ad me: "Intellege, fili hominis, quoniam in tempore finis complebitur visio ".
DAN|8|18|Cumque loqueretur ad me, collapsus sum pronus in terram, et tetigit me et statuit me in gradu meo
DAN|8|19|dixitque: " Ecce ego ostendam tibi, quae futura sint in novissimo maledictionis, quoniam in tempore erit finis.
DAN|8|20|Aries, quem vidisti habere cornua, reges Medorum est atque Persarum;
DAN|8|21|porro hircus caprarum rex Graecorum est, et cornu grande, quod erat inter oculos eius, ipse est rex primus.
DAN|8|22|Quod autem, fracto illo, surrexerunt quattuor pro eo, quattuor regna de gente eius consurgent sed non in fortitudine eius.
DAN|8|23|Et post regnum eorum, cum creverint iniquitate, consurget rex impudens facie et intellegens propositiones;
DAN|8|24|et roborabitur fortitudo eius sed non in viribus suis, et supra quam credi potest universa vastabit et prosperabitur et faciet et interficiet robustos et populum sanctorum,
DAN|8|25|et secundum sapientiam suam prosperabitur dolus in manu eius, et in corde suo magnificabitur et in tranquillitate occidet plurimos et contra principem principum consurget et sine manu conteretur.
DAN|8|26|Et visio vespere et mane, quae dicta est, vera est; tu ergo signa visionem, quia post dies multos erit ".
DAN|8|27|Et ego Daniel langui et aegrotavi per dies; cumque surrexissem, faciebam opera regis et stupebam ad visionem, et non erat qui intellegeret.
DAN|9|1|In anno primo Darii filii Asueri de semine Medorum, qui impe ravit super regnum Chaldaeorum,
DAN|9|2|anno uno regni eius, ego Daniel intellexi in libris numerum annorum, de quo factus est sermo Domini ad Ieremiam prophetam, ut complerentur desolationes Ierusalem, septuaginta anni;
DAN|9|3|et posui faciem meam ad Dominum Deum meum, ut quaererem rogationem et deprecationem in ieiuniis, sacco et cinere.
DAN|9|4|Et oravi Dominum Deum et confessus sum et dixi: Obsecro, Domine, Deus magne et terribilis, custodiens pactum et misericordiam diligentibus eum et custodientibus mandata eius;
DAN|9|5|peccavimus, inique fecimus, impie egimus et recessimus et declinavimus a mandatis tuis ac iudiciis tuis;
DAN|9|6|non oboedivimus servis tuis prophetis, qui locuti sunt in nomine tuo regibus nostris, principibus nostris, patribus nostris omnique populo terrae.
DAN|9|7|Tibi, Domine, iustitia; nobis autem confusio faciei, sicut est hodie viro Iudae et habitatoribus Ierusalem et omni Israel, his qui prope sunt et his qui procul in universis terris, ad quas eiecisti eos propter iniquitates eorum, in quibus peccaverunt in te.
DAN|9|8|Domine, nobis confusio faciei, regibus nostris, principibus nostris et patribus nostris, quia peccavimus tibi;
DAN|9|9|Domino autem, Deo nostro, misericordia et propitiatio, quia recessimus a te.
DAN|9|10|Et non audivimus vocem Domini Dei nostri, ut ambularemus in lege eius, quam posuit nobis per servos suos prophetas;
DAN|9|11|et omnis Israel praevaricati sunt legem tuam et declinaverunt, ne audirent vocem tuam, et stillavit super nos maledictio et detestatio, quae scripta est in libro Moysis servi Dei, quia peccavimus ei.
DAN|9|12|Et statuit sermones suos, quos locutus est super nos et super iudices nostros, qui iudicaverunt nos, ut superducerent in nos magnum malum, quale numquam fuit sub omni caelo, secundum quod factum est in Ierusalem.
DAN|9|13|Sicut scriptum est in lege Moysis, omne malum hoc venit super nos, et non rogavimus faciem Domini Dei nostri, ut reverteremur ab iniquitatibus nostris et cogitaremus veritatem tuam.
DAN|9|14|Et vigilavit Dominus super malitiam et adduxit eam super nos, quia iustus Dominus Deus noster in omnibus operibus suis, quae fecit; non enim audivimus vocem eius.
DAN|9|15|Et nunc, Domine Deus noster, qui eduxisti populum tuum de terra Aegypti in manu forti et fecisti tibi nomen secundum diem hanc, peccavimus, iniquitatem fecimus,
DAN|9|16|Domine, in omnem iustitiam tuam; avertatur, obsecro, ira tua et furor tuus a civitate tua Ierusalem et monte sancto tuo; propter peccata enim nostra et iniquitates patrum nostrorum Ierusalem et populus tuus in opprobrium sunt omnibus per circuitum nostrum.
DAN|9|17|Nunc ergo exaudi, Deus noster, orationem servi tui et preces eius et ostende faciem tuam super sanctuarium tuum, quod desertum est, propter temetipsum.
DAN|9|18|Inclina, Deus meus, aurem tuam et audi; aperi oculos tuos et vide desolationem nostram et civitatem, super quam invocatum est nomen tuum; neque enim in iustificationibus nostris prosternimus preces ante faciem tuam sed in miserationibus tuis multis.
DAN|9|19|Exaudi, Domine! Placare, Domine! Attende et fac! Ne moreris propter temetipsum, Deus meus, quia nomen tuum invocatum est super civitatem et super populum tuum ".
DAN|9|20|Cumque adhuc loquerer et orarem et confiterer peccata mea et peccata populi mei Israel et prosternerem preces meas in conspectu Dei mei pro monte sancto Dei mei,
DAN|9|21|adhuc me loquente in oratione, ecce vir Gabriel, quem videram in visione principio, cito volans tetigit me in tempore sacrificii vespertini;
DAN|9|22|et docuit me et locutus est mihi dixitque: "Daniel, nunc egressus sum, ut docerem te, et intellegeres.
DAN|9|23|Ab exordio precum tuarum egressus est sermo; ego autem veni, ut indicarem, quia vir desideriorum es tu; ergo animadverte sermonem et intellege visionem.
DAN|9|24|Septuaginta hebdomades decretae suntsuper populum tuum et super urbem sanctam tuam,ut consummetur praevaricatio,et finem accipiat peccatum,et deleatur iniquitas,et adducatur iustitia sempiterna,et impleatur visio et prophetes,et ungatur Sanctus sanctorum.
DAN|9|25|Scito ergo et animadverte:ab exitu sermonisut iterum aedificetur Ierusalemusque ad christum ducem,hebdomades septem.Et hebdomades sexaginta duae erunt;et rursum aedificabitur platea et muriin angustia temporum.
DAN|9|26|Et post hebdomades sexaginta duasoccidetur christus;et nihil erit ei.Et civitatem et sanctuarium dissipabitpopulus ducis venturi,et finis eius vastitas,et usque ad finem bellistatuta desolatio.
DAN|9|27|Confirmabit autem pactum multishebdomade una;et in dimidio hebdomadideficiet hostia et sacrificium,et erit super alam abominationis vastator,et usquedum consummatio et decretumeffundantur super vastatorem ".
DAN|10|1|Anno tertio Cyri regis Per sarum verbum revelatum est Danieli cognomento Baltassar, et verum verbum et acies magna; intellexitque sermonem, intellegentia enim fuit ei in visione.
DAN|10|2|In diebus illis ego Daniel lugebam tribus hebdomadis dierum,
DAN|10|3|panem desiderabilem non comedi, et caro et vinum non introierunt in os meum, sed neque unguento unctus sum, donec complerentur tres hebdomades dierum.
DAN|10|4|Die autem vicesima et quarta mensis primi eram iuxta fluvium magnum, qui est Tigris,
DAN|10|5|et levavi oculos meos et vidi: et ecce vir unus vestitus lineis, et renes eius accincti auro obryzo;
DAN|10|6|et corpus eius quasi chrysolithus, et facies eius velut species fulgoris, et oculi eius ut lampas ardens, et brachia eius et, quae deorsum sunt usque ad pedes, quasi species aeris candentis, et vox sermonum eius ut vox multitudinis.
DAN|10|7|Vidi autem ego Daniel solus visionem; porro viri, qui erant mecum, visionem non viderunt, sed terror nimius irruit super eos, et fugerunt in absconditum.
DAN|10|8|Ego autem relictus solus vidi visionem grandem hanc, et non remansit in me fortitudo, sed et species mea immutata est in me usque ad dissipationem, nec habui quidquam virium.
DAN|10|9|Et audivi vocem sermonum eius; et audiens vocem sermonum eius iacebam consternatus super faciem meam, et vultus meus haerebat terrae.
DAN|10|10|Et ecce manus tetigit me et erexit me super genua mea et super palmas manuum mearum,
DAN|10|11|et dixit ad me: " Daniel, vir desideriorum, intellege verba, quae ego loquor ad te, et sta in gradu tuo; nunc enim sum missus ad te ". Cumque dixisset mihi sermonem istum, steti tremens.
DAN|10|12|Et ait ad me: " Noli metuere, Daniel, quia ex die primo, quo posuisti cor tuum ad intellegendum et ad humiliandum te in conspectu Dei tui, exaudita sunt verba tua; et ego veni propter sermones tuos.
DAN|10|13|Princeps autem regni Persarum restitit mihi viginti et uno diebus; et ecce Michael, unus de principibus primis, venit in adiutorium meum; et ego remansi ibi iuxta regem Persarum.
DAN|10|14|Veni autem, ut docerem te, quae ventura sunt populo tuo in novissimis diebus, quoniam adhuc visio in dies ".
DAN|10|15|Cumque loqueretur mihi huiuscemodi verbis, deieci vultum meum ad terram et tacui.
DAN|10|16|Et ecce quasi similitudo filiorum hominis tetigit labia mea; et aperiens os meum locutus sum et dixi ad eum, qui stabat contra me: " Domine mi, in visione angustiae venerunt super me, et nihil in me remansit virium.
DAN|10|17|Et quomodo poterit servus domini mei loqui cum hoc domino meo? Nihil enim in me remansit virium, et halitus meus non remansit in me ".
DAN|10|18|Rursum ergo tetigit me quasi visio hominis et confortavit me
DAN|10|19|et dixit: "Noli timere, vir desideriorum; pax tibi, confortare et esto robustus ". Cumque loqueretur mecum, convalui et dixi: " Loquere, domine mi, quia confortasti me ".
DAN|10|20|Et ait: " Numquid scis, quare venerim ad te? Et nunc revertar, ut proelier adversum principem Persarum. Et ego egrediar, et ecce princeps Graecorum veniens.
DAN|10|21|Verumtamen annuntiabo tibi, quod expressum est in scriptura veritatis; et nemo est adiutor meus adversus hos, nisi Michael princeps vester.
DAN|11|1|Ego autem ab anno primo Darii Medi astabam ei, ut confortaretur et roboraretur.
DAN|11|2|Et nunc veritatem annuntiabo tibi: Ecce adhuc tres reges stabunt pro Perside, et quartus ditabitur opibus nimis super omnes et, cum invaluerit divitiis suis, concitabit omnia adversum regnum Graeciae.
DAN|11|3|Surget vero rex fortis et dominabitur dominatione multa et faciet, quod placuerit ei;
DAN|11|4|et cum steterit, conteretur regnum eius et dividetur in quattuor ventos caeli, sed non in posteros eius neque secundum potentiam illius, qua dominatus est; lacerabitur enim regnum eius etiam ad alios, exceptis his.
DAN|11|5|Et confortabitur rex austri, et unus de principibus eius praevalebit super eum et dominabitur dominatione super dominationem eius.
DAN|11|6|Et post finem annorum foederabuntur; filiaque regis austri veniet ad regem aquilonis facere amicitiam. Et non obtinebit fortitudinem brachii, nec stabit brachium eius; et tradetur ipsa, et qui adduxerunt eam, et adulescens eius, et qui confortabat eam in temporibus.
DAN|11|7|Et stabit de germine radicum eius plantatio loco eius et veniet ad exercitum et ingredietur oppidum regis aquilonis; et faciet adversus eos et confortabitur.
DAN|11|8|Insuper et deos eorum cum sculptilibus eorum et vasis pretiosis argenti et auri captivos ducet in Aegyptum: ipse per aliquot annos praevalebit adversus regem aquilonis.
DAN|11|9|Et intrabit in regnum regis austri et revertetur ad terram suam.
DAN|11|10|Filii autem eius provocabuntur et congregabunt multitudinem exercituum plurimorum; et veniet properans et inundans et revertetur et concitabitur et congredietur usque ad oppidum eius.
DAN|11|11|Et provocabitur rex austri et egredietur et pugnabit adversus eum, adversus regem aquilonis; et praeparabit multitudinem nimiam, et dabitur multitudo in manu eius.
DAN|11|12|Et tolletur multitudo, et exaltabitur cor eius, et deiciet multa milia, sed non praevalebit.
DAN|11|13|Revertetur enim rex aquilonis et praeparabit multitudinem maiorem quam prius; et in fine temporum annorumque veniet properans cum exercitu magno et opibus nimis.
DAN|11|14|Et in temporibus illis multi consurgent adversus regem austri, filii quoque praevaricatorum populi tui extollentur, ut impleant visionem, et corruent.
DAN|11|15|Et veniet rex aquilonis et comportabit aggerem et capiet urbem munitissimam; et brachia austri non sustinebunt, et populo electorum eius non erit fortitudo ad resistendum.
DAN|11|16|Et faciet veniens super eum iuxta placitum suum, et non erit qui stet contra faciem eius; et stabit in terra inclita, et consumptio in manu eius.
DAN|11|17|Et ponet faciem suam, ut veniat ad tenendum universum regnum eius, et recta faciet cum eo et filiam feminarum dabit ei, ut evertat illud; et non stabit nec illius erit.
DAN|11|18|Et convertet faciem suam ad insulas et capiet multas, et cessare faciet princeps opprobrium eius, et opprobrium eius convertetur in eum.
DAN|11|19|Et convertet faciem suam ad oppida terrae suae et impinget et corruet, et non invenietur.
DAN|11|20|Et stabit in loco eius, qui mittat exactorem in decus regni; et in paucis diebus conteretur, non in furore nec in proelio.
DAN|11|21|Et stabit in loco eius despectus, et non tribuetur ei honor regius; et veniet clam et obtinebit regnum in fraudulentia.
DAN|11|22|Et brachia pugnantis expugnabuntur a facie eius et conterentur; insuper et dux foederis.
DAN|11|23|Et post amicitias, cum eo faciet dolum et ascendet et superabit in modico populo.
DAN|11|24|In prosperitate uberes urbes ingredietur et faciet, quae non fecerunt patres eius et patres patrum eius: rapinas et praedam et divitias eorum dissipabit et contra oppida cogitationes inibit, et hoc usque ad tempus.
DAN|11|25|Et concitabitur fortitudo eius et cor eius adversum regem austri in exercitu magno; et rex austri provocabitur ad bellum multis auxiliis et fortibus nimis, et non stabit, quia inibunt adversus eum consilia.
DAN|11|26|Et comedentes panem cum eo conterent illum; exercitusque eius opprimetur, et cadent interfecti plurimi.
DAN|11|27|Duorum quoque regum cor erit, ut malefaciant et ad mensam unam mendacium loquentur et non proficient, quia adhuc finis in aliud tempus.
DAN|11|28|Et revertetur in terram suam cum opibus multis, et cor eius adversum testamentum sanctum; et faciet et revertetur in terram suam.
DAN|11|29|Statuto tempore revertetur et veniet ad austrum, et non erit priori simile novissimum.
DAN|11|30|Et venient super eum trieres, Romani; et percutietur et revertetur et indignabitur contra testamentum sanctum et faciet reverteturque et cogitabit adversum eos, qui dereliquerunt testamentum sanctum.
DAN|11|31|Et brachia ex eo stabunt et polluent sanctuarium fortitudinis et auferent iuge sacrificium et dabunt abominationem vastatoris.
DAN|11|32|Et impios in testamentum errare faciet fraudulenter; populus autem scientium Deum suum obtinebit et faciet.
DAN|11|33|Et docti in populo docebunt plurimos; et ruent in gladio et in flamma et in captivitate et in rapina per dies.
DAN|11|34|Cumque corruerint, sublevabuntur auxilio parvulo, et applicabuntur eis plurimi fraudulenter.
DAN|11|35|Et de eruditis ruent, ut aliqui eorum conflentur et purgentur et dealbentur usque ad tempus praefinitum, quia adhuc aliud tempus erit.
DAN|11|36|Et faciet iuxta voluntatem suam rex et elevabitur et magnificabitur adversus omnem deum et adversus Deum deorum loquetur magnifica et prosperabitur, donec compleatur iracundia; perpetrata quippe est definitio.
DAN|11|37|Et deos patrum suorum non reputabit neque concupiscentiam feminarum nec quemquam deorum curabit, quia super universa magnificabit se;
DAN|11|38|deum autem oppidorum in loco suo venerabitur et deum, quem ignoraverunt patres eius, colet auro et argento et lapide pretioso rebusque pretiosis
DAN|11|39|et faciet adversus oppida munita cum deo alieno; qui cognoverit eum, multiplicabit gloriam eius et dabit eis potestatem in multis et terram dividet pretio.
DAN|11|40|Et in tempore praefinito proeliabitur adversus eum rex austri, et quasi tempestas veniet contra illum rex aquilonis in curribus et in equitibus et in classe magna, et ingredietur terras et conteret et pertransiet.
DAN|11|41|Et introibit in terram gloriosam, et multae corruent; hae autem solae salvabuntur de manu eius: Edom et Moab et principium filiorum Ammon.
DAN|11|42|Et mittet manum suam in terras, et terra Aegypti non effugiet;
DAN|11|43|et dominabitur thesaurorum auri et argenti et in omnibus pretiosis Aegypti, et Libyes et Aethiopes in vestigia eius transibunt.
DAN|11|44|Et fama turbabit eum ab oriente et ab aquilone; et veniet in ira magna, ut conterat et interficiat plurimos,
DAN|11|45|et figet tabernacula palatii sui inter maria super montem sanctum decoris; et veniet usque ad summitatem eius, et nemo auxiliabitur ei.
DAN|12|1|In tempore autem illo con surget Michael, princeps magnus, qui stat pro filiis populi tui, et erit tempus angustiae, quale non fuit ab eo, quo gentes esse coeperunt, usque ad tempus illud. Et in tempore illo salvabitur populus tuus, omnis, qui inventus fuerit scriptus in libro.
DAN|12|2|Et multi de his, qui dormiunt in terra pulveris, evigilabunt: alii in vitam aeternam, et alii in opprobrium sempiternum.
DAN|12|3|Qui autem docti fuerint, fulgebunt quasi splendor firmamenti; et, qui ad iustitiam erudierint multos, quasi stellae in perpetuas aeternitates.
DAN|12|4|Tu autem, Daniel, claude sermones et signa librum usque ad tempus finis; pertransibunt plurimi, et multiplex erit scientia ".
DAN|12|5|Et vidi ego Daniel: et ecce duo alii stabant, unus hinc super ripam fluminis, et alius inde ex altera ripa fluminis.
DAN|12|6|Et dixit viro, qui indutus erat lineis, qui stabat super aquas fluminis: Usquequo finis horum mirabilium? ".
DAN|12|7|Et audivi virum, qui indutus erat lineis, qui stabat super aquas fluminis, cum levasset dexteram et sinistram suam in caelum et iurasset per Viventem in aeternum: " Quia in tempus, tempora et dimidium temporis; et cum completa fuerit dispersio manus populi sancti, complebuntur universa haec ".
DAN|12|8|Et ego audivi et non intellexi et dixi: " Domine mi, quid erit finis horum? ".
DAN|12|9|Et ait: " Vade, Daniel, quia clausi sunt signatique sermones usque ad tempus praefinitum.
DAN|12|10|Purificabuntur et dealbabuntur et probabuntur multi, et impie agent impii, neque intellegent omnes impii; porro docti intellegent.
DAN|12|11|Et a tempore, cum ablatum fuerit iuge sacrificium, et posita fuerit abominatio vastatoris, dies mille ducenti nonaginta.
DAN|12|12|Beatus, qui exspectat et pervenit usque ad dies mille trecentos triginta quinque.
DAN|12|13|Tu autem vade ad finem et requiesce; et stabis in sorte tua in fine dierum ".Hucusque Daniel in Hebraeo volumine legimus. Cetera, quae sequuntur usque ad finem libri, de Theodotionis editione translata sunt).
DAN|13|1|Et erat vir habitans in Ba bylone, et nomen eius Ioa chim;
DAN|13|2|et accepit uxorem nomine Susannam, filiam Helciae, pulchram nimis et timentem Dominum;
DAN|13|3|parentes enim illius, cum essent iusti, erudierunt filiam suam secundum legem Moysis.
DAN|13|4|Erat autem Ioachim dives valde, et erat ei pomerium vicinum domui suae; et ad ipsum confluebant Iudaei, eo quod esset honorabilior omnium.
DAN|13|5|Et constituti sunt de populo duo senes iudices in anno illo, de quibus locutus est Dominus quia egressa est iniquitas de Babylone a senibus iudicibus, qui videbantur regere populum.
DAN|13|6|Isti frequentabant domum Ioachim, et veniebant ad eos omnes, qui habebant iudicia.
DAN|13|7|Cum autem populus revertisset per meridiem, ingrediebatur Susanna et deambulabat in pomerio viri sui.
DAN|13|8|Et videbant eam duo senes cotidie ingredientem et deambulantem et facti sunt in concupiscentia eius
DAN|13|9|et everterunt sensum suum et declinaverunt oculos suos, ut non viderent caelum neque recordarentur iudiciorum iustorum.
DAN|13|10|Erant ergo ambo vulnerati amore eius nec indicaverunt sibi vicissim dolorem suum;
DAN|13|11|erubescebant enim indicare concupiscentiam suam, volentes concumbere cum ea.
DAN|13|12|Et observabant cotidie sollicitius videre eam. Dixitque alter ad alterum:
DAN|13|13|" Eamus domum, quia prandi hora est ". Et egressi recesserunt a se.
DAN|13|14|Cumque revertissent, venerunt in unum et, sciscitantes ab invicem causam, confessi sunt concupiscentiam suam; et tunc in commune statuerunt tempus, quando eam possent invenire solam.
DAN|13|15|Factum est autem, cum observarent diem aptum, ingressa est aliquando sicut heri et nudiustertius cum duabus solis puellis voluitque lavari in pomerio, aestus quippe erat.
DAN|13|16|Et non erat ibi quisquam, praeter duos senes absconditos et contemplantes eam.
DAN|13|17|Dixit ergo puellis: " Afferte mihi oleum et smegmata et ostia pomerii claudite, ut laver ".
DAN|13|18|Et fecerunt, sicut praeceperat; clauseruntque ostia pomerii et egressae sunt per posticium, ut afferrent, quae iusserat; nesciebantque senes intus esse absconditos.
DAN|13|19|Cum autem egressae essent puellae, surrexerunt duo senes et accurrerunt ad eam et dixerunt:
DAN|13|20|" Ecce ostia pomerii clausa sunt, et nemo nos videt, et in concupiscentia tui sumus; quam ob rem assentire nobis et commiscere nobiscum.
DAN|13|21|Quod si nolueris, dicemus testimonium contra te, quod fuerit tecum iuvenis et ob hanc causam emiseris puellas a te ".
DAN|13|22|Ingemuit Susanna et ait: " Angustiae sunt mihi undique: si enim hoc egero, mors mihi est; si autem non egero, non effugiam manus vestras;
DAN|13|23|sed melius mihi est absque opere incidere in manus vestras quam peccare in conspectu Domini ".
DAN|13|24|Et exclamavit voce magna Susanna; exclamaverunt autem et senes adversus eam,
DAN|13|25|et, cum cucurrisset unus, aperuit ostia pomerii.
DAN|13|26|Cum ergo audissent clamorem in pomerio famuli domus, irruerunt per posticam, ut viderent quidnam esset ei.
DAN|13|27|Postquam autem senes locuti sunt sermones suos, erubuerunt servi vehementer, quia numquam dictus fuerat sermo huiuscemodi de Susanna. Et factum est die crastina,
DAN|13|28|cum venisset populus ad virum eius Ioachim, venerunt et duo presbyteri pleni iniqua cogitatione adversum Susannam, ut interficerent eam;
DAN|13|29|et dixerunt coram populo: " Mittite ad Susannam, filiam Helciae, quae est uxor Ioachim "; et miserunt.
DAN|13|30|Et venit cum parentibus et filiis et universis cognatis suis.
DAN|13|31|Porro Susanna erat delicata nimis et pulchra specie.
DAN|13|32|At iniqui illi iusserunt, ut discooperiretur - erat enim cooperta - ut satiarentur decore eius.
DAN|13|33|Flebant igitur sui et omnes, qui videbant eam.
DAN|13|34|Consurgentes autem duo presbyteri in medio populi, posuerunt manus super caput eius;
DAN|13|35|quae flens suspexit ad caelum: erat enim cor eius fiduciam habens in Domino.
DAN|13|36|Et dixerunt presbyteri: " Cum deambularemus in pomerio soli, ingressa est haec cum duabus puellis et clausit ostia pomerii et dimisit puellas;
DAN|13|37|venitque ad eam adulescens, qui erat absconditus, et concubuit cum ea.
DAN|13|38|Porro nos cum essemus in angulo pomerii, videntes iniquitatem cucurrimus ad eos et vidimus eos commisceri.
DAN|13|39|Et illum quidem non quivimus comprehendere, quia fortior nobis erat et, apertis ostiis, exilivit.
DAN|13|40|Hanc autem cum apprehendissemus, interrogavimus, quisnam esset adulescens, et noluit indicare nobis. Huius rei testes sumus ".
DAN|13|41|Credidit eis multitudo quasi senibus populi et iudicibus, et condemnaverunt eam ad mortem.
DAN|13|42|Exclamavit autem voce magna Susanna et dixit: " Deus aeterne, qui absconditorum es cognitor, qui nosti omnia antequam fiant,
DAN|13|43|tu scis quoniam falsum contra me tulerunt testimonium; et ecce morior, cum nihil horum fecerim, quae isti malitiose composuerunt adversum me ".
DAN|13|44|Exaudivit autem Dominus vocem eius.
DAN|13|45|Cumque duceretur ad mortem, suscitavit Deus spiritum sanctum pueri iunioris, cuius nomen Daniel;
DAN|13|46|et exclamavit voce magna: " Innocens ego sum a sanguine huius ".
DAN|13|47|Et conversus omnis populus ad eum dixit: " Quis est iste sermo, quem tu locutus es? ".
DAN|13|48|Qui cum staret in medio eorum, ait: " Sic fatui, filii Israel? Non iudicantes neque, quod verum est, cognoscentes, condemnastis filiam Israel!
DAN|13|49|Revertimini ad iudicium, quia falsum testimonium locuti sunt adversum eam ".
DAN|13|50|Reversus est ergo omnis populus cum festinatione, et dixerunt ei senes: Veni et sede in medio nostrum et indica nobis, quia tibi dedit Deus honorem senectutis ".
DAN|13|51|Et dixit ad eos Daniel: " Separate illos ab invicem procul, et diiudicabo eos ".
DAN|13|52|Cum ergo divisi essent alter ab altero, vocavit unum de eis et dixit ad eum: " Inveterate dierum malorum, nunc venerunt peccata tua, quae operabaris prius,
DAN|13|53|iudicans iudicia iniusta, innocentes opprimens et dimittens noxios, dicente Domino: "Innocentem et iustum non interficies".
DAN|13|54|Nunc ergo, si vidisti eam, dic sub qua arbore videris eos loquentes sibi ". Qui ait: " Sub schino ".
DAN|13|55|Dixit autem Daniel: " Recte mentitus es in caput tuum; ecce enim angelus Dei, accepta sententia a Deo, scindet te medium ".
DAN|13|56|Et amoto eo, iussit adduci alium et dixit ei: " Semen Chanaan et non Iudae, species decepit te, et concupiscentia subvertit cor tuum.
DAN|13|57|Sic faciebatis filiabus Israel, et illae timentes loquebantur vobis, sed non filia Iudae sustinuit iniquitatem vestram.
DAN|13|58|Nunc ergo dic mihi sub qua arbore comprehenderis eos colloquentes sibi.Qui ait: " Sub prino ".
DAN|13|59|Dixit autem ei Daniel: " Recte mentitus es et tu in caput tuum; manet enim angelus Dei, gladium habens, ut secet te medium et interficiat vos ".
DAN|13|60|Exclamavit itaque omnis coetus voce magna et benedixerunt Deo, qui salvat sperantes in se.
DAN|13|61|Et consurrexerunt adversum duos presbyteros - convicerat enim eos Daniel ex ore suo falsum dixisse testimonium - feceruntque eis, sicut male egerant adversum proximum,
DAN|13|62|ut facerent secundum legem Moysis; et interfecerunt eos, et salvatus est sanguis innoxius in die illa.
DAN|13|63|Helcias autem et uxor eius laudaverunt Deum pro filia sua Susanna, cum Ioachim marito eius et cognatis omnibus, quia non esset inventa in ea res turpis.
DAN|13|64|Daniel autem factus est magnus in conspectu populi a die illa et deinceps.
DAN|14|1|Et rex Astyages appositus est ad patres suos, et suscepit Cyrus Perses regnum eius.
DAN|14|2|Erat autem Daniel conviva regis et honoratus super omnes amicos eius.
DAN|14|3|Erat quoque idolum nomine Bel apud Babylonios, ct impendebantur in eo per dies singulos similae artabae duodecim et oves quadraginta vinique metretae sex.
DAN|14|4|Rex quoque colebat eum et ibat per singulos dies adorare eum; porro Daniel adorabat Deum suum. Dixitque ei rex: " Quare non adoras Bel? ".
DAN|14|5|Qui respondens ait ei: " Quia non colo idola manufacta sed viventem Deum, qui creavit caelum et terram et habet potestatem omnis carnis ".
DAN|14|6|Et dixit ad eum rex: "Non tibi videtur esse Bel vivens deus? An non vides, quanta comedat et bibat cotidie? ".
DAN|14|7|Et ait Daniel arridens: " Ne erres, rex; iste enim intrinsecus luteus est et forinsecus aereus, neque comedit neque bibit aliquando ".
DAN|14|8|Et iratus rex vocavit sacerdotes eius et ait eis: " Nisi dixeritis mihi, quis est qui comedat impensas has, moriemini;
DAN|14|9|si autem ostenderitis quoniam Bel comedat haec, morietur Daniel, quia blasphemavit in Bel ". Et dixit Daniel regi: " Fiat iuxta verbum tuum ".
DAN|14|10|Erant autem sacerdotes Bel septuaginta, exceptis uxoribus et parvulis et filiis. Et venit rex cum Daniele in templum Belis.
DAN|14|11|Et dixerunt sacerdotes Belis: " Ecce nos egredimur foras; et tu, rex, affer escas et vinum miscens pone et claude ostium et signa anulo tuo;
DAN|14|12|et, cum ingressus fueris mane, nisi inveneris omnia comesta a Bel, morte moriemur, vel Daniel, qui mentitus est adversum nos ".
DAN|14|13|Contemnebant autem, quia fecerant sub mensa absconditum introitum et per illum ingrediebantur semper et devorabant ea.
DAN|14|14|Factum est igitur, postquam egressi sunt illi, et rex posuit cibos ante Bel; et praecepit Daniel pueris suis, et attulerunt cinerem et cribraverunt per totum templum coram rege solo et egressi clauserunt ostium et signantes anulo regis abierunt.
DAN|14|15|Sacerdotes autem ingressi sunt nocte iuxta consuetudinem suam et uxores et filii eorum et comederunt omnia et biberunt.
DAN|14|16|Surrexit autem rex primo diluculo, et Daniel cum eo;
DAN|14|17|et ait rex: " Salvane sunt signa, Daniel? ". Qui respondit: " Salva, rex ".
DAN|14|18|Statimque cum aperuisset ostium, intuitus rex mensam, exclamavit voce magna: " Magnus es, Bel, et non est apud te dolus quisquam ".
DAN|14|19|Et risit Daniel et tenuit regem, ne ingrederetur intro, et dixit: " Ecce pavimentum; animadverte, cuius vestigia sunt haec ".
DAN|14|20|Et dixit rex: " Video vestigia virorum et mulierum et infantium ". Et iratus est rex.
DAN|14|21|Tunc apprehendit sacerdotes et uxores et filios eorum, et ostenderunt ei abscondita ostiola, per quae ingrediebantur et consumebant, quae erant super mensam.
DAN|14|22|Occidit ergo illos rex et tradidit Bel in potestate Danieli, qui subvertit eum et templum eius.
DAN|14|23|Et erat draco magnus, et colebant eum Babylonii.
DAN|14|24|Et dixit rex Danieli: " Non potes dicere quia iste non sit deus vivens; adora ergo eum ".
DAN|14|25|Dixitque Daniel: " Dominum Deum meum adoro, quia ipse est Deus vivens.
DAN|14|26|Tu autem, rex, da mihi potestatem, et interficiam draconem absque gladio et fuste ". Et ait rex: " Do tibi ".
DAN|14|27|Tulit ergo Daniel picem et adipem et pilos et coxit pariter; fecitque massas et dedit in os draconis et, cum comedisset, diruptus est draco. Et dixit: " Ecce quae colebatis ".
DAN|14|28|Cum audissent Babylonii, indignati sunt vehementer et congregati adversum regem dixerunt: "Iudaeus factus est rex; Bel destruxit, draconem interfecit et sacerdotes occidit ".
DAN|14|29|Et dixerunt, cum venissent ad regem: " Trade nobis Danielem; alioquin interficiemus te et domum tuam ".
DAN|14|30|Vidit ergo rex quod irruerent in eum vehementer et, necessitate compulsus, tradidit eis Danielem.
DAN|14|31|Qui miserunt eum in lacum leonum, et erat ibi diebus sex.
DAN|14|32|Porro in lacu erant septem leones, et dabantur eis cotidie duo corpora et duae oves; et tunc non data sunt eis, ut devorarent Danielem.
DAN|14|33|Erat autem Abacuc propheta in Iudaea et ipse coxerat pulmentum et intriverat panes in alveolo et ibat in campum, ut ferret messoribus.
DAN|14|34|Dixitque angelus Domini ad Abacuc: " Fer prandium, quod habes, in Babylonem Danieli, qui est in lacu leonum ".
DAN|14|35|Et dixit Abacuc: " Domine, Babylonem non vidi et lacum nescio ".
DAN|14|36|Et apprehendit eum angelus Domini in vertice eius et portavit eum capillo capitis sui posuitque eum in Babylone supra lacum in impetu spiritus sui.
DAN|14|37|Et clamavit Abacuc dicens: " Daniel, Daniel, tolle prandium, quod misit tibi Deus ".
DAN|14|38|Et ait Daniel: "Recordatus es enim mei, Deus, et non dereliquisti diligentes te ".
DAN|14|39|Surgensque Daniel comedit. Porro angelus Dei restituit Abacuc confestim in loco suo.
DAN|14|40|Venit ergo rex die septima, ut lugeret Danielem; et venit ad lacum et introspexit, et ecce Daniel sedens.
DAN|14|41|Et exclamavit rex voce magna dicens: "Magnus es, Domine, Deus Danielis, et non est alius praeter te ".
DAN|14|42|Porro illos, qui perditionis eius causa fuerant, intromisit in lacum; et devorati sunt in momento coram eo.
