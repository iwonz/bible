GAL|1|1|Paulus apostolus, non ab ho minibus neque per hominem, sed per Iesum Christum et Deum Patrem, qui suscitavit eum a mortuis,
GAL|1|2|et, qui mecum sunt, omnes fratres ecclesiis Galatiae:
GAL|1|3|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo,
GAL|1|4|qui dedit semetipsum pro peccatis nostris, ut eriperet nos de praesenti saeculo nequam secundum voluntatem Dei et Patris nostri,
GAL|1|5|cui gloria in saecula saeculorum. Amen.
GAL|1|6|Miror quod tam cito transferimini ab eo, qui vos vocavit in gratia Christi, in aliud evangelium;
GAL|1|7|quod non est aliud, nisi sunt aliqui, qui vos conturbant et volunt convertere evangelium Christi.
GAL|1|8|Sed licet nos aut angelus de caelo evangelizet vobis praeterquam quod evangelizavimus vobis, anathema sit!
GAL|1|9|Sicut praediximus, et nunc iterum dico: Si quis vobis evangelizaverit praeter id, quod accepistis, anathema sit!
GAL|1|10|Modo enim hominibus suadeo aut Deo? Aut quaero hominibus placere? Si adhuc hominibus placerem, Christi servus non essem!
GAL|1|11|Notum enim vobis facio, fratres, evangelium, quod evangelizatum est a me, quia non est secundum hominem;
GAL|1|12|neque enim ego ab homine accepi illud neque didici sed per revelationem Iesu Christi.
GAL|1|13|Audistis enim conversationem meam aliquando in Iudaismo, quoniam supra modum persequebar ecclesiam Dei et expugnabam illam;
GAL|1|14|et proficiebam in Iudaismo supra multos coaetaneos in genere meo, abundantius aemulator exsistens paternarum mearum traditionum.
GAL|1|15|Cum autem placuit Deo, qui me segregavit de utero matris meae et vocavit per gratiam suam,
GAL|1|16|ut revelaret Filium suum in me, ut evangelizarem illum in gentibus, continuo non contuli cum carne et sanguine
GAL|1|17|neque ascendi Hierosolymam ad antecessores meos apostolos; sed abii in Arabiam et iterum reversus sum Damascum.
GAL|1|18|Deinde post annos tres, ascendi Hierosolymam videre Cepham et mansi apud eum diebus quindecim;
GAL|1|19|alium autem apostolorum non vidi, nisi Iacobum fratrem Domini.
GAL|1|20|Quae autem scribo vobis, ecce coram Deo quia non mentior.
GAL|1|21|Deinde veni in partes Syriae et Ciliciae.
GAL|1|22|Eram autem ignotus facie ecclesiis Iudaeae, quae sunt in Christo;
GAL|1|23|tantum autem auditum habebant: " Qui persequebatur nos aliquando, nunc evangelizat fidem, quam aliquando expugnabat ",
GAL|1|24|et in me glorificabant Deum.
GAL|2|1|Deinde post annos quattuor decim, iterum ascendi Hieroso lymam cum Barnaba, assumpto et Tito;
GAL|2|2|ascendi autem secundum revelationem; et contuli cum illis evangelium, quod praedico in gentibus, seorsum autem his, qui observabantur, ne forte in vacuum currerem aut cucurrissem.
GAL|2|3|Sed neque Titus, qui mecum erat, cum esset Graecus, compulsus est circumcidi.
GAL|2|4|Sed propter subintroductos falsos fratres, qui subintroierunt explorare libertatem nostram, quam habemus in Christo Iesu, ut nos in servitutem redigerent;
GAL|2|5|quibus neque ad horam cessimus subicientes nos, ut veritas evangelii permaneat apud vos.
GAL|2|6|Ab his autem, qui videbantur esse aliquid - quales aliquando fuerint, nihil mea interest; Deus personam hominis non accipit - mihi enim, qui observabantur, nihil contulerunt,
GAL|2|7|sed e contra, cum vidissent quod creditum est mihi evangelium praeputii, sicut Petro circumcisionis
GAL|2|8|- qui enim operatus est Petro in apostolatum circumcisionis, operatus est et mihi inter gentes -
GAL|2|9|et cum cognovissent gratiam, quae data est mihi, Iacobus et Cephas et Ioannes, qui videbantur columnae esse, dexteras dederunt mihi et Barnabae communionis, ut nos in gentes, ipsi autem in circumcisionem;
GAL|2|10|tantum ut pauperum memores essemus, quod etiam sollicitus fui hoc ipsum facere.
GAL|2|11|Cum autem venisset Cephas Antiochiam, in faciem ei restiti, quia reprehensibilis erat.
GAL|2|12|Prius enim quam venirent quidam ab Iacobo, cum gentibus comedebat; cum autem venissent, subtrahebat et segregabat se, timens eos, qui ex circumcisione erant.
GAL|2|13|Et simulationi eius consenserunt ceteri Iudaei, ita ut et Barnabas simul abduceretur illorum simulatione.
GAL|2|14|Sed cum vidissem quod non recte ambularent ad veritatem evangelii, dixi Cephae coram omnibus: " Si tu, cum Iudaeus sis, gentiliter et non Iudaice vivis, quomodo gentes cogis iudaizare? ".
GAL|2|15|Nos natura Iudaei et non ex gentibus peccatores,
GAL|2|16|scientes autem quod non iustificatur homo ex operibus legis, nisi per fidem Iesu Christi, et nos in Christum Iesum credidimus, ut iustificemur ex fide Christi et non ex operibus legis, quoniam ex operibus legis non iustificabitur omnis caro.
GAL|2|17|Quodsi quaerentes iustificari in Christo, inventi sumus et ipsi peccatores, numquid Christus peccati minister est? Absit!
GAL|2|18|Si enim, quae destruxi, haec iterum aedifico, praevaricatorem me constituo.
GAL|2|19|Ego enim per legem legi mortuus sum, ut Deo vivam. Christo confixus sum cruci;
GAL|2|20|vivo autem iam non ego, vivit vero in me Christus; quod autem nunc vivo in carne, in fide vivo Filii Dei, qui dilexit me et tradidit seipsum pro me.
GAL|2|21|Non irritam facio gratiam Dei; si enim per legem iustitia, ergo Christus gratis mortuus est.
GAL|3|1|O insensati Galatae, quis vos fascinavit, ante quorum oculos Iesus Christus descriptus est crucifixus?
GAL|3|2|Hoc solum volo a vobis discere: Ex operibus legis Spiritum accepistis an ex auditu fidei?
GAL|3|3|Sic stulti estis? Cum Spiritu coeperitis, nunc carne consummamini?
GAL|3|4|Tanta passi estis sine causa? Si tamen et sine causa!
GAL|3|5|Qui ergo tribuit vobis Spiritum et operatur virtutes in vobis, ex operibus legis an ex auditu fidei?
GAL|3|6|Sicut Abraham credidit Deo, et reputatum est ei ad iustitiam.
GAL|3|7|Cognoscitis ergo quia qui ex fide sunt, hi sunt filii Abrahae.
GAL|3|8|Providens autem Scriptura, quia ex fide iustificat gentes Deus, praenuntiavit Abrahae: "Benedicentur in te omnes gentes".
GAL|3|9|Igitur, qui ex fide sunt, benedi cuntur cum fideli Abraham.
GAL|3|10|Quicumque enim ex operibus legis sunt, sub maledicto sunt; scriptum est enim: " Maledictus omnis, qui non permanserit in omnibus, quae scripta sunt in libro legis, ut faciat ea ".
GAL|3|11|Quoniam autem in lege nemo iustificatur apud Deum manifestum est, quia iustus ex fide vivet;
GAL|3|12|lex autem non est ex fide; sed, qui fecerit ea, vivet in illis.
GAL|3|13|Christus nos redemit de maledicto legis factus pro nobis maledictum, quia scriptum est: " Maledictus omnis, qui pendet in ligno ",
GAL|3|14|ut in gentes benedictio Abrahae fieret in Christo Iesu, ut promissionem Spiritus accipiamus per fidem.
GAL|3|15|Fratres, secundum hominem dico, tamen hominis confirmatum testamentum nemo irritum facit aut superordinat.
GAL|3|16|Abrahae autem dictae sunt promissiones et semini eius. Non dicit: " Et seminibus ", quasi in multis, sed quasi in uno: "Et semini tuo", qui est Christus.
GAL|3|17|Hoc autem dico: Testamentum confirmatum a Deo, quae post quadringentos et triginta annos facta est lex, non irritum facit ad evacuandam promissionem.
GAL|3|18|Nam si ex lege hereditas, iam non ex promissione; Abrahae autem per promissionem donavit Deus.
GAL|3|19|Quid igitur lex? Propter transgressiones apposita est, donec veniret semen, cui promissum est, ordinata per angelos in manu mediatoris.
GAL|3|20|Mediator autem unius non est, Deus autem unus est.
GAL|3|21|Lex ergo adversus promissa Dei? Absit. Si enim data esset lex, quae posset vivificare, vere ex lege esset iustitia.
GAL|3|22|Sed conclusit Scriptura omnia sub peccato, ut promissio ex fide Iesu Christi daretur credentibus.
GAL|3|23|Prius autem quam veniret fides, sub lege custodiebamur conclusi in eam fidem, quae revelanda erat.
GAL|3|24|Itaque lex paedagogus noster fuit in Christum, ut ex fide iustificemur;
GAL|3|25|at ubi venit fides, iam non sumus sub paedagogo.
GAL|3|26|Omnes enim filii Dei estis per fidem in Christo Iesu.
GAL|3|27|Quicumque enim in Christum baptizati estis, Christum induistis:
GAL|3|28|non est Iudaeus neque Graecus, non est servus neque liber, non est masculus et femina; omnes enim vos unus estis in Christo Iesu.
GAL|3|29|Si autem vos Christi, ergo Abrahae semen estis, secundum promissionem heredes.
GAL|4|1|Dico autem: Quanto tempore heres parvulus est, nihil differt a servo, cum sit dominus omnium,
GAL|4|2|sed sub tutoribus est et actoribus usque ad praefinitum tempus a patre.
GAL|4|3|Ita et nos, cum essemus parvuli, sub elementis mundi eramus servientes;
GAL|4|4|at ubi venit plenitudo temporis, misit Deus Filium suum, factum ex muliere, factum sub lege,
GAL|4|5|ut eos, qui sub lege erant, redimeret, ut adoptionem filiorum reciperemus.
GAL|4|6|Quoniam autem estis filii, misit Deus Spiritum Filii sui in corda nostra clamantem: " Abba, Pater! ".
GAL|4|7|Itaque iam non es servus sed filius; quod si filius, et heres per Deum.
GAL|4|8|Sed tunc quidem ignorantes Deum, his, qui natura non sunt dii, servistis;
GAL|4|9|nunc autem, cum cognoveritis Deum, immo cogniti sitis a Deo, quomodo convertimini iterum ad infirma et egena elementa, quibus rursus ut antea servire vultis?
GAL|4|10|Dies observatis et menses et tempora et annos!
GAL|4|11|Timeo vos, ne forte sine causa laboraverim in vobis.
GAL|4|12|Estote sicut ego, quia et ego sicut vos; fratres, obsecro vos. Nihil me laesistis;
GAL|4|13|scitis autem quia per infirmitatem carnis pridem vobis evangelizavi,
GAL|4|14|et tentationem vestram in carne mea non sprevistis neque respuistis, sed sicut angelum Dei excepistis me, sicut Christum Iesum.
GAL|4|15|Ubi est ergo beatitudo vestra? Testimonium enim perhibeo vobis, quia, si fieri posset, oculos vestros eruissetis et dedissetis mihi.
GAL|4|16|Ergo inimicus vobis factus sum, verum dicens vobis?
GAL|4|17|Aemulantur vos non bene, sed excludere vos volunt, ut illos aemulemini.
GAL|4|18|Bonum est autem aemulari in bono semper, et non tantum cum praesens sum apud vos,
GAL|4|19|filioli mei, quos iterum parturio, donec formetur Christus in vobis!
GAL|4|20|Vellem autem esse apud vos modo et mutare vocem meam, quoniam incertus sum in vobis.
GAL|4|21|Dicite mihi, qui sub lege vultis esse: Legem non auditis?
GAL|4|22|Scriptum est enim quoniam Abraham duos filios habuit, unum de ancilla et unum de libera.
GAL|4|23|Sed qui de ancilla, secundum carnem natus est; qui autem de libera, per promissionem.
GAL|4|24|Quae sunt per allegoriam dicta; ipsae enim sunt duo Testamenta, unum quidem a monte Sinai, in servitutem generans, quod est Agar.
GAL|4|25|Illud vero Agar mons est Sinai in Arabia, respondet autem Ierusalem, quae nunc est; servit enim cum filiis suis.
GAL|4|26|Illa autem, quae sursum est Ierusalem, libera est, quae est mater nostra;
GAL|4|27|scriptum est enim: Laetare, sterilis, quae non paris,erumpe et exclama, quae non parturis,quia multi filii desertaemagis quam eius, quae habet virum ".
GAL|4|28|Vos autem, fratres, secundum Isaac promissionis filii estis.
GAL|4|29|Sed quomodo tunc, qui secundum carnem natus fuerat, persequebatur eum, qui secundum spiritum, ita et nunc.
GAL|4|30|Sed quid dicit Scriptura? " Eice ancillam et filium eius; non enim heres erit filius ancillae cum filio liberae ".
GAL|4|31|Itaque, fratres, non sumus ancillae filii sed liberae.
GAL|5|1|Hac libertate nos Christus liberavit; state igitur et nolite iterum iugo servitutis detineri.
GAL|5|2|Ecce ego Paulus dico vobis quoniam, si circumcidamini, Christus vobis nihil proderit.
GAL|5|3|Testificor autem rursum omni homini circumcidenti se quoniam debitor est universae legis faciendae.
GAL|5|4|Evacuati estis a Christo, qui in lege iustificamini, a gratia excidistis.
GAL|5|5|Nos enim Spiritu ex fide spem iustitiae exspectamus.
GAL|5|6|Nam in Christo Iesu neque circumcisio aliquid valet neque praeputium, sed fides, quae per caritatem operatur.
GAL|5|7|Currebatis bene; quis vos impedivit veritati non oboedire?
GAL|5|8|Haec persuasio non est ex eo, qui vocat vos.
GAL|5|9|Modicum fermentum totam massam corrumpit.
GAL|5|10|Ego confido in vobis in Domino, quod nihil aliud sapietis; qui autem conturbat vos, portabit iudicium, quicumque est ille.
GAL|5|11|Ego autem, fratres, si circumcisionem adhuc praedico, quid adhuc persecutionem patior? Ergo evacuatum est scandalum crucis.
GAL|5|12|Utinam et abscidantur, qui vos conturbant!
GAL|5|13|Vos enim in libertatem vocati estis, fratres; tantum ne libertatem in occasionem detis carni, sed per caritatem servite invicem.
GAL|5|14|Omnis enim lex in uno sermone impletur, in hoc: Diliges proximum tuum sicut teipsum.
GAL|5|15|Quod si invicem mordetis et devoratis, videte, ne ab invicem consumamini!
GAL|5|16|Dico autem: Spiritu ambulate et concupiscentiam carnis ne perfeceritis.
GAL|5|17|Caro enim concupiscit adversus Spiritum, Spiritus autem adversus carnem; haec enim invicem adversantur, ut non, quaecumque vultis, illa faciatis.
GAL|5|18|Quod si Spiritu ducimini, non estis sub lege.
GAL|5|19|Manifesta autem sunt opera carnis, quae sunt fornicatio, immunditia, luxuria,
GAL|5|20|idolorum servitus, veneficia, inimicitiae, contentiones, aemulationes, irae, rixae, dissensiones, sectae,
GAL|5|21|invidiae, ebrietates, comissationes et his similia; quae praedico vobis, sicut praedixi, quoniam, qui talia agunt, regnum Dei non consequentur.
GAL|5|22|Fructus autem Spiritus est caritas, gaudium, pax, longanimitas, benignitas, bonitas, fides,
GAL|5|23|mansuetudo, continentia; adversus huiusmodi non est lex.
GAL|5|24|Qui autem sunt Christi Iesu, carnem crucifixerunt cum vitiis et concupiscentiis.
GAL|5|25|Si vivimus Spiritu, Spiritu et ambulemus.
GAL|5|26|Non efficiamur inanis gloriae cupidi, invicem provocantes, invicem invidentes.
GAL|6|1|Fratres, et si praeoccupatus fuerit homo in aliquo delicto, vos, qui spiritales estis, huiusmodi instruite in spiritu lenitatis, considerans teipsum, ne et tu tenteris.
GAL|6|2|Alter alterius onera portate et sic adimplebitis legem Christi.
GAL|6|3|Nam si quis existimat se aliquid esse, cum sit nihil, ipse se seducit;
GAL|6|4|opus autem suum probet unusquisque et sic in semetipso tantum gloriationem habebit et non in altero.
GAL|6|5|Unusquisque enim onus suum portabit.
GAL|6|6|Communicet autem is, qui catechizatur verbum, ei qui se catechizat, in omnibus bonis.
GAL|6|7|Nolite errare: Deus non irridetur. Quae enim seminaverit homo, haec et metet;
GAL|6|8|quoniam, qui seminat in carne sua, de carne metet corruptionem; qui autem seminat in Spiritu, de Spiritu metet vitam aeternam.
GAL|6|9|Bonum autem facientes infatigabiles, tempore enim suo metemus non deficientes.
GAL|6|10|Ergo dum tempus habemus, operemur bonum ad omnes, maxime autem ad domesticos fidei.
GAL|6|11|Videte qualibus litteris scripsi vobis mea manu.
GAL|6|12|Quicumque volunt placere in carne, hi cogunt vos circumcidi, tantum ut crucis Christi persecutionem non patiantur;
GAL|6|13|neque enim, qui circumciduntur, legem custodiunt, sed volunt vos circumcidi, ut in carne vestra glorientur.
GAL|6|14|Mihi autem absit gloriari, nisi in cruce Domini nostri Iesu Christi, per quem mihi mundus crucifixus est, et ego mundo.
GAL|6|15|Neque enim circumcisio aliquid est neque praeputium sed nova creatura.
GAL|6|16|Et quicumque hanc regulam secuti fuerint, pax super illos et misericordia et super Israel Dei.
GAL|6|17|De cetero nemo mihi molestus sit; ego enim stigmata Iesu in super corpore meo porto.
GAL|6|18|Gratia Domini nostri Iesu Christi cum spiritu vestro, fratres. Amen.
