GEN|1|1|in principio creavit Deus caelum et terram
GEN|1|2|terra autem erat inanis et vacua et tenebrae super faciem abyssi et spiritus Dei ferebatur super aquas
GEN|1|3|dixitque Deus fiat lux et facta est lux
GEN|1|4|et vidit Deus lucem quod esset bona et divisit lucem ac tenebras
GEN|1|5|appellavitque lucem diem et tenebras noctem factumque est vespere et mane dies unus
GEN|1|6|dixit quoque Deus fiat firmamentum in medio aquarum et dividat aquas ab aquis
GEN|1|7|et fecit Deus firmamentum divisitque aquas quae erant sub firmamento ab his quae erant super firmamentum et factum est ita
GEN|1|8|vocavitque Deus firmamentum caelum et factum est vespere et mane dies secundus
GEN|1|9|dixit vero Deus congregentur aquae quae sub caelo sunt in locum unum et appareat arida factumque est ita
GEN|1|10|et vocavit Deus aridam terram congregationesque aquarum appellavit maria et vidit Deus quod esset bonum
GEN|1|11|et ait germinet terra herbam virentem et facientem semen et lignum pomiferum faciens fructum iuxta genus suum cuius semen in semet ipso sit super terram et factum est ita
GEN|1|12|et protulit terra herbam virentem et adferentem semen iuxta genus suum lignumque faciens fructum et habens unumquodque sementem secundum speciem suam et vidit Deus quod esset bonum
GEN|1|13|factumque est vespere et mane dies tertius
GEN|1|14|dixit autem Deus fiant luminaria in firmamento caeli ut dividant diem ac noctem et sint in signa et tempora et dies et annos
GEN|1|15|ut luceant in firmamento caeli et inluminent terram et factum est ita
GEN|1|16|fecitque Deus duo magna luminaria luminare maius ut praeesset diei et luminare minus ut praeesset nocti et stellas
GEN|1|17|et posuit eas in firmamento caeli ut lucerent super terram
GEN|1|18|et praeessent diei ac nocti et dividerent lucem ac tenebras et vidit Deus quod esset bonum
GEN|1|19|et factum est vespere et mane dies quartus
GEN|1|20|dixit etiam Deus producant aquae reptile animae viventis et volatile super terram sub firmamento caeli
GEN|1|21|creavitque Deus cete grandia et omnem animam viventem atque motabilem quam produxerant aquae in species suas et omne volatile secundum genus suum et vidit Deus quod esset bonum
GEN|1|22|benedixitque eis dicens crescite et multiplicamini et replete aquas maris avesque multiplicentur super terram
GEN|1|23|et factum est vespere et mane dies quintus
GEN|1|24|dixit quoque Deus producat terra animam viventem in genere suo iumenta et reptilia et bestias terrae secundum species suas factumque est ita
GEN|1|25|et fecit Deus bestias terrae iuxta species suas et iumenta et omne reptile terrae in genere suo et vidit Deus quod esset bonum
GEN|1|26|et ait faciamus hominem ad imaginem et similitudinem nostram et praesit piscibus maris et volatilibus caeli et bestiis universaeque terrae omnique reptili quod movetur in terra
GEN|1|27|et creavit Deus hominem ad imaginem suam ad imaginem Dei creavit illum masculum et feminam creavit eos
GEN|1|28|benedixitque illis Deus et ait crescite et multiplicamini et replete terram et subicite eam et dominamini piscibus maris et volatilibus caeli et universis animantibus quae moventur super terram
GEN|1|29|dixitque Deus ecce dedi vobis omnem herbam adferentem semen super terram et universa ligna quae habent in semet ipsis sementem generis sui ut sint vobis in escam
GEN|1|30|et cunctis animantibus terrae omnique volucri caeli et universis quae moventur in terra et in quibus est anima vivens ut habeant ad vescendum et factum est ita
GEN|1|31|viditque Deus cuncta quae fecit et erant valde bona et factum est vespere et mane dies sextus
GEN|2|1|igitur perfecti sunt caeli et terra et omnis ornatus eorum
GEN|2|2|conplevitque Deus die septimo opus suum quod fecerat et requievit die septimo ab universo opere quod patrarat
GEN|2|3|et benedixit diei septimo et sanctificavit illum quia in ipso cessaverat ab omni opere suo quod creavit Deus ut faceret
GEN|2|4|istae generationes caeli et terrae quando creatae sunt in die quo fecit Dominus Deus caelum et terram
GEN|2|5|et omne virgultum agri antequam oreretur in terra omnemque herbam regionis priusquam germinaret non enim pluerat Dominus Deus super terram et homo non erat qui operaretur terram
GEN|2|6|sed fons ascendebat e terra inrigans universam superficiem terrae
GEN|2|7|formavit igitur Dominus Deus hominem de limo terrae et inspiravit in faciem eius spiraculum vitae et factus est homo in animam viventem
GEN|2|8|plantaverat autem Dominus Deus paradisum voluptatis a principio in quo posuit hominem quem formaverat
GEN|2|9|produxitque Dominus Deus de humo omne lignum pulchrum visu et ad vescendum suave lignum etiam vitae in medio paradisi lignumque scientiae boni et mali
GEN|2|10|et fluvius egrediebatur de loco voluptatis ad inrigandum paradisum qui inde dividitur in quattuor capita
GEN|2|11|nomen uni Phison ipse est qui circuit omnem terram Evilat ubi nascitur aurum
GEN|2|12|et aurum terrae illius optimum est ibique invenitur bdellium et lapis onychinus
GEN|2|13|et nomen fluvio secundo Geon ipse est qui circuit omnem terram Aethiopiae
GEN|2|14|nomen vero fluminis tertii Tigris ipse vadit contra Assyrios fluvius autem quartus ipse est Eufrates
GEN|2|15|tulit ergo Dominus Deus hominem et posuit eum in paradiso voluptatis ut operaretur et custodiret illum
GEN|2|16|praecepitque ei dicens ex omni ligno paradisi comede
GEN|2|17|de ligno autem scientiae boni et mali ne comedas in quocumque enim die comederis ex eo morte morieris
GEN|2|18|dixit quoque Dominus Deus non est bonum esse hominem solum faciamus ei adiutorium similem sui
GEN|2|19|formatis igitur Dominus Deus de humo cunctis animantibus terrae et universis volatilibus caeli adduxit ea ad Adam ut videret quid vocaret ea omne enim quod vocavit Adam animae viventis ipsum est nomen eius
GEN|2|20|appellavitque Adam nominibus suis cuncta animantia et universa volatilia caeli et omnes bestias terrae Adam vero non inveniebatur adiutor similis eius
GEN|2|21|inmisit ergo Dominus Deus soporem in Adam cumque obdormisset tulit unam de costis eius et replevit carnem pro ea
GEN|2|22|et aedificavit Dominus Deus costam quam tulerat de Adam in mulierem et adduxit eam ad Adam
GEN|2|23|dixitque Adam hoc nunc os ex ossibus meis et caro de carne mea haec vocabitur virago quoniam de viro sumpta est
GEN|2|24|quam ob rem relinquet homo patrem suum et matrem et adherebit uxori suae et erunt duo in carne una
GEN|2|25|erant autem uterque nudi Adam scilicet et uxor eius et non erubescebant
GEN|3|1|sed et serpens erat callidior cunctis animantibus terrae quae fecerat Dominus Deus qui dixit ad mulierem cur praecepit vobis Deus ut non comederetis de omni ligno paradisi
GEN|3|2|cui respondit mulier de fructu lignorum quae sunt in paradiso vescemur
GEN|3|3|de fructu vero ligni quod est in medio paradisi praecepit nobis Deus ne comederemus et ne tangeremus illud ne forte moriamur
GEN|3|4|dixit autem serpens ad mulierem nequaquam morte moriemini
GEN|3|5|scit enim Deus quod in quocumque die comederitis ex eo aperientur oculi vestri et eritis sicut dii scientes bonum et malum
GEN|3|6|vidit igitur mulier quod bonum esset lignum ad vescendum et pulchrum oculis aspectuque delectabile et tulit de fructu illius et comedit deditque viro suo qui comedit
GEN|3|7|et aperti sunt oculi amborum cumque cognovissent esse se nudos consuerunt folia ficus et fecerunt sibi perizomata
GEN|3|8|et cum audissent vocem Domini Dei deambulantis in paradiso ad auram post meridiem abscondit se Adam et uxor eius a facie Domini Dei in medio ligni paradisi
GEN|3|9|vocavitque Dominus Deus Adam et dixit ei ubi es
GEN|3|10|qui ait vocem tuam audivi in paradiso et timui eo quod nudus essem et abscondi me
GEN|3|11|cui dixit quis enim indicavit tibi quod nudus esses nisi quod ex ligno de quo tibi praeceperam ne comederes comedisti
GEN|3|12|dixitque Adam mulier quam dedisti sociam mihi dedit mihi de ligno et comedi
GEN|3|13|et dixit Dominus Deus ad mulierem quare hoc fecisti quae respondit serpens decepit me et comedi
GEN|3|14|et ait Dominus Deus ad serpentem quia fecisti hoc maledictus es inter omnia animantia et bestias terrae super pectus tuum gradieris et terram comedes cunctis diebus vitae tuae
GEN|3|15|inimicitias ponam inter te et mulierem et semen tuum et semen illius ipsa conteret caput tuum et tu insidiaberis calcaneo eius
GEN|3|16|mulieri quoque dixit multiplicabo aerumnas tuas et conceptus tuos in dolore paries filios et sub viri potestate eris et ipse dominabitur tui
GEN|3|17|ad Adam vero dixit quia audisti vocem uxoris tuae et comedisti de ligno ex quo praeceperam tibi ne comederes maledicta terra in opere tuo in laboribus comedes eam cunctis diebus vitae tuae
GEN|3|18|spinas et tribulos germinabit tibi et comedes herbas terrae
GEN|3|19|in sudore vultus tui vesceris pane donec revertaris in terram de qua sumptus es quia pulvis es et in pulverem reverteris
GEN|3|20|et vocavit Adam nomen uxoris suae Hava eo quod mater esset cunctorum viventium
GEN|3|21|fecit quoque Dominus Deus Adam et uxori eius tunicas pellicias et induit eos
GEN|3|22|et ait ecce Adam factus est quasi unus ex nobis sciens bonum et malum nunc ergo ne forte mittat manum suam et sumat etiam de ligno vitae et comedat et vivat in aeternum
GEN|3|23|emisit eum Dominus Deus de paradiso voluptatis ut operaretur terram de qua sumptus est
GEN|3|24|eiecitque Adam et conlocavit ante paradisum voluptatis cherubin et flammeum gladium atque versatilem ad custodiendam viam ligni vitae
GEN|4|1|Adam vero cognovit Havam uxorem suam quae concepit et peperit Cain dicens possedi hominem per Dominum
GEN|4|2|rursusque peperit fratrem eius Abel fuit autem Abel pastor ovium et Cain agricola
GEN|4|3|factum est autem post multos dies ut offerret Cain de fructibus terrae munera Domino
GEN|4|4|Abel quoque obtulit de primogenitis gregis sui et de adipibus eorum et respexit Dominus ad Abel et ad munera eius
GEN|4|5|ad Cain vero et ad munera illius non respexit iratusque est Cain vehementer et concidit vultus eius
GEN|4|6|dixitque Dominus ad eum quare maestus es et cur concidit facies tua
GEN|4|7|nonne si bene egeris recipies sin autem male statim in foribus peccatum aderit sed sub te erit appetitus eius et tu dominaberis illius
GEN|4|8|dixitque Cain ad Abel fratrem suum egrediamur foras cumque essent in agro consurrexit Cain adversus Abel fratrem suum et interfecit eum
GEN|4|9|et ait Dominus ad Cain ubi est Abel frater tuus qui respondit nescio num custos fratris mei sum
GEN|4|10|dixitque ad eum quid fecisti vox sanguinis fratris tui clamat ad me de terra
GEN|4|11|nunc igitur maledictus eris super terram quae aperuit os suum et suscepit sanguinem fratris tui de manu tua
GEN|4|12|cum operatus fueris eam non dabit tibi fructus suos vagus et profugus eris super terram
GEN|4|13|dixitque Cain ad Dominum maior est iniquitas mea quam ut veniam merear
GEN|4|14|ecce eicis me hodie a facie terrae et a facie tua abscondar et ero vagus et profugus in terra omnis igitur qui invenerit me occidet me
GEN|4|15|dixitque ei Dominus nequaquam ita fiet sed omnis qui occiderit Cain septuplum punietur posuitque Dominus Cain signum ut non eum interficeret omnis qui invenisset eum
GEN|4|16|egressusque Cain a facie Domini habitavit in terra profugus ad orientalem plagam Eden
GEN|4|17|cognovit autem Cain uxorem suam quae concepit et peperit Enoch et aedificavit civitatem vocavitque nomen eius ex nomine filii sui Enoch
GEN|4|18|porro Enoch genuit Irad et Irad genuit Maviahel et Maviahel genuit Matusahel et Matusahel genuit Lamech
GEN|4|19|qui accepit uxores duas nomen uni Ada et nomen alteri Sella
GEN|4|20|genuitque Ada Iabel qui fuit pater habitantium in tentoriis atque pastorum
GEN|4|21|et nomen fratris eius Iubal ipse fuit pater canentium cithara et organo
GEN|4|22|Sella quoque genuit Thubalcain qui fuit malleator et faber in cuncta opera aeris et ferri soror vero Thubalcain Noemma
GEN|4|23|dixitque Lamech uxoribus suis Adae et Sellae audite vocem meam uxores Lamech auscultate sermonem meum quoniam occidi virum in vulnus meum et adulescentulum in livorem meum
GEN|4|24|septuplum ultio dabitur de Cain de Lamech vero septuagies septies
GEN|4|25|cognovit quoque adhuc Adam uxorem suam et peperit filium vocavitque nomen eius Seth dicens posuit mihi Deus semen aliud pro Abel quem occidit Cain
GEN|4|26|sed et Seth natus est filius quem vocavit Enos iste coepit invocare nomen Domini
GEN|5|1|hic est liber generationis Adam in die qua creavit Deus hominem ad similitudinem Dei fecit illum
GEN|5|2|masculum et feminam creavit eos et benedixit illis et vocavit nomen eorum Adam in die qua creati sunt
GEN|5|3|vixit autem Adam centum triginta annis et genuit ad similitudinem et imaginem suam vocavitque nomen eius Seth
GEN|5|4|et facti sunt dies Adam postquam genuit Seth octingenti anni genuitque filios et filias
GEN|5|5|et factum est omne tempus quod vixit Adam anni nongenti triginta et mortuus est
GEN|5|6|vixit quoque Seth centum quinque annos et genuit Enos
GEN|5|7|vixitque Seth postquam genuit Enos octingentis septem annis genuitque filios et filias
GEN|5|8|et facti sunt omnes dies Seth nongentorum duodecim annorum et mortuus est
GEN|5|9|vixit vero Enos nonaginta annis et genuit Cainan
GEN|5|10|post cuius ortum vixit octingentis quindecim annis et genuit filios et filias
GEN|5|11|factique sunt omnes dies Enos nongentorum quinque annorum et mortuus est
GEN|5|12|vixit quoque Cainan septuaginta annis et genuit Malalehel
GEN|5|13|et vixit Cainan postquam genuit Malalehel octingentos quadraginta annos genuitque filios et filias
GEN|5|14|et facti sunt omnes dies Cainan nongenti decem anni et mortuus est
GEN|5|15|vixit autem Malalehel sexaginta quinque annos et genuit Iared
GEN|5|16|et vixit Malalehel postquam genuit Iared octingentis triginta annis et genuit filios et filias
GEN|5|17|et facti sunt omnes dies Malalehel octingenti nonaginta quinque anni et mortuus est
GEN|5|18|vixitque Iared centum sexaginta duobus annis et genuit Enoch
GEN|5|19|et vixit Iared postquam genuit Enoch octingentos annos et genuit filios et filias
GEN|5|20|et facti sunt omnes dies Iared nongenti sexaginta duo anni et mortuus est
GEN|5|21|porro Enoch vixit sexaginta quinque annis et genuit Mathusalam
GEN|5|22|et ambulavit Enoch cum Deo postquam genuit Mathusalam trecentis annis et genuit filios et filias
GEN|5|23|et facti sunt omnes dies Enoch trecenti sexaginta quinque anni
GEN|5|24|ambulavitque cum Deo et non apparuit quia tulit eum Deus
GEN|5|25|vixit quoque Mathusalam centum octoginta septem annos et genuit Lamech
GEN|5|26|et vixit Mathusalam postquam genuit Lamech septingentos octoginta duos annos et genuit filios et filias
GEN|5|27|et facti sunt omnes dies Mathusalae nongenti sexaginta novem anni et mortuus est
GEN|5|28|vixit autem Lamech centum octoginta duobus annis et genuit filium
GEN|5|29|vocavitque nomen eius Noe dicens iste consolabitur nos ab operibus et laboribus manuum nostrarum in terra cui maledixit Dominus
GEN|5|30|vixitque Lamech postquam genuit Noe quingentos nonaginta quinque annos et genuit filios et filias
GEN|5|31|et facti sunt omnes dies Lamech septingenti septuaginta septem anni et mortuus est
GEN|5|32|Noe vero cum quingentorum esset annorum genuit Sem et Ham et Iafeth
GEN|6|1|cumque coepissent homines multiplicari super terram et filias procreassent
GEN|6|2|videntes filii Dei filias eorum quod essent pulchrae acceperunt uxores sibi ex omnibus quas elegerant
GEN|6|3|dixitque Deus non permanebit spiritus meus in homine in aeternum quia caro est eruntque dies illius centum viginti annorum
GEN|6|4|gigantes autem erant super terram in diebus illis postquam enim ingressi sunt filii Dei ad filias hominum illaeque genuerunt isti sunt potentes a saeculo viri famosi
GEN|6|5|videns autem Deus quod multa malitia hominum esset in terra et cuncta cogitatio cordis intenta esset ad malum omni tempore
GEN|6|6|paenituit eum quod hominem fecisset in terra et tactus dolore cordis intrinsecus
GEN|6|7|delebo inquit hominem quem creavi a facie terrae ab homine usque ad animantia a reptili usque ad volucres caeli paenitet enim me fecisse eos
GEN|6|8|Noe vero invenit gratiam coram Domino
GEN|6|9|hae generationes Noe Noe vir iustus atque perfectus fuit in generationibus suis cum Deo ambulavit
GEN|6|10|et genuit tres filios Sem Ham et Iafeth
GEN|6|11|corrupta est autem terra coram Deo et repleta est iniquitate
GEN|6|12|cumque vidisset Deus terram esse corruptam omnis quippe caro corruperat viam suam super terram
GEN|6|13|dixit ad Noe finis universae carnis venit coram me repleta est terra iniquitate a facie eorum et ego disperdam eos cum terra
GEN|6|14|fac tibi arcam de lignis levigatis mansiunculas in arca facies et bitumine linies intrinsecus et extrinsecus
GEN|6|15|et sic facies eam trecentorum cubitorum erit longitudo arcae quinquaginta cubitorum latitudo et triginta cubitorum altitudo illius
GEN|6|16|fenestram in arca facies et in cubito consummabis summitatem ostium autem arcae pones ex latere deorsum cenacula et tristega facies in ea
GEN|6|17|ecce ego adducam diluvii aquas super terram ut interficiam omnem carnem in qua spiritus vitae est subter caelum universa quae in terra sunt consumentur
GEN|6|18|ponamque foedus meum tecum et ingredieris arcam tu et filii tui uxor tua et uxores filiorum tuorum tecum
GEN|6|19|et ex cunctis animantibus universae carnis bina induces in arcam ut vivant tecum masculini sexus et feminini
GEN|6|20|de volucribus iuxta genus suum et de iumentis in genere suo et ex omni reptili terrae secundum genus suum bina de omnibus ingredientur tecum ut possint vivere
GEN|6|21|tolles igitur tecum ex omnibus escis quae mandi possunt et conportabis apud te et erunt tam tibi quam illis in cibum
GEN|6|22|fecit ergo Noe omnia quae praeceperat illi Deus
GEN|7|1|dixitque Dominus ad eum ingredere tu et omnis domus tua arcam te enim vidi iustum coram me in generatione hac
GEN|7|2|ex omnibus animantibus mundis tolle septena septena masculum et feminam de animantibus vero non mundis duo duo masculum et feminam
GEN|7|3|sed et de volatilibus caeli septena septena masculum et feminam ut salvetur semen super faciem universae terrae
GEN|7|4|adhuc enim et post dies septem ego pluam super terram quadraginta diebus et quadraginta noctibus et delebo omnem substantiam quam feci de superficie terrae
GEN|7|5|fecit ergo Noe omnia quae mandaverat ei Dominus
GEN|7|6|eratque sescentorum annorum quando diluvii aquae inundaverunt super terram
GEN|7|7|et ingressus est Noe et filii eius uxor eius et uxores filiorum eius cum eo in arcam propter aquas diluvii
GEN|7|8|de animantibus quoque mundis et inmundis et de volucribus et ex omni quod movetur super terram
GEN|7|9|duo et duo ingressa sunt ad Noe in arcam masculus et femina sicut praeceperat Deus Noe
GEN|7|10|cumque transissent septem dies aquae diluvii inundaverunt super terram
GEN|7|11|anno sescentesimo vitae Noe mense secundo septimodecimo die mensis rupti sunt omnes fontes abyssi magnae et cataractae caeli apertae sunt
GEN|7|12|et facta est pluvia super terram quadraginta diebus et quadraginta noctibus
GEN|7|13|in articulo diei illius ingressus est Noe et Sem et Ham et Iafeth filii eius uxor illius et tres uxores filiorum eius cum eis in arcam
GEN|7|14|ipsi et omne animal secundum genus suum universaque iumenta in genus suum et omne quod movetur super terram in genere suo cunctumque volatile secundum genus suum universae aves omnesque volucres
GEN|7|15|ingressae sunt ad Noe in arcam bina et bina ex omni carne in qua erat spiritus vitae
GEN|7|16|et quae ingressa sunt masculus et femina ex omni carne introierunt sicut praeceperat ei Deus et inclusit eum Dominus de foris
GEN|7|17|factumque est diluvium quadraginta diebus super terram et multiplicatae sunt aquae et elevaverunt arcam in sublime a terra
GEN|7|18|vehementer inundaverunt et omnia repleverunt in superficie terrae porro arca ferebatur super aquas
GEN|7|19|et aquae praevaluerunt nimis super terram opertique sunt omnes montes excelsi sub universo caelo
GEN|7|20|quindecim cubitis altior fuit aqua super montes quos operuerat
GEN|7|21|consumptaque est omnis caro quae movebatur super terram volucrum animantium bestiarum omniumque reptilium quae reptant super terram universi homines
GEN|7|22|et cuncta in quibus spiraculum vitae est in terra mortua sunt
GEN|7|23|et delevit omnem substantiam quae erat super terram ab homine usque ad pecus tam reptile quam volucres caeli et deleta sunt de terra remansit autem solus Noe et qui cum eo erant in arca
GEN|7|24|obtinueruntque aquae terras centum quinquaginta diebus
GEN|8|1|recordatus autem Deus Noe cunctarumque animantium et omnium iumentorum quae erant cum eo in arca adduxit spiritum super terram et inminutae sunt aquae
GEN|8|2|et clausi sunt fontes abyssi et cataractae caeli et prohibitae sunt pluviae de caelo
GEN|8|3|reversaeque aquae de terra euntes et redeuntes et coeperunt minui post centum quinquaginta dies
GEN|8|4|requievitque arca mense septimo vicesima septima die mensis super montes Armeniae
GEN|8|5|at vero aquae ibant et decrescebant usque ad decimum mensem decimo enim mense prima die mensis apparuerunt cacumina montium
GEN|8|6|cumque transissent quadraginta dies aperiens Noe fenestram arcae quam fecerat dimisit corvum
GEN|8|7|qui egrediebatur et revertebatur donec siccarentur aquae super terram
GEN|8|8|emisit quoque columbam post eum ut videret si iam cessassent aquae super faciem terrae
GEN|8|9|quae cum non invenisset ubi requiesceret pes eius reversa est ad eum in arcam aquae enim erant super universam terram extenditque manum et adprehensam intulit in arcam
GEN|8|10|expectatis autem ultra septem diebus aliis rursum dimisit columbam ex arca
GEN|8|11|at illa venit ad eum ad vesperam portans ramum olivae virentibus foliis in ore suo intellexit ergo Noe quod cessassent aquae super terram
GEN|8|12|expectavitque nihilominus septem alios dies et emisit columbam quae non est reversa ultra ad eum
GEN|8|13|igitur sescentesimo primo anno primo mense prima die mensis inminutae sunt aquae super terram et aperiens Noe tectum arcae aspexit viditque quod exsiccata esset superficies terrae
GEN|8|14|mense secundo septima et vicesima die mensis arefacta est terra
GEN|8|15|locutus est autem Deus ad Noe dicens
GEN|8|16|egredere de arca tu et uxor tua filii tui et uxores filiorum tuorum tecum
GEN|8|17|cuncta animantia quae sunt apud te ex omni carne tam in volatilibus quam in bestiis et in universis reptilibus quae reptant super terram educ tecum et ingredimini super terram crescite et multiplicamini super eam
GEN|8|18|egressus est ergo Noe et filii eius uxor illius et uxores filiorum eius cum eo
GEN|8|19|sed et omnia animantia iumenta et reptilia quae repunt super terram secundum genus suum arcam egressa sunt
GEN|8|20|aedificavit autem Noe altare Domino et tollens de cunctis pecoribus et volucribus mundis obtulit holocausta super altare
GEN|8|21|odoratusque est Dominus odorem suavitatis et ait ad eum nequaquam ultra maledicam terrae propter homines sensus enim et cogitatio humani cordis in malum prona sunt ab adulescentia sua non igitur ultra percutiam omnem animantem sicut feci
GEN|8|22|cunctis diebus terrae sementis et messis frigus et aestus aestas et hiemps nox et dies non requiescent
GEN|9|1|benedixitque Deus Noe et filiis eius et dixit ad eos crescite et multiplicamini et implete terram
GEN|9|2|et terror vester ac tremor sit super cuncta animalia terrae et super omnes volucres caeli cum universis quae moventur in terra omnes pisces maris manui vestrae traditi sunt
GEN|9|3|et omne quod movetur et vivit erit vobis in cibum quasi holera virentia tradidi vobis omnia
GEN|9|4|excepto quod carnem cum sanguine non comedetis
GEN|9|5|sanguinem enim animarum vestrarum requiram de manu cunctarum bestiarum et de manu hominis de manu viri et fratris eius requiram animam hominis
GEN|9|6|quicumque effuderit humanum sanguinem fundetur sanguis illius ad imaginem quippe Dei factus est homo
GEN|9|7|vos autem crescite et multiplicamini et ingredimini super terram et implete eam
GEN|9|8|haec quoque dixit Deus ad Noe et ad filios eius cum eo
GEN|9|9|ecce ego statuam pactum meum vobiscum et cum semine vestro post vos
GEN|9|10|et ad omnem animam viventem quae est vobiscum tam in volucribus quam in iumentis et pecudibus terrae cunctis quae egressa sunt de arca et universis bestiis terrae
GEN|9|11|statuam pactum meum vobiscum et nequaquam ultra interficietur omnis caro aquis diluvii neque erit deinceps diluvium dissipans terram
GEN|9|12|dixitque Deus hoc signum foederis quod do inter me et vos et ad omnem animam viventem quae est vobiscum in generationes sempiternas
GEN|9|13|arcum meum ponam in nubibus et erit signum foederis inter me et inter terram
GEN|9|14|cumque obduxero nubibus caelum apparebit arcus meus in nubibus
GEN|9|15|et recordabor foederis mei vobiscum et cum omni anima vivente quae carnem vegetat et non erunt ultra aquae diluvii ad delendam universam carnem
GEN|9|16|eritque arcus in nubibus et videbo illum et recordabor foederis sempiterni quod pactum est inter Deum et inter omnem animam viventem universae carnis quae est super terram
GEN|9|17|dixitque Deus Noe hoc erit signum foederis quod constitui inter me et inter omnem carnem super terram
GEN|9|18|erant igitur filii Noe qui egressi sunt de arca Sem Ham et Iafeth porro Ham ipse est pater Chanaan
GEN|9|19|tres isti sunt filii Noe et ab his disseminatum est omne hominum genus super universam terram
GEN|9|20|coepitque Noe vir agricola exercere terram et plantavit vineam
GEN|9|21|bibensque vinum inebriatus est et nudatus in tabernaculo suo
GEN|9|22|quod cum vidisset Ham pater Chanaan verenda scilicet patris sui esse nuda nuntiavit duobus fratribus suis foras
GEN|9|23|at vero Sem et Iafeth pallium inposuerunt umeris suis et incedentes retrorsum operuerunt verecunda patris sui faciesque eorum aversae erant et patris virilia non viderunt
GEN|9|24|evigilans autem Noe ex vino cum didicisset quae fecerat ei filius suus minor
GEN|9|25|ait maledictus Chanaan servus servorum erit fratribus suis
GEN|9|26|dixitque benedictus Dominus Deus Sem sit Chanaan servus eius
GEN|9|27|dilatet Deus Iafeth et habitet in tabernaculis Sem sitque Chanaan servus eius
GEN|9|28|vixit autem Noe post diluvium trecentis quinquaginta annis
GEN|9|29|et impleti sunt omnes dies eius nongentorum quinquaginta annorum et mortuus est
GEN|10|1|hae generationes filiorum Noe Sem Ham Iafeth natique sunt eis filii post diluvium
GEN|10|2|filii Iafeth Gomer Magog et Madai Iavan et Thubal et Mosoch et Thiras
GEN|10|3|porro filii Gomer Aschenez et Rifath et Thogorma
GEN|10|4|filii autem Iavan Elisa et Tharsis Cetthim et Dodanim
GEN|10|5|ab his divisae sunt insulae gentium in regionibus suis unusquisque secundum linguam et familias in nationibus suis
GEN|10|6|filii autem Ham Chus et Mesraim et Fut et Chanaan
GEN|10|7|filii Chus Saba et Hevila et Sabatha et Regma et Sabathaca filii Regma Saba et Dadan
GEN|10|8|porro Chus genuit Nemrod ipse coepit esse potens in terra
GEN|10|9|et erat robustus venator coram Domino ab hoc exivit proverbium quasi Nemrod robustus venator coram Domino
GEN|10|10|fuit autem principium regni eius Babylon et Arach et Archad et Chalanne in terra Sennaar
GEN|10|11|de terra illa egressus est Assur et aedificavit Nineven et plateas civitatis et Chale
GEN|10|12|Resen quoque inter Nineven et Chale haec est civitas magna
GEN|10|13|at vero Mesraim genuit Ludim et Anamim et Laabim Nepthuim
GEN|10|14|et Phetrusim et Cesluim de quibus egressi sunt Philisthim et Capthurim
GEN|10|15|Chanaan autem genuit Sidonem primogenitum suum Ettheum
GEN|10|16|et Iebuseum et Amorreum Gergeseum
GEN|10|17|Eveum et Araceum Sineum
GEN|10|18|et Aradium Samariten et Amatheum et post haec disseminati sunt populi Chananeorum
GEN|10|19|factique sunt termini Chanaan venientibus a Sidone Geraram usque Gazam donec ingrediaris Sodomam et Gomorram et Adama et Seboim usque Lesa
GEN|10|20|hii filii Ham in cognationibus et linguis et generationibus terrisque et gentibus suis
GEN|10|21|de Sem quoque nati sunt patre omnium filiorum Eber fratre Iafeth maiore
GEN|10|22|filii Sem Aelam et Assur et Arfaxad et Lud et Aram
GEN|10|23|filii Aram Us et Hul et Gether et Mes
GEN|10|24|at vero Arfaxad genuit Sala de quo ortus est Eber
GEN|10|25|natique sunt Eber filii duo nomen uni Faleg eo quod in diebus eius divisa sit terra et nomen fratris eius Iectan
GEN|10|26|qui Iectan genuit Helmodad et Saleph et Asarmoth Iare
GEN|10|27|et Aduram et Uzal Decla
GEN|10|28|et Ebal et Abimahel Saba
GEN|10|29|et Ophir et Evila et Iobab omnes isti filii Iectan
GEN|10|30|et facta est habitatio eorum de Messa pergentibus usque Sephar montem orientalem
GEN|10|31|isti filii Sem secundum cognationes et linguas et regiones in gentibus suis
GEN|10|32|hae familiae Noe iuxta populos et nationes suas ab his divisae sunt gentes in terra post diluvium
GEN|11|1|erat autem terra labii unius et sermonum eorundem
GEN|11|2|cumque proficiscerentur de oriente invenerunt campum in terra Sennaar et habitaverunt in eo
GEN|11|3|dixitque alter ad proximum suum venite faciamus lateres et coquamus eos igni habueruntque lateres pro saxis et bitumen pro cemento
GEN|11|4|et dixerunt venite faciamus nobis civitatem et turrem cuius culmen pertingat ad caelum et celebremus nomen nostrum antequam dividamur in universas terras
GEN|11|5|descendit autem Dominus ut videret civitatem et turrem quam aedificabant filii Adam
GEN|11|6|et dixit ecce unus est populus et unum labium omnibus coeperuntque hoc facere nec desistent a cogitationibus suis donec eas opere conpleant
GEN|11|7|venite igitur descendamus et confundamus ibi linguam eorum ut non audiat unusquisque vocem proximi sui
GEN|11|8|atque ita divisit eos Dominus ex illo loco in universas terras et cessaverunt aedificare civitatem
GEN|11|9|et idcirco vocatum est nomen eius Babel quia ibi confusum est labium universae terrae et inde dispersit eos Dominus super faciem cunctarum regionum
GEN|11|10|hae generationes Sem Sem centum erat annorum quando genuit Arfaxad biennio post diluvium
GEN|11|11|vixitque Sem postquam genuit Arfaxad quingentos annos et genuit filios et filias
GEN|11|12|porro Arfaxad vixit triginta quinque annos et genuit Sale
GEN|11|13|vixitque Arfaxad postquam genuit Sale trecentis tribus annis et genuit filios et filias
GEN|11|14|Sale quoque vixit triginta annis et genuit Eber
GEN|11|15|vixitque Sale postquam genuit Eber quadringentis tribus annis et genuit filios et filias
GEN|11|16|vixit autem Eber triginta quattuor annis et genuit Faleg
GEN|11|17|et vixit Eber postquam genuit Faleg quadringentis triginta annis et genuit filios et filias
GEN|11|18|vixit quoque Faleg triginta annis et genuit Reu
GEN|11|19|vixitque Faleg postquam genuit Reu ducentis novem annis et genuit filios et filias
GEN|11|20|vixit autem Reu triginta duobus annis et genuit Sarug
GEN|11|21|vixitque Reu postquam genuit Sarug ducentis septem annis et genuit filios et filias
GEN|11|22|vixit vero Sarug triginta annis et genuit Nahor
GEN|11|23|vixitque Sarug postquam genuit Nahor ducentos annos et genuit filios et filias
GEN|11|24|vixit autem Nahor viginti novem annis et genuit Thare
GEN|11|25|vixitque Nahor postquam genuit Thare centum decem et novem annos et genuit filios et filias
GEN|11|26|vixitque Thare septuaginta annis et genuit Abram et Nahor et Aran
GEN|11|27|hae sunt autem generationes Thare Thare genuit Abram et Nahor et Aran porro Aran genuit Loth
GEN|11|28|mortuusque est Aran ante Thare patrem suum in terra nativitatis suae in Ur Chaldeorum
GEN|11|29|duxerunt autem Abram et Nahor uxores nomen autem uxoris Abram Sarai et nomen uxoris Nahor Melcha filia Aran patris Melchae et patris Ieschae
GEN|11|30|erat autem Sarai sterilis nec habebat liberos
GEN|11|31|tulit itaque Thare Abram filium suum et Loth filium Aran filium filii sui et Sarai nurum suam uxorem Abram filii sui et eduxit eos de Ur Chaldeorum ut irent in terram Chanaan veneruntque usque Haran et habitaverunt ibi
GEN|11|32|et facti sunt dies Thare ducentorum quinque annorum et mortuus est in Haran
GEN|12|1|dixit autem Dominus ad Abram egredere de terra tua et de cognatione tua et de domo patris tui in terram quam monstrabo tibi
GEN|12|2|faciamque te in gentem magnam et benedicam tibi et magnificabo nomen tuum erisque benedictus
GEN|12|3|benedicam benedicentibus tibi et maledicam maledicentibus tibi atque in te benedicentur universae cognationes terrae
GEN|12|4|egressus est itaque Abram sicut praeceperat ei Dominus et ivit cum eo Loth septuaginta quinque annorum erat Abram cum egrederetur de Haran
GEN|12|5|tulitque Sarai uxorem suam et Loth filium fratris sui universamque substantiam quam possederant et animas quas fecerant in Haran et egressi sunt ut irent in terram Chanaan cumque venissent in eam
GEN|12|6|pertransivit Abram terram usque ad locum Sychem usque ad convallem Inlustrem Chananeus autem tunc erat in terra
GEN|12|7|apparuitque Dominus Abram et dixit ei semini tuo dabo terram hanc qui aedificavit ibi altare Domino qui apparuerat ei
GEN|12|8|et inde transgrediens ad montem qui erat contra orientem Bethel tetendit ibi tabernaculum suum ab occidente habens Bethel et ab oriente Ai aedificavit quoque ibi altare Domino et invocavit nomen eius
GEN|12|9|perrexitque Abram vadens et ultra progrediens ad meridiem
GEN|12|10|facta est autem fames in terra descenditque Abram in Aegyptum ut peregrinaretur ibi praevaluerat enim fames in terra
GEN|12|11|cumque prope esset ut ingrederetur Aegyptum dixit Sarai uxori suae novi quod pulchra sis mulier
GEN|12|12|et quod cum viderint te Aegyptii dicturi sunt uxor ipsius est et interficient me et te reservabunt
GEN|12|13|dic ergo obsecro te quod soror mea sis ut bene sit mihi propter te et vivat anima mea ob gratiam tui
GEN|12|14|cum itaque ingressus esset Abram Aegyptum viderunt Aegyptii mulierem quod esset pulchra nimis
GEN|12|15|et nuntiaverunt principes Pharaoni et laudaverunt eam apud illum et sublata est mulier in domum Pharaonis
GEN|12|16|Abram vero bene usi sunt propter illam fueruntque ei oves et boves et asini et servi et famulae et asinae et cameli
GEN|12|17|flagellavit autem Dominus Pharaonem plagis maximis et domum eius propter Sarai uxorem Abram
GEN|12|18|vocavitque Pharao Abram et dixit ei quidnam est quod fecisti mihi quare non indicasti quod uxor tua esset
GEN|12|19|quam ob causam dixisti esse sororem tuam ut tollerem eam mihi in uxorem nunc igitur ecce coniux tua accipe eam et vade
GEN|12|20|praecepitque Pharao super Abram viris et deduxerunt eum et uxorem illius et omnia quae habebat
GEN|13|1|ascendit ergo Abram de Aegypto ipse et uxor eius et omnia quae habebat et Loth cum eo ad australem plagam
GEN|13|2|erat autem dives valde in possessione argenti et auri
GEN|13|3|reversusque est per iter quo venerat a meridie in Bethel usque ad locum ubi prius fixerat tabernaculum inter Bethel et Ai
GEN|13|4|in loco altaris quod fecerat prius et invocavit ibi nomen Domini
GEN|13|5|sed et Loth qui erat cum Abram fuerunt greges ovium et armenta et tabernacula
GEN|13|6|nec poterat eos capere terra ut habitarent simul erat quippe substantia eorum multa et non quibant habitare communiter
GEN|13|7|unde et facta est rixa inter pastores gregum Abram et Loth eo autem tempore Chananeus et Ferezeus habitabant in illa terra
GEN|13|8|dixit ergo Abram ad Loth ne quaeso sit iurgium inter me et te et inter pastores meos et pastores tuos fratres enim sumus
GEN|13|9|ecce universa terra coram te est recede a me obsecro si ad sinistram ieris ego ad dexteram tenebo si tu dexteram elegeris ego ad sinistram pergam
GEN|13|10|elevatis itaque Loth oculis vidit omnem circa regionem Iordanis quae universa inrigabatur antequam subverteret Dominus Sodomam et Gomorram sicut paradisus Domini et sicut Aegyptus venientibus in Segor
GEN|13|11|elegitque sibi Loth regionem circa Iordanem et recessit ab oriente divisique sunt alterutrum a fratre suo
GEN|13|12|Abram habitavit in terra Chanaan Loth moratus est in oppidis quae erant circa Iordanem et habitavit in Sodomis
GEN|13|13|homines autem Sodomitae pessimi erant et peccatores coram Domino nimis
GEN|13|14|dixitque Dominus ad Abram postquam divisus est Loth ab eo leva oculos tuos et vide a loco in quo nunc es ad aquilonem et ad meridiem ad orientem et ad occidentem
GEN|13|15|omnem terram quam conspicis tibi dabo et semini tuo usque in sempiternum
GEN|13|16|faciamque semen tuum sicut pulverem terrae si quis potest hominum numerare pulverem semen quoque tuum numerare poterit
GEN|13|17|surge et perambula terram in longitudine et in latitudine sua quia tibi daturus sum eam
GEN|13|18|movens igitur Abram tabernaculum suum venit et habitavit iuxta convallem Mambre quod est in Hebron aedificavitque ibi altare Domino
GEN|14|1|factum est autem in illo tempore ut Amrafel rex Sennaar et Arioch rex Ponti et Chodorlahomor rex Aelamitarum et Thadal rex Gentium
GEN|14|2|inirent bellum contra Bara regem Sodomorum et contra Bersa regem Gomorrae et contra Sennaab regem Adamae et contra Semeber regem Seboim contraque regem Balae ipsa est Segor
GEN|14|3|omnes hii convenerunt in vallem Silvestrem quae nunc est mare Salis
GEN|14|4|duodecim enim annis servierant Chodorlahomor et tertiodecimo anno recesserunt ab eo
GEN|14|5|igitur anno quartodecimo venit Chodorlahomor et reges qui erant cum eo percusseruntque Rafaim in Astharothcarnaim et Zuzim cum eis et Emim in Savecariathaim
GEN|14|6|et Chorreos in montibus Seir usque ad campestria Pharan quae est in solitudine
GEN|14|7|reversique sunt et venerunt ad fontem Mesfat ipsa est Cades et percusserunt omnem regionem Amalechitarum et Amorreum qui habitabat in Asasonthamar
GEN|14|8|et egressi sunt rex Sodomorum et rex Gomorrae rexque Adamae et rex Seboim necnon et rex Balae quae est Segor et direxerunt contra eos aciem in valle Silvestri
GEN|14|9|scilicet adversum Chodorlahomor regem Aelamitarum et Thadal regem Gentium et Amrafel regem Sennaar et Arioch regem Ponti quattuor reges adversus quinque
GEN|14|10|vallis autem Silvestris habebat puteos multos bituminis itaque rex Sodomorum et Gomorrae terga verterunt cecideruntque ibi et qui remanserant fugerunt ad montem
GEN|14|11|tulerunt autem omnem substantiam Sodomorum et Gomorrae et universa quae ad cibum pertinent et abierunt
GEN|14|12|necnon et Loth et substantiam eius filium fratris Abram qui habitabat in Sodomis
GEN|14|13|et ecce unus qui evaserat nuntiavit Abram Hebraeo qui habitabat in convalle Mambre Amorrei fratris Eschol et fratris Aner hii enim pepigerant foedus cum Abram
GEN|14|14|quod cum audisset Abram captum videlicet Loth fratrem suum numeravit expeditos vernaculos suos trecentos decem et octo et persecutus est eos usque Dan
GEN|14|15|et divisis sociis inruit super eos nocte percussitque eos et persecutus est usque Hoba quae est ad levam Damasci
GEN|14|16|reduxitque omnem substantiam et Loth fratrem suum cum substantia illius mulieres quoque et populum
GEN|14|17|egressus est autem rex Sodomorum in occursum eius postquam reversus est a caede Chodorlahomor et regum qui cum eo erant in valle Save quae est vallis Regis
GEN|14|18|at vero Melchisedech rex Salem proferens panem et vinum erat enim sacerdos Dei altissimi
GEN|14|19|benedixit ei et ait benedictus Abram Deo excelso qui creavit caelum et terram
GEN|14|20|et benedictus Deus excelsus quo protegente hostes in manibus tuis sunt et dedit ei decimas ex omnibus
GEN|14|21|dixit autem rex Sodomorum ad Abram da mihi animas cetera tolle tibi
GEN|14|22|qui respondit ei levo manum meam ad Dominum Deum excelsum possessorem caeli et terrae
GEN|14|23|quod a filo subteminis usque ad corrigiam caligae non accipiam ex omnibus quae tua sunt ne dicas ego ditavi Abram
GEN|14|24|exceptis his quae comederunt iuvenes et partibus virorum qui venerunt mecum Aner Eschol et Mambre isti accipient partes suas
GEN|15|1|his itaque transactis factus est sermo Domini ad Abram per visionem dicens noli timere Abram ego protector tuus sum et merces tua magna nimis
GEN|15|2|dixitque Abram Domine Deus quid dabis mihi ego vadam absque liberis et filius procuratoris domus meae iste Damascus Eliezer
GEN|15|3|addiditque Abram mihi autem non dedisti semen et ecce vernaculus meus heres meus erit
GEN|15|4|statimque sermo Domini factus est ad eum dicens non erit hic heres tuus sed qui egredietur de utero tuo ipsum habebis heredem
GEN|15|5|eduxitque eum foras et ait illi suspice caelum et numera stellas si potes et dixit ei sic erit semen tuum
GEN|15|6|credidit Domino et reputatum est ei ad iustitiam
GEN|15|7|dixitque ad eum ego Dominus qui eduxi te de Ur Chaldeorum ut darem tibi terram istam et possideres eam
GEN|15|8|at ille ait Domine Deus unde scire possum quod possessurus sim eam
GEN|15|9|respondens Dominus sume inquit mihi vaccam triennem et capram trimam et arietem annorum trium turturem quoque et columbam
GEN|15|10|qui tollens universa haec divisit per medium et utrasque partes contra se altrinsecus posuit aves autem non divisit
GEN|15|11|descenderuntque volucres super cadavera et abigebat eas Abram
GEN|15|12|cumque sol occumberet sopor inruit super Abram et horror magnus et tenebrosus invasit eum
GEN|15|13|dictumque est ad eum scito praenoscens quod peregrinum futurum sit semen tuum in terra non sua et subicient eos servituti et adfligent quadringentis annis
GEN|15|14|verumtamen gentem cui servituri sunt ego iudicabo et post haec egredientur cum magna substantia
GEN|15|15|tu autem ibis ad patres tuos in pace sepultus in senectute bona
GEN|15|16|generatione autem quarta revertentur huc necdum enim conpletae sunt iniquitates Amorreorum usque ad praesens tempus
GEN|15|17|cum ergo occubuisset sol facta est caligo tenebrosa et apparuit clibanus fumans et lampas ignis transiens inter divisiones illas
GEN|15|18|in die illo pepigit Dominus cum Abram foedus dicens semini tuo dabo terram hanc a fluvio Aegypti usque ad fluvium magnum flumen Eufraten
GEN|15|19|Cineos et Cenezeos et Cedmoneos
GEN|15|20|et Hettheos et Ferezeos Rafaim quoque
GEN|15|21|et Amorreos et Chananeos et Gergeseos et Iebuseos
GEN|16|1|igitur Sarai uxor Abram non genuerat liberos sed habens ancillam aegyptiam nomine Agar
GEN|16|2|dixit marito suo ecce conclusit me Dominus ne parerem ingredere ad ancillam meam si forte saltem ex illa suscipiam filios cumque ille adquiesceret deprecanti
GEN|16|3|tulit Agar Aegyptiam ancillam suam post annos decem quam habitare coeperant in terra Chanaan et dedit eam viro suo uxorem
GEN|16|4|qui ingressus est ad eam at illa concepisse se videns despexit dominam suam
GEN|16|5|dixitque Sarai ad Abram inique agis contra me ego dedi ancillam meam in sinum tuum quae videns quod conceperit despectui me habet iudicet Dominus inter me et te
GEN|16|6|cui respondens Abram ecce ait ancilla tua in manu tua est utere ea ut libet adfligente igitur eam Sarai fugam iniit
GEN|16|7|cumque invenisset illam angelus Domini iuxta fontem aquae in solitudine qui est in via Sur
GEN|16|8|dixit ad eam Agar ancilla Sarai unde venis et quo vadis quae respondit a facie Sarai dominae meae ego fugio
GEN|16|9|dixitque ei angelus Domini revertere ad dominam tuam et humiliare sub manibus ipsius
GEN|16|10|et rursum multiplicans inquit multiplicabo semen tuum et non numerabitur prae multitudine
GEN|16|11|ac deinceps ecce ait concepisti et paries filium vocabisque nomen eius Ismahel eo quod audierit Dominus adflictionem tuam
GEN|16|12|hic erit ferus homo manus eius contra omnes et manus omnium contra eum et e regione universorum fratrum suorum figet tabernacula
GEN|16|13|vocavit autem nomen Domini qui loquebatur ad eam Tu Deus qui vidisti me dixit enim profecto hic vidi posteriora videntis me
GEN|16|14|propterea appellavit puteum illum puteum Viventis et videntis me ipse est inter Cades et Barad
GEN|16|15|peperitque Abrae filium qui vocavit nomen eius Ismahel
GEN|16|16|octoginta et sex annorum erat quando peperit ei Agar Ismahelem
GEN|17|1|postquam vero nonaginta et novem annorum esse coeperat apparuit ei Dominus dixitque ad eum ego Deus omnipotens ambula coram me et esto perfectus
GEN|17|2|ponamque foedus meum inter me et te et multiplicabo te vehementer nimis
GEN|17|3|cecidit Abram pronus in faciem
GEN|17|4|dixitque ei Deus ego sum et pactum meum tecum erisque pater multarum gentium
GEN|17|5|nec ultra vocabitur nomen tuum Abram sed appellaberis Abraham quia patrem multarum gentium constitui te
GEN|17|6|faciamque te crescere vehementissime et ponam in gentibus regesque ex te egredientur
GEN|17|7|et statuam pactum meum inter me et te et inter semen tuum post te in generationibus suis foedere sempiterno ut sim Deus tuus et seminis tui post te
GEN|17|8|daboque tibi et semini tuo terram peregrinationis tuae omnem terram Chanaan in possessionem aeternam eroque Deus eorum
GEN|17|9|dixit iterum Deus ad Abraham et tu ergo custodies pactum meum et semen tuum post te in generationibus suis
GEN|17|10|hoc est pactum quod observabitis inter me et vos et semen tuum post te circumcidetur ex vobis omne masculinum
GEN|17|11|et circumcidetis carnem praeputii vestri ut sit in signum foederis inter me et vos
GEN|17|12|infans octo dierum circumcidetur in vobis omne masculinum in generationibus vestris tam vernaculus quam empticius circumcidetur et quicumque non fuerit de stirpe vestra
GEN|17|13|eritque pactum meum in carne vestra in foedus aeternum
GEN|17|14|masculus cuius praeputii caro circumcisa non fuerit delebitur anima illa de populo suo quia pactum meum irritum fecit
GEN|17|15|dixit quoque Deus ad Abraham Sarai uxorem tuam non vocabis Sarai sed Sarram
GEN|17|16|et benedicam ei et ex illa dabo tibi filium cui benedicturus sum eritque in nationes et reges populorum orientur ex eo
GEN|17|17|cecidit Abraham in faciem et risit dicens in corde suo putasne centenario nascetur filius et Sarra nonagenaria pariet
GEN|17|18|dixitque ad Deum utinam Ismahel vivat coram te
GEN|17|19|et ait Deus ad Abraham Sarra uxor tua pariet tibi filium vocabisque nomen eius Isaac et constituam pactum meum illi in foedus sempiternum et semini eius post eum
GEN|17|20|super Ismahel quoque exaudivi te ecce benedicam ei et augebo et multiplicabo eum valde duodecim duces generabit et faciam illum in gentem magnam
GEN|17|21|pactum vero meum statuam ad Isaac quem pariet tibi Sarra tempore isto in anno altero
GEN|17|22|cumque finitus esset sermo loquentis cum eo ascendit Deus ab Abraham
GEN|17|23|tulit autem Abraham Ismahelem filium suum et omnes vernaculos domus suae universosque quos emerat cunctos mares ex omnibus viris domus suae et circumcidit carnem praeputii eorum statim in ipsa die sicut praeceperat ei Deus
GEN|17|24|nonaginta novem erat annorum quando circumcidit carnem praeputii sui
GEN|17|25|et Ismahel filius eius tredecim annos impleverat tempore circumcisionis suae
GEN|17|26|eadem die circumcisus est Abraham et Ismahel filius eius
GEN|17|27|et omnes viri domus illius tam vernaculi quam empticii et alienigenae pariter circumcisi sunt
GEN|18|1|apparuit autem ei Dominus in convalle Mambre sedenti in ostio tabernaculi sui in ipso fervore diei
GEN|18|2|cumque elevasset oculos apparuerunt ei tres viri stantes propter eum quos cum vidisset cucurrit in occursum eorum de ostio tabernaculi et adoravit in terra
GEN|18|3|et dixit Domine si inveni gratiam in oculis tuis ne transeas servum tuum
GEN|18|4|sed adferam pauxillum aquae et lavate pedes vestros et requiescite sub arbore
GEN|18|5|ponam buccellam panis et confortate cor vestrum postea transibitis idcirco enim declinastis ad servum vestrum qui dixerunt fac ut locutus es
GEN|18|6|festinavit Abraham in tabernaculum ad Sarram dixitque ei adcelera tria sata similae commisce et fac subcinericios panes
GEN|18|7|ipse vero ad armentum cucurrit et tulit inde vitulum tenerrimum et optimum deditque puero qui festinavit et coxit illum
GEN|18|8|tulit quoque butyrum et lac et vitulum quem coxerat et posuit coram eis ipse vero stabat iuxta eos sub arbore
GEN|18|9|cumque comedissent dixerunt ad eum ubi est Sarra uxor tua ille respondit ecce in tabernaculo est
GEN|18|10|cui dixit revertens veniam ad te tempore isto vita comite et habebit filium Sarra uxor tua quo audito Sarra risit post ostium tabernaculi
GEN|18|11|erant autem ambo senes provectaeque aetatis et desierant Sarrae fieri muliebria
GEN|18|12|quae risit occulte dicens postquam consenui et dominus meus vetulus est voluptati operam dabo
GEN|18|13|dixit autem Dominus ad Abraham quare risit Sarra dicens num vere paritura sum anus
GEN|18|14|numquid Deo est quicquam difficile iuxta condictum revertar ad te hoc eodem tempore vita comite et habebit Sarra filium
GEN|18|15|negavit Sarra dicens non risi timore perterrita Dominus autem non est inquit ita sed risisti
GEN|18|16|cum ergo surrexissent inde viri direxerunt oculos suos contra Sodomam et Abraham simul gradiebatur deducens eos
GEN|18|17|dixitque Dominus num celare potero Abraham quae gesturus sum
GEN|18|18|cum futurus sit in gentem magnam ac robustissimam et benedicendae sint in illo omnes nationes terrae
GEN|18|19|scio enim quod praecepturus sit filiis suis et domui suae post se ut custodiant viam Domini et faciant iustitiam et iudicium ut adducat Dominus propter Abraham omnia quae locutus est ad eum
GEN|18|20|dixit itaque Dominus clamor Sodomorum et Gomorrae multiplicatus est et peccatum earum adgravatum est nimis
GEN|18|21|descendam et videbo utrum clamorem qui venit ad me opere conpleverint an non est ita ut sciam
GEN|18|22|converteruntque se inde et abierunt Sodomam Abraham vero adhuc stabat coram Domino
GEN|18|23|et adpropinquans ait numquid perdes iustum cum impio
GEN|18|24|si fuerint quinquaginta iusti in civitate peribunt simul et non parces loco illi propter quinquaginta iustos si fuerint in eo
GEN|18|25|absit a te ut rem hanc facias et occidas iustum cum impio fiatque iustus sicut impius non est hoc tuum qui iudicas omnem terram nequaquam facies iudicium
GEN|18|26|dixitque Dominus ad eum si invenero Sodomis quinquaginta iustos in medio civitatis dimittam omni loco propter eos
GEN|18|27|respondens Abraham ait quia semel coepi loquar ad Dominum meum cum sim pulvis et cinis
GEN|18|28|quid si minus quinquaginta iustis quinque fuerint delebis propter quinque universam urbem et ait non delebo si invenero ibi quadraginta quinque
GEN|18|29|rursumque locutus est ad eum sin autem quadraginta inventi fuerint quid facies ait non percutiam propter quadraginta
GEN|18|30|ne quaeso inquit indigneris Domine si loquar quid si inventi fuerint ibi triginta respondit non faciam si invenero ibi triginta
GEN|18|31|quia semel ait coepi loquar ad Dominum meum quid si inventi fuerint ibi viginti dixit non interficiam propter viginti
GEN|18|32|obsecro inquit ne irascaris Domine si loquar adhuc semel quid si inventi fuerint ibi decem dixit non delebo propter decem
GEN|18|33|abiit Dominus postquam cessavit loqui ad Abraham et ille reversus est in locum suum
GEN|19|1|veneruntque duo angeli Sodomam vespere sedente Loth in foribus civitatis qui cum vidisset surrexit et ivit obviam eis adoravitque pronus in terra
GEN|19|2|et dixit obsecro domini declinate in domum pueri vestri et manete ibi lavate pedes vestros et mane proficiscimini in viam vestram qui dixerunt minime sed in platea manebimus
GEN|19|3|conpulit illos oppido ut deverterent ad eum ingressisque domum illius fecit convivium coxit azyma et comederunt
GEN|19|4|prius autem quam irent cubitum viri civitatis vallaverunt domum a puero usque ad senem omnis populus simul
GEN|19|5|vocaveruntque Loth et dixerunt ei ubi sunt viri qui introierunt ad te nocte educ illos huc ut cognoscamus eos
GEN|19|6|egressus ad eos Loth post tergum adcludens ostium ait
GEN|19|7|nolite quaeso fratres mei nolite malum hoc facere
GEN|19|8|habeo duas filias quae necdum cognoverunt virum educam eas ad vos et abutimini eis sicut placuerit vobis dummodo viris istis nihil faciatis mali quia ingressi sunt sub umbraculum tegminis mei
GEN|19|9|at illi dixerunt recede illuc et rursus ingressus es inquiunt ut advena numquid ut iudices te ergo ipsum magis quam hos adfligemus vimque faciebant Loth vehementissime iam prope erat ut refringerent fores
GEN|19|10|et ecce miserunt manum viri et introduxerunt ad se Loth cluseruntque ostium
GEN|19|11|et eos qui erant foris percusserunt caecitate a minimo usque ad maximum ita ut ostium invenire non possent
GEN|19|12|dixerunt autem ad Loth habes hic tuorum quempiam generum aut filios aut filias omnes qui tui sunt educ de urbe hac
GEN|19|13|delebimus enim locum istum eo quod increverit clamor eorum coram Domino qui misit nos ut perdamus illos
GEN|19|14|egressus itaque Loth locutus est ad generos suos qui accepturi erant filias eius et dixit surgite egredimini de loco isto quia delebit Dominus civitatem hanc et visus est eis quasi ludens loqui
GEN|19|15|cumque esset mane cogebant eum angeli dicentes surge et tolle uxorem tuam et duas filias quas habes ne et tu pariter pereas in scelere civitatis
GEN|19|16|dissimulante illo adprehenderunt manum eius et manum uxoris ac duarum filiarum eius eo quod parceret Dominus illi
GEN|19|17|et eduxerunt eum posueruntque extra civitatem ibi locutus est ad eum salva animam tuam noli respicere post tergum nec stes in omni circa regione sed in monte salvum te fac ne et tu simul pereas
GEN|19|18|dixitque Loth ad eos quaeso Domine mi
GEN|19|19|quia invenit servus tuus gratiam coram te et magnificasti misericordiam tuam quam fecisti mecum ut salvares animam meam nec possum in monte salvari ne forte adprehendat me malum et moriar
GEN|19|20|est civitas haec iuxta ad quam possum fugere parva et salvabor in ea numquid non modica est et vivet anima mea
GEN|19|21|dixitque ad eum ecce etiam in hoc suscepi preces tuas ut non subvertam urbem pro qua locutus es
GEN|19|22|festina et salvare ibi quia non potero facere quicquam donec ingrediaris illuc idcirco vocatum est nomen urbis illius Segor
GEN|19|23|sol egressus est super terram et Loth ingressus est in Segor
GEN|19|24|igitur Dominus pluit super Sodomam et Gomorram sulphur et ignem a Domino de caelo
GEN|19|25|et subvertit civitates has et omnem circa regionem universos habitatores urbium et cuncta terrae virentia
GEN|19|26|respiciensque uxor eius post se versa est in statuam salis
GEN|19|27|Abraham autem consurgens mane ubi steterat prius cum Domino
GEN|19|28|intuitus est Sodomam et Gomorram et universam terram regionis illius viditque ascendentem favillam de terra quasi fornacis fumum
GEN|19|29|cum enim subverteret Deus civitates regionis illius recordatus est Abrahae et liberavit Loth de subversione urbium in quibus habitaverat
GEN|19|30|ascenditque Loth de Segor et mansit in monte duae quoque filiae eius cum eo timuerat enim manere in Segor et mansit in spelunca ipse et duae filiae eius
GEN|19|31|dixitque maior ad minorem pater noster senex est et nullus virorum remansit in terra qui possit ingredi ad nos iuxta morem universae terrae
GEN|19|32|veni inebriemus eum vino dormiamusque cum eo ut servare possimus ex patre nostro semen
GEN|19|33|dederunt itaque patri suo bibere vinum nocte illa et ingressa est maior dormivitque cum patre at ille non sensit nec quando accubuit filia nec quando surrexit
GEN|19|34|altera quoque die dixit maior ad minorem ecce dormivi heri cum patre meo demus ei bibere vinum etiam hac nocte et dormies cum eo ut salvemus semen de patre nostro
GEN|19|35|dederunt et illa nocte patri vinum ingressaque minor filia dormivit cum eo et nec tunc quidem sensit quando concubuerit vel quando illa surrexerit
GEN|19|36|conceperunt ergo duae filiae Loth de patre suo
GEN|19|37|peperitque maior filium et vocavit nomen eius Moab ipse est pater Moabitarum usque in praesentem diem
GEN|19|38|minor quoque peperit filium et vocavit nomen eius Ammon id est filius populi mei ipse est pater Ammanitarum usque hodie
GEN|20|1|profectus inde Abraham in terram australem habitavit inter Cades et Sur et peregrinatus est in Geraris
GEN|20|2|dixitque de Sarra uxore sua soror mea est misit ergo Abimelech rex Gerarae et tulit eam
GEN|20|3|venit autem Deus ad Abimelech per somnium noctis et ait ei en morieris propter mulierem quam tulisti habet enim virum
GEN|20|4|Abimelech vero non tetigerat eam et ait Domine num gentem ignorantem et iustam interficies
GEN|20|5|nonne ipse dixit mihi soror mea est et ipsa ait frater meus est in simplicitate cordis mei et munditia manuum mearum feci hoc
GEN|20|6|dixitque ad eum Deus et ego scio quod simplici corde feceris et ideo custodivi te ne peccares in me et non dimisi ut tangeres eam
GEN|20|7|nunc igitur redde uxorem viro suo quia propheta est et orabit pro te et vives si autem nolueris reddere scito quod morte morieris tu et omnia quae tua sunt
GEN|20|8|statimque de nocte consurgens Abimelech vocavit omnes servos suos et locutus est universa verba haec in auribus eorum timueruntque omnes viri valde
GEN|20|9|vocavit autem Abimelech etiam Abraham et dixit ei quid fecisti nobis quid peccavimus in te quia induxisti super me et super regnum meum peccatum grande quae non debuisti facere fecisti nobis
GEN|20|10|rursusque expostulans ait quid vidisti ut hoc faceres
GEN|20|11|respondit Abraham cogitavi mecum dicens forsitan non est timor Dei in loco isto et interficient me propter uxorem meam
GEN|20|12|alias autem et vere soror mea est filia patris mei et non filia matris meae et duxi eam uxorem
GEN|20|13|postquam autem eduxit me Deus de domo patris mei dixi ad eam hanc misericordiam facies mecum in omni loco ad quem ingrediemur dices quod frater tuus sim
GEN|20|14|tulit igitur Abimelech oves et boves et servos et ancillas et dedit Abraham reddiditque illi Sarram uxorem suam
GEN|20|15|et ait terra coram vobis est ubicumque tibi placuerit habita
GEN|20|16|Sarrae autem dixit ecce mille argenteos dedi fratri tuo hoc erit tibi in velamen oculorum ad omnes qui tecum sunt et quocumque perrexeris mementoque te deprehensam
GEN|20|17|orante autem Abraham sanavit Deus Abimelech et uxorem ancillasque eius et pepererunt
GEN|20|18|concluserat enim Deus omnem vulvam domus Abimelech propter Sarram uxorem Abraham
GEN|21|1|visitavit autem Dominus Sarram sicut promiserat et implevit quae locutus est
GEN|21|2|concepitque et peperit filium in senectute sua tempore quo praedixerat ei Deus
GEN|21|3|vocavitque Abraham nomen filii sui quem genuit ei Sarra Isaac
GEN|21|4|et circumcidit eum octavo die sicut praeceperat ei Deus
GEN|21|5|cum centum esset annorum hac quippe aetate patris natus est Isaac
GEN|21|6|dixitque Sarra risum fecit mihi Deus quicumque audierit conridebit mihi
GEN|21|7|rursumque ait quis auditurum crederet Abraham quod Sarra lactaret filium quem peperit ei iam seni
GEN|21|8|crevit igitur puer et ablactatus est fecitque Abraham grande convivium in die ablactationis eius
GEN|21|9|cumque vidisset Sarra filium Agar Aegyptiae ludentem dixit ad Abraham
GEN|21|10|eice ancillam hanc et filium eius non enim erit heres filius ancillae cum filio meo Isaac
GEN|21|11|dure accepit hoc Abraham pro filio suo
GEN|21|12|cui dixit Deus non tibi videatur asperum super puero et super ancilla tua omnia quae dixerit tibi Sarra audi vocem eius quia in Isaac vocabitur tibi semen
GEN|21|13|sed et filium ancillae faciam in gentem magnam quia semen tuum est
GEN|21|14|surrexit itaque Abraham mane et tollens panem et utrem aquae inposuit scapulae eius tradiditque puerum et dimisit eam quae cum abisset errabat in solitudine Bersabee
GEN|21|15|cumque consumpta esset aqua in utre abiecit puerum subter unam arborum quae ibi erant
GEN|21|16|et abiit seditque e regione procul quantum potest arcus iacere dixit enim non videbo morientem puerum et sedens contra levavit vocem suam et flevit
GEN|21|17|exaudivit autem Deus vocem pueri vocavitque angelus Domini Agar de caelo dicens quid agis Agar noli timere exaudivit enim Deus vocem pueri de loco in quo est
GEN|21|18|surge tolle puerum et tene manum illius quia in gentem magnam faciam eum
GEN|21|19|aperuitque oculos eius Deus quae videns puteum aquae abiit et implevit utrem deditque puero bibere
GEN|21|20|et fuit cum eo qui crevit et moratus est in solitudine et factus est iuvenis sagittarius
GEN|21|21|habitavitque in deserto Pharan et accepit illi mater sua uxorem de terra Aegypti
GEN|21|22|eodem tempore dixit Abimelech et Fichol princeps exercitus eius ad Abraham Deus tecum est in universis quae agis
GEN|21|23|iura ergo per Dominum ne noceas mihi et posteris meis stirpique meae sed iuxta misericordiam quam feci tibi facies mihi et terrae in qua versatus es advena
GEN|21|24|dixitque Abraham ego iurabo
GEN|21|25|et increpavit Abimelech propter puteum aquae quem vi abstulerant servi illius
GEN|21|26|respondit Abimelech nescivi quis fecerit hanc rem sed et tu non indicasti mihi et ego non audivi praeter hodie
GEN|21|27|tulit itaque Abraham oves et boves et dedit Abimelech percusseruntque ambo foedus
GEN|21|28|et statuit Abraham septem agnas gregis seorsum
GEN|21|29|cui dixit Abimelech quid sibi volunt septem agnae istae quas stare fecisti seorsum
GEN|21|30|at ille septem inquit agnas accipies de manu mea ut sint in testimonium mihi quoniam ego fodi puteum istum
GEN|21|31|idcirco vocatus est locus ille Bersabee quia ibi uterque iuraverunt
GEN|21|32|et inierunt foedus pro puteo Iuramenti
GEN|21|33|surrexit autem Abimelech et Fichol princeps militiae eius reversique sunt in terram Palestinorum Abraham vero plantavit nemus in Bersabee et invocavit ibi nomen Domini Dei aeterni
GEN|21|34|et fuit colonus terrae Philisthinorum diebus multis
GEN|22|1|quae postquam gesta sunt temptavit Deus Abraham et dixit ad eum Abraham ille respondit adsum
GEN|22|2|ait ei tolle filium tuum unigenitum quem diligis Isaac et vade in terram Visionis atque offer eum ibi holocaustum super unum montium quem monstravero tibi
GEN|22|3|igitur Abraham de nocte consurgens stravit asinum suum ducens secum duos iuvenes et Isaac filium suum cumque concidisset ligna in holocaustum abiit ad locum quem praeceperat ei Deus
GEN|22|4|die autem tertio elevatis oculis vidit locum procul
GEN|22|5|dixitque ad pueros suos expectate hic cum asino ego et puer illuc usque properantes postquam adoraverimus revertemur ad vos
GEN|22|6|tulit quoque ligna holocausti et inposuit super Isaac filium suum ipse vero portabat in manibus ignem et gladium cumque duo pergerent simul
GEN|22|7|dixit Isaac patri suo pater mi at ille respondit quid vis fili ecce inquit ignis et ligna ubi est victima holocausti
GEN|22|8|dixit Abraham Deus providebit sibi victimam holocausti fili mi pergebant ergo pariter
GEN|22|9|veneruntque ad locum quem ostenderat ei Deus in quo aedificavit altare et desuper ligna conposuit cumque conligasset Isaac filium suum posuit eum in altari super struem lignorum
GEN|22|10|extenditque manum et arripuit gladium ut immolaret filium
GEN|22|11|et ecce angelus Domini de caelo clamavit dicens Abraham Abraham qui respondit adsum
GEN|22|12|dixitque ei non extendas manum tuam super puerum neque facias illi quicquam nunc cognovi quod timeas Dominum et non peperceris filio tuo unigenito propter me
GEN|22|13|levavit Abraham oculos viditque post tergum arietem inter vepres herentem cornibus quem adsumens obtulit holocaustum pro filio
GEN|22|14|appellavitque nomen loci illius Dominus videt unde usque hodie dicitur in monte Dominus videbit
GEN|22|15|vocavit autem angelus Domini Abraham secundo de caelo dicens
GEN|22|16|per memet ipsum iuravi dicit Dominus quia fecisti rem hanc et non pepercisti filio tuo unigenito
GEN|22|17|benedicam tibi et multiplicabo semen tuum sicut stellas caeli et velut harenam quae est in litore maris possidebit semen tuum portas inimicorum suorum
GEN|22|18|et benedicentur in semine tuo omnes gentes terrae quia oboedisti voci meae
GEN|22|19|reversus est Abraham ad pueros suos abieruntque Bersabee simul et habitavit ibi
GEN|22|20|his itaque gestis nuntiatum est Abraham quod Melcha quoque genuisset filios Nahor fratri suo
GEN|22|21|Hus primogenitum et Buz fratrem eius Camuhel patrem Syrorum
GEN|22|22|et Chased et Azau Pheldas quoque et Iedlaph
GEN|22|23|ac Bathuel de quo nata est Rebecca octo istos genuit Melcha Nahor fratri Abraham
GEN|22|24|concubina vero illius nomine Roma peperit Tabee et Gaom et Thaas et Maacha
GEN|23|1|vixit autem Sarra centum viginti septem annis
GEN|23|2|et mortua est in civitate Arbee quae est Hebron in terra Chanaan venitque Abraham ut plangeret et fleret eam
GEN|23|3|cumque surrexisset ab officio funeris locutus est ad filios Heth dicens
GEN|23|4|advena sum et peregrinus apud vos date mihi ius sepulchri vobiscum ut sepeliam mortuum meum
GEN|23|5|responderuntque filii Heth
GEN|23|6|audi nos domine princeps Dei es apud nos in electis sepulchris nostris sepeli mortuum tuum nullusque prohibere te poterit quin in monumento eius sepelias mortuum tuum
GEN|23|7|surrexit Abraham et adoravit populum terrae filios videlicet Heth
GEN|23|8|dixitque ad eos si placet animae vestrae ut sepeliam mortuum meum audite me et intercedite apud Ephron filium Soor
GEN|23|9|ut det mihi speluncam duplicem quam habet in extrema parte agri sui pecunia digna tradat mihi eam coram vobis in possessionem sepulchri
GEN|23|10|habitabat autem Ephron in medio filiorum Heth responditque ad Abraham cunctis audientibus qui ingrediebantur portam civitatis illius dicens
GEN|23|11|nequaquam ita fiat domine mi sed magis ausculta quod loquor agrum trado tibi et speluncam quae in eo est praesentibus filiis populi mei sepeli mortuum tuum
GEN|23|12|adoravit Abraham coram populo terrae
GEN|23|13|et locutus est ad Ephron circumstante plebe quaeso ut audias me dabo pecuniam pro agro suscipe eam et sic sepeliam mortuum meum in eo
GEN|23|14|respondit Ephron
GEN|23|15|domine mi audi terram quam postulas quadringentis argenti siclis valet istud est pretium inter me et te sed quantum est hoc sepeli mortuum tuum
GEN|23|16|quod cum audisset Abraham adpendit pecuniam quam Ephron postulaverat audientibus filiis Heth quadringentos siclos argenti et probati monetae publicae
GEN|23|17|confirmatusque est ager quondam Ephronis in quo erat spelunca duplex respiciens Mambre tam ipse quam spelunca et omnes arbores eius in cunctis terminis per circuitum
GEN|23|18|Abrahae in possessionem videntibus filiis Heth et cunctis qui intrabant portam civitatis illius
GEN|23|19|atque ita sepelivit Abraham Sarram uxorem suam in spelunca agri duplici qui respiciebat Mambre haec est Hebron in terra Chanaan
GEN|23|20|et confirmatus est ager et antrum quod erat in eo Abrahae in possessionem monumenti a filiis Heth
GEN|24|1|erat autem Abraham senex dierumque multorum et Dominus in cunctis benedixerat ei
GEN|24|2|dixitque ad servum seniorem domus suae qui praeerat omnibus quae habebat pone manum tuam subter femur meum
GEN|24|3|ut adiurem te per Dominum Deum caeli et terrae ut non accipias uxorem filio meo de filiabus Chananeorum inter quos habito
GEN|24|4|sed ad terram et ad cognationem meam proficiscaris et inde accipias uxorem filio meo Isaac
GEN|24|5|respondit servus si noluerit mulier venire mecum in terram hanc num reducere debeo filium tuum ad locum de quo egressus es
GEN|24|6|dixit Abraham cave nequando reducas illuc filium meum
GEN|24|7|Dominus Deus caeli qui tulit me de domo patris mei et de terra nativitatis meae qui locutus est mihi et iuravit dicens semini tuo dabo terram hanc ipse mittet angelum suum coram te et accipies inde uxorem filio meo
GEN|24|8|sin autem noluerit mulier sequi te non teneberis iuramento filium tantum meum ne reducas illuc
GEN|24|9|posuit ergo servus manum sub femore Abraham domini sui et iuravit illi super sermone hoc
GEN|24|10|tulitque decem camelos de grege domini sui et abiit ex omnibus bonis eius portans secum profectusque perrexit Mesopotamiam ad urbem Nahor
GEN|24|11|cumque camelos fecisset accumbere extra oppidum iuxta puteum aquae vespere eo tempore quo solent mulieres egredi ad hauriendam aquam dixit
GEN|24|12|Domine Deus domini mei Abraham occurre obsecro hodie mihi et fac misericordiam cum domino meo Abraham
GEN|24|13|ecce ego sto propter fontem aquae et filiae habitatorum huius civitatis egredientur ad hauriendam aquam
GEN|24|14|igitur puella cui ego dixero inclina hydriam tuam ut bibam et illa responderit bibe quin et camelis tuis dabo potum ipsa est quam praeparasti servo tuo Isaac et per hoc intellegam quod feceris misericordiam cum domino meo
GEN|24|15|necdum intra se verba conpleverat et ecce Rebecca egrediebatur filia Bathuel filii Melchae uxoris Nahor fratris Abraham habens hydriam in scapula
GEN|24|16|puella decora nimis virgoque pulcherrima et incognita viro descenderat autem ad fontem et impleverat hydriam ac revertebatur
GEN|24|17|occurritque ei servus et ait pauxillum mihi ad sorbendum praebe aquae de hydria tua
GEN|24|18|quae respondit bibe domine mi celeriterque deposuit hydriam super ulnam suam et dedit ei potum
GEN|24|19|cumque ille bibisset adiecit quin et camelis tuis hauriam aquam donec cuncti bibant
GEN|24|20|effundensque hydriam in canalibus recurrit ad puteum ut hauriret aquam et haustam omnibus camelis dedit
GEN|24|21|ille autem contemplabatur eam tacitus scire volens utrum prosperum fecisset iter suum Dominus an non
GEN|24|22|postquam ergo biberunt cameli protulit vir inaures aureas adpendentes siclos duos et armillas totidem pondo siclorum decem
GEN|24|23|dixitque ad eam cuius es filia indica mihi est in domo patris tui locus ad manendum
GEN|24|24|quae respondit filia Bathuelis sum filii Melchae quem peperit Nahor
GEN|24|25|et addidit dicens palearum quoque et faeni plurimum est apud nos et locus spatiosus ad manendum
GEN|24|26|inclinavit se homo et adoravit Dominum
GEN|24|27|dicens benedictus Dominus Deus domini mei Abraham qui non abstulit misericordiam et veritatem suam a domino meo et recto me itinere perduxit in domum fratris domini mei
GEN|24|28|cucurrit itaque puella et nuntiavit in domum matris suae omnia quae audierat
GEN|24|29|habebat autem Rebecca fratrem nomine Laban qui festinus egressus est ad hominem ubi erat fons
GEN|24|30|cumque vidisset inaures et armillas in manibus sororis suae et audisset cuncta verba referentis haec locutus est mihi homo venit ad virum qui stabat iuxta camelos et propter fontem aquae
GEN|24|31|dixitque ad eum ingredere benedicte Domini cur foris stas praeparavi domum et locum camelis
GEN|24|32|et introduxit eum hospitium ac destravit camelos deditque paleas et faenum et aquam ad lavandos pedes camelorum et virorum qui venerant cum eo
GEN|24|33|et adpositus est in conspectu eius panis qui ait non comedam donec loquar sermones meos respondit ei loquere
GEN|24|34|at ille servus inquit Abraham sum
GEN|24|35|et Dominus benedixit domino meo valde magnificatusque est et dedit ei oves et boves argentum et aurum servos et ancillas camelos et asinos
GEN|24|36|et peperit Sarra uxor domini mei filium domino meo in senectute sua deditque illi omnia quae habuerat
GEN|24|37|et adiuravit me dominus meus dicens non accipies uxorem filio meo de filiabus Chananeorum in quorum terra habito
GEN|24|38|sed ad domum patris mei perges et de cognatione mea accipies uxorem filio meo
GEN|24|39|ego vero respondi domino meo quid si noluerit venire mecum mulier
GEN|24|40|Dominus ait in cuius conspectu ambulo mittet angelum suum tecum et diriget viam tuam accipiesque uxorem filio meo de cognatione mea et de domo patris mei
GEN|24|41|innocens eris a maledictione mea cum veneris ad propinquos meos et non dederint tibi
GEN|24|42|veni ergo hodie ad fontem et dixi Domine Deus domini mei Abraham si direxisti viam meam in qua nunc ambulo
GEN|24|43|ecce sto iuxta fontem aquae et virgo quae egredietur ad hauriendam aquam audierit a me da mihi pauxillum aquae ad bibendum ex hydria tua
GEN|24|44|et dixerit mihi et tu bibe et camelis tuis hauriam ipsa est mulier quam praeparavit Dominus filio domini mei
GEN|24|45|dum haec mecum tacitus volverem apparuit Rebecca veniens cum hydria quam portabat in scapula descenditque ad fontem et hausit aquam et aio ad eam da mihi paululum bibere
GEN|24|46|quae festina deposuit hydriam de umero et dixit mihi et tu bibe et camelis tuis potum tribuam bibi et adaquavit camelos
GEN|24|47|interrogavique eam et dixi cuius es filia quae respondit filia Bathuelis sum filii Nahor quem peperit illi Melcha suspendi itaque inaures ad ornandam faciem eius et armillas posui in manibus
GEN|24|48|pronusque adoravi Dominum benedicens Domino Deo domini mei Abraham qui perduxisset me recto itinere ut sumerem filiam fratris domini mei filio eius
GEN|24|49|quam ob rem si facitis misericordiam et veritatem cum domino meo indicate mihi sin autem aliud placet et hoc dicite ut vadam ad dextram sive ad sinistram
GEN|24|50|responderunt Laban et Bathuel a Domino egressus est sermo non possumus extra placitum eius quicquam aliud tecum loqui
GEN|24|51|en Rebecca coram te est tolle eam et proficiscere et sit uxor filii domini tui sicut locutus est Dominus
GEN|24|52|quod cum audisset puer Abraham adoravit in terra Dominum
GEN|24|53|prolatisque vasis argenteis et aureis ac vestibus dedit ea Rebeccae pro munere fratribus quoque eius et matri dona obtulit
GEN|24|54|initoque convivio vescentes pariter et bibentes manserunt ibi surgens autem mane locutus est puer dimittite me ut vadam ad dominum meum
GEN|24|55|responderunt fratres eius et mater maneat puella saltem decem dies apud nos et postea proficiscetur
GEN|24|56|nolite ait me retinere quia Dominus direxit viam meam dimittite me ut pergam ad dominum meum
GEN|24|57|dixerunt vocemus puellam et quaeramus ipsius voluntatem
GEN|24|58|cumque vocata venisset sciscitati sunt vis ire cum homine isto quae ait vadam
GEN|24|59|dimiserunt ergo eam et nutricem illius servumque Abraham et comites eius
GEN|24|60|inprecantes prospera sorori suae atque dicentes soror nostra es crescas in mille milia et possideat semen tuum portas inimicorum suorum
GEN|24|61|igitur Rebecca et puellae illius ascensis camelis secutae sunt virum qui festinus revertebatur ad dominum suum
GEN|24|62|eo tempore Isaac deambulabat per viam quae ducit ad puteum cuius nomen est Viventis et videntis habitabat enim in terra australi
GEN|24|63|et egressus fuerat ad meditandum in agro inclinata iam die cumque levasset oculos vidit camelos venientes procul
GEN|24|64|Rebecca quoque conspecto Isaac descendit de camelo
GEN|24|65|et ait ad puerum quis est ille homo qui venit per agrum in occursum nobis dixit ei ipse est dominus meus at illa tollens cito pallium operuit se
GEN|24|66|servus autem cuncta quae gesserat narravit Isaac
GEN|24|67|qui introduxit eam in tabernaculum Sarrae matris suae et accepit uxorem et in tantum dilexit ut dolorem qui ex morte matris acciderat temperaret
GEN|25|1|Abraham vero aliam duxit uxorem nomine Cetthuram
GEN|25|2|quae peperit ei Zamram et Iexan et Madan et Madian et Iesboch et Sue
GEN|25|3|Iexan quoque genuit Saba et Dadan filii Dadan fuerunt Assurim et Lathusim et Loommim
GEN|25|4|at vero ex Madian ortus est Epha et Opher et Enoch et Abida et Eldaa omnes hii filii Cetthurae
GEN|25|5|deditque Abraham cuncta quae possederat Isaac
GEN|25|6|filiis autem concubinarum largitus est munera et separavit eos ab Isaac filio suo dum adhuc ipse viveret ad plagam orientalem
GEN|25|7|fuerunt autem dies vitae eius centum septuaginta quinque anni
GEN|25|8|et deficiens mortuus est in senectute bona provectaeque aetatis et plenus dierum congregatusque est ad populum suum
GEN|25|9|et sepelierunt eum Isaac et Ismahel filii sui in spelunca duplici quae sita est in agro Ephron filii Soor Hetthei e regione Mambre
GEN|25|10|quem emerat a filiis Heth ibi sepultus est ipse et Sarra uxor eius
GEN|25|11|et post obitum illius benedixit Deus Isaac filio eius qui habitabat iuxta puteum nomine Viventis et videntis
GEN|25|12|hae sunt generationes Ismahel filii Abraham quem peperit ei Agar Aegyptia famula Sarrae
GEN|25|13|et haec nomina filiorum eius in vocabulis et generationibus suis primogenitus Ismahelis Nabaioth dein Cedar et Abdeel et Mabsam
GEN|25|14|Masma quoque et Duma et Massa
GEN|25|15|Adad et Thema Itur et Naphis et Cedma
GEN|25|16|isti sunt filii Ismahel et haec nomina per castella et oppida eorum duodecim principes tribuum suarum
GEN|25|17|anni vitae Ismahel centum triginta septem deficiens mortuus est et adpositus ad populum suum
GEN|25|18|habitavit autem ab Evila usque Sur quae respicit Aegyptum introeuntibus Assyrios coram cunctis fratribus suis obiit
GEN|25|19|hae quoque sunt generationes Isaac filii Abraham Abraham genuit Isaac
GEN|25|20|qui cum quadraginta esset annorum duxit uxorem Rebeccam filiam Bathuel Syri de Mesopotamiam sororem Laban
GEN|25|21|deprecatusque est Dominum pro uxore sua eo quod esset sterilis qui exaudivit eum et dedit conceptum Rebeccae
GEN|25|22|sed conlidebantur in utero eius parvuli quae ait si sic mihi futurum erat quid necesse fuit concipere perrexitque ut consuleret Dominum
GEN|25|23|qui respondens ait duae gentes in utero tuo sunt et duo populi ex ventre tuo dividentur populusque populum superabit et maior minori serviet
GEN|25|24|iam tempus pariendi venerat et ecce gemini in utero repperti sunt
GEN|25|25|qui primus egressus est rufus erat et totus in morem pellis hispidus vocatumque est nomen eius Esau protinus alter egrediens plantam fratris tenebat manu et idcirco appellavit eum Iacob
GEN|25|26|sexagenarius erat Isaac quando nati sunt parvuli
GEN|25|27|quibus adultis factus est Esau vir gnarus venandi et homo agricola Iacob autem vir simplex habitabat in tabernaculis
GEN|25|28|Isaac amabat Esau eo quod de venationibus illius vesceretur et Rebecca diligebat Iacob
GEN|25|29|coxit autem Iacob pulmentum ad quem cum venisset Esau de agro lassus
GEN|25|30|ait da mihi de coctione hac rufa quia oppido lassus sum quam ob causam vocatum est nomen eius Edom
GEN|25|31|cui dixit Iacob vende mihi primogenita tua
GEN|25|32|ille respondit en morior quid mihi proderunt primogenita
GEN|25|33|ait Iacob iura ergo mihi iuravit Esau et vendidit primogenita
GEN|25|34|et sic accepto pane et lentis edulio comedit et bibit et abiit parvipendens quod primogenita vendidisset
GEN|26|1|orta autem fame super terram post eam sterilitatem quae acciderat in diebus Abraham abiit Isaac ad Abimelech regem Palestinorum in Gerara
GEN|26|2|apparuitque ei Dominus et ait ne descendas in Aegyptum sed quiesce in terra quam dixero tibi
GEN|26|3|et peregrinare in ea eroque tecum et benedicam tibi tibi enim et semini tuo dabo universas regiones has conplens iuramentum quod spopondi Abraham patri tuo
GEN|26|4|et multiplicabo semen tuum sicut stellas caeli daboque posteris tuis universas regiones has et benedicentur in semine tuo omnes gentes terrae
GEN|26|5|eo quod oboedierit Abraham voci meae et custodierit praecepta et mandata mea et caerimonias legesque servaverit
GEN|26|6|mansit itaque Isaac in Geraris
GEN|26|7|qui cum interrogaretur a viris loci illius super uxore sua respondit soror mea est timuerat enim confiteri quod sibi esset sociata coniugio reputans ne forte interficerent eum propter illius pulchritudinem
GEN|26|8|cumque pertransissent dies plurimi et ibi demoraretur prospiciens Abimelech Palestinorum rex per fenestram vidit eum iocantem cum Rebecca uxore sua
GEN|26|9|et accersito ait perspicuum est quod uxor tua sit cur mentitus es sororem tuam esse respondit timui ne morerer propter eam
GEN|26|10|dixitque Abimelech quare inposuisti nobis potuit coire quispiam de populo cum uxore tua et induxeras super nos grande peccatum praecepitque omni populo dicens
GEN|26|11|qui tetigerit hominis huius uxorem morte morietur
GEN|26|12|seruit autem Isaac in terra illa et invenit in ipso anno centuplum benedixitque ei Dominus
GEN|26|13|et locupletatus est homo et ibat proficiens atque succrescens donec magnus vehementer effectus est
GEN|26|14|habuit quoque possessionem ovium et armentorum et familiae plurimum ob haec invidentes ei Palestini
GEN|26|15|omnes puteos quos foderant servi patris illius Abraham illo tempore obstruxerunt implentes humo
GEN|26|16|in tantum ut ipse Abimelech diceret ad Isaac recede a nobis quoniam potentior nostri factus es valde
GEN|26|17|et ille discedens veniret ad torrentem Gerarae habitaretque ibi
GEN|26|18|rursum fodit alios puteos quos foderant servi patris sui Abraham et quos illo mortuo olim obstruxerant Philisthim appellavitque eos hisdem nominibus quibus ante pater vocaverat
GEN|26|19|foderunt in torrente et reppererunt aquam vivam
GEN|26|20|sed et ibi iurgium fuit pastorum Gerarae adversum pastores Isaac dicentium nostra est aqua quam ob rem nomen putei ex eo quod acciderat vocavit Calumniam
GEN|26|21|foderunt et alium et pro illo quoque rixati sunt appellavitque eum Inimicitias
GEN|26|22|profectus inde fodit alium puteum pro quo non contenderunt itaque vocavit nomen illius Latitudo dicens nunc dilatavit nos Dominus et fecit crescere super terram
GEN|26|23|ascendit autem ex illo loco in Bersabee
GEN|26|24|ubi apparuit ei Dominus in ipsa nocte dicens ego sum Deus Abraham patris tui noli metuere quia tecum sum benedicam tibi et multiplicabo semen tuum propter servum meum Abraham
GEN|26|25|itaque aedificavit ibi altare et invocato nomine Domini extendit tabernaculum praecepitque servis suis ut foderent puteum
GEN|26|26|ad quem locum cum venissent de Geraris Abimelech et Ochozath amicus illius et Fichol dux militum
GEN|26|27|locutus est eis Isaac quid venistis ad me hominem quem odistis et expulistis a vobis
GEN|26|28|qui responderunt vidimus tecum esse Dominum et idcirco nunc diximus sit iuramentum inter nos et ineamus foedus
GEN|26|29|ut non facias nobis quicquam mali sicut et nos nihil tuorum adtigimus nec fecimus quod te laederet sed cum pace dimisimus auctum benedictione Domini
GEN|26|30|fecit ergo eis convivium et post cibum et potum
GEN|26|31|surgentes mane iuraverunt sibi mutuo dimisitque eos Isaac pacifice in locum suum
GEN|26|32|ecce autem venerunt in ipso die servi Isaac adnuntiantes ei de puteo quem foderant atque dicentes invenimus aquam
GEN|26|33|unde appellavit eum Abundantiam et nomen urbi inpositum est Bersabee usque in praesentem diem
GEN|26|34|Esau vero quadragenarius duxit uxores Iudith filiam Beeri Hetthei et Basemath filiam Helon eiusdem loci
GEN|26|35|quae ambae offenderant animum Isaac et Rebeccae
GEN|27|1|senuit autem Isaac et caligaverunt oculi eius et videre non poterat vocavitque Esau filium suum maiorem et dixit ei fili mi qui respondit adsum
GEN|27|2|cui pater vides inquit quod senuerim et ignorem diem mortis meae
GEN|27|3|sume arma tua faretram et arcum et egredere foras cumque venatu aliquid adprehenderis
GEN|27|4|fac mihi inde pulmentum sicut velle me nosti et adfer ut comedam et benedicat tibi anima mea antequam moriar
GEN|27|5|quod cum audisset Rebecca et ille abisset in agrum ut iussionem patris expleret
GEN|27|6|dixit filio suo Iacob audivi patrem tuum loquentem cum Esau fratre tuo et dicentem ei
GEN|27|7|adfer mihi venationem tuam et fac cibos ut comedam et benedicam tibi coram Domino antequam moriar
GEN|27|8|nunc ergo fili mi adquiesce consiliis meis
GEN|27|9|et pergens ad gregem adfer mihi duos hedos optimos ut faciam ex eis escas patri tuo quibus libenter vescitur
GEN|27|10|quas cum intuleris et comederit benedicat tibi priusquam moriatur
GEN|27|11|cui ille respondit nosti quod Esau frater meus homo pilosus sit et ego lenis
GEN|27|12|si adtractaverit me pater meus et senserit timeo ne putet sibi voluisse inludere et inducat super me maledictionem pro benedictione
GEN|27|13|ad quem mater in me sit ait ista maledictio fili mi tantum audi vocem meam et perge adferque quae dixi
GEN|27|14|abiit et adtulit deditque matri paravit illa cibos sicut noverat velle patrem illius
GEN|27|15|et vestibus Esau valde bonis quas apud se habebat domi induit eum
GEN|27|16|pelliculasque hedorum circumdedit manibus et colli nuda protexit
GEN|27|17|dedit pulmentum et panes quos coxerat tradidit
GEN|27|18|quibus inlatis dixit pater mi et ille respondit audio quis tu es fili mi
GEN|27|19|dixitque Iacob ego sum Esau primogenitus tuus feci sicut praecepisti mihi surge sede et comede de venatione mea ut benedicat mihi anima tua
GEN|27|20|rursum Isaac ad filium suum quomodo inquit tam cito invenire potuisti fili mi qui respondit voluntatis Dei fuit ut cito mihi occurreret quod volebam
GEN|27|21|dixitque Isaac accede huc ut tangam te fili mi et probem utrum tu sis filius meus Esau an non
GEN|27|22|accessit ille ad patrem et palpato eo dixit Isaac vox quidem vox Iacob est sed manus manus sunt Esau
GEN|27|23|et non cognovit eum quia pilosae manus similitudinem maioris expresserant benedicens ergo illi
GEN|27|24|ait tu es filius meus Esau respondit ego sum
GEN|27|25|at ille offer inquit mihi cibos de venatione tua fili mi ut benedicat tibi anima mea quos cum oblatos comedisset obtulit ei etiam vinum quo hausto
GEN|27|26|dixit ad eum accede ad me et da mihi osculum fili mi
GEN|27|27|accessit et osculatus est eum statimque ut sensit vestimentorum illius flagrantiam benedicens ait ecce odor filii mei sicut odor agri cui benedixit Dominus
GEN|27|28|det tibi Deus de rore caeli et de pinguedine terrae abundantiam frumenti et vini
GEN|27|29|et serviant tibi populi et adorent te tribus esto dominus fratrum tuorum et incurventur ante te filii matris tuae qui maledixerit tibi sit maledictus et qui benedixerit benedictionibus repleatur
GEN|27|30|vix Isaac sermonem impleverat et egresso Iacob foras venit Esau
GEN|27|31|coctosque de venatione cibos intulit patri dicens surge pater mi et comede de venatione filii tui ut benedicat mihi anima tua
GEN|27|32|dixitque illi Isaac quis enim es tu qui respondit ego sum primogenitus filius tuus Esau
GEN|27|33|expavit Isaac stupore vehementi et ultra quam credi potest admirans ait quis igitur ille est qui dudum captam venationem adtulit mihi et comedi ex omnibus priusquam tu venires benedixique ei et erit benedictus
GEN|27|34|auditis Esau sermonibus patris inrugiit clamore magno et consternatus ait benedic etiam mihi pater mi
GEN|27|35|qui ait venit germanus tuus fraudulenter et accepit benedictionem tuam
GEN|27|36|at ille subiunxit iuste vocatum est nomen eius Iacob subplantavit enim me en altera vice primogenita mea ante tulit et nunc secundo subripuit benedictionem meam rursumque ad patrem numquid non reservasti ait et mihi benedictionem
GEN|27|37|respondit Isaac dominum tuum illum constitui et omnes fratres eius servituti illius subiugavi frumento et vino stabilivi eum tibi post haec fili mi ultra quid faciam
GEN|27|38|cui Esau num unam inquit tantum benedictionem habes pater mihi quoque obsecro ut benedicas cumque heiulatu magno fleret
GEN|27|39|motus Isaac dixit ad eum in pinguedine terrae et in rore caeli desuper
GEN|27|40|erit benedictio tua vives gladio et fratri tuo servies tempusque veniet cum excutias et solvas iugum eius de cervicibus tuis
GEN|27|41|oderat ergo semper Esau Iacob pro benedictione qua benedixerat ei pater dixitque in corde suo veniant dies luctus patris mei ut occidam Iacob fratrem meum
GEN|27|42|nuntiata sunt haec Rebeccae quae mittens et vocans Iacob filium suum dixit ad eum ecce Esau frater tuus minatur ut occidat te
GEN|27|43|nunc ergo fili audi vocem meam et consurgens fuge ad Laban fratrem meum in Haran
GEN|27|44|habitabisque cum eo dies paucos donec requiescat furor fratris tui
GEN|27|45|et cesset indignatio eius obliviscaturque eorum quae fecisti in eum postea mittam et adducam te inde huc cur utroque orbabor filio in una die
GEN|27|46|dixit quoque Rebecca ad Isaac taedet me vitae meae propter filias Heth si acceperit Iacob uxorem de stirpe huius terrae nolo vivere
GEN|28|1|vocavit itaque Isaac Iacob et benedixit praecepitque ei dicens noli accipere coniugem de genere Chanaan
GEN|28|2|sed vade et proficiscere in Mesopotamiam Syriae ad domum Bathuel patrem matris tuae et accipe tibi inde uxorem de filiabus Laban avunculi tui
GEN|28|3|Deus autem omnipotens benedicat tibi et crescere te faciat atque multiplicet ut sis in turbas populorum
GEN|28|4|et det tibi benedictiones Abraham et semini tuo post te ut possideas terram peregrinationis tuae quam pollicitus est avo tuo
GEN|28|5|cumque dimisisset eum Isaac profectus venit in Mesopotamiam Syriae ad Laban filium Bathuel Syri fratrem Rebeccae matris suae
GEN|28|6|videns autem Esau quod benedixisset pater suus Iacob et misisset eum in Mesopotamiam Syriae ut inde uxorem duceret et quod post benedictionem praecepisset ei dicens non accipies coniugem de filiabus Chanaan
GEN|28|7|quodque oboediens Iacob parentibus isset in Syriam
GEN|28|8|probans quoque quod non libenter aspiceret filias Chanaan pater suus
GEN|28|9|ivit ad Ismahelem et duxit uxorem absque his quas prius habebat Maeleth filiam Ismahel filii Abraham sororem Nabaioth
GEN|28|10|igitur egressus Iacob de Bersabee pergebat Haran
GEN|28|11|cumque venisset ad quendam locum et vellet in eo requiescere post solis occubitum tulit de lapidibus qui iacebant et subponens capiti suo dormivit in eodem loco
GEN|28|12|viditque in somnis scalam stantem super terram et cacumen illius tangens caelum angelos quoque Dei ascendentes et descendentes per eam
GEN|28|13|et Dominum innixum scalae dicentem sibi ego sum Dominus Deus Abraham patris tui et Deus Isaac terram in qua dormis tibi dabo et semini tuo
GEN|28|14|eritque germen tuum quasi pulvis terrae dilataberis ad occidentem et orientem septentrionem et meridiem et benedicentur in te et in semine tuo cunctae tribus terrae
GEN|28|15|et ero custos tuus quocumque perrexeris et reducam te in terram hanc nec dimittam nisi conplevero universa quae dixi
GEN|28|16|cumque evigilasset Iacob de somno ait vere Dominus est in loco isto et ego nesciebam
GEN|28|17|pavensque quam terribilis inquit est locus iste non est hic aliud nisi domus Dei et porta caeli
GEN|28|18|surgens ergo mane tulit lapidem quem subposuerat capiti suo et erexit in titulum fundens oleum desuper
GEN|28|19|appellavitque nomen urbis Bethel quae prius Luza vocabatur
GEN|28|20|vovit etiam votum dicens si fuerit Deus mecum et custodierit me in via per quam ambulo et dederit mihi panem ad vescendum et vestem ad induendum
GEN|28|21|reversusque fuero prospere ad domum patris mei erit mihi Dominus in Deum
GEN|28|22|et lapis iste quem erexi in titulum vocabitur Domus Dei cunctorumque quae dederis mihi decimas offeram tibi
GEN|29|1|profectus ergo Iacob venit ad terram orientalem
GEN|29|2|et vidit puteum in agro tresque greges ovium accubantes iuxta eum nam ex illo adaquabantur pecora et os eius grandi lapide claudebatur
GEN|29|3|morisque erat ut cunctis ovibus congregatis devolverent lapidem et refectis gregibus rursum super os putei ponerent
GEN|29|4|dixitque ad pastores fratres unde estis qui responderunt de Haran
GEN|29|5|quos interrogans numquid ait nostis Laban filium Nahor dixerunt novimus
GEN|29|6|sanusne est inquit valet inquiunt et ecce Rahel filia eius venit cum grege suo
GEN|29|7|dixitque Iacob adhuc multum diei superest nec est tempus ut reducantur ad caulas greges date ante potum ovibus et sic ad pastum eas reducite
GEN|29|8|qui responderunt non possumus donec omnia pecora congregentur et amoveamus lapidem de ore putei ut adaquemus greges
GEN|29|9|adhuc loquebantur et ecce Rahel veniebat cum ovibus patris sui nam gregem ipsa pascebat
GEN|29|10|quam cum vidisset Iacob et sciret consobrinam suam ovesque Laban avunculi sui amovit lapidem quo puteus claudebatur
GEN|29|11|et adaquato grege osculatus est eam elevataque voce flevit
GEN|29|12|et indicavit ei quod frater esset patris eius et filius Rebeccae at illa festinans nuntiavit patri suo
GEN|29|13|qui cum audisset venisse Iacob filium sororis suae cucurrit obviam conplexusque eum et in oscula ruens duxit in domum suam auditis autem causis itineris
GEN|29|14|respondit os meum es et caro mea et postquam expleti sunt dies mensis unius
GEN|29|15|dixit ei num quia frater meus es gratis servies mihi dic quid mercedis accipias
GEN|29|16|habebat vero filias duas nomen maioris Lia minor appellabatur Rahel
GEN|29|17|sed Lia lippis erat oculis Rahel decora facie et venusto aspectu
GEN|29|18|quam diligens Iacob ait serviam tibi pro Rahel filia tua minore septem annis
GEN|29|19|respondit Laban melius est ut tibi eam dem quam viro alteri mane apud me
GEN|29|20|servivit igitur Iacob pro Rahel septem annis et videbantur illi pauci dies prae amoris magnitudine
GEN|29|21|dixitque ad Laban da mihi uxorem meam quia iam tempus expletum est ut ingrediar ad eam
GEN|29|22|qui vocatis multis amicorum turbis ad convivium fecit nuptias
GEN|29|23|et vespere filiam suam Liam introduxit ad eum
GEN|29|24|dans ancillam filiae Zelpham nomine ad quam cum ex more Iacob fuisset ingressus facto mane vidit Liam
GEN|29|25|et dixit ad socerum quid est quod facere voluisti nonne pro Rahel servivi tibi quare inposuisti mihi
GEN|29|26|respondit Laban non est in loco nostro consuetudinis ut minores ante tradamus ad nuptias
GEN|29|27|imple ebdomadem dierum huius copulae et hanc quoque dabo tibi pro opere quo serviturus es mihi septem annis aliis
GEN|29|28|adquievit placito et ebdomade transacta Rahel duxit uxorem
GEN|29|29|cui pater servam Balam dederat
GEN|29|30|tandemque potitus optatis nuptiis amorem sequentis priori praetulit serviens apud eum septem annis aliis
GEN|29|31|videns autem Dominus quod despiceret Liam aperuit vulvam eius sorore sterili permanente
GEN|29|32|quae conceptum genuit filium vocavitque nomen eius Ruben dicens vidit Dominus humilitatem meam nunc amabit me vir meus
GEN|29|33|rursumque concepit et peperit filium et ait quoniam audivit Dominus haberi me contemptui dedit etiam istum mihi vocavitque nomen illius Symeon
GEN|29|34|concepit tertio et genuit alium dixitque nunc quoque copulabitur mihi maritus meus eo quod pepererim illi tres filios et idcirco appellavit nomen eius Levi
GEN|29|35|quarto concepit et peperit filium et ait modo confitebor Domino et ob hoc vocavit eum Iudam cessavitque parere
GEN|30|1|cernens autem Rahel quod infecunda esset invidit sorori et ait marito suo da mihi liberos alioquin moriar
GEN|30|2|cui iratus respondit Iacob num pro Deo ego sum qui privavit te fructu ventris tui
GEN|30|3|at illa habeo inquit famulam Balam ingredere ad eam ut pariat super genua mea et habeam ex ea filios
GEN|30|4|deditque illi Balam in coniugium quae
GEN|30|5|ingresso ad se viro concepit et peperit filium
GEN|30|6|dixitque Rahel iudicavit mihi Dominus et exaudivit vocem meam dans mihi filium et idcirco appellavit nomen illius Dan
GEN|30|7|rursumque Bala concipiens peperit alterum
GEN|30|8|pro quo ait Rahel conparavit me Deus cum sorore mea et invalui vocavitque eum Nepthalim
GEN|30|9|sentiens Lia quod parere desisset Zelpham ancillam suam marito tradidit
GEN|30|10|qua post conceptum edente filium
GEN|30|11|dixit feliciter et idcirco vocavit nomen eius Gad
GEN|30|12|peperit quoque Zelpha alterum
GEN|30|13|dixitque Lia hoc pro beatitudine mea beatam quippe me dicent mulieres propterea appellavit eum Aser
GEN|30|14|egressus autem Ruben tempore messis triticeae in agro repperit mandragoras quos matri Liae detulit dixitque Rahel da mihi partem de mandragoris filii tui
GEN|30|15|illa respondit parumne tibi videtur quod praeripueris maritum mihi nisi etiam mandragoras filii mei tuleris ait Rahel dormiat tecum hac nocte pro mandragoris filii tui
GEN|30|16|redeuntique ad vesperam de agro Iacob egressa est in occursum Lia et ad me inquit intrabis quia mercede conduxi te pro mandragoris filii mei dormivit cum ea nocte illa
GEN|30|17|et exaudivit Deus preces eius concepitque et peperit filium quintum
GEN|30|18|et ait dedit Deus mercedem mihi quia dedi ancillam meam viro meo appellavitque nomen illius Isachar
GEN|30|19|rursum Lia concipiens peperit sextum filium
GEN|30|20|et ait ditavit me Deus dote bona etiam hac vice mecum erit maritus meus eo quod genuerim ei sex filios et idcirco appellavit nomen eius Zabulon
GEN|30|21|post quem peperit filiam nomine Dinam
GEN|30|22|recordatus quoque Dominus Rahelis exaudivit eam et aperuit vulvam illius
GEN|30|23|quae concepit et peperit filium dicens abstulit Deus obprobrium meum
GEN|30|24|et vocavit nomen illius Ioseph dicens addat mihi Dominus filium alterum
GEN|30|25|nato autem Ioseph dixit Iacob socero suo dimitte me ut revertar in patriam et ad terram meam
GEN|30|26|da mihi uxores et liberos meos pro quibus servivi tibi ut abeam tu nosti servitutem qua servivi tibi
GEN|30|27|ait ei Laban inveniam gratiam in conspectu tuo experimento didici quod benedixerit mihi Deus propter te
GEN|30|28|constitue mercedem tuam quam dem tibi
GEN|30|29|at ille respondit tu nosti quomodo servierim tibi et quanta in manibus meis fuerit possessio tua
GEN|30|30|modicum habuisti antequam venirem et nunc dives effectus es benedixitque tibi Dominus ad introitum meum iustum est igitur ut aliquando provideam etiam domui meae
GEN|30|31|dixitque Laban quid dabo tibi at ille ait nihil volo sed si feceris quod postulo iterum pascam et custodiam pecora tua
GEN|30|32|gyra omnes greges tuos et separa cunctas oves varias et sparso vellere et quodcumque furvum et maculosum variumque fuerit tam in ovibus quam in capris erit merces mea
GEN|30|33|respondebitque mihi cras iustitia mea quando placiti tempus advenerit coram te et omnia quae non fuerint varia et maculosa et furva tam in ovibus quam in capris furti me arguent
GEN|30|34|dixit Laban gratum habeo quod petis
GEN|30|35|et separavit in die illo capras et oves hircos et arietes varios atque maculosos cunctum autem gregem unicolorem id est albi et nigri velleris tradidit in manu filiorum suorum
GEN|30|36|et posuit spatium itineris inter se et generum dierum trium qui pascebat reliquos greges eius
GEN|30|37|tollens ergo Iacob virgas populeas virides et amigdalinas et ex platanis ex parte decorticavit eas detractisque corticibus in his quae spoliata fuerant candor apparuit illa vero quae integra erant viridia permanserunt atque in hunc modum color effectus est varius
GEN|30|38|posuitque eas in canalibus ubi effundebatur aqua ut cum venissent greges ad bibendum ante oculos haberent virgas et in aspectu earum conciperent
GEN|30|39|factumque est ut in ipso calore coitus oves intuerentur virgas et parerent maculosa et varia et diverso colore respersa
GEN|30|40|divisitque gregem Iacob et posuit virgas ante oculos arietum erant autem alba quaeque et nigra Laban cetera vero Iacob separatis inter se gregibus
GEN|30|41|igitur quando primo tempore ascendebantur oves ponebat Iacob virgas in canalibus aquarum ante oculos arietum et ovium ut in earum contemplatione conciperent
GEN|30|42|quando vero serotina admissura erat et conceptus extremus non ponebat eas factaque sunt ea quae erant serotina Laban et quae primi temporis Iacob
GEN|30|43|ditatusque est homo ultra modum et habuit greges multos ancillas et servos camelos et asinos
GEN|31|1|postquam autem audivit verba filiorum Laban dicentium tulit Iacob omnia quae fuerunt patris nostri et de illius facultate ditatus factus est inclitus
GEN|31|2|animadvertit quoque faciem Laban quod non esset erga se sicut heri et nudius tertius
GEN|31|3|maxime dicente sibi Domino revertere in terram patrum tuorum et ad generationem tuam eroque tecum
GEN|31|4|misit et vocavit Rahel et Liam in agrum ubi pascebat greges
GEN|31|5|dixitque eis video faciem patris vestri quod non sit erga me sicut heri et nudius tertius Deus autem patris mei fuit mecum
GEN|31|6|et ipsae nostis quod totis viribus meis servierim patri vestro
GEN|31|7|sed pater vester circumvenit me et mutavit mercedem meam decem vicibus et tamen non dimisit eum Deus ut noceret mihi
GEN|31|8|si quando dixit variae erunt mercedes tuae pariebant omnes oves varios fetus quando vero e contrario ait alba quaeque accipies pro mercede omnes greges alba pepererunt
GEN|31|9|tulitque Deus substantiam patris vestri et dedit mihi
GEN|31|10|postquam enim conceptus ovium tempus advenerat levavi oculos meos et vidi in somnis ascendentes mares super feminas varios et maculosos et diversorum colorum
GEN|31|11|dixitque angelus Dei ad me in somnis Iacob et ego respondi adsum
GEN|31|12|qui ait leva oculos tuos et vide universos masculos ascendentes super feminas varios respersos atque maculosos vidi enim omnia quae fecit tibi Laban
GEN|31|13|ego sum Deus Bethel ubi unxisti lapidem et votum vovisti mihi nunc ergo surge et egredere de terra hac revertens in terram nativitatis tuae
GEN|31|14|responderunt Rahel et Lia numquid habemus residui quicquam in facultatibus et hereditate domus patris nostri
GEN|31|15|nonne quasi alienas reputavit nos et vendidit comeditque pretium nostrum
GEN|31|16|sed Deus tulit opes patris nostri et nobis eas tradidit ac filiis nostris unde omnia quae praecepit fac
GEN|31|17|surrexit itaque Iacob et inpositis liberis et coniugibus suis super camelos abiit
GEN|31|18|tulitque omnem substantiam et greges et quicquid in Mesopotamiam quaesierat pergens ad Isaac patrem suum in terram Chanaan
GEN|31|19|eo tempore Laban ierat ad tondendas oves et Rahel furata est idola patris sui
GEN|31|20|noluitque Iacob confiteri socero quod fugeret
GEN|31|21|cumque abisset tam ipse quam omnia quae iuris eius erant et amne transmisso pergeret contra montem Galaad
GEN|31|22|nuntiatum est Laban die tertio quod fugeret Iacob
GEN|31|23|qui adsumptis fratribus suis persecutus est eum diebus septem et conprehendit in monte Galaad
GEN|31|24|viditque in somnis dicentem sibi Dominum cave ne quicquam aspere loquaris contra Iacob
GEN|31|25|iamque Iacob extenderat in monte tabernaculum cum ille consecutus eum cum fratribus suis in eodem monte Galaad fixit tentorium
GEN|31|26|et dixit ad Iacob quare ita egisti ut clam me abigeres filias meas quasi captivas gladio
GEN|31|27|cur ignorante me fugere voluisti nec indicare mihi ut prosequerer te cum gaudio et canticis et tympanis et cithara
GEN|31|28|non es passus ut oscularer filios meos ac filias stulte operatus es et nunc
GEN|31|29|valet quidem manus mea reddere tibi malum sed Deus patris vestri heri dixit mihi cave ne loquaris cum Iacob quicquam durius
GEN|31|30|esto ad tuos ire cupiebas et desiderio tibi erat domus patris tui cur furatus es deos meos
GEN|31|31|respondit Iacob quod inscio te profectus sum timui ne violenter auferres filias tuas
GEN|31|32|quod autem furti arguis apud quemcumque inveneris deos tuos necetur coram fratribus nostris scrutare quicquid tuorum apud me inveneris et aufer haec dicens ignorabat quod Rahel furata esset idola
GEN|31|33|ingressus itaque Laban tabernaculum Iacob et Liae et utriusque famulae non invenit cumque intrasset tentorium Rahelis
GEN|31|34|illa festinans abscondit idola subter stramen cameli et sedit desuper scrutantique omne tentorium et nihil invenienti
GEN|31|35|ait ne irascatur dominus meus quod coram te adsurgere nequeo quia iuxta consuetudinem feminarum nunc accidit mihi sic delusa sollicitudo quaerentis est
GEN|31|36|tumensque Iacob cum iurgio ait quam ob culpam meam et ob quod peccatum sic exarsisti post me
GEN|31|37|et scrutatus es omnem supellectilem meam quid invenisti de cuncta substantia domus tuae pone hic coram fratribus meis et fratribus tuis et iudicent inter me et te
GEN|31|38|idcirco viginti annis fui tecum oves tuae et caprae steriles non fuerunt arietes gregis tui non comedi
GEN|31|39|nec captum a bestia ostendi tibi ego damnum omne reddebam quicquid furto perierat a me exigebas
GEN|31|40|die noctuque aestu urebar et gelu fugiebat somnus ab oculis meis
GEN|31|41|sic per viginti annos in domo tua servivi tibi quattuordecim pro filiabus et sex pro gregibus tuis inmutasti quoque mercedem meam decem vicibus
GEN|31|42|nisi Deus patris mei Abraham et Timor Isaac adfuisset mihi forsitan modo nudum me dimisisses adflictionem meam et laborem manuum mearum respexit Deus et arguit te heri
GEN|31|43|respondit ei Laban filiae et filii et greges tui et omnia quae cernis mea sunt quid possum facere filiis et nepotibus meis
GEN|31|44|veni ergo et ineamus foedus ut sit testimonium inter me et te
GEN|31|45|tulit itaque Iacob lapidem et erexit illum in titulum
GEN|31|46|dixitque fratribus suis adferte lapides qui congregantes fecerunt tumulum comederuntque super eum
GEN|31|47|quem vocavit Laban tumulus Testis et Iacob acervum Testimonii uterque iuxta proprietatem linguae suae
GEN|31|48|dixitque Laban tumulus iste testis erit inter me et te hodie et idcirco appellatum est nomen eius Galaad id est tumulus Testis
GEN|31|49|intueatur Dominus et iudicet inter nos quando recesserimus a nobis
GEN|31|50|si adflixeris filias meas et si introduxeris uxores alias super eas nullus sermonis nostri testis est absque Deo qui praesens respicit
GEN|31|51|dixitque rursus ad Iacob en tumulus hic et lapis quem erexi inter me et te
GEN|31|52|testis erit tumulus inquam iste et lapis sint in testimonio si aut ego transiero illum pergens ad te aut tu praeterieris malum mihi cogitans
GEN|31|53|Deus Abraham et Deus Nahor iudicet inter nos Deus patris eorum iuravit Iacob per Timorem patris sui Isaac
GEN|31|54|immolatisque victimis in monte vocavit fratres suos ut ederent panem qui cum comedissent manserunt ibi
GEN|31|55|Laban vero de nocte consurgens osculatus est filios et filias suas et benedixit illis reversus in locum suum
GEN|32|1|Iacob quoque abiit itinere quo coeperat fueruntque ei obviam angeli Dei
GEN|32|2|quos cum vidisset ait castra Dei sunt haec et appellavit nomen loci illius Manaim id est Castra
GEN|32|3|misit autem et nuntios ante se ad Esau fratrem suum in terram Seir regionis Edom
GEN|32|4|praecepitque eis dicens sic loquimini domino meo Esau haec dicit frater tuus Iacob apud Laban peregrinatus sum et fui usque in praesentem diem
GEN|32|5|habeo boves et asinos oves et servos atque ancillas mittoque nunc legationem ad dominum meum ut inveniam gratiam in conspectu tuo
GEN|32|6|reversi sunt nuntii ad Iacob dicentes venimus ad Esau fratrem tuum et ecce properat in occursum tibi cum quadringentis viris
GEN|32|7|timuit Iacob valde et perterritus divisit populum qui secum erat greges quoque et oves et boves et camelos in duas turmas
GEN|32|8|dicens si venerit Esau ad unam turmam et percusserit eam alia turma quae reliqua est salvabitur
GEN|32|9|dixitque Iacob Deus patris mei Abraham et Deus patris mei Isaac Domine qui dixisti mihi revertere in terram tuam et in locum nativitatis tuae et benefaciam tibi
GEN|32|10|minor sum cunctis miserationibus et veritate quam explesti servo tuo in baculo meo transivi Iordanem istum et nunc cum duabus turmis regredior
GEN|32|11|erue me de manu fratris mei de manu Esau quia valde eum timeo ne forte veniens percutiat matrem cum filiis
GEN|32|12|tu locutus es quod bene mihi faceres et dilatares semen meum sicut harenam maris quae prae multitudine numerari non potest
GEN|32|13|cumque dormisset ibi nocte illa separavit de his quae habebat munera Esau fratri suo
GEN|32|14|capras ducentas hircos viginti oves ducentas arietes viginti
GEN|32|15|camelos fetas cum pullis suis triginta vaccas quadraginta et tauros viginti asinas viginti et pullos earum decem
GEN|32|16|et misit per manus servorum suorum singulos seorsum greges dixitque pueris suis antecedite me et sit spatium inter gregem et gregem
GEN|32|17|et praecepit priori dicens si obvium habueris Esau fratrem meum et interrogaverit te cuius es et quo vadis et cuius sunt ista quae sequeris
GEN|32|18|respondebis servi tui Iacob munera misit domino meo Esau ipse quoque post nos venit
GEN|32|19|similiter mandata dedit secundo ac tertio et cunctis qui sequebantur greges dicens hisdem verbis loquimini ad Esau cum inveneritis eum
GEN|32|20|et addetis ipse quoque servus tuus Iacob iter nostrum insequitur dixit enim placabo illum muneribus quae praecedunt et postea videbo forsitan propitiabitur mihi
GEN|32|21|praecesserunt itaque munera ante eum ipse vero mansit nocte illa in Castris
GEN|32|22|cumque mature surrexisset tulit duas uxores suas et totidem famulas cum undecim filiis et transivit vadum Iaboc
GEN|32|23|transductisque omnibus quae ad se pertinebant
GEN|32|24|remansit solus et ecce vir luctabatur cum eo usque mane
GEN|32|25|qui cum videret quod eum superare non posset tetigit nervum femoris eius et statim emarcuit
GEN|32|26|dixitque ad eum dimitte me iam enim ascendit aurora respondit non dimittam te nisi benedixeris mihi
GEN|32|27|ait ergo quod nomen est tibi respondit Iacob
GEN|32|28|at ille nequaquam inquit Iacob appellabitur nomen tuum sed Israhel quoniam si contra Deum fortis fuisti quanto magis contra homines praevalebis
GEN|32|29|interrogavit eum Iacob dic mihi quo appellaris nomine respondit cur quaeris nomen meum et benedixit ei in eodem loco
GEN|32|30|vocavitque Iacob nomen loci illius Phanuhel dicens vidi Deum facie ad faciem et salva facta est anima mea
GEN|32|31|ortusque est ei statim sol postquam transgressus est Phanuhel ipse vero claudicabat pede
GEN|32|32|quam ob causam non comedunt filii Israhel nervum qui emarcuit in femore Iacob usque in praesentem diem eo quod tetigerit nervum femoris eius et obstipuerit
GEN|33|1|levans autem Iacob oculos suos vidit venientem Esau et cum eo quadringentos viros divisitque filios Liae et Rahel ambarumque famularum
GEN|33|2|et posuit utramque ancillam et liberos earum in principio Liam vero et filios eius in secundo loco Rahel autem et Ioseph novissimos
GEN|33|3|et ipse praegrediens adoravit pronus in terram septies donec adpropinquaret frater eius
GEN|33|4|currens itaque Esau obviam fratri suo amplexatus est eum stringensque collum et osculans flevit
GEN|33|5|levatisque oculis vidit mulieres et parvulos earum et ait quid sibi volunt isti et si ad te pertinent respondit parvuli sunt quos donavit mihi Deus servo tuo
GEN|33|6|et adpropinquantes ancillae et filii earum incurvati sunt
GEN|33|7|accessitque Lia cum liberis suis et cum similiter adorassent extremi Ioseph et Rahel adoraverunt
GEN|33|8|quaenam sunt inquit istae turmae quas obvias habui respondit ut invenirem gratiam coram domino meo
GEN|33|9|et ille habeo ait plurima frater mi sint tua tibi
GEN|33|10|dixit Iacob noli ita obsecro sed si inveni gratiam in oculis tuis accipe munusculum de manibus meis sic enim vidi faciem tuam quasi viderim vultum Dei esto mihi propitius
GEN|33|11|et suscipe benedictionem quam adtuli tibi et quam donavit mihi Deus tribuens omnia vix fratre conpellente suscipiens
GEN|33|12|ait gradiamur simul eroque socius itineris tui
GEN|33|13|dixit Iacob nosti domine mi quod parvulos habeam teneros et oves ac boves fetas mecum quas si plus in ambulando fecero laborare morientur una die cuncti greges
GEN|33|14|praecedat dominus meus ante servum suum et ego sequar paulatim vestigia eius sicut videro posse parvulos meos donec veniam ad dominum meum in Seir
GEN|33|15|respondit Esau oro te ut de populo qui mecum est saltem socii remaneant viae tuae non est inquit necesse hoc uno indigeo ut inveniam gratiam in conspectu domini mei
GEN|33|16|reversus est itaque illo die Esau itinere quo venerat in Seir
GEN|33|17|et Iacob venit in Soccoth ubi aedificata domo et fixis tentoriis appellavit nomen loci illius Soccoth id est Tabernacula
GEN|33|18|transivitque in Salem urbem Sycimorum quae est in terra Chanaan postquam regressus est de Mesopotamiam Syriae et habitavit iuxta oppidum
GEN|33|19|emitque partem agri in qua fixerat tabernaculum a filiis Emor patris Sychem centum agnis
GEN|33|20|et erecto ibi altari invocavit super illud Fortissimum Deum Israhel
GEN|34|1|egressa est autem Dina filia Liae ut videret mulieres regionis illius
GEN|34|2|quam cum vidisset Sychem filius Emor Evei princeps terrae illius adamavit et rapuit et dormivit cum illa vi opprimens virginem
GEN|34|3|et conglutinata est anima eius cum ea tristemque blanditiis delinivit
GEN|34|4|et pergens ad Emor patrem suum accipe mihi inquit puellam hanc coniugem
GEN|34|5|quod cum audisset Iacob absentibus filiis et in pastu occupatis pecorum siluit donec redirent
GEN|34|6|egresso autem Emor patre Sychem ut loqueretur ad Iacob
GEN|34|7|ecce filii eius veniebant de agro auditoque quod acciderat irati sunt valde eo quod foedam rem esset operatus in Israhel et violata filia Iacob rem inlicitam perpetrasset
GEN|34|8|locutus est itaque Emor ad eos Sychem filii mei adhesit anima filiae vestrae date eam illi uxorem
GEN|34|9|et iungamus vicissim conubia filias vestras tradite nobis et filias nostras accipite
GEN|34|10|et habitate nobiscum terra in potestate vestra est exercete negotiamini et possidete eam
GEN|34|11|sed et Sychem ad patrem et ad fratres eius ait inveniam gratiam coram vobis et quaecumque statueritis dabo
GEN|34|12|augete dotem munera postulate libens tribuam quod petieritis tantum date mihi puellam hanc uxorem
GEN|34|13|responderunt filii Iacob Sychem et patri eius in dolo saevientes ob stuprum sororis
GEN|34|14|non possumus facere quod petitis nec dare sororem nostram homini incircumciso quod inlicitum et nefarium est apud nos
GEN|34|15|sed in hoc valebimus foederari si esse volueritis nostri similes et circumcidatur in vobis omne masculini sexus
GEN|34|16|tunc dabimus et accipiemus mutuo filias nostras ac vestras et habitabimus vobiscum erimusque unus populus
GEN|34|17|sin autem circumcidi nolueritis tollemus filiam nostram et recedemus
GEN|34|18|placuit oblatio eorum Emor et Sychem filio eius
GEN|34|19|nec distulit adulescens quin statim quod petebatur expleret amabat enim puellam valde et ipse erat inclitus in omni domo patris sui
GEN|34|20|ingressique portam urbis locuti sunt populo
GEN|34|21|viri isti pacifici sunt et volunt habitare nobiscum negotientur in terra et exerceant eam quae spatiosa et lata cultoribus indiget filias eorum accipiemus uxores et nostras illis dabimus
GEN|34|22|unum est quod differtur tantum bonum si circumcidamus masculos nostros ritum gentis imitantes
GEN|34|23|et substantia eorum et pecora et cuncta quae possident nostra erunt tantum in hoc adquiescamus et habitantes simul unum efficiemus populum
GEN|34|24|adsensi sunt omnes circumcisis cunctis maribus
GEN|34|25|et ecce die tertio quando gravissimus vulnerum dolor est arreptis duo Iacob filii Symeon et Levi fratres Dinae gladiis ingressi sunt urbem confidenter interfectisque omnibus masculis
GEN|34|26|Emor et Sychem pariter necaverunt tollentes Dinam de domo Sychem sororem suam
GEN|34|27|quibus egressis inruerunt super occisos ceteri filii Iacob et depopulati sunt urbem in ultionem stupri
GEN|34|28|oves eorum et armenta et asinos cunctaque vastantes quae in domibus et in agris erant
GEN|34|29|parvulos quoque et uxores eorum duxere captivas
GEN|34|30|quibus patratis audacter Iacob dixit ad Symeon et Levi turbastis me et odiosum fecistis Chananeis et Ferezeis habitatoribus terrae huius nos pauci sumus illi congregati percutient me et delebor ego et domus mea
GEN|34|31|responderunt numquid ut scorto abuti debuere sorore nostra
GEN|35|1|interea locutus est Deus ad Iacob surge et ascende Bethel et habita ibi facque altare Deo qui apparuit tibi quando fugiebas Esau fratrem tuum
GEN|35|2|Iacob vero convocata omni domo sua ait abicite deos alienos qui in medio vestri sunt et mundamini ac mutate vestimenta vestra
GEN|35|3|surgite et ascendamus in Bethel ut faciamus ibi altare Deo qui exaudivit me in die tribulationis meae et fuit socius itineris mei
GEN|35|4|dederunt ergo ei omnes deos alienos quos habebant et inaures quae erant in auribus eorum at ille infodit ea subter terebinthum quae est post urbem Sychem
GEN|35|5|cumque profecti essent terror Dei invasit omnes per circuitum civitates et non sunt ausi persequi recedentes
GEN|35|6|venit igitur Iacob Luzam quae est in terra Chanaan cognomento Bethel ipse et omnis populus cum eo
GEN|35|7|aedificavitque ibi altare et appellavit nomen loci Domus Dei ibi enim apparuit ei Deus cum fugeret fratrem suum
GEN|35|8|eodem tempore mortua est Debbora nutrix Rebeccae et sepulta ad radices Bethel subter quercum vocatumque est nomen loci quercus Fletus
GEN|35|9|apparuit autem iterum Deus Iacob postquam reversus est de Mesopotamiam Syriae benedixitque ei
GEN|35|10|dicens non vocaberis ultra Iacob sed Israhel erit nomen tuum et appellavit eum Israhel
GEN|35|11|dixitque ei ego Deus omnipotens cresce et multiplicare gentes et populi nationum erunt ex te reges de lumbis tuis egredientur
GEN|35|12|terramque quam dedi Abraham et Isaac dabo tibi et semini tuo post te
GEN|35|13|et recessit ab eo
GEN|35|14|ille vero erexit titulum lapideum in loco quo locutus ei fuerat Deus libans super eum libamina et effundens oleum
GEN|35|15|vocansque nomen loci Bethel
GEN|35|16|egressus inde venit verno tempore ad terram quae ducit Efratham in qua cum parturiret Rahel
GEN|35|17|ob difficultatem partus periclitari coepit dixitque ei obsetrix noli timere quia et hunc habebis filium
GEN|35|18|egrediente autem anima prae dolore et inminente iam morte vocavit nomen filii sui Benoni id est filius doloris mei pater vero appellavit eum Beniamin id est filius dexterae
GEN|35|19|mortua est ergo Rahel et sepulta in via quae ducit Efratham haec est Bethleem
GEN|35|20|erexitque Iacob titulum super sepulchrum eius hic est titulus monumenti Rahel usque in praesentem diem
GEN|35|21|egressus inde fixit tabernaculum trans turrem Gregis
GEN|35|22|cumque habitaret in illa regione abiit Ruben et dormivit cum Bala concubina patris sui quod illum minime latuit erant autem filii Iacob duodecim
GEN|35|23|filii Liae primogenitus Ruben et Symeon et Levi et Iudas et Isachar et Zabulon
GEN|35|24|filii Rahel Ioseph et Beniamin
GEN|35|25|filii Balae ancillae Rahelis Dan et Nepthalim
GEN|35|26|filii Zelphae ancillae Liae Gad et Aser hii filii Iacob qui nati sunt ei in Mesopotamiam Syriae
GEN|35|27|venit etiam ad Isaac patrem suum in Mambre civitatem Arbee haec est Hebron in qua peregrinatus est Abraham et Isaac
GEN|35|28|et conpleti sunt dies Isaac centum octoginta annorum
GEN|35|29|consumptusque aetate mortuus est et adpositus populo suo senex et plenus dierum et sepelierunt eum Esau et Iacob filii sui
GEN|36|1|hae sunt autem generationes Esau ipse est Edom
GEN|36|2|Esau accepit uxores de filiabus Chanaan Ada filiam Elom Hetthei et Oolibama filiam Anae filiae Sebeon Evei
GEN|36|3|Basemath quoque filiam Ismahel sororem Nabaioth
GEN|36|4|peperit autem Ada Eliphaz Basemath genuit Rauhel
GEN|36|5|Oolibama edidit Hieus et Hielom et Core hii filii Esau qui nati sunt ei in terra Chanaan
GEN|36|6|tulit autem Esau uxores suas et filios et filias et omnem animam domus suae et substantiam et pecora et cuncta quae habere poterat in terra Chanaan et abiit in alteram regionem recessitque a fratre suo Iacob
GEN|36|7|divites enim erant valde et simul habitare non poterant nec sustinebat eos terra peregrinationis eorum prae multitudine gregum
GEN|36|8|habitavitque Esau in monte Seir ipse est Edom
GEN|36|9|hae sunt generationes Esau patris Edom in monte Seir
GEN|36|10|et haec nomina filiorum eius Eliphaz filius Ada uxoris Esau Rauhel quoque filius Basemath uxoris eius
GEN|36|11|fueruntque filii Eliphaz Theman Omar Sephu et Gatham et Cenez
GEN|36|12|erat autem Thamna concubina Eliphaz filii Esau quae peperit ei Amalech hii sunt filii Adae uxoris Esau
GEN|36|13|filii autem Rauhel Naath et Zara Semma et Meza hii filii Basemath uxoris Esau
GEN|36|14|isti quoque erant filii Oolibama filiae Ana filiae Sebeon uxoris Esau quos genuit ei Hieus et Hielom et Core
GEN|36|15|hii duces filiorum Esau filii Eliphaz primogeniti Esau dux Theman dux Omar dux Sephu dux Cenez
GEN|36|16|dux Core dux Gatham dux Amalech hii filii Eliphaz in terra Edom et hii filii Adae
GEN|36|17|hii quoque filii Rauhel filii Esau dux Naath dux Zara dux Semma dux Meza hii duces Rauhel in terra Edom isti filii Basemath uxoris Esau
GEN|36|18|hii autem filii Oolibama uxoris Esau dux Hieus dux Hielom dux Core hii duces Oolibama filiae Ana uxoris Esau
GEN|36|19|isti filii Esau et hii duces eorum ipse est Edom
GEN|36|20|isti filii Seir Horrei habitatores terrae Lotham et Sobal et Sebeon et Anan
GEN|36|21|Dison et Eser et Disan hii duces Horrei filii Seir in terra Edom
GEN|36|22|facti sunt autem filii Lotham Horrei et Heman erat autem soror Lotham Thamna
GEN|36|23|et isti filii Sobal Alvam et Maneeth et Hebal Sephi et Onam
GEN|36|24|et hii filii Sebeon Ahaia et Anam iste est Ana qui invenit aquas calidas in solitudine cum pasceret asinos Sebeon patris sui
GEN|36|25|habuitque filium Disan et filiam Oolibama
GEN|36|26|et isti filii Disan Amdan et Esban et Iethran et Charan
GEN|36|27|hii quoque filii Eser Balaan et Zevan et Acham
GEN|36|28|habuit autem filios Disan Hus et Aran
GEN|36|29|isti duces Horreorum dux Lothan dux Sobal dux Sebeon dux Ana
GEN|36|30|dux Dison dux Eser dux Disan isti duces Horreorum qui imperaverunt in terra Seir
GEN|36|31|reges autem qui regnaverunt in terra Edom antequam haberent regem filii Israhel fuerunt hii
GEN|36|32|Bale filius Beor nomenque urbis eius Denaba
GEN|36|33|mortuus est autem Bale et regnavit pro eo Iobab filius Zare de Bosra
GEN|36|34|cumque mortuus esset Iobab regnavit pro eo Husan de terra Themanorum
GEN|36|35|hoc quoque mortuo regnavit pro eo Adad filius Badadi qui percussit Madian in regione Moab et nomen urbis eius Ahuith
GEN|36|36|cumque mortuus esset Adad regnavit pro eo Semla de Maserecha
GEN|36|37|hoc quoque mortuo regnavit pro eo Saul de fluvio Rooboth
GEN|36|38|cumque et hic obisset successit in regnum Baalanam filius Achobor
GEN|36|39|isto quoque mortuo regnavit pro eo Adad nomenque urbis eius Phau et appellabatur uxor illius Meezabel filia Matred filiae Mizaab
GEN|36|40|haec ergo nomina Esau in cognationibus et locis et vocabulis suis dux Thamna dux Alva dux Ietheth
GEN|36|41|dux Oolibama dux Ela dux Phinon
GEN|36|42|dux Cenez dux Theman dux Mabsar
GEN|36|43|dux Mabdiel dux Iram hii duces Edom habitantes in terra imperii sui ipse est Esau pater Idumeorum
GEN|37|1|habitavit autem Iacob in terra Chanaan in qua peregrinatus est pater suus
GEN|37|2|et hae sunt generationes eius Ioseph cum sedecim esset annorum pascebat gregem cum fratribus suis adhuc puer et erat cum filiis Balae et Zelphae uxorum patris sui accusavitque fratres suos apud patrem crimine pessimo
GEN|37|3|Israhel autem diligebat Ioseph super omnes filios suos eo quod in senectute genuisset eum fecitque ei tunicam polymitam
GEN|37|4|videntes autem fratres eius quod a patre plus cunctis filiis amaretur oderant eum nec poterant ei quicquam pacificum loqui
GEN|37|5|accidit quoque ut visum somnium referret fratribus quae causa maioris odii seminarium fuit
GEN|37|6|dixitque ad eos audite somnium meum quod vidi
GEN|37|7|putabam ligare nos manipulos in agro et quasi consurgere manipulum meum et stare vestrosque manipulos circumstantes adorare manipulum meum
GEN|37|8|responderunt fratres eius numquid rex noster eris aut subiciemur dicioni tuae haec ergo causa somniorum atque sermonum invidiae et odii fomitem ministravit
GEN|37|9|aliud quoque vidit somnium quod narrans fratribus ait vidi per somnium quasi solem et lunam et stellas undecim adorare me
GEN|37|10|quod cum patri suo et fratribus rettulisset increpavit eum pater et dixit quid sibi vult hoc somnium quod vidisti num ego et mater tua et fratres adorabimus te super terram
GEN|37|11|invidebant igitur ei fratres sui pater vero rem tacitus considerabat
GEN|37|12|cumque fratres illius in pascendis gregibus patris morarentur in Sychem
GEN|37|13|dixit ad eum Israhel fratres tui pascunt oves in Sycimis veni mittam te ad eos quo respondente
GEN|37|14|praesto sum ait vade et vide si cuncta prospera sint erga fratres tuos et pecora et renuntia mihi quid agatur missus de valle Hebron venit in Sychem
GEN|37|15|invenitque eum vir errantem in agro et interrogavit quid quaereret
GEN|37|16|at ille respondit fratres meos quaero indica mihi ubi pascant greges
GEN|37|17|dixitque ei vir recesserunt de loco isto audivi autem eos dicentes eamus in Dothain perrexit ergo Ioseph post fratres suos et invenit eos in Dothain
GEN|37|18|qui cum vidissent eum procul antequam accederet ad eos cogitaverunt illum occidere
GEN|37|19|et mutuo loquebantur ecce somniator venit
GEN|37|20|venite occidamus eum et mittamus in cisternam veterem dicemusque fera pessima devoravit eum et tunc apparebit quid illi prosint somnia sua
GEN|37|21|audiens hoc Ruben nitebatur liberare eum de manibus eorum et dicebat
GEN|37|22|non interficiamus animam eius nec effundatis sanguinem sed proicite eum in cisternam hanc quae est in solitudine manusque vestras servate innoxias hoc autem dicebat volens eripere eum de manibus eorum et reddere patri suo
GEN|37|23|confestim igitur ut pervenit ad fratres nudaverunt eum tunica talari et polymita
GEN|37|24|miseruntque in cisternam quae non habebat aquam
GEN|37|25|et sedentes ut comederent panem viderunt viatores Ismahelitas venire de Galaad et camelos eorum portare aromata et resinam et stacten in Aegyptum
GEN|37|26|dixit ergo Iudas fratribus suis quid nobis prodest si occiderimus fratrem nostrum et celaverimus sanguinem ipsius
GEN|37|27|melius est ut vendatur Ismahelitis et manus nostrae non polluantur frater enim et caro nostra est adquieverunt fratres sermonibus eius
GEN|37|28|et praetereuntibus Madianitis negotiatoribus extrahentes eum de cisterna vendiderunt Ismahelitis viginti argenteis qui duxerunt eum in Aegyptum
GEN|37|29|reversusque Ruben ad cisternam non invenit puerum
GEN|37|30|et scissis vestibus pergens ad fratres ait puer non conparet et ego quo ibo
GEN|37|31|tulerunt autem tunicam eius et in sanguinem hedi quem occiderant tinxerunt
GEN|37|32|mittentes qui ferrent ad patrem et dicerent hanc invenimus vide utrum tunica filii tui sit an non
GEN|37|33|quam cum agnovisset pater ait tunica filii mei est fera pessima comedit eum bestia devoravit Ioseph
GEN|37|34|scissisque vestibus indutus est cilicio lugens filium multo tempore
GEN|37|35|congregatis autem cunctis liberis eius ut lenirent dolorem patris noluit consolationem recipere et ait descendam ad filium meum lugens in infernum et illo perseverante in fletu
GEN|37|36|Madianei vendiderunt Ioseph in Aegypto Putiphar eunucho Pharaonis magistro militiae
GEN|38|1|eo tempore descendens Iudas a fratribus suis divertit ad virum odollamitem nomine Hiram
GEN|38|2|viditque ibi filiam hominis chananei vocabulo Suae et uxore accepta ingressus est ad eam
GEN|38|3|quae concepit et peperit filium vocavitque nomen eius Her
GEN|38|4|rursum concepto fetu natum filium nominavit Onam
GEN|38|5|tertium quoque peperit quem appellavit Sela quo nato parere ultra cessavit
GEN|38|6|dedit autem Iudas uxorem primogenito suo Her nomine Thamar
GEN|38|7|fuitque Her primogenitus Iudae nequam in conspectu Domini et ab eo occisus est
GEN|38|8|dixit ergo Iudas ad Onam filium suum ingredere ad uxorem fratris tui et sociare illi ut suscites semen fratri tuo
GEN|38|9|ille sciens non sibi nasci filios introiens ad uxorem fratris sui semen fundebat in terram ne liberi fratris nomine nascerentur
GEN|38|10|et idcirco percussit eum Dominus quod rem detestabilem faceret
GEN|38|11|quam ob rem dixit Iudas Thamar nurui suae esto vidua in domo patris tui donec crescat Sela filius meus timebat enim ne et ipse moreretur sicut fratres eius quae abiit et habitavit in domo patris sui
GEN|38|12|evolutis autem multis diebus mortua est filia Suae uxor Iudae qui post luctum consolatione suscepta ascendebat ad tonsores ovium suarum ipse et Hiras opilio gregis Odollamita in Thamnas
GEN|38|13|nuntiatumque est Thamar quod socer illius ascenderet in Thamnas ad tondendas oves
GEN|38|14|quae depositis viduitatis vestibus adsumpsit theristrum et mutato habitu sedit in bivio itineris quod ducit Thamnam eo quod crevisset Sela et non eum accepisset maritum
GEN|38|15|quam cum vidisset Iudas suspicatus est esse meretricem operuerat enim vultum suum ne cognosceretur
GEN|38|16|ingrediensque ad eam ait dimitte me ut coeam tecum nesciebat enim quod nurus sua esset qua respondente quid mihi dabis ut fruaris concubitu meo
GEN|38|17|dixit mittam tibi hedum de gregibus rursum illa dicente patiar quod vis si dederis mihi arrabonem donec mittas quod polliceris
GEN|38|18|ait Iudas quid vis tibi pro arrabone dari respondit anulum tuum et armillam et baculum quem manu tenes ad unum igitur coitum concepit mulier
GEN|38|19|et surgens abiit depositoque habitu quem adsumpserat induta est viduitatis vestibus
GEN|38|20|misit autem Iudas hedum per pastorem suum Odollamitem ut reciperet pignus quod dederat mulieri qui cum non invenisset eam
GEN|38|21|interrogavit homines loci illius ubi est mulier quae sedebat in bivio respondentibus cunctis non fuit in loco isto meretrix
GEN|38|22|reversus est ad Iudam et dixit ei non inveni eam sed et homines loci illius dixerunt mihi numquam ibi sedisse scortum
GEN|38|23|ait Iudas habeat sibi certe mendacii nos arguere non poterit ego misi hedum quem promiseram et tu non invenisti eam
GEN|38|24|ecce autem post tres menses nuntiaverunt Iudae dicentes fornicata est Thamar nurus tua et videtur uterus illius intumescere dixit Iudas producite eam ut conburatur
GEN|38|25|quae cum educeretur ad poenam misit ad socerum suum dicens de viro cuius haec sunt concepi cognosce cuius sit anulus et armilla et baculus
GEN|38|26|qui agnitis muneribus ait iustior me est quia non tradidi eam Sela filio meo attamen ultra non cognovit illam
GEN|38|27|instante autem partu apparuerunt gemini in utero atque in ipsa effusione infantum unus protulit manum in qua obsetrix ligavit coccinum dicens
GEN|38|28|iste egreditur prior
GEN|38|29|illo vero retrahente manum egressus est alter dixitque mulier quare divisa est propter te maceria et ob hanc causam vocavit nomen eius Phares
GEN|38|30|postea egressus est frater in cuius manu erat coccinum quem appellavit Zara
GEN|39|1|igitur Ioseph ductus est in Aegyptum emitque eum Putiphar eunuchus Pharaonis princeps exercitus vir aegyptius de manu Ismahelitarum a quibus perductus erat
GEN|39|2|fuitque Dominus cum eo et erat vir in cunctis prospere agens habitabatque in domo domini sui
GEN|39|3|qui optime noverat esse Dominum cum eo et omnia quae gereret ab eo dirigi in manu illius
GEN|39|4|invenitque Ioseph gratiam coram domino suo et ministrabat ei a quo praepositus omnibus gubernabat creditam sibi domum et universa quae tradita fuerant
GEN|39|5|benedixitque Dominus domui Aegyptii propter Ioseph et multiplicavit tam in aedibus quam in agris cunctam eius substantiam
GEN|39|6|nec quicquam aliud noverat nisi panem quo vescebatur erat autem Ioseph pulchra facie et decorus aspectu
GEN|39|7|post multos itaque dies iecit domina oculos suos in Ioseph et ait dormi mecum
GEN|39|8|qui nequaquam adquiescens operi nefario dixit ad eam ecce dominus meus omnibus mihi traditis ignorat quid habeat in domo sua
GEN|39|9|nec quicquam est quod non in mea sit potestate vel non tradiderit mihi praeter te quae uxor eius es quomodo ergo possum malum hoc facere et peccare in Deum meum
GEN|39|10|huiuscemodi verbis per singulos dies et mulier molesta erat adulescenti et ille recusabat stuprum
GEN|39|11|accidit autem ut quadam die intraret Ioseph domum et operis quippiam absque arbitris faceret
GEN|39|12|et illa adprehensa lacinia vestimenti eius diceret dormi mecum qui relicto in manu illius pallio fugit et egressus est foras
GEN|39|13|cumque vidisset mulier vestem in manibus suis et se esse contemptam
GEN|39|14|vocavit homines domus suae et ait ad eos en introduxit virum hebraeum ut inluderet nobis ingressus est ad me ut coiret mecum cumque ego succlamassem
GEN|39|15|et audisset vocem meam reliquit pallium quod tenebam et fugit foras
GEN|39|16|in argumentum ergo fidei retentum pallium ostendit marito revertenti domum
GEN|39|17|et ait ingressus est ad me servus hebraeus quem adduxisti ut inluderet mihi
GEN|39|18|cumque vidisset me clamare reliquit pallium et fugit foras
GEN|39|19|his auditis dominus et nimium credulus verbis coniugis iratus est valde
GEN|39|20|tradiditque Ioseph in carcerem ubi vincti regis custodiebantur et erat ibi clausus
GEN|39|21|fuit autem Dominus cum Ioseph et misertus illius dedit ei gratiam in conspectu principis carceris
GEN|39|22|qui tradidit in manu ipsius universos vinctos qui in custodia tenebantur et quicquid fiebat sub ipso erat
GEN|39|23|nec noverat aliquid cunctis ei creditis Dominus enim erat cum illo et omnia eius opera dirigebat
GEN|40|1|his ita gestis accidit ut peccarent duo eunuchi pincerna regis Aegypti et pistor domino suo
GEN|40|2|iratusque Pharao contra eos nam alter pincernis praeerat alter pistoribus
GEN|40|3|misit eos in carcerem principis militum in quo erat vinctus et Ioseph
GEN|40|4|at custos carceris tradidit eos Ioseph qui et ministrabat eis aliquantum temporis fluxerat et illi in custodia tenebantur
GEN|40|5|videruntque ambo somnium nocte una iuxta interpretationem congruam sibi
GEN|40|6|ad quos cum introisset Ioseph mane et vidisset eos tristes
GEN|40|7|sciscitatus est dicens cur tristior est hodie solito facies vestra
GEN|40|8|qui responderunt somnium vidimus et non est qui interpretetur nobis dixitque ad eos Ioseph numquid non Dei est interpretatio referte mihi quid videritis
GEN|40|9|narravit prior praepositus pincernarum somnium videbam coram me vitem
GEN|40|10|in qua erant tres propagines crescere paulatim gemmas et post flores uvas maturescere
GEN|40|11|calicemque Pharaonis in manu mea tuli ergo uvas et expressi in calicem quem tenebam et tradidi poculum Pharaoni
GEN|40|12|respondit Ioseph haec est interpretatio somnii tres propagines tres adhuc dies sunt
GEN|40|13|post quos recordabitur Pharao magisterii tui et restituet te in gradum pristinum dabisque ei calicem iuxta officium tuum sicut facere ante consueveras
GEN|40|14|tantum memento mei cum tibi bene fuerit et facies mecum misericordiam ut suggeras Pharaoni et educat me de isto carcere
GEN|40|15|quia furto sublatus sum de terra Hebraeorum et hic innocens in lacum missus sum
GEN|40|16|videns pistorum magister quod prudenter somnium dissolvisset ait et ego vidi somnium quod haberem tria canistra farinae super caput meum
GEN|40|17|et in uno canistro quod erat excelsius portare me omnes cibos qui fiunt arte pistoria avesque comedere ex eo
GEN|40|18|respondit Ioseph haec est interpretatio somnii tria canistra tres adhuc dies sunt
GEN|40|19|post quos auferet Pharao caput tuum ac suspendet te in cruce et lacerabunt volucres carnes tuas
GEN|40|20|exin dies tertius natalicius Pharaonis erat qui faciens grande convivium pueris suis recordatus est inter epulas magistri pincernarum et pistorum principis
GEN|40|21|restituitque alterum in locum suum ut porrigeret regi poculum
GEN|40|22|alterum suspendit in patibulo ut coniectoris veritas probaretur
GEN|40|23|et tamen succedentibus prosperis praepositus pincernarum oblitus est interpretis sui
GEN|41|1|post duos annos vidit Pharao somnium putabat se stare super fluvium
GEN|41|2|de quo ascendebant septem boves pulchrae et crassae nimis et pascebantur in locis palustribus
GEN|41|3|aliae quoque septem emergebant de flumine foedae confectaeque macie et pascebantur in ipsa amnis ripa in locis virentibus
GEN|41|4|devoraveruntque eas quarum mira species et habitudo corporum erat expergefactus Pharao
GEN|41|5|rursum dormivit et vidit alterum somnium septem spicae pullulabant in culmo uno plenae atque formonsae
GEN|41|6|aliae quoque totidem spicae tenues et percussae uredine oriebantur
GEN|41|7|devorantes omnem priorum pulchritudinem evigilans post quietem
GEN|41|8|et facto mane pavore perterritus misit ad coniectores Aegypti cunctosque sapientes et accersitis narravit somnium nec erat qui interpretaretur
GEN|41|9|tunc demum reminiscens pincernarum magister ait confiteor peccatum meum
GEN|41|10|iratus rex servis suis me et magistrum pistorum retrudi iussit in carcerem principis militum
GEN|41|11|ubi una nocte uterque vidimus somnium praesagum futurorum
GEN|41|12|erat ibi puer hebraeus eiusdem ducis militum famulus cui narrantes somnia
GEN|41|13|audivimus quicquid postea rei probavit eventus ego enim redditus sum officio meo et ille suspensus est in cruce
GEN|41|14|protinus ad regis imperium eductum de carcere Ioseph totonderunt ac veste mutata obtulerunt ei
GEN|41|15|cui ille ait vidi somnia nec est qui edisserat quae audivi te prudentissime conicere
GEN|41|16|respondit Ioseph absque me Deus respondebit prospera Pharaoni
GEN|41|17|narravit ergo ille quod viderat putabam me stare super ripam fluminis
GEN|41|18|et septem boves de amne conscendere pulchras nimis et obesis carnibus quae in pastu paludis virecta carpebant
GEN|41|19|et ecce has sequebantur aliae septem boves in tantum deformes et macilentae ut numquam tales in terra Aegypti viderim
GEN|41|20|quae devoratis et consumptis prioribus
GEN|41|21|nullum saturitatis dedere vestigium sed simili macie et squalore torpebant evigilans rursum sopore depressus
GEN|41|22|vidi somnium septem spicae pullulabant in culmo uno plenae atque pulcherrimae
GEN|41|23|aliae quoque septem tenues et percussae uredine oriebantur stipula
GEN|41|24|quae priorum pulchritudinem devorarunt narravi coniectoribus somnium et nemo est qui edisserat
GEN|41|25|respondit Ioseph somnium regis unum est quae facturus est Deus ostendit Pharaoni
GEN|41|26|septem boves pulchrae et septem spicae plenae septem ubertatis anni sunt eandemque vim somnii conprehendunt
GEN|41|27|septem quoque boves tenues atque macilentae quae ascenderunt post eas et septem spicae tenues et vento urente percussae septem anni sunt venturae famis
GEN|41|28|qui hoc ordine conplebuntur
GEN|41|29|ecce septem anni venient fertilitatis magnae in universa terra Aegypti
GEN|41|30|quos sequentur septem anni alii tantae sterilitatis ut oblivioni tradatur cuncta retro abundantia consumptura est enim fames omnem terram
GEN|41|31|et ubertatis magnitudinem perditura inopiae magnitudo
GEN|41|32|quod autem vidisti secundo ad eandem rem pertinens somnium firmitatis indicium est eo quod fiat sermo Dei et velocius impleatur
GEN|41|33|nunc ergo provideat rex virum sapientem et industrium et praeficiat eum terrae Aegypti
GEN|41|34|qui constituat praepositos per singulas regiones et quintam partem fructuum per septem annos fertilitatis
GEN|41|35|qui iam nunc futuri sunt congreget in horrea et omne frumentum sub Pharaonis potestate condatur serveturque in urbibus
GEN|41|36|et paretur futurae septem annorum fami quae pressura est Aegyptum et non consumetur terra inopia
GEN|41|37|placuit Pharaoni consilium et cunctis ministris eius
GEN|41|38|locutusque est ad eos num invenire poterimus talem virum qui spiritu Dei plenus sit
GEN|41|39|dixit ergo ad Ioseph quia ostendit Deus tibi omnia quae locutus es numquid sapientiorem et similem tui invenire potero
GEN|41|40|tu eris super domum meam et ad tui oris imperium cunctus populus oboediet uno tantum regni solio te praecedam
GEN|41|41|dicens quoque rursum Pharao ad Ioseph ecce constitui te super universam terram Aegypti
GEN|41|42|tulit anulum de manu sua et dedit in manu eius vestivitque eum stola byssina et collo torquem auream circumposuit
GEN|41|43|fecitque ascendere super currum suum secundum clamante praecone ut omnes coram eo genuflecterent et praepositum esse scirent universae terrae Aegypti
GEN|41|44|dixit quoque rex ad Ioseph ego sum Pharao absque tuo imperio non movebit quisquam manum aut pedem in omni terra Aegypti
GEN|41|45|vertitque nomen illius et vocavit eum lingua aegyptiaca Salvatorem mundi dedit quoque illi uxorem Aseneth filiam Putiphare sacerdotis Heliopoleos egressus itaque Ioseph ad terram Aegypti
GEN|41|46|triginta autem erat annorum quando stetit in conspectu regis Pharaonis circuivit omnes regiones Aegypti
GEN|41|47|venitque fertilitas septem annorum et in manipulos redactae segetes congregatae sunt in horrea Aegypti
GEN|41|48|omnis etiam frugum abundantia in singulis urbibus condita est
GEN|41|49|tantaque fuit multitudo tritici ut harenae maris coaequaretur et copia mensuram excederet
GEN|41|50|nati sunt autem Ioseph filii duo antequam veniret fames quos ei peperit Aseneth filia Putiphare sacerdotis Heliopoleos
GEN|41|51|vocavitque nomen primogeniti Manasse dicens oblivisci me fecit Deus omnium laborum meorum et domum patris mei
GEN|41|52|nomen quoque secundi appellavit Ephraim dicens crescere me fecit Deus in terra paupertatis meae
GEN|41|53|igitur transactis septem annis ubertatis qui fuerant in Aegypto
GEN|41|54|coeperunt venire septem anni inopiae quos praedixerat Ioseph et in universo orbe fames praevaluit in cuncta autem terra Aegypti erat panis
GEN|41|55|qua esuriente clamavit populus ad Pharaonem alimenta petens quibus ille respondit ite ad Ioseph et quicquid vobis dixerit facite
GEN|41|56|crescebat autem cotidie fames in omni terra aperuitque Ioseph universa horrea et vendebat Aegyptiis nam et illos oppresserat fames
GEN|41|57|omnesque provinciae veniebant in Aegyptum ut emerent escas et malum inopiae temperarent
GEN|42|1|audiens autem Iacob quod alimenta venderentur in Aegypto dixit filiis suis quare neglegitis
GEN|42|2|audivi quod triticum venundetur in Aegypto descendite et emite nobis necessaria ut possimus vivere et non consumamur inopia
GEN|42|3|descendentes igitur fratres Ioseph decem ut emerent frumenta in Aegypto
GEN|42|4|Beniamin domi retento ab Iacob qui dixerat fratribus eius ne forte in itinere quicquam patiatur mali
GEN|42|5|ingressi sunt terram Aegypti cum aliis qui pergebant ad emendum erat autem fames in terra Chanaan
GEN|42|6|et Ioseph princeps Aegypti atque ad illius nutum frumenta populis vendebantur cumque adorassent eum fratres sui
GEN|42|7|et agnovisset eos quasi ad alienos durius loquebatur interrogans eos unde venistis qui responderunt de terra Chanaan ut emamus victui necessaria
GEN|42|8|et tamen fratres ipse cognoscens non est agnitus ab eis
GEN|42|9|recordatusque somniorum quae aliquando viderat ait exploratores estis ut videatis infirmiora terrae venistis
GEN|42|10|qui dixerunt non est ita domine sed servi tui venerunt ut emerent cibos
GEN|42|11|omnes filii unius viri sumus pacifici venimus nec quicquam famuli tui machinantur mali
GEN|42|12|quibus ille respondit aliter est inmunita terrae huius considerare venistis
GEN|42|13|et illi duodecim inquiunt servi tui fratres sumus filii viri unius in terra Chanaan minimus cum patre nostro est alius non est super
GEN|42|14|hoc est ait quod locutus sum exploratores estis
GEN|42|15|iam nunc experimentum vestri capiam per salutem Pharaonis non egrediemini hinc donec veniat frater vester minimus
GEN|42|16|mittite e vobis unum et adducat eum vos autem eritis in vinculis donec probentur quae dixistis utrum falsa an vera sint alioquin per salutem Pharaonis exploratores estis
GEN|42|17|tradidit ergo eos custodiae tribus diebus
GEN|42|18|die autem tertio eductis de carcere ait facite quod dixi et vivetis Deum enim timeo
GEN|42|19|si pacifici estis frater vester unus ligetur in carcere vos autem abite et ferte frumenta quae emistis in domos vestras
GEN|42|20|et fratrem vestrum minimum ad me adducite ut possim vestros probare sermones et non moriamini fecerunt ut dixerat
GEN|42|21|et locuti sunt invicem merito haec patimur quia peccavimus in fratrem nostrum videntes angustiam animae illius cum deprecaretur nos et non audivimus idcirco venit super nos ista tribulatio
GEN|42|22|e quibus unus Ruben ait numquid non dixi vobis nolite peccare in puerum et non audistis me en sanguis eius exquiritur
GEN|42|23|nesciebant autem quod intellegeret Ioseph eo quod per interpretem loquebatur ad eos
GEN|42|24|avertitque se parumper et flevit et reversus locutus est ad eos
GEN|42|25|tollens Symeon et ligans illis praesentibus iussitque ministris ut implerent saccos eorum tritico et reponerent pecunias singulorum in sacculis suis datis supra cibariis in via qui fecerunt ita
GEN|42|26|at illi portantes frumenta in asinis profecti sunt
GEN|42|27|apertoque unus sacco ut daret iumento pabulum in diversorio contemplatus pecuniam in ore sacculi
GEN|42|28|dixit fratribus suis reddita est mihi pecunia en habetur in sacco et obstupefacti turbatique dixerunt mutuo quidnam est hoc quod fecit nobis Deus
GEN|42|29|veneruntque ad Iacob patrem suum in terra Chanaan et narraverunt ei omnia quae accidissent sibi dicentes
GEN|42|30|locutus est nobis dominus terrae dure et putavit nos exploratores provinciae
GEN|42|31|cui respondimus pacifici sumus nec ullas molimur insidias
GEN|42|32|duodecim fratres uno patre geniti sumus unus non est super minimus cum patre versatur in terra Chanaan
GEN|42|33|qui ait nobis sic probabo quod pacifici sitis fratrem vestrum unum dimittite apud me et cibaria domibus vestris necessaria sumite et abite
GEN|42|34|fratremque vestrum minimum adducite ad me ut sciam quod non sitis exploratores et istum qui tenetur in vinculis recipere possitis ac deinceps emendi quae vultis habeatis licentiam
GEN|42|35|his dictis cum frumenta effunderent singuli reppererunt in ore saccorum ligatas pecunias exterritisque simul omnibus
GEN|42|36|dixit pater Iacob absque liberis me esse fecistis Ioseph non est super Symeon tenetur in vinculis Beniamin auferetis in me haec mala omnia reciderunt
GEN|42|37|cui respondit Ruben duos filios meos interfice si non reduxero illum tibi trade in manu mea et ego eum restituam
GEN|42|38|at ille non descendet inquit filius meus vobiscum frater eius mortuus est ipse solus remansit si quid ei adversi acciderit in terra ad quam pergitis deducetis canos meos cum dolore ad inferos
GEN|43|1|interim fames omnem terram vehementer premebat
GEN|43|2|consumptisque cibis quos ex Aegypto detulerant dixit Iacob ad filios suos revertimini et emite pauxillum escarum
GEN|43|3|respondit Iudas denuntiavit nobis vir ille sub testificatione iurandi dicens non videbitis faciem meam nisi fratrem vestrum minimum adduxeritis vobiscum
GEN|43|4|si ergo vis mittere eum nobiscum pergemus pariter et ememus tibi necessaria
GEN|43|5|si autem non vis non ibimus vir enim ut saepe diximus denuntiavit nobis dicens non videbitis faciem meam absque fratre vestro minimo
GEN|43|6|dixit eis Israhel in meam hoc fecistis miseriam ut indicaretis ei et alium habere vos fratrem
GEN|43|7|at illi responderunt interrogavit nos homo per ordinem nostram progeniem si pater viveret si haberemus fratrem et nos respondimus ei consequenter iuxta id quod fuerat sciscitatus numquid scire poteramus quod dicturus esset adducite vobiscum fratrem vestrum
GEN|43|8|Iudas quoque dixit patri suo mitte puerum mecum ut proficiscamur et possimus vivere ne moriamur nos et parvuli nostri
GEN|43|9|ego suscipio puerum de manu mea require illum nisi reduxero et tradidero eum tibi ero peccati in te reus omni tempore
GEN|43|10|si non intercessisset dilatio iam vice altera venissemus
GEN|43|11|igitur Israhel pater eorum dixit ad eos si sic necesse est facite quod vultis sumite de optimis terrae fructibus in vasis vestris et deferte viro munera modicum resinae et mellis et styracis et stactes et terebinthi et amigdalarum
GEN|43|12|pecuniamque duplicem ferte vobiscum et illam quam invenistis in sacculis reportate ne forte errore factum sit
GEN|43|13|sed et fratrem vestrum tollite et ite ad virum
GEN|43|14|Deus autem meus omnipotens faciat vobis eum placabilem et remittat vobiscum fratrem vestrum quem tenet et hunc Beniamin ego autem quasi orbatus absque liberis ero
GEN|43|15|tulerunt ergo viri munera et pecuniam duplicem et Beniamin descenderuntque in Aegyptum et steterunt coram Ioseph
GEN|43|16|quos cum ille vidisset et Beniamin simul praecepit dispensatori domus suae dicens introduc viros domum et occide victimas et instrue convivium quoniam mecum sunt comesuri meridie
GEN|43|17|fecit ille sicut fuerat imperatum et introduxit viros domum
GEN|43|18|ibique exterriti dixerunt mutuo propter pecuniam quam rettulimus prius in saccis nostris introducti sumus ut devolvat in nos calumniam et violenter subiciat servituti et nos et asinos nostros
GEN|43|19|quam ob rem in ipsis foribus accedentes ad dispensatorem
GEN|43|20|locuti sunt oramus domine ut audias iam ante descendimus ut emeremus escas
GEN|43|21|quibus emptis cum venissemus ad diversorium aperuimus sacculos nostros et invenimus pecuniam in ore saccorum quam nunc eodem pondere reportamus
GEN|43|22|sed et aliud adtulimus argentum ut emamus quae necessaria sunt non est in nostra conscientia quis eam posuerit in marsuppiis nostris
GEN|43|23|at ille respondit pax vobiscum nolite timere Deus vester et Deus patris vestri dedit vobis thesauros in sacculis vestris nam pecuniam quam dedistis mihi probatam ego habeo eduxitque ad eos Symeon
GEN|43|24|et introductis domum adtulit aquam et laverunt pedes suos deditque pabula asinis eorum
GEN|43|25|illi vero parabant munera donec ingrederetur Ioseph meridie audierant enim quod ibi comesuri essent panem
GEN|43|26|igitur ingressus est Ioseph domum suam obtuleruntque ei munera tenentes in manibus et adoraverunt proni in terram
GEN|43|27|at ille clementer resalutatis eis interrogavit dicens salvusne est pater vester senex de quo dixeratis mihi adhuc vivit
GEN|43|28|qui responderunt sospes est servus tuus pater noster adhuc vivit et incurvati adoraverunt eum
GEN|43|29|adtollens autem oculos Ioseph vidit Beniamin fratrem suum uterinum et ait iste est frater vester parvulus de quo dixeratis mihi et rursum Deus inquit misereatur tui fili mi
GEN|43|30|festinavitque quia commota fuerant viscera eius super fratre suo et erumpebant lacrimae et introiens cubiculum flevit
GEN|43|31|rursusque lota facie egressus continuit se et ait ponite panes
GEN|43|32|quibus adpositis seorsum Ioseph et seorsum fratribus Aegyptiis quoque qui vescebantur simul seorsum inlicitum est enim Aegyptiis comedere cum Hebraeis et profanum putant huiuscemodi convivium
GEN|43|33|sederunt coram eo primogenitus iuxta primogenita sua et minimus iuxta aetatem suam et mirabantur nimis
GEN|43|34|sumptis partibus quas ab eo acceperant maiorque pars venit Beniamin ita ut quinque partibus excederet biberuntque et inebriati sunt cum eo
GEN|44|1|praecepit autem Ioseph dispensatori domus suae dicens imple saccos eorum frumento quantum possunt capere et pone pecuniam singulorum in summitate sacci
GEN|44|2|scyphum autem meum argenteum et pretium quod dedit tritici pone in ore sacci iunioris factumque est ita
GEN|44|3|et orto mane dimissi sunt cum asinis suis
GEN|44|4|iamque urbem exierant et processerant paululum tum Ioseph arcessito dispensatore domus surge inquit persequere viros et adprehensis dicito quare reddidistis malum pro bono
GEN|44|5|scyphum quem furati estis ipse est in quo bibit dominus meus et in quo augurari solet pessimam rem fecistis
GEN|44|6|fecit ille ut iusserat et adprehensis per ordinem locutus est
GEN|44|7|qui responderunt quare sic loquitur dominus noster ut servi tui tantum flagitii commiserint
GEN|44|8|pecuniam quam invenimus in summitate saccorum reportavimus ad te de terra Chanaan et quomodo consequens est ut furati simus de domo domini tui aurum vel argentum
GEN|44|9|apud quemcumque fuerit inventum servorum tuorum quod quaeris moriatur et nos servi erimus domini nostri
GEN|44|10|qui dixit fiat iuxta vestram sententiam apud quem fuerit inventum ipse sit servus meus vos autem eritis innoxii
GEN|44|11|itaque festinato deponentes in terram saccos aperuerunt singuli
GEN|44|12|quos scrutatus incipiens a maiore usque ad minimum invenit scyphum in sacco Beniamin
GEN|44|13|at illi scissis vestibus oneratisque rursum asinis reversi sunt in oppidum
GEN|44|14|primusque Iudas cum fratribus ingressus est ad Ioseph necdum enim de loco abierat omnesque ante eum in terra pariter corruerunt
GEN|44|15|quibus ille ait cur sic agere voluistis an ignoratis quod non sit similis mei in augurandi scientia
GEN|44|16|cui Iudas quid respondebimus inquit domino meo vel quid loquemur aut iusti poterimus obtendere Deus invenit iniquitatem servorum tuorum en omnes servi sumus domini mei et nos et apud quem inventus est scyphus
GEN|44|17|respondit Ioseph absit a me ut sic agam qui furatus est scyphum ipse sit servus meus vos autem abite liberi ad patrem vestrum
GEN|44|18|accedens propius Iudas confidenter ait oro domine mi loquatur servus tuus verbum in auribus tuis et ne irascaris famulo tuo tu es enim post Pharaonem
GEN|44|19|dominus meus interrogasti prius servos tuos habetis patrem aut fratrem
GEN|44|20|et nos respondimus tibi domino meo est nobis pater senex et puer parvulus qui in senecta illius natus est cuius uterinus frater est mortuus et ipsum solum habet mater sua pater vero tenere diligit eum
GEN|44|21|dixistique servis tuis adducite eum ad me et ponam oculos meos super illum
GEN|44|22|suggessimus domino meo non potest puer relinquere patrem suum si enim illum dimiserit morietur
GEN|44|23|et dixisti servis tuis nisi venerit frater vester minimus vobiscum non videbitis amplius faciem meam
GEN|44|24|cum ergo ascendissemus ad famulum tuum patrem nostrum narravimus ei omnia quae locutus est dominus meus
GEN|44|25|et dixit pater noster revertimini et emite nobis parum tritici
GEN|44|26|cui diximus ire non possumus si frater noster minimus descendet nobiscum proficiscemur simul alioquin illo absente non audemus videre faciem viri
GEN|44|27|atque ille respondit vos scitis quod duos genuerit mihi uxor mea
GEN|44|28|egressus est unus et dixistis bestia devoravit eum et hucusque non conparet
GEN|44|29|si tuleritis et istum et aliquid ei in via contigerit deducetis canos meos cum maerore ad inferos
GEN|44|30|igitur si intravero ad servum tuum patrem nostrum et puer defuerit cum anima illius ex huius anima pendeat
GEN|44|31|videritque eum non esse nobiscum morietur et deducent famuli tui canos eius cum dolore ad inferos
GEN|44|32|ego proprie servus tuus qui in meam hunc recepi fidem et spopondi dicens nisi reduxero eum peccati reus ero in patrem meum omni tempore
GEN|44|33|manebo itaque servus tuus pro puero in ministerium domini mei et puer ascendat cum fratribus suis
GEN|44|34|non enim possum redire ad patrem absente puero ne calamitatis quae oppressura est patrem meum testis adsistam
GEN|45|1|non se poterat ultra cohibere Ioseph multis coram adstantibus unde praecepit ut egrederentur cuncti foras et nullus interesset alienus agnitioni mutuae
GEN|45|2|elevavitque vocem cum fletu quam audierunt Aegyptii omnisque domus Pharaonis
GEN|45|3|et dixit fratribus suis ego sum Ioseph adhuc pater meus vivit nec poterant respondere fratres nimio timore perterriti
GEN|45|4|ad quos ille clementer accedite inquit ad me et cum accessissent prope ego sum ait Ioseph frater vester quem vendidistis in Aegypto
GEN|45|5|nolite pavere nec vobis durum esse videatur quod vendidistis me in his regionibus pro salute enim vestra misit me Deus ante vos in Aegyptum
GEN|45|6|biennium est quod fames esse coepit in terra et adhuc quinque anni restant quibus nec arari poterit nec meti
GEN|45|7|praemisitque me Deus ut reservemini super terram et escas ad vivendum habere possitis
GEN|45|8|non vestro consilio sed Dei huc voluntate missus sum qui fecit me quasi patrem Pharaonis et dominum universae domus eius ac principem in omni terra Aegypti
GEN|45|9|festinate et ascendite ad patrem meum et dicetis ei haec mandat filius tuus Ioseph Deus me fecit dominum universae terrae Aegypti descende ad me ne moreris
GEN|45|10|et habita in terra Gessen erisque iuxta me tu et filii tui et filii filiorum tuorum oves tuae et armenta tua et universa quae possides
GEN|45|11|ibique te pascam adhuc enim quinque anni residui sunt famis ne et tu pereas et domus tua et omnia quae possides
GEN|45|12|en oculi vestri et oculi fratris mei Beniamin vident quod os meum loquatur ad vos
GEN|45|13|nuntiate patri meo universam gloriam meam et cuncta quae vidistis in Aegypto festinate et adducite eum ad me
GEN|45|14|cumque amplexatus recidisset in collum Beniamin fratris sui flevit illo quoque flente similiter super collum eius
GEN|45|15|osculatusque est Ioseph omnes fratres suos et ploravit super singulos post quae ausi sunt loqui ad eum
GEN|45|16|auditumque est et celebri sermone vulgatum in aula regis venerunt fratres Ioseph et gavisus est Pharao atque omnis familia eius
GEN|45|17|dixitque ad Ioseph ut imperaret fratribus suis dicens onerantes iumenta ite in terram Chanaan
GEN|45|18|et tollite inde patrem vestrum et cognationem et venite ad me et ego dabo vobis omnia bona Aegypti ut comedatis medullam terrae
GEN|45|19|praecipe etiam ut tollant plaustra de terra Aegypti ad subvectionem parvulorum suorum et coniugum ac dicito tollite patrem vestrum et properate quantocius venientes
GEN|45|20|ne dimittatis quicquam de supellectili vestra quia omnes opes Aegypti vestrae erunt
GEN|45|21|fecerunt filii Israhel ut eis mandatum fuerat quibus dedit Ioseph plaustra secundum Pharaonis imperium et cibaria in itinere
GEN|45|22|singulisque proferri iussit binas stolas Beniamin vero dedit trecentos argenteos cum quinque stolis optimis
GEN|45|23|tantundem pecuniae et vestium mittens patri suo addens eis asinos decem qui subveherent ex omnibus divitiis Aegypti et totidem asinas triticum in itinere panesque portantes
GEN|45|24|dimisit ergo fratres suos et proficiscentibus ait ne irascamini in via
GEN|45|25|qui ascendentes ex Aegypto venerunt in terram Chanaan ad patrem suum Iacob
GEN|45|26|et nuntiaverunt ei dicentes Ioseph vivit et ipse dominatur in omni terra Aegypti quo audito quasi de gravi somno evigilans tamen non credebat eis
GEN|45|27|illi contra referebant omnem ordinem rei cumque vidisset plaustra et universa quae miserat revixit spiritus eius
GEN|45|28|et ait sufficit mihi si adhuc Ioseph filius meus vivit vadam et videbo illum antequam moriar
GEN|46|1|profectusque Israhel cum omnibus quae habebat venit ad puteum Iuramenti et mactatis ibi victimis Deo patris sui Isaac
GEN|46|2|audivit eum per visionem nocte vocantem se et dicentem sibi Iacob Iacob cui respondit ecce adsum
GEN|46|3|ait illi Deus ego sum Fortissimus Deus patris tui noli timere et descende in Aegyptum quia in gentem magnam faciam te ibi
GEN|46|4|ego descendam tecum illuc et ego inde adducam te revertentem Ioseph quoque ponet manum suam super oculos tuos
GEN|46|5|surrexit Iacob a puteo Iuramenti tuleruntque eum filii cum parvulis et uxoribus suis in plaustris quae miserat Pharao ad portandum senem
GEN|46|6|et omnia quae possederat in terra Chanaan venitque in Aegyptum cum omni semine suo
GEN|46|7|filii eius et nepotes filiae et cuncta simul progenies
GEN|46|8|haec sunt autem nomina filiorum Israhel qui ingressi sunt in Aegyptum ipse cum liberis suis primogenitus Ruben
GEN|46|9|filii Ruben Enoch et Phallu et Esrom et Charmi
GEN|46|10|filii Symeon Iemuhel et Iamin et Ahod et Iachin et Saher et Saul filius Chananitidis
GEN|46|11|filii Levi Gerson Caath et Merari
GEN|46|12|filii Iuda Her et Onan et Sela et Phares et Zara mortui sunt autem Her et Onan in terra Chanaan natique sunt filii Phares Esrom et Amul
GEN|46|13|filii Isachar Thola et Phua et Iob et Semron
GEN|46|14|filii Zabulon Sared et Helon et Iahelel
GEN|46|15|hii filii Liae quos genuit in Mesopotamiam Syriae cum Dina filia sua omnes animae filiorum eius et filiarum triginta tres
GEN|46|16|filii Gad Sephion et Haggi Suni et Esebon Heri et Arodi et Areli
GEN|46|17|filii Aser Iamne et Iesua et Iesui et Beria Sara quoque soror eorum filii Beria Heber et Melchihel
GEN|46|18|hii filii Zelphae quam dedit Laban Liae filiae suae et hos genuit Iacob sedecim animas
GEN|46|19|filii Rahel uxoris Iacob Ioseph et Beniamin
GEN|46|20|natique sunt Ioseph filii in terra Aegypti quos genuit ei Aseneth filia Putiphare sacerdotis Heliopoleos Manasses et Ephraim
GEN|46|21|filii Beniamin Bela et Bechor et Asbel Gera et Naaman et Ehi et Ros Mophim et Opphim et Ared
GEN|46|22|hii filii Rahel quos genuit Iacob omnes animae quattuordecim
GEN|46|23|filii Dan Usim
GEN|46|24|filii Nepthalim Iasihel et Guni et Hieser et Sallem
GEN|46|25|hii filii Balae quam dedit Laban Raheli filiae suae et hos genuit Iacob omnes animae septem
GEN|46|26|cunctae animae quae ingressae sunt cum Iacob in Aegyptum et egressae de femore illius absque uxoribus filiorum sexaginta sex
GEN|46|27|filii autem Ioseph qui nati sunt ei in terra Aegypti animae duae omnis anima domus Iacob quae ingressa est Aegyptum fuere septuaginta
GEN|46|28|misit autem Iudam ante se ad Ioseph ut nuntiaret ei et ille occurreret in Gessen
GEN|46|29|quo cum pervenisset iuncto Ioseph curru suo ascendit obviam patri ad eundem locum vidensque eum inruit super collum eius et inter amplexus flevit
GEN|46|30|dixitque pater ad Ioseph iam laetus moriar quia vidi faciem tuam et superstitem te relinquo
GEN|46|31|et ille locutus est ad fratres et ad omnem domum patris sui ascendam et nuntiabo Pharaoni dicamque ei fratres mei et domus patris mei qui erant in terra Chanaan venerunt ad me
GEN|46|32|et sunt viri pastores ovium curamque habent alendorum gregum pecora sua et armenta et omnia quae habere potuerunt adduxerunt secum
GEN|46|33|cumque vocaverit vos et dixerit quod est opus vestrum
GEN|46|34|respondebitis viri pastores sumus servi tui ab infantia nostra usque in praesens et nos et patres nostri haec autem dicetis ut habitare possitis in terra Gessen quia detestantur Aegyptii omnes pastores ovium
GEN|47|1|ingressus ergo Ioseph nuntiavit Pharaoni dicens pater meus et fratres oves eorum et armenta et cuncta quae possident venerunt de terra Chanaan et ecce consistunt in terra Gessen
GEN|47|2|extremos quoque fratrum suorum quinque viros statuit coram rege
GEN|47|3|quos ille interrogavit quid habetis operis responderunt pastores ovium sumus servi tui et nos et patres nostri
GEN|47|4|ad peregrinandum in terra tua venimus quoniam non est herba gregibus servorum tuorum ingravescente fame in regione Chanaan petimusque ut esse nos iubeas servos tuos in terra Gessen
GEN|47|5|dixit itaque rex ad Ioseph pater tuus et fratres tui venerunt ad te
GEN|47|6|terra Aegypti in conspectu tuo est in optimo loco fac habitare eos et trade eis terram Gessen quod si nosti esse in eis viros industrios constitue illos magistros pecorum meorum
GEN|47|7|post haec introduxit Ioseph patrem suum ad regem et statuit eum coram eo qui benedicens illi
GEN|47|8|et interrogatus ab eo quot sunt dies annorum vitae tuae
GEN|47|9|respondit dies peregrinationis vitae meae centum triginta annorum sunt parvi et mali et non pervenerunt usque ad dies patrum meorum quibus peregrinati sunt
GEN|47|10|et benedicto rege egressus est foras
GEN|47|11|Ioseph vero patri et fratribus suis dedit possessionem in Aegypto in optimo loco terrae solo Ramesses ut praeceperat Pharao
GEN|47|12|et alebat eos omnemque domum patris sui praebens cibaria singulis
GEN|47|13|in toto enim orbe panis deerat et oppresserat fames terram maxime Aegypti et Chanaan
GEN|47|14|e quibus omnem pecuniam congregavit pro venditione frumenti et intulit eam in aerarium regis
GEN|47|15|cumque defecisset emptoris pretium venit cuncta Aegyptus ad Ioseph dicens da nobis panes quare morimur coram te deficiente pecunia
GEN|47|16|quibus ille respondit adducite pecora vestra et dabo vobis pro eis cibos si pretium non habetis
GEN|47|17|quae cum adduxissent dedit eis alimenta pro equis et ovibus et bubus et asinis sustentavitque eos illo anno pro commutatione pecorum
GEN|47|18|veneruntque anno secundo et dixerunt ei non celamus dominum nostrum quod deficiente pecunia pecora simul defecerint nec clam te est quod absque corporibus et terra nihil habeamus
GEN|47|19|cur ergo morimur te vidente et nos et terra nostra tui erimus eme nos in servitutem regiam et praebe semina ne pereunte cultore redigatur terra in solitudinem
GEN|47|20|emit igitur Ioseph omnem terram Aegypti vendentibus singulis possessiones suas prae magnitudine famis subiecitque eam Pharaoni
GEN|47|21|et cunctos populos eius a novissimis terminis Aegypti usque ad extremos fines eius
GEN|47|22|praeter terram sacerdotum quae a rege tradita fuerat eis quibus et statuta cibaria ex horreis publicis praebebantur et idcirco non sunt conpulsi vendere possessiones suas
GEN|47|23|dixit ergo Ioseph ad populos en ut cernitis et vos et terram vestram Pharao possidet accipite semina et serite agros
GEN|47|24|ut fruges habere possitis quintam partem regi dabitis quattuor reliquas permitto vobis in sementem et in cibos famulis et liberis vestris
GEN|47|25|qui responderunt salus nostra in manu tua est respiciat nos tantum dominus noster et laeti serviemus regi
GEN|47|26|ex eo tempore usque in praesentem diem in universa terra Aegypti regibus quinta pars solvitur et factum est quasi in legem absque terra sacerdotali quae libera ab hac condicione fuit
GEN|47|27|habitavit ergo Israhel in Aegypto id est in terra Gessen et possedit eam auctusque est et multiplicatus nimis
GEN|47|28|et vixit in ea decem et septem annis factique sunt omnes dies vitae illius centum quadraginta septem annorum
GEN|47|29|cumque adpropinquare cerneret mortis diem vocavit filium suum Ioseph et dixit ad eum si inveni gratiam in conspectu tuo pone manum sub femore meo et facies mihi misericordiam et veritatem ut non sepelias me in Aegypto
GEN|47|30|sed dormiam cum patribus meis et auferas me de hac terra condasque in sepulchro maiorum cui respondit Ioseph ego faciam quod iussisti
GEN|47|31|et ille iura ergo inquit mihi quo iurante adoravit Israhel Deum conversus ad lectuli caput
GEN|48|1|his ita transactis nuntiatum est Ioseph quod aegrotaret pater eius qui adsumptis duobus filiis Manasse et Ephraim ire perrexit
GEN|48|2|dictumque est seni ecce filius tuus Ioseph venit ad te qui confortatus sedit in lectulo
GEN|48|3|et ingresso ad se ait Deus omnipotens apparuit mihi in Luza quae est in terra Chanaan benedixitque mihi
GEN|48|4|et ait ego te augebo et multiplicabo et faciam in turbas populorum daboque tibi terram hanc et semini tuo post te in possessionem sempiternam
GEN|48|5|duo igitur filii tui qui nati sunt tibi in terra Aegypti antequam huc venirem ad te mei erunt Ephraim et Manasses sicut Ruben et Symeon reputabuntur mihi
GEN|48|6|reliquos autem quos genueris post eos tui erunt et nomine fratrum suorum vocabuntur in possessionibus suis
GEN|48|7|mihi enim quando veniebam de Mesopotamiam mortua est Rahel in terra Chanaan in ipso itinere eratque vernum tempus et ingrediebar Ephratam et sepelivi eam iuxta viam Ephratae quae alio nomine appellatur Bethleem
GEN|48|8|videns autem filios eius dixit ad eum qui sunt isti
GEN|48|9|respondit filii mei sunt quos dedit mihi Deus in hoc loco adduc inquit eos ad me ut benedicam illis
GEN|48|10|oculi enim Israhel caligabant prae nimia senectute et clare videre non poterat adplicitosque ad se deosculatus et circumplexus
GEN|48|11|dixit ad filium non sum fraudatus aspectu tuo insuper ostendit mihi Deus semen tuum
GEN|48|12|cumque tulisset eos Ioseph de gremio patris adoravit pronus in terram
GEN|48|13|et posuit Ephraim ad dexteram suam id est ad sinistram Israhel Manassen vero in sinistra sua ad dexteram scilicet patris adplicuitque ambos ad eum
GEN|48|14|qui extendens manum dextram posuit super caput Ephraim iunioris fratris sinistram autem super caput Manasse qui maior natu erat commutans manus
GEN|48|15|benedixitque Ioseph filio suo et ait Deus in cuius conspectu ambulaverunt patres mei Abraham et Isaac Deus qui pascit me ab adulescentia mea usque in praesentem diem
GEN|48|16|angelus qui eruit me de cunctis malis benedicat pueris et invocetur super eos nomen meum nomina quoque patrum meorum Abraham et Isaac et crescant in multitudinem super terram
GEN|48|17|videns autem Ioseph quod posuisset pater suus dexteram manum super caput Ephraim graviter accepit et adprehensam patris manum levare conatus est de capite Ephraim et transferre super caput Manasse
GEN|48|18|dixitque ad patrem non ita convenit pater quia hic est primogenitus pone dexteram tuam super caput eius
GEN|48|19|qui rennuens ait scio fili mi scio et iste quidem erit in populos et multiplicabitur sed frater eius iunior maior illo erit et semen illius crescet in gentes
GEN|48|20|benedixitque eis in ipso tempore dicens in te benedicetur Israhel atque dicetur faciat tibi Deus sicut Ephraim et sicut Manasse constituitque Ephraim ante Manassen
GEN|48|21|et ait ad Ioseph filium suum en ego morior et erit Deus vobiscum reducetque vos ad terram patrum vestrorum
GEN|48|22|do tibi partem unam extra fratres tuos quam tuli de manu Amorrei in gladio et arcu meo
GEN|49|1|vocavit autem Iacob filios suos et ait eis congregamini ut adnuntiem quae ventura sunt vobis diebus novissimis
GEN|49|2|congregamini et audite filii Iacob audite Israhel patrem vestrum
GEN|49|3|Ruben primogenitus meus tu fortitudo mea et principium doloris mei prior in donis maior imperio
GEN|49|4|effusus es sicut aqua non crescas quia ascendisti cubile patris tui et maculasti stratum eius
GEN|49|5|Symeon et Levi fratres vasa iniquitatis bellantia
GEN|49|6|in consilio eorum ne veniat anima mea et in coetu illorum non sit gloria mea quia in furore suo occiderunt virum et in voluntate sua suffoderunt murum
GEN|49|7|maledictus furor eorum quia pertinax et indignatio illorum quia dura dividam eos in Iacob et dispergam illos in Israhel
GEN|49|8|Iuda te laudabunt fratres tui manus tua in cervicibus inimicorum tuorum adorabunt te filii patris tui
GEN|49|9|catulus leonis Iuda a praeda fili mi ascendisti requiescens accubuisti ut leo et quasi leaena quis suscitabit eum
GEN|49|10|non auferetur sceptrum de Iuda et dux de femoribus eius donec veniat qui mittendus est et ipse erit expectatio gentium
GEN|49|11|ligans ad vineam pullum suum et ad vitem o fili mi asinam suam lavabit vino stolam suam et sanguine uvae pallium suum
GEN|49|12|pulchriores oculi eius vino et dentes lacte candidiores
GEN|49|13|Zabulon in litore maris habitabit et in statione navium pertingens usque ad Sidonem
GEN|49|14|Isachar asinus fortis accubans inter terminos
GEN|49|15|vidit requiem quod esset bona et terram quod optima et subposuit umerum suum ad portandum factusque est tributis serviens
GEN|49|16|Dan iudicabit populum suum sicut et alia tribus Israhel
GEN|49|17|fiat Dan coluber in via cerastes in semita mordens ungulas equi ut cadat ascensor eius retro
GEN|49|18|salutare tuum expectabo Domine
GEN|49|19|Gad accinctus proeliabitur ante eum et ipse accingetur retrorsum
GEN|49|20|Aser pinguis panis eius et praebebit delicias regibus
GEN|49|21|Nepthalim cervus emissus et dans eloquia pulchritudinis
GEN|49|22|filius adcrescens Ioseph filius adcrescens et decorus aspectu filiae discurrerunt super murum
GEN|49|23|sed exasperaverunt eum et iurgati sunt invideruntque illi habentes iacula
GEN|49|24|sedit in forti arcus eius et dissoluta sunt vincula brachiorum et manuum illius per manus potentis Iacob inde pastor egressus est lapis Israhel
GEN|49|25|Deus patris tui erit adiutor tuus et Omnipotens benedicet tibi benedictionibus caeli desuper benedictionibus abyssi iacentis deorsum benedictionibus uberum et vulvae
GEN|49|26|benedictiones patris tui confortatae sunt benedictionibus patrum eius donec veniret desiderium collium aeternorum fiant in capite Ioseph et in vertice nazarei inter fratres suos
GEN|49|27|Beniamin lupus rapax mane comedet praedam et vespere dividet spolia
GEN|49|28|omnes hii in tribubus Israhel duodecim haec locutus est eis pater suus benedixitque singulis benedictionibus propriis
GEN|49|29|et praecepit eis dicens ego congregor ad populum meum sepelite me cum patribus meis in spelunca duplici quae est in agro Ephron Hetthei
GEN|49|30|contra Mambre in terra Chanaan quam emit Abraham cum agro ab Ephron Hettheo in possessionem sepulchri
GEN|49|31|ibi sepelierunt eum et Sarram uxorem eius ibi sepultus est Isaac cum Rebecca coniuge ibi et Lia condita iacet
GEN|49|32|finitisque mandatis quibus filios instruebat collegit pedes suos super lectulum et obiit adpositusque est ad populum suum
GEN|49|33|
GEN|50|1|quod cernens Ioseph ruit super faciem patris flens et deosculans eum
GEN|50|2|praecepitque servis suis medicis ut aromatibus condirent patrem
GEN|50|3|quibus iussa explentibus transierunt quadraginta dies iste quippe mos erat cadaverum conditorum flevitque eum Aegyptus septuaginta diebus
GEN|50|4|et expleto planctus tempore locutus est Ioseph ad familiam Pharaonis si inveni gratiam in conspectu vestro loquimini in auribus Pharaonis
GEN|50|5|eo quod pater meus adiuraverit me dicens en morior in sepulchro meo quod fodi mihi in terra Chanaan sepelies me ascendam igitur et sepeliam patrem meum ac revertar
GEN|50|6|dixitque ei Pharao ascende et sepeli patrem tuum sicut adiuratus es
GEN|50|7|quo ascendente ierunt cum eo omnes senes domus Pharaonis cunctique maiores natu terrae Aegypti
GEN|50|8|domus Ioseph cum fratribus suis absque parvulis et gregibus atque armentis quae dereliquerant in terra Gessen
GEN|50|9|habuit quoque in comitatu currus et equites et facta est turba non modica
GEN|50|10|veneruntque ad aream Atad quae sita est trans Iordanem ubi celebrantes exequias planctu magno atque vehementi impleverunt septem dies
GEN|50|11|quod cum vidissent habitatores terrae Chanaan dixerunt planctus magnus est iste Aegyptiis et idcirco appellaverunt nomen loci illius Planctus Aegypti
GEN|50|12|fecerunt ergo filii Iacob sicut praeceperat eis
GEN|50|13|et portantes eum in terram Chanaan sepelierunt in spelunca duplici quam emerat Abraham cum agro in possessionem sepulchri ab Ephron Hettheo contra faciem Mambre
GEN|50|14|reversusque est Ioseph in Aegyptum cum fratribus suis et omni comitatu sepulto patre
GEN|50|15|quo mortuo timentes fratres eius et mutuo conloquentes ne forte memor sit iniuriae quam passus est et reddat nobis malum omne quod fecimus
GEN|50|16|mandaverunt ei pater tuus praecepit nobis antequam moreretur
GEN|50|17|ut haec tibi verbis illius diceremus obsecro ut obliviscaris sceleris fratrum tuorum et peccati atque malitiae quam exercuerunt in te nos quoque oramus ut servis Dei patris tui dimittas iniquitatem hanc quibus auditis flevit Ioseph
GEN|50|18|veneruntque ad eum fratres sui et proni in terram dixerunt servi tui sumus
GEN|50|19|quibus ille respondit nolite timere num Dei possumus rennuere voluntatem
GEN|50|20|vos cogitastis de me malum et Deus vertit illud in bonum ut exaltaret me sicut inpraesentiarum cernitis et salvos faceret multos populos
GEN|50|21|nolite metuere ego pascam vos et parvulos vestros consolatusque est eos et blande ac leniter est locutus
GEN|50|22|et habitavit in Aegypto cum omni domo patris sui vixitque centum decem annis et vidit Ephraim filios usque ad tertiam generationem filii quoque Machir filii Manasse nati sunt in genibus Ioseph
GEN|50|23|quibus transactis locutus est fratribus suis post mortem meam Deus visitabit vos et ascendere faciet de terra ista ad terram quam iuravit Abraham Isaac et Iacob
GEN|50|24|cumque adiurasset eos atque dixisset Deus visitabit vos asportate vobiscum ossa mea de loco isto
GEN|50|25|mortuus est expletis centum decem vitae suae annis et conditus aromatibus repositus est in loculo in Aegypto
GEN|50|26|
