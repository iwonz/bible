ROM|1|1|Павел, раб Иисуса Христа, призванный Апостол, избранный к благовестию Божию,
ROM|1|2|которое Бог прежде обещал через пророков Своих, в святых писаниях,
ROM|1|3|о Сыне Своем, Который родился от семени Давидова по плоти
ROM|1|4|и открылся Сыном Божиим в силе, по духу святыни, через воскресение из мертвых, о Иисусе Христе Господе нашем,
ROM|1|5|через Которого мы получили благодать и апостольство, чтобы во имя Его покорять вере все народы,
ROM|1|6|между которыми находитесь и вы, призванные Иисусом Христом, –
ROM|1|7|всем находящимся в Риме возлюбленным Божиим, призванным святым: благодать вам и мир от Бога отца нашего и Господа Иисуса Христа.
ROM|1|8|Прежде всего благодарю Бога моего через Иисуса Христа за всех вас, что вера ваша возвещается во всем мире.
ROM|1|9|Свидетель мне Бог, Которому служу духом моим в благовествовании Сына Его, что непрестанно воспоминаю о вас,
ROM|1|10|всегда прося в молитвах моих, чтобы воля Божия когда–нибудь благопоспешила мне придти к вам,
ROM|1|11|ибо я весьма желаю увидеть вас, чтобы преподать вам некое дарование духовное к утверждению вашему,
ROM|1|12|то есть утешиться с вами верою общею, вашею и моею.
ROM|1|13|Не хочу, братия, [оставить] вас в неведении, что я многократно намеревался придти к вам (но встречал препятствия даже доныне), чтобы иметь некий плод и у вас, как и у прочих народов.
ROM|1|14|Я должен и Еллинам и варварам, мудрецам и невеждам.
ROM|1|15|Итак, что до меня, я готов благовествовать и вам, находящимся в Риме.
ROM|1|16|Ибо я не стыжусь благовествования Христова, потому что [оно] есть сила Божия ко спасению всякому верующему, во–первых, Иудею, [потом] и Еллину.
ROM|1|17|В нем открывается правда Божия от веры в веру, как написано: праведный верою жив будет.
ROM|1|18|Ибо открывается гнев Божий с неба на всякое нечестие и неправду человеков, подавляющих истину неправдою.
ROM|1|19|Ибо, что можно знать о Боге, явно для них, потому что Бог явил им.
ROM|1|20|Ибо невидимое Его, вечная сила Его и Божество, от создания мира через рассматривание творений видимы, так что они безответны.
ROM|1|21|Но как они, познав Бога, не прославили Его, как Бога, и не возблагодарили, но осуетились в умствованиях своих, и омрачилось несмысленное их сердце;
ROM|1|22|называя себя мудрыми, обезумели,
ROM|1|23|и славу нетленного Бога изменили в образ, подобный тленному человеку, и птицам, и четвероногим, и пресмыкающимся, –
ROM|1|24|то и предал их Бог в похотях сердец их нечистоте, так что они сквернили сами свои тела.
ROM|1|25|Они заменили истину Божию ложью, и поклонялись, и служили твари вместо Творца, Который благословен во веки, аминь.
ROM|1|26|Потому предал их Бог постыдным страстям: женщины их заменили естественное употребление противоестественным;
ROM|1|27|подобно и мужчины, оставив естественное употребление женского пола, разжигались похотью друг на друга, мужчины на мужчинах делая срам и получая в самих себе должное возмездие за свое заблуждение.
ROM|1|28|И как они не заботились иметь Бога в разуме, то предал их Бог превратному уму – делать непотребства,
ROM|1|29|так что они исполнены всякой неправды, блуда, лукавства, корыстолюбия, злобы, исполнены зависти, убийства, распрей, обмана, злонравия,
ROM|1|30|злоречивы, клеветники, богоненавистники, обидчики, самохвалы, горды, изобретательны на зло, непослушны родителям,
ROM|1|31|безрассудны, вероломны, нелюбовны, непримиримы, немилостивы.
ROM|1|32|Они знают праведный [суд] Божий, что делающие такие [дела] достойны смерти; однако не только [их] делают, но и делающих одобряют.
ROM|2|1|Итак, неизвинителен ты, всякий человек, судящий [другого], ибо тем же судом, каким судишь другого, осуждаешь себя, потому что, судя [другого], делаешь то же.
ROM|2|2|А мы знаем, что поистине есть суд Божий на делающих такие [дела].
ROM|2|3|Неужели думаешь ты, человек, что избежишь суда Божия, осуждая делающих такие [дела] и (сам) делая то же?
ROM|2|4|Или пренебрегаешь богатство благости, кротости и долготерпения Божия, не разумея, что благость Божия ведет тебя к покаянию?
ROM|2|5|Но, по упорству твоему и нераскаянному сердцу, ты сам себе собираешь гнев на день гнева и откровения праведного суда от Бога,
ROM|2|6|Который воздаст каждому по делам его:
ROM|2|7|тем, которые постоянством в добром деле ищут славы, чести и бессмертия, – жизнь вечную;
ROM|2|8|а тем, которые упорствуют и не покоряются истине, но предаются неправде, – ярость и гнев.
ROM|2|9|Скорбь и теснота всякой душе человека, делающего злое, во–первых, Иудея, [потом] и Еллина!
ROM|2|10|Напротив, слава и честь и мир всякому, делающему доброе, во–первых, Иудею, [потом] и Еллину!
ROM|2|11|Ибо нет лицеприятия у Бога.
ROM|2|12|Те, которые, не [имея] закона, согрешили, вне закона и погибнут; а те, которые под законом согрешили, по закону осудятся
ROM|2|13|(потому что не слушатели закона праведны пред Богом, но исполнители закона оправданы будут,
ROM|2|14|ибо когда язычники, не имеющие закона, по природе законное делают, то, не имея закона, они сами себе закон:
ROM|2|15|они показывают, что дело закона у них написано в сердцах, о чем свидетельствует совесть их и мысли их, то обвиняющие, то оправдывающие одна другую)
ROM|2|16|в день, когда, по благовествованию моему, Бог будет судить тайные [дела] человеков через Иисуса Христа.
ROM|2|17|Вот, ты называешься Иудеем, и успокаиваешь себя законом, и хвалишься Богом,
ROM|2|18|и знаешь волю [Его], и разумеешь лучшее, научаясь из закона,
ROM|2|19|и уверен о себе, что ты путеводитель слепых, свет для находящихся во тьме,
ROM|2|20|наставник невежд, учитель младенцев, имеющий в законе образец ведения и истины:
ROM|2|21|как же ты, уча другого, не учишь себя самого?
ROM|2|22|Проповедуя не красть, крадешь? говоря: "не прелюбодействуй", прелюбодействуешь? гнушаясь идолов, святотатствуешь?
ROM|2|23|Хвалишься законом, а преступлением закона бесчестишь Бога?
ROM|2|24|Ибо ради вас, как написано, имя Божие хулится у язычников.
ROM|2|25|Обрезание полезно, если исполняешь закон; а если ты преступник закона, то обрезание твое стало необрезанием.
ROM|2|26|Итак, если необрезанный соблюдает постановления закона, то его необрезание не вменится ли ему в обрезание?
ROM|2|27|И необрезанный по природе, исполняющий закон, не осудит ли тебя, преступника закона при Писании и обрезании?
ROM|2|28|Ибо не тот Иудей, кто [таков] по наружности, и не то обрезание, которое наружно, на плоти;
ROM|2|29|но [тот] Иудей, кто внутренно [таков], и [то] обрезание, [которое] в сердце, по духу, [а] не по букве: ему и похвала не от людей, но от Бога.
ROM|3|1|Итак, какое преимущество [быть] Иудеем, или какая польза от обрезания?
ROM|3|2|Великое преимущество во всех отношениях, а наипаче [в том], что им вверено слово Божие.
ROM|3|3|Ибо что же? если некоторые и неверны были, неверность их уничтожит ли верность Божию?
ROM|3|4|Никак. Бог верен, а всякий человек лжив, как написано: Ты праведен в словах Твоих и победишь в суде Твоем.
ROM|3|5|Если же наша неправда открывает правду Божию, то что скажем? не будет ли Бог несправедлив, когда изъявляет гнев? (говорю по человеческому [рассуждению]).
ROM|3|6|Никак. Ибо [иначе] как Богу судить мир?
ROM|3|7|Ибо, если верность Божия возвышается моею неверностью к славе Божией, за что еще меня же судить, как грешника?
ROM|3|8|И не делать ли нам зло, чтобы вышло добро, как некоторые злословят нас и говорят, будто мы так учим? Праведен суд на таковых.
ROM|3|9|Итак, что же? имеем ли мы преимущество? Нисколько. Ибо мы уже доказали, что как Иудеи, так и Еллины, все под грехом,
ROM|3|10|как написано: нет праведного ни одного;
ROM|3|11|нет разумевающего; никто не ищет Бога;
ROM|3|12|все совратились с пути, до одного негодны; нет делающего добро, нет ни одного.
ROM|3|13|Гортань их – открытый гроб; языком своим обманывают; яд аспидов на губах их.
ROM|3|14|Уста их полны злословия и горечи.
ROM|3|15|Ноги их быстры на пролитие крови;
ROM|3|16|разрушение и пагуба на путях их;
ROM|3|17|они не знают пути мира.
ROM|3|18|Нет страха Божия перед глазами их.
ROM|3|19|Но мы знаем, что закон, если что говорит, говорит к состоящим под законом, так что заграждаются всякие уста, и весь мир становится виновен пред Богом,
ROM|3|20|потому что делами закона не оправдается пред Ним никакая плоть; ибо законом познается грех.
ROM|3|21|Но ныне, независимо от закона, явилась правда Божия, о которой свидетельствуют закон и пророки,
ROM|3|22|правда Божия через веру в Иисуса Христа во всех и на всех верующих, ибо нет различия,
ROM|3|23|потому что все согрешили и лишены славы Божией,
ROM|3|24|получая оправдание даром, по благодати Его, искуплением во Христе Иисусе,
ROM|3|25|которого Бог предложил в жертву умилостивления в Крови Его через веру, для показания правды Его в прощении грехов, соделанных прежде,
ROM|3|26|во [время] долготерпения Божия, к показанию правды Его в настоящее время, да [явится] Он праведным и оправдывающим верующего в Иисуса.
ROM|3|27|Где же то, чем бы хвалиться? уничтожено. Каким законом? [законом] дел? Нет, но законом веры.
ROM|3|28|Ибо мы признаем, что человек оправдывается верою, независимо от дел закона.
ROM|3|29|Неужели Бог [есть Бог] Иудеев только, а не и язычников? Конечно, и язычников,
ROM|3|30|потому что один Бог, Который оправдает обрезанных по вере и необрезанных через веру.
ROM|3|31|Итак, мы уничтожаем закон верою? Никак; но закон утверждаем.
ROM|4|1|Что же, скажем, Авраам, отец наш, приобрел по плоти?
ROM|4|2|Если Авраам оправдался делами, он имеет похвалу, но не пред Богом.
ROM|4|3|Ибо что говорит Писание? Поверил Авраам Богу, и это вменилось ему в праведность.
ROM|4|4|Воздаяние делающему вменяется не по милости, но по долгу.
ROM|4|5|А не делающему, но верующему в Того, Кто оправдывает нечестивого, вера его вменяется в праведность.
ROM|4|6|Так и Давид называет блаженным человека, которому Бог вменяет праведность независимо от дел:
ROM|4|7|Блаженны, чьи беззакония прощены и чьи грехи покрыты.
ROM|4|8|Блажен человек, которому Господь не вменит греха.
ROM|4|9|Блаженство сие [относится] к обрезанию, или к необрезанию? Мы говорим, что Аврааму вера вменилась в праведность.
ROM|4|10|Когда вменилась? по обрезании или до обрезания? Не по обрезании, а до обрезания.
ROM|4|11|И знак обрезания он получил, [как] печать праведности через веру, которую [имел] в необрезании, так что он стал отцом всех верующих в необрезании, чтобы и им вменилась праведность,
ROM|4|12|и отцом обрезанных, не только [принявших] обрезание, но и ходящих по следам веры отца нашего Авраама, которую [имел он] в необрезании.
ROM|4|13|Ибо не законом [даровано] Аврааму, или семени его, обетование – быть наследником мира, но праведностью веры.
ROM|4|14|Если утверждающиеся на законе суть наследники, то тщетна вера, бездейственно обетование;
ROM|4|15|ибо закон производит гнев, потому что, где нет закона, нет и преступления.
ROM|4|16|Итак по вере, чтобы [было] по милости, дабы обетование было непреложно для всех, не только по закону, но и по вере потомков Авраама, который есть отец всем нам
ROM|4|17|(как написано: Я поставил тебя отцом многих народов) пред Богом, Которому он поверил, животворящим мертвых и называющим несуществующее, как существующее.
ROM|4|18|Он, сверх надежды, поверил с надеждою, через что сделался отцом многих народов, по сказанному: "так [многочисленно] будет семя твое".
ROM|4|19|И, не изнемогши в вере, он не помышлял, что тело его, почти столетнего, уже омертвело, и утроба Саррина в омертвении;
ROM|4|20|не поколебался в обетовании Божием неверием, но пребыл тверд в вере, воздав славу Богу
ROM|4|21|и будучи вполне уверен, что Он силен и исполнить обещанное.
ROM|4|22|Потому и вменилось ему в праведность.
ROM|4|23|А впрочем не в отношении к нему одному написано, что вменилось ему,
ROM|4|24|но и в отношении к нам; вменится и нам, верующим в Того, Кто воскресил из мертвых Иисуса Христа, Господа нашего,
ROM|4|25|Который предан за грехи наши и воскрес для оправдания нашего.
ROM|5|1|Итак, оправдавшись верою, мы имеем мир с Богом через Господа нашего Иисуса Христа,
ROM|5|2|через Которого верою и получили мы доступ к той благодати, в которой стоим и хвалимся надеждою славы Божией.
ROM|5|3|И не сим только, но хвалимся и скорбями, зная, что от скорби происходит терпение,
ROM|5|4|от терпения опытность, от опытности надежда,
ROM|5|5|а надежда не постыжает, потому что любовь Божия излилась в сердца наши Духом Святым, данным нам.
ROM|5|6|Ибо Христос, когда еще мы были немощны, в определенное время умер за нечестивых.
ROM|5|7|Ибо едва ли кто умрет за праведника; разве за благодетеля, может быть, кто и решится умереть.
ROM|5|8|Но Бог Свою любовь к нам доказывает тем, что Христос умер за нас, когда мы были еще грешниками.
ROM|5|9|Посему тем более ныне, будучи оправданы Кровию Его, спасемся Им от гнева.
ROM|5|10|Ибо если, будучи врагами, мы примирились с Богом смертью Сына Его, то тем более, примирившись, спасемся жизнью Его.
ROM|5|11|И не довольно сего, но и хвалимся Богом чрез Господа нашего Иисуса Христа, посредством Которого мы получили ныне примирение.
ROM|5|12|Посему, как одним человеком грех вошел в мир, и грехом смерть, так и смерть перешла во всех человеков, [потому что] в нем все согрешили.
ROM|5|13|Ибо [и] до закона грех был в мире; но грех не вменяется, когда нет закона.
ROM|5|14|Однако же смерть царствовала от Адама до Моисея и над несогрешившими подобно преступлению Адама, который есть образ будущего.
ROM|5|15|Но дар благодати не как преступление. Ибо если преступлением одного подверглись смерти многие, то тем более благодать Божия и дар по благодати одного Человека, Иисуса Христа, преизбыточествуют для многих.
ROM|5|16|И дар не как [суд] за одного согрешившего; ибо суд за одно [преступление] – к осуждению; а дар благодати – к оправданию от многих преступлений.
ROM|5|17|Ибо если преступлением одного смерть царствовала посредством одного, то тем более приемлющие обилие благодати и дар праведности будут царствовать в жизни посредством единого Иисуса Христа.
ROM|5|18|Посему, как преступлением одного всем человекам осуждение, так правдою одного всем человекам оправдание к жизни.
ROM|5|19|Ибо, как непослушанием одного человека сделались многие грешными, так и послушанием одного сделаются праведными многие.
ROM|5|20|Закон же пришел после, и таким образом умножилось преступление. А когда умножился грех, стала преизобиловать благодать,
ROM|5|21|дабы, как грех царствовал к смерти, так и благодать воцарилась через праведность к жизни вечной Иисусом Христом, Господом нашим.
ROM|6|1|Что же скажем? оставаться ли нам в грехе, чтобы умножилась благодать? Никак.
ROM|6|2|Мы умерли для греха: как же нам жить в нем?
ROM|6|3|Неужели не знаете, что все мы, крестившиеся во Христа Иисуса, в смерть Его крестились?
ROM|6|4|Итак мы погреблись с Ним крещением в смерть, дабы, как Христос воскрес из мертвых славою Отца, так и нам ходить в обновленной жизни.
ROM|6|5|Ибо если мы соединены с Ним подобием смерти Его, то должны быть [соединены] и [подобием] воскресения,
ROM|6|6|зная то, что ветхий наш человек распят с Ним, чтобы упразднено было тело греховное, дабы нам не быть уже рабами греху;
ROM|6|7|ибо умерший освободился от греха.
ROM|6|8|Если же мы умерли со Христом, то веруем, что и жить будем с Ним,
ROM|6|9|зная, что Христос, воскреснув из мертвых, уже не умирает: смерть уже не имеет над Ним власти.
ROM|6|10|Ибо, что Он умер, то умер однажды для греха; а что живет, то живет для Бога.
ROM|6|11|Так и вы почитайте себя мертвыми для греха, живыми же для Бога во Христе Иисусе, Господе нашем.
ROM|6|12|Итак да не царствует грех в смертном вашем теле, чтобы вам повиноваться ему в похотях его;
ROM|6|13|и не предавайте членов ваших греху в орудия неправды, но представьте себя Богу, как оживших из мертвых, и члены ваши Богу в орудия праведности.
ROM|6|14|Грех не должен над вами господствовать, ибо вы не под законом, но под благодатью.
ROM|6|15|Что же? станем ли грешить, потому что мы не под законом, а под благодатью? Никак.
ROM|6|16|Неужели вы не знаете, что, кому вы отдаете себя в рабы для послушания, того вы и рабы, кому повинуетесь, или [рабы] греха к смерти, или послушания к праведности?
ROM|6|17|Благодарение Богу, что вы, быв прежде рабами греха, от сердца стали послушны тому образу учения, которому предали себя.
ROM|6|18|Освободившись же от греха, вы стали рабами праведности.
ROM|6|19|Говорю по [рассуждению] человеческому, ради немощи плоти вашей. Как предавали вы члены ваши в рабы нечистоте и беззаконию на [дела] беззаконные, так ныне представьте члены ваши в рабы праведности на [дела] святые.
ROM|6|20|Ибо, когда вы были рабами греха, тогда были свободны от праведности.
ROM|6|21|Какой же плод вы имели тогда? [Такие дела], каких ныне сами стыдитесь, потому что конец их – смерть.
ROM|6|22|Но ныне, когда вы освободились от греха и стали рабами Богу, плод ваш есть святость, а конец – жизнь вечная.
ROM|6|23|Ибо возмездие за грех – смерть, а дар Божий – жизнь вечная во Христе Иисусе, Господе нашем.
ROM|7|1|Разве вы не знаете, братия (ибо говорю знающим закон), что закон имеет власть над человеком, пока он жив?
ROM|7|2|Замужняя женщина привязана законом к живому мужу; а если умрет муж, она освобождается от закона замужества.
ROM|7|3|Посему, если при живом муже выйдет за другого, называется прелюбодейцею; если же умрет муж, она свободна от закона, и не будет прелюбодейцею, выйдя за другого мужа.
ROM|7|4|Так и вы, братия мои, умерли для закона телом Христовым, чтобы принадлежать другому, Воскресшему из мертвых, да приносим плод Богу.
ROM|7|5|Ибо, когда мы жили по плоти, тогда страсти греховные, [обнаруживаемые] законом, действовали в членах наших, чтобы приносить плод смерти;
ROM|7|6|но ныне, умерши для закона, которым были связаны, мы освободились от него, чтобы нам служить Богу в обновлении духа, а не по ветхой букве.
ROM|7|7|Что же скажем? Неужели [от] закона грех? Никак. Но я не иначе узнал грех, как посредством закона. Ибо я не понимал бы и пожелания, если бы закон не говорил: не пожелай.
ROM|7|8|Но грех, взяв повод от заповеди, произвел во мне всякое пожелание: ибо без закона грех мертв.
ROM|7|9|Я жил некогда без закона; но когда пришла заповедь, то грех ожил,
ROM|7|10|а я умер; и таким образом заповедь, [данная] для жизни, послужила мне к смерти,
ROM|7|11|потому что грех, взяв повод от заповеди, обольстил меня и умертвил ею.
ROM|7|12|Посему закон свят, и заповедь свята и праведна и добра.
ROM|7|13|Итак, неужели доброе сделалось мне смертоносным? Никак; но грех, оказывающийся грехом потому, что посредством доброго причиняет мне смерть, так что грех становится крайне грешен посредством заповеди.
ROM|7|14|Ибо мы знаем, что закон духовен, а я плотян, продан греху.
ROM|7|15|Ибо не понимаю, что делаю: потому что не то делаю, что хочу, а что ненавижу, то делаю.
ROM|7|16|Если же делаю то, чего не хочу, то соглашаюсь с законом, что он добр,
ROM|7|17|а потому уже не я делаю то, но живущий во мне грех.
ROM|7|18|Ибо знаю, что не живет во мне, то есть в плоти моей, доброе; потому что желание добра есть во мне, но чтобы сделать оное, того не нахожу.
ROM|7|19|Доброго, которого хочу, не делаю, а злое, которого не хочу, делаю.
ROM|7|20|Если же делаю то, чего не хочу, уже не я делаю то, но живущий во мне грех.
ROM|7|21|Итак я нахожу закон, что, когда хочу делать доброе, прилежит мне злое.
ROM|7|22|Ибо по внутреннему человеку нахожу удовольствие в законе Божием;
ROM|7|23|но в членах моих вижу иной закон, противоборствующий закону ума моего и делающий меня пленником закона греховного, находящегося в членах моих.
ROM|7|24|Бедный я человек! кто избавит меня от сего тела смерти?
ROM|7|25|Благодарю Бога моего Иисусом Христом, Господом нашим. Итак тот же самый я умом моим служу закону Божию, а плотию закону греха.
ROM|8|1|Итак нет ныне никакого осуждения тем, которые во Христе Иисусе живут не по плоти, но по духу,
ROM|8|2|потому что закон духа жизни во Христе Иисусе освободил меня от закона греха и смерти.
ROM|8|3|Как закон, ослабленный плотию, был бессилен, то Бог послал Сына Своего в подобии плоти греховной [в жертву] за грех и осудил грех во плоти,
ROM|8|4|чтобы оправдание закона исполнилось в нас, живущих не по плоти, но по духу.
ROM|8|5|Ибо живущие по плоти о плотском помышляют, а живущие по духу – о духовном.
ROM|8|6|Помышления плотские суть смерть, а помышления духовные – жизнь и мир,
ROM|8|7|потому что плотские помышления суть вражда против Бога; ибо закону Божию не покоряются, да и не могут.
ROM|8|8|Посему живущие по плоти Богу угодить не могут.
ROM|8|9|Но вы не по плоти живете, а по духу, если только Дух Божий живет в вас. Если же кто Духа Христова не имеет, тот [и] не Его.
ROM|8|10|А если Христос в вас, то тело мертво для греха, но дух жив для праведности.
ROM|8|11|Если же Дух Того, Кто воскресил из мертвых Иисуса, живет в вас, то Воскресивший Христа из мертвых оживит и ваши смертные тела Духом Своим, живущим в вас.
ROM|8|12|Итак, братия, мы не должники плоти, чтобы жить по плоти;
ROM|8|13|ибо если живете по плоти, то умрете, а если духом умерщвляете дела плотские, то живы будете.
ROM|8|14|Ибо все, водимые Духом Божиим, суть сыны Божии.
ROM|8|15|Потому что вы не приняли духа рабства, [чтобы] опять [жить] в страхе, но приняли Духа усыновления, Которым взываем: "Авва, Отче!"
ROM|8|16|Сей самый Дух свидетельствует духу нашему, что мы – дети Божии.
ROM|8|17|А если дети, то и наследники, наследники Божии, сонаследники же Христу, если только с Ним страдаем, чтобы с Ним и прославиться.
ROM|8|18|Ибо думаю, что нынешние временные страдания ничего не стоят в сравнении с тою славою, которая откроется в нас.
ROM|8|19|Ибо тварь с надеждою ожидает откровения сынов Божиих,
ROM|8|20|потому что тварь покорилась суете не добровольно, но по воле покорившего ее, в надежде,
ROM|8|21|что и сама тварь освобождена будет от рабства тлению в свободу славы детей Божиих.
ROM|8|22|Ибо знаем, что вся тварь совокупно стенает и мучится доныне;
ROM|8|23|и не только [она], но и мы сами, имея начаток Духа, и мы в себе стенаем, ожидая усыновления, искупления тела нашего.
ROM|8|24|Ибо мы спасены в надежде. Надежда же, когда видит, не есть надежда; ибо если кто видит, то чего ему и надеяться?
ROM|8|25|Но когда надеемся того, чего не видим, тогда ожидаем в терпении.
ROM|8|26|Также и Дух подкрепляет нас в немощах наших; ибо мы не знаем, о чем молиться, как должно, но Сам Дух ходатайствует за нас воздыханиями неизреченными.
ROM|8|27|Испытующий же сердца знает, какая мысль у Духа, потому что Он ходатайствует за святых по [воле] Божией.
ROM|8|28|Притом знаем, что любящим Бога, призванным по [Его] изволению, все содействует ко благу.
ROM|8|29|Ибо кого Он предузнал, тем и предопределил быть подобными образу Сына Своего, дабы Он был первородным между многими братиями.
ROM|8|30|А кого Он предопределил, тех и призвал, а кого призвал, тех и оправдал; а кого оправдал, тех и прославил.
ROM|8|31|Что же сказать на это? Если Бог за нас, кто против нас?
ROM|8|32|Тот, Который Сына Своего не пощадил, но предал Его за всех нас, как с Ним не дарует нам и всего?
ROM|8|33|Кто будет обвинять избранных Божиих? Бог оправдывает [их].
ROM|8|34|Кто осуждает? Христос Иисус умер, но и воскрес: Он и одесную Бога, Он и ходатайствует за нас.
ROM|8|35|Кто отлучит нас от любви Божией: скорбь, или теснота, или гонение, или голод, или нагота, или опасность, или меч? как написано:
ROM|8|36|за Тебя умерщвляют нас всякий день, считают нас за овец, [обреченных] на заклание.
ROM|8|37|Но все сие преодолеваем силою Возлюбившего нас.
ROM|8|38|Ибо я уверен, что ни смерть, ни жизнь, ни Ангелы, ни Начала, ни Силы, ни настоящее, ни будущее,
ROM|8|39|ни высота, ни глубина, ни другая какая тварь не может отлучить нас от любви Божией во Христе Иисусе, Господе нашем.
ROM|9|1|Истину говорю во Христе, не лгу, свидетельствует мне совесть моя в Духе Святом,
ROM|9|2|что великая для меня печаль и непрестанное мучение сердцу моему:
ROM|9|3|я желал бы сам быть отлученным от Христа за братьев моих, родных мне по плоти,
ROM|9|4|то есть Израильтян, которым принадлежат усыновление и слава, и заветы, и законоположение, и богослужение, и обетования;
ROM|9|5|их и отцы, и от них Христос по плоти, сущий над всем Бог, благословенный во веки, аминь.
ROM|9|6|Но не то, чтобы слово Божие не сбылось: ибо не все те Израильтяне, которые от Израиля;
ROM|9|7|и не все дети Авраама, которые от семени его, но сказано: в Исааке наречется тебе семя.
ROM|9|8|То есть не плотские дети суть дети Божии, но дети обетования признаются за семя.
ROM|9|9|А слово обетования таково: в это же время приду, и у Сарры будет сын.
ROM|9|10|И не одно это; но [так было] и с Ревеккою, когда она зачала в одно время [двух сыновей] от Исаака, отца нашего.
ROM|9|11|Ибо, когда они еще не родились и не сделали ничего доброго или худого (дабы изволение Божие в избрании происходило
ROM|9|12|не от дел, но от Призывающего), сказано было ей: больший будет в порабощении у меньшего,
ROM|9|13|как и написано: Иакова Я возлюбил, а Исава возненавидел.
ROM|9|14|Что же скажем? Неужели неправда у Бога? Никак.
ROM|9|15|Ибо Он говорит Моисею: кого миловать, помилую; кого жалеть, пожалею.
ROM|9|16|Итак [помилование зависит] не от желающего и не от подвизающегося, но от Бога милующего.
ROM|9|17|Ибо Писание говорит фараону: для того самого Я и поставил тебя, чтобы показать над тобою силу Мою и чтобы проповедано было имя Мое по всей земле.
ROM|9|18|Итак, кого хочет, милует; а кого хочет, ожесточает.
ROM|9|19|Ты скажешь мне: "за что же еще обвиняет? Ибо кто противостанет воле Его?"
ROM|9|20|А ты кто, человек, что споришь с Богом? Изделие скажет ли сделавшему его: "зачем ты меня так сделал?"
ROM|9|21|Не властен ли горшечник над глиною, чтобы из той же смеси сделать один сосуд для почетного [употребления], а другой для низкого?
ROM|9|22|Что же, если Бог, желая показать гнев и явить могущество Свое, с великим долготерпением щадил сосуды гнева, готовые к погибели,
ROM|9|23|дабы вместе явить богатство славы Своей над сосудами милосердия, которые Он приготовил к славе,
ROM|9|24|над нами, которых Он призвал не только из Иудеев, но и из язычников?
ROM|9|25|Как и у Осии говорит: не Мой народ назову Моим народом, и не возлюбленную – возлюбленною.
ROM|9|26|И на том месте, где сказано им: вы не Мой народ, там названы будут сынами Бога живаго.
ROM|9|27|А Исаия провозглашает об Израиле: хотя бы сыны Израилевы были числом, как песок морской, [только] остаток спасется;
ROM|9|28|ибо дело оканчивает и скоро решит по правде, дело решительное совершит Господь на земле.
ROM|9|29|И, как предсказал Исаия: если бы Господь Саваоф не оставил нам семени, то мы сделались бы, как Содом, и были бы подобны Гоморре.
ROM|9|30|Что же скажем? Язычники, не искавшие праведности, получили праведность, праведность от веры.
ROM|9|31|А Израиль, искавший закона праведности, не достиг до закона праведности.
ROM|9|32|Почему? потому что [искали] не в вере, а в делах закона. Ибо преткнулись о камень преткновения,
ROM|9|33|как написано: вот, полагаю в Сионе камень преткновения и камень соблазна; но всякий, верующий в Него, не постыдится.
ROM|10|1|Братия! желание моего сердца и молитва к Богу об Израиле во спасение.
ROM|10|2|Ибо свидетельствую им, что имеют ревность по Боге, но не по рассуждению.
ROM|10|3|Ибо, не разумея праведности Божией и усиливаясь поставить собственную праведность, они не покорились праведности Божией,
ROM|10|4|потому что конец закона – Христос, к праведности всякого верующего.
ROM|10|5|Моисей пишет о праведности от закона: исполнивший его человек жив будет им.
ROM|10|6|А праведность от веры так говорит: не говори в сердце твоем: кто взойдет на небо? то есть Христа свести.
ROM|10|7|Или кто сойдет в бездну? то есть Христа из мертвых возвести.
ROM|10|8|Но что говорит Писание? Близко к тебе слово, в устах твоих и в сердце твоем, то есть слово веры, которое проповедуем.
ROM|10|9|Ибо если устами твоими будешь исповедывать Иисуса Господом и сердцем твоим веровать, что Бог воскресил Его из мертвых, то спасешься,
ROM|10|10|потому что сердцем веруют к праведности, а устами исповедуют ко спасению.
ROM|10|11|Ибо Писание говорит: всякий, верующий в Него, не постыдится.
ROM|10|12|Здесь нет различия между Иудеем и Еллином, потому что один Господь у всех, богатый для всех, призывающих Его.
ROM|10|13|Ибо всякий, кто призовет имя Господне, спасется.
ROM|10|14|Но как призывать [Того], в Кого не уверовали? как веровать [в] [Того], о Ком не слыхали? как слышать без проповедующего?
ROM|10|15|И как проповедывать, если не будут посланы? как написано: как прекрасны ноги благовествующих мир, благовествующих благое!
ROM|10|16|Но не все послушались благовествования. Ибо Исаия говорит: Господи! кто поверил слышанному от нас?
ROM|10|17|Итак вера от слышания, а слышание от слова Божия.
ROM|10|18|Но спрашиваю: разве они не слышали? Напротив, по всей земле прошел голос их, и до пределов вселенной слова их.
ROM|10|19|Еще спрашиваю: разве Израиль не знал? Но первый Моисей говорит: Я возбужу в вас ревность не народом, раздражу вас народом несмысленным.
ROM|10|20|А Исаия смело говорит: Меня нашли не искавшие Меня; Я открылся не вопрошавшим о Мне.
ROM|10|21|Об Израиле же говорит: целый день Я простирал руки Мои к народу непослушному и упорному.
ROM|11|1|Итак, спрашиваю: неужели Бог отверг народ Свой? Никак. Ибо и я Израильтянин, от семени Авраамова, из колена Вениаминова.
ROM|11|2|Не отверг Бог народа Своего, который Он наперед знал. Или не знаете, что говорит Писание в [повествовании об] Илии? как он жалуется Богу на Израиля, говоря:
ROM|11|3|Господи! пророков Твоих убили, жертвенники Твои разрушили; остался я один, и моей души ищут.
ROM|11|4|Что же говорит ему Божеский ответ? Я соблюл Себе семь тысяч человек, которые не преклонили колени перед Ваалом.
ROM|11|5|Так и в нынешнее время, по избранию благодати, сохранился остаток.
ROM|11|6|Но если по благодати, то не по делам; иначе благодать не была бы уже благодатью. А если по делам, то это уже не благодать; иначе дело не есть уже дело.
ROM|11|7|Что же? Израиль, чего искал, того не получил; избранные же получили, а прочие ожесточились,
ROM|11|8|как написано: Бог дал им дух усыпления, глаза, которыми не видят, и уши, которыми не слышат, даже до сего дня.
ROM|11|9|И Давид говорит: да будет трапеза их сетью, тенетами и петлею в возмездие им;
ROM|11|10|да помрачатся глаза их, чтобы не видеть, и хребет их да будет согбен навсегда.
ROM|11|11|Итак спрашиваю: неужели они преткнулись, чтобы [совсем] пасть? Никак. Но от их падения спасение язычникам, чтобы возбудить в них ревность.
ROM|11|12|Если же падение их – богатство миру, и оскудение их – богатство язычникам, то тем более полнота их.
ROM|11|13|Вам говорю, язычникам. Как Апостол язычников, я прославляю служение мое.
ROM|11|14|Не возбужу ли ревность в [сродниках] моих по плоти и не спасу ли некоторых из них?
ROM|11|15|Ибо если отвержение их – примирение мира, то что [будет] принятие, как не жизнь из мертвых?
ROM|11|16|Если начаток свят, то и целое; и если корень свят, то и ветви.
ROM|11|17|Если же некоторые из ветвей отломились, а ты, дикая маслина, привился на место их и стал общником корня и сока маслины,
ROM|11|18|то не превозносись перед ветвями. Если же превозносишься, [то] [вспомни, что] не ты корень держишь, но корень тебя.
ROM|11|19|Скажешь: "ветви отломились, чтобы мне привиться".
ROM|11|20|Хорошо. Они отломились неверием, а ты держишься верою: не гордись, но бойся.
ROM|11|21|Ибо если Бог не пощадил природных ветвей, то смотри, пощадит ли и тебя.
ROM|11|22|Итак видишь благость и строгость Божию: строгость к отпадшим, а благость к тебе, если пребудешь в благости [Божией]; иначе и ты будешь отсечен.
ROM|11|23|Но и те, если не пребудут в неверии, привьются, потому что Бог силен опять привить их.
ROM|11|24|Ибо если ты отсечен от дикой по природе маслины и не по природе привился к хорошей маслине, то тем более сии природные привьются к своей маслине.
ROM|11|25|Ибо не хочу оставить вас, братия, в неведении о тайне сей, – чтобы вы не мечтали о себе, – что ожесточение произошло в Израиле отчасти, [до времени], пока войдет полное [число] язычников;
ROM|11|26|и так весь Израиль спасется, как написано: придет от Сиона Избавитель, и отвратит нечестие от Иакова.
ROM|11|27|И сей завет им от Меня, когда сниму с них грехи их.
ROM|11|28|В отношении к благовестию, они враги ради вас; а в отношении к избранию, возлюбленные [Божии] ради отцов.
ROM|11|29|Ибо дары и призвание Божие непреложны.
ROM|11|30|Как и вы некогда были непослушны Богу, а ныне помилованы, по непослушанию их,
ROM|11|31|так и они теперь непослушны для помилования вас, чтобы и сами они были помилованы.
ROM|11|32|Ибо всех заключил Бог в непослушание, чтобы всех помиловать.
ROM|11|33|О, бездна богатства и премудрости и ведения Божия! Как непостижимы судьбы Его и неисследимы пути Его!
ROM|11|34|Ибо кто познал ум Господень? Или кто был советником Ему?
ROM|11|35|Или кто дал Ему наперед, чтобы Он должен был воздать?
ROM|11|36|Ибо все из Него, Им и к Нему. Ему слава во веки, аминь.
ROM|12|1|Итак умоляю вас, братия, милосердием Божиим, представьте тела ваши в жертву живую, святую, благоугодную Богу, [для] разумного служения вашего,
ROM|12|2|и не сообразуйтесь с веком сим, но преобразуйтесь обновлением ума вашего, чтобы вам познавать, что есть воля Божия, благая, угодная и совершенная.
ROM|12|3|По данной мне благодати, всякому из вас говорю: не думайте [о] [себе] более, нежели должно думать; но думайте скромно, по мере веры, какую каждому Бог уделил.
ROM|12|4|Ибо, как в одном теле у нас много членов, но не у всех членов одно и то же дело,
ROM|12|5|так мы, многие, составляем одно тело во Христе, а порознь один для другого члены.
ROM|12|6|И как, по данной нам благодати, имеем различные дарования, [то], [имеешь ли] пророчество, [пророчествуй] по мере веры;
ROM|12|7|[имеешь ли] служение, [пребывай] в служении; учитель ли, – в учении;
ROM|12|8|увещатель ли, увещевай; раздаватель ли, [раздавай] в простоте; начальник ли, [начальствуй] с усердием; благотворитель ли, [благотвори] с радушием.
ROM|12|9|Любовь [да будет] непритворна; отвращайтесь зла, прилепляйтесь к добру;
ROM|12|10|будьте братолюбивы друг к другу с нежностью; в почтительности друг друга предупреждайте;
ROM|12|11|в усердии не ослабевайте; духом пламенейте; Господу служите;
ROM|12|12|утешайтесь надеждою; в скорби [будьте] терпеливы, в молитве постоянны;
ROM|12|13|в нуждах святых принимайте участие; ревнуйте о странноприимстве.
ROM|12|14|Благословляйте гонителей ваших; благословляйте, а не проклинайте.
ROM|12|15|Радуйтесь с радующимися и плачьте с плачущими.
ROM|12|16|Будьте единомысленны между собою; не высокомудрствуйте, но последуйте смиренным; не мечтайте о себе;
ROM|12|17|никому не воздавайте злом за зло, но пекитесь о добром перед всеми человеками.
ROM|12|18|Если возможно с вашей стороны, будьте в мире со всеми людьми.
ROM|12|19|Не мстите за себя, возлюбленные, но дайте место гневу [Божию]. Ибо написано: Мне отмщение, Я воздам, говорит Господь.
ROM|12|20|Итак, если враг твой голоден, накорми его; если жаждет, напой его: ибо, делая сие, ты соберешь ему на голову горящие уголья.
ROM|12|21|Не будь побежден злом, но побеждай зло добром.
ROM|13|1|Всякая душа да будет покорна высшим властям, ибо нет власти не от Бога; существующие же власти от Бога установлены.
ROM|13|2|Посему противящийся власти противится Божию установлению. А противящиеся сами навлекут на себя осуждение.
ROM|13|3|Ибо начальствующие страшны не для добрых дел, но для злых. Хочешь ли не бояться власти? Делай добро, и получишь похвалу от нее,
ROM|13|4|ибо [начальник] есть Божий слуга, тебе на добро. Если же делаешь зло, бойся, ибо он не напрасно носит меч: он Божий слуга, отмститель в наказание делающему злое.
ROM|13|5|И потому надобно повиноваться не только из [страха] наказания, но и по совести.
ROM|13|6|Для сего вы и подати платите, ибо они Божии служители, сим самым постоянно занятые.
ROM|13|7|Итак отдавайте всякому должное: кому подать, подать; кому оброк, оброк; кому страх, страх; кому честь, честь.
ROM|13|8|Не оставайтесь должными никому ничем, кроме взаимной любви; ибо любящий другого исполнил закон.
ROM|13|9|Ибо заповеди: не прелюбодействуй, не убивай, не кради, не лжесвидетельствуй, не пожелай [чужого] и все другие заключаются в сем слове: люби ближнего твоего, как самого себя.
ROM|13|10|Любовь не делает ближнему зла; итак любовь есть исполнение закона.
ROM|13|11|Так [поступайте], зная время, что наступил уже час пробудиться нам от сна. Ибо ныне ближе к нам спасение, нежели когда мы уверовали.
ROM|13|12|Ночь прошла, а день приблизился: итак отвергнем дела тьмы и облечемся в оружия света.
ROM|13|13|Как днем, будем вести себя благочинно, не [предаваясь] ни пированиям и пьянству, ни сладострастию и распутству, ни ссорам и зависти;
ROM|13|14|но облекитесь в Господа нашего Иисуса Христа, и попечения о плоти не превращайте в похоти.
ROM|14|1|Немощного в вере принимайте без споров о мнениях.
ROM|14|2|Ибо иной уверен, [что можно] есть все, а немощный ест овощи.
ROM|14|3|Кто ест, не уничижай того, кто не ест; и кто не ест, не осуждай того, кто ест, потому что Бог принял его.
ROM|14|4|Кто ты, осуждающий чужого раба? Перед своим Господом стоит он, или падает. И будет восставлен, ибо силен Бог восставить его.
ROM|14|5|Иной отличает день от дня, а другой судит о всяком дне [равно]. Всякий [поступай] по удостоверению своего ума.
ROM|14|6|Кто различает дни, для Господа различает; и кто не различает дней, для Господа не различает. Кто ест, для Господа ест, ибо благодарит Бога; и кто не ест, для Господа не ест, и благодарит Бога.
ROM|14|7|Ибо никто из нас не живет для себя, и никто не умирает для себя;
ROM|14|8|а живем ли – для Господа живем; умираем ли – для Господа умираем: и потому, живем ли или умираем, – [всегда] Господни.
ROM|14|9|Ибо Христос для того и умер, и воскрес, и ожил, чтобы владычествовать и над мертвыми и над живыми.
ROM|14|10|А ты что осуждаешь брата твоего? Или и ты, что унижаешь брата твоего? Все мы предстанем на суд Христов.
ROM|14|11|Ибо написано: живу Я, говорит Господь, предо Мною преклонится всякое колено, и всякий язык будет исповедывать Бога.
ROM|14|12|Итак каждый из нас за себя даст отчет Богу.
ROM|14|13|Не станем же более судить друг друга, а лучше судите о том, как бы не подавать брату [случая к] преткновению или соблазну.
ROM|14|14|Я знаю и уверен в Господе Иисусе, что нет ничего в себе самом нечистого; только почитающему что–либо нечистым, тому нечисто.
ROM|14|15|Если же за пищу огорчается брат твой, то ты уже не по любви поступаешь. Не губи твоею пищею того, за кого Христос умер.
ROM|14|16|Да не хулится ваше доброе.
ROM|14|17|Ибо Царствие Божие не пища и питие, но праведность и мир и радость во Святом Духе.
ROM|14|18|Кто сим служит Христу, тот угоден Богу и [достоин] одобрения от людей.
ROM|14|19|Итак будем искать того, что служит к миру и ко взаимному назиданию.
ROM|14|20|Ради пищи не разрушай дела Божия. Все чисто, но худо человеку, который ест на соблазн.
ROM|14|21|Лучше не есть мяса, не пить вина и не [делать] ничего [такого], отчего брат твой претыкается, или соблазняется, или изнемогает.
ROM|14|22|Ты имеешь веру? имей ее сам в себе, пред Богом. Блажен, кто не осуждает себя в том, что избирает.
ROM|14|23|А сомневающийся, если ест, осуждается, потому что не по вере; а все, что не по вере, грех.
ROM|14|24|Могущему же утвердить вас, по благовествованию моему и проповеди Иисуса Христа, по откровению тайны, о которой от вечных времен было умолчано,
ROM|14|25|но которая ныне явлена, и через писания пророческие, по повелению вечного Бога, возвещена всем народам для покорения их вере,
ROM|14|26|Единому Премудрому Богу, через Иисуса Христа, слава во веки. Аминь.
ROM|15|1|Мы, сильные, должны сносить немощи бессильных и не себе угождать.
ROM|15|2|Каждый из нас должен угождать ближнему, во благо, к назиданию.
ROM|15|3|Ибо и Христос не Себе угождал, но, как написано: злословия злословящих Тебя пали на Меня.
ROM|15|4|А все, что писано было прежде, написано нам в наставление, чтобы мы терпением и утешением из Писаний сохраняли надежду.
ROM|15|5|Бог же терпения и утешения да дарует вам быть в единомыслии между собою, по [учению] Христа Иисуса,
ROM|15|6|дабы вы единодушно, едиными устами славили Бога и Отца Господа нашего Иисуса Христа.
ROM|15|7|Посему принимайте друг друга, как и Христос принял вас в славу Божию.
ROM|15|8|Разумею то, что Иисус Христос сделался служителем для обрезанных – ради истины Божией, чтобы исполнить обещанное отцам,
ROM|15|9|а для язычников – из милости, чтобы славили Бога, как написано: за то буду славить Тебя, (Господи,) между язычниками, и буду петь имени Твоему.
ROM|15|10|И еще сказано: возвеселитесь, язычники, с народом Его.
ROM|15|11|И еще: хвалите Господа, все язычники, и прославляйте Его, все народы.
ROM|15|12|Исаия также говорит: будет корень Иессеев, и восстанет владеть народами; на Него язычники надеяться будут.
ROM|15|13|Бог же надежды да исполнит вас всякой радости и мира в вере, дабы вы, силою Духа Святаго, обогатились надеждою.
ROM|15|14|И сам я уверен о вас, братия мои, что и вы полны благости, исполнены всякого познания и можете наставлять друг друга;
ROM|15|15|но писал вам, братия, с некоторою смелостью, отчасти как бы в напоминание вам, по данной мне от Бога благодати
ROM|15|16|быть служителем Иисуса Христа у язычников и [совершать] священнодействие благовествования Божия, дабы сие приношение язычников, будучи освящено Духом Святым, было благоприятно [Богу].
ROM|15|17|Итак я могу похвалиться в Иисусе Христе в том, что [относится] к Богу,
ROM|15|18|ибо не осмелюсь сказать что–нибудь такое, чего не совершил Христос через меня, в покорении язычников [вере], словом и делом,
ROM|15|19|силою знамений и чудес, силою Духа Божия, так что благовествование Христово распространено мною от Иерусалима и окрестности до Иллирика.
ROM|15|20|Притом я старался благовествовать не там, где [уже] было известно имя Христово, дабы не созидать на чужом основании,
ROM|15|21|но как написано: не имевшие о Нем известия увидят, и не слышавшие узнают.
ROM|15|22|Сие–то много раз и препятствовало мне придти к вам.
ROM|15|23|Ныне же, не имея [такого] места в сих странах, а с давних лет имея желание придти к вам,
ROM|15|24|как только предприму путь в Испанию, приду к вам. Ибо надеюсь, что, проходя, увижусь с вами и что вы проводите меня туда, как скоро наслажусь [общением] с вами, хотя отчасти.
ROM|15|25|А теперь я иду в Иерусалим, чтобы послужить святым,
ROM|15|26|ибо Македония и Ахаия усердствуют некоторым подаянием для бедных между святыми в Иерусалиме.
ROM|15|27|Усердствуют, да и должники они перед ними. Ибо если язычники сделались участниками в их духовном, то должны и им послужить в телесном.
ROM|15|28|Исполнив это и верно доставив им сей плод [усердия], я отправлюсь через ваши [места] в Испанию,
ROM|15|29|и уверен, что когда приду к вам, то приду с полным благословением благовествования Христова.
ROM|15|30|Между тем умоляю вас, братия, Господом нашим Иисусом Христом и любовью Духа, подвизаться со мною в молитвах за меня к Богу,
ROM|15|31|чтобы избавиться мне от неверующих в Иудее и чтобы служение мое для Иерусалима было благоприятно святым,
ROM|15|32|дабы мне в радости, если Богу угодно, придти к вам и успокоиться с вами.
ROM|15|33|Бог же мира да будет со всеми вами, аминь.
ROM|16|1|Представляю вам Фиву, сестру нашу, диакониссу церкви Кенхрейской.
ROM|16|2|Примите ее для Господа, как прилично святым, и помогите ей, в чем она будет иметь нужду у вас, ибо и она была помощницею многим и мне самому.
ROM|16|3|Приветствуйте Прискиллу и Акилу, сотрудников моих во Христе Иисусе
ROM|16|4|(которые голову свою полагали за мою душу, которых не я один благодарю, но и все церкви из язычников), и домашнюю их церковь.
ROM|16|5|Приветствуйте возлюбленного моего Епенета, который есть начаток Ахаии для Христа.
ROM|16|6|Приветствуйте Мариам, которая много трудилась для нас.
ROM|16|7|Приветствуйте Андроника и Юнию, сродников моих и узников со мною, прославившихся между Апостолами и прежде меня еще уверовавших во Христа.
ROM|16|8|Приветствуйте Амплия, возлюбленного мне в Господе.
ROM|16|9|Приветствуйте Урбана, сотрудника нашего во Христе, и Стахия, возлюбленного мне.
ROM|16|10|Приветствуйте Апеллеса, испытанного во Христе. Приветствуйте [верных] из дома Аристовулова.
ROM|16|11|Приветствуйте Иродиона, сродника моего. Приветствуйте из домашних Наркисса тех, которые в Господе.
ROM|16|12|Приветствуйте Трифену и Трифосу, трудящихся о Господе. Приветствуйте Персиду возлюбленную, которая много потрудилась о Господе.
ROM|16|13|Приветствуйте Руфа, избранного в Господе, и матерь его и мою.
ROM|16|14|Приветствуйте Асинкрита, Флегонта, Ерма, Патрова, Ермия и других с ними братьев.
ROM|16|15|Приветствуйте Филолога и Юлию, Нирея и сестру его, и Олимпана, и всех с ними святых.
ROM|16|16|Приветствуйте друг друга с целованием святым. Приветствуют вас все церкви Христовы.
ROM|16|17|Умоляю вас, братия, остерегайтесь производящих разделения и соблазны, вопреки учению, которому вы научились, и уклоняйтесь от них;
ROM|16|18|ибо такие [люди] служат не Господу нашему Иисусу Христу, а своему чреву, и ласкательством и красноречием обольщают сердца простодушных.
ROM|16|19|Ваша покорность [вере] всем известна; посему я радуюсь за вас, но желаю, чтобы вы были мудры на добро и просты на зло.
ROM|16|20|Бог же мира сокрушит сатану под ногами вашими вскоре. Благодать Господа нашего Иисуса Христа с вами! Аминь.
ROM|16|21|Приветствуют вас Тимофей, сотрудник мой, и Луций, Иасон и Сосипатр, сродники мои.
ROM|16|22|Приветствую вас в Господе и я, Тертий, писавший сие послание.
ROM|16|23|Приветствует вас Гаий, странноприимец мой и всей церкви. Приветствует вас Ераст, городской казнохранитель, и брат Кварт.
ROM|16|24|Благодать Господа нашего Иисуса Христа со всеми вами. Аминь.
