1COR|1|1|Павел, волею Божиею призванный Апостол Иисуса Христа, и Сосфен брат,
1COR|1|2|церкви Божией, находящейся в Коринфе, освященным во Христе Иисусе, призванным святым, со всеми призывающими имя Господа нашего Иисуса Христа, во всяком месте, у них и у нас:
1COR|1|3|благодать вам и мир от Бога Отца нашего и Господа Иисуса Христа.
1COR|1|4|Непрестанно благодарю Бога моего за вас, ради благодати Божией, дарованной вам во Христе Иисусе,
1COR|1|5|потому что в Нем вы обогатились всем, всяким словом и всяким познанием, –
1COR|1|6|ибо свидетельство Христово утвердилось в вас, –
1COR|1|7|так что вы не имеете недостатка ни в каком даровании, ожидая явления Господа нашего Иисуса Христа,
1COR|1|8|Который и утвердит вас до конца, [чтобы вам быть] неповинными в день Господа нашего Иисуса Христа.
1COR|1|9|Верен Бог, Которым вы призваны в общение Сына Его Иисуса Христа, Господа нашего.
1COR|1|10|Умоляю вас, братия, именем Господа нашего Иисуса Христа, чтобы все вы говорили одно, и не было между вами разделений, но чтобы вы соединены были в одном духе и в одних мыслях.
1COR|1|11|Ибо от [домашних] Хлоиных сделалось мне известным о вас, братия мои, что между вами есть споры.
1COR|1|12|Я разумею то, что у вас говорят: "я Павлов"; "я Аполлосов"; "я Кифин"; "а я Христов".
1COR|1|13|Разве разделился Христос? разве Павел распялся за вас? или во имя Павла вы крестились?
1COR|1|14|Благодарю Бога, что я никого из вас не крестил, кроме Криспа и Гаия,
1COR|1|15|дабы не сказал кто, что я крестил в мое имя.
1COR|1|16|Крестил я также Стефанов дом; а крестил ли еще кого, не знаю.
1COR|1|17|Ибо Христос послал меня не крестить, а благовествовать, не в премудрости слова, чтобы не упразднить креста Христова.
1COR|1|18|Ибо слово о кресте для погибающих юродство есть, а для нас, спасаемых, – сила Божия.
1COR|1|19|Ибо написано: погублю мудрость мудрецов, и разум разумных отвергну.
1COR|1|20|Где мудрец? где книжник? где совопросник века сего? Не обратил ли Бог мудрость мира сего в безумие?
1COR|1|21|Ибо когда мир [своею] мудростью не познал Бога в премудрости Божией, то благоугодно было Богу юродством проповеди спасти верующих.
1COR|1|22|Ибо и Иудеи требуют чудес, и Еллины ищут мудрости;
1COR|1|23|а мы проповедуем Христа распятого, для Иудеев соблазн, а для Еллинов безумие,
1COR|1|24|для самих же призванных, Иудеев и Еллинов, Христа, Божию силу и Божию премудрость;
1COR|1|25|потому что немудрое Божие премудрее человеков, и немощное Божие сильнее человеков.
1COR|1|26|Посмотрите, братия, кто вы, призванные: не много [из вас] мудрых по плоти, не много сильных, не много благородных;
1COR|1|27|но Бог избрал немудрое мира, чтобы посрамить мудрых, и немощное мира избрал Бог, чтобы посрамить сильное;
1COR|1|28|и незнатное мира и уничиженное и ничего не значащее избрал Бог, чтобы упразднить значащее, –
1COR|1|29|для того, чтобы никакая плоть не хвалилась пред Богом.
1COR|1|30|От Него и вы во Христе Иисусе, Который сделался для нас премудростью от Бога, праведностью и освящением и искуплением,
1COR|1|31|чтобы [было], как написано: хвалящийся хвались Господом.
1COR|2|1|И когда я приходил к вам, братия, приходил возвещать вам свидетельство Божие не в превосходстве слова или мудрости,
1COR|2|2|ибо я рассудил быть у вас незнающим ничего, кроме Иисуса Христа, и притом распятого,
1COR|2|3|и был я у вас в немощи и в страхе и в великом трепете.
1COR|2|4|И слово мое и проповедь моя не в убедительных словах человеческой мудрости, но в явлении духа и силы,
1COR|2|5|чтобы вера ваша [утверждалась] не на мудрости человеческой, но на силе Божией.
1COR|2|6|Мудрость же мы проповедуем между совершенными, но мудрость не века сего и не властей века сего преходящих,
1COR|2|7|но проповедуем премудрость Божию, тайную, сокровенную, которую предназначил Бог прежде веков к славе нашей,
1COR|2|8|которой никто из властей века сего не познал; ибо если бы познали, то не распяли бы Господа славы.
1COR|2|9|Но, как написано: не видел того глаз, не слышало ухо, и не приходило то на сердце человеку, что приготовил Бог любящим Его.
1COR|2|10|А нам Бог открыл [это] Духом Своим; ибо Дух все проницает, и глубины Божии.
1COR|2|11|Ибо кто из человеков знает, что в человеке, кроме духа человеческого, живущего в нем? Так и Божьего никто не знает, кроме Духа Божия.
1COR|2|12|Но мы приняли не духа мира сего, а Духа от Бога, дабы знать дарованное нам от Бога,
1COR|2|13|что и возвещаем не от человеческой мудрости изученными словами, но изученными от Духа Святаго, соображая духовное с духовным.
1COR|2|14|Душевный человек не принимает того, что от Духа Божия, потому что он почитает это безумием; и не может разуметь, потому что о сем [надобно] судить духовно.
1COR|2|15|Но духовный судит о всем, а о нем судить никто не может.
1COR|2|16|Ибо кто познал ум Господень, чтобы [мог] судить его? А мы имеем ум Христов.
1COR|3|1|И я не мог говорить с вами, братия, как с духовными, но как с плотскими, как с младенцами во Христе.
1COR|3|2|Я питал вас молоком, а не [твердою] пищею, ибо вы были еще не в силах, да и теперь не в силах,
1COR|3|3|потому что вы еще плотские. Ибо если между вами зависть, споры и разногласия, то не плотские ли вы? и не по человеческому ли [обычаю] поступаете?
1COR|3|4|Ибо когда один говорит: "я Павлов", а другой: "я Аполлосов", то не плотские ли вы?
1COR|3|5|Кто Павел? кто Аполлос? Они только служители, через которых вы уверовали, и притом поскольку каждому дал Господь.
1COR|3|6|Я насадил, Аполлос поливал, но возрастил Бог;
1COR|3|7|посему и насаждающий и поливающий есть ничто, а [все] Бог возращающий.
1COR|3|8|Насаждающий же и поливающий суть одно; но каждый получит свою награду по своему труду.
1COR|3|9|Ибо мы соработники у Бога, [а] вы Божия нива, Божие строение.
1COR|3|10|Я, по данной мне от Бога благодати, как мудрый строитель, положил основание, а другой строит на [нем]; но каждый смотри, как строит.
1COR|3|11|Ибо никто не может положить другого основания, кроме положенного, которое есть Иисус Христос.
1COR|3|12|Строит ли кто на этом основании из золота, серебра, драгоценных камней, дерева, сена, соломы, –
1COR|3|13|каждого дело обнаружится; ибо день покажет, потому что в огне открывается, и огонь испытает дело каждого, каково оно есть.
1COR|3|14|У кого дело, которое он строил, устоит, тот получит награду.
1COR|3|15|А у кого дело сгорит, тот потерпит урон; впрочем сам спасется, но так, как бы из огня.
1COR|3|16|Разве не знаете, что вы храм Божий, и Дух Божий живет в вас?
1COR|3|17|Если кто разорит храм Божий, того покарает Бог: ибо храм Божий свят; а этот [храм] – вы.
1COR|3|18|Никто не обольщай самого себя. Если кто из вас думает быть мудрым в веке сем, тот будь безумным, чтобы быть мудрым.
1COR|3|19|Ибо мудрость мира сего есть безумие пред Богом, как написано: уловляет мудрых в лукавстве их.
1COR|3|20|И еще: Господь знает умствования мудрецов, что они суетны.
1COR|3|21|Итак никто не хвались человеками, ибо все ваше:
1COR|3|22|Павел ли, или Аполлос, или Кифа, или мир, или жизнь, или смерть, или настоящее, или будущее, – все ваше;
1COR|3|23|вы же – Христовы, а Христос – Божий.
1COR|4|1|Итак каждый должен разуметь нас, как служителей Христовых и домостроителей таин Божиих.
1COR|4|2|От домостроителей же требуется, чтобы каждый оказался верным.
1COR|4|3|Для меня очень мало значит, как судите обо мне вы или [как] [судят] другие люди; я и сам не сужу о себе.
1COR|4|4|Ибо [хотя] я ничего не знаю за собою, но тем не оправдываюсь; судия же мне Господь.
1COR|4|5|Посему не судите никак прежде времени, пока не придет Господь, Который и осветит скрытое во мраке и обнаружит сердечные намерения, и тогда каждому будет похвала от Бога.
1COR|4|6|Это, братия, приложил я к себе и Аполлосу ради вас, чтобы вы научились от нас не мудрствовать сверх того, что написано, и не превозносились один перед другим.
1COR|4|7|Ибо кто отличает тебя? Что ты имеешь, чего бы не получил? А если получил, что хвалишься, как будто не получил?
1COR|4|8|Вы уже пресытились, вы уже обогатились, вы стали царствовать без нас. О, если бы вы [и в самом деле] царствовали, чтобы и нам с вами царствовать!
1COR|4|9|Ибо я думаю, что нам, последним посланникам, Бог судил быть как бы приговоренными к смерти, потому что мы сделались позорищем для мира, для Ангелов и человеков.
1COR|4|10|Мы безумны Христа ради, а вы мудры во Христе; мы немощны, а вы крепки; вы в славе, а мы в бесчестии.
1COR|4|11|Даже доныне терпим голод и жажду, и наготу и побои, и скитаемся,
1COR|4|12|и трудимся, работая своими руками. Злословят нас, мы благословляем; гонят нас, мы терпим;
1COR|4|13|хулят нас, мы молим; мы как сор для мира, [как] прах, всеми [попираемый] доныне.
1COR|4|14|Не к постыжению вашему пишу сие, но вразумляю вас, как возлюбленных детей моих.
1COR|4|15|Ибо, хотя у вас тысячи наставников во Христе, но не много отцов; я родил вас во Христе Иисусе благовествованием.
1COR|4|16|Посему умоляю вас: подражайте мне, как я Христу.
1COR|4|17|Для сего я послал к вам Тимофея, моего возлюбленного и верного в Господе сына, который напомнит вам о путях моих во Христе, как я учу везде во всякой церкви.
1COR|4|18|Как я не иду к вам, то некоторые [у вас] возгордились;
1COR|4|19|но я скоро приду к вам, если угодно будет Господу, и испытаю не слова возгордившихся, а силу,
1COR|4|20|ибо Царство Божие не в слове, а в силе.
1COR|4|21|Чего вы хотите? с жезлом придти к вам, или с любовью и духом кротости?
1COR|5|1|Есть верный слух, что у вас [появилось] блудодеяние, и притом такое блудодеяние, какого не слышно даже у язычников, что некто [вместо] [жены] имеет жену отца своего.
1COR|5|2|И вы возгордились, вместо того, чтобы лучше плакать, дабы изъят был из среды вас сделавший такое дело.
1COR|5|3|А я, отсутствуя телом, но присутствуя [у вас] духом, уже решил, как бы находясь у вас: сделавшего такое дело,
1COR|5|4|в собрании вашем во имя Господа нашего Иисуса Христа, обще с моим духом, силою Господа нашего Иисуса Христа,
1COR|5|5|предать сатане во измождение плоти, чтобы дух был спасен в день Господа нашего Иисуса Христа.
1COR|5|6|Нечем вам хвалиться. Разве не знаете, что малая закваска квасит все тесто?
1COR|5|7|Итак очистите старую закваску, чтобы быть вам новым тестом, так как вы бесквасны, ибо Пасха наша, Христос, заклан за нас.
1COR|5|8|Посему станем праздновать не со старою закваскою, не с закваскою порока и лукавства, но с опресноками чистоты и истины.
1COR|5|9|Я писал вам в послании – не сообщаться с блудниками;
1COR|5|10|впрочем не вообще с блудниками мира сего, или лихоимцами, или хищниками, или идолослужителями, ибо иначе надлежало бы вам выйти из мира [сего].
1COR|5|11|Но я писал вам не сообщаться с тем, кто, называясь братом, остается блудником, или лихоимцем, или идолослужителем, или злоречивым, или пьяницею, или хищником; с таким даже и не есть вместе.
1COR|5|12|Ибо что мне судить и внешних? Не внутренних ли вы судите?
1COR|5|13|Внешних же судит Бог. Итак, извергните развращенного из среды вас.
1COR|6|1|Как смеет кто у вас, имея дело с другим, судиться у нечестивых, а не у святых?
1COR|6|2|Разве не знаете, что святые будут судить мир? Если же вами будет судим мир, то неужели вы недостойны судить маловажные [дела]?
1COR|6|3|Разве не знаете, что мы будем судить ангелов, не тем ли более [дела] житейские?
1COR|6|4|А вы, когда имеете житейские тяжбы, поставляете [своими судьями] ничего не значащих в церкви.
1COR|6|5|К стыду вашему говорю: неужели нет между вами ни одного разумного, который мог бы рассудить между братьями своими?
1COR|6|6|Но брат с братом судится, и притом перед неверными.
1COR|6|7|И то уже весьма унизительно для вас, что вы имеете тяжбы между собою. Для чего бы вам лучше не оставаться обиженными? для чего бы вам лучше не терпеть лишения?
1COR|6|8|Но вы [сами] обижаете и отнимаете, и притом у братьев.
1COR|6|9|Или не знаете, что неправедные Царства Божия не наследуют? Не обманывайтесь: ни блудники, ни идолослужители, ни прелюбодеи, ни малакии, ни мужеложники,
1COR|6|10|ни воры, ни лихоимцы, ни пьяницы, ни злоречивые, ни хищники – Царства Божия не наследуют.
1COR|6|11|И такими были некоторые из вас; но омылись, но освятились, но оправдались именем Господа нашего Иисуса Христа и Духом Бога нашего.
1COR|6|12|Все мне позволительно, но не все полезно; все мне позволительно, но ничто не должно обладать мною.
1COR|6|13|Пища для чрева, и чрево для пищи; но Бог уничтожит и то и другое. Тело же не для блуда, но для Господа, и Господь для тела.
1COR|6|14|Бог воскресил Господа, воскресит и нас силою Своею.
1COR|6|15|Разве не знаете, что тела ваши суть члены Христовы? Итак отниму ли члены у Христа, чтобы сделать [их] членами блудницы? Да не будет!
1COR|6|16|Или не знаете, что совокупляющийся с блудницею становится одно тело [с нею]? ибо сказано: два будут одна плоть.
1COR|6|17|А соединяющийся с Господом есть один дух с Господом.
1COR|6|18|Бегайте блуда; всякий грех, какой делает человек, есть вне тела, а блудник грешит против собственного тела.
1COR|6|19|Не знаете ли, что тела ваши суть храм живущего в вас Святаго Духа, Которого имеете вы от Бога, и вы не свои?
1COR|6|20|Ибо вы куплены [дорогою] ценою. Посему прославляйте Бога и в телах ваших и в душах ваших, которые суть Божии.
1COR|7|1|А о чем вы писали ко мне, то хорошо человеку не касаться женщины.
1COR|7|2|Но, [во избежание] блуда, каждый имей свою жену, и каждая имей своего мужа.
1COR|7|3|Муж оказывай жене должное благорасположение; подобно и жена мужу.
1COR|7|4|Жена не властна над своим телом, но муж; равно и муж не властен над своим телом, но жена.
1COR|7|5|Не уклоняйтесь друг от друга, разве по согласию, на время, для упражнения в посте и молитве, а [потом] опять будьте вместе, чтобы не искушал вас сатана невоздержанием вашим.
1COR|7|6|Впрочем это сказано мною как позволение, а не как повеление.
1COR|7|7|Ибо желаю, чтобы все люди были, как и я; но каждый имеет свое дарование от Бога, один так, другой иначе.
1COR|7|8|Безбрачным же и вдовам говорю: хорошо им оставаться, как я.
1COR|7|9|Но если не [могут] воздержаться, пусть вступают в брак; ибо лучше вступить в брак, нежели разжигаться.
1COR|7|10|А вступившим в брак не я повелеваю, а Господь: жене не разводиться с мужем, –
1COR|7|11|если же разведется, то должна оставаться безбрачною, или примириться с мужем своим, – и мужу не оставлять жены [своей].
1COR|7|12|Прочим же я говорю, а не Господь: если какой брат имеет жену неверующую, и она согласна жить с ним, то он не должен оставлять ее;
1COR|7|13|и жена, которая имеет мужа неверующего, и он согласен жить с нею, не должна оставлять его.
1COR|7|14|Ибо неверующий муж освящается женою верующею, и жена неверующая освящается мужем верующим. Иначе дети ваши были бы нечисты, а теперь святы.
1COR|7|15|Если же неверующий [хочет] развестись, пусть разводится; брат или сестра в таких [случаях] не связаны; к миру призвал нас Господь.
1COR|7|16|Почему ты знаешь, жена, не спасешь ли мужа? Или ты, муж, почему знаешь, не спасешь ли жены?
1COR|7|17|Только каждый поступай так, как Бог ему определил, и каждый, как Господь призвал. Так я повелеваю по всем церквам.
1COR|7|18|Призван ли кто обрезанным, не скрывайся; призван ли кто необрезанным, не обрезывайся.
1COR|7|19|Обрезание ничто и необрезание ничто, но [все] в соблюдении заповедей Божиих.
1COR|7|20|Каждый оставайся в том звании, в котором призван.
1COR|7|21|Рабом ли ты призван, не смущайся; но если и можешь сделаться свободным, то лучшим воспользуйся.
1COR|7|22|Ибо раб, призванный в Господе, есть свободный Господа; равно и призванный свободным есть раб Христов.
1COR|7|23|Вы куплены [дорогою] ценою; не делайтесь рабами человеков.
1COR|7|24|В каком [звании] кто призван, братия, в том каждый и оставайся пред Богом.
1COR|7|25|Относительно девства я не имею повеления Господня, а даю совет, как получивший от Господа милость быть [Ему] верным.
1COR|7|26|По настоящей нужде за лучшее признаю, что хорошо человеку оставаться так.
1COR|7|27|Соединен ли ты с женой? не ищи развода. Остался ли без жены? не ищи жены.
1COR|7|28|Впрочем, если и женишься, не согрешишь; и если девица выйдет замуж, не согрешит. Но таковые будут иметь скорби по плоти; а мне вас жаль.
1COR|7|29|Я вам сказываю, братия: время уже коротко, так что имеющие жен должны быть, как не имеющие;
1COR|7|30|и плачущие, как не плачущие; и радующиеся, как не радующиеся; и покупающие, как не приобретающие;
1COR|7|31|и пользующиеся миром сим, как не пользующиеся; ибо проходит образ мира сего.
1COR|7|32|А я хочу, чтобы вы были без забот. Неженатый заботится о Господнем, как угодить Господу;
1COR|7|33|а женатый заботится о мирском, как угодить жене. Есть разность между замужнею и девицею:
1COR|7|34|незамужняя заботится о Господнем, как угодить Господу, чтобы быть святою и телом и духом; а замужняя заботится о мирском, как угодить мужу.
1COR|7|35|Говорю это для вашей же пользы, не с тем, чтобы наложить на вас узы, но чтобы вы благочинно и непрестанно [служили] Господу без развлечения.
1COR|7|36|Если же кто почитает неприличным для своей девицы то, чтобы она, будучи в зрелом возрасте, оставалась так, тот пусть делает, как хочет: не согрешит; пусть [таковые] выходят замуж.
1COR|7|37|Но кто непоколебимо тверд в сердце своем и, не будучи стесняем нуждою, но будучи властен в своей воле, решился в сердце своем соблюдать свою деву, тот хорошо поступает.
1COR|7|38|Посему выдающий замуж свою девицу поступает хорошо; а не выдающий поступает лучше.
1COR|7|39|Жена связана законом, доколе жив муж ее; если же муж ее умрет, свободна выйти, за кого хочет, только в Господе.
1COR|7|40|Но она блаженнее, если останется так, по моему совету; а думаю, и я имею Духа Божия.
1COR|8|1|О идоложертвенных [яствах] мы знаем, потому что мы все имеем знание; но знание надмевает, а любовь назидает.
1COR|8|2|Кто думает, что он знает что–нибудь, тот ничего еще не знает так, как должно знать.
1COR|8|3|Но кто любит Бога, тому дано знание от Него.
1COR|8|4|Итак об употреблении в пищу идоложертвенного мы знаем, что идол в мире ничто, и что нет иного Бога, кроме Единого.
1COR|8|5|Ибо хотя и есть так называемые боги, или на небе, или на земле, так как есть много богов и господ много, –
1COR|8|6|но у нас один Бог Отец, из Которого все, и мы для Него, и один Господь Иисус Христос, Которым все, и мы Им.
1COR|8|7|Но не у всех [такое] знание: некоторые и доныне с совестью, [признающею] идолов, едят [идоложертвенное] как жертвы идольские, и совесть их, будучи немощна, оскверняется.
1COR|8|8|Пища не приближает нас к Богу: ибо, едим ли мы, ничего не приобретаем; не едим ли, ничего не теряем.
1COR|8|9|Берегитесь однако же, чтобы эта свобода ваша не послужила соблазном для немощных.
1COR|8|10|Ибо если кто–нибудь увидит, что ты, имея знание, сидишь за столом в капище, то совесть его, как немощного, не расположит ли и его есть идоложертвенное?
1COR|8|11|И от знания твоего погибнет немощный брат, за которого умер Христос.
1COR|8|12|А согрешая таким образом против братьев и уязвляя немощную совесть их, вы согрешаете против Христа.
1COR|8|13|И потому, если пища соблазняет брата моего, не буду есть мяса вовек, чтобы не соблазнить брата моего.
1COR|9|1|Не Апостол ли я? Не свободен ли я? Не видел ли я Иисуса Христа, Господа нашего? Не мое ли дело вы в Господе?
1COR|9|2|Если для других я не Апостол, то для вас [Апостол]; ибо печать моего апостольства – вы в Господе.
1COR|9|3|Вот мое защищение против осуждающих меня.
1COR|9|4|Или мы не имеем власти есть и пить?
1COR|9|5|Или не имеем власти иметь спутницею сестру жену, как и прочие Апостолы, и братья Господни, и Кифа?
1COR|9|6|Или один я и Варнава не имеем власти не работать?
1COR|9|7|Какой воин служит когда–либо на своем содержании? Кто, насадив виноград, не ест плодов его? Кто, пася стадо, не ест молока от стада?
1COR|9|8|По человеческому ли только [рассуждению] я это говорю? Не то же ли говорит и закон?
1COR|9|9|Ибо в Моисеевом законе написано: не заграждай рта у вола молотящего. О волах ли печется Бог?
1COR|9|10|Или, конечно, для нас говорится? Так, для нас это написано; ибо, кто пашет, должен пахать с надеждою, и кто молотит, [должен молотить] с надеждою получить ожидаемое.
1COR|9|11|Если мы посеяли в вас духовное, велико ли то, если пожнем у вас телесное?
1COR|9|12|Если другие имеют у вас власть, не паче ли мы? Однако мы не пользовались сею властью, но все переносим, дабы не поставить какой преграды благовествованию Христову.
1COR|9|13|Разве не знаете, что священнодействующие питаются от святилища? что служащие жертвеннику берут долю от жертвенника?
1COR|9|14|Так и Господь повелел проповедующим Евангелие жить от благовествования.
1COR|9|15|Но я не пользовался ничем таковым. И написал это не для того, чтобы так было для меня. Ибо для меня лучше умереть, нежели чтобы кто уничтожил похвалу мою.
1COR|9|16|Ибо если я благовествую, то нечем мне хвалиться, потому что это необходимая [обязанность] моя, и горе мне, если не благовествую!
1COR|9|17|Ибо если делаю это добровольно, то [буду] иметь награду; а если недобровольно, то [исполняю только] вверенное мне служение.
1COR|9|18|За что же мне награда? За то, что, проповедуя Евангелие, благовествую о Христе безмездно, не пользуясь моею властью в благовествовании.
1COR|9|19|Ибо, будучи свободен от всех, я всем поработил себя, дабы больше приобрести:
1COR|9|20|для Иудеев я был как Иудей, чтобы приобрести Иудеев; для подзаконных был как подзаконный, чтобы приобрести подзаконных;
1COR|9|21|для чуждых закона – как чуждый закона, – не будучи чужд закона пред Богом, но подзаконен Христу, – чтобы приобрести чуждых закона;
1COR|9|22|для немощных был как немощный, чтобы приобрести немощных. Для всех я сделался всем, чтобы спасти по крайней мере некоторых.
1COR|9|23|Сие же делаю для Евангелия, чтобы быть соучастником его.
1COR|9|24|Не знаете ли, что бегущие на ристалище бегут все, но один получает награду? Так бегите, чтобы получить.
1COR|9|25|Все подвижники воздерживаются от всего: те для получения венца тленного, а мы – нетленного.
1COR|9|26|И потому я бегу не так, как на неверное, бьюсь не так, чтобы только бить воздух;
1COR|9|27|но усмиряю и порабощаю тело мое, дабы, проповедуя другим, самому не остаться недостойным.
1COR|10|1|Не хочу оставить вас, братия, в неведении, что отцы наши все были под облаком, и все прошли сквозь море;
1COR|10|2|и все крестились в Моисея в облаке и в море;
1COR|10|3|и все ели одну и ту же духовную пищу;
1COR|10|4|и все пили одно и то же духовное питие: ибо пили из духовного последующего камня; камень же был Христос.
1COR|10|5|Но не о многих из них благоволил Бог, ибо они поражены были в пустыне.
1COR|10|6|А это были образы для нас, чтобы мы не были похотливы на злое, как они были похотливы.
1COR|10|7|Не будьте также идолопоклонниками, как некоторые из них, о которых написано: народ сел есть и пить, и встал играть.
1COR|10|8|Не станем блудодействовать, как некоторые из них блудодействовали, и в один день погибло их двадцать три тысячи.
1COR|10|9|Не станем искушать Христа, как некоторые из них искушали и погибли от змей.
1COR|10|10|Не ропщите, как некоторые из них роптали и погибли от истребителя.
1COR|10|11|Все это происходило с ними, [как] образы; а описано в наставление нам, достигшим последних веков.
1COR|10|12|Посему, кто думает, что он стоит, берегись, чтобы не упасть.
1COR|10|13|Вас постигло искушение не иное, как человеческое; и верен Бог, Который не попустит вам быть искушаемыми сверх сил, но при искушении даст и облегчение, так чтобы вы могли перенести.
1COR|10|14|Итак, возлюбленные мои, убегайте идолослужения.
1COR|10|15|Я говорю [вам] как рассудительным; сами рассудите о том, что говорю.
1COR|10|16|Чаша благословения, которую благословляем, не есть ли приобщение Крови Христовой? Хлеб, который преломляем, не есть ли приобщение Тела Христова?
1COR|10|17|Один хлеб, и мы многие одно тело; ибо все причащаемся от одного хлеба.
1COR|10|18|Посмотрите на Израиля по плоти: те, которые едят жертвы, не участники ли жертвенника?
1COR|10|19|Что же я говорю? То ли, что идол есть что–нибудь, или идоложертвенное значит что–нибудь?
1COR|10|20|[Нет], но что язычники, принося жертвы, приносят бесам, а не Богу. Но я не хочу, чтобы вы были в общении с бесами.
1COR|10|21|Не можете пить чашу Господню и чашу бесовскую; не можете быть участниками в трапезе Господней и в трапезе бесовской.
1COR|10|22|Неужели мы [решимся] раздражать Господа? Разве мы сильнее Его?
1COR|10|23|Все мне позволительно, но не все полезно; все мне позволительно, но не все назидает.
1COR|10|24|Никто не ищи своего, но каждый [пользы] другого.
1COR|10|25|Все, что продается на торгу, ешьте без всякого исследования, для [спокойствия] совести;
1COR|10|26|ибо Господня земля, и что наполняет ее.
1COR|10|27|Если кто из неверных позовет вас, и вы захотите пойти, то все, предлагаемое вам, ешьте без всякого исследования, для [спокойствия] совести.
1COR|10|28|Но если кто скажет вам: это идоложертвенное, – то не ешьте ради того, кто объявил вам, и ради совести. Ибо Господня земля, и что наполняет ее.
1COR|10|29|Совесть же разумею не свою, а другого: ибо для чего моей свободе быть судимой чужою совестью?
1COR|10|30|Если я с благодарением принимаю [пищу], то для чего порицать меня за то, за что я благодарю?
1COR|10|31|Итак, едите ли, пьете ли, или иное что делаете, все делайте в славу Божию.
1COR|10|32|Не подавайте соблазна ни Иудеям, ни Еллинам, ни церкви Божией,
1COR|10|33|так, как и я угождаю всем во всем, ища не своей пользы, но [пользы] многих, чтобы они спаслись.
1COR|11|1|Будьте подражателями мне, как я Христу.
1COR|11|2|Хвалю вас, братия, что вы все мое помните и держите предания так, как я передал вам.
1COR|11|3|Хочу также, чтобы вы знали, что всякому мужу глава Христос, жене глава – муж, а Христу глава – Бог.
1COR|11|4|Всякий муж, молящийся или пророчествующий с покрытою головою, постыжает свою голову.
1COR|11|5|И всякая жена, молящаяся или пророчествующая с открытою головою, постыжает свою голову, ибо [это] то же, как если бы она была обритая.
1COR|11|6|Ибо если жена не хочет покрываться, то пусть и стрижется; а если жене стыдно быть остриженной или обритой, пусть покрывается.
1COR|11|7|Итак муж не должен покрывать голову, потому что он есть образ и слава Божия; а жена есть слава мужа.
1COR|11|8|Ибо не муж от жены, но жена от мужа;
1COR|11|9|и не муж создан для жены, но жена для мужа.
1COR|11|10|Посему жена и должна иметь на голове своей [знак] власти [над] [нею], для Ангелов.
1COR|11|11|Впрочем ни муж без жены, ни жена без мужа, в Господе.
1COR|11|12|Ибо как жена от мужа, так и муж через жену; все же – от Бога.
1COR|11|13|Рассудите сами, прилично ли жене молиться Богу с непокрытою [головою]?
1COR|11|14|Не сама ли природа учит вас, что если муж растит волосы, то это бесчестье для него,
1COR|11|15|но если жена растит волосы, для нее это честь, так как волосы даны ей вместо покрывала?
1COR|11|16|А если бы кто захотел спорить, то мы не имеем такого обычая, ни церкви Божии.
1COR|11|17|Но, предлагая сие, не хвалю [вас], что вы собираетесь не на лучшее, а на худшее.
1COR|11|18|Ибо, во–первых, слышу, что, когда вы собираетесь в церковь, между вами бывают разделения, чему отчасти и верю.
1COR|11|19|Ибо надлежит быть и разномыслиям между вами, дабы открылись между вами искусные.
1COR|11|20|Далее, вы собираетесь, [так, что это] не значит вкушать вечерю Господню;
1COR|11|21|ибо всякий поспешает прежде [других] есть свою пищу, [так] [что] иной бывает голоден, а иной упивается.
1COR|11|22|Разве у вас нет домов на то, чтобы есть и пить? Или пренебрегаете церковь Божию и унижаете неимущих? Что сказать вам? похвалить ли вас за это? Не похвалю.
1COR|11|23|Ибо я от [Самого] Господа принял то, что и вам передал, что Господь Иисус в ту ночь, в которую предан был, взял хлеб
1COR|11|24|и, возблагодарив, преломил и сказал: приимите, ядите, сие есть Тело Мое, за вас ломимое; сие творите в Мое воспоминание.
1COR|11|25|Также и чашу после вечери, и сказал: сия чаша есть новый завет в Моей Крови; сие творите, когда только будете пить, в Мое воспоминание.
1COR|11|26|Ибо всякий раз, когда вы едите хлеб сей и пьете чашу сию, смерть Господню возвещаете, доколе Он придет.
1COR|11|27|Посему, кто будет есть хлеб сей или пить чашу Господню недостойно, виновен будет против Тела и Крови Господней.
1COR|11|28|Да испытывает же себя человек, и таким образом пусть ест от хлеба сего и пьет из чаши сей.
1COR|11|29|Ибо, кто ест и пьет недостойно, тот ест и пьет осуждение себе, не рассуждая о Теле Господнем.
1COR|11|30|От того многие из вас немощны и больны и немало умирает.
1COR|11|31|Ибо если бы мы судили сами себя, то не были бы судимы.
1COR|11|32|Будучи же судимы, наказываемся от Господа, чтобы не быть осужденными с миром.
1COR|11|33|Посему, братия мои, собираясь на вечерю, друг друга ждите.
1COR|11|34|А если кто голоден, пусть ест дома, чтобы собираться вам не на осуждение. Прочее устрою, когда приду.
1COR|12|1|Не хочу оставить вас, братия, в неведении и о [дарах] духовных.
1COR|12|2|Знаете, что когда вы были язычниками, то ходили к безгласным идолам, так, как бы вели вас.
1COR|12|3|Потому сказываю вам, что никто, говорящий Духом Божиим, не произнесет анафемы на Иисуса, и никто не может назвать Иисуса Господом, как только Духом Святым.
1COR|12|4|Дары различны, но Дух один и тот же;
1COR|12|5|и служения различны, а Господь один и тот же;
1COR|12|6|и действия различны, а Бог один и тот же, производящий все во всех.
1COR|12|7|Но каждому дается проявление Духа на пользу.
1COR|12|8|Одному дается Духом слово мудрости, другому слово знания, тем же Духом;
1COR|12|9|иному вера, тем же Духом; иному дары исцелений, тем же Духом;
1COR|12|10|иному чудотворения, иному пророчество, иному различение духов, иному разные языки, иному истолкование языков.
1COR|12|11|Все же сие производит один и тот же Дух, разделяя каждому особо, как Ему угодно.
1COR|12|12|Ибо, как тело одно, но имеет многие члены, и все члены одного тела, хотя их и много, составляют одно тело, – так и Христос.
1COR|12|13|Ибо все мы одним Духом крестились в одно тело, Иудеи или Еллины, рабы или свободные, и все напоены одним Духом.
1COR|12|14|Тело же не из одного члена, но из многих.
1COR|12|15|Если нога скажет: я не принадлежу к телу, потому что я не рука, то неужели она потому не принадлежит к телу?
1COR|12|16|И если ухо скажет: я не принадлежу к телу, потому что я не глаз, то неужели оно потому не принадлежит к телу?
1COR|12|17|Если все тело глаз, то где слух? Если все слух, то где обоняние?
1COR|12|18|Но Бог расположил члены, каждый в [составе] тела, как Ему было угодно.
1COR|12|19|А если бы все были один член, то где [было бы] тело?
1COR|12|20|Но теперь членов много, а тело одно.
1COR|12|21|Не может глаз сказать руке: ты мне не надобна; или также голова ногам: вы мне не нужны.
1COR|12|22|Напротив, члены тела, которые кажутся слабейшими, гораздо нужнее,
1COR|12|23|и которые нам кажутся менее благородными в теле, о тех более прилагаем попечения;
1COR|12|24|и неблагообразные наши более благовидно покрываются, а благообразные наши не имеют [в том] нужды. Но Бог соразмерил тело, внушив о менее совершенном большее попечение,
1COR|12|25|дабы не было разделения в теле, а все члены одинаково заботились друг о друге.
1COR|12|26|Посему, страдает ли один член, страдают с ним все члены; славится ли один член, с ним радуются все члены.
1COR|12|27|И вы – тело Христово, а порознь – члены.
1COR|12|28|И иных Бог поставил в Церкви, во–первых, Апостолами, во–вторых, пророками, в–третьих, учителями; далее, [иным дал] силы [чудодейственные], также дары исцелений, вспоможения, управления, разные языки.
1COR|12|29|Все ли Апостолы? Все ли пророки? Все ли учители? Все ли чудотворцы?
1COR|12|30|Все ли имеют дары исцелений? Все ли говорят языками? Все ли истолкователи?
1COR|12|31|Ревнуйте о дарах больших, и я покажу вам путь еще превосходнейший.
1COR|13|1|Если я говорю языками человеческими и ангельскими, а любви не имею, то я – медь звенящая или кимвал звучащий.
1COR|13|2|Если имею [дар] пророчества, и знаю все тайны, и имею всякое познание и всю веру, так что [могу] и горы переставлять, а не имею любви, – то я ничто.
1COR|13|3|И если я раздам все имение мое и отдам тело мое на сожжение, а любви не имею, нет мне в том никакой пользы.
1COR|13|4|Любовь долготерпит, милосердствует, любовь не завидует, любовь не превозносится, не гордится,
1COR|13|5|не бесчинствует, не ищет своего, не раздражается, не мыслит зла,
1COR|13|6|не радуется неправде, а сорадуется истине;
1COR|13|7|все покрывает, всему верит, всего надеется, все переносит.
1COR|13|8|Любовь никогда не перестает, хотя и пророчества прекратятся, и языки умолкнут, и знание упразднится.
1COR|13|9|Ибо мы отчасти знаем, и отчасти пророчествуем;
1COR|13|10|когда же настанет совершенное, тогда то, что отчасти, прекратится.
1COR|13|11|Когда я был младенцем, то по–младенчески говорил, по–младенчески мыслил, по–младенчески рассуждал; а как стал мужем, то оставил младенческое.
1COR|13|12|Теперь мы видим как бы сквозь [тусклое] стекло, гадательно, тогда же лицем к лицу; теперь знаю я отчасти, а тогда познаю, подобно как я познан.
1COR|13|13|А теперь пребывают сии три: вера, надежда, любовь; но любовь из них больше.
1COR|14|1|Достигайте любви; ревнуйте о [дарах] духовных, особенно же о том, чтобы пророчествовать.
1COR|14|2|Ибо кто говорит на [незнакомом] языке, тот говорит не людям, а Богу; потому что никто не понимает [его], он тайны говорит духом;
1COR|14|3|а кто пророчествует, тот говорит людям в назидание, увещание и утешение.
1COR|14|4|Кто говорит на [незнакомом] языке, тот назидает себя; а кто пророчествует, тот назидает церковь.
1COR|14|5|Желаю, чтобы вы все говорили языками; но лучше, чтобы вы пророчествовали; ибо пророчествующий превосходнее того, кто говорит языками, разве он притом будет и изъяснять, чтобы церковь получила назидание.
1COR|14|6|Теперь, если я приду к вам, братия, и стану говорить на [незнакомых] языках, то какую принесу вам пользу, когда не изъяснюсь вам или откровением, или познанием, или пророчеством, или учением?
1COR|14|7|И бездушные [вещи], издающие звук, свирель или гусли, если не производят раздельных тонов, как распознать то, что играют на свирели или на гуслях?
1COR|14|8|И если труба будет издавать неопределенный звук, кто станет готовиться к сражению?
1COR|14|9|Так если и вы языком произносите невразумительные слова, то как узнают, что вы говорите? Вы будете говорить на ветер.
1COR|14|10|Сколько, например, различных слов в мире, и ни одного из них нет без значения.
1COR|14|11|Но если я не разумею значения слов, то я для говорящего чужестранец, и говорящий для меня чужестранец.
1COR|14|12|Так и вы, ревнуя о [дарах] духовных, старайтесь обогатиться [ими] к назиданию церкви.
1COR|14|13|А потому, говорящий на [незнакомом] языке, молись о даре истолкования.
1COR|14|14|Ибо когда я молюсь на [незнакомом] языке, то хотя дух мой и молится, но ум мой остается без плода.
1COR|14|15|Что же делать? Стану молиться духом, стану молиться и умом; буду петь духом, буду петь и умом.
1COR|14|16|Ибо если ты будешь благословлять духом, то стоящий на месте простолюдина как скажет: "аминь" при твоем благодарении? Ибо он не понимает, что ты говоришь.
1COR|14|17|Ты хорошо благодаришь, но другой не назидается.
1COR|14|18|Благодарю Бога моего: я более всех вас говорю языками;
1COR|14|19|но в церкви хочу лучше пять слов сказать умом моим, чтобы и других наставить, нежели тьму слов на [незнакомом] языке.
1COR|14|20|Братия! не будьте дети умом: на злое будьте младенцы, а по уму будьте совершеннолетни.
1COR|14|21|В законе написано: иными языками и иными устами буду говорить народу сему; но и тогда не послушают Меня, говорит Господь.
1COR|14|22|Итак языки суть знамение не для верующих, а для неверующих; пророчество же не для неверующих, а для верующих.
1COR|14|23|Если вся церковь сойдется вместе, и все станут говорить [незнакомыми] языками, и войдут к вам незнающие или неверующие, то не скажут ли, что вы беснуетесь?
1COR|14|24|Но когда все пророчествуют, и войдет кто неверующий или незнающий, то он всеми обличается, всеми судится.
1COR|14|25|И таким образом тайны сердца его обнаруживаются, и он падет ниц, поклонится Богу и скажет: истинно с вами Бог.
1COR|14|26|Итак что же, братия? Когда вы сходитесь, и у каждого из вас есть псалом, есть поучение, есть язык, есть откровение, есть истолкование, – все сие да будет к назиданию.
1COR|14|27|Если кто говорит на [незнакомом] языке, [говорите] двое, или много трое, и то порознь, а один изъясняй.
1COR|14|28|Если же не будет истолкователя, то молчи в церкви, а говори себе и Богу.
1COR|14|29|И пророки пусть говорят двое или трое, а прочие пусть рассуждают.
1COR|14|30|Если же другому из сидящих будет откровение, то первый молчи.
1COR|14|31|Ибо все один за другим можете пророчествовать, чтобы всем поучаться и всем получать утешение.
1COR|14|32|И духи пророческие послушны пророкам,
1COR|14|33|потому что Бог не есть [Бог] неустройства, но мира. Так [бывает] во всех церквах у святых.
1COR|14|34|Жены ваши в церквах да молчат, ибо не позволено им говорить, а быть в подчинении, как и закон говорит.
1COR|14|35|Если же они хотят чему научиться, пусть спрашивают [о том] дома у мужей своих; ибо неприлично жене говорить в церкви.
1COR|14|36|Разве от вас вышло слово Божие? Или до вас одних достигло?
1COR|14|37|Если кто почитает себя пророком или духовным, тот да разумеет, что я пишу вам, ибо это заповеди Господни.
1COR|14|38|А кто не разумеет, пусть не разумеет.
1COR|14|39|Итак, братия, ревнуйте о том, чтобы пророчествовать, но не запрещайте говорить и языками;
1COR|14|40|только все должно быть благопристойно и чинно.
1COR|15|1|Напоминаю вам, братия, Евангелие, которое я благовествовал вам, которое вы и приняли, в котором и утвердились,
1COR|15|2|которым и спасаетесь, если преподанное удерживаете так, как я благовествовал вам, если только не тщетно уверовали.
1COR|15|3|Ибо я первоначально преподал вам, что и [сам] принял, [то] [есть], что Христос умер за грехи наши, по Писанию,
1COR|15|4|и что Он погребен был, и что воскрес в третий день, по Писанию,
1COR|15|5|и что явился Кифе, потом двенадцати;
1COR|15|6|потом явился более нежели пятистам братий в одно время, из которых большая часть доныне в живых, а некоторые и почили;
1COR|15|7|потом явился Иакову, также всем Апостолам;
1COR|15|8|а после всех явился и мне, как некоему извергу.
1COR|15|9|Ибо я наименьший из Апостолов, и недостоин называться Апостолом, потому что гнал церковь Божию.
1COR|15|10|Но благодатию Божиею есмь то, что есмь; и благодать Его во мне не была тщетна, но я более всех их потрудился: не я, впрочем, а благодать Божия, которая со мною.
1COR|15|11|Итак я ли, они ли, мы так проповедуем, и вы так уверовали.
1COR|15|12|Если же о Христе проповедуется, что Он воскрес из мертвых, то как некоторые из вас говорят, что нет воскресения мертвых?
1COR|15|13|Если нет воскресения мертвых, то и Христос не воскрес;
1COR|15|14|а если Христос не воскрес, то и проповедь наша тщетна, тщетна и вера ваша.
1COR|15|15|Притом мы оказались бы и лжесвидетелями о Боге, потому что свидетельствовали бы о Боге, что Он воскресил Христа, Которого Он не воскрешал, если, [то есть], мертвые не воскресают;
1COR|15|16|ибо если мертвые не воскресают, то и Христос не воскрес.
1COR|15|17|А если Христос не воскрес, то вера ваша тщетна: вы еще во грехах ваших.
1COR|15|18|Поэтому и умершие во Христе погибли.
1COR|15|19|И если мы в этой только жизни надеемся на Христа, то мы несчастнее всех человеков.
1COR|15|20|Но Христос воскрес из мертвых, первенец из умерших.
1COR|15|21|Ибо, как смерть через человека, [так] через человека и воскресение мертвых.
1COR|15|22|Как в Адаме все умирают, так во Христе все оживут,
1COR|15|23|каждый в своем порядке: первенец Христос, потом Христовы, в пришествие Его.
1COR|15|24|А затем конец, когда Он предаст Царство Богу и Отцу, когда упразднит всякое начальство и всякую власть и силу.
1COR|15|25|Ибо Ему надлежит царствовать, доколе низложит всех врагов под ноги Свои.
1COR|15|26|Последний же враг истребится – смерть,
1COR|15|27|потому что все покорил под ноги Его. Когда же сказано, что [Ему] все покорено, то ясно, что кроме Того, Который покорил Ему все.
1COR|15|28|Когда же все покорит Ему, тогда и Сам Сын покорится Покорившему все Ему, да будет Бог все во всем.
1COR|15|29|Иначе, что делают крестящиеся для мертвых? Если мертвые совсем не воскресают, то для чего и крестятся для мертвых?
1COR|15|30|Для чего и мы ежечасно подвергаемся бедствиям?
1COR|15|31|Я каждый день умираю: свидетельствуюсь в том похвалою вашею, братия, которую я имею во Христе Иисусе, Господе нашем.
1COR|15|32|По [рассуждению] человеческому, когда я боролся со зверями в Ефесе, какая мне польза, если мертвые не воскресают? Станем есть и пить, ибо завтра умрем!
1COR|15|33|Не обманывайтесь: худые сообщества развращают добрые нравы.
1COR|15|34|Отрезвитесь, как должно, и не грешите; ибо, к стыду вашему скажу, некоторые из вас не знают Бога.
1COR|15|35|Но скажет кто–нибудь: как воскреснут мертвые? и в каком теле придут?
1COR|15|36|Безрассудный! то, что ты сеешь, не оживет, если не умрет.
1COR|15|37|И когда ты сеешь, то сеешь не тело будущее, а голое зерно, какое случится, пшеничное или другое какое;
1COR|15|38|но Бог дает ему тело, как хочет, и каждому семени свое тело.
1COR|15|39|Не всякая плоть такая же плоть; но иная плоть у человеков, иная плоть у скотов, иная у рыб, иная у птиц.
1COR|15|40|Есть тела небесные и тела земные; но иная слава небесных, иная земных.
1COR|15|41|Иная слава солнца, иная слава луны, иная звезд; и звезда от звезды разнится в славе.
1COR|15|42|Так и при воскресении мертвых: сеется в тлении, восстает в нетлении;
1COR|15|43|сеется в уничижении, восстает в славе; сеется в немощи, восстает в силе;
1COR|15|44|сеется тело душевное, восстает тело духовное. Есть тело душевное, есть тело и духовное.
1COR|15|45|Так и написано: первый человек Адам стал душею живущею; а последний Адам есть дух животворящий.
1COR|15|46|Но не духовное прежде, а душевное, потом духовное.
1COR|15|47|Первый человек – из земли, перстный; второй человек – Господь с неба.
1COR|15|48|Каков перстный, таковы и перстные; и каков небесный, таковы и небесные.
1COR|15|49|И как мы носили образ перстного, будем носить и образ небесного.
1COR|15|50|Но то скажу [вам], братия, что плоть и кровь не могут наследовать Царствия Божия, и тление не наследует нетления.
1COR|15|51|Говорю вам тайну: не все мы умрем, но все изменимся
1COR|15|52|вдруг, во мгновение ока, при последней трубе; ибо вострубит, и мертвые воскреснут нетленными, а мы изменимся.
1COR|15|53|Ибо тленному сему надлежит облечься в нетление, и смертному сему облечься в бессмертие.
1COR|15|54|Когда же тленное сие облечется в нетление и смертное сие облечется в бессмертие, тогда сбудется слово написанное: поглощена смерть победою.
1COR|15|55|Смерть! где твое жало? ад! где твоя победа?
1COR|15|56|Жало же смерти – грех; а сила греха – закон.
1COR|15|57|Благодарение Богу, даровавшему нам победу Господом нашим Иисусом Христом!
1COR|15|58|Итак, братия мои возлюбленные, будьте тверды, непоколебимы, всегда преуспевайте в деле Господнем, зная, что труд ваш не тщетен пред Господом.
1COR|16|1|При сборе же для святых поступайте так, как я установил в церквах Галатийских.
1COR|16|2|В первый день недели каждый из вас пусть отлагает у себя и сберегает, сколько позволит ему состояние, чтобы не делать сборов, когда я приду.
1COR|16|3|Когда же приду, то, которых вы изберете, тех отправлю с письмами, для доставления вашего подаяния в Иерусалим.
1COR|16|4|А если прилично будет и мне отправиться, то они со мной пойдут.
1COR|16|5|Я приду к вам, когда пройду Македонию; ибо я иду через Македонию.
1COR|16|6|У вас же, может быть, поживу, или и перезимую, чтобы вы меня проводили, куда пойду.
1COR|16|7|Ибо я не хочу видеться с вами теперь мимоходом, а надеюсь пробыть у вас несколько времени, если Господь позволит.
1COR|16|8|В Ефесе же я пробуду до Пятидесятницы,
1COR|16|9|ибо для меня отверста великая и широкая дверь, и противников много.
1COR|16|10|Если же придет к вам Тимофей, смотрите, чтобы он был у вас безопасен; ибо он делает дело Господне, как и я.
1COR|16|11|Посему никто не пренебрегай его, но проводите его с миром, чтобы он пришел ко мне, ибо я жду его с братиями.
1COR|16|12|А что до брата Аполлоса, я очень просил его, чтобы он с братиями пошел к вам; но он никак не хотел идти ныне, а придет, когда ему будет удобно.
1COR|16|13|Бодрствуйте, стойте в вере, будьте мужественны, тверды.
1COR|16|14|Все у вас да будет с любовью.
1COR|16|15|Прошу вас, братия (вы знаете семейство Стефаново, что оно есть начаток Ахаии и что они посвятили себя на служение святым),
1COR|16|16|будьте и вы почтительны к таковым и ко всякому содействующему и трудящемуся.
1COR|16|17|Я рад прибытию Стефана, Фортуната и Ахаика: они восполнили для меня отсутствие ваше,
1COR|16|18|ибо они мой и ваш дух успокоили. Почитайте таковых.
1COR|16|19|Приветствуют вас церкви Асийские; приветствуют вас усердно в Господе Акила и Прискилла с домашнею их церковью.
1COR|16|20|Приветствуют вас все братия. Приветствуйте друг друга святым целованием.
1COR|16|21|Мое, Павлово, приветствие собственноручно.
1COR|16|22|Кто не любит Господа Иисуса Христа, анафема, маранафа.
1COR|16|23|Благодать Господа нашего Иисуса Христа с вами,
1COR|16|24|и любовь моя со всеми вами во Христе Иисусе. Аминь.
