2THESS|1|1|Павел и Силуан и Тимофей – Фессалоникской церкви в Боге Отце нашем и Господе Иисусе Христе:
2THESS|1|2|благодать вам и мир от Бога Отца нашего и Господа Иисуса Христа.
2THESS|1|3|Всегда по справедливости мы должны благодарить Бога за вас, братия, потому что возрастает вера ваша, и умножается любовь каждого друг ко другу между всеми вами,
2THESS|1|4|так что мы сами хвалимся вами в церквах Божиих, терпением вашим и верою во всех гонениях и скорбях, переносимых вами
2THESS|1|5|в доказательство того, что будет праведный суд Божий, чтобы вам удостоиться Царствия Божия, для которого и страдаете.
2THESS|1|6|Ибо праведно пред Богом – оскорбляющим вас воздать скорбью,
2THESS|1|7|а вам, оскорбляемым, отрадою вместе с нами, в явление Господа Иисуса с неба, с Ангелами силы Его,
2THESS|1|8|в пламенеющем огне совершающего отмщение не познавшим Бога и не покоряющимся благовествованию Господа нашего Иисуса Христа,
2THESS|1|9|которые подвергнутся наказанию, вечной погибели, от лица Господа и от славы могущества Его,
2THESS|1|10|когда Он приидет прославиться во святых Своих и явиться дивным в день оный во всех веровавших, так как вы поверили нашему свидетельству.
2THESS|1|11|Для сего и молимся всегда за вас, чтобы Бог наш соделал вас достойными звания и совершил всякое благоволение благости и дело веры в силе,
2THESS|1|12|да прославится имя Господа нашего Иисуса Христа в вас, и вы в Нем, по благодати Бога нашего и Господа Иисуса Христа.
2THESS|2|1|Молим вас, братия, о пришествии Господа нашего Иисуса Христа и нашем собрании к Нему,
2THESS|2|2|не спешить колебаться умом и смущаться ни от духа, ни от слова, ни от послания, как бы нами посланного, будто уже наступает день Христов.
2THESS|2|3|Да не обольстит вас никто никак: [ибо день тот не] [придет], доколе не придет прежде отступление и не откроется человек греха, сын погибели,
2THESS|2|4|противящийся и превозносящийся выше всего, называемого Богом или святынею, так что в храме Божием сядет он, как Бог, выдавая себя за Бога.
2THESS|2|5|Не помните ли, что я, еще находясь у вас, говорил вам это?
2THESS|2|6|И ныне вы знаете, что не допускает открыться ему в свое время.
2THESS|2|7|Ибо тайна беззакония уже в действии, только [не совершится] до тех пор, пока не будет взят от среды удерживающий теперь.
2THESS|2|8|И тогда откроется беззаконник, которого Господь Иисус убьет духом уст Своих и истребит явлением пришествия Своего
2THESS|2|9|того, которого пришествие, по действию сатаны, будет со всякою силою и знамениями и чудесами ложными,
2THESS|2|10|и со всяким неправедным обольщением погибающих за то, что они не приняли любви истины для своего спасения.
2THESS|2|11|И за сие пошлет им Бог действие заблуждения, так что они будут верить лжи,
2THESS|2|12|да будут осуждены все, не веровавшие истине, но возлюбившие неправду.
2THESS|2|13|Мы же всегда должны благодарить Бога за вас, возлюбленные Господом братия, что Бог от начала, через освящение Духа и веру истине, избрал вас ко спасению,
2THESS|2|14|к которому и призвал вас благовествованием нашим, для достижения славы Господа нашего Иисуса Христа.
2THESS|2|15|Итак, братия, стойте и держите предания, которым вы научены или словом или посланием нашим.
2THESS|2|16|Сам же Господь наш Иисус Христос и Бог и Отец наш, возлюбивший нас и давший утешение вечное и надежду благую во благодати,
2THESS|2|17|да утешит ваши сердца и да утвердит вас во всяком слове и деле благом.
2THESS|3|1|Итак молитесь за нас, братия, чтобы слово Господне распространялось и прославлялось, как и у вас,
2THESS|3|2|и чтобы нам избавиться от беспорядочных и лукавых людей, ибо не во всех вера.
2THESS|3|3|Но верен Господь, Который утвердит вас и сохранит от лукавого.
2THESS|3|4|Мы уверены о вас в Господе, что вы исполняете и будете исполнять то, что мы вам повелеваем.
2THESS|3|5|Господь же да управит сердца ваши в любовь Божию и в терпение Христово.
2THESS|3|6|Завещеваем же вам, братия, именем Господа нашего Иисуса Христа, удаляться от всякого брата, поступающего бесчинно, а не по преданию, которое приняли от нас,
2THESS|3|7|ибо вы сами знаете, как должны вы подражать нам; ибо мы не бесчинствовали у вас,
2THESS|3|8|ни у кого не ели хлеба даром, но занимались трудом и работою ночь и день, чтобы не обременить кого из вас, –
2THESS|3|9|не потому, чтобы мы не имели власти, но чтобы себя самих дать вам в образец для подражания нам.
2THESS|3|10|Ибо когда мы были у вас, то завещевали вам сие: если кто не хочет трудиться, тот и не ешь.
2THESS|3|11|Но слышим, что некоторые у вас поступают бесчинно, ничего не делают, а суетятся.
2THESS|3|12|Таковых увещеваем и убеждаем Господом нашим Иисусом Христом, чтобы они, работая в безмолвии, ели свой хлеб.
2THESS|3|13|Вы же, братия, не унывайте, делая добро.
2THESS|3|14|Если же кто не послушает слова нашего в сем послании, того имейте на замечании и не сообщайтесь с ним, чтобы устыдить его.
2THESS|3|15|Но не считайте его за врага, а вразумляйте, как брата.
2THESS|3|16|Сам же Господь мира да даст вам мир всегда во всем. Господь со всеми вами!
2THESS|3|17|Приветствие моею рукою, Павловою, что служит знаком во всяком послании; пишу я так:
2THESS|3|18|благодать Господа нашего Иисуса Христа со всеми вами. Аминь.
