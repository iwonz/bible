MARK|1|1|initium evangelii Iesu Christi Filii Dei
MARK|1|2|sicut scriptum est in Esaia propheta ecce mitto angelum meum ante faciem tuam qui praeparabit viam tuam
MARK|1|3|vox clamantis in deserto parate viam Domini rectas facite semitas eius
MARK|1|4|fuit Iohannes in deserto baptizans et praedicans baptismum paenitentiae in remissionem peccatorum
MARK|1|5|et egrediebatur ad illum omnis Iudaeae regio et Hierosolymitae universi et baptizabantur ab illo in Iordane flumine confitentes peccata sua
MARK|1|6|et erat Iohannes vestitus pilis cameli et zona pellicia circa lumbos eius et lucustas et mel silvestre edebat
MARK|1|7|et praedicabat dicens venit fortior me post me cuius non sum dignus procumbens solvere corrigiam calciamentorum eius
MARK|1|8|ego baptizavi vos aqua ille vero baptizabit vos Spiritu Sancto
MARK|1|9|et factum est in diebus illis venit Iesus a Nazareth Galilaeae et baptizatus est in Iordane ab Iohanne
MARK|1|10|et statim ascendens de aqua vidit apertos caelos et Spiritum tamquam columbam descendentem et manentem in ipso
MARK|1|11|et vox facta est de caelis tu es Filius meus dilectus in te conplacui
MARK|1|12|et statim Spiritus expellit eum in desertum
MARK|1|13|et erat in deserto quadraginta diebus et quadraginta noctibus et temptabatur a Satana eratque cum bestiis et angeli ministrabant illi
MARK|1|14|postquam autem traditus est Iohannes venit Iesus in Galilaeam praedicans evangelium regni Dei
MARK|1|15|et dicens quoniam impletum est tempus et adpropinquavit regnum Dei paenitemini et credite evangelio
MARK|1|16|et praeteriens secus mare Galilaeae vidit Simonem et Andream fratrem eius mittentes retia in mare erant enim piscatores
MARK|1|17|et dixit eis Iesus venite post me et faciam vos fieri piscatores hominum
MARK|1|18|et protinus relictis retibus secuti sunt eum
MARK|1|19|et progressus inde pusillum vidit Iacobum Zebedaei et Iohannem fratrem eius et ipsos in navi conponentes retia
MARK|1|20|et statim vocavit illos et relicto patre suo Zebedaeo in navi cum mercennariis secuti sunt eum
MARK|1|21|et ingrediuntur Capharnaum et statim sabbatis ingressus synagogam docebat eos
MARK|1|22|et stupebant super doctrina eius erat enim docens eos quasi potestatem habens et non sicut scribae
MARK|1|23|et erat in synagoga eorum homo in spiritu inmundo et exclamavit
MARK|1|24|dicens quid nobis et tibi Iesu Nazarene venisti perdere nos scio qui sis Sanctus Dei
MARK|1|25|et comminatus est ei Iesus dicens obmutesce et exi de homine
MARK|1|26|et discerpens eum spiritus inmundus et exclamans voce magna exivit ab eo
MARK|1|27|et mirati sunt omnes ita ut conquirerent inter se dicentes quidnam est hoc quae doctrina haec nova quia in potestate et spiritibus inmundis imperat et oboediunt ei
MARK|1|28|et processit rumor eius statim in omnem regionem Galilaeae
MARK|1|29|et protinus egredientes de synagoga venerunt in domum Simonis et Andreae cum Iacobo et Iohanne
MARK|1|30|decumbebat autem socrus Simonis febricitans et statim dicunt ei de illa
MARK|1|31|et accedens elevavit eam adprehensa manu eius et continuo dimisit eam febris et ministrabat eis
MARK|1|32|vespere autem facto cum occidisset sol adferebant ad eum omnes male habentes et daemonia habentes
MARK|1|33|et erat omnis civitas congregata ad ianuam
MARK|1|34|et curavit multos qui vexabantur variis languoribus et daemonia multa eiciebat et non sinebat loqui ea quoniam sciebant eum
MARK|1|35|et diluculo valde surgens egressus abiit in desertum locum ibique orabat
MARK|1|36|et persecutus est eum Simon et qui cum illo erant
MARK|1|37|et cum invenissent eum dixerunt ei quia omnes quaerunt te
MARK|1|38|et ait illis eamus in proximos vicos et civitates ut et ibi praedicem ad hoc enim veni
MARK|1|39|et erat praedicans in synagogis eorum et omni Galilaea et daemonia eiciens
MARK|1|40|et venit ad eum leprosus deprecans eum et genu flexo dixit si vis potes me mundare
MARK|1|41|Iesus autem misertus eius extendit manum suam et tangens eum ait illi volo mundare
MARK|1|42|et cum dixisset statim discessit ab eo lepra et mundatus est
MARK|1|43|et comminatus ei statim eiecit illum
MARK|1|44|et dicit ei vide nemini dixeris sed vade ostende te principi sacerdotum et offer pro emundatione tua quae praecepit Moses in testimonium illis
MARK|1|45|at ille egressus coepit praedicare et diffamare sermonem ita ut iam non posset manifeste in civitatem introire sed foris in desertis locis esse et conveniebant ad eum undique
MARK|2|1|et iterum intravit Capharnaum post dies
MARK|2|2|et auditum est quod in domo esset et convenerunt multi ita ut non caperet neque ad ianuam et loquebatur eis verbum
MARK|2|3|et venerunt ferentes ad eum paralyticum qui a quattuor portabatur
MARK|2|4|et cum non possent offerre eum illi prae turba nudaverunt tectum ubi erat et patefacientes submiserunt grabattum in quo paralyticus iacebat
MARK|2|5|cum vidisset autem Iesus fidem illorum ait paralytico fili dimittuntur tibi peccata
MARK|2|6|erant autem illic quidam de scribis sedentes et cogitantes in cordibus suis
MARK|2|7|quid hic sic loquitur blasphemat quis potest dimittere peccata nisi solus Deus
MARK|2|8|quo statim cognito Iesus spiritu suo quia sic cogitarent intra se dicit illis quid ista cogitatis in cordibus vestris
MARK|2|9|quid est facilius dicere paralytico dimittuntur tibi peccata an dicere surge et tolle grabattum tuum et ambula
MARK|2|10|ut autem sciatis quia potestatem habet Filius hominis in terra dimittendi peccata ait paralytico
MARK|2|11|tibi dico surge tolle grabattum tuum et vade in domum tuam
MARK|2|12|et statim ille surrexit et sublato grabatto abiit coram omnibus ita ut admirarentur omnes et honorificarent Deum dicentes quia numquam sic vidimus
MARK|2|13|et egressus est rursus ad mare omnisque turba veniebat ad eum et docebat eos
MARK|2|14|et cum praeteriret vidit Levin Alphei sedentem ad teloneum et ait illi sequere me et surgens secutus est eum
MARK|2|15|et factum est cum accumberet in domo illius multi publicani et peccatores simul discumbebant cum Iesu et discipulis eius erant enim multi qui et sequebantur eum
MARK|2|16|et scribae et Pharisaei videntes quia manducaret cum peccatoribus et publicanis dicebant discipulis eius quare cum publicanis et peccatoribus manducat et bibit magister vester
MARK|2|17|hoc audito Iesus ait illis non necesse habent sani medicum sed qui male habent non enim veni vocare iustos sed peccatores
MARK|2|18|et erant discipuli Iohannis et Pharisaei ieiunantes et veniunt et dicunt illi cur discipuli Iohannis et Pharisaeorum ieiunant tui autem discipuli non ieiunant
MARK|2|19|et ait illis Iesus numquid possunt filii nuptiarum quamdiu sponsus cum illis est ieiunare quanto tempore habent secum sponsum non possunt ieiunare
MARK|2|20|venient autem dies cum auferetur ab eis sponsus et tunc ieiunabunt in illa die
MARK|2|21|nemo adsumentum panni rudis adsuit vestimento veteri alioquin aufert supplementum novum a veteri et maior scissura fit
MARK|2|22|et nemo mittit vinum novellum in utres veteres alioquin disrumpet vinum utres et vinum effunditur et utres peribunt sed vinum novum in utres novos mitti debet
MARK|2|23|et factum est iterum cum sabbatis ambularet per sata et discipuli eius coeperunt praegredi et vellere spicas
MARK|2|24|Pharisaei autem dicebant ei ecce quid faciunt sabbatis quod non licet
MARK|2|25|et ait illis numquam legistis quid fecerit David quando necessitatem habuit et esuriit ipse et qui cum eo erant
MARK|2|26|quomodo introiit in domum Dei sub Abiathar principe sacerdotum et panes propositionis manducavit quos non licet manducare nisi sacerdotibus et dedit eis qui cum eo erant
MARK|2|27|et dicebat eis sabbatum propter hominem factum est et non homo propter sabbatum
MARK|2|28|itaque dominus est Filius hominis etiam sabbati
MARK|3|1|et introivit iterum synagogam et erat ibi homo habens manum aridam
MARK|3|2|et observabant eum si sabbatis curaret ut accusarent illum
MARK|3|3|et ait homini habenti manum aridam surge in medium
MARK|3|4|et dicit eis licet sabbatis bene facere an male animam salvam facere an perdere at illi tacebant
MARK|3|5|et circumspiciens eos cum ira contristatus super caecitatem cordis eorum dicit homini extende manum tuam et extendit et restituta est manus illi
MARK|3|6|exeuntes autem statim Pharisaei cum Herodianis consilium faciebant adversus eum quomodo eum perderent
MARK|3|7|et Iesus cum discipulis suis secessit ad mare et multa turba a Galilaea et Iudaea secuta est eum
MARK|3|8|et ab Hierosolymis et ab Idumea et trans Iordanen et qui circa Tyrum et Sidonem multitudo magna audientes quae faciebat venerunt ad eum
MARK|3|9|et dixit discipulis suis ut navicula sibi deserviret propter turbam ne conprimerent eum
MARK|3|10|multos enim sanabat ita ut inruerent in eum ut illum tangerent quotquot habebant plagas
MARK|3|11|et spiritus inmundi cum illum videbant procidebant ei et clamabant dicentes
MARK|3|12|tu es Filius Dei et vehementer comminabatur eis ne manifestarent illum
MARK|3|13|et ascendens in montem vocavit ad se quos voluit ipse et venerunt ad eum
MARK|3|14|et fecit ut essent duodecim cum illo et ut mitteret eos praedicare
MARK|3|15|et dedit illis potestatem curandi infirmitates et eiciendi daemonia
MARK|3|16|et inposuit Simoni nomen Petrus
MARK|3|17|et Iacobum Zebedaei et Iohannem fratrem Iacobi et inposuit eis nomina Boanerges quod est Filii tonitrui
MARK|3|18|et Andream et Philippum et Bartholomeum et Mattheum et Thomam et Iacobum Alphei et Thaddeum et Simonem Cananeum
MARK|3|19|et Iudam Scarioth qui et tradidit illum
MARK|3|20|et veniunt ad domum et convenit iterum turba ita ut non possent neque panem manducare
MARK|3|21|et cum audissent sui exierunt tenere eum dicebant enim quoniam in furorem versus est
MARK|3|22|et scribae qui ab Hierosolymis descenderant dicebant quoniam Beelzebub habet et quia in principe daemonum eicit daemonia
MARK|3|23|et convocatis eis in parabolis dicebat illis quomodo potest Satanas Satanan eicere
MARK|3|24|et si regnum in se dividatur non potest stare regnum illud
MARK|3|25|et si domus super semet ipsam dispertiatur non poterit domus illa stare
MARK|3|26|et si Satanas consurrexit in semet ipsum dispertitus est et non potest stare sed finem habet
MARK|3|27|nemo potest vasa fortis ingressus in domum diripere nisi prius fortem alliget et tunc domum eius diripiet
MARK|3|28|amen dico vobis quoniam omnia dimittentur filiis hominum peccata et blasphemiae quibus blasphemaverint
MARK|3|29|qui autem blasphemaverit in Spiritum Sanctum non habet remissionem in aeternum sed reus erit aeterni delicti
MARK|3|30|quoniam dicebant spiritum inmundum habet
MARK|3|31|et veniunt mater eius et fratres et foris stantes miserunt ad eum vocantes eum
MARK|3|32|et sedebat circa eum turba et dicunt ei ecce mater tua et fratres tui foris quaerunt te
MARK|3|33|et respondens eis ait quae est mater mea et fratres mei
MARK|3|34|et circumspiciens eos qui in circuitu eius sedebant ait ecce mater mea et fratres mei
MARK|3|35|qui enim fecerit voluntatem Dei hic frater meus et soror mea et mater est
MARK|4|1|et iterum coepit docere ad mare et congregata est ad eum turba multa ita ut in navem ascendens sederet in mari et omnis turba circa mare super terram erat
MARK|4|2|et docebat eos in parabolis multa et dicebat illis in doctrina sua
MARK|4|3|audite ecce exiit seminans ad seminandum
MARK|4|4|et dum seminat aliud cecidit circa viam et venerunt volucres et comederunt illud
MARK|4|5|aliud vero cecidit super petrosa ubi non habuit terram multam et statim exortum est quoniam non habebat altitudinem terrae
MARK|4|6|et quando exortus est sol exaestuavit et eo quod non haberet radicem exaruit
MARK|4|7|et aliud cecidit in spinas et ascenderunt spinae et offocaverunt illud et fructum non dedit
MARK|4|8|et aliud cecidit in terram bonam et dabat fructum ascendentem et crescentem et adferebat unum triginta et unum sexaginta et unum centum
MARK|4|9|et dicebat qui habet aures audiendi audiat
MARK|4|10|et cum esset singularis interrogaverunt eum hii qui cum eo erant cum duodecim parabolas
MARK|4|11|et dicebat eis vobis datum est mysterium regni Dei illis autem qui foris sunt in parabolis omnia fiunt
MARK|4|12|ut videntes videant et non videant et audientes audiant et non intellegant nequando convertantur et dimittantur eis peccata
MARK|4|13|et ait illis nescitis parabolam hanc et quomodo omnes parabolas cognoscetis
MARK|4|14|qui seminat verbum seminat
MARK|4|15|hii autem sunt qui circa viam ubi seminatur verbum et cum audierint confestim venit Satanas et aufert verbum quod seminatum est in corda eorum
MARK|4|16|et hii sunt similiter qui super petrosa seminantur qui cum audierint verbum statim cum gaudio accipiunt illud
MARK|4|17|et non habent radicem in se sed temporales sunt deinde orta tribulatione et persecutione propter verbum confestim scandalizantur
MARK|4|18|et alii sunt qui in spinis seminantur hii sunt qui verbum audiunt
MARK|4|19|et aerumnae saeculi et deceptio divitiarum et circa reliqua concupiscentiae introeuntes suffocant verbum et sine fructu efficitur
MARK|4|20|et hii sunt qui super terram bonam seminati sunt qui audiunt verbum et suscipiunt et fructificant unum triginta et unum sexaginta et unum centum
MARK|4|21|et dicebat illis numquid venit lucerna ut sub modio ponatur aut sub lecto nonne ut super candelabrum ponatur
MARK|4|22|non enim est aliquid absconditum quod non manifestetur nec factum est occultum sed ut in palam veniat
MARK|4|23|si quis habet aures audiendi audiat
MARK|4|24|et dicebat illis videte quid audiatis in qua mensura mensi fueritis remetietur vobis et adicietur vobis
MARK|4|25|qui enim habet dabitur illi et qui non habet etiam quod habet auferetur ab illo
MARK|4|26|et dicebat sic est regnum Dei quemadmodum si homo iaciat sementem in terram
MARK|4|27|et dormiat et exsurgat nocte ac die et semen germinet et increscat dum nescit ille
MARK|4|28|ultro enim terra fructificat primum herbam deinde spicam deinde plenum frumentum in spica
MARK|4|29|et cum se produxerit fructus statim mittit falcem quoniam adest messis
MARK|4|30|et dicebat cui adsimilabimus regnum Dei aut cui parabolae conparabimus illud
MARK|4|31|sicut granum sinapis quod cum seminatum fuerit in terra minus est omnibus seminibus quae sunt in terra
MARK|4|32|et cum seminatum fuerit ascendit et fit maius omnibus holeribus et facit ramos magnos ita ut possint sub umbra eius aves caeli habitare
MARK|4|33|et talibus multis parabolis loquebatur eis verbum prout poterant audire
MARK|4|34|sine parabola autem non loquebatur eis seorsum autem discipulis suis disserebat omnia
MARK|4|35|et ait illis illa die cum sero esset factum transeamus contra
MARK|4|36|et dimittentes turbam adsumunt eum ita ut erat in navi et aliae naves erant cum illo
MARK|4|37|et facta est procella magna venti et fluctus mittebat in navem ita ut impleretur navis
MARK|4|38|et erat ipse in puppi supra cervical dormiens et excitant eum et dicunt ei magister non ad te pertinet quia perimus
MARK|4|39|et exsurgens comminatus est vento et dixit mari tace obmutesce et cessavit ventus et facta est tranquillitas magna
MARK|4|40|et ait illis quid timidi estis necdum habetis fidem et timuerunt magno timore et dicebant ad alterutrum quis putas est iste quia et ventus et mare oboediunt ei
MARK|5|1|et venerunt trans fretum maris in regionem Gerasenorum
MARK|5|2|et exeunti ei de navi statim occurrit ei de monumentis homo in spiritu inmundo
MARK|5|3|qui domicilium habebat in monumentis et neque catenis iam quisquam eum poterat ligare
MARK|5|4|quoniam saepe conpedibus et catenis vinctus disrupisset catenas et conpedes comminuisset et nemo poterat eum domare
MARK|5|5|et semper nocte ac die in monumentis et in montibus erat clamans et concidens se lapidibus
MARK|5|6|videns autem Iesum a longe cucurrit et adoravit eum
MARK|5|7|et clamans voce magna dicit quid mihi et tibi Iesu Fili Dei summi adiuro te per Deum ne me torqueas
MARK|5|8|dicebat enim illi exi spiritus inmunde ab homine
MARK|5|9|et interrogabat eum quod tibi nomen est et dicit ei Legio nomen mihi est quia multi sumus
MARK|5|10|et deprecabatur eum multum ne se expelleret extra regionem
MARK|5|11|erat autem ibi circa montem grex porcorum magnus pascens
MARK|5|12|et deprecabantur eum spiritus dicentes mitte nos in porcos ut in eos introeamus
MARK|5|13|et concessit eis statim Iesus et exeuntes spiritus inmundi introierunt in porcos et magno impetu grex praecipitatus est in mare ad duo milia et suffocati sunt in mare
MARK|5|14|qui autem pascebant eos fugerunt et nuntiaverunt in civitatem et in agros et egressi sunt videre quid esset facti
MARK|5|15|et veniunt ad Iesum et vident illum qui a daemonio vexabatur sedentem vestitum et sanae mentis et timuerunt
MARK|5|16|et narraverunt illis qui viderant qualiter factum esset ei qui daemonium habuerat et de porcis
MARK|5|17|et rogare eum coeperunt ut discederet de finibus eorum
MARK|5|18|cumque ascenderet navem coepit illum deprecari qui daemonio vexatus fuerat ut esset cum illo
MARK|5|19|et non admisit eum sed ait illi vade in domum tuam ad tuos et adnuntia illis quanta tibi Dominus fecerit et misertus sit tui
MARK|5|20|et abiit et coepit praedicare in Decapoli quanta sibi fecisset Iesus et omnes mirabantur
MARK|5|21|et cum transcendisset Iesus in navi rursus trans fretum convenit turba multa ad illum et erat circa mare
MARK|5|22|et venit quidam de archisynagogis nomine Iairus et videns eum procidit ad pedes eius
MARK|5|23|et deprecabatur eum multum dicens quoniam filia mea in extremis est veni inpone manus super eam ut salva sit et vivat
MARK|5|24|et abiit cum illo et sequebatur eum turba multa et conprimebant illum
MARK|5|25|et mulier quae erat in profluvio sanguinis annis duodecim
MARK|5|26|et fuerat multa perpessa a conpluribus medicis et erogaverat omnia sua nec quicquam profecerat sed magis deterius habebat
MARK|5|27|cum audisset de Iesu venit in turba retro et tetigit vestimentum eius
MARK|5|28|dicebat enim quia si vel vestimentum eius tetigero salva ero
MARK|5|29|et confestim siccatus est fons sanguinis eius et sensit corpore quod sanata esset a plaga
MARK|5|30|et statim Iesus cognoscens in semet ipso virtutem quae exierat de eo conversus ad turbam aiebat quis tetigit vestimenta mea
MARK|5|31|et dicebant ei discipuli sui vides turbam conprimentem te et dicis quis me tetigit
MARK|5|32|et circumspiciebat videre eam quae hoc fecerat
MARK|5|33|mulier autem timens et tremens sciens quod factum esset in se venit et procidit ante eum et dixit ei omnem veritatem
MARK|5|34|ille autem dixit ei filia fides tua te salvam fecit vade in pace et esto sana a plaga tua
MARK|5|35|adhuc eo loquente veniunt ab archisynagogo dicentes quia filia tua mortua est quid ultra vexas magistrum
MARK|5|36|Iesus autem verbo quod dicebatur audito ait archisynagogo noli timere tantummodo crede
MARK|5|37|et non admisit quemquam sequi se nisi Petrum et Iacobum et Iohannem fratrem Iacobi
MARK|5|38|et veniunt in domum archisynagogi et videt tumultum et flentes et heiulantes multum
MARK|5|39|et ingressus ait eis quid turbamini et ploratis puella non est mortua sed dormit
MARK|5|40|et inridebant eum ipse vero eiectis omnibus adsumit patrem et matrem puellae et qui secum erant et ingreditur ubi erat puella iacens
MARK|5|41|et tenens manum puellae ait illi talitha cumi quod est interpretatum puella tibi dico surge
MARK|5|42|et confestim surrexit puella et ambulabat erat autem annorum duodecim et obstipuerunt stupore maximo
MARK|5|43|et praecepit illis vehementer ut nemo id sciret et dixit dari illi manducare
MARK|6|1|et egressus inde abiit in patriam suam et sequebantur illum discipuli sui
MARK|6|2|et facto sabbato coepit in synagoga docere et multi audientes admirabantur in doctrina eius dicentes unde huic haec omnia et quae est sapientia quae data est illi et virtutes tales quae per manus eius efficiuntur
MARK|6|3|nonne iste est faber filius Mariae frater Iacobi et Ioseph et Iudae et Simonis nonne et sorores eius hic nobiscum sunt et scandalizabantur in illo
MARK|6|4|et dicebat eis Iesus quia non est propheta sine honore nisi in patria sua et in cognatione sua et in domo sua
MARK|6|5|et non poterat ibi virtutem ullam facere nisi paucos infirmos inpositis manibus curavit
MARK|6|6|et mirabatur propter incredulitatem eorum
MARK|6|7|et circumibat castella in circuitu docens et convocavit duodecim et coepit eos mittere binos et dabat illis potestatem spirituum inmundorum
MARK|6|8|et praecepit eis ne quid tollerent in via nisi virgam tantum non peram non panem neque in zona aes
MARK|6|9|sed calciatos sandaliis et ne induerentur duabus tunicis
MARK|6|10|et dicebat eis quocumque introieritis in domum illic manete donec exeatis inde
MARK|6|11|et quicumque non receperint vos nec audierint vos exeuntes inde excutite pulverem de pedibus vestris in testimonium illis
MARK|6|12|et exeuntes praedicabant ut paenitentiam agerent
MARK|6|13|et daemonia multa eiciebant et unguebant oleo multos aegrotos et sanabant
MARK|6|14|et audivit Herodes rex manifestum enim factum est nomen eius et dicebat quia Iohannes Baptista resurrexit a mortuis et propterea inoperantur virtutes in illo
MARK|6|15|alii autem dicebant quia Helias est alii vero dicebant propheta est quasi unus ex prophetis
MARK|6|16|quo audito Herodes ait quem ego decollavi Iohannem hic a mortuis resurrexit
MARK|6|17|ipse enim Herodes misit ac tenuit Iohannem et vinxit eum in carcere propter Herodiadem uxorem Philippi fratris sui quia duxerat eam
MARK|6|18|dicebat enim Iohannes Herodi non licet tibi habere uxorem fratris tui
MARK|6|19|Herodias autem insidiabatur illi et volebat occidere eum nec poterat
MARK|6|20|Herodes enim metuebat Iohannem sciens eum virum iustum et sanctum et custodiebat eum et audito eo multa faciebat et libenter eum audiebat
MARK|6|21|et cum dies oportunus accidisset Herodes natalis sui cenam fecit principibus et tribunis et primis Galilaeae
MARK|6|22|cumque introisset filia ipsius Herodiadis et saltasset et placuisset Herodi simulque recumbentibus rex ait puellae pete a me quod vis et dabo tibi
MARK|6|23|et iuravit illi quia quicquid petieris dabo tibi licet dimidium regni mei
MARK|6|24|quae cum exisset dixit matri suae quid petam et illa dixit caput Iohannis Baptistae
MARK|6|25|cumque introisset statim cum festinatione ad regem petivit dicens volo ut protinus des mihi in disco caput Iohannis Baptistae
MARK|6|26|et contristatus rex propter iusiurandum et propter simul recumbentes noluit eam contristare
MARK|6|27|sed misso speculatore praecepit adferri caput eius in disco et decollavit eum in carcere
MARK|6|28|et adtulit caput eius in disco et dedit illud puellae et puella dedit matri suae
MARK|6|29|quo audito discipuli eius venerunt et tulerunt corpus eius et posuerunt illud in monumento
MARK|6|30|et convenientes apostoli ad Iesum renuntiaverunt illi omnia quae egerant et docuerant
MARK|6|31|et ait illis venite seorsum in desertum locum et requiescite pusillum erant enim qui veniebant et rediebant multi et nec manducandi spatium habebant
MARK|6|32|et ascendentes in navi abierunt in desertum locum seorsum
MARK|6|33|et viderunt eos abeuntes et cognoverunt multi et pedestre et de omnibus civitatibus concurrerunt illuc et praevenerunt eos
MARK|6|34|et exiens vidit multam turbam Iesus et misertus est super eos quia erant sicut oves non habentes pastorem et coepit docere illos multa
MARK|6|35|et cum iam hora multa fieret accesserunt discipuli eius dicentes desertus est locus hic et iam hora praeterivit
MARK|6|36|dimitte illos ut euntes in proximas villas et vicos emant sibi cibos quos manducent
MARK|6|37|et respondens ait illis date illis manducare et dixerunt ei euntes emamus denariis ducentis panes et dabimus eis manducare
MARK|6|38|et dicit eis quot panes habetis ite et videte et cum cognovissent dicunt quinque et duos pisces
MARK|6|39|et praecepit illis ut accumbere facerent omnes secundum contubernia super viride faenum
MARK|6|40|et discubuerunt in partes per centenos et per quinquagenos
MARK|6|41|et acceptis quinque panibus et duobus piscibus intuens in caelum benedixit et fregit panes et dedit discipulis suis ut ponerent ante eos et duos pisces divisit omnibus
MARK|6|42|et manducaverunt omnes et saturati sunt
MARK|6|43|et sustulerunt reliquias fragmentorum duodecim cofinos plenos et de piscibus
MARK|6|44|erant autem qui manducaverunt quinque milia virorum
MARK|6|45|et statim coegit discipulos suos ascendere navem ut praecederent eum trans fretum ad Bethsaidam dum ipse dimitteret populum
MARK|6|46|et cum dimisisset eos abiit in montem orare
MARK|6|47|et cum sero esset erat navis in medio mari et ipse solus in terra
MARK|6|48|et videns eos laborantes in remigando erat enim ventus contrarius eis et circa quartam vigiliam noctis venit ad eos ambulans super mare et volebat praeterire eos
MARK|6|49|at illi ut viderunt eum ambulantem super mare putaverunt fantasma esse et exclamaverunt
MARK|6|50|omnes enim eum viderunt et conturbati sunt et statim locutus est cum eis et dixit illis confidite ego sum nolite timere
MARK|6|51|et ascendit ad illos in navem et cessavit ventus et plus magis intra se stupebant
MARK|6|52|non enim intellexerant de panibus erat enim cor illorum obcaecatum
MARK|6|53|et cum transfretassent pervenerunt in terram Gennesareth et adplicuerunt
MARK|6|54|cumque egressi essent de navi continuo cognoverunt eum
MARK|6|55|et percurrentes universam regionem illam coeperunt in grabattis eos qui se male habebant circumferre ubi audiebant eum esse
MARK|6|56|et quocumque introibat in vicos vel in villas aut civitates in plateis ponebant infirmos et deprecabantur eum ut vel fimbriam vestimenti eius tangerent et quotquot tangebant eum salvi fiebant
MARK|7|1|et conveniunt ad eum Pharisaei et quidam de scribis venientes ab Hierosolymis
MARK|7|2|et cum vidissent quosdam ex discipulis eius communibus manibus id est non lotis manducare panes vituperaverunt
MARK|7|3|Pharisaei enim et omnes Iudaei nisi crebro lavent manus non manducant tenentes traditionem seniorum
MARK|7|4|et a foro nisi baptizentur non comedunt et alia multa sunt quae tradita sunt illis servare baptismata calicum et urceorum et aeramentorum et lectorum
MARK|7|5|et interrogant eum Pharisaei et scribae quare discipuli tui non ambulant iuxta traditionem seniorum sed communibus manibus manducant panem
MARK|7|6|at ille respondens dixit eis bene prophetavit Esaias de vobis hypocritis sicut scriptum est populus hic labiis me honorat cor autem eorum longe est a me
MARK|7|7|in vanum autem me colunt docentes doctrinas praecepta hominum
MARK|7|8|relinquentes enim mandatum Dei tenetis traditionem hominum baptismata urceorum et calicum et alia similia his facitis multa
MARK|7|9|et dicebat illis bene irritum facitis praeceptum Dei ut traditionem vestram servetis
MARK|7|10|Moses enim dixit honora patrem tuum et matrem tuam et qui maledixerit patri aut matri morte moriatur
MARK|7|11|vos autem dicitis si dixerit homo patri aut matri corban quod est donum quodcumque ex me tibi profuerit
MARK|7|12|et ultra non dimittitis eum quicquam facere patri suo aut matri
MARK|7|13|rescindentes verbum Dei per traditionem vestram quam tradidistis et similia huiusmodi multa facitis
MARK|7|14|et advocans iterum turbam dicebat illis audite me omnes et intellegite
MARK|7|15|nihil est extra hominem introiens in eum quod possit eum coinquinare sed quae de homine procedunt illa sunt quae communicant hominem
MARK|7|16|si quis habet aures audiendi audiat
MARK|7|17|et cum introisset in domum a turba interrogabant eum discipuli eius parabolam
MARK|7|18|et ait illis sic et vos inprudentes estis non intellegitis quia omne extrinsecus introiens in hominem non potest eum communicare
MARK|7|19|quia non introit in cor eius sed in ventrem et in secessum exit purgans omnes escas
MARK|7|20|dicebat autem quoniam quae de homine exeunt illa communicant hominem
MARK|7|21|ab intus enim de corde hominum cogitationes malae procedunt adulteria fornicationes homicidia
MARK|7|22|furta avaritiae nequitiae dolus inpudicitia oculus malus blasphemia superbia stultitia
MARK|7|23|omnia haec mala ab intus procedunt et communicant hominem
MARK|7|24|et inde surgens abiit in fines Tyri et Sidonis et ingressus domum neminem voluit scire et non potuit latere
MARK|7|25|mulier enim statim ut audivit de eo cuius habebat filia spiritum inmundum intravit et procidit ad pedes eius
MARK|7|26|erat autem mulier gentilis Syrophoenissa genere et rogabat eum ut daemonium eiceret de filia eius
MARK|7|27|qui dixit illi sine prius saturari filios non est enim bonum sumere panem filiorum et mittere canibus
MARK|7|28|at illa respondit et dicit ei utique Domine nam et catelli sub mensa comedunt de micis puerorum
MARK|7|29|et ait illi propter hunc sermonem vade exiit daemonium de filia tua
MARK|7|30|et cum abisset domum suam invenit puellam iacentem supra lectum et daemonium exisse
MARK|7|31|et iterum exiens de finibus Tyri venit per Sidonem ad mare Galilaeae inter medios fines Decapoleos
MARK|7|32|et adducunt ei surdum et mutum et deprecantur eum ut inponat illi manum
MARK|7|33|et adprehendens eum de turba seorsum misit digitos suos in auriculas et expuens tetigit linguam eius
MARK|7|34|et suspiciens in caelum ingemuit et ait illi eppheta quod est adaperire
MARK|7|35|et statim apertae sunt aures eius et solutum est vinculum linguae eius et loquebatur recte
MARK|7|36|et praecepit illis ne cui dicerent quanto autem eis praecipiebat tanto magis plus praedicabant
MARK|7|37|et eo amplius admirabantur dicentes bene omnia fecit et surdos facit audire et mutos loqui
MARK|8|1|in illis diebus iterum cum turba multa esset nec haberent quod manducarent convocatis discipulis ait illis
MARK|8|2|misereor super turba quia ecce iam triduo sustinent me nec habent quod manducent
MARK|8|3|et si dimisero eos ieiunos in domum suam deficient in via quidam enim ex eis de longe venerunt
MARK|8|4|et responderunt ei discipuli sui unde istos poterit quis hic saturare panibus in solitudine
MARK|8|5|et interrogavit eos quot panes habetis qui dixerunt septem
MARK|8|6|et praecepit turbae discumbere supra terram et accipiens septem panes gratias agens fregit et dabat discipulis suis ut adponerent et adposuerunt turbae
MARK|8|7|et habebant pisciculos paucos et ipsos benedixit et iussit adponi
MARK|8|8|et manducaverunt et saturati sunt et sustulerunt quod superaverat de fragmentis septem sportas
MARK|8|9|erant autem qui manducaverunt quasi quattuor milia et dimisit eos
MARK|8|10|et statim ascendens navem cum discipulis suis venit in partes Dalmanutha
MARK|8|11|et exierunt Pharisaei et coeperunt conquirere cum eo quaerentes ab illo signum de caelo temptantes eum
MARK|8|12|et ingemescens spiritu ait quid generatio ista quaerit signum amen dico vobis si dabitur generationi isti signum
MARK|8|13|et dimittens eos ascendens iterum abiit trans fretum
MARK|8|14|et obliti sunt sumere panes et nisi unum panem non habebant secum in navi
MARK|8|15|et praecipiebat eis dicens videte cavete a fermento Pharisaeorum et fermento Herodis
MARK|8|16|et cogitabant ad alterutrum dicentes quia panes non habemus
MARK|8|17|quo cognito Iesus ait illis quid cogitatis quia panes non habetis nondum cognoscitis nec intellegitis adhuc caecatum habetis cor vestrum
MARK|8|18|oculos habentes non videtis et aures habentes non auditis nec recordamini
MARK|8|19|quando quinque panes fregi in quinque milia et quot cofinos fragmentorum plenos sustulistis dicunt ei duodecim
MARK|8|20|quando et septem panes in quattuor milia quot sportas fragmentorum tulistis et dicunt ei septem
MARK|8|21|et dicebat eis quomodo nondum intellegitis
MARK|8|22|et veniunt Bethsaida et adducunt ei caecum et rogabant eum ut illum tangeret
MARK|8|23|et adprehendens manum caeci eduxit eum extra vicum et expuens in oculos eius inpositis manibus suis interrogavit eum si aliquid videret
MARK|8|24|et aspiciens ait video homines velut arbores ambulantes
MARK|8|25|deinde iterum inposuit manus super oculos eius et coepit videre et restitutus est ita ut videret clare omnia
MARK|8|26|et misit illum in domum suam dicens vade in domum tuam et si in vicum introieris nemini dixeris
MARK|8|27|et egressus est Iesus et discipuli eius in castella Caesareae Philippi et in via interrogabat discipulos suos dicens eis quem me dicunt esse homines
MARK|8|28|qui responderunt illi dicentes Iohannem Baptistam alii Heliam alii vero quasi unum de prophetis
MARK|8|29|tunc dicit illis vos vero quem me dicitis esse respondens Petrus ait ei tu es Christus
MARK|8|30|et comminatus est eis ne cui dicerent de illo
MARK|8|31|et coepit docere illos quoniam oportet Filium hominis multa pati et reprobari a senioribus et a summis sacerdotibus et scribis et occidi et post tres dies resurgere
MARK|8|32|et palam verbum loquebatur et adprehendens eum Petrus coepit increpare eum
MARK|8|33|qui conversus et videns discipulos suos comminatus est Petro dicens vade retro me Satana quoniam non sapis quae Dei sunt sed quae sunt hominum
MARK|8|34|et convocata turba cum discipulis suis dixit eis si quis vult post me sequi deneget se ipsum et tollat crucem suam et sequatur me
MARK|8|35|qui enim voluerit animam suam salvam facere perdet eam qui autem perdiderit animam suam propter me et evangelium salvam eam faciet
MARK|8|36|quid enim proderit homini si lucretur mundum totum et detrimentum faciat animae suae
MARK|8|37|aut quid dabit homo commutationem pro anima sua
MARK|8|38|qui enim me confusus fuerit et mea verba in generatione ista adultera et peccatrice et Filius hominis confundetur eum cum venerit in gloria Patris sui cum angelis sanctis
MARK|8|39|et dicebat illis amen dico vobis quia sunt quidam de hic stantibus qui non gustabunt mortem donec videant regnum Dei veniens in virtute
MARK|9|1|et post dies sex adsumit Iesus Petrum et Iacobum et Iohannem et ducit illos in montem excelsum seorsum solos et transfiguratus est coram ipsis
MARK|9|2|et vestimenta eius facta sunt splendentia candida nimis velut nix qualia fullo super terram non potest candida facere
MARK|9|3|et apparuit illis Helias cum Mose et erant loquentes cum Iesu
MARK|9|4|et respondens Petrus ait Iesu rabbi bonum est hic nos esse et faciamus tria tabernacula tibi unum et Mosi unum et Heliae unum
MARK|9|5|non enim sciebat quid diceret erant enim timore exterriti
MARK|9|6|et facta est nubes obumbrans eos et venit vox de nube dicens hic est Filius meus carissimus audite illum
MARK|9|7|et statim circumspicientes neminem amplius viderunt nisi Iesum tantum secum
MARK|9|8|et descendentibus illis de monte praecepit illis ne cui quae vidissent narrarent nisi cum Filius hominis a mortuis resurrexerit
MARK|9|9|et verbum continuerunt apud se conquirentes quid esset cum a mortuis resurrexerit
MARK|9|10|et interrogabant eum dicentes quid ergo dicunt Pharisaei et scribae quia Heliam oporteat venire primum
MARK|9|11|qui respondens ait illis Helias cum venerit primo restituet omnia et quomodo scriptum est in Filium hominis ut multa patiatur et contemnatur
MARK|9|12|sed dico vobis quia et Helias venit et fecerunt illi quaecumque voluerunt sicut scriptum est de eo
MARK|9|13|et veniens ad discipulos suos vidit turbam magnam circa eos et scribas conquirentes cum illis
MARK|9|14|et confestim omnis populus videns eum stupefactus est et adcurrentes salutabant eum
MARK|9|15|et interrogavit eos quid inter vos conquiritis
MARK|9|16|et respondens unus de turba dixit magister adtuli filium meum ad te habentem spiritum mutum
MARK|9|17|qui ubicumque eum adprehenderit adlidit eum et spumat et stridet dentibus et arescit et dixi discipulis tuis ut eicerent illum et non potuerunt
MARK|9|18|qui respondens eis dicit o generatio incredula quamdiu apud vos ero quamdiu vos patiar adferte illum ad me
MARK|9|19|et adtulerunt eum et cum vidisset illum statim spiritus conturbavit eum et elisus in terram volutabatur spumans
MARK|9|20|et interrogavit patrem eius quantum temporis est ex quo hoc ei accidit at ille ait ab infantia
MARK|9|21|et frequenter eum et in ignem et in aquas misit ut eum perderet sed si quid potes adiuva nos misertus nostri
MARK|9|22|Iesus autem ait illi si potes credere omnia possibilia credenti
MARK|9|23|et continuo exclamans pater pueri cum lacrimis aiebat credo adiuva incredulitatem meam
MARK|9|24|et cum videret Iesus concurrentem turbam comminatus est spiritui inmundo dicens illi surde et mute spiritus ego tibi praecipio exi ab eo et amplius ne introeas in eum
MARK|9|25|et clamans et multum discerpens eum exiit ab eo et factus est sicut mortuus ita ut multi dicerent quia mortuus est
MARK|9|26|Iesus autem tenens manum eius elevavit illum et surrexit
MARK|9|27|et cum introisset in domum discipuli eius secreto interrogabant eum quare nos non potuimus eicere eum
MARK|9|28|et dixit illis hoc genus in nullo potest exire nisi in oratione et ieiunio
MARK|9|29|et inde profecti praetergrediebantur Galilaeam nec volebat quemquam scire
MARK|9|30|docebat autem discipulos suos et dicebat illis quoniam Filius hominis tradetur in manus hominum et occident eum et occisus tertia die resurget
MARK|9|31|at illi ignorabant verbum et timebant eum interrogare
MARK|9|32|et venerunt Capharnaum qui cum domi esset interrogabat eos quid in via tractabatis
MARK|9|33|at illi tacebant siquidem inter se in via disputaverant quis esset illorum maior
MARK|9|34|et residens vocavit duodecim et ait illis si quis vult primus esse erit omnium novissimus et omnium minister
MARK|9|35|et accipiens puerum statuit eum in medio eorum quem cum conplexus esset ait illis
MARK|9|36|quisquis unum ex huiusmodi pueris receperit in nomine meo me recipit et quicumque me susceperit non me suscipit sed eum qui me misit
MARK|9|37|respondit illi Iohannes dicens magister vidimus quendam in nomine tuo eicientem daemonia qui non sequitur nos et prohibuimus eum
MARK|9|38|Iesus autem ait nolite prohibere eum nemo est enim qui faciat virtutem in nomine meo et possit cito male loqui de me
MARK|9|39|qui enim non est adversum vos pro vobis est
MARK|9|40|quisquis enim potum dederit vobis calicem aquae in nomine meo quia Christi estis amen dico vobis non perdet mercedem suam
MARK|9|41|et quisquis scandalizaverit unum ex his pusillis credentibus in me bonum est ei magis si circumdaretur mola asinaria collo eius et in mare mitteretur
MARK|9|42|et si scandalizaverit te manus tua abscide illam bonum est tibi debilem introire in vitam quam duas manus habentem ire in gehennam in ignem inextinguibilem
MARK|9|43|ubi vermis eorum non moritur et ignis non extinguitur
MARK|9|44|et si pes tuus te scandalizat amputa illum bonum est tibi claudum introire in vitam aeternam quam duos pedes habentem mitti in gehennam ignis inextinguibilis
MARK|9|45|ubi vermis eorum non moritur et ignis non extinguitur
MARK|9|46|quod si oculus tuus scandalizat te eice eum bonum est tibi luscum introire in regnum Dei quam duos oculos habentem mitti in gehennam ignis
MARK|9|47|ubi vermis eorum non moritur et ignis non extinguitur
MARK|9|48|omnis enim igne sallietur et omnis victima sallietur
MARK|9|49|bonum est sal quod si sal insulsum fuerit in quo illud condietis habete in vobis sal et pacem habete inter vos
MARK|9|50|
MARK|10|1|et inde exsurgens venit in fines Iudaeae ultra Iordanen et conveniunt iterum turbae ad eum et sicut consueverat iterum docebat illos
MARK|10|2|et accedentes Pharisaei interrogabant eum si licet viro uxorem dimittere temptantes eum
MARK|10|3|at ille respondens dixit eis quid vobis praecepit Moses
MARK|10|4|qui dixerunt Moses permisit libellum repudii scribere et dimittere
MARK|10|5|quibus respondens Iesus ait ad duritiam cordis vestri scripsit vobis praeceptum istud
MARK|10|6|ab initio autem creaturae masculum et feminam fecit eos Deus
MARK|10|7|propter hoc relinquet homo patrem suum et matrem et adherebit ad uxorem suam
MARK|10|8|et erunt duo in carne una itaque iam non sunt duo sed una caro
MARK|10|9|quod ergo Deus iunxit homo non separet
MARK|10|10|et in domo iterum discipuli eius de eodem interrogaverunt eum
MARK|10|11|et dicit illis quicumque dimiserit uxorem suam et aliam duxerit adulterium committit super eam
MARK|10|12|et si uxor dimiserit virum suum et alii nupserit moechatur
MARK|10|13|et offerebant illi parvulos ut tangeret illos discipuli autem comminabantur offerentibus
MARK|10|14|quos cum videret Iesus indigne tulit et ait illis sinite parvulos venire ad me et ne prohibueritis eos talium est enim regnum Dei
MARK|10|15|amen dico vobis quisque non receperit regnum Dei velut parvulus non intrabit in illud
MARK|10|16|et conplexans eos et inponens manus super illos benedicebat eos
MARK|10|17|et cum egressus esset in viam procurrens quidam genu flexo ante eum rogabat eum magister bone quid faciam ut vitam aeternam percipiam
MARK|10|18|Iesus autem dixit ei quid me dicis bonum nemo bonus nisi unus Deus
MARK|10|19|praecepta nosti ne adulteres ne occidas ne fureris ne falsum testimonium dixeris ne fraudem feceris honora patrem tuum et matrem
MARK|10|20|et ille respondens ait illi magister omnia haec conservavi a iuventute mea
MARK|10|21|Iesus autem intuitus eum dilexit eum et dixit illi unum tibi deest vade quaecumque habes vende et da pauperibus et habebis thesaurum in caelo et veni sequere me
MARK|10|22|qui contristatus in verbo abiit maerens erat enim habens possessiones multas
MARK|10|23|et circumspiciens Iesus ait discipulis suis quam difficile qui pecunias habent in regnum Dei introibunt
MARK|10|24|discipuli autem obstupescebant in verbis eius at Iesus rursus respondens ait illis filioli quam difficile est confidentes in pecuniis regnum Dei introire
MARK|10|25|facilius est camelum per foramen acus transire quam divitem intrare in regnum Dei
MARK|10|26|qui magis admirabantur dicentes ad semet ipsos et quis potest salvus fieri
MARK|10|27|et intuens illos Iesus ait apud homines inpossibile est sed non apud Deum omnia enim possibilia sunt apud Deum
MARK|10|28|coepit Petrus ei dicere ecce nos dimisimus omnia et secuti sumus te
MARK|10|29|respondens Iesus ait amen dico vobis nemo est qui reliquerit domum aut fratres aut sorores aut matrem aut patrem aut filios aut agros propter me et propter evangelium
MARK|10|30|qui non accipiat centies tantum nunc in tempore hoc domos et fratres et sorores et matres et filios et agros cum persecutionibus et in saeculo futuro vitam aeternam
MARK|10|31|multi autem erunt primi novissimi et novissimi primi
MARK|10|32|erant autem in via ascendentes in Hierosolyma et praecedebat illos Iesus et stupebant et sequentes timebant et adsumens iterum duodecim coepit illis dicere quae essent ei ventura
MARK|10|33|quia ecce ascendimus in Hierosolyma et Filius hominis tradetur principibus sacerdotum et scribis et senioribus et damnabunt eum morti et tradent eum gentibus
MARK|10|34|et inludent ei et conspuent eum et flagellabunt eum et interficient eum et tertia die resurget
MARK|10|35|et accedunt ad illum Iacobus et Iohannes filii Zebedaei dicentes magister volumus ut quodcumque petierimus facias nobis
MARK|10|36|at ille dixit eis quid vultis ut faciam vobis
MARK|10|37|et dixerunt da nobis ut unus ad dexteram tuam et alius ad sinistram tuam sedeamus in gloria tua
MARK|10|38|Iesus autem ait eis nescitis quid petatis potestis bibere calicem quem ego bibo aut baptismum quo ego baptizor baptizari
MARK|10|39|at illi dixerunt ei possumus Iesus autem ait eis calicem quidem quem ego bibo bibetis et baptismum quo ego baptizor baptizabimini
MARK|10|40|sedere autem ad dexteram meam vel ad sinistram non est meum dare sed quibus paratum est
MARK|10|41|et audientes decem coeperunt indignari de Iacobo et Iohanne
MARK|10|42|Iesus autem vocans eos ait illis scitis quia hii qui videntur principari gentibus dominantur eis et principes eorum potestatem habent ipsorum
MARK|10|43|non ita est autem in vobis sed quicumque voluerit fieri maior erit vester minister
MARK|10|44|et quicumque voluerit in vobis primus esse erit omnium servus
MARK|10|45|nam et Filius hominis non venit ut ministraretur ei sed ut ministraret et daret animam suam redemptionem pro multis
MARK|10|46|et veniunt Hierichum et proficiscente eo de Hiericho et discipulis eius et plurima multitudine filius Timei Bartimeus caecus sedebat iuxta viam mendicans
MARK|10|47|qui cum audisset quia Iesus Nazarenus est coepit clamare et dicere Fili David Iesu miserere mei
MARK|10|48|et comminabantur illi multi ut taceret at ille multo magis clamabat Fili David miserere mei
MARK|10|49|et stans Iesus praecepit illum vocari et vocant caecum dicentes ei animaequior esto surge vocat te
MARK|10|50|qui proiecto vestimento suo exiliens venit ad eum
MARK|10|51|et respondens illi Iesus dixit quid vis tibi faciam caecus autem dixit ei rabboni ut videam
MARK|10|52|Iesus autem ait illi vade fides tua te salvum fecit et confestim vidit et sequebatur eum in via
MARK|11|1|et cum adpropinquarent Hierosolymae et Bethaniae ad montem Olivarum mittit duos ex discipulis suis
MARK|11|2|et ait illis ite in castellum quod est contra vos et statim introeuntes illuc invenietis pullum ligatum super quem nemo adhuc hominum sedit solvite illum et adducite
MARK|11|3|et si quis vobis dixerit quid facitis dicite quia Domino necessarius est et continuo illum dimittet huc
MARK|11|4|et abeuntes invenerunt pullum ligatum ante ianuam foris in bivio et solvunt eum
MARK|11|5|et quidam de illic stantibus dicebant illis quid facitis solventes pullum
MARK|11|6|qui dixerunt eis sicut praeceperat illis Iesus et dimiserunt eis
MARK|11|7|et duxerunt pullum ad Iesum et inponunt illi vestimenta sua et sedit super eo
MARK|11|8|multi autem vestimenta sua straverunt in via alii autem frondes caedebant de arboribus et sternebant in via
MARK|11|9|et qui praeibant et qui sequebantur clamabant dicentes osanna benedictus qui venit in nomine Domini
MARK|11|10|benedictum quod venit regnum patris nostri David osanna in excelsis
MARK|11|11|et introivit Hierosolyma in templum et circumspectis omnibus cum iam vespera esset hora exivit in Bethania cum duodecim
MARK|11|12|et alia die cum exirent a Bethania esuriit
MARK|11|13|cumque vidisset a longe ficum habentem folia venit si quid forte inveniret in ea et cum venisset ad eam nihil invenit praeter folia non enim erat tempus ficorum
MARK|11|14|et respondens dixit ei iam non amplius in aeternum quisquam fructum ex te manducet et audiebant discipuli eius
MARK|11|15|et veniunt Hierosolymam et cum introisset templum coepit eicere vendentes et ementes in templo et mensas nummulariorum et cathedras vendentium columbas evertit
MARK|11|16|et non sinebat ut quisquam vas transferret per templum
MARK|11|17|et docebat dicens eis non scriptum est quia domus mea domus orationis vocabitur omnibus gentibus vos autem fecistis eam speluncam latronum
MARK|11|18|quo audito principes sacerdotum et scribae quaerebant quomodo eum perderent timebant enim eum quoniam universa turba admirabatur super doctrina eius
MARK|11|19|et cum vespera facta esset egrediebatur de civitate
MARK|11|20|et cum mane transirent viderunt ficum aridam factam a radicibus
MARK|11|21|et recordatus Petrus dicit ei rabbi ecce ficus cui maledixisti aruit
MARK|11|22|et respondens Iesus ait illis habete fidem Dei
MARK|11|23|amen dico vobis quicumque dixerit huic monti tollere et mittere in mare et non haesitaverit in corde suo sed crediderit quia quodcumque dixerit fiat fiet ei
MARK|11|24|propterea dico vobis omnia quaecumque orantes petitis credite quia accipietis et veniet vobis
MARK|11|25|et cum stabitis ad orandum dimittite si quid habetis adversus aliquem ut et Pater vester qui in caelis est dimittat vobis peccata vestra
MARK|11|26|quod si vos non dimiseritis nec Pater vester qui in caelis est dimittet vobis peccata vestra
MARK|11|27|et veniunt rursus Hierosolymam et cum ambularet in templo accedunt ad eum summi sacerdotes et scribae et seniores
MARK|11|28|et dicunt illi in qua potestate haec facis et quis tibi dedit hanc potestatem ut ista facias
MARK|11|29|Iesus autem respondens ait illis interrogabo vos et ego unum verbum et respondete mihi et dicam vobis in qua potestate haec faciam
MARK|11|30|baptismum Iohannis de caelo erat an ex hominibus respondete mihi
MARK|11|31|at illi cogitabant secum dicentes si dixerimus de caelo dicet quare ergo non credidistis ei
MARK|11|32|sed dicemus ex hominibus timebant populum omnes enim habebant Iohannem quia vere propheta esset
MARK|11|33|et respondentes dicunt Iesu nescimus respondens Iesus ait illis neque ego dico vobis in qua potestate haec faciam
MARK|12|1|et coepit illis in parabolis loqui vineam pastinavit homo et circumdedit sepem et fodit lacum et aedificavit turrem et locavit eam agricolis et peregre profectus est
MARK|12|2|et misit ad agricolas in tempore servum ut ab agricolis acciperet de fructu vineae
MARK|12|3|qui adprehensum eum ceciderunt et dimiserunt vacuum
MARK|12|4|et iterum misit ad illos alium servum et illum capite vulneraverunt et contumeliis adfecerunt
MARK|12|5|et rursum alium misit et illum occiderunt et plures alios quosdam caedentes alios vero occidentes
MARK|12|6|adhuc ergo unum habens filium carissimum et illum misit ad eos novissimum dicens quia reverebuntur filium meum
MARK|12|7|coloni autem dixerunt ad invicem hic est heres venite occidamus eum et nostra erit hereditas
MARK|12|8|et adprehendentes eum occiderunt et eiecerunt extra vineam
MARK|12|9|quid ergo faciet dominus vineae veniet et perdet colonos et dabit vineam aliis
MARK|12|10|nec scripturam hanc legistis lapidem quem reprobaverunt aedificantes hic factus est in caput anguli
MARK|12|11|a Domino factum est istud et est mirabile in oculis nostris
MARK|12|12|et quaerebant eum tenere et timuerunt turbam cognoverunt enim quoniam ad eos parabolam hanc dixerit et relicto eo abierunt
MARK|12|13|et mittunt ad eum quosdam ex Pharisaeis et Herodianis ut eum caperent in verbo
MARK|12|14|qui venientes dicunt ei magister scimus quoniam verax es et non curas quemquam nec enim vides in faciem hominis sed in veritate viam Dei doces licet dari tributum Caesari an non dabimus
MARK|12|15|qui sciens versutiam eorum ait illis quid me temptatis adferte mihi denarium ut videam
MARK|12|16|at illi adtulerunt et ait illis cuius est imago haec et inscriptio dicunt illi Caesaris
MARK|12|17|respondens autem Iesus dixit illis reddite igitur quae sunt Caesaris Caesari et quae sunt Dei Deo et mirabantur super eo
MARK|12|18|et venerunt ad eum Sadducaei qui dicunt resurrectionem non esse et interrogabant eum dicentes
MARK|12|19|magister Moses nobis scripsit ut si cuius frater mortuus fuerit et dimiserit uxorem et filios non reliquerit accipiat frater eius uxorem ipsius et resuscitet semen fratri suo
MARK|12|20|septem ergo fratres erant et primus accepit uxorem et mortuus est non relicto semine
MARK|12|21|et secundus accepit eam et mortuus est et nec iste reliquit semen et tertius similiter
MARK|12|22|et acceperunt eam similiter septem et non reliquerunt semen novissima omnium defuncta est et mulier
MARK|12|23|in resurrectione ergo cum resurrexerint cuius de his erit uxor septem enim habuerunt eam uxorem
MARK|12|24|et respondens Iesus ait illis non ideo erratis non scientes scripturas neque virtutem Dei
MARK|12|25|cum enim a mortuis resurrexerint neque nubent neque nubentur sed sunt sicut angeli in caelis
MARK|12|26|de mortuis autem quod resurgant non legistis in libro Mosi super rubum quomodo dixerit illi Deus inquiens ego sum Deus Abraham et Deus Isaac et Deus Iacob
MARK|12|27|non est Deus mortuorum sed vivorum vos ergo multum erratis
MARK|12|28|et accessit unus de scribis qui audierat illos conquirentes et videns quoniam bene illis responderit interrogavit eum quod esset primum omnium mandatum
MARK|12|29|Iesus autem respondit ei quia primum omnium mandatum est audi Israhel Dominus Deus noster Deus unus est
MARK|12|30|et diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex tota mente tua et ex tota virtute tua hoc est primum mandatum
MARK|12|31|secundum autem simile illi diliges proximum tuum tamquam te ipsum maius horum aliud mandatum non est
MARK|12|32|et ait illi scriba bene magister in veritate dixisti quia unus est et non est alius praeter eum
MARK|12|33|et ut diligatur ex toto corde et ex toto intellectu et ex tota anima et ex tota fortitudine et diligere proximum tamquam se ipsum maius est omnibus holocaustomatibus et sacrificiis
MARK|12|34|Iesus autem videns quod sapienter respondisset dixit illi non es longe a regno Dei et nemo iam audebat eum interrogare
MARK|12|35|et respondens Iesus dicebat docens in templo quomodo dicunt scribae Christum Filium esse David
MARK|12|36|ipse enim David dicit in Spiritu Sancto dixit Dominus Domino meo sede a dextris meis donec ponam inimicos tuos scabillum pedum tuorum
MARK|12|37|ipse ergo David dicit eum Dominum et unde est filius eius et multa turba eum libenter audivit
MARK|12|38|et dicebat eis in doctrina sua cavete a scribis qui volunt in stolis ambulare et salutari in foro
MARK|12|39|et in primis cathedris sedere in synagogis et primos discubitus in cenis
MARK|12|40|qui devorant domos viduarum sub obtentu prolixae orationis hii accipient prolixius iudicium
MARK|12|41|et sedens Iesus contra gazofilacium aspiciebat quomodo turba iactaret aes in gazofilacium et multi divites iactabant multa
MARK|12|42|cum venisset autem una vidua pauper misit duo minuta quod est quadrans
MARK|12|43|et convocans discipulos suos ait illis amen dico vobis quoniam vidua haec pauper plus omnibus misit qui miserunt in gazofilacium
MARK|12|44|omnes enim ex eo quod abundabat illis miserunt haec vero de penuria sua omnia quae habuit misit totum victum suum
MARK|13|1|et cum egrederetur de templo ait illi unus ex discipulis suis magister aspice quales lapides et quales structurae
MARK|13|2|et respondens Iesus ait illi vides has omnes magnas aedificationes non relinquetur lapis super lapidem qui non destruatur
MARK|13|3|et cum sederet in montem Olivarum contra templum interrogabant eum separatim Petrus et Iacobus et Iohannes et Andreas
MARK|13|4|dic nobis quando ista fient et quod signum erit quando haec omnia incipient consummari
MARK|13|5|et respondens Iesus coepit dicere illis videte ne quis vos seducat
MARK|13|6|multi enim venient in nomine meo dicentes quia ego sum et multos seducent
MARK|13|7|cum audieritis autem bella et opiniones bellorum ne timueritis oportet enim fieri sed nondum finis
MARK|13|8|exsurget autem gens super gentem et regnum super regnum et erunt terraemotus per loca et fames initium dolorum haec
MARK|13|9|videte autem vosmet ipsos tradent enim vos conciliis et in synagogis vapulabitis et ante praesides et reges stabitis propter me in testimonium illis
MARK|13|10|et in omnes gentes primum oportet praedicari evangelium
MARK|13|11|et cum duxerint vos tradentes nolite praecogitare quid loquamini sed quod datum vobis fuerit in illa hora id loquimini non enim estis vos loquentes sed Spiritus Sanctus
MARK|13|12|tradet autem frater fratrem in mortem et pater filium et consurgent filii in parentes et morte adficient eos
MARK|13|13|et eritis odio omnibus propter nomen meum qui autem sustinuerit in finem hic salvus erit
MARK|13|14|cum autem videritis abominationem desolationis stantem ubi non debet qui legit intellegat tunc qui in Iudaea sunt fugiant in montes
MARK|13|15|et qui super tectum ne descendat in domum nec introeat ut tollat quid de domo sua
MARK|13|16|et qui in agro erit non revertatur retro tollere vestimentum suum
MARK|13|17|vae autem praegnatibus et nutrientibus in illis diebus
MARK|13|18|orate vero ut hieme non fiant
MARK|13|19|erunt enim dies illi tribulationes tales quales non fuerunt ab initio creaturae quam condidit Deus usque nunc neque fient
MARK|13|20|et nisi breviasset Dominus dies non fuisset salva omnis caro sed propter electos quos elegit breviavit dies
MARK|13|21|et tunc si quis vobis dixerit ecce hic est Christus ecce illic ne credideritis
MARK|13|22|exsurgent enim pseudochristi et pseudoprophetae et dabunt signa et portenta ad seducendos si potest fieri etiam electos
MARK|13|23|vos ergo videte ecce praedixi vobis omnia
MARK|13|24|sed in illis diebus post tribulationem illam sol contenebrabitur et luna non dabit splendorem suum
MARK|13|25|et erunt stellae caeli decidentes et virtutes quae sunt in caelis movebuntur
MARK|13|26|et tunc videbunt Filium hominis venientem in nubibus cum virtute multa et gloria
MARK|13|27|et tunc mittet angelos suos et congregabit electos suos a quattuor ventis a summo terrae usque ad summum caeli
MARK|13|28|a ficu autem discite parabolam cum iam ramus eius tener fuerit et nata fuerint folia cognoscitis quia in proximo sit aestas
MARK|13|29|sic et vos cum videritis haec fieri scitote quod in proximo sit in ostiis
MARK|13|30|amen dico vobis quoniam non transiet generatio haec donec omnia ista fiant
MARK|13|31|caelum et terra transibunt verba autem mea non transibunt
MARK|13|32|de die autem illo vel hora nemo scit neque angeli in caelo neque Filius nisi Pater
MARK|13|33|videte vigilate et orate nescitis enim quando tempus sit
MARK|13|34|sicut homo qui peregre profectus reliquit domum suam et dedit servis suis potestatem cuiusque operis et ianitori praecipiat ut vigilet
MARK|13|35|vigilate ergo nescitis enim quando dominus domus veniat sero an media nocte an galli cantu an mane
MARK|13|36|ne cum venerit repente inveniat vos dormientes
MARK|13|37|quod autem vobis dico omnibus dico vigilate
MARK|14|1|erat autem pascha et azyma post biduum et quaerebant summi sacerdotes et scribae quomodo eum dolo tenerent et occiderent
MARK|14|2|dicebant enim non in die festo ne forte tumultus fieret populi
MARK|14|3|et cum esset Bethaniae in domo Simonis leprosi et recumberet venit mulier habens alabastrum unguenti nardi spicati pretiosi et fracto alabastro effudit super caput eius
MARK|14|4|erant autem quidam indigne ferentes intra semet ipsos et dicentes ut quid perditio ista unguenti facta est
MARK|14|5|poterat enim unguentum istud veniri plus quam trecentis denariis et dari pauperibus et fremebant in eam
MARK|14|6|Iesus autem dixit sinite eam quid illi molesti estis bonum opus operata est in me
MARK|14|7|semper enim pauperes habetis vobiscum et cum volueritis potestis illis benefacere me autem non semper habetis
MARK|14|8|quod habuit haec fecit praevenit unguere corpus meum in sepulturam
MARK|14|9|amen dico vobis ubicumque praedicatum fuerit evangelium istud in universum mundum et quod fecit haec narrabitur in memoriam eius
MARK|14|10|et Iudas Scariotis unus de duodecim abiit ad summos sacerdotes ut proderet eum illis
MARK|14|11|qui audientes gavisi sunt et promiserunt ei pecuniam se daturos et quaerebat quomodo illum oportune traderet
MARK|14|12|et primo die azymorum quando pascha immolabant dicunt ei discipuli quo vis eamus et paremus tibi ut manduces pascha
MARK|14|13|et mittit duos ex discipulis suis et dicit eis ite in civitatem et occurret vobis homo laguenam aquae baiulans sequimini eum
MARK|14|14|et quocumque introierit dicite domino domus quia magister dicit ubi est refectio mea ubi pascha cum discipulis meis manducem
MARK|14|15|et ipse vobis demonstrabit cenaculum grande stratum et illic parate nobis
MARK|14|16|et abierunt discipuli eius et venerunt in civitatem et invenerunt sicut dixerat illis et praeparaverunt pascha
MARK|14|17|vespere autem facto venit cum duodecim
MARK|14|18|et discumbentibus eis et manducantibus ait Iesus amen dico vobis quia unus ex vobis me tradet qui manducat mecum
MARK|14|19|at illi coeperunt contristari et dicere ei singillatim numquid ego
MARK|14|20|qui ait illis unus ex duodecim qui intinguit mecum in catino
MARK|14|21|et Filius quidem hominis vadit sicut scriptum est de eo vae autem homini illi per quem Filius hominis traditur bonum ei si non esset natus homo ille
MARK|14|22|et manducantibus illis accepit Iesus panem et benedicens fregit et dedit eis et ait sumite hoc est corpus meum
MARK|14|23|et accepto calice gratias agens dedit eis et biberunt ex illo omnes
MARK|14|24|et ait illis hic est sanguis meus novi testamenti qui pro multis effunditur
MARK|14|25|amen dico vobis quod iam non bibam de genimine vitis usque in diem illum cum illud bibam novum in regno Dei
MARK|14|26|et hymno dicto exierunt in montem Olivarum
MARK|14|27|et ait eis Iesus omnes scandalizabimini in nocte ista quia scriptum est percutiam pastorem et dispergentur oves
MARK|14|28|sed posteaquam resurrexero praecedam vos in Galilaeam
MARK|14|29|Petrus autem ait ei et si omnes scandalizati fuerint sed non ego
MARK|14|30|et ait illi Iesus amen dico tibi quia tu hodie in nocte hac priusquam bis gallus vocem dederit ter me es negaturus
MARK|14|31|at ille amplius loquebatur et si oportuerit me simul conmori tibi non te negabo similiter autem et omnes dicebant
MARK|14|32|et veniunt in praedium cui nomen Gethsemani et ait discipulis suis sedete hic donec orem
MARK|14|33|et adsumit Petrum et Iacobum et Iohannem secum et coepit pavere et taedere
MARK|14|34|et ait illis tristis est anima mea usque ad mortem sustinete hic et vigilate
MARK|14|35|et cum processisset paululum procidit super terram et orabat ut si fieri posset transiret ab eo hora
MARK|14|36|et dixit Abba Pater omnia possibilia tibi sunt transfer calicem hunc a me sed non quod ego volo sed quod tu
MARK|14|37|et venit et invenit eos dormientes et ait Petro Simon dormis non potuisti una hora vigilare
MARK|14|38|vigilate et orate ut non intretis in temptationem spiritus quidem promptus caro vero infirma
MARK|14|39|et iterum abiens oravit eundem sermonem dicens
MARK|14|40|et reversus denuo invenit eos dormientes erant enim oculi illorum ingravati et ignorabant quid responderent ei
MARK|14|41|et venit tertio et ait illis dormite iam et requiescite sufficit venit hora ecce traditur Filius hominis in manus peccatorum
MARK|14|42|surgite eamus ecce qui me tradit prope est
MARK|14|43|et adhuc eo loquente venit Iudas Scarioth unus ex duodecim et cum illo turba cum gladiis et lignis a summis sacerdotibus et a scribis et a senioribus
MARK|14|44|dederat autem traditor eius signum eis dicens quemcumque osculatus fuero ipse est tenete eum et ducite
MARK|14|45|et cum venisset statim accedens ad eum ait rabbi et osculatus est eum
MARK|14|46|at illi manus iniecerunt in eum et tenuerunt eum
MARK|14|47|unus autem quidam de circumstantibus educens gladium percussit servum summi sacerdotis et amputavit illi auriculam
MARK|14|48|et respondens Iesus ait illis tamquam ad latronem existis cum gladiis et lignis conprehendere me
MARK|14|49|cotidie eram apud vos in templo docens et non me tenuistis sed ut adimpleantur scripturae
MARK|14|50|tunc discipuli eius relinquentes eum omnes fugerunt
MARK|14|51|adulescens autem quidam sequebatur illum amictus sindone super nudo et tenuerunt eum
MARK|14|52|at ille reiecta sindone nudus profugit ab eis
MARK|14|53|et adduxerunt Iesum ad summum sacerdotem et conveniunt omnes sacerdotes et scribae et seniores
MARK|14|54|Petrus autem a longe secutus est eum usque intro in atrium summi sacerdotis et sedebat cum ministris et calefaciebat se ad ignem
MARK|14|55|summi vero sacerdotes et omne concilium quaerebant adversum Iesum testimonium ut eum morti traderent nec inveniebant
MARK|14|56|multi enim testimonium falsum dicebant adversus eum et convenientia testimonia non erant
MARK|14|57|et quidam surgentes falsum testimonium ferebant adversus eum dicentes
MARK|14|58|quoniam nos audivimus eum dicentem ego dissolvam templum hoc manufactum et per triduum aliud non manufactum aedificabo
MARK|14|59|et non erat conveniens testimonium illorum
MARK|14|60|et exsurgens summus sacerdos in medium interrogavit Iesum dicens non respondes quicquam ad ea quae tibi obiciuntur ab his
MARK|14|61|ille autem tacebat et nihil respondit rursum summus sacerdos interrogabat eum et dicit ei tu es Christus Filius Benedicti
MARK|14|62|Iesus autem dixit illi ego sum et videbitis Filium hominis a dextris sedentem Virtutis et venientem cum nubibus caeli
MARK|14|63|summus autem sacerdos scindens vestimenta sua ait quid adhuc desideramus testes
MARK|14|64|audistis blasphemiam quid vobis videtur qui omnes condemnaverunt eum esse reum mortis
MARK|14|65|et coeperunt quidam conspuere eum et velare faciem eius et colaphis eum caedere et dicere ei prophetiza et ministri alapis eum caedebant
MARK|14|66|et cum esset Petrus in atrio deorsum venit una ex ancillis summi sacerdotis
MARK|14|67|et cum vidisset Petrum calefacientem se aspiciens illum ait et tu cum Iesu Nazareno eras
MARK|14|68|at ille negavit dicens neque scio neque novi quid dicas et exiit foras ante atrium et gallus cantavit
MARK|14|69|rursus autem cum vidisset illum ancilla coepit dicere circumstantibus quia hic ex illis est
MARK|14|70|at ille iterum negavit et post pusillum rursus qui adstabant dicebant Petro vere ex illis es nam et Galilaeus es
MARK|14|71|ille autem coepit anathematizare et iurare quia nescio hominem istum quem dicitis
MARK|14|72|et statim iterum gallus cantavit et recordatus est Petrus verbi quod dixerat ei Iesus priusquam gallus cantet bis ter me negabis et coepit flere
MARK|15|1|et confestim mane consilium facientes summi sacerdotes cum senioribus et scribis et universo concilio vincientes Iesum duxerunt et tradiderunt Pilato
MARK|15|2|et interrogavit eum Pilatus tu es rex Iudaeorum at ille respondens ait illi tu dicis
MARK|15|3|et accusabant eum summi sacerdotes in multis
MARK|15|4|Pilatus autem rursum interrogavit eum dicens non respondes quicquam vide in quantis te accusant
MARK|15|5|Iesus autem amplius nihil respondit ita ut miraretur Pilatus
MARK|15|6|per diem autem festum dimittere solebat illis unum ex vinctis quemcumque petissent
MARK|15|7|erat autem qui dicebatur Barabbas qui cum seditiosis erat vinctus qui in seditione fecerant homicidium
MARK|15|8|et cum ascendisset turba coepit rogare sicut semper faciebat illis
MARK|15|9|Pilatus autem respondit eis et dixit vultis dimittam vobis regem Iudaeorum
MARK|15|10|sciebat enim quod per invidiam tradidissent eum summi sacerdotes
MARK|15|11|pontifices autem concitaverunt turbam ut magis Barabban dimitteret eis
MARK|15|12|Pilatus autem iterum respondens ait illis quid ergo vultis faciam regi Iudaeorum
MARK|15|13|at illi iterum clamaverunt crucifige eum
MARK|15|14|Pilatus vero dicebat eis quid enim mali fecit at illi magis clamabant crucifige eum
MARK|15|15|Pilatus autem volens populo satisfacere dimisit illis Barabban et tradidit Iesum flagellis caesum ut crucifigeretur
MARK|15|16|milites autem duxerunt eum intro in atrium praetorii et convocant totam cohortem
MARK|15|17|et induunt eum purpuram et inponunt ei plectentes spineam coronam
MARK|15|18|et coeperunt salutare eum have rex Iudaeorum
MARK|15|19|et percutiebant caput eius harundine et conspuebant eum et ponentes genua adorabant eum
MARK|15|20|et postquam inluserunt ei exuerunt illum purpuram et induerunt eum vestimentis suis et educunt illum ut crucifigerent eum
MARK|15|21|et angariaverunt praetereuntem quempiam Simonem Cyreneum venientem de villa patrem Alexandri et Rufi ut tolleret crucem eius
MARK|15|22|et perducunt illum in Golgotha locum quod est interpretatum Calvariae locus
MARK|15|23|et dabant ei bibere murratum vinum et non accepit
MARK|15|24|et crucifigentes eum diviserunt vestimenta eius mittentes sortem super eis quis quid tolleret
MARK|15|25|erat autem hora tertia et crucifixerunt eum
MARK|15|26|et erat titulus causae eius inscriptus rex Iudaeorum
MARK|15|27|et cum eo crucifigunt duos latrones unum a dextris et alium a sinistris eius
MARK|15|28|et adimpleta est scriptura quae dicit et cum iniquis reputatus est
MARK|15|29|et praetereuntes blasphemabant eum moventes capita sua et dicentes va qui destruit templum et in tribus diebus aedificat
MARK|15|30|salvum fac temet ipsum descendens de cruce
MARK|15|31|similiter et summi sacerdotes ludentes ad alterutrum cum scribis dicebant alios salvos fecit se ipsum non potest salvum facere
MARK|15|32|Christus rex Israhel descendat nunc de cruce ut videamus et credamus et qui cum eo crucifixi erant conviciabantur ei
MARK|15|33|et facta hora sexta tenebrae factae sunt per totam terram usque in horam nonam
MARK|15|34|et hora nona exclamavit Iesus voce magna dicens Heloi Heloi lama sabacthani quod est interpretatum Deus meus Deus meus ut quid dereliquisti me
MARK|15|35|et quidam de circumstantibus audientes dicebant ecce Heliam vocat
MARK|15|36|currens autem unus et implens spongiam aceto circumponensque calamo potum dabat ei dicens sinite videamus si veniat Helias ad deponendum eum
MARK|15|37|Iesus autem emissa voce magna exspiravit
MARK|15|38|et velum templi scissum est in duo a sursum usque deorsum
MARK|15|39|videns autem centurio qui ex adverso stabat quia sic clamans exspirasset ait vere homo hic Filius Dei erat
MARK|15|40|erant autem et mulieres de longe aspicientes inter quas et Maria Magdalene et Maria Iacobi minoris et Ioseph mater et Salome
MARK|15|41|et cum esset in Galilaea sequebantur eum et ministrabant ei et aliae multae quae simul cum eo ascenderant Hierosolyma
MARK|15|42|et cum iam sero esset factum quia erat parasceve quod est ante sabbatum
MARK|15|43|venit Ioseph ab Arimathia nobilis decurio qui et ipse erat expectans regnum Dei et audacter introiit ad Pilatum et petiit corpus Iesu
MARK|15|44|Pilatus autem mirabatur si iam obisset et accersito centurione interrogavit eum si iam mortuus esset
MARK|15|45|et cum cognovisset a centurione donavit corpus Ioseph
MARK|15|46|Ioseph autem mercatus sindonem et deponens eum involvit sindone et posuit eum in monumento quod erat excisum de petra et advolvit lapidem ad ostium monumenti
MARK|15|47|Maria autem Magdalene et Maria Ioseph aspiciebant ubi poneretur
MARK|16|1|et cum transisset sabbatum Maria Magdalene et Maria Iacobi et Salome emerunt aromata ut venientes unguerent eum
MARK|16|2|et valde mane una sabbatorum veniunt ad monumentum orto iam sole
MARK|16|3|et dicebant ad invicem quis revolvet nobis lapidem ab ostio monumenti
MARK|16|4|et respicientes vident revolutum lapidem erat quippe magnus valde
MARK|16|5|et introeuntes in monumento viderunt iuvenem sedentem in dextris coopertum stola candida et obstipuerunt
MARK|16|6|qui dicit illis nolite expavescere Iesum quaeritis Nazarenum crucifixum surrexit non est hic ecce locus ubi posuerunt eum
MARK|16|7|sed ite et dicite discipulis eius et Petro quia praecedit vos in Galilaeam ibi eum videbitis sicut dixit vobis
MARK|16|8|at illae exeuntes fugerunt de monumento invaserat enim eas tremor et pavor et nemini quicquam dixerunt timebant enim
MARK|16|9|surgens autem mane prima sabbati apparuit primo Mariae Magdalenae de qua eiecerat septem daemonia
MARK|16|10|illa vadens nuntiavit his qui cum eo fuerant lugentibus et flentibus
MARK|16|11|et illi audientes quia viveret et visus esset ab ea non crediderunt
MARK|16|12|post haec autem duobus ex eis ambulantibus ostensus est in alia effigie euntibus in villam
MARK|16|13|et illi euntes nuntiaverunt ceteris nec illis crediderunt
MARK|16|14|novissime recumbentibus illis undecim apparuit et exprobravit incredulitatem illorum et duritiam cordis quia his qui viderant eum resurrexisse non crediderant
MARK|16|15|et dixit eis euntes in mundum universum praedicate evangelium omni creaturae
MARK|16|16|qui crediderit et baptizatus fuerit salvus erit qui vero non crediderit condemnabitur
MARK|16|17|signa autem eos qui crediderint haec sequentur in nomine meo daemonia eicient linguis loquentur novis
MARK|16|18|serpentes tollent et si mortiferum quid biberint non eos nocebit super aegrotos manus inponent et bene habebunt
MARK|16|19|et Dominus quidem postquam locutus est eis adsumptus est in caelum et sedit a dextris Dei
MARK|16|20|illi autem profecti praedicaverunt ubique Domino cooperante et sermonem confirmante sequentibus signis
