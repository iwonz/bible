HAG|1|1|In anno secundo Darii regis, in mense sexto, in die prima men sis, factum est verbum Domini in manu Aggaei prophetae ad Zorobabel filium Salathiel ducem Iudae et ad Iesua filium Iosedec sacerdotem magnum dicens:
HAG|1|2|" Haec ait Dominus exercituum dicens: Populus iste dicit: "Nondum venit tempus domus Domini aedificandae" ".
HAG|1|3|Et factum est verbum Domini in manu Aggaei prophetae dicens:
HAG|1|4|" Numquid tempus vobis est, ut habitetis in domibus laqueatis, et domus ista deserta?
HAG|1|5|Et nunc haec dicit Dominus exercituum: Ponite corda vestra super vias vestras:
HAG|1|6|seminastis multum et intulistis parum, comedistis et non estis satiati, bibistis et non estis inebriati, operuistis vos et non estis calefacti, et, qui pro mercede operatus est, misit eam in sacculum pertusum.
HAG|1|7|Haec dicit Dominus exercituum: Ponite corda vestra super vias vestras.
HAG|1|8|Ascendite in montem, portate lignum et aedificate domum, et acceptabilis mihi erit et glorificabor, dicit Dominus.
HAG|1|9|Respexistis ad amplius, et ecce factum est minus; et intulistis in domum, et exsufflavi illud. Quam ob causam?, dicit Dominus exercituum. Quia domus mea deserta est, et vos festinatis unusquisque in domum suam.
HAG|1|10|Propter hoc super vos prohibiti sunt caeli, ne darent rorem, et terra prohibita est, ne daret fructum suum.
HAG|1|11|Et vocavi siccitatem super terram et super montes et super triticum et super vinum et super oleum et, quaecumque profert humus, et super homines et super iumenta et super omnem laborem manuum ".
HAG|1|12|Et audivit Zorobabel filius Salathiel et Iesua filius Iosedec sacerdos magnus et omnes reliquiae populi vocem Domini Dei sui et verba Aggaei prophetae, sicut misit eum Dominus Deus eorum ad ipsos; et timuit populus a facie Domini.
HAG|1|13|Et dixit Aggaeus nuntius Domini secundum mandatum Domini populo dicens: Ego vobiscum, dicit Dominus ".
HAG|1|14|Et suscitavit Dominus spiritum Zorobabel filii Salathiel ducis Iudae et spiritum Iesua filii Iosedec sacerdotis magni et spiritum reliquorum omnium de populo; et ingressi sunt et faciebant opus in domo Domini exercituum Dei sui.
HAG|1|15|In die vicesima et quarta mensis, in sexto mense, in anno secundo Darii regis.
HAG|2|1|In septimo mense, vicesima et prima mensis, factum est ver bum Domini in manu Aggaei prophetae dicens:
HAG|2|2|" Loquere ad Zorobabel filium Salathiel ducem Iudae et ad Iesua filium Iosedec sacerdotem magnum et ad reliquos populi dicens:
HAG|2|3|Quis in vobis est derelictus, qui vidit domum istam in gloria sua prima? Et quid vos videtis eam nunc? Numquid non ita est quasi non sit in oculis vestris?
HAG|2|4|Sed et nunc confortare, Zorobabel, dicit Dominus, et confortare, Iesua fili Iosedec sacerdos magne, et confortare, omnis popule terrae, dicit Dominus exercituum; et facite, quoniam ego vobiscum sum, dicit Dominus exercituum.
HAG|2|5|Verbum quod pepigi vobiscum, cum egrederemini de terra Aegypti, et spiritus meus stat in medio vestrum; nolite timere.
HAG|2|6|Quia haec dicit Dominus exercituum: Adhuc unum modicum est, et ego commovebo caelum et terram et mare et aridam.
HAG|2|7|Et movebo omnes gentes, et venient thesauri cunctarum gentium, et implebo domum istam gloria, dicit Dominus exercituum.
HAG|2|8|Meum est argentum et meum est aurum, dicit Dominus exercituum.
HAG|2|9|Maior erit gloria domus istius novissima plus quam prima, dicit Dominus exercituum; et in loco isto dabo pacem, dicit Dominus exercituum ".
HAG|2|10|In vicesima et quarta noni mensis, in anno secundo Darii, factum est verbum Domini ad Aggaeum prophetam dicens:
HAG|2|11|" Haec dicit Dominus exercituum: Interroga sacerdotes legem dicens:
HAG|2|12|Si tulerit homo carnem sanctificatam in ora vestimenti sui et tetigerit de summitate eius panem aut pulmentum aut vinum aut oleum aut omnem cibum, numquid sanctificabitur? ". Respondentes autem sacerdotes dixerunt: " Non.
HAG|2|13|Et dixit Aggaeus: " Si tetigerit pollutus cadavere omnia haec, numquid contaminabuntur? ". Et responderunt sacerdotes et dixerunt: " Contaminabuntur ".
HAG|2|14|Et respondit Aggaeus et dixit: " Sic populus iste et sic gens ista ante faciem meam, dicit Dominus, et sic omne opus manuum eorum et omnia, quae offerunt ibi, contaminata sunt.
HAG|2|15|Et nunc ponite corda vestra a die hac et supra: Antequam poneretur lapis super lapidem in templo Domini,
HAG|2|16|quid fuistis? Cum accederetis ad acervum viginti modiorum, erant decem; cum intraretis ad torcular, ut hauriretis quinquaginta lagenas, erant viginti.
HAG|2|17|Percussi vos ariditate et rubigine et grandine omnia opera manuum vestrarum, et non fuit in vobis qui reverteretur ad me, dicit Dominus.
HAG|2|18|Ponite corda vestra ex die ista et in futurum, a die vicesima et quarta noni mensis, a die, qua fundamenta iacta sunt templi Domini, ponite super cor vestrum.
HAG|2|19|Numquid adhuc semen in horreo est, et adhuc vinea et ficus et malogranatum et lignum olivae non portavit fructum? Ex die hac benedicam.
HAG|2|20|Et factum est verbum Domini secundo ad Aggaeum in vicesima et quarta mensis dicens:
HAG|2|21|" Loquere ad Zorobabel ducem Iudae dicens: Ego movebo caelum pariter et terram
HAG|2|22|et subvertam solium regnorum et conteram fortitudinem regnorum gentium et subvertam quadrigam et ascensores eius; et descendent equi et ascensores eorum, unusquisque percussus gladio fratris sui.
HAG|2|23|In die illo, dicit Dominus exercituum, assumam te, Zorobabel fili Salathiel, serve meus, dicit Dominus, et ponam te quasi signaculum, quia te elegi ", dicit Dominus exercituum.
