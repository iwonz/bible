JER|1|1|verba Hieremiae filii Helciae de sacerdotibus qui fuerunt in Anathoth in terra Beniamin
JER|1|2|quod factum est verbum Domini ad eum in diebus Iosiae filii Amon regis Iuda in tertiodecimo anno regni eius
JER|1|3|et factum est in diebus Ioachim filii Iosiae regis Iuda usque ad consummationem undecimi anni Sedeciae filii Iosiae regis Iuda usque ad transmigrationem Hierusalem in mense quinto
JER|1|4|et factum est verbum Domini ad me dicens
JER|1|5|priusquam te formarem in utero novi te et antequam exires de vulva sanctificavi te prophetam gentibus dedi te
JER|1|6|et dixi a a a Domine Deus ecce nescio loqui quia puer ego sum
JER|1|7|et dixit Dominus ad me noli dicere puer sum quoniam ad omnia quae mittam te ibis et universa quaecumque mandavero tibi loqueris
JER|1|8|ne timeas a facie eorum quia tecum ego sum ut eruam te dicit Dominus
JER|1|9|et misit Dominus manum suam et tetigit os meum et dixit Dominus ad me ecce dedi verba mea in ore tuo
JER|1|10|ecce constitui te hodie super gentes et super regna ut evellas et destruas et disperdas et dissipes et aedifices et plantes
JER|1|11|et factum est verbum Domini ad me dicens quid tu vides Hieremia et dixi virgam vigilantem ego video
JER|1|12|et dixit Dominus ad me bene vidisti quia vigilabo ego super verbo meo ut faciam illud
JER|1|13|et factum est verbum Domini secundo ad me dicens quid tu vides et dixi ollam succensam ego video et faciem eius a facie aquilonis
JER|1|14|et dixit Dominus ad me ab aquilone pandetur malum super omnes habitatores terrae
JER|1|15|quia ecce ego convocabo omnes cognationes regnorum aquilonis ait Dominus et venient et ponent unusquisque solium suum in introitu portarum Hierusalem et super omnes muros eius in circuitu et super universas urbes Iuda
JER|1|16|et loquar iudicia mea cum eis super omni malitia eorum qui dereliquerunt me et libaverunt diis alienis et adoraverunt opus manuum suarum
JER|1|17|tu ergo accinge lumbos tuos et surge et loquere ad eos omnia quae ego praecipio tibi ne formides a facie eorum nec enim timere te faciam vultum eorum
JER|1|18|ego quippe dedi te hodie in civitatem munitam et in columnam ferream et in murum aereum super omnem terram regibus Iuda principibus eius et sacerdotibus et populo terrae
JER|1|19|et bellabunt adversum te et non praevalebunt quia tecum ego sum ait Dominus ut liberem te
JER|2|1|et factum est verbum Domini ad me dicens
JER|2|2|vade et clama in auribus Hierusalem dicens haec dicit Dominus recordatus sum tui miserans adulescentiam tuam et caritatem disponsationis tuae quando secuta me es in deserto in terra quae non seminatur
JER|2|3|sanctus Israhel Domino primitiae frugum eius omnes qui devorant eum delinquunt mala venient super eos dicit Dominus
JER|2|4|audite verbum Domini domus Iacob et omnes cognationes domus Israhel
JER|2|5|haec dicit Dominus quid invenerunt patres vestri in me iniquitatis quia elongaverunt a me et ambulaverunt post vanitatem et vani facti sunt
JER|2|6|et non dixerunt ubi est Dominus qui ascendere nos fecit de terra Aegypti qui transduxit nos per desertum per terram inhabitabilem et inviam per terram sitis et imaginem mortis per terram in qua non ambulavit vir neque habitavit homo
JER|2|7|et induxi vos in terram Carmeli ut comederetis fructum eius et optima illius et ingressi contaminastis terram meam et hereditatem meam posuistis in abominationem
JER|2|8|sacerdotes non dixerunt ubi est Dominus et tenentes legem nescierunt me et pastores praevaricati sunt in me et prophetae prophetaverunt in Baal et idola secuti sunt
JER|2|9|propterea adhuc iudicio contendam vobiscum ait Dominus et cum filiis vestris disceptabo
JER|2|10|transite ad insulas Cetthim et videte et in Cedar mittite et considerate vehementer et videte si factum est huiuscemodi
JER|2|11|si mutavit gens deos et certe ipsi non sunt dii populus vero meus mutavit Gloriam suam in idolum
JER|2|12|obstupescite caeli super hoc et portae eius desolamini vehementer dicit Dominus
JER|2|13|duo enim mala fecit populus meus me dereliquerunt fontem aquae vivae ut foderent sibi cisternas cisternas dissipatas quae continere non valent aquas
JER|2|14|numquid servus est Israhel aut vernaculus quare ergo est factus in praedam
JER|2|15|super eum rugierunt leones et dederunt vocem suam posuerunt terram eius in solitudinem civitates eius exustae sunt et non est qui habitet in eis
JER|2|16|filii quoque Memfeos et Tafnes constupraverunt te usque ad verticem
JER|2|17|numquid non istud factum est tibi quia dereliquisti Dominum Deum tuum eo tempore quo ducebat te per viam
JER|2|18|et nunc quid tibi vis in via Aegypti ut bibas aquam turbidam et quid tibi cum via Assyriorum ut bibas aquam Fluminis
JER|2|19|arguet te malitia tua et aversio tua increpabit te scito et vide quia malum et amarum est reliquisse te Dominum Deum tuum et non esse timorem mei apud te dicit Dominus Deus exercituum
JER|2|20|a saeculo confregisti iugum meum rupisti vincula mea et dixisti non serviam in omni enim colle sublimi et sub omni ligno frondoso tu prosternebaris meretrix
JER|2|21|ego autem plantavi te vineam electam omne semen verum quomodo ergo conversa es in pravum vinea aliena
JER|2|22|si laveris te nitro et multiplicaveris tibi herbam borith maculata es in iniquitate tua coram me dicit Dominus Deus
JER|2|23|quomodo dicis non sum polluta post Baalim non ambulavi vide vias tuas in convalle scito quid feceris cursor levis explicans vias tuas
JER|2|24|onager adsuetus in solitudine in desiderio animae suae adtraxit ventum amoris sui nullus avertet eam omnes qui quaerunt eam non deficient in menstruis eius invenient eam
JER|2|25|prohibe pedem tuum a nuditate et guttur tuum a siti et dixisti desperavi nequaquam faciam adamavi quippe alienos et post eos ambulabo
JER|2|26|quomodo confunditur fur quando deprehenditur sic confusi sunt domus Israhel ipsi et reges eorum principes et sacerdotes et prophetae eorum
JER|2|27|dicentes ligno pater meus es tu et lapidi tu me genuisti verterunt ad me tergum et non faciem et in tempore adflictionis suae dicent surge et libera nos
JER|2|28|ubi sunt dii tui quos fecisti tibi surgant et liberent te in tempore adflictionis tuae secundum numerum quippe civitatum tuarum erant dii tui Iuda
JER|2|29|quid vultis mecum iudicio contendere omnes dereliquistis me dicit Dominus
JER|2|30|frustra percussi filios vestros disciplinam non receperunt devoravit gladius vester prophetas vestros quasi leo vastator
JER|2|31|generatio vestra videte verbum Domini numquid solitudo factus sum Israheli aut terra serotina quare ergo dixit populus meus recessimus non veniemus ultra ad te
JER|2|32|numquid obliviscitur virgo ornamenti sui sponsa fasciae pectoralis suae populus vero meus oblitus est mei diebus innumeris
JER|2|33|quid niteris bonam ostendere viam tuam ad quaerendam dilectionem quae insuper et malitias tuas docuisti vias tuas
JER|2|34|et in alis tuis inventus est sanguis animarum pauperum et innocentium non in fossis inveni eos sed in omnibus quae supra memoravi
JER|2|35|et dixisti absque peccato et innocens ego sum et propterea avertatur furor tuus a me ecce ego iudicio contendam tecum eo quod dixeris non peccavi
JER|2|36|quam vilis es facta nimis iterans vias tuas et ab Aegypto confunderis sicut confusa es ab Assur
JER|2|37|nam et ab ista egredieris et manus tuae erunt super caput tuum quoniam obtrivit Dominus confidentiam tuam et nihil habebis prosperum
JER|3|1|vulgo dicitur si dimiserit vir uxorem suam et recedens ab eo duxerit virum alterum numquid revertetur ad eam ultra numquid non polluta et contaminata erit mulier illa tu autem fornicata es cum amatoribus multis tamen revertere ad me dicit Dominus
JER|3|2|leva oculos tuos in directum et vide ubi non prostrata sis in viis sedebas expectans eos quasi latro in solitudine et polluisti terram in fornicationibus tuis et in malitiis tuis
JER|3|3|quam ob rem prohibitae sunt stillae pluviarum et serotinus imber non fuit frons mulieris meretricis facta est tibi noluisti erubescere
JER|3|4|ergo saltim amodo voca me pater meus dux virginitatis meae tu es
JER|3|5|numquid irasceris in perpetuum aut perseverabis in finem ecce locuta es et fecisti mala et potuisti
JER|3|6|et dixit Dominus ad me in diebus Iosiae regis numquid vidisti quae fecerit aversatrix Israhel abiit sibimet super omnem montem excelsum et sub omne lignum frondosum et fornicata est ibi
JER|3|7|et dixi cum fecisset haec omnia ad me convertere et non est reversa et vidit praevaricatrix soror eius Iuda
JER|3|8|quia pro eo quod moechata esset aversatrix Israhel dimisissem eam et dedissem ei libellum repudii et non timuit praevaricatrix Iuda soror eius sed abiit et fornicata est etiam ipsa
JER|3|9|et facilitate fornicationis suae contaminavit terram et moechata est cum lapide et cum ligno
JER|3|10|et in omnibus his non est reversa ad me praevaricatrix soror eius Iuda in toto corde suo sed in mendacio ait Dominus
JER|3|11|et dixit Dominus ad me iustificavit animam suam aversatrix Israhel conparatione praevaricatricis Iuda
JER|3|12|vade et clama sermones istos contra aquilonem et dices revertere aversatrix Israhel ait Dominus et non avertam faciem meam a vobis quia sanctus ego sum dicit Dominus et non irascar in perpetuum
JER|3|13|tamen scito iniquitatem tuam quia in Dominum Deum tuum praevaricata es et dispersisti vias tuas alienis sub omni ligno frondoso et vocem meam non audisti ait Dominus
JER|3|14|convertimini filii revertentes dicit Dominus quia ego vir vester et adsumam vos unum de civitate et duos de cognatione et introducam vos in Sion
JER|3|15|et dabo vobis pastores iuxta cor meum et pascent vos scientia et doctrina
JER|3|16|cumque multiplicati fueritis et creveritis in terra in diebus illis ait Dominus non dicent ultra arca testamenti Domini neque ascendet super cor neque recordabuntur illius nec visitabitur nec fiet ultra
JER|3|17|in tempore illo vocabunt Hierusalem solium Domini et congregabuntur ad eam omnes gentes in nomine Domini in Hierusalem et non ambulabunt post pravitatem cordis sui pessimi
JER|3|18|in diebus illis ibit domus Iuda ad domum Israhel et venient simul de terra aquilonis ad terram quam dedi patribus vestris
JER|3|19|ego autem dixi quomodo ponam te in filiis et tribuam tibi terram desiderabilem hereditatem praeclaram exercituum gentium et dixi patrem vocabis me et post me ingredi non cessabis
JER|3|20|sed quomodo si contemnat mulier amatorem suum sic contempsit me domus Israhel dicit Dominus
JER|3|21|vox in viis audita est ploratus et ululatus filiorum Israhel quoniam iniquam fecerunt viam suam obliti sunt Domini Dei sui
JER|3|22|convertimini filii revertentes et sanabo aversiones vestras ecce nos venimus ad te tu enim es Dominus Deus noster
JER|3|23|vere mendaces erant colles multitudo montium vere in Domino Deo nostro salus Israhel
JER|3|24|confusio comedit laborem patrum nostrorum ab adulescentia nostra greges eorum et armenta eorum filios eorum et filias eorum
JER|3|25|dormiemus in confusione nostra et operiet nos ignominia nostra quoniam Domino Deo nostro peccavimus nos et patres nostri ab adulescentia nostra usque ad hanc diem et non audivimus vocem Domini Dei nostri
JER|4|1|si converteris Israhel ait Dominus ad me convertere si abstuleris offendicula tua a facie mea non commoveberis
JER|4|2|et iurabis vivit Dominus in veritate et in iudicio et in iustitia et benedicent eum gentes ipsumque laudabunt
JER|4|3|haec enim dicit Dominus viro Iuda et Hierusalem novate vobis novale et nolite serere super spinas
JER|4|4|circumcidimini Domino et auferte praeputia cordium vestrorum vir Iuda et habitatores Hierusalem ne forte egrediatur ut ignis indignatio mea et succendatur et non sit qui extinguat propter malitiam cogitationum vestrarum
JER|4|5|adnuntiate in Iuda et in Hierusalem auditum facite loquimini et canite tuba in terra clamate fortiter dicite congregamini et ingrediamur civitates munitas
JER|4|6|levate signum in Sion confortamini nolite stare quia malum ego adduco ab aquilone et contritionem magnam
JER|4|7|ascendit leo de cubili suo et praedo gentium se levavit egressus est de loco suo ut ponat terram tuam in desolationem civitates tuae vastabuntur remanentes absque habitatore
JER|4|8|super hoc accingite vos ciliciis plangite et ululate quia non est aversa ira furoris Domini a nobis
JER|4|9|et erit in die illa dicit Dominus peribit cor regis et cor principum et obstupescent sacerdotes et prophetae consternabuntur
JER|4|10|et dixi heu heu heu Domine Deus ergone decepisti populum istum et Hierusalem dicens pax erit vobis et ecce pervenit gladius usque ad animam
JER|4|11|in tempore illo dicetur populo huic et Hierusalem ventus urens in viis quae sunt in deserto viae filiae populi mei non ad ventilandum et ad purgandum
JER|4|12|spiritus plenus ex his veniet mihi et nunc ego sed loquar iudicia mea cum eis
JER|4|13|ecce quasi nubes ascendet et quasi tempestas currus eius velociores aquilis equi illius vae nobis quoniam vastati sumus
JER|4|14|lava a malitia cor tuum Hierusalem ut salva fias usquequo morabuntur in te cogitationes noxiae
JER|4|15|vox enim adnuntiantis a Dan et notum facientis idolum de monte Ephraim
JER|4|16|concitate gentes ecce auditum est in Hierusalem custodes venire de terra longinqua et dare super civitates Iuda vocem suam
JER|4|17|quasi custodes agrorum facti sunt super eam in gyro quia me ad iracundiam provocavit ait Dominus
JER|4|18|viae tuae et cogitationes tuae fecerunt haec tibi ista malitia tua quia amara quia tetigit cor tuum
JER|4|19|ventrem meum ventrem meum doleo sensus cordis mei turbati sunt in me non tacebo quoniam vocem bucinae audivit anima mea clamorem proelii
JER|4|20|contritio super contritionem vocata est et vastata est omnis terra repente vastata sunt tabernacula mea subito pelles meae
JER|4|21|usquequo videbo fugientem audiam vocem bucinae
JER|4|22|quia stultus populus meus me non cognovit filii insipientes sunt et vecordes sapientes sunt ut faciant mala bene autem facere nescierunt
JER|4|23|aspexi terram et ecce vacua erat et nihili et caelos et non erat lux in eis
JER|4|24|vidi montes et ecce movebantur et omnes colles conturbati sunt
JER|4|25|intuitus sum et non erat homo et omne volatile caeli recessit
JER|4|26|aspexi et ecce Carmelus desertus et omnes urbes eius destructae sunt a facie Domini et a facie irae furoris eius
JER|4|27|haec enim dicit Dominus deserta erit omnis terra sed tamen consummationem non faciam
JER|4|28|lugebit terra et maerebunt caeli desuper eo quod locutus sum cogitavi et non paenituit me nec aversus sum ab eo
JER|4|29|a voce equitis et mittentis sagittam fugit omnis civitas ingressi sunt ardua et ascenderunt rupes universae urbes derelictae sunt et non habitat in eis homo
JER|4|30|tu autem vastata quid facies cum vestieris te coccino cum ornata fueris monili aureo et pinxeris stibio oculos tuos frustra conponeris contempserunt te amatores tui animam tuam quaerent
JER|4|31|vocem enim quasi parturientis audivi angustias ut puerperae vox filiae Sion intermorientis expandentisque manus suas vae mihi quia defecit anima mea propter interfectos
JER|5|1|circuite vias Hierusalem et aspicite et considerate et quaerite in plateis eius an inveniatis virum facientem iudicium et quaerentem fidem et propitius ero eius
JER|5|2|quod si etiam vivit Dominus dixerint et hoc falso iurabunt
JER|5|3|Domine oculi tui respiciunt fidem percussisti eos et non doluerunt adtrivisti eos et rennuerunt accipere disciplinam induraverunt facies suas super petram noluerunt reverti
JER|5|4|ego autem dixi forsitan pauperes sunt et stulti ignorantes viam Domini iudicium Dei sui
JER|5|5|ibo igitur ad optimates et loquar eis ipsi enim cognoverunt viam Domini iudicium Dei sui et ecce magis hii simul confregerunt iugum ruperunt vincula
JER|5|6|idcirco percussit eos leo de silva lupus ad vesperam vastavit eos pardus vigilans super civitates eorum omnis qui egressus fuerit ex eis capietur quia multiplicatae sunt praevaricationes eorum confortatae sunt aversiones eorum
JER|5|7|super quo propitius tibi esse potero filii tui dereliquerunt me et iurant in his qui non sunt dii saturavi eos et moechati sunt et in domo meretricis luxuriabantur
JER|5|8|equi amatores et admissarii facti sunt unusquisque ad uxorem proximi sui hinniebat
JER|5|9|numquid super his non visitabo dicit Dominus et in gente tali non ulciscetur anima mea
JER|5|10|ascendite muros eius et dissipate consummationem autem nolite facere auferte propagines eius quia non sunt Domini
JER|5|11|praevaricatione enim praevaricata est in me domus Israhel et domus Iuda ait Dominus
JER|5|12|negaverunt Dominum et dixerunt non est ipse neque veniet super nos malum gladium et famem non videbimus
JER|5|13|prophetae fuerunt in ventum et responsum non fuit in eis haec ergo evenient illis
JER|5|14|haec dicit Dominus Deus exercituum quia locuti estis verbum istud ecce ego do verba mea in ore tuo in ignem et populum istum ligna et vorabit eos
JER|5|15|ecce ego adducam super vos gentem de longinquo domus Israhel ait Dominus gentem robustam gentem antiquam gentem cuius ignorabis linguam nec intelleges quid loquatur
JER|5|16|faretra eius quasi sepulchrum patens universi fortes
JER|5|17|et comedet segetes tuas et panem tuum devorabit filios tuos et filias tuas comedet gregem tuum et armenta tua comedet vineam tuam et ficum tuam et conteret urbes munitas tuas in quibus tu habes fiduciam gladio
JER|5|18|verumtamen et diebus illis ait Dominus non faciam vos in consummationem
JER|5|19|quod si dixeritis quare fecit Dominus Deus noster nobis haec omnia dices ad eos sicut dereliquistis me et servistis deo alieno in terra vestra sic servietis alienis in terra non vestra
JER|5|20|adnuntiate hoc domui Iacob et auditum facite in Iuda dicentes
JER|5|21|audi populus stulte qui non habes cor qui habentes oculos non videtis et aures et non auditis
JER|5|22|me ergo non timebitis ait Dominus et a facie mea non dolebitis qui posui harenam terminum mari praeceptum sempiternum quod non praeteribit et commovebuntur et non poterunt et intumescent fluctus eius et non transibunt illud
JER|5|23|populo autem huic factum est cor incredulum et exasperans recesserunt et abierunt
JER|5|24|et non dixerunt in corde suo metuamus Dominum Deum nostrum qui dat nobis pluviam temporaneam et serotinam in tempore suo plenitudinem annuae messis custodientem nobis
JER|5|25|iniquitates nostrae declinaverunt haec et peccata nostra prohibuerunt bonum a nobis
JER|5|26|quia inventi sunt in populo meo impii insidiantes quasi aucupes laqueos ponentes et pedicas ad capiendos viros
JER|5|27|sicut decipula plena avibus sic domus eorum plenae dolo ideo magnificati sunt et ditati
JER|5|28|incrassati sunt et inpinguati et praeterierunt sermones meos pessime causam non iudicaverunt causam pupilli non direxerunt et iudicium pauperum non iudicaverunt
JER|5|29|numquid super his non visitabo dicit Dominus aut super gentem huiuscemodi non ulciscetur anima mea
JER|5|30|stupor et mirabilia facta sunt in terra
JER|5|31|prophetae prophetabant mendacium et sacerdotes adplaudebant manibus suis et populus meus dilexit talia quid igitur fiet in novissimo eius
JER|6|1|confortamini filii Beniamin in medio Hierusalem et in Thecua clangite bucina et super Bethaccharem levate vexillum quia malum visum est ab aquilone et contritio magna
JER|6|2|speciosae et delicatae adsimilavi filiam Sion
JER|6|3|ad eam venient pastores et greges eorum fixerunt in ea tentoria in circuitu pascet unusquisque eos qui sub manu sua sunt
JER|6|4|sanctificate super eam bellum consurgite et ascendamus in meridie vae nobis quia declinavit dies quia longiores factae sunt umbrae vesperi
JER|6|5|surgite et ascendamus in nocte et dissipemus domos eius
JER|6|6|quia haec dicit Dominus exercituum caedite lignum eius et fundite circa Hierusalem aggerem haec est civitas visitationis omnis calumnia in medio eius
JER|6|7|sicut frigidam facit cisterna aquam suam sic frigidam fecit malitiam suam iniquitas et vastitas audietur in ea coram me semper infirmitas et plaga
JER|6|8|erudire Hierusalem ne forte recedat anima mea a te ne forte ponam te desertam terram inhabitabilem
JER|6|9|haec dicit Dominus exercituum usque ad racemum colligent quasi in vinea reliquias Israhel converte manum tuam quasi vindemiator ad cartallum
JER|6|10|cui loquar et quem contestabor ut audiant ecce incircumcisae aures eorum et audire non possunt ecce verbum Domini factum est eis in obprobrium et non suscipient illud
JER|6|11|idcirco furore Domini plenus sum laboravi sustinens effunde super parvulum foris et super concilium iuvenum simul vir enim cum muliere capietur senex cum pleno dierum
JER|6|12|et transibunt domus eorum ad alteros agri et uxores pariter quia extendam manum meam super habitantes terram dicit Dominus
JER|6|13|a minore quippe usque ad maiorem omnes avaritiae student et a propheta usque ad sacerdotem cuncti faciunt dolum
JER|6|14|et curabant contritionem filiae populi mei cum ignominia dicentes pax pax et non erat pax
JER|6|15|confusi sunt quia abominationem fecerunt quin potius confusione non sunt confusi et erubescere nescierunt quam ob rem cadent inter ruentes in tempore visitationis suae corruent dicit Dominus
JER|6|16|haec dicit Dominus state super vias et videte et interrogate de semitis antiquis quae sit via bona et ambulate in ea et invenietis refrigerium animabus vestris et dixerunt non ambulabimus
JER|6|17|et constitui super vos speculatores audite vocem tubae et dixerunt non audiemus
JER|6|18|ideo audite gentes et cognosce congregatio quanta ego faciam eis
JER|6|19|audi terra ecce ego adducam mala super populum istum fructum cogitationum eius quia verba mea non audierunt et legem meam proiecerunt
JER|6|20|ut quid mihi tus de Saba adfertis et calamum suave olentem de terra longinqua holocaustomata vestra non sunt accepta et victimae vestrae non placuerunt mihi
JER|6|21|propterea haec dicit Dominus ecce ego dabo in populum istum ruinas et ruent in eis patres et filii simul vicinus et proximus et peribunt
JER|6|22|haec dicit Dominus ecce populus venit de terra aquilonis et gens magna consurget a finibus terrae
JER|6|23|sagittam et scutum arripiet crudelis est et non miserebitur vox eius quasi mare sonabit et super equos ascendent praeparati quasi vir ad proelium adversum te filia Sion
JER|6|24|audivimus famam eius dissolutae sunt manus nostrae tribulatio adprehendit nos dolores ut parturientem
JER|6|25|nolite exire ad agros et in via ne ambuletis quoniam gladius inimici pavor in circuitu
JER|6|26|filia populi mei accingere cilicio et conspergere cinere luctum unigeniti fac tibi planctum amarum quia repente veniet vastator super nos
JER|6|27|probatorem dedi te in populo meo robustum et scies et probabis viam eorum
JER|6|28|omnes isti principes declinantum ambulantes fraudulenter aes et ferrum universi corrupti sunt
JER|6|29|defecit sufflatorium in igne consumptum est plumbum frustra conflavit conflator malitiae enim eorum non sunt consumptae
JER|6|30|argentum reprobum vocate eos quia Dominus proiecit illos
JER|7|1|verbum quod factum est ad Hieremiam a Domino dicens
JER|7|2|sta in porta domus Domini et praedica ibi verbum istud et dic audite verbum Domini omnis Iuda qui ingredimini per portas has ut adoretis Dominum
JER|7|3|haec dicit Dominus exercituum Deus Israhel bonas facite vias vestras et studia vestra et habitabo vobiscum in loco isto
JER|7|4|nolite confidere in verbis mendacii dicentes templum Domini templum Domini templum Domini est
JER|7|5|quoniam si bene direxeritis vias vestras et studia vestra si feceritis iudicium inter virum et proximum eius
JER|7|6|advenae et pupillo et viduae non feceritis calumniam nec sanguinem innocentem effuderitis in loco hoc et post deos alienos non ambulaveritis in malum vobismet ipsis
JER|7|7|habitabo vobiscum in loco isto in terra quam dedi patribus vestris a saeculo usque in saeculum
JER|7|8|ecce vos confiditis vobis in sermonibus mendacii qui non proderunt vobis
JER|7|9|furari occidere adulterare iurare mendaciter libare Baali et ire post deos alienos quos ignoratis
JER|7|10|et venistis et stetistis coram me in domo hac in qua invocatum est nomen meum et dixistis liberati sumus eo quod fecerimus omnes abominationes istas
JER|7|11|ergo spelunca latronum facta est domus ista in qua invocatum est nomen meum in oculis vestris ego ego sum ego vidi dicit Dominus
JER|7|12|ite ad locum meum in Silo ubi habitavit nomen meum a principio et videte quae fecerim ei propter malitiam populi mei Israhel
JER|7|13|et nunc quia fecistis omnia opera haec dicit Dominus et locutus sum ad vos mane consurgens et loquens et non audistis et vocavi vos et non respondistis
JER|7|14|faciam domui huic in qua invocatum est nomen meum et in qua vos habetis fiduciam et loco quem dedi vobis et patribus vestris sicut feci Silo
JER|7|15|et proiciam vos a facie mea sicut proieci omnes fratres vestros universum semen Ephraim
JER|7|16|tu ergo noli orare pro populo hoc nec adsumas pro eis laudem et orationem et non obsistas mihi quia non exaudiam te
JER|7|17|nonne vides quid isti faciant in civitatibus Iuda et in plateis Hierusalem
JER|7|18|filii colligunt ligna et patres succendunt ignem et mulieres conspergunt adipem ut faciant placentas Reginae caeli et libent diis alienis et me ad iracundiam provocent
JER|7|19|numquid me ad iracundiam provocant dicit Dominus nonne semet ipsos in confusionem vultus sui
JER|7|20|ideo haec dicit Dominus Deus ecce furor meus et indignatio mea conflatur super locum istum super viros et super iumenta et super lignum regionis et super fruges terrae et succendetur et non extinguetur
JER|7|21|haec dicit Dominus exercituum Deus Israhel holocaustomata vestra addite victimis vestris et comedite carnes
JER|7|22|quia non sum locutus cum patribus vestris et non praecepi eis in die qua eduxi eos de terra Aegypti de verbo holocaustomatum et victimarum
JER|7|23|sed hoc verbum praecepi eis dicens audite vocem meam et ero vobis Deus et vos eritis mihi populus et ambulate in omni via quam mandavi vobis ut bene sit vobis
JER|7|24|et non audierunt nec inclinaverunt aurem suam sed abierunt in voluntatibus et pravitate cordis sui mali factique sunt retrorsum et non in ante
JER|7|25|a die qua egressi sunt patres eorum de terra Aegypti usque ad diem hanc et misi ad vos omnes servos meos prophetas per diem consurgens diluculo et mittens
JER|7|26|et non audierunt me nec inclinaverunt aurem suam sed induraverunt cervicem et peius operati sunt quam patres eorum
JER|7|27|et loqueris ad eos omnia verba haec et non audient te et vocabis eos et non respondebunt tibi
JER|7|28|et dices ad eos haec est gens quae non audivit vocem Domini Dei sui nec recepit disciplinam periit fides et ablata est de ore eorum
JER|7|29|tonde capillum tuum et proice et sume in directum planctum quia proiecit Dominus et reliquit generationem furoris sui
JER|7|30|quia fecerunt filii Iuda malum in oculis meis dicit Dominus posuerunt offendicula sua in domo in qua invocatum est nomen meum ut polluerent eam
JER|7|31|et aedificaverunt excelsa Thofeth qui est in valle filii Ennom ut incenderent filios suos et filias suas igni quae non praecepi nec cogitavi in corde meo
JER|7|32|ideo ecce dies venient dicit Dominus et non dicetur amplius Thofeth et vallis filii Ennom sed vallis Interfectionis et sepelient in Thofeth eo quod non sit locus
JER|7|33|et erit morticinum populi huius in cibum volucribus caeli et bestiis terrae et non erit qui abigat
JER|7|34|et quiescere faciam de urbibus Iuda et de plateis Hierusalem vocem gaudii et vocem laetitiae vocem sponsi et vocem sponsae in desolatione enim erit terra
JER|8|1|in tempore illo ait Dominus eicient ossa regis Iuda et ossa principum eius et ossa sacerdotum et ossa prophetarum et ossa eorum qui habitaverunt Hierusalem de sepulchris suis
JER|8|2|et pandent ea ad solem et lunam et omnem militiam caeli quae dilexerunt et quibus servierunt et post quae ambulaverunt et quae quaesierunt et adoraverunt non colligentur et non sepelientur in sterquilinium super faciem terrae erunt
JER|8|3|et eligent magis mortem quam vitam omnes qui residui fuerint de cognatione hac pessima in universis locis quae derelicta sunt ad quae eieci eos dicit Dominus exercituum
JER|8|4|et dices ad eos haec dicit Dominus numquid qui cadet non resurget et qui aversus est non revertetur
JER|8|5|quare ergo aversus est populus iste in Hierusalem aversione contentiosa adprehenderunt mendacium et noluerunt reverti
JER|8|6|adtendi et auscultavi nemo quod bonum est loquitur nullus est qui agat paenitentiam super peccato suo dicens quid feci omnes conversi sunt ad cursum suum quasi equus impetu vadens in proelio
JER|8|7|milvus in caelo cognovit tempus suum turtur et hirundo et ciconia custodierunt tempus adventus sui populus autem meus non cognovit iudicium Domini
JER|8|8|quomodo dicitis sapientes nos sumus et lex Domini nobiscum est vere mendacium operatus est stilus mendax scribarum
JER|8|9|confusi sunt sapientes perterriti et capti sunt verbum enim Domini proiecerunt et sapientia nulla est in eis
JER|8|10|propterea dabo mulieres eorum exteris agros eorum heredibus quia a minimo usque ad maximum omnes avaritiam sequuntur a propheta usque ad sacerdotem cuncti faciunt mendacium
JER|8|11|et sanabant contritionem filiae populi mei ad ignominiam dicentes pax pax cum non esset pax
JER|8|12|confusi sunt quia abominationem fecerunt quinimmo confusione non sunt confusi et erubescere nescierunt idcirco cadent inter corruentes in tempore visitationis suae corruent dicit Dominus
JER|8|13|congregans congregabo eos ait Dominus non est uva in vitibus et non sunt ficus in ficulnea folium defluxit et dedi eis quae praetergressa sunt
JER|8|14|quare sedemus convenite et ingrediamur civitatem munitam et sileamus ibi quia Dominus noster silere nos fecit et potum dedit nobis aquam fellis peccavimus enim Domino
JER|8|15|expectavimus pacem et non erat bonum tempus medellae et ecce formido
JER|8|16|a Dan auditus est fremitus equorum eius a voce hinnituum pugnatorum eius commota est omnis terra et venerunt et devoraverunt terram et plenitudinem eius urbem et habitatores eius
JER|8|17|quia ecce ego mittam vobis serpentes regulos quibus non est incantatio et mordebunt vos ait Dominus
JER|8|18|dolor meus super dolorem in me cor meum maerens
JER|8|19|ecce vox clamoris filiae populi mei de terra longinqua numquid Dominus non est in Sion aut rex eius non est in ea quare ergo me ad iracundiam concitaverunt in sculptilibus suis et in vanitatibus alienis
JER|8|20|transiit messis finita est aestas et nos salvati non sumus
JER|8|21|super contritionem filiae populi mei contritus sum et contristatus stupor obtinuit me
JER|8|22|numquid resina non est in Galaad aut medicus non est ibi quare igitur non est obducta cicatrix filiae populi mei
JER|9|1|quis dabit capiti meo aquam et oculis meis fontem lacrimarum et plorabo die et nocte interfectos filiae populi mei
JER|9|2|quis dabit me in solitudine diversorium viatorum et derelinquam populum meum et recedam ab eis quia omnes adulteri sunt coetus praevaricatorum
JER|9|3|et extenderunt linguam suam quasi arcum mendacii et non veritatis confortati sunt in terra quia de malo ad malum egressi sunt et me non cognoverunt dicit Dominus
JER|9|4|unusquisque se a proximo suo custodiat et in omni fratre suo non habeat fiduciam quia omnis frater subplantans subplantabit et omnis amicus fraudulenter incedet
JER|9|5|et vir fratrem suum deridebit et veritatem non loquentur docuerunt enim linguam suam loqui mendacium ut inique agerent laboraverunt
JER|9|6|habitatio tua in medio doli in dolo rennuerunt scire me dicit Dominus
JER|9|7|propterea haec dicit Dominus exercituum ecce ego conflabo et probabo eos quid enim aliud faciam a facie filiae populi mei
JER|9|8|sagitta vulnerans lingua eorum dolum locuta est in ore suo pacem cum amico suo loquitur et occulte ponit ei insidias
JER|9|9|numquid super his non visitabo dicit Dominus aut in gentem huiuscemodi non ulciscetur anima mea
JER|9|10|super montes adsumam fletum ac lamentum et super speciosa deserti planctum quoniam incensa sunt eo quod non sit vir pertransiens et non audierunt vocem possidentis a volucre caeli usque ad pecora transmigraverunt et recesserunt
JER|9|11|et dabo Hierusalem in acervos harenae et cubilia draconum et civitates Iuda dabo in desolationem eo quod non sit habitator
JER|9|12|quis est vir sapiens qui intellegat hoc et ad quem verbum oris Domini fiat ut adnuntiet istud quare perierit terra exusta sit quasi desertum eo quod non sit qui pertranseat
JER|9|13|et dixit Dominus quia dereliquerunt legem meam quam dedi eis et non audierunt vocem meam et non ambulaverunt in ea
JER|9|14|et abierunt post pravitatem cordis sui et post Baalim quos didicerunt a patribus suis
JER|9|15|idcirco haec dicit Dominus exercituum Deus Israhel ecce ego cibabo eos populum istum absinthio et potum dabo eis aquam fellis
JER|9|16|et dispergam eos in gentibus quas non noverunt ipsi et patres eorum et mittam post eos gladium donec consumantur
JER|9|17|haec dicit Dominus exercituum contemplamini et vocate lamentatrices et veniant et ad eas quae sapientes sunt mittite et properent
JER|9|18|festinent et adsumant super nos lamentum deducant oculi nostri lacrimas et palpebrae nostrae defluant aquis
JER|9|19|quia vox lamentationis audita est de Sion quomodo vastati sumus et confusi vehementer quia dereliquimus terram quoniam deiecta sunt tabernacula nostra
JER|9|20|audite ergo mulieres verbum Domini et adsumat auris vestra sermonem oris eius et docete filias vestras lamentum et unaquaeque proximam suam planctum
JER|9|21|quia ascendit mors per fenestras nostras ingressa est domos nostras disperdere parvulos de foris iuvenes de plateis
JER|9|22|loquere haec dicit Dominus et cadet morticinum hominis quasi stercus super faciem regionis et quasi faenum post tergum metentis et non est qui colligat
JER|9|23|haec dicit Dominus non glorietur sapiens in sapientia sua et non glorietur fortis in fortitudine sua et non glorietur dives in divitiis suis
JER|9|24|sed in hoc glorietur qui gloriatur scire et nosse me quia ego sum Dominus qui facio misericordiam et iudicium et iustitiam in terra haec enim placent mihi ait Dominus
JER|9|25|ecce dies veniunt dicit Dominus et visitabo super omnem qui circumcisum habet praeputium
JER|9|26|super Aegyptum et super Iudam et super Edom et super filios Ammon et super Moab et super omnes qui adtonsi sunt in comam habitantes in deserto quia omnes gentes habent praeputium omnis autem domus Israhel incircumcisi sunt corde
JER|10|1|audite verbum quod locutus est Dominus super vos domus Israhel
JER|10|2|haec dicit Dominus iuxta vias gentium nolite discere et a signis caeli nolite metuere quae timent gentes
JER|10|3|quia leges populorum vanae sunt quia lignum de saltu praecidit opus manuum artificis in ascia
JER|10|4|argento et auro decoravit illud clavis et malleis conpegit ut non dissolvatur
JER|10|5|in similitudinem palmae fabricata sunt et non loquentur portata tollentur quia incedere non valent nolite ergo timere ea quia nec male possunt facere nec bene
JER|10|6|non est similis tui Domine magnus tu et magnum nomen tuum in fortitudine
JER|10|7|quis non timebit te o rex gentium tuum est enim decus inter cunctos sapientes gentium et in universis regnis eorum nullus est similis tui
JER|10|8|pariter insipientes et fatui probabuntur doctrina vanitatis eorum lignum est
JER|10|9|argentum involutum de Tharsis adfertur et aurum de Ofaz opus artificis et manus aerarii hyacinthus et purpura indumentum eorum opus artificum universa haec
JER|10|10|Dominus autem Deus verus est ipse Deus vivens et rex sempiternus ab indignatione eius commovebitur terra et non sustinebunt gentes comminationem eius
JER|10|11|sic ergo dicetis eis dii qui caelos et terram non fecerunt pereant de terra et de his quae sub caelis sunt
JER|10|12|qui facit terram in fortitudine sua praeparat orbem in sapientia sua et prudentia sua extendit caelos
JER|10|13|ad vocem suam dat multitudinem aquarum in caelo et elevat nebulas ab extremitatibus terrae fulgura in pluviam facit et educit ventum de thesauris suis
JER|10|14|stultus factus est omnis homo ab scientia confusus est omnis artifex in sculptili quoniam falsum est quod conflavit et non est spiritus in eis
JER|10|15|vana sunt et opus risu dignum in tempore visitationis suae peribunt
JER|10|16|non est his similis pars Iacob qui enim formavit omnia ipse est et Israhel virga hereditatis eius Dominus exercituum nomen illi
JER|10|17|congrega de terra confusionem tuam quae habitas in obsidione
JER|10|18|quia haec dicit Dominus ecce ego longe proiciam habitatores terrae in hac vice et tribulabo eos ita ut inveniantur
JER|10|19|vae mihi super contritione mea pessima plaga mea ego autem dixi plane haec infirmitas mea est et portabo illam
JER|10|20|tabernaculum meum vastatum est omnes funiculi mei disrupti sunt filii mei exierunt a me et non subsistunt non est qui extendat ultra tentorium meum et erigat pelles meas
JER|10|21|quia stulte egerunt pastores et Dominum non quaesierunt propterea non intellexerunt et omnis grex eorum dispersus est
JER|10|22|vox auditionis ecce venit et commotio magna de terra aquilonis ut ponat civitates Iuda solitudinem et habitaculum draconum
JER|10|23|scio Domine quia non est hominis via eius nec viri est ut ambulet et dirigat gressus suos
JER|10|24|corripe me Domine verumtamen in iudicio et non in furore tuo ne forte ad nihilum redigas me
JER|10|25|effunde indignationem tuam super gentes quae non cognoverunt te et super provincias quae nomen tuum non invocaverunt quia comederunt Iacob et devoraverunt eum et consumpserunt illum et decus eius dissipaverunt
JER|11|1|verbum quod factum est ad Hieremiam a Domino dicens
JER|11|2|audite verba pacti huius et loquimini ad viros Iuda et habitatores Hierusalem
JER|11|3|et dices ad eos haec dicit Dominus Deus Israhel maledictus vir qui non audierit verba pacti huius
JER|11|4|quod praecepi patribus vestris in die qua eduxi eos de terra Aegypti de fornace ferrea dicens audite vocem meam et facite omnia quae praecipio vobis et eritis mihi in populum et ego ero vobis in Deum
JER|11|5|ut suscitem iuramentum quod iuravi patribus vestris daturum me eis terram fluentem lacte et melle sicut est dies haec et respondi et dixi amen Domine
JER|11|6|et dixit Dominus ad me vociferare omnia verba haec in civitatibus Iuda et foris Hierusalem dicens audite verba pacti huius et facite illa
JER|11|7|quia contestans contestatus sum patres vestros in die qua eduxi eos de terra Aegypti usque ad diem hanc mane surgens contestatus sum et dixi audite vocem meam
JER|11|8|et non audierunt nec inclinaverunt aurem suam sed abierunt unusquisque in pravitate cordis sui mali et induxi super eos omnia verba pacti huius quod praecepi ut facerent et non fecerunt
JER|11|9|et dixit Dominus ad me inventa est coniuratio in viris Iuda et in habitatoribus Hierusalem
JER|11|10|reversi sunt ad iniquitates patrum suorum priores qui noluerunt audire verba mea et hii ergo abierunt post deos alienos ut servirent eis irritum fecerunt domus Israhel et domus Iuda pactum meum quod pepigi cum patribus eorum
JER|11|11|quam ob rem haec dicit Dominus ecce ego inducam super eos mala de quibus exire non poterunt et clamabunt ad me et non exaudiam eos
JER|11|12|et ibunt civitates Iuda et habitatores Hierusalem et clamabunt ad deos quibus libant et non salvabunt eos in tempore adflictionis eorum
JER|11|13|secundum numerum enim civitatum tuarum erant dii tui Iuda et secundum numerum viarum Hierusalem posuistis aras confusionis aras ad libandum Baali
JER|11|14|tu ergo noli orare pro populo hoc et ne adsumas pro eis laudem et orationem quia non exaudiam in tempore clamoris eorum ad me in tempore adflictionis eorum
JER|11|15|quid est quod dilectus meus in domo mea fecit scelera multa numquid carnes sanctae auferent a te malitias tuas in quibus gloriata es
JER|11|16|olivam uberem pulchram fructiferam speciosam vocavit Dominus nomen tuum ad vocem loquellae grandis exarsit ignis in ea et conbusta sunt frutecta eius
JER|11|17|et Dominus exercituum qui plantavit te locutus est super te malum pro malis domus Israhel et domus Iuda quae fecerunt sibi ad inritandum me libantes Baali
JER|11|18|tu autem Domine demonstrasti mihi et cognovi tunc ostendisti mihi studia eorum
JER|11|19|et ego quasi agnus mansuetus qui portatur ad victimam et non cognovi quia super me cogitaverunt consilia mittamus lignum in panem eius et eradamus eum de terra viventium et nomen eius non memoretur amplius
JER|11|20|tu autem Domine Sabaoth qui iudicas iuste et probas renes et cor videam ultionem tuam ex eis tibi enim revelavi causam meam
JER|11|21|propterea haec dicit Dominus ad viros Anathoth qui quaerunt animam tuam et dicunt non prophetabis in nomine Domini et non morieris in manibus nostris
JER|11|22|propterea haec dicit Dominus exercituum ecce ego visitabo super eos iuvenes morientur in gladio filii eorum et filiae eorum morientur in fame
JER|11|23|et reliquiae non erunt ex eis inducam enim malum super viros Anathoth annum visitationis eorum
JER|12|1|iustus quidem tu es Domine si disputem tecum verumtamen iusta loquar ad te quare via impiorum prosperatur bene est omnibus qui praevaricantur et inique agunt
JER|12|2|plantasti eos et radicem miserunt proficiunt et faciunt fructum prope es tu ori eorum et longe a renibus eorum
JER|12|3|et tu Domine nosti me vidisti me et probasti cor meum tecum congrega eos quasi gregem ad victimam et sanctifica eos in die occisionis
JER|12|4|usquequo lugebit terra et herba omnis regionis siccabitur propter malitiam habitantium in ea consumptum est animal et volucre quoniam dixerunt non videbit novissima nostra
JER|12|5|si cum peditibus currens laborasti quomodo contendere poteris cum equis cum autem in terra pacis secura fueris quid facies in superbia Iordanis
JER|12|6|nam et fratres tui et domus patris tui etiam ipsi pugnaverunt adversum te et clamaverunt post te plena voce ne credas eis cum locuti fuerint tibi bona
JER|12|7|reliqui domum meam dimisi hereditatem meam dedi dilectam animam meam in manu inimicorum eius
JER|12|8|facta est mihi hereditas mea quasi leo in silva dedit contra me vocem ideo odivi eam
JER|12|9|numquid avis discolor hereditas mea mihi numquid avis tincta per totum venite congregamini omnes bestiae terrae properate ad devorandum
JER|12|10|pastores multi demoliti sunt vineam meam conculcaverunt partem meam dederunt portionem meam desiderabilem in desertum solitudinis
JER|12|11|posuerunt eam in dissipationem luxitque super me desolatione desolata est omnis terra quia nullus est qui recogitet corde
JER|12|12|super omnes vias deserti venerunt vastatores quia gladius Domini devoravit ab extremo terrae usque ad extremum eius non est pax universae carni
JER|12|13|seminaverunt triticum et spinas messuerunt hereditatem acceperunt et non eis proderit confundemini a fructibus vestris propter iram furoris Domini
JER|12|14|haec dicit Dominus adversum omnes vicinos meos pessimos qui tangunt hereditatem quam distribui populo meo Israhel ecce ego evellam eos de terra eorum et domum Iuda evellam de medio eorum
JER|12|15|et cum evellero eos convertar et miserebor eorum et reducam eos virum ad hereditatem suam et virum in terram suam
JER|12|16|et erit si eruditi didicerint vias populi mei ut iurent in nomine meo vivit Dominus sicut docuerunt populum meum iurare in Baal aedificabuntur in medio populi mei
JER|12|17|quod si non audierint evellam gentem illam evulsione et perditione ait Dominus
JER|13|1|haec dicit Dominus ad me vade et posside tibi lumbare lineum et pones illud super lumbos tuos et in aquam non inferes illud
JER|13|2|et possedi lumbare iuxta verbum Domini et posui circa lumbos meos
JER|13|3|et factus est sermo Domini ad me secundo dicens
JER|13|4|tolle lumbare quod possedisti quod est circa lumbos tuos et surgens vade ad Eufraten et absconde illud ibi in foramine petrae
JER|13|5|et abii et abscondi illud in Eufraten sicut praeceperat mihi Dominus
JER|13|6|et factum est post dies plurimos dixit Dominus ad me surge vade ad Eufraten et tolle inde lumbare quod praecepi tibi ut absconderes illud ibi
JER|13|7|et abii ad Eufraten et fodi et tuli lumbare de loco ubi absconderam illud et ecce conputruerat lumbare ita ut nullo usui aptum esset
JER|13|8|et factum est verbum Domini ad me dicens
JER|13|9|haec dicit Dominus sic putrescere faciam superbiam Iuda et superbiam Hierusalem multam
JER|13|10|populum istum pessimum qui nolunt audire verba mea et ambulant in pravitate cordis sui abieruntque post deos alienos ut servirent eis et adorarent eos et erunt sicut lumbare istud quod nullo usui aptum est
JER|13|11|sicut enim adheret lumbare ad lumbos viri sic adglutinavi mihi omnem domum Israhel et omnem domum Iuda dicit Dominus ut esset mihi in populum et in nomen et in laudem et in gloriam et non audierunt
JER|13|12|dices ergo ad eos sermonem istum haec dicit Dominus Deus Israhel omnis laguncula implebitur vino et dicent ad te numquid ignoramus quia omnis laguncula implebitur vino
JER|13|13|et dices ad eos haec dicit Dominus ecce ego implebo omnes habitatores terrae huius et reges qui sedent de stirpe David super thronum eius et sacerdotes et prophetas et omnes habitatores Hierusalem ebrietate
JER|13|14|et dispergam eos virum a fratre suo et patres et filios pariter ait Dominus non parcam et non concedam neque miserebor ut non disperdam eos
JER|13|15|audite et auribus percipite nolite elevari quia Dominus locutus est
JER|13|16|date Domino Deo vestro gloriam antequam contenebrescat et antequam offendant pedes vestri ad montes caligosos expectabitis lucem et ponet eam in umbram mortis et in caliginem
JER|13|17|quod si hoc non audieritis in abscondito plorabit anima mea a facie superbiae plorans plorabit et deducet oculus meus lacrimam quia captus est grex Domini
JER|13|18|dic regi et dominatrici humiliamini sedete quoniam descendit de capite vestro corona gloriae vestrae
JER|13|19|civitates austri clausae sunt et non est qui aperiat translata est omnis Iudaea transmigratione perfecta
JER|13|20|levate oculos vestros et videte qui venitis ab aquilone ubi est grex qui datus est tibi pecus inclitum tuum
JER|13|21|quid dices cum visitaverit te tu enim docuisti eos adversum te et erudisti in caput tuum numquid non dolores adprehendent te quasi mulierem parturientem
JER|13|22|quod si dixeris in corde tuo quare venerunt mihi haec propter multitudinem iniquitatis tuae revelata sunt verecundiora tua pollutae sunt plantae tuae
JER|13|23|si mutare potest Aethiops pellem suam aut pardus varietates suas et vos poteritis bene facere cum didiceritis malum
JER|13|24|et disseminabo eos quasi stipulam quae vento raptatur in deserto
JER|13|25|haec sors tua parsque mensurae tuae a me dicit Dominus quia oblita es mei et confisa es in mendacio
JER|13|26|unde et ego nudavi femora tua contra faciem tuam et apparuit ignominia tua
JER|13|27|adulteria tua et hinnitus tuus scelus fornicationis tuae super colles in agro vidi abominationes tuas vae tibi Hierusalem non mundaberis post me usquequo adhuc
JER|14|1|quod factum est verbum Domini ad Hieremiam de sermonibus siccitatis
JER|14|2|luxit Iudaea et portae eius corruerunt et obscuratae sunt in terra et clamor Hierusalem ascendit
JER|14|3|maiores miserunt minores suos ad aquam venerunt ad hauriendum non invenerunt aquam reportaverunt vasa sua vacua confusi sunt et adflicti et operuerunt capita sua
JER|14|4|propter terrae vastitatem quia non venit pluvia in terra confusi sunt agricolae operuerunt capita sua
JER|14|5|nam et cerva in agro peperit et reliquit quia non erat herba
JER|14|6|et onagri steterunt in rupibus traxerunt ventum quasi dracones defecerunt oculi eorum quia non erat herba
JER|14|7|si iniquitates nostrae responderunt nobis Domine fac propter nomen tuum quoniam multae sunt aversiones nostrae tibi peccavimus
JER|14|8|expectatio Israhel salvator eius in tempore tribulationis quare quasi colonus futurus es in terra et quasi viator declinans ad manendum
JER|14|9|quare futurus es velut vir vagus ut fortis qui non potest salvare tu autem in nobis es Domine et nomen tuum super nos invocatum est ne derelinquas nos
JER|14|10|haec dicit Dominus populo huic qui dilexit movere pedes suos et non quievit et Domino non placuit nunc recordabitur iniquitatum eorum et visitabit peccata eorum
JER|14|11|et dixit Dominus ad me noli orare pro populo isto in bonum
JER|14|12|cum ieiunaverint non exaudiam preces eorum et si obtulerint holocaustomata et victimas non suscipiam ea quoniam gladio et fame et peste ego consumam eos
JER|14|13|et dixi a a a Domine Deus prophetae dicunt eis non videbitis gladium et famis non erit in vobis sed pacem veram dabit vobis in loco isto
JER|14|14|et dixit Dominus ad me falso prophetae vaticinantur in nomine meo non misi eos et non praecepi eis neque locutus sum ad eos visionem mendacem et divinationem et fraudulentiam et seductionem cordis sui prophetant vobis
JER|14|15|ideo haec dicit Dominus de prophetis qui prophetant in nomine meo quos ego non misi dicentes gladius et famis non erit in terra hac in gladio et fame consumentur prophetae illi
JER|14|16|et populi quibus prophetant erunt proiecti in viis Hierusalem prae fame et gladio et non erit qui sepeliat eos ipsi et uxores eorum filii et filiae eorum et effundam super eos malum suum
JER|14|17|et dices ad eos verbum istud deducant oculi mei lacrimam per noctem et diem et non taceant quoniam contritione magna contrita est virgo filia populi mei plaga pessima vehementer
JER|14|18|si egressus fuero ad agros ecce occisi gladio et si introiero in civitatem ecce adtenuati fame propheta quoque et sacerdos abierunt in terram quam ignorabant
JER|14|19|numquid proiciens abiecisti Iudam aut Sion abominata est anima tua quare ergo percussisti nos ita ut nulla sit sanitas expectavimus pacem et non est bonum et tempus curationis et ecce turbatio
JER|14|20|cognovimus Domine impietates nostras iniquitatem patrum nostrorum quia peccavimus tibi
JER|14|21|ne nos des in obprobrium propter nomen tuum neque facias nobis contumeliam solii gloriae tuae recordare ne irritum facias foedus tuum nobiscum
JER|14|22|numquid sunt in sculptilibus gentium qui pluant aut caeli possunt dare imbres nonne tu es Domine Deus noster quem expectavimus tu enim fecisti omnia haec
JER|15|1|et dixit Dominus ad me si steterit Moses et Samuhel coram me non est anima mea ad populum istum eice illos a facie mea et egrediantur
JER|15|2|quod si dixerint ad te quo egrediemur dices ad eos haec dicit Dominus qui ad mortem ad mortem et qui ad gladium ad gladium et qui ad famem ad famem et qui ad captivitatem ad captivitatem
JER|15|3|et visitabo super eos quattuor species dicit Dominus gladium ad occisionem et canes ad lacerandum et volatilia caeli et bestias terrae ad devorandum et dissipandum
JER|15|4|et dabo eos in fervorem universis regnis terrae propter Manassem filium Ezechiae regis Iuda super omnibus quae fecit in Hierusalem
JER|15|5|quis enim miserebitur tui Hierusalem aut quis contristabitur pro te aut quis ibit ad rogandum pro pace tua
JER|15|6|tu reliquisti me dicit Dominus retrorsum abisti et extendam manum meam super te et interficiam te laboravi rogans
JER|15|7|et dispergam eos ventilabro in portis terrae interfeci et perdidi populum meum et tamen a viis suis non sunt reversi
JER|15|8|multiplicatae sunt mihi viduae eius super harenam maris induxi eis super matrem adulescentis vastatorem meridie misi super civitates repente terrorem
JER|15|9|infirmata est quae peperit septem defecit anima eius occidit ei sol cum adhuc esset dies confusa est et erubuit et residuos eius in gladium dabo in conspectu inimicorum eorum ait Dominus
JER|15|10|vae mihi mater mea quare genuisti me virum rixae virum discordiae in universa terra non feneravi nec feneravit mihi quisquam omnes maledicunt mihi
JER|15|11|dicit Dominus si non reliquiae tuae in bonum si non occurri tibi in tempore adflictionis et in tempore tribulationis adversum inimicum
JER|15|12|numquid foederabitur ferrum ferro ab aquilone et aes
JER|15|13|divitias tuas et thesauros tuos in direptionem dabo gratis in omnibus peccatis tuis et in omnibus terminis tuis
JER|15|14|et adducam inimicos tuos de terra qua nescis quia ignis succensus est in furore meo super vos ardebit
JER|15|15|tu scis Domine recordare mei et visita me et tuere me ab his qui persequuntur me noli in patientia tua suscipere me scito quoniam sustinui pro te obprobrium
JER|15|16|inventi sunt sermones tui et comedi eos et factum est mihi verbum tuum in gaudium et in laetitiam cordis mei quoniam invocatum est nomen tuum super me Domine Deus exercituum
JER|15|17|non sedi in concilio ludentium et gloriatus sum a facie manus tuae solus sedebam quoniam comminatione replesti me
JER|15|18|quare factus est dolor meus perpetuus et plaga mea desperabilis rennuit curari facta est mihi quasi mendacium aquarum infidelium
JER|15|19|propter hoc haec dicit Dominus si converteris convertam te et ante faciem meam stabis et si separaveris pretiosum a vili quasi os meum eris convertentur ipsi ad te et tu non converteris ad eos
JER|15|20|et dabo te populo huic in murum aereum fortem et bellabunt adversum te et non praevalebunt quia ego tecum sum ut salvem te et eruam dicit Dominus
JER|15|21|et liberabo te de manu pessimorum et redimam te de manu fortium
JER|16|1|et factum est verbum Domini ad me dicens
JER|16|2|non accipies uxorem et non erunt tibi filii et filiae in loco isto
JER|16|3|quia haec dicit Dominus super filios et filias qui generantur in loco isto et super matres eorum quae genuerunt eos et super patres eorum de quorum stirpe sunt nati in terra hac
JER|16|4|mortibus aegrotationum morientur non plangentur et non sepelientur in sterquilinium super faciem terrae erunt et gladio et fame consumentur et erit cadaver eorum in escam volatilibus caeli et bestiis terrae
JER|16|5|haec enim dicit Dominus ne ingrediaris domum convivii neque vadas ad plangendum neque consoleris eos quia abstuli pacem meam a populo isto dicit Dominus misericordiam et miserationes
JER|16|6|et morientur grandes et parvi in terra ista non sepelientur neque plangentur et non se incident neque calvitium fiet pro eis
JER|16|7|et non frangent inter eos lugenti panem ad consolandum super mortuo et non dabunt eis potum calicis ad consolandum super patre suo et matre
JER|16|8|et domum convivii non ingredieris ut sedeas cum eis et comedas et bibas
JER|16|9|quia haec dicit Dominus exercituum Deus Israhel ecce ego auferam de loco isto in oculis vestris et in diebus vestris vocem gaudii et vocem laetitiae vocem sponsi et vocem sponsae
JER|16|10|et cum adnuntiaveris populo huic omnia verba haec et dixerint tibi quare locutus est Dominus super nos omne malum grande istud quae iniquitas nostra et quod peccatum nostrum quod peccavimus Domino Deo nostro
JER|16|11|dices ad eos quia dereliquerunt patres vestri me ait Dominus et abierunt post deos alienos et servierunt eis et adoraverunt eos et me dereliquerunt et legem meam non custodierunt
JER|16|12|sed et vos peius operati estis quam patres vestri ecce enim ambulat unusquisque post pravitatem cordis sui mali ut me non audiat
JER|16|13|et eiciam vos de terra hac in terram quam ignoratis vos et patres vestri et servietis ibi diis alienis die ac nocte qui non dabunt vobis requiem
JER|16|14|propterea ecce dies veniunt dicit Dominus et non dicetur ultra vivit Dominus qui eduxit filios Israhel de terra Aegypti
JER|16|15|sed vivit Dominus qui eduxit filios Israhel de terra aquilonis et de universis terris ad quas eieci eos et reducam eos in terram suam quam dedi patribus eorum
JER|16|16|ecce ego mittam piscatores multos dicit Dominus et piscabuntur eos et post haec mittam eis multos venatores et venabuntur eos de omni monte et de omni colle et de cavernis petrarum
JER|16|17|quia oculi mei super omnes vias eorum non sunt absconditae a facie mea et non fuit occulta iniquitas eorum ab oculis meis
JER|16|18|et reddam primum duplices iniquitates et peccata eorum quia contaminaverunt terram meam in morticinis idolorum suorum et abominationibus suis impleverunt hereditatem meam
JER|16|19|Domine fortitudo mea et robur meum et refugium meum in die tribulationis ad te gentes venient ab extremis terrae et dicent vere mendacium possederunt patres nostri vanitatem quae eis non profuit
JER|16|20|numquid faciet sibi homo deos et ipsi non sunt dii
JER|16|21|idcirco ecce ego ostendam eis per vicem hanc ostendam eis manum meam et virtutem meam et scient quia nomen mihi Dominus
JER|17|1|peccatum Iuda scriptum est stilo ferreo in ungue adamantino exaratum super latitudinem cordis eorum et in cornibus ararum eorum
JER|17|2|cum recordati fuerint filii eorum ararum suarum et lucorum lignorumque frondentium in montibus excelsis
JER|17|3|sacrificantes in agro fortitudinem tuam et omnes thesauros tuos in direptionem dabo excelsa tua propter peccata in universis finibus tuis
JER|17|4|et relinqueris sola ab hereditate tua quam dedi tibi et servire te faciam inimicis tuis in terra quam ignoras quoniam ignem succendisti in furore meo usque in aeternum ardebit
JER|17|5|haec dicit Dominus maledictus homo qui confidit in homine et ponit carnem brachium suum et a Domino recedit cor eius
JER|17|6|erit enim quasi myrice in deserto et non videbit cum venerit bonum sed habitabit in siccitate in deserto in terra salsuginis et inhabitabili
JER|17|7|benedictus vir qui confidit in Domino et erit Dominus fiducia eius
JER|17|8|et erit quasi lignum quod transplantatur super aquas quod ad humorem mittit radices suas et non timebit cum venerit aestus et erit folium eius viride et in tempore siccitatis non erit sollicitum nec aliquando desinet facere fructum
JER|17|9|pravum est cor omnium et inscrutabile quis cognoscet illud
JER|17|10|ego Dominus scrutans cor et probans renes qui do unicuique iuxta viam et iuxta fructum adinventionum suarum
JER|17|11|perdix fovit quae non peperit fecit divitias et non in iudicio in dimidio dierum suorum derelinquet eas et in novissimo suo erit insipiens
JER|17|12|solium gloriae altitudinis a principio locus sanctificationis nostrae
JER|17|13|expectatio Israhel Domine omnes qui te derelinquunt confundentur recedentes in terra scribentur quoniam dereliquerunt venam aquarum viventium Dominum
JER|17|14|sana me Domine et sanabor salvum me fac et salvus ero quoniam laus mea tu es
JER|17|15|ecce ipsi dicunt ad me ubi est verbum Domini veniat
JER|17|16|et ego non sum turbatus te pastorem sequens et diem hominis non desideravi tu scis quod egressum est de labiis meis rectum in conspectu tuo fuit
JER|17|17|non sis mihi tu formidini spes mea tu in die adflictionis
JER|17|18|confundantur qui persequuntur me et non confundar ego paveant illi et non paveam ego induc super eos diem adflictionis et duplici contritione contere eos
JER|17|19|haec dicit Dominus ad me vade et sta in porta filiorum populi per quam ingrediuntur reges Iuda et egrediuntur et in cunctis portis Hierusalem
JER|17|20|et dices ad eos audite verbum Domini reges Iuda et omnis Iudaea cunctique habitatores Hierusalem qui ingredimini per portas istas
JER|17|21|haec dicit Dominus custodite animas vestras et nolite portare pondera in die sabbati nec inferatis per portas Hierusalem
JER|17|22|et nolite eicere onera de domibus vestris in die sabbati et omne opus non facietis sanctificate diem sabbati sicut praecepi patribus vestris
JER|17|23|et non audierunt nec inclinaverunt aurem suam sed induraverunt cervicem suam ne audirent me et ne acciperent disciplinam
JER|17|24|et erit si audieritis me dicit Dominus ut non inferatis onera per portas civitatis huius in die sabbati et si sanctificaveritis diem sabbati ne faciatis in ea omne opus
JER|17|25|ingredientur per portas civitatis huius reges et principes sedentes super solium David et ascendentes in curribus et equis ipsi et principes eorum vir Iuda et habitatores Hierusalem et habitabitur civitas haec in sempiternum
JER|17|26|et venient de civitate Iuda et de circuitu Hierusalem et de terra Beniamin et de campestribus et de montuosis et ab austro portantes holocaustum et victimam et sacrificium et tus et inferent oblationem in domum Domini
JER|17|27|si autem non audieritis me ut sanctificetis diem sabbati et ne portetis onus et ne inferatis per portas Hierusalem in die sabbati succendam ignem in portis eius et devorabit domos Hierusalem et non extinguetur
JER|18|1|verbum quod factum est ad Hieremiam a Domino dicens
JER|18|2|surge et descende in domum figuli et ibi audies verba mea
JER|18|3|et descendi in domum figuli et ecce ipse faciebat opus super rotam
JER|18|4|et dissipatum est vas quod ipse faciebat e luto manibus suis conversusque fecit illud vas alterum sicut placuerat in oculis eius ut faceret
JER|18|5|et factum est verbum Domini ad me dicens
JER|18|6|numquid sicut figulus iste non potero facere vobis domus Israhel ait Dominus ecce sicut lutum in manu figuli sic vos in manu mea domus Israhel
JER|18|7|repente loquar adversum gentem et adversum regnum ut eradicem et destruam et disperdam illud
JER|18|8|si paenitentiam egerit gens illa a malo suo quod locutus sum adversum eam agam et ego paenitentiam super malo quod cogitavi ut facerem ei
JER|18|9|et subito loquar de gente et regno ut aedificem et ut plantem illud
JER|18|10|si fecerit malum in oculis meis ut non audiat vocem meam paenitentiam agam super bono quod locutus sum ut facerem ei
JER|18|11|nunc ergo dic viro Iudae et habitatoribus Hierusalem dicens haec dicit Dominus ecce ego fingo contra vos malum et cogito contra vos cogitationem revertatur unusquisque a via sua mala et dirigite vias vestras et studia vestra
JER|18|12|qui dixerunt desperavimus post cogitationes enim nostras ibimus et unusquisque pravitatem cordis sui mali faciemus
JER|18|13|ideo haec dicit Dominus interrogate gentes quis audivit talia horribilia quae fecit nimis virgo Israhel
JER|18|14|numquid deficiet de petra agri nix Libani aut evelli possunt aquae erumpentes frigidae et defluentes
JER|18|15|quia oblitus est mei populus meus frustra libantes et inpingentes in viis suis in semitis saeculi ut ambularent per eas in itinere non trito
JER|18|16|ut fieret terra eorum in desolationem et in sibilum sempiternum omnis qui praeterit per eam obstupescet et movebit caput suum
JER|18|17|sicut ventus urens dispergam eos coram inimico dorsum et non faciem ostendam eis in die perditionis eorum
JER|18|18|et dixerunt venite et cogitemus contra Hieremiam cogitationes non enim peribit lex a sacerdote neque consilium a sapiente nec sermo a propheta venite et percutiamus eum lingua et non adtendamus ad universos sermones eius
JER|18|19|adtende Domine ad me et audi vocem adversariorum meorum
JER|18|20|numquid redditur pro bono malum quia foderunt foveam animae meae recordare quod steterim in conspectu tuo ut loquerer pro eis bonum et averterem indignationem tuam ab eis
JER|18|21|propterea da filios eorum in famem et deduc eos in manus gladii fiant uxores eorum absque liberis et viduae et viri earum interficiantur morte iuvenes eorum confodiantur gladio in proelio
JER|18|22|audiatur clamor de domibus eorum adduces enim super eos latronem repente quia foderunt foveam ut caperent me et laqueos absconderunt pedibus meis
JER|18|23|tu autem Domine scis omne consilium eorum adversum me in mortem ne propitieris iniquitati eorum et peccatum eorum a facie tua non deleatur fiant corruentes in conspectu tuo in tempore furoris tui abutere eis
JER|19|1|haec dicit Dominus vade et accipe lagunculam figuli testeam a senioribus populi et a senioribus sacerdotum
JER|19|2|et egredere ad vallem filii Ennom quae est iuxta introitum portae Fictilis et praedicabis ibi verba quae ego loquar ad te
JER|19|3|et dices audite verbum Domini reges Iuda et habitatores Hierusalem haec dicit Dominus exercituum Deus Israhel ecce ego inducam adflictionem super locum istum ita ut omnis qui audierit illam tinniant aures eius
JER|19|4|eo quod dereliquerint me et alienum fecerint locum istum et libaverint in eo diis alienis quos nescierunt ipsi et patres eorum et reges Iuda et repleverunt locum istum sanguine innocentium
JER|19|5|et aedificaverunt excelsa Baali ad conburendos filios suos igni in holocaustum Baali quae non praecepi nec locutus sum nec ascenderunt in cor meum
JER|19|6|propterea ecce dies veniunt dicit Dominus et non vocabitur locus iste amplius Thofeth et vallis filii Ennom sed vallis Occisionis
JER|19|7|et dissipabo consilium Iudae et Hierusalem in loco isto et subvertam eos gladio in conspectu inimicorum suorum et in manu quaerentium animas eorum et dabo cadavera eorum escam volatilibus caeli et bestiis terrae
JER|19|8|et ponam civitatem hanc in stuporem et in sibilum omnis qui praeterierit per eam obstupescet et sibilabit super universa plaga eius
JER|19|9|et cibabo eos carnibus filiorum suorum et carnibus filiarum suarum et unusquisque carnes amici sui comedet in obsidione et in angustia in qua concludent eos inimici eorum et qui quaerunt animas eorum
JER|19|10|et conteres lagunculam in oculis virorum qui ibunt tecum
JER|19|11|et dices ad eos haec dicit Dominus exercituum sic conteram populum istum et civitatem istam sicut conteritur vas figuli quod non potest ultra instaurari et in Thofeth sepelientur eo quod non sit alius locus ad sepeliendum
JER|19|12|sic faciam loco huic ait Dominus et habitatoribus eius ut ponam civitatem istam sicut Thofeth
JER|19|13|et erunt domus Hierusalem et domus regum Iuda sicut locus Thofeth inmundae omnes domus in quarum domatibus sacrificaverunt omni militiae caeli et libaverunt libamina diis alienis
JER|19|14|venit autem Hieremias de Thofeth quo miserat eum Dominus ad prophetandum et stetit in atrio domus Domini et dixit ad omnem populum
JER|19|15|haec dicit Dominus exercituum Deus Israhel ecce ego inducam super civitatem hanc et super omnes urbes eius universa mala quae locutus sum adversum eam quoniam induraverunt cervicem suam ut non audirent sermones meos
JER|20|1|et audivit Phassur filius Emmer sacerdos qui constitutus erat princeps in domo Domini Hieremiam prophetantem sermones istos
JER|20|2|et percussit Phassur Hieremiam prophetam et misit eum in nervum quod erat in porta Beniamin superiori in domo Domini
JER|20|3|cumque inluxisset in crastinum eduxit Phassur Hieremiam de nervo et dixit ad eum Hieremias non Phassur vocavit Dominus nomen tuum sed Pavorem undique
JER|20|4|quia haec dicit Dominus ecce ego dabo te in pavorem te et omnes amicos tuos et corruent gladio inimicorum suorum et oculi tui videbunt et omnem Iudam dabo in manu regis Babylonis et traducet eos in Babylonem et percutiet eos gladio
JER|20|5|et dabo universam substantiam civitatis huius et omnem laborem eius omneque pretium et cunctos thesauros regum Iuda dabo in manu inimicorum eorum et diripient eos et tollent et ducent in Babylonem
JER|20|6|tu autem Phassur et omnes habitatores domus tuae ibitis in captivitatem et in Babylonem venies et ibi morieris ibique sepelieris tu et omnes amici tui quibus prophetasti mendacium
JER|20|7|seduxisti me Domine et seductus sum fortior me fuisti et invaluisti factus sum in derisum tota die omnes subsannant me
JER|20|8|quia iam olim loquor vociferans iniquitatem et vastitatem clamito et factus est mihi sermo Domini in obprobrium et in derisum tota die
JER|20|9|et dixi non recordabor eius neque loquar ultra in nomine illius et factus est in corde meo quasi ignis exaestuans claususque in ossibus meis et defeci ferre non sustinens
JER|20|10|audivi enim contumelias multorum et terrorem in circuitu persequimini et persequamur eum ab omnibus viris qui erant pacifici mei et custodientes latus meum si quo modo decipiatur et praevaleamus adversus eum et consequamur ultionem ex eo
JER|20|11|Dominus autem mecum est quasi bellator fortis idcirco qui persequuntur me cadent et infirmi erunt confundentur vehementer quia non intellexerunt obprobrium sempiternum quod numquam delebitur
JER|20|12|et tu Domine exercituum probator iusti qui vides renes et cor videam quaeso ultionem tuam ex eis tibi enim revelavi causam meam
JER|20|13|cantate Domino laudate Dominum quia liberavit animam pauperis de manu malorum
JER|20|14|maledicta dies in qua natus sum dies in qua peperit me mater mea non sit benedicta
JER|20|15|maledictus vir qui adnuntiavit patri meo dicens natus est tibi puer masculus et quasi gaudio laetificavit eum
JER|20|16|sit homo ille ut sunt civitates quas subvertit Dominus et non paenituit eum audiat clamorem mane et ululatum in tempore meridiano
JER|20|17|qui non me interfecit a vulva ut fieret mihi mater mea sepulchrum et vulva eius conceptus aeternus
JER|20|18|quare de vulva egressus sum ut viderem laborem et dolorem et consumerentur in confusione dies mei
JER|21|1|verbum quod factum est ad Hieremiam a Domino quando misit ad eum rex Sedecias Phassur filium Melchiae et Sophoniam filium Maasiae sacerdotem dicens
JER|21|2|interroga pro nobis Dominum quia Nabuchodonosor rex Babylonis proeliatur adversum nos si forte faciat Dominus nobiscum secundum omnia mirabilia sua et recedat a nobis
JER|21|3|et dixit Hieremias ad eos sic dicetis Sedeciae
JER|21|4|haec dicit Dominus Deus Israhel ecce ego convertam vasa belli quae in manibus vestris sunt et quibus vos pugnatis adversum regem Babylonis et Chaldeos qui obsident vos in circuitu murorum et congregabo ea in medio civitatis huius
JER|21|5|et debellabo ego vos in manu extenta et brachio forti et in furore et in indignatione et in ira grandi
JER|21|6|et percutiam habitatores civitatis huius homines et bestiae pestilentia magna morientur
JER|21|7|et post haec ait Dominus dabo Sedeciam regem Iuda et servos eius et populum eius et qui derelicti sunt in civitate hac a peste et gladio et fame in manu Nabuchodonosor regis Babylonis et in manu inimicorum eorum et in manu quaerentium animam eorum et percutiet eos in ore gladii et non movebitur neque parcet nec miserebitur
JER|21|8|et ad populum hunc dices haec dicit Dominus ecce ego do coram vobis viam vitae et viam mortis
JER|21|9|qui habitaverit in urbe hac morietur gladio et fame et peste qui autem egressus fuerit et transfugerit ad Chaldeos qui obsident vos vivet et erit ei anima sua quasi spolium
JER|21|10|posui enim faciem meam super civitatem hanc in malum et non in bonum ait Dominus in manu regis Babylonis dabitur et exuret eam igni
JER|21|11|et domui regis Iuda audite verbum Domini
JER|21|12|domus David haec dicit Dominus iudicate mane iudicium et eruite vi oppressum de manu calumniantis ne forte egrediatur ut ignis indignatio mea et succendatur et non sit qui extinguat propter malitiam studiorum vestrorum
JER|21|13|ecce ego ad te habitatricem vallis solidae atque campestris ait Dominus qui dicitis quis percutiet nos et quis ingredietur domos nostras
JER|21|14|et visitabo super vos iuxta fructum studiorum vestrorum dicit Dominus et succendam ignem in saltu eius et devorabit omnia in circuitu eius
JER|22|1|haec dicit Dominus descende in domum regis Iuda et loqueris ibi verbum hoc
JER|22|2|et dices audi verbum Domini rex Iuda qui sedes super solium David tu et servi tui et populus tuus qui ingredimini per portas istas
JER|22|3|haec dicit Dominus facite iudicium et iustitiam et liberate vi oppressum de manu calumniatoris et advenam et pupillum et viduam nolite contristare neque opprimatis inique et sanguinem innocentem ne effundatis in loco isto
JER|22|4|si enim facientes feceritis verbum istud ingredientur per portas domus huius reges sedentes de genere David super thronum eius et ascendentes currus et equos ipsi et servi et populus eorum
JER|22|5|quod si non audieritis verba haec in memet ipso iuravi dicit Dominus quia in solitudinem erit domus haec
JER|22|6|quia haec dicit Dominus super domum regis Iuda Galaad tu mihi caput Libani si non posuero te solitudinem urbes inhabitabiles
JER|22|7|et sanctificabo super te interficientem virum et arma eius et succident electam cedrum tuam et praecipitabunt in ignem
JER|22|8|et pertransibunt gentes multae per civitatem hanc et dicet unusquisque proximo suo quare fecit Dominus sic civitati huic grandi
JER|22|9|et respondebunt eo quod dereliquerint pactum Domini Dei sui et adoraverint deos alienos et servierint eis
JER|22|10|nolite flere mortuum neque lugeatis super eum fletu plangite eum qui egreditur quia non revertetur ultra nec videbit terram nativitatis suae
JER|22|11|quia haec dicit Dominus ad Sellum filium Iosiae regem Iuda qui regnavit pro Iosia patre suo qui egressus est de loco isto non revertetur huc amplius
JER|22|12|sed in loco ad quem transtuli eum ibi morietur et terram istam non videbit amplius
JER|22|13|vae qui aedificat domum suam in iniustitia et cenacula sua non in iudicio amicum suum opprimet frustra et mercedem eius non reddet ei
JER|22|14|qui dicit aedificabo mihi domum latam et cenacula spatiosa qui aperit sibi fenestras et facit laquearia cedrina pingitque sinopide
JER|22|15|numquid regnabis quoniam confers te cedro pater tuus numquid non comedit et bibit et fecit iudicium et iustitiam tunc cum bene erat ei
JER|22|16|iudicavit causam pauperis et egeni in bonum suum numquid non ideo quia cognovit me dicit Dominus
JER|22|17|tui vero oculi et cor ad avaritiam et ad sanguinem innocentem fundendum et ad calumniam et ad cursum mali operis
JER|22|18|propterea haec dicit Dominus ad Ioachim filium Iosiae regem Iuda non plangent eum vae frater et vae fratres non concrepabunt ei vae domine et vae inclite
JER|22|19|sepultura asini sepelietur putrefactus et proiectus extra portas Hierusalem
JER|22|20|ascende Libanum et clama et in Basan da vocem tuam et clama ad transeuntes quia contriti sunt omnes amatores tui
JER|22|21|locutus sum ad te in abundantia tua dixisti non audiam haec est via tua ab adulescentia tua quia non audisti vocem meam
JER|22|22|omnes pastores tuos pascet ventus et amatores tui in captivitatem ibunt et tunc confunderis et erubesces ab omni malitia tua
JER|22|23|quae sedes in Libano et nidificas in cedris quomodo congemuisti cum venissent tibi dolores quasi dolores parturientis
JER|22|24|vivo ego dicit Dominus quia si fuerit Iechonias filius Ioachim regis Iuda anulus in manu dextera mea inde avellam eum
JER|22|25|et dabo te in manu quaerentium animam tuam et in manu quorum tu formidas faciem et in manu Nabuchodonosor regis Babylonis et in manu Chaldeorum
JER|22|26|et mittam te et matrem tuam quae genuit te in terram alienam in qua nati non estis ibique moriemini
JER|22|27|et in terram ad quam ipsi levant animam suam ut revertantur illuc non revertentur
JER|22|28|numquid vas fictile atque contritum vir iste Iechonias numquid vas absque omni voluptate quare abiecti sunt ipse et semen eius et proiecti in terram quam ignoraverunt
JER|22|29|terra terra terra audi sermonem Domini
JER|22|30|haec dicit Dominus scribe virum istum sterilem virum qui in diebus suis non prosperabitur nec enim erit de semine eius vir qui sedeat super solium David et potestatem habeat ultra in Iuda
JER|23|1|vae pastoribus qui disperdunt et dilacerant gregem pascuae meae dicit Dominus
JER|23|2|ideo haec dicit Dominus Deus Israhel ad pastores qui pascunt populum meum vos dispersistis gregem meum eiecistis eos et non visitastis eos ecce ego visitabo super vos malitiam studiorum vestrorum ait Dominus
JER|23|3|et ego congregabo reliquias gregis mei de omnibus terris ad quas eiecero eos illuc et convertam eos ad rura sua et crescent et multiplicabuntur
JER|23|4|et suscitabo super eos pastores et pascent eos non formidabunt ultra et non pavebunt et nullus quaeretur ex numero dicit Dominus
JER|23|5|ecce dies veniunt ait Dominus et suscitabo David germen iustum et regnabit rex et sapiens erit et faciet iudicium et iustitiam in terra
JER|23|6|in diebus illius salvabitur Iuda et Israhel habitabit confidenter et hoc est nomen quod vocabunt eum Dominus iustus noster
JER|23|7|propter hoc ecce dies veniunt dicit Dominus et non dicent ultra vivit Dominus qui eduxit filios Israhel de terra Aegypti
JER|23|8|sed vivit Dominus qui eduxit et adduxit semen domus Israhel de terra aquilonis et de cunctis terris ad quas eieceram eos illuc et habitabunt in terra sua
JER|23|9|ad prophetas contritum est cor meum in medio mei contremuerunt omnia ossa mea factus sum quasi vir ebrius et quasi homo madidus a vino a facie Domini et a facie verborum sanctorum eius
JER|23|10|quia adulteris repleta est terra quia a facie maledictionis luxit terra arefacta sunt arva deserti factus est cursus eorum malus et fortitudo eorum dissimilis
JER|23|11|propheta namque et sacerdos polluti sunt et in domo mea inveni malum eorum ait Dominus
JER|23|12|idcirco via eorum erit quasi lubricum in tenebris inpellentur enim et corruent in ea adferam enim super eos mala annum visitationis eorum ait Dominus
JER|23|13|et in prophetis Samariae vidi fatuitatem prophetabant in Baal et decipiebant populum meum Israhel
JER|23|14|et in prophetis Hierusalem vidi similitudinem adulterium et iter mendacii et confortaverunt manus pessimorum ut non converteretur unusquisque a malitia sua facti sunt mihi omnes Sodoma et habitatores eius quasi Gomorra
JER|23|15|propterea haec dicit Dominus exercituum ad prophetas ecce ego cibabo eos absinthio et potabo eos felle a prophetis enim Hierusalem est egressa pollutio super omnem terram
JER|23|16|haec dicit Dominus exercituum nolite audire verba prophetarum qui prophetant vobis et decipiunt vos visionem cordis sui loquuntur non de ore Domini
JER|23|17|dicunt his qui blasphemant me locutus est Dominus pax erit vobis et omni qui ambulat in pravitate cordis sui dixerunt non veniet super vos malum
JER|23|18|quis enim adfuit in consilio Domini et vidit et audivit sermonem eius quis consideravit verbum illius et audivit
JER|23|19|ecce turbo dominicae indignationis egredietur et tempestas erumpens super caput impiorum veniet
JER|23|20|non revertetur furor Domini usque dum faciat et usque dum conpleat cogitationem cordis sui in novissimis diebus intellegetis consilium eius
JER|23|21|non mittebam prophetas et ipsi currebant non loquebar ad eos et ipsi prophetabant
JER|23|22|si stetissent in consilio meo et nota fecissent verba mea populo meo avertissem utique eos a via sua mala et a pessimis cogitationibus suis
JER|23|23|putasne Deus e vicino ego sum dicit Dominus et non Deus de longe
JER|23|24|si occultabitur vir in absconditis et ego non videbo eum dicit Dominus numquid non caelum et terram ego impleo ait Dominus
JER|23|25|audivi quae dixerunt prophetae prophetantes in nomine meo mendacium atque dicentes somniavi somniavi
JER|23|26|usquequo istud in corde est prophetarum vaticinantium mendacium et prophetantium seductiones cordis sui
JER|23|27|qui volunt facere ut obliviscatur populus meus nominis mei propter somnia eorum quae narrant unusquisque ad proximum suum sicut obliti sunt patres eorum nominis mei propter Baal
JER|23|28|propheta qui habet somnium narret somnium et qui habet sermonem meum loquatur sermonem meum vere quid paleis ad triticum dicit Dominus
JER|23|29|numquid non verba mea sunt quasi ignis ait Dominus et quasi malleus conterens petram
JER|23|30|propterea ecce ego ad prophetas ait Dominus qui furantur verba mea unusquisque a proximo suo
JER|23|31|ecce ego ad prophetas ait Dominus qui adsumunt linguas suas et aiunt dicit Dominus
JER|23|32|ecce ego ad prophetas somniantes mendacium ait Dominus qui narraverunt ea et seduxerunt populum meum in mendacio suo et in miraculis suis cum ego non misissem eos nec mandassem eis qui nihil profuerunt populo huic dicit Dominus
JER|23|33|si igitur interrogaverit te populus iste vel propheta aut sacerdos dicens quod est onus Domini dices ad eos ut quid vobis onus proiciam quippe vos dicit Dominus
JER|23|34|et prophetes et sacerdos et populus qui dicit onus Domini visitabo super virum illum et super domum eius
JER|23|35|haec dicetis unusquisque ad proximum et ad fratrem suum quid respondit Dominus et quid locutus est Dominus
JER|23|36|et onus Domini ultra non memorabitur quia onus erit unicuique sermo suus et pervertitis verba Dei viventis Domini exercituum Dei nostri
JER|23|37|haec dices ad prophetam quid respondit tibi Dominus et quid locutus est Dominus
JER|23|38|si autem onus Domini dixeritis propter hoc haec dicit Dominus quia dixistis sermonem istum onus Domini et misi ad vos dicens nolite dicere onus Domini
JER|23|39|propterea ecce ego tollam vos portans et derelinquam vos et civitatem quam dedi vobis et patribus vestris a facie mea
JER|23|40|et dabo vos in obprobrium sempiternum et in ignominiam aeternam quae numquam oblivione delebitur
JER|24|1|ostendit mihi Dominus et ecce duo calathi pleni ficis positi ante templum Domini postquam transtulit Nabuchodonosor rex Babylonis Iechoniam filium Ioachim regem Iuda et principes eius et fabrum et inclusorem de Hierusalem et adduxit eos in Babylonem
JER|24|2|calathus unus ficus bonas habebat nimis ut solent ficus esse primi temporis et calathus unus ficus habebat malas nimis quae comedi non poterant eo quod essent malae
JER|24|3|et dixit Dominus ad me quid tu vides Hieremia et dixi ficus ficus bonas bonas valde et malas malas valde quae comedi non possunt eo quod sint malae
JER|24|4|et factum est verbum Domini ad me dicens
JER|24|5|haec dicit Dominus Deus Israhel sicut ficus hae bonae sic cognoscam transmigrationem Iuda quam emisi de loco isto in terram Chaldeorum in bonum
JER|24|6|et ponam oculos meos super eos ad placandum et reducam eos in terram hanc et aedificabo eos et non destruam et plantabo eos et non evellam
JER|24|7|et dabo eis cor ut sciant me quia ego sum Dominus et erunt mihi in populum et ego ero eis in Deum quia revertentur ad me in toto corde suo
JER|24|8|et sicut ficus pessimae quae comedi non possunt eo quod sint malae haec dicit Dominus sic dabo Sedeciam regem Iuda et principes eius et reliquos de Hierusalem qui remanserunt in urbe hac et qui habitant in terra Aegypti
JER|24|9|et dabo eos in vexationem adflictionemque omnibus regnis terrae in obprobrium et in parabolam et in proverbium et in maledictionem in universis locis ad quos eieci eos
JER|24|10|et mittam in eis gladium et famem et pestem donec consumantur de terra quam dedi eis et patribus eorum
JER|25|1|verbum quod factum est ad Hieremiam de omni populo Iudae in anno quarto Ioachim filii Iosiae regis Iuda ipse est annus primus Nabuchodonosor regis Babylonis
JER|25|2|quae locutus est Hieremias propheta ad omnem populum Iuda et ad universos habitatores Hierusalem dicens
JER|25|3|a tertiodecimo anno Iosiae filii Amon regis Iuda usque ad diem hanc iste est tertius et vicesimus annus factum est verbum Domini ad me et locutus sum ad vos de nocte consurgens et loquens et non audistis
JER|25|4|et misit Dominus ad vos omnes servos suos prophetas consurgens diluculo mittensque et non audistis neque inclinastis aures vestras ut audiretis
JER|25|5|cum diceret revertimini unusquisque a via sua mala et a pessimis cogitationibus vestris et habitabitis in terram quam dedit Dominus vobis et patribus vestris a saeculo et usque in saeculum
JER|25|6|et nolite ire post deos alienos ut serviatis eis adoretisque eos neque me ad iracundiam provocetis in operibus manuum vestrarum et non adfligam vos
JER|25|7|et non audistis me dicit Dominus ut me ad iracundiam provocaretis in operibus manuum vestrarum in malum vestrum
JER|25|8|propterea haec dicit Dominus exercituum pro eo quod non audistis verba mea
JER|25|9|ecce ego mittam et adsumam universas cognationes aquilonis ait Dominus et ad Nabuchodonosor regem Babylonis servum meum et adducam eos super terram istam et super habitatores eius et super omnes nationes quae in circuitu illius sunt et interficiam eos et ponam eos in stuporem et in sibilum et in solitudines sempiternas
JER|25|10|perdamque ex eis vocem gaudii et vocem laetitiae vocem sponsae et vocem sponsi vocem molae et lumen lucernae
JER|25|11|et erit universa terra eius in solitudinem et in stuporem et servient omnes gentes istae regi Babylonis septuaginta annis
JER|25|12|cumque impleti fuerint anni septuaginta visitabo super regem Babylonis et super gentem illam dicit Dominus iniquitatem eorum et super terram Chaldeorum et ponam illam in solitudines sempiternas
JER|25|13|et adducam super terram illam omnia verba mea quae locutus sum contra eam omne quod scriptum est in libro isto quaecumque prophetavit Hieremias adversum omnes gentes
JER|25|14|quia servierunt eis cum essent gentes multae et reges magni et reddam eis secundum opera eorum et secundum facta manuum suarum
JER|25|15|quia sic dicit Dominus exercituum Deus Israhel sume calicem vini furoris huius de manu mea et propinabis de illo cunctis gentibus ad quas ego mittam te
JER|25|16|et bibent et turbabuntur et insanient a facie gladii quem ego mittam inter eos
JER|25|17|et accepi calicem de manu Domini et propinavi cunctis gentibus ad quas misit me Dominus
JER|25|18|Hierusalem et civitatibus Iudae et regibus eius et principibus eius ut darem eos in solitudinem et in stuporem in sibilum et in maledictionem sicut est dies ista
JER|25|19|Pharaoni regi Aegypti et servis eius et principibus eius et omni populo eius
JER|25|20|et universis generaliter cunctis regibus terrae Ausitidis et cunctis regibus terrae Philisthim et Ascaloni et Gazae et Accaroni et reliquiis Azoti
JER|25|21|Idumeae et Moab et filiis Ammon
JER|25|22|et cunctis regibus Tyri et cunctis regibus Sidonis et regibus terrae insularum qui sunt trans mare
JER|25|23|et Dedan et Theman et Buz et universis qui adtonsi sunt in comam
JER|25|24|et cunctis regibus Arabiae et cunctis regibus occidentis qui habitant in deserto
JER|25|25|et cunctis regibus Zambri et cunctis regibus Aelam et cunctis regibus Medorum
JER|25|26|et cunctis regibus aquilonis de prope et de longe unicuique contra fratrem suum et omnibus regnis terrae quae super faciem eius sunt et rex Sesach bibet post eos
JER|25|27|et dices ad eos haec dicit Dominus exercituum Deus Israhel bibite et inebriamini et vomite et cadite neque surgatis a facie gladii quem ego mittam inter vos
JER|25|28|cumque noluerint accipere calicem de manu ut bibant dices ad eos haec dicit Dominus exercituum bibentes bibetis
JER|25|29|quia ecce in civitate in qua invocatum est nomen meum ego incipio adfligere et vos quasi innocentes inmunes eritis non eritis inmunes gladium enim ego voco super omnes habitatores terrae dicit Dominus exercituum
JER|25|30|et tu prophetabis ad eos omnia verba haec et dices ad illos Dominus de excelso rugiet et de habitaculo sancto suo dabit vocem suam rugiens rugiet super decorem suum celeuma quasi calcantium concinetur adversus omnes habitatores terrae
JER|25|31|pervenit sonitus usque ad extrema terrae quia iudicium Domino cum gentibus iudicatur ipse cum omni carne impios tradidit gladio dicit Dominus
JER|25|32|haec dicit Dominus exercituum ecce adflictio egredietur de gente in gentem et turbo magnus egredietur a summitatibus terrae
JER|25|33|et erunt interfecti Domini in die illa a summo terrae usque ad summum eius non plangentur et non colligentur neque sepelientur in sterquilinium super faciem terrae iacebunt
JER|25|34|ululate pastores et clamate et aspergite vos cinere optimates gregis quia conpleti sunt dies vestri ut interficiamini et dissipationes vestrae et cadetis quasi vasa pretiosa
JER|25|35|et peribit fuga a pastoribus et salvatio ab optimatibus gregis
JER|25|36|vox clamoris pastorum et ululatus optimatium gregis quia vastavit Dominus pascuam eorum
JER|25|37|et conticuerunt arva pacis a facie irae furoris Domini
JER|25|38|dereliquit quasi leo umbraculum suum facta est terra eorum in desolationem a facie irae columbae et a facie irae furoris Domini
JER|26|1|in principio regis Ioachim filii Iosiae regis Iuda factum est verbum istud a Domino dicens
JER|26|2|haec dicit Dominus sta in atrio domus Domini et loqueris ad omnes civitates Iuda de quibus veniunt ut adorent in domo Domini universos sermones quos ego mandavi tibi ut loquaris ad eos noli subtrahere verbum
JER|26|3|si forte audiant et convertantur unusquisque a via sua mala et paeniteat me mali quod cogito facere eis propter malitias studiorum eorum
JER|26|4|et dices ad eos haec dicit Dominus si non audieritis me ut ambuletis in lege mea quam dedi vobis
JER|26|5|ut audiatis sermones servorum meorum prophetarum quos ego misi ad vos de nocte consurgens et dirigens et non audistis
JER|26|6|dabo domum istam sicut Silo et urbem hanc dabo in maledictionem cunctis gentibus terrae
JER|26|7|et audierunt sacerdotes et prophetae et omnis populus Hieremiam loquentem verba haec in domo Domini
JER|26|8|cumque conplesset Hieremias loquens omnia quae praeceperat ei Dominus ut loqueretur ad universum populum adprehenderunt eum sacerdotes et prophetae et omnis populus dicens morte morietur
JER|26|9|quare prophetavit in nomine Domini dicens sicut Silo erit domus haec et urbs ista desolabitur eo quod non sit habitator et congregatus est omnis populus adversum Hieremiam in domum Domini
JER|26|10|et audierunt principes Iuda verba haec et ascenderunt de domo regis in domum Domini et sederunt in introitu portae Domini novae
JER|26|11|et locuti sunt sacerdotes et prophetae ad principes et ad omnem populum dicentes iudicium mortis est viro huic quia prophetavit adversum civitatem istam sicut audistis auribus vestris
JER|26|12|et ait Hieremias ad omnes principes et ad universum populum dicens Dominus misit me ut prophetarem ad domum istam et ad civitatem hanc omnia verba quae audistis
JER|26|13|nunc ergo bonas facite vias vestras et studia vestra et audite vocem Domini Dei vestri et paenitebit Dominum mali quod locutus est adversum vos
JER|26|14|ego autem ecce in manibus vestris sum facite mihi ut bonum et rectum est in oculis vestris
JER|26|15|verumtamen scitote et cognoscite quod si occideritis me sanguinem innocentem traditis contra vosmet ipsos et contra civitatem istam et habitatores eius in veritate enim misit me Dominus ad vos ut loquerer in auribus vestris omnia verba haec
JER|26|16|et dixerunt principes et omnis populus ad sacerdotes et prophetas non est viro huic iudicium mortis quia in nomine Domini Dei nostri locutus est ad nos
JER|26|17|surrexerunt ergo viri de senioribus terrae et dixerunt ad omnem coetum populi loquentes
JER|26|18|Michas de Morasthim fuit propheta in diebus Ezechiae regis Iudae et ait ad omnem populum Iudae dicens haec dicit Dominus exercituum Sion quasi ager arabitur et Hierusalem in acervum lapidum erit et mons domus in excelsa silvarum
JER|26|19|numquid morte condemnavit eum Ezechias rex Iuda et omnis Iuda numquid non timuerunt Dominum et deprecati sunt faciem Domini et paenituit Dominum mali quod locutus erat adversum eos itaque nos facimus malum grande contra animas nostras
JER|26|20|fuit quoque vir prophetans in nomine Domini Urias filius Semei de Cariathiarim et prophetavit adversum civitatem istam et adversum terram hanc iuxta universa verba Hieremiae
JER|26|21|et audivit rex Ioachim et omnes potentes et principes eius verba haec et quaesivit rex interficere eum et audivit Urias et timuit fugitque et ingressus est Aegyptum
JER|26|22|et misit rex Ioachim viros in Aegyptum Elnathan filium Achobor et viros cum eo in Aegyptum
JER|26|23|et eduxerunt Uriam de Aegypto et adduxerunt eum ad regem Ioachim et percussit eum gladio et proiecit cadaver eius in sepulchris vulgi ignobilis
JER|26|24|igitur manus Ahicam filii Saphan fuit cum Hieremia ut non traderetur in manu populi et interficerent eum
JER|27|1|in principio regni Ioachim filii Iosiae regis Iuda factum est verbum istud ad Hieremiam a Domino dicens
JER|27|2|haec dicit Dominus ad me fac tibi vincula et catenas et pones eas in collo tuo
JER|27|3|et mittes eas ad regem Edom et ad regem Moab et ad regem filiorum Ammon et ad regem Tyri et ad regem Sidonis in manu nuntiorum qui venerunt Hierusalem ad Sedeciam regem Iuda
JER|27|4|et praecipies eis ut ad dominos suos loquantur haec dicit Dominus exercituum Deus Israhel haec dicetis ad dominos vestros
JER|27|5|ego feci terram et hominem et iumenta quae sunt super faciem terrae in fortitudine mea magna et in brachio meo extento et dedi eam ei qui placuit in oculis meis
JER|27|6|et nunc itaque ego dedi omnes terras istas in manu Nabuchodonosor regis Babylonis servi mei insuper et bestias agri dedi ei ut serviant illi
JER|27|7|et servient ei omnes gentes et filio eius et filio filii eius donec veniat tempus terrae eius et ipsius et servient ei gentes multae et reges magni
JER|27|8|gens autem et regnum quod non servierit Nabuchodonosor regi Babylonis et quicumque non curvaverit collum suum sub iugo regis Babylonis in gladio et in fame et in peste visitabo super gentem illam ait Dominus donec consumam eos in manu eius
JER|27|9|vos ergo nolite audire prophetas vestros et divinos et somniatores et augures et maleficos qui dicunt vobis non servietis regi Babylonis
JER|27|10|quia mendacium prophetant vobis ut longe faciant vos de terra vestra et eiciant vos et pereatis
JER|27|11|porro gens quae subiecerit cervicem suam sub iugo regis Babylonis et servierit ei dimittam eam in terra sua dicit Dominus et colet eam et habitabit in ea
JER|27|12|et ad Sedeciam regem Iuda locutus sum secundum omnia verba haec dicens subicite colla vestra sub iugo regis Babylonis et servite ei et populo eius et vivetis
JER|27|13|quare moriemini tu et populus tuus gladio fame et peste sicut locutus est Dominus ad gentem quae servire noluerit regi Babylonis
JER|27|14|nolite audire verba prophetarum dicentium vobis non servietis regi Babylonis quia mendacium ipsi loquuntur vobis
JER|27|15|quia non misi eos ait Dominus et ipsi prophetant in nomine meo mendaciter ut eiciant vos et pereatis tam vos quam prophetae qui vaticinantur vobis
JER|27|16|et ad sacerdotes et ad populum istum locutus sum dicens haec dicit Dominus nolite audire verba prophetarum vestrorum qui prophetant vobis dicentes ecce vasa Domini revertentur de Babylone nunc cito mendacium enim prophetant vobis
JER|27|17|nolite ergo audire eos sed servite regi Babylonis ut vivatis quare datur haec civitas in solitudinem
JER|27|18|et si prophetae sunt et est verbum Domini in eis occurrant Domino exercituum ut non veniant vasa quae derelicta fuerant in domum Domini et in domum regis Iuda et in Hierusalem in Babylonem
JER|27|19|quia haec dicit Dominus exercituum ad columnas et ad mare et ad bases et ad reliqua vasorum quae remanserunt in civitate hac
JER|27|20|quae non tulit Nabuchodonosor rex Babylonis cum transferret Iechoniam filium Ioachim regem Iuda de Hierusalem in Babylonem et omnes optimates Iuda et Hierusalem
JER|27|21|quia haec dicit Dominus exercituum Deus Israhel ad vasa quae derelicta sunt in domum Domini et in domum regis Iuda et Hierusalem
JER|27|22|in Babylonem transferentur et ibi erunt usque ad diem visitationis suae dicit Dominus et adferri faciam ea et restitui in loco isto
JER|28|1|et factum est in anno illo in principio regni Sedeciae regis Iuda in anno quarto in mense quinto dixit ad me Ananias filius Azur propheta de Gabaon in domo Domini coram sacerdotibus et omni populo dicens
JER|28|2|haec dicit Dominus exercituum Deus Israhel contrivi iugum regis Babylonis
JER|28|3|adhuc duo anni dierum et ego referri faciam ad locum istum omnia vasa Domini quae tulit Nabuchodonosor rex Babylonis de loco isto et transtulit ea in Babylonem
JER|28|4|et Iechoniam filium Ioachim regem Iuda et omnem transmigrationem Iudae qui ingressi sunt in Babylonem ego convertam ad locum istum ait Dominus conteram enim iugum regis Babylonis
JER|28|5|et dixit Hieremias propheta ad Ananiam prophetam in oculis sacerdotum et in oculis omnis populi qui stabant in domo Domini
JER|28|6|et ait Hieremias propheta amen sic faciat Dominus suscitet Dominus verba tua quae prophetasti ut referantur vasa in domum Domini et omnis transmigratio de Babylone ad locum istum
JER|28|7|verumtamen audi verbum hoc quod ego loquor in auribus tuis et in auribus universi populi
JER|28|8|prophetae qui fuerunt ante me et te ab initio et prophetaverunt super terras multas et super regna magna de proelio et de adflictione et de fame
JER|28|9|propheta qui vaticinatus est pacem cum venerit verbum eius scietur propheta quem misit Dominus in veritate
JER|28|10|et tulit Ananias propheta catenam de collo Hieremiae prophetae et confregit eam
JER|28|11|et ait Ananias in conspectu omnis populi dicens haec dicit Dominus sic confringam iugum Nabuchodonosor regis Babylonis post duos annos dierum de collo omnium gentium
JER|28|12|et abiit Hieremias prophetes in viam suam et factum est verbum Domini ad Hieremiam postquam confregit Ananias propheta catenam de collo Hieremiae prophetae dicens
JER|28|13|vade et dices Ananiae haec dicit Dominus catenas ligneas contrivisti et facies pro eis catenas ferreas
JER|28|14|quia haec dicit Dominus exercituum Deus Israhel iugum ferreum posui super collum cunctarum gentium istarum ut serviant Nabuchodonosor regi Babylonis et servient ei insuper et bestias terrae dedi ei
JER|28|15|et dixit Hieremias propheta ad Ananiam prophetam audi Anania non misit te Dominus et tu confidere fecisti populum istum in mendacio
JER|28|16|idcirco haec dicit Dominus ecce emittam te a facie terrae hoc anno morieris adversum Dominum enim locutus es
JER|28|17|et mortuus est Ananias propheta in anno illo mense septimo
JER|29|1|et haec sunt verba libri quae misit Hieremias propheta de Hierusalem ad reliquias seniorum transmigrationis et ad sacerdotes et ad prophetas et ad omnem populum quem transduxerat Nabuchodonosor de Hierusalem in Babylonem
JER|29|2|postquam egressus est Iechonias rex et domina et eunuchi et principes Iuda et Hierusalem et faber et inclusor de Hierusalem
JER|29|3|in manu Ellasa filii Saphan et Gamaliae filii Helciae quos misit Sedecias rex Iuda ad Nabuchodonosor regem Babylonis in Babylonem dicens
JER|29|4|haec dicit Dominus exercituum Deus Israhel omni transmigrationi quam transtuli de Hierusalem in Babylonem
JER|29|5|aedificate domos et habitate et plantate hortos et comedite fructum eorum
JER|29|6|accipite uxores et generate filios et filias date filiis vestris uxores et filias vestras date viris et pariant filios et filias et multiplicamini ibi et nolite esse pauci numero
JER|29|7|et quaerite pacem civitatis ad quam transmigrare vos feci et orate pro ea ad Dominum quia in pace illius erit pax vobis
JER|29|8|haec enim dicit Dominus exercituum Deus Israhel non vos inducant prophetae vestri qui sunt in medio vestrum et divini vestri et ne adtendatis ad somnia vestra quae vos somniatis
JER|29|9|quia falso ipsi prophetant vobis in nomine meo et non misi eos dicit Dominus
JER|29|10|quia haec dicit Dominus cum coeperint impleri in Babylone septuaginta anni visitabo vos et suscitabo super vos verbum meum bonum ut reducam vos ad locum istum
JER|29|11|ego enim scio cogitationes quas cogito super vos ait Dominus cogitationes pacis et non adflictionis ut dem vobis finem et patientiam
JER|29|12|et invocabitis me et ibitis et orabitis me et exaudiam vos
JER|29|13|quaeretis me et invenietis cum quaesieritis me in toto corde vestro
JER|29|14|et inveniar a vobis ait Dominus et reducam captivitatem vestram et congregabo vos de universis gentibus et de cunctis locis ad quae expuli vos dicit Dominus et reverti vos faciam de loco ad quem transmigrare vos feci
JER|29|15|quia dixistis suscitavit nobis Dominus prophetas in Babylone
JER|29|16|quia haec dicit Dominus ad regem qui sedet super solium David et ad omnem populum habitatorem urbis huius ad fratres vestros qui non sunt egressi vobiscum in transmigrationem
JER|29|17|haec dicit Dominus exercituum ecce mittam in eis gladium et famem et pestem et ponam eos quasi ficus malas quae comedi non possunt eo quod pessimae sint
JER|29|18|et persequar eos in gladio in fame et in pestilentia et dabo eos in vexationem universis regnis terrae in maledictionem et in stuporem et in sibilum et in obprobrium cunctis gentibus ad quas ego eieci eos
JER|29|19|eo quod non audierint verba mea dicit Dominus quae misi ad eos per servos meos prophetas de nocte consurgens et mittens et non audistis dicit Dominus
JER|29|20|vos ergo audite verbum Domini omnis transmigratio quam emisi de Hierusalem in Babylonem
JER|29|21|haec dicit Dominus exercituum Deus Israhel ad Ahab filium Culia et ad Sedeciam filium Maasiae qui prophetant vobis in nomine meo mendaciter ecce ego tradam eos in manu Nabuchodonosor regis Babylonis et percutiet eos in oculis vestris
JER|29|22|et adsumetur ex eis maledictio omni transmigrationi Iuda quae est in Babylone dicentium ponat te Dominus sicut Sedeciam et sicut Ahab quos frixit rex Babylonis in igne
JER|29|23|pro eo quod fecerint stultitiam in Israhel et moechati sunt in uxores amicorum suorum et locuti sunt verbum in nomine meo mendaciter quod non mandavi eis ego sum iudex et testis dicit Dominus
JER|29|24|et ad Semeiam Neelamiten dices
JER|29|25|haec dicit Dominus exercituum Deus Israhel pro eo quod misisti in nomine tuo libros ad omnem populum qui est in Hierusalem et ad Sophoniam filium Maasiae sacerdotem et ad universos sacerdotes dicens
JER|29|26|Dominus dedit te sacerdotem pro Ioiadae sacerdote ut sis dux in domo Domini super omnem virum arrepticium et prophetantem ut mittas eum in nervum et in carcerem
JER|29|27|et nunc quare non increpasti Hieremiam Anathothiten qui prophetat vobis
JER|29|28|quia super hoc misit ad nos in Babylonem dicens longum est aedificate domos et habitate et plantate hortos et comedite fructum eorum
JER|29|29|legit ergo Sophonias sacerdos librum istum in auribus Hieremiae prophetae
JER|29|30|et factum est verbum Domini ad Hieremiam dicens
JER|29|31|mitte ad omnem transmigrationem dicens haec dicit Dominus ad Semeiam Neelamiten pro eo quod prophetavit vobis Semeias et ego non misi eum et fecit vos confidere in mendacio
JER|29|32|idcirco haec dicit Dominus ecce ego visitabo super Semeiam Neelamiten et super semen eius non erit ei vir sedens in medio populi huius et non videbit bonum quod ego faciam populo meo ait Dominus quia praevaricationem locutus est adversum Dominum
JER|30|1|hoc verbum quod factum est ad Hieremiam a Domino dicens
JER|30|2|haec dicit Dominus Deus Israhel dicens scribe tibi omnia verba quae locutus sum ad te in libro
JER|30|3|ecce enim dies veniunt dicit Dominus et convertam conversionem populi mei Israhel et Iuda ait Dominus et convertam eos ad terram quam dedi patribus eorum et possidebunt eam
JER|30|4|et haec verba quae locutus est Dominus ad Israhel et ad Iudam
JER|30|5|quoniam haec dicit Dominus vocem terroris audivimus formido et non est pax
JER|30|6|interrogate et videte si generat masculus quare ergo vidi omnis viri manum super lumbum suum quasi parientis et conversae sunt universae facies in auruginem
JER|30|7|vae quia magna dies illa nec est similis eius tempusque tribulationis est Iacob et ex ipso salvabitur
JER|30|8|et erit in die illa ait Dominus exercituum conteram iugum eius de collo tuo et vincula illius disrumpam et non dominabuntur ei amplius alieni
JER|30|9|sed servient Domino Deo suo et David regi suo quem suscitabo eis
JER|30|10|tu ergo ne timeas serve meus Iacob ait Dominus neque paveas Israhel quia ecce ego salvo te de terra longinqua et semen tuum de terra captivitatis eorum et revertetur Iacob et quiescet et cunctis affluet et non erit quem formidet
JER|30|11|quoniam tecum ego sum ait Dominus ut salvem te faciam enim consummationem in cunctis gentibus in quibus dispersi te te autem non faciam in consummationem sed castigabo te in iudicio ut non tibi videaris innoxius
JER|30|12|quia haec dicit Dominus insanabilis fractura tua pessima plaga tua
JER|30|13|non est qui iudicet iudicium tuum ad alligandum curationum utilitas non est tibi
JER|30|14|omnes amatores tui obliti sunt tui te non quaerent plaga enim inimici percussi te castigatione crudeli propter multitudinem iniquitatis tuae dura facta sunt peccata tua
JER|30|15|quid clamas super contritione tua insanabilis est dolor tuus propter multitudinem iniquitatis tuae et dura peccata tua feci haec tibi
JER|30|16|propterea omnes qui comedunt te devorabuntur et universi hostes tui in captivitatem ducentur et qui te vastant vastabuntur cunctosque praedatores tuos dabo in praedam
JER|30|17|obducam enim cicatricem tibi et a vulneribus tuis sanabo te dicit Dominus quia Eiectam vocaverunt te Sion haec est quae non habebat requirentem
JER|30|18|haec dicit Dominus ecce ego convertam conversionem tabernaculorum Iacob et tectis eius miserebor et aedificabitur civitas in excelso suo et templum iuxta ordinem suum fundabitur
JER|30|19|et egredietur de eis laus voxque ludentium et multiplicabo eos et non inminuentur et glorificabo eos et non adtenuabuntur
JER|30|20|et erunt filii eius sicut a principio et coetus eius coram me permanebit et visitabo adversum omnes qui tribulant eum
JER|30|21|et erit dux eius ex eo et princeps de medio eius producetur et adplicabo eum et accedet ad me quis enim iste est qui adplicet cor suum ut adpropinquet mihi ait Dominus
JER|30|22|et eritis mihi in populum et ego ero vobis in Deum
JER|30|23|ecce turbo Domini furor egrediens procella ruens in capite impiorum conquiescet
JER|30|24|non avertet iram indignationis Dominus donec faciat et conpleat cogitationem cordis sui in novissimo dierum intellegetis ea
JER|31|1|in tempore illo dicit Dominus ero Deus universis cognationibus Israhel et ipsi erunt mihi in populum
JER|31|2|haec dicit Dominus invenit gratiam in deserto populus qui remanserat gladio vadet ad requiem suam Israhel
JER|31|3|longe Dominus apparuit mihi et in caritate perpetua dilexi te ideo adtraxi te miserans
JER|31|4|rursumque aedificabo te et aedificaberis virgo Israhel adhuc ornaberis tympanis tuis et egredieris in choro ludentium
JER|31|5|adhuc plantabis vineas in montibus Samariae plantabunt plantantes et donec tempus veniat non vindemiabunt
JER|31|6|quia erit dies in qua clamabunt custodes in monte Ephraim surgite et ascendamus in Sion ad Dominum Deum nostrum
JER|31|7|quia haec dicit Dominus exultate in laetitia Iacob et hinnite contra caput gentium personate canite et dicite salva Domine populum tuum reliquias Israhel
JER|31|8|ecce ego adducam eos de terra aquilonis et congregabo eos ab extremis terrae inter quos erunt caecus et claudus et praegnans et pariens simul coetus magnus revertentium huc
JER|31|9|in fletu venient et in precibus deducam eos et adducam eos per torrentes aquarum in via recta et non inpingent in ea quia factus sum Israheli pater et Ephraim primogenitus meus est
JER|31|10|audite verbum Domini gentes et adnuntiate insulis quae procul sunt et dicite qui dispersit Israhel congregabit eum et custodiet eum sicut pastor gregem suum
JER|31|11|redemit enim Dominus Iacob et liberavit eum de manu potentioris
JER|31|12|et venient et laudabunt in monte Sion et confluent ad bona Domini super frumento et vino et oleo et fetu pecorum et armentorum eritque anima eorum quasi hortus inriguus et ultra non esurient
JER|31|13|tunc laetabitur virgo in choro iuvenes et senes simul et convertam luctum eorum in gaudium et consolabor eos et laetificabo a dolore suo
JER|31|14|et inebriabo animam sacerdotum pinguedine et populus meus bonis meis adimplebitur ait Dominus
JER|31|15|haec dicit Dominus vox in excelso audita est lamentationis fletus et luctus Rachel plorantis filios suos et nolentis consolari super eis quia non sunt
JER|31|16|haec dicit Dominus quiescat vox tua a ploratu et oculi tui a lacrimis quia est merces operi tuo ait Dominus et revertentur de terra inimici
JER|31|17|et est spes novissimis tuis ait Dominus et revertentur filii ad terminos suos
JER|31|18|audiens audivi Ephraim transmigrantem castigasti me et eruditus sum quasi iuvenculus indomitus converte me et revertar quia tu Dominus Deus meus
JER|31|19|postquam enim convertisti me egi paenitentiam et postquam ostendisti mihi percussi femur meum confusus sum et erubui quoniam sustinui obprobrium adulescentiae meae
JER|31|20|si filius honorabilis mihi Ephraim si puer delicatus quia ex quo locutus sum de eo adhuc recordabor eius idcirco conturbata sunt viscera mea super eum miserans miserebor eius ait Dominus
JER|31|21|statue tibi speculam pone tibi amaritudines dirige cor tuum in viam directam in qua ambulasti revertere virgo Israhel revertere ad civitates tuas istas
JER|31|22|usquequo deliciis dissolveris filia vaga quia creavit Dominus novum super terram femina circumdabit virum
JER|31|23|haec dicit Dominus exercituum Deus Israhel adhuc dicent verbum istud in terra Iuda et in urbibus eius cum convertero captivitatem eorum benedicat tibi Dominus pulchritudo iustitiae mons sanctus
JER|31|24|et habitabunt in eo Iudas et omnes civitates eius simul agricolae et minantes greges
JER|31|25|quia inebriavi animam lassam et omnem animam esurientem saturavi
JER|31|26|ideo quasi de somno suscitatus sum et vidi et somnus meus dulcis mihi
JER|31|27|ecce dies veniunt dicit Dominus et seminabo domum Israhel et domum Iuda semine hominis et semine iumentorum
JER|31|28|et sicut vigilavi super eos ut evellerem et demolirer et dissiparem et disperderem et adfligerem sic vigilabo super eos ut aedificem et plantem ait Dominus
JER|31|29|in diebus illis non dicent ultra patres comederunt uvam acerbam et dentes filiorum obstipuerunt
JER|31|30|sed unusquisque in iniquitate sua morietur omnis homo qui comederit uvam acerbam obstupescent dentes eius
JER|31|31|ecce dies veniunt dicit Dominus et feriam domui Israhel et domui Iuda foedus novum
JER|31|32|non secundum pactum quod pepigi cum patribus vestris in die qua adprehendi manum eorum ut educerem eos de terra Aegypti pactum quod irritum fecerunt et ego dominatus sum eorum dicit Dominus
JER|31|33|sed hoc erit pactum quod feriam cum domo Israhel post dies illos dicit Dominus dabo legem meam in visceribus eorum et in corde eorum scribam eam et ero eis in Deum et ipsi erunt mihi in populum
JER|31|34|et non docebunt ultra vir proximum suum et vir fratrem suum dicens cognoscite Dominum omnes enim cognoscent me a minimo eorum usque ad maximum ait Dominus quia propitiabor iniquitati eorum et peccati eorum non ero memor amplius
JER|31|35|haec dicit Dominus qui dat solem in lumine diei ordinem lunae et stellarum in lumine noctis qui turbat mare et sonant fluctus eius Dominus exercituum nomen illi
JER|31|36|si defecerint leges istae coram me dicit Dominus tunc et semen Israhel deficiet ut non sit gens coram me cunctis diebus
JER|31|37|haec dicit Dominus si mensurari potuerint caeli sursum et investigari fundamenta terrae deorsum et ego abiciam universum semen Israhel propter omnia quae fecerunt dicit Dominus
JER|31|38|ecce dies veniunt dicit Dominus et aedificabitur civitas Domino a turre Ananehel usque ad portam Anguli
JER|31|39|et exibit ultra norma mensurae in conspectu eius super collem Gareb et circuibit Goatha
JER|31|40|et omnem vallem cadaverum et cineris et universam regionem mortis usque ad torrentem Cedron et usque ad angulum portae Equorum orientalis sanctum Domini non evelletur et non destruetur ultra in perpetuum
JER|32|1|verbum quod factum est ad Hieremiam a Domino in anno decimo Sedeciae regis Iuda ipse est annus octavusdecimus Nabuchodonosor
JER|32|2|tunc exercitus regis Babylonis obsidebat Hierusalem et Hieremias propheta erat clausus in atrio carceris qui erat in domo regis Iuda
JER|32|3|clauserat enim eum Sedecias rex Iuda dicens quare vaticinaris dicens haec dicit Dominus ecce ego dabo civitatem istam in manu regis Babylonis et capiet eam
JER|32|4|et Sedecias rex Iuda non effugiet de manu Chaldeorum sed tradetur in manu regis Babylonis et loquetur os eius cum ore illius et oculi eius oculos illius videbunt
JER|32|5|et in Babylonem ducet Sedeciam et ibi erit donec visitem eum ait Dominus si autem dimicaveritis adversum Chaldeos nihil prosperum habebitis
JER|32|6|et dixit Hieremias factum est verbum Domini ad me dicens
JER|32|7|ecce Anamehel filius Sellum patruelis tuus veniet ad te dicens eme tibi agrum meum qui est in Anathoth tibi enim conpetit ex propinquitate ut emas
JER|32|8|et venit ad me Anamehel filius patrui mei secundum verbum Domini ad vestibulum carceris et ait ad me posside agrum meum qui est in Anathoth in terra Beniamin quia tibi conpetit hereditas et tu propinquus ut possideas intellexi autem quod verbum Domini esset
JER|32|9|et emi agrum ab Anamehel filio patrui mei qui est in Anathoth et adpendi ei argentum septem stateres et decem argenteos
JER|32|10|et scripsi in libro et signavi et adhibui testes et adpendi argentum in statera
JER|32|11|et accepi librum possessionis signatum stipulationes et rata et signa forinsecus
JER|32|12|et dedi librum possessionis Baruch filio Neri filii Maasiae in oculis Anamehel patruelis mei et in oculis testium qui scripti erant in libro emptionis in oculis omnium Iudaeorum qui sedebant in atrio carceris
JER|32|13|et praecepi Baruch coram eis dicens
JER|32|14|haec dicit Dominus exercituum Deus Israhel sume libros istos librum emptionis hunc signatum et librum hunc qui apertus est et pones illos in vase fictili ut permanere possint diebus multis
JER|32|15|haec enim dicit Dominus exercituum Deus Israhel adhuc possidebuntur domus et agri et vineae in terra ista
JER|32|16|et oravi ad Dominum postquam tradidi librum possessionis Baruch filio Neri dicens
JER|32|17|heu heu heu Domine Deus ecce tu fecisti caelum et terram in fortitudine tua magna et in brachio tuo extento non erit tibi difficile omne verbum
JER|32|18|qui facis misericordiam in milibus et reddes iniquitatem patrum in sinu filiorum eorum post eos fortissime magne potens Dominus exercituum nomen tibi
JER|32|19|magnus consilio et inconprehensibilis cogitatu cuius oculi aperti sunt super omnes vias filiorum Adam ut reddas unicuique secundum vias suas et secundum fructum adinventionum eius
JER|32|20|qui posuisti signa et portenta in terra Aegypti usque ad diem hanc et in Israhel et in hominibus et fecisti tibi nomen sicut est dies haec
JER|32|21|et eduxisti populum tuum Israhel de terra Aegypti in signis et in portentis et in manu robusta et in brachio extento et in terrore magno
JER|32|22|et dedisti eis terram hanc quam iurasti patribus eorum ut dares eis terram fluentem lacte et melle
JER|32|23|et ingressi sunt et possederunt eam et non oboedierunt voci tuae et in lege tua non ambulaverunt omnia quae mandasti eis ut facerent non fecerunt et evenerunt eis omnia mala haec
JER|32|24|ecce munitiones extructae sunt adversum civitatem ut capiatur et urbs data est in manu Chaldeorum qui proeliantur adversum eam a facie gladii et famis et pestilentiae et quaecumque locutus es acciderunt ut ipse tu cernis
JER|32|25|et tu dicis mihi Domine Deus eme agrum argento et adhibe testes cum urbs data sit in manu Chaldeorum
JER|32|26|et factum est verbum Domini ad Hieremiam dicens
JER|32|27|ecce ego Dominus Deus universae carnis numquid mihi difficile erit omne verbum
JER|32|28|propterea haec dicit Dominus ecce ego tradam civitatem istam in manu Chaldeorum et in manu regis Babylonis et capiet eam
JER|32|29|et venient Chaldei proeliantes adversum urbem hanc et succendent eam igni et conburent eam et domos in quarum domatibus sacrificabant Baal et libabant diis alienis libamina ad inritandum me
JER|32|30|erant enim filii Israhel et filii Iuda iugiter facientes malum in oculis meis ab adulescentia sua filii Israhel qui usque nunc exacerbant me in opere manuum suarum dicit Dominus
JER|32|31|quia in furore et in indignatione mea facta est mihi civitas haec a die qua aedificaverunt eam usque ad diem istam qua aufertur de conspectu meo
JER|32|32|propter malitiam filiorum Israhel et filiorum Iuda quam fecerunt ad iracundiam me provocantes ipsi et reges eorum principes eorum et sacerdotes et prophetae eorum vir Iuda et habitatores Hierusalem
JER|32|33|et verterunt ad me terga et non facies cum docerem eos diluculo et erudirem et nollent audire ut acciperent disciplinam
JER|32|34|et posuerunt idola sua in domo in qua invocatum est nomen meum ut polluerent eam
JER|32|35|et aedificaverunt excelsa Baal quae sunt in valle filii Ennom ut initiarent filios suos et filias suas Moloch quod non mandavi eis nec ascendit in cor meum ut facerent abominationem hanc et in peccatum deducerent Iudam
JER|32|36|et nunc propter ista haec dicit Dominus Deus Israhel ad civitatem hanc de qua vos dicitis quod tradatur in manu regis Babylonis in gladio et in fame et in peste
JER|32|37|ecce ego congregabo eos de universis terris ad quas eieci eos in furore meo et in ira mea et in indignatione grandi et reducam eos ad locum istum et habitare eos faciam confidenter
JER|32|38|et erunt mihi in populum et ego ero eis in Deum
JER|32|39|et dabo eis cor unum et viam unam ut timeant me universis diebus et bene sit eis et filiis eorum post eos
JER|32|40|et feriam eis pactum sempiternum et non desinam eis benefacere et timorem meum dabo in corde eorum ut non recedant a me
JER|32|41|et laetabor super eis cum bene eis fecero et plantabo eos in terra ista in veritate in toto corde meo et in tota anima mea
JER|32|42|quia haec dicit Dominus sicut adduxi super populum istum omne malum hoc grande sic adducam super eos omne bonum quod ego loquor ad eos
JER|32|43|et possidebuntur agri in terra ista de qua vos dicitis quod deserta sit eo quod non remanserit homo et iumentum et data sit in manu Chaldeorum
JER|32|44|agri pecunia ementur et scribentur in libro et inprimetur signum et testis adhibebitur in terra Beniamin et in circuitu Hierusalem in civitatibus Iuda et in civitatibus montanis et in civitatibus campestribus et in civitatibus quae ad austrum sunt quia convertam captivitatem eorum ait Dominus
JER|33|1|et factum est verbum Domini ad Hieremiam secundo cum adhuc clausus esset in atrio carceris dicens
JER|33|2|haec dicit Dominus qui facturus est Dominus et formaturus illud et paraturus Dominus nomen eius
JER|33|3|clama ad me et exaudiam te et adnuntiabo tibi grandia et firma quae nescis
JER|33|4|quia haec dicit Dominus Deus Israhel ad domos urbis huius et ad domos regis Iuda quae destructae sunt et ad munitiones et gladium
JER|33|5|venientium ut dimicent cum Chaldeis et impleant eas cadaveribus hominum quas percussi in furore meo et in indignatione mea abscondens faciem meam a civitate hac propter omnem malitiam eorum
JER|33|6|ecce ego obducam ei cicatricem et sanitatem et curabo eos et revelabo illis deprecationem pacis et veritatis
JER|33|7|et convertam conversionem Iuda et conversionem Hierusalem et aedificabo eos sicut a principio
JER|33|8|et emundabo illos ab omni iniquitate sua in qua peccaverunt mihi et propitius ero cunctis iniquitatibus eorum in quibus deliquerunt mihi et spreverunt me
JER|33|9|et erit mihi in nomen et in gaudium et in laudem et in exultationem cunctis gentibus terrae quae audierint omnia bona quae ego facturus sum eis et pavebunt et turbabuntur in universis bonis et in omni pace quam ego faciam ei
JER|33|10|haec dicit Dominus adhuc audietur in loco isto quem vos dicitis esse desertum eo quod non sit homo et iumentum in civitatibus Iuda et foris Hierusalem quae desolatae sunt absque homine et absque habitatore et absque pecore
JER|33|11|vox gaudii et vox laetitiae vox sponsi et vox sponsae vox dicentium confitemini Domino exercituum quoniam bonus Dominus quoniam in aeternum misericordia eius et portantium vota in domum Domini reducam enim conversionem terrae sicut a principio dicit Dominus
JER|33|12|haec dicit Dominus exercituum adhuc erit in loco isto deserto absque homine et absque iumento et in cunctis civitatibus eius habitaculum pastorum accubantium gregum
JER|33|13|in civitatibus montuosis et in civitatibus campestribus et in civitatibus quae ad austrum sunt et in terra Beniamin et in circuitu Hierusalem et in civitatibus Iuda adhuc transibunt greges ad manum numerantis ait Dominus
JER|33|14|ecce dies veniunt dicit Dominus et suscitabo verbum bonum quod locutus sum ad domum Israhel et ad domum Iuda
JER|33|15|in diebus illis et in tempore illo germinare faciam David germen iustitiae et faciet iudicium et iustitiam in terra
JER|33|16|in diebus illis salvabitur Iuda et Hierusalem habitabit confidenter et hoc est quod vocabit eam Dominus iustus noster
JER|33|17|quia haec dicit Dominus non interibit de David vir qui sedeat super thronum domus Israhel
JER|33|18|et de sacerdotibus et Levitis non interibit vir a facie mea qui offerat holocaustomata et incendat sacrificium et caedat victimas cunctis diebus
JER|33|19|et factum est verbum Domini ad Hieremiam dicens
JER|33|20|haec dicit Dominus si irritum fieri potest pactum meum cum die et pactum meum cum nocte ut non sit dies et nox in tempore suo
JER|33|21|et pactum meum irritum esse poterit cum David servo meo ut non sit ex eo filius qui regnet in throno eius et Levitae et sacerdotes ministri mei
JER|33|22|sicuti numerari non possunt stellae caeli et metiri harena maris sic multiplicabo semen David servi mei et Levitas ministros meos
JER|33|23|et factum est verbum Domini ad Hieremiam dicens
JER|33|24|numquid non vidisti quid populus hic locutus sit dicens duae cognationes quas elegerat Dominus abiectae sunt et populum meum despexerunt eo quod non sit ultra gens coram eis
JER|33|25|haec dicit Dominus si pactum meum inter diem et noctem et leges caelo et terrae non posui
JER|33|26|equidem et semen Iacob et David servi mei proiciam ut non adsumam de semine eius principes seminis Abraham et Isaac et Iacob reducam enim conversionem eorum et miserebor eis
JER|34|1|verbum quod factum est ad Hieremiam a Domino quando Nabuchodonosor rex Babylonis et omnis exercitus eius universaque regna terrae quae erant sub potestate manus eius et omnes populi bellabant contra Hierusalem et contra omnes urbes eius dicens
JER|34|2|haec dicit Dominus Deus Israhel vade et loquere ad Sedeciam regem Iuda et dices ad eum haec dicit Dominus ecce ego tradam civitatem hanc in manu regis Babylonis et succendet eam igni
JER|34|3|et tu non effugies de manu eius sed conprehensione capieris et in manu eius traderis et oculi tui oculos regis Babylonis videbunt et os eius cum ore tuo loquetur et Babylonem introibis
JER|34|4|attamen audi verbum Domini Sedecia rex Iuda haec dicit Dominus ad te non morieris in gladio
JER|34|5|sed in pace morieris et secundum conbustiones patrum tuorum regum priorum qui fuerunt ante te sic conburent te et vae domine plangent te quia verbum ego locutus sum dicit Dominus
JER|34|6|et locutus est Hieremias propheta ad Sedeciam regem Iuda universa verba haec in Hierusalem
JER|34|7|et exercitus regis Babylonis pugnabat contra Hierusalem et contra omnes civitates Iuda quae reliquae erant contra Lachis et contra Azeca haec enim supererant de civitatibus Iuda urbes munitae
JER|34|8|verbum quod factum est ad Hieremiam a Domino postquam percussit rex Sedecias foedus cum omni populo in Hierusalem praedicans
JER|34|9|ut dimitteret unusquisque servum suum et unusquisque ancillam suam hebraeum et hebraeam liberos et nequaquam dominarentur eis id est in Iudaeo et fratre suo
JER|34|10|audierunt ergo omnes principes et universus populus qui inierant pactum ut dimitteret unusquisque servum suum et unusquisque ancillam suam liberos et ultra non dominarentur in eis audierunt igitur et dimiserunt
JER|34|11|et conversi sunt deinceps et retraxerunt servos et ancillas suas quos dimiserant liberos et subiugaverunt in famulos et in famulas
JER|34|12|et factum est verbum Domini ad Hieremiam a Domino dicens
JER|34|13|haec dicit Dominus Deus Israhel ego percussi foedus cum patribus vestris in die qua eduxi eos de terra Aegypti de domo servitutis dicens
JER|34|14|cum conpleti fuerint septem anni dimittat unusquisque fratrem suum hebraeum qui venditus est ei et serviet tibi sex annis et dimittes eum a te liberum et non audierunt patres vestri me nec inclinaverunt aurem suam
JER|34|15|et conversi estis vos hodie et fecistis quod rectum est in oculis meis ut praedicaretis libertatem unusquisque ad amicum suum et inistis pactum in conspectu meo in domo in qua invocatum est nomen meum super eam
JER|34|16|et reversi estis et commaculastis nomen meum et reduxistis unusquisque servum suum et unusquisque ancillam suam quos dimiseratis ut essent liberi et suae potestatis et subiugastis eos ut sint vobis servi et ancillae
JER|34|17|propterea haec dicit Dominus vos non audistis me ut praedicaretis libertatem unusquisque fratri suo et unusquisque amico suo ecce ego praedico libertatem ait Dominus ad gladium et pestem et famem et dabo vos in commotionem cunctis regnis terrae
JER|34|18|et dabo viros qui praevaricantur foedus meum et non observaverunt verba foederis quibus adsensi sunt in conspectu meo vitulum quem ceciderunt in duas partes et transierunt inter divisiones eius
JER|34|19|principes Iuda et principes Hierusalem eunuchi et sacerdotes et omnis populus terrae qui transierunt inter divisiones vituli
JER|34|20|et dabo eos in manu inimicorum suorum et in manu quaerentium animam eorum et erit morticinum eorum in escam volucribus caeli et bestiis terrae
JER|34|21|et Sedeciam regem Iuda et principes eius dabo in manu inimicorum suorum et in manu quaerentium animam eorum et in manu exercituum regis Babylonis qui recesserunt a vobis
JER|34|22|ecce ego praecipio dicit Dominus et reducam eos in civitatem hanc et proeliabuntur adversum eam et capient eam et incendent igni et civitates Iuda dabo in solitudinem eo quod non sit habitator
JER|35|1|verbum quod factum est ad Hieremiam a Domino in diebus Ioachim filii Iosiae regis Iuda dicens
JER|35|2|vade ad domum Rechabitarum et loquere eis et introduces eos in domum Domini in unam exedram thesaurorum et dabis eis bibere vinum
JER|35|3|et adsumpsi Iezoniam filium Hieremiae filii Absaniae et fratres eius et omnes filios eius et universam domum Rechabitarum
JER|35|4|et introduxi eos in domum Domini ad gazofilacium filiorum Anan filii Hiegedeliae hominis Dei quod erat iuxta gazofilacium principum super thesaurum Maasiae filii Sellum qui erat custos vestibuli
JER|35|5|et posui coram filiis domus Rechabitarum scyphos plenos vino et calices et dixi ad eos bibite vinum
JER|35|6|qui responderunt non bibemus vinum quia Ionadab filius Rechab pater noster praecepit nobis dicens non bibetis vinum vos et filii vestri usque in sempiternum
JER|35|7|et domum non aedificabitis et sementem non seretis et vineas non plantabitis nec habebitis sed in tabernaculis habitabitis cunctis diebus vestris ut vivatis diebus multis super faciem terrae in qua vos peregrinamini
JER|35|8|oboedivimus ergo voci Ionadab filii Rechab patris nostri in omnibus quae praecepit nobis ita ut non biberemus vinum cunctis diebus nostris nos et mulieres nostrae filii et filiae nostrae
JER|35|9|et non aedificaremus domos ad habitandum et vineam et agrum et sementem non habuimus
JER|35|10|sed habitavimus in tabernaculis et oboedientes fecimus iuxta omnia quae praecepit nobis Ionadab pater noster
JER|35|11|cum autem ascendisset Nabuchodonosor rex Babylonis ad terram nostram diximus venite et ingrediamur Hierusalem a facie exercitus Chaldeorum et a facie exercitus Syriae et mansimus in Hierusalem
JER|35|12|et factum est verbum Domini ad Hieremiam dicens
JER|35|13|haec dicit Dominus exercituum Deus Israhel vade et dic viris Iuda et habitatoribus Hierusalem numquid non recipietis disciplinam ut oboediatis verbis meis dicit Dominus
JER|35|14|praevaluerunt sermones Ionadab filii Rechab quos praecepit filiis suis ut non biberent vinum et non biberunt usque ad diem hanc quia oboedierunt praecepto patris sui ego autem locutus sum ad vos de mane consurgens et loquens et non oboedistis mihi
JER|35|15|misique ad vos omnes servos meos prophetas consurgens diluculo mittensque et dicens convertimini unusquisque a via sua pessima et bona facite studia vestra et nolite sequi deos alienos neque colatis eos et habitabitis in terra quam dedi vobis et patribus vestris et non inclinastis aurem vestram neque audistis me
JER|35|16|firmaverunt igitur filii Ionadab filii Rechab praeceptum patris sui quod praeceperat eis populus autem iste non oboedivit mihi
JER|35|17|idcirco haec dicit Dominus exercituum Deus Israhel ecce ego adduco super Iudam et super omnes habitatores Hierusalem universam adflictionem quam locutus sum adversum eos eo quod locutus sum ad illos et non audierunt vocavi illos et non responderunt mihi
JER|35|18|domui autem Rechabitarum dixit Hieremias haec dicit Dominus exercituum Deus Israhel pro eo quod oboedistis praecepto Ionadab patris vestri et custodistis omnia mandata eius et fecistis universa quae praecepit vobis
JER|35|19|propterea haec dicit Dominus exercituum Deus Israhel non deficiet vir de stirpe Ionadab filii Rechab stans in conspectu meo cunctis diebus
JER|36|1|et factum est in anno quarto Ioachim filii Iosiae regis Iuda factum est verbum hoc ad Hieremiam a Domino dicens
JER|36|2|tolle volumen libri et scribes in eo omnia verba quae locutus sum tibi adversum Israhel et Iudam et adversum omnes gentes a die qua locutus sum ad te ex diebus Iosiae usque ad diem hanc
JER|36|3|si forte audiente domo Iuda universa mala quae ego cogito facere eis revertatur unusquisque a via sua pessima et propitius ero iniquitati et peccato eorum
JER|36|4|vocavit ergo Hieremias Baruch filium Neriae et scripsit Baruch ex ore Hieremiae omnes sermones Domini quos locutus est ad eum in volumine libri
JER|36|5|et praecepit Hieremias Baruch dicens ego clausus sum nec valeo ingredi domum Domini
JER|36|6|ingredere ergo tu et lege de volumine in quo scripsisti ex ore meo verba Domini audiente populo in domo Domini in die ieiunii insuper et audiente universo Iuda qui veniunt de civitatibus suis leges eis
JER|36|7|si forte cadat oratio eorum in conspectu Domini et revertatur unusquisque a via sua pessima quoniam magnus furor et indignatio quam locutus est Dominus adversum populum hunc
JER|36|8|et fecit Baruch filius Neriae iuxta omnia quae praeceperat ei Hieremias propheta legens ex volumine sermones Domini in domo Domini
JER|36|9|factum est autem in anno quinto Ioachim filii Iosiae regis Iuda in mense nono praedicaverunt ieiunium in conspectu Domini omni populo in Hierusalem et universae multitudini quae confluxerat de civitatibus Iuda in Hierusalem
JER|36|10|legitque Baruch ex volumine sermones Hieremiae in domo Domini in gazofilacio Gamariae filii Saphan scribae in vestibulo superiori in introitu portae novae domus Domini audiente omni populo
JER|36|11|cumque audisset Micheas filius Gamariae filii Saphan omnes sermones Domini ex libro
JER|36|12|descendit in domum regis ad gazofilacium scribae et ecce ibi omnes principes sedebant Elisama scriba et Dalaias filius Semeiae et Elnathan filius Achobor et Gamarias filius Saphan et Sedecias filius Ananiae et universi principes
JER|36|13|et nuntiavit eis Micheas omnia verba quae audivit legente Baruch ex volumine in auribus populi
JER|36|14|miserunt itaque omnes principes ad Baruch Iudi filium Nathaniae filii Selemiae filii Chusi dicentes volumen ex quo legisti audiente populo sume in manu tua et veni tulit ergo Baruch filius Neriae volumen in manu sua et venit ad eos
JER|36|15|et dixerunt ad eum sede et lege haec in auribus nostris et legit Baruch in auribus eorum
JER|36|16|igitur cum audissent omnia verba obstipuerunt unusquisque ad proximum suum et dixerunt ad Baruch nuntiare debemus regi omnes sermones istos
JER|36|17|et interrogaverunt eum dicentes indica nobis quomodo scripsisti omnes sermones istos ex ore eius
JER|36|18|dixit autem eis Baruch ex ore suo loquebatur quasi legens ad me omnes sermones istos et ego scribebam in volumine atramento
JER|36|19|et dixerunt principes ad Baruch vade et abscondere tu et Hieremias et nemo sciat ubi sitis
JER|36|20|et ingressi sunt ad regem in atrium porro volumen commendaverunt in gazofilacio Elisamae scribae et nuntiaverunt audiente rege omnes sermones
JER|36|21|misitque rex Iudi ut sumeret volumen qui tollens illud de gazofilacio Elisamae scribae legit audiente rege et universis principibus qui stabant circa regem
JER|36|22|rex autem sedebat in domo hiemali in mense nono et posita erat arula coram eo plena prunis
JER|36|23|cumque legisset Iudi tres pagellas vel quattuor scidit illud scalpello scribae et proiecit in igne qui erat super arulam donec consumeretur omne volumen igni qui erat in arula
JER|36|24|et non timuerunt neque sciderunt vestimenta sua rex et omnes servi eius qui audierunt universos sermones istos
JER|36|25|verumtamen Elnathan et Dalaias et Gamarias contradixerunt regi ne conbureret librum et non audivit eos
JER|36|26|et praecepit rex Hieremahel filio Ammelech et Saraiae filio Ezrihel et Selemiae filio Abdehel ut conprehenderent Baruch scribam et Hieremiam prophetam abscondit autem eos Dominus
JER|36|27|et factum est verbum Domini ad Hieremiam postquam conbuserat rex volumen et sermones quos scripserat Baruch ex ore Hieremiae dicens
JER|36|28|rursum tolle volumen aliud et scribe in eo omnes sermones priores qui erant in volumine primo quod conbusit Ioachim rex Iuda
JER|36|29|et ad Ioachim regem Iuda dices haec dicit Dominus tu conbusisti volumen illud dicens quare scripsisti in eo adnuntians festinus veniet rex Babylonis et vastabit terram hanc et cessare faciet ex illa hominem et iumentum
JER|36|30|propterea haec dicit Dominus contra Ioachim regem Iuda non erit ex eo qui sedeat super solium David et cadaver eius proicietur ad aestum per diem et ad gelu per noctem
JER|36|31|et visitabo contra eum et contra semen eius et contra servos eius iniquitates suas et adducam super eos et super habitatores Hierusalem et super viros Iuda omne malum quod locutus sum ad eos et non audierunt
JER|36|32|Hieremias autem tulit volumen aliud et dedit illud Baruch filio Neriae scribae qui scripsit in eo ex ore Hieremiae omnes sermones libri quem conbuserat Ioachim rex Iuda igni et insuper additi sunt sermones multo plures quam ante fuerant
JER|37|1|et regnavit rex Sedecias filius Iosiae pro Iechonia filio Ioachim quem constituit regem Nabuchodonosor rex Babylonis in terra Iuda
JER|37|2|et non oboedivit ipse et servi eius et populus terrae verbis Domini quae locutus est in manu Hieremiae prophetae
JER|37|3|et misit rex Sedecias Iuchal filium Selemiae et Sophoniam filium Maasiae sacerdotem ad Hieremiam prophetam dicens ora pro nobis Dominum Deum nostrum
JER|37|4|Hieremias autem libere ambulabat in medio populi non enim miserant eum in custodiam carceris igitur exercitus Pharao egressus est Aegyptum et audientes Chaldei qui obsidebant Hierusalem huiuscemodi nuntium recesserunt ab Hierusalem
JER|37|5|et factum est verbum Domini ad Hieremiam prophetam dicens
JER|37|6|haec dicit Dominus Deus Israhel sic dicetis regi Iuda qui misit vos ad me ad interrogandum ecce exercitus Pharaonis qui egressus est vobis in auxilium revertetur in terram suam in Aegyptum
JER|37|7|et redient Chaldei et bellabunt contra civitatem hanc et capient eam et incendent igni
JER|37|8|haec dicit Dominus nolite decipere animas vestras dicentes euntes abibunt et recedent a nobis Chaldei quia non abibunt
JER|37|9|sed et si percusseritis omnem exercitum Chaldeorum qui proeliantur adversum vos et derelicti fuerint ex eis aliqui vulnerati singuli de tentorio suo consurgent et incendent civitatem hanc igni
JER|37|10|ergo cum recessisset exercitus Chaldeorum ab Hierusalem propter exercitum Pharaonis
JER|37|11|egressus est Hieremias de Hierusalem ut iret in terram Beniamin et divideret ibi possessionem in conspectu civium
JER|37|12|cumque pervenisset ad portam Beniamin erat ibi custos portae per vices nomine Hierias filius Selemiae filii Ananiae et adprehendit Hieremiam prophetam dicens ad Chaldeos profugis
JER|37|13|et respondit Hieremias falsum est non fugio ad Chaldeos et non audivit eum sed conprehendit Hierias Hieremiam et adduxit eum ad principes
JER|37|14|quam ob rem irati principes contra Hieremiam caesum eum miserunt in carcerem qui erat in domo Ionathan scribae ipse enim praepositus erat super carcerem
JER|37|15|itaque ingressus est Hieremias in domum laci et in ergastula et sedit ibi Hieremias diebus multis
JER|37|16|mittens autem rex Sedecias tulit eum et interrogavit in domo sua abscondite et dixit putasne est sermo a Domino et dixit Hieremias est et ait in manu regis Babylonis traderis
JER|37|17|et dixit Hieremias ad regem Sedeciam quid peccavi tibi et servis tuis et populo tuo quia misisti me in domum carceris
JER|37|18|ubi sunt prophetae vestri qui prophetabant vobis et dicebant non veniet rex Babylonis super vos et super terram hanc
JER|37|19|nunc ergo audi obsecro domine mi rex valeat deprecatio mea in conspectu tuo et ne me remittas in domum Ionathan scribae ne moriar ibi
JER|37|20|praecepit ergo rex Sedecias ut traderetur Hieremias in vestibulo carceris et daretur ei torta panis cotidie excepto pulmento donec consumerentur omnes panes de civitate et mansit Hieremias in vestibulo carceris
JER|38|1|audivit autem Saphatias filius Matthan et Gedelias filius Phassur et Iuchal filius Selemiae et Phassur filius Melchiae sermones quos Hieremias loquebatur ad omnem populum dicens
JER|38|2|haec dicit Dominus quicumque manserit in civitate hac morietur gladio et fame et peste qui autem profugerit ad Chaldeos vivet et erit anima eius sospes et vivens
JER|38|3|haec dicit Dominus tradenda tradetur civitas haec in manu exercitus regis Babylonis et capiet eam
JER|38|4|et dixerunt principes regi rogamus ut occidatur homo iste de industria enim dissolvit manus virorum bellantium qui remanserunt in civitate hac et manus universi populi loquens ad eos iuxta verba haec siquidem homo hic non quaerit pacem populi huius sed malum
JER|38|5|et dixit rex Sedecias ecce ipse in manibus vestris est nec enim fas est regem vobis quicquam negare
JER|38|6|tulerunt ergo Hieremiam et proiecerunt eum in lacu Melchiae filii Ammelech qui erat in vestibulo carceris et submiserunt Hieremiam in funibus et in lacum non erat aqua sed lutum descendit itaque Hieremias in caenum
JER|38|7|audivit autem Abdemelech Aethiops vir eunuchus qui erat in domo regis quod misissent Hieremiam in lacum porro rex sedebat in porta Beniamin
JER|38|8|et egressus est Abdemelech de domo regis et locutus est ad regem dicens
JER|38|9|domine mi rex malefecerunt viri isti omnia quaecumque perpetrarunt contra Hieremiam prophetam mittentes eum in lacum ut moriatur ibi fame non sunt enim panes ultra in civitate
JER|38|10|praecepit itaque rex Abdemelech Aethiopi dicens tolle tecum hinc triginta viros et leva Hieremiam prophetam de lacu antequam moriatur
JER|38|11|adsumptis ergo Abdemelech secum viris ingressus est domum regis quae erat sub cellario et tulit inde veteres pannos et antiqua quae conputruerant et submisit ea ad Hieremiam in lacum per funiculos
JER|38|12|dixitque Abdemelech Aethiops ad Hieremiam pone veteres pannos et haec scissa et putrida sub cubitu manuum tuarum et subter funes fecit ergo Hieremias sic
JER|38|13|et extraxerunt Hieremiam funibus et eduxerunt eum de lacu mansit autem Hieremias in vestibulo carceris
JER|38|14|et misit rex Sedecias et tulit ad se Hieremiam prophetam ad ostium tertium quod erat in domo Domini et dixit rex ad Hieremiam interrogo ego te sermonem ne abscondas a me aliquid
JER|38|15|dixit autem Hieremias ad Sedeciam si adnuntiavero tibi numquid non interficies me et si consilium tibi dedero non me audies
JER|38|16|iuravit ergo rex Sedecias Hieremiae clam dicens vivit Dominus qui fecit nobis animam hanc si occidero te et si tradidero te in manu virorum istorum qui quaerunt animam tuam
JER|38|17|et dixit Hieremias ad Sedeciam haec dicit Dominus exercituum Deus Israhel si profectus exieris ad principes regis Babylonis vivet anima tua et civitas haec non succendetur igni et salvus eris tu et domus tua
JER|38|18|si autem non exieris ad principes regis Babylonis tradetur civitas haec in manu Chaldeorum et succendent eam igni et tu non effugies de manu eorum
JER|38|19|et dixit rex Sedecias ad Hieremiam sollicitus sum propter Iudaeos qui transfugerunt ad Chaldeos ne forte tradar in manus eorum et inludant mihi
JER|38|20|respondit autem Hieremias non te tradent audi quaeso vocem Domini quam ego loquor ad te et bene tibi erit et vivet anima tua
JER|38|21|quod si nolueris egredi iste est sermo quem ostendit mihi Dominus
JER|38|22|ecce omnes mulieres quae remanserunt in domo regis Iuda educentur ad principes regis Babylonis et ipsae dicent seduxerunt te et praevaluerunt adversum te viri pacifici tui demerserunt in caeno et lubrico pedes tuos et recesserunt a te
JER|38|23|et omnes uxores tuae et filii tui educentur ad Chaldeos et non effugies manus eorum sed in manu regis Babylonis capieris et civitatem hanc conburet igni
JER|38|24|dixit ergo Sedecias ad Hieremiam nullus sciat verba haec et non morieris
JER|38|25|si autem audierint principes quia locutus sum tecum et venerint ad te et dixerint tibi indica nobis quid locutus sis cum rege ne celes nos et non te interficiemus et quid locutus est tecum rex
JER|38|26|dices ad eos prostravi ego preces meas coram rege ne me reduci iuberet in domum Ionathan et ibi morerer
JER|38|27|venerunt ergo omnes principes ad Hieremiam et interrogaverunt eum et locutus est eis iuxta omnia verba quae praeceperat ei rex et cessaverunt ab eo nihil enim fuerat auditum
JER|38|28|mansit vero Hieremias in vestibulo carceris usque ad diem quo capta est Hierusalem et factum est ut caperetur Hierusalem
JER|39|1|anno nono Sedeciae regis Iuda mense decimo venit Nabuchodonosor rex Babylonis et omnis exercitus eius ad Hierusalem et obsidebant eam
JER|39|2|undecimo autem anno Sedeciae mense quarto quinta mensis aperta est civitas
JER|39|3|et ingressi sunt omnes principes regis Babylonis et sederunt in porta media Neregel Sereser Semegar Nabu Sarsachim Rabsares Neregel Sereser Rebmag et omnes reliqui principes regis Babylonis
JER|39|4|cumque vidisset eos Sedecias rex Iuda et omnes viri bellatores fugerunt et egressi sunt nocte de civitate per viam horti regis et per portam quae erat inter duos muros et egressi sunt ad viam deserti
JER|39|5|persecutus est autem eos exercitus Chaldeorum et conprehenderunt Sedeciam in campo solitudinis hiericuntinae et captum adduxerunt ad Nabuchodonosor regem Babylonis in Reblatha quae est in terra Emath et locutus est ad eum iudicia
JER|39|6|et occidit rex Babylonis filios Sedeciae in Reblatha in oculis eius et omnes nobiles Iuda occidit rex Babylonis
JER|39|7|oculos quoque Sedeciae eruit et vinxit eum conpedibus ut duceretur in Babylonem
JER|39|8|domum quoque regis et domum vulgi succenderunt Chaldei igni et murum Hierusalem subverterunt
JER|39|9|et reliquias populi quae remanserunt in civitate et perfugas qui transfugerant ad eum et superfluos vulgi qui remanserant transtulit Nabuzardan magister militum in Babylonem
JER|39|10|et de plebe pauperum qui nihil penitus habebant dimisit Nabuzardan magister militum in terra Iuda et dedit eis vineas et cisternas in die illa
JER|39|11|praeceperat autem Nabuchodonosor rex Babylonis de Hieremia Nabuzardan magistro militiae dicens
JER|39|12|tolle illum et pone super eum oculos tuos nihilque ei mali facias sed ut voluerit sic facies ei
JER|39|13|misit ergo Nabuzardan princeps militiae et Nabu et Sesban et Rabsares et Neregel et Sereser et Rebmag et omnes optimates regis Babylonis
JER|39|14|miserunt et tulerunt Hieremiam de vestibulo carceris et tradiderunt eum Godoliae filio Ahicam filii Saphan ut intraret domum et habitaret in populo
JER|39|15|ad Hieremiam autem factus fuerat sermo Domini cum clausus esset in vestibulo carceris dicens
JER|39|16|vade et dic Abdemelech Aethiopi dicens haec dicit Dominus exercituum Deus Israhel ecce ego inducam sermones meos super civitatem hanc in malum et non in bonum et erunt in conspectu tuo in die illa
JER|39|17|et liberabo te in die illa ait Dominus et non traderis in manus virorum quos tu formidas
JER|39|18|sed eruens liberabo te et gladio non cades sed erit tibi anima tua in salutem quia in me habuisti fiduciam ait Dominus
JER|40|1|sermo qui factus est ad Hieremiam a Domino postquam dimissus est a Nabuzardan magistro militiae de Rama quando tulit eum vinctum catenis in medio omnium qui migrabant de Hierusalem et Iuda et ducebantur in Babylonem
JER|40|2|tollens ergo princeps militiae Hieremiam dixit ad eum Dominus Deus tuus locutus est malum hoc super locum istum
JER|40|3|et adduxit et fecit Dominus sicut locutus est quia peccastis Domino et non audistis vocem eius et factus est vobis sermo hic
JER|40|4|nunc ergo ecce solvi te hodie de catenis quae sunt in manibus tuis si placet tibi ut venias mecum in Babylonem veni et ponam oculos meos super te si autem displicet tibi venire mecum in Babylonem reside ecce omnis terra in conspectu tuo quod elegeris et quo placuerit tibi ut vadas illuc perge
JER|40|5|et mecum noli venire sed habita apud Godoliam filium Ahicam filii Saphan quem praeposuit rex Babylonis civitatibus Iudaeae habita ergo cum eo in medio populi vel quocumque placuerit tibi ut vadas vade dedit quoque ei magister militiae cibaria et munuscula et dimisit eum
JER|40|6|venit autem Hieremias ad Godoliam filium Ahicam in Masphat et habitavit cum eo in medio populi qui relictus fuerat in terra
JER|40|7|cum ergo audissent omnes principes exercitus qui dispersi fuerant per regiones ipsi et socii eorum quod praefecisset rex Babylonis Godoliam filium Ahicam terrae et quod commendasset ei viros et mulieres et parvulos et de pauperibus terrae qui non fuerant translati in Babylonem
JER|40|8|venerunt ad Godoliam in Masphat et Ismahel filius Nathaniae et Iohanan et Ionathan filii Caree et Sareas filius Thenoemeth et filii Offi qui erat de Nethophathi et Iezonias filius Maachathi ipsi et viri eorum
JER|40|9|et iuravit eis Godolias filius Ahicam filii Saphan et comitibus eorum dicens nolite timere servire Chaldeis habitate in terra et servite regi Babylonis et bene erit vobis
JER|40|10|ecce ego habito in Masphat ut respondeam praecepto Chaldeorum qui mittuntur ad nos vos autem colligite vindemiam et messem et oleum et condite in vasis vestris et manete in urbibus vestris quas tenetis
JER|40|11|sed et omnes Iudaei qui erant in Moab et in filiis Ammon et in Idumea et in universis regionibus audito quod dedisset rex Babylonis reliquias in Iudaeam et quod praeposuisset super eos Godoliam filium Ahicam filii Saphan
JER|40|12|reversi sunt inquam omnes Iudaei de universis locis ad quae profugerant et venerunt in terram Iuda ad Godoliam in Masphat et collegerunt vinum et messem multam nimis
JER|40|13|Iohanan autem filius Caree et omnes principes exercitus qui dispersi erant in regionibus venerunt ad Godoliam in Masphat
JER|40|14|et dixerunt ei scito quia Baalis rex filiorum Ammon misit Ismahel filium Nathaniae percutere animam tuam et non credidit eis Godolias filius Ahicam
JER|40|15|Iohanan vero filius Caree dixit ad Godoliam seorsum in Masphat loquens ibo et percutiam Ismahel filium Nathaniae nullo sciente ne interficiat animam tuam et dissipentur omnes Iudaei qui congregati sunt ad te et peribunt reliquiae Iuda
JER|40|16|et ait Godolias filius Ahicam ad Iohanan filium Caree noli facere verbum hoc falsum enim tu loqueris de Ismahel
JER|41|1|et factum est in mense septimo venit Ismahel filius Nathaniae filii Elisama de semine regali et optimates regis et decem viri cum eo ad Godoliam filium Ahicam in Masphat et comederunt ibi panes simul in Masphat
JER|41|2|surrexit autem Ismahel filius Nathaniae et decem viri qui erant cum eo et percusserunt Godoliam filium Ahicam filii Saphan gladio et interfecerunt eum quem praefecerat rex Babylonis terrae
JER|41|3|omnes quoque Iudaeos qui erant cum Godolia in Masphat et Chaldeos qui repperti sunt ibi et viros bellatores percussit Ismahel
JER|41|4|secundo autem die postquam occiderat Godoliam nullo adhuc sciente
JER|41|5|venerunt viri de Sychem et de Silo et de Samaria octoginta viri rasi barbam et scissis vestibus et squalentes munera et tus habebant in manu ut offerrent in domo Domini
JER|41|6|egressus ergo Ismahel filius Nathaniae in occursum eorum de Masphat incedens et plorans ibat cum autem occurrisset eis dixit ad eos venite ad Godoliam filium Ahicam
JER|41|7|qui cum venissent ad medium civitatis interfecit eos Ismahel filius Nathaniae circa medium laci ipse et viri qui erant cum eo
JER|41|8|decem autem viri repperti sunt inter eos qui dixerunt ad Ismahel noli occidere nos quia habemus thesauros in agro frumenti et hordei et olei et mellis et cessavit et non interfecit eos cum fratribus suis
JER|41|9|lacus autem in quem proiecerat Ismahel omnia cadavera virorum quos percussit propter Godoliam ipse est quem fecit rex Asa propter Baasa regem Israhel ipsum replevit Ismahel filius Nathaniae occisis
JER|41|10|et captivas duxit Ismahel omnes reliquias populi qui erant in Masphat filias regis et universum populum qui remanserat in Masphat quos commendarat Nabuzardan princeps militiae Godoliae filio Ahicam et cepit eos Ismahel filius Nathaniae et abiit ut transiret ad filios Ammon
JER|41|11|audivit autem Iohanan filius Caree et omnes principes bellatorum qui erant cum eo omne malum quod fecerat Ismahel filius Nathaniae
JER|41|12|et adsumptis universis viris profecti sunt ut bellarent adversum Ismahel filium Nathaniae et invenerunt eum ad aquas Multas quae sunt in Gabaon
JER|41|13|cumque vidisset omnis populus qui erat cum Ismahel Iohanan filium Caree et universos principes bellatorum qui erant cum eo laetati sunt
JER|41|14|et reversus est omnis populus quem ceperat Ismahel in Masphat reversusque abiit ad Iohanan filium Caree
JER|41|15|Ismahel autem filius Nathaniae fugit cum octo viris a facie Iohanan et abiit ad filios Ammon
JER|41|16|tulit ergo Iohanan filius Caree et omnes principes bellatorum qui erant cum eo universas reliquias vulgi quas reduxerat ab Ismahel filio Nathaniae de Masphat postquam percussit Godoliam filium Ahicam fortes viros ad proelium et mulieres et pueros et eunuchos quos reduxerat de Gabaon
JER|41|17|et abierunt et sederunt peregrinantes in Chamaam quae est iuxta Bethleem ut pergerent et introirent Aegyptum
JER|41|18|a facie Chaldeorum timebant enim eos quia percusserat Ismahel filius Nathaniae Godoliam filium Ahicam quem praeposuerat rex Babylonis in terra Iuda
JER|42|1|et accesserunt omnes principes bellatorum et Iohanan filius Caree et Iezonias filius Osaiae et reliquum vulgus a parvo usque ad magnum
JER|42|2|dixeruntque ad Hieremiam prophetam cadat oratio nostra in conspectu tuo et ora pro nobis ad Dominum Deum tuum pro universis reliquiis istis quia derelicti sumus pauci de pluribus sicut oculi tui nos intuentur
JER|42|3|et adnuntiet nobis Dominus Deus tuus viam per quam pergamus et verbum quod faciamus
JER|42|4|dixit autem ad eos Hieremias propheta audivi ecce ego oro ad Dominum Deum vestrum secundum verba vestra omne verbum quodcumque responderit mihi indicabo vobis nec celabo vos quicquam
JER|42|5|et illi dixerunt ad Hieremiam sit Dominus inter nos testis veritatis et fidei si non iuxta omne verbum in quo miserit te Dominus Deus tuus ad nos sic faciemus
JER|42|6|sive bonum est sive malum voci Domini Dei nostri ad quem mittimus te oboediemus ut bene sit nobis cum audierimus vocem Domini Dei nostri
JER|42|7|cum autem conpleti essent decem dies factum est verbum Domini ad Hieremiam
JER|42|8|vocavitque Iohanan filium Caree et omnes principes bellatorum qui erant cum eo et universum populum a minimo usque ad magnum
JER|42|9|et dixit ad eos haec dicit Dominus Deus Israhel ad quem misistis me ut prosternerem preces vestras in conspectu eius
JER|42|10|si quiescentes manseritis in terra hac aedificabo vos et non destruam plantabo et non evellam iam enim placatus sum super malo quod feci vobis
JER|42|11|nolite timere a facie regis Babylonis quem vos pavidi formidatis nolite eum metuere dicit Dominus quia vobiscum sum ego ut salvos faciam vos et eruam de manu eius
JER|42|12|et dabo vobis misericordiam et miserebor vestri et habitare vos faciam in terra vestra
JER|42|13|si autem dixeritis vos non habitabimus in terra ista nec audiemus vocem Domini Dei nostri
JER|42|14|dicentes nequaquam sed ad terram Aegypti pergemus ubi non videbimus bellum et clangorem tubae non audiemus et famem non sustinebimus et ibi habitabimus
JER|42|15|propter hoc nunc audite verbum Domini reliquiae Iuda haec dicit Dominus exercituum Deus Israhel si posueritis faciem vestram ut ingrediamini Aegyptum et intraveritis ut ibi habitetis
JER|42|16|gladium quem vos formidatis ibi conprehendet vos in terra Aegypti et fames pro qua estis solliciti adherebit vobis in Aegypto et ibi moriemini
JER|42|17|omnesque viri qui posuerint faciem suam ut ingrediantur Aegyptum et habitent ibi morientur gladio et fame et peste nullus de eis remanebit nec effugient a facie mali quod ego adferam super eos
JER|42|18|quia haec dicit Dominus exercituum Deus Israhel sicut conflatus est furor meus et indignatio mea super habitatores Hierusalem sic conflabitur indignatio mea super vos cum ingressi fueritis Aegyptum et eritis in iusiurandum et in stuporem et in maledictum et in obprobrium et nequaquam ultra videbitis locum istum
JER|42|19|verbum Domini super vos reliquiae Iuda nolite intrare Aegyptum scientes scietis quia obtestatus sum vobis hodie
JER|42|20|quia decepistis animas vestras vos enim misistis me ad Dominum Deum nostrum dicentes ora pro nobis ad Dominum Deum nostrum et iuxta omnia quaecumque dixerit tibi Dominus Deus noster sic adnuntia nobis et faciemus
JER|42|21|et adnuntiavi vobis hodie et non audistis vocem Domini Dei vestri super universis pro quibus misit me ad vos
JER|42|22|nunc ergo scientes scietis quia gladio et fame et peste moriemini in loco ad quem voluistis intrare ut habitaretis ibi
JER|43|1|factum est autem cum conplesset Hieremias loquens ad populum universos sermones Domini Dei eorum pro quibus miserat eum Dominus Deus eorum ad illos omnia verba haec
JER|43|2|dixit Azarias filius Osaiae et Iohanan filius Caree et omnes viri superbi dicentes ad Hieremiam mendacium tu loqueris non misit te Dominus Deus noster dicens ne ingrediamini Aegyptum ut habitetis illuc
JER|43|3|sed Baruch filius Neriae incitat te adversum nos ut tradat nos in manibus Chaldeorum ut interficiat nos et transduci faciat in Babylonem
JER|43|4|et non audivit Iohanan filius Caree et omnes principes bellatorum et universus populus vocem Domini ut maneret in terra Iuda
JER|43|5|sed tollens Iohanan filius Caree et universi principes bellatorum universos reliquiarum Iuda qui reversi fuerant de cunctis gentibus ad quas fuerant ante dispersi ut habitarent in terra Iuda
JER|43|6|viros et mulieres et parvulos et filias regis et omnem animam quam reliquerat Nabuzardan princeps militiae cum Godolia filio Ahicam filii Saphan et Hieremiam prophetam et Baruch filium Neriae
JER|43|7|et ingressi sunt terram Aegypti quia non oboedierunt voci Domini et venerunt usque ad Tafnas
JER|43|8|et factus est sermo Domini ad Hieremiam in Tafnis dicens
JER|43|9|sume in manu tua lapides grandes et absconde eos in crypta quae est sub muro latericio in porta domus Pharaonis in Tafnis cernentibus viris iudaeis
JER|43|10|et dices ad eos haec dicit Dominus exercituum Deus Israhel ecce ego mittam et adsumam Nabuchodonosor regem Babylonis servum meum et ponam thronum eius super lapides istos quos abscondi et statuet solium suum super eos
JER|43|11|veniensque percutiet terram Aegypti quos in morte in morte et quos in captivitate in captivitate et quos in gladio in gladio
JER|43|12|et succendet ignem in delubris deorum Aegypti et conburet ea et captivos ducet illos et amicietur terra Aegypti sicut amicitur pastor pallio suo et egredietur inde in pace
JER|43|13|et conteret statuas domus Solis quae sunt in terra Aegypti et delubra deorum Aegypti conburet igni
JER|44|1|verbum quod factum est ad Hieremiam ad omnes Iudaeos qui habitant in terra Aegypti habitantes in Magdolo et in Tafnis et in Memphis et in terra Fatures dicens
JER|44|2|haec dicit Dominus exercituum Deus Israhel vos vidistis omne malum istud quod adduxi super Hierusalem et super omnes urbes Iuda et ecce sunt desertae hodie et non est in eis habitator
JER|44|3|propter malitiam quam fecerunt ut me ad iracundiam provocarent et irent et sacrificarent et colerent deos alienos quos nesciebant et illi et vos et patres vestri
JER|44|4|et misi ad vos omnes servos meos prophetas de nocte consurgens mittensque et dicens nolite facere verbum abominationis huius quam odi
JER|44|5|et non audierunt nec inclinaverunt aurem suam ut converterentur a malis suis et non sacrificarent diis alienis
JER|44|6|et conflata est indignatio mea et furor meus et succensa est in civitatibus Iuda et in plateis Hierusalem et versae sunt in solitudinem et vastitatem secundum diem hanc
JER|44|7|et nunc haec dicit Dominus exercituum Deus Israhel quare vos facitis malum grande contra animas vestras ut intereat ex vobis vir et mulier parvulus et lactans de medio Iudae nec relinquatur vobis quicquam residuum
JER|44|8|provocantes me in operibus manuum vestrarum sacrificando diis alienis in terra Aegypti in quam ingressi estis ut habitetis ibi et dispereatis et sitis in maledictionem et in obprobrium cunctis gentibus terrae
JER|44|9|numquid obliti estis mala patrum vestrorum et mala regum Iuda et mala uxorum eius et mala vestra et mala uxorum vestrarum quae fecerunt in terra Iuda et in regionibus Hierusalem
JER|44|10|non sunt mundati usque ad diem hanc et non timuerunt et non ambulaverunt in lege et in praeceptis meis quae dedi coram vobis et coram patribus vestris
JER|44|11|ideo haec dicit Dominus exercituum Deus Israhel ecce ego pono faciem meam in vobis in malum et disperdam omnem Iudam
JER|44|12|et adsumam reliquias Iudae qui posuerunt facies suas ut ingrederentur terram Aegypti et habitarent ibi et consumentur omnes in terra Aegypti cadent in gladio et in fame consumentur a minimo usque ad maximum in gladio et in fame morientur et erunt in iusiurandum et in miraculum et in maledictionem et in obprobrium
JER|44|13|et visitabo habitatores terrae Aegypti sicut visitavi super Hierusalem in gladio et in fame et in peste
JER|44|14|et non erit qui effugiat et sit residuus de reliquiis Iudaeorum qui vadunt ut peregrinentur in terra Aegypti et revertantur in terram Iuda ad quam ipsi elevant animas suas ut revertantur et habitent ibi non revertentur nisi qui fugerint
JER|44|15|responderunt autem Hieremiae omnes viri scientes quod sacrificarent uxores eorum diis alienis et universae mulieres quarum stabat multitudo grandis et omnis populus habitantium in terra Aegypti in Fatures dicens
JER|44|16|sermonem quem locutus es ad nos in nomine Domini non audiemus ex te
JER|44|17|sed facientes faciemus omne verbum quod egreditur de ore nostro ut sacrificemus Reginae caeli et libemus ei libamina sicut fecimus nos et patres nostri reges nostri et principes nostri in urbibus Iuda et in plateis Hierusalem et saturati sumus panibus et bene nobis erat malumque non vidimus
JER|44|18|ex eo autem quo cessavimus sacrificare Reginae caeli et libare ei libamina indigemus omnibus et gladio et fame consumpti sumus
JER|44|19|quod si nos sacrificamus Reginae caeli et libamus ei libamina numquid sine viris nostris fecimus ei placentas ad colendum eam et liba libandi
JER|44|20|et dixit Hieremias ad omnem populum adversum viros et adversum mulieres et adversum universam plebem qui responderant ei verbum dicens
JER|44|21|numquid non sacrificium quod sacrificastis in civitatibus Iuda et in plateis Hierusalem vos et patres vestri reges vestri et principes vestri et populus terrae horum recordatus est Dominus et ascendit super cor eius
JER|44|22|et non poterat Dominus ultra portare propter malitiam studiorum vestrorum et propter abominationes quas fecistis et facta est terra vestra in desolationem et in stuporem et in maledictum eo quod non sit habitator sicut est dies haec
JER|44|23|propterea quod sacrificaveritis idolis et peccaveritis Domino et non audieritis vocem Domini et in lege et in praeceptis et in testimoniis eius non ambulaveritis idcirco evenerunt vobis mala haec sicut est dies haec
JER|44|24|dixit autem Hieremias ad omnem populum et ad universas mulieres audite verbum Domini omnis Iuda qui estis in terra Aegypti
JER|44|25|haec inquit Dominus exercituum Deus Israhel dicens vos et uxores vestrae locuti estis ore vestro et manibus vestris implestis dicentes faciamus vota nostra quae vovimus ut sacrificemus Reginae caeli et libemus ei libamina implestis vota vestra et opere perpetrastis ea
JER|44|26|ideo audite verbum Domini omnis Iuda qui habitatis in terra Aegypti ecce ego iuravi in nomine meo magno ait Dominus quia nequaquam ultra nomen meum vocabitur ex ore omnis viri iudaei dicentis vivit Dominus Deus in omni terra Aegypti
JER|44|27|ecce ego vigilabo super eos in malum et non in bonum et consumentur omnes viri Iuda qui sunt in terra Aegypti gladio et fame donec penitus consumantur
JER|44|28|et qui fugerint gladium revertentur de terra Aegypti in terram Iuda viri pauci et scient omnes reliquiae Iuda ingredientium terram Aegypti ut habitent ibi cuius sermo conpleatur meus an illorum
JER|44|29|et hoc vobis signum ait Dominus quod visitem ego super vos in loco isto ut sciatis quia vere conplebuntur sermones mei contra vos in malum
JER|44|30|haec dicit Dominus ecce ego tradam Pharaonem Efree regem Aegypti in manu inimicorum eius et in manu quaerentium animam illius sicut tradidi Sedeciam regem Iuda in manu Nabuchodonosor regis Babylonis inimici sui et quaerentis animam eius
JER|45|1|verbum quod locutus est Hieremias propheta ad Baruch filium Neri cum scripsisset verba haec in libro de ore Hieremiae anno quarto Ioachim filii Iosiae regis Iuda dicens
JER|45|2|haec dicit Dominus Deus Israhel ad te Baruch
JER|45|3|dixisti vae misero mihi quoniam addidit Dominus dolorem dolori meo laboravi in gemitu meo et requiem non inveni
JER|45|4|haec dices ad eum sic dicit Dominus ecce quos aedificavi ego destruo et quos plantavi ego evello et universam terram hanc
JER|45|5|et tu quaeris tibi grandia noli quaerere quia ecce ego adducam malum super omnem carnem ait Dominus et dabo tibi animam tuam in salutem in omnibus locis ad quaecumque perrexeris
JER|46|1|quod factum est verbum Domini ad Hieremiam prophetam contra gentes
JER|46|2|ad Aegyptum adversum exercitum Pharaonis Nechao regis Aegypti qui erat iuxta flumen Eufraten in Charchamis quem percussit Nabuchodonosor rex Babylonis in quarto anno Ioachim filii Iosiae regis Iuda
JER|46|3|praeparate scutum et clypeum et procedite ad bellum
JER|46|4|iungite equos et ascendite equites state in galeis polite lanceas induite vos loricis
JER|46|5|quid igitur vidi ipsos pavidos et terga vertentes fortes eorum caesos fugerunt conciti nec respexerunt terror undique ait Dominus
JER|46|6|non fugiat velox nec salvari se putet fortis ad aquilonem iuxta flumen Eufraten victi sunt et ruerunt
JER|46|7|quis est iste qui quasi flumen ascendit et veluti fluviorum intumescunt gurgites eius
JER|46|8|Aegyptus fluminis instar ascendet et velut flumina movebuntur fluctus eius et dicet ascendens operiam terram perdam civitatem et habitatores eius
JER|46|9|ascendite equos et exultate in curribus et procedant fortes Aethiopia et Lybies tenentes scutum et Lydii arripientes et iacientes sagittas
JER|46|10|dies autem ille Domini Dei exercituum dies ultionis ut sumat vindictam de inimicis suis devorabit gladius et saturabitur et inebriabitur sanguine eorum victima enim Domini exercituum in terra aquilonis iuxta flumen Eufraten
JER|46|11|ascende in Galaad et tolle resinam virgo filia Aegypti frustra multiplicas medicamina sanitas non erit tibi
JER|46|12|audierunt gentes ignominiam tuam et ululatus tuus replevit terram quia fortis inpegit in fortem ambo pariter conciderunt
JER|46|13|verbum quod locutus est Dominus ad Hieremiam prophetam super eo quod venturus esset Nabuchodonosor rex Babylonis et percussurus terram Aegypti
JER|46|14|adnuntiate Aegypto et auditum facite Magdolo et resonet in Memphis et in Tafnis dicite sta et praepara te quia devoravit gladius ea quae per circuitum tuum sunt
JER|46|15|quare conputruit fortis tuus non stetit quoniam Dominus subvertit eum
JER|46|16|multiplicavit ruentes ceciditque vir ad proximum suum et dicent surge et revertamur ad populum nostrum et ad terram nativitatis nostrae a facie gladii columbae
JER|46|17|vocate nomen Pharao regis Aegypti Tumultum adduxit tempus
JER|46|18|vivo ego inquit Rex Dominus exercituum nomen eius quoniam sicut Thabor in montibus et sicut Carmelus in mari veniet
JER|46|19|vasa transmigrationis fac tibi habitatrix filia Aegypti quia Memphis in solitudinem erit et deseretur inhabitabilis
JER|46|20|vitula eligans atque formonsa Aegyptus stimulator ab aquilone veniet ei
JER|46|21|mercennarii quoque eius qui versabantur in medio eius quasi vituli saginati versi sunt et fugerunt simul nec stare potuerunt quia dies interfectionis eorum venit super eos tempus visitationis eorum
JER|46|22|vox eius quasi aeris sonabit quoniam cum exercitu properabunt et cum securibus venient ei quasi ligna caedentes
JER|46|23|succiderunt saltum eius ait Dominus qui supputari non potest multiplicati sunt super lucustas et non est eis numerus
JER|46|24|confusa est filia Aegypti et tradita in manu populi aquilonis
JER|46|25|dixit Dominus exercituum Deus Israhel ecce ego visitabo super tumultum Alexandriae et super Pharao et super Aegyptum et super deos eius et super reges eius et super Pharao et super eos qui confidunt in eo
JER|46|26|et dabo eos in manu quaerentium animam eorum et in manu Nabuchodonosor regis Babylonis et in manu servorum eius et post haec habitabitur sicut diebus pristinis ait Dominus
JER|46|27|et tu ne timeas serve meus Iacob et ne paveas Israhel quia ecce ego salvum te faciam de longinquo et semen tuum de terra captivitatis suae et revertetur Iacob et quiescet et prosperabitur et non erit qui exterreat eum
JER|46|28|et tu noli timere serve meus Iacob ait Dominus quia tecum ego sum quia consumam ego cunctas gentes ad quas eieci te te vero non consumam sed castigabo te in iudicio nec quasi innocenti parcam tibi
JER|47|1|quod factum est verbum Domini ad Hieremiam prophetam contra Palestinos antequam percuteret Pharao Gazam
JER|47|2|haec dicit Dominus ecce aquae ascendunt ab aquilone et erunt quasi torrens inundans et operient terram et plenitudinem eius urbem et habitatores eius clamabunt homines et ululabit omnis habitator terrae
JER|47|3|ab strepitu pompae armorum et bellatorum eius a commotione quadrigarum eius et multitudine rotarum illius non respexerunt patres filios manibus dissolutis
JER|47|4|pro adventu diei in quo vastabuntur omnes Philisthim et dissipabitur Tyrus et Sidon cum omnibus reliquis auxiliis suis depopulatus est enim Dominus Palestinos reliquias insulae Cappadociae
JER|47|5|venit calvitium super Gazam conticuit Ascalon et reliquiae vallis earum usquequo concideris
JER|47|6|o mucro Domini usquequo non quiescis ingredere in vaginam tuam refrigerare et sile
JER|47|7|quomodo quiescet cum Dominus praeceperit ei adversus Ascalonem et adversus maritimas eius regiones ibique condixerit illi
JER|48|1|ad Moab haec dicit Dominus exercituum Deus Israhel vae super Nabo quoniam vastata est et confusa capta est Cariathaim confusa est fortis et tremuit
JER|48|2|non est ultra exultatio in Moab contra Esebon cogitaverunt malum venite et disperdamus eam de gente ergo silens conticesces sequeturque te gladius
JER|48|3|vox clamoris de Oronaim vastitas et contritio magna
JER|48|4|contrita est Moab adnuntiate clamorem parvulis eius
JER|48|5|per ascensum enim Luaith plorans ascendet in fletu quoniam in descensu Oronaim hostes ululatum contritionis audierunt
JER|48|6|fugite salvate animas vestras et eritis quasi myrice in deserto
JER|48|7|pro eo enim quod habuisti fiduciam in munitionibus tuis et in thesauris tuis tu quoque capieris et ibit Chamos in transmigrationem sacerdotes eius et principes eius simul
JER|48|8|et veniet praedo ad omnem urbem et urbs nulla salvabitur et peribit vallis et dissipabuntur campestria quoniam dixit Dominus
JER|48|9|date florem Moab quia floriens egredietur et civitates eius desertae erunt et inhabitabiles
JER|48|10|maledictus qui facit opus Domini fraudulenter et maledictus qui prohibet gladium suum a sanguine
JER|48|11|fertilis fuit Moab ab adulescentia sua et requievit in fecibus suis nec transfusus est de vase in vas et in transmigrationem non abiit idcirco permansit gustus eius in eo et odor eius non est inmutatus
JER|48|12|propterea ecce dies veniunt dicit Dominus et mittam ei ordinatores et stratores laguncularum et sternent eum et vasa eius exhaurient et lagoenas eorum conlident
JER|48|13|et confundetur Moab a Chamos sicut confusa est domus Israhel a Bethel in qua habebat fiduciam
JER|48|14|quomodo dicitis fortes sumus et viri robusti ad proeliandum
JER|48|15|vastata est Moab et civitates illius ascenderunt et electi iuvenes eius descenderunt in occisionem ait Rex Dominus exercituum nomen ei
JER|48|16|prope est interitus Moab ut veniat et malum eius velociter adcurret nimis
JER|48|17|consolamini eum omnes qui estis in circuitu eius et universi qui scitis nomen eius dicite quomodo confracta est virga fortis baculus gloriosus
JER|48|18|descende de gloria et sede in siti habitatio filiae Dibon quoniam vastator Moab ascendet ad te dissipabit munitiones tuas
JER|48|19|in via sta et prospice habitatio Aroer interroga fugientem et eum qui evasit dic quid accidit
JER|48|20|confusus est Moab quoniam victus est ululate et clamate adnuntiate in Arnon quoniam vastata est Moab
JER|48|21|et iudicium venit ad terram campestrem super Helon et super Iaesa et super Mefath
JER|48|22|et super Dibon et super Nabo et super domum Deblathaim
JER|48|23|et super Cariathaim et super Bethgamul et super Bethmaon
JER|48|24|et super Carioth et super Bosra et super omnes civitates terrae Moab quae longe et quae prope sunt
JER|48|25|abscisum est cornu Moab et brachium eius contritum est ait Dominus
JER|48|26|inebriate eum quoniam contra Dominum erectus est et adlidet manum Moab in vomitu suo et erit in derisum etiam ipse
JER|48|27|fuit enim in derisum tibi Israhel quasi inter fures repperisses eum propter verba ergo tua quae adversum illum locutus es captivus duceris
JER|48|28|relinquite civitates et habitate in petra habitatores Moab et estote quasi columba nidificans in summo ore foraminis
JER|48|29|audivimus superbiam Moab superbus est valde sublimitatem eius et arrogantiam et superbiam et altitudinem cordis illius
JER|48|30|ego scio ait Dominus iactantiam eius et quod non sit iuxta eam virtus eius nec iuxta quod poterat conata sit facere
JER|48|31|ideo super Moab heiulabo et ad Moab universam clamabo ad viros muri fictilis lamentantes
JER|48|32|de planctu Iazer plorabo tibi vinea Sobema propagines tuae transierunt mare usque ad mare Iazer pervenerunt super messem tuam et vindemiam tuam praedo inruit
JER|48|33|ablata est laetitia et exultatio de Carmelo et de terra Moab et vinum de torcularibus sustuli nequaquam calcator uvae solitum celeuma cantabit
JER|48|34|de clamore Esebon usque Eleale et Iaesa dederunt vocem suam a Segor usque ad Oronaim vitula conternante aquae quoque Namrim pessimae erunt
JER|48|35|et auferam de Moab ait Dominus offerentem in excelsis et sacrificantem diis eius
JER|48|36|propterea cor meum ad Moab quasi tibiae resonabit et cor meum ad viros muri fictilis dabit sonitum tibiarum quia plus fecit quam potuit idcirco perierunt
JER|48|37|omne enim caput calvitium et omnis barba rasa erit in cunctis manibus conligatio et super omne dorsum cilicium
JER|48|38|super omnia tecta Moab et in plateis eius omnis planctus quia contrivi Moab sicut vas inutile ait Dominus
JER|48|39|quomodo victa est et ululaverunt quomodo deiecit cervicem Moab et confusus est eritque Moab in derisum et in exemplum omnibus in circuitu suo
JER|48|40|haec dicit Dominus ecce quasi aquila evolabit et extendet alas suas ad Moab
JER|48|41|capta est Carioth et munitiones conprehensae sunt et erit cor fortium Moab in die illa sicut cor mulieris parturientis
JER|48|42|et cessabit Moab esse populus quoniam contra Dominum gloriatus est
JER|48|43|pavor et fovea et laqueus super te o habitator Moab ait Dominus
JER|48|44|qui fugit a facie pavoris cadet in foveam et qui conscenderit de fovea capietur laqueo adducam enim super Moab annum visitationis eorum dicit Dominus
JER|48|45|in umbra Esebon steterunt de laqueo fugientes quia ignis egressus est de Esebon et flamma de medio Seon et devorabit partem Moab et verticem filiorum tumultus
JER|48|46|vae tibi Moab peristi popule Chamos quia conprehensi sunt filii tui et filiae tuae in captivitatem
JER|48|47|et convertam captivitatem Moab in novissimis diebus ait Dominus hucusque iudicia Moab
JER|49|1|ad filios Ammon haec dicit Dominus numquid filii non sunt Israhel aut heres non est ei cur igitur hereditate possedit Melchom Gad et populus eius in urbibus eius habitavit
JER|49|2|ideo ecce dies veniunt dicit Dominus et auditum faciam super Rabbath filiorum Ammon fremitum proelii et erit in tumulum dissipata filiaeque eius igni succendentur et possidebit Israhel possessores suos dicit Dominus
JER|49|3|ulula Esebon quoniam vastata est Ahi clamate filiae Rabbath accingite vos ciliciis plangite et circuite per sepes quia Melchom in transmigratione ducetur sacerdotes eius et principes eius simul
JER|49|4|quid gloriaris in vallibus defluxit vallis tua filia delicata quae confidebas in thesauris tuis et dicebas quis veniet ad me
JER|49|5|ecce ego inducam super te terrorem ait Dominus Deus exercituum ab omnibus qui sunt in circuitu tuo et dispergemini singuli a conspectu vestro nec erit qui congreget fugientem
JER|49|6|et post haec reverti faciam captivos filiorum Ammon ait Dominus
JER|49|7|ad Idumeam haec dicit Dominus exercituum numquid non est ultra sapientia in Theman periit consilium a filiis inutilis facta est sapientia eorum
JER|49|8|fugite terga vertite descendite in voragine habitatores Dedan quoniam perditionem Esau adduxi super eum tempus visitationis eius
JER|49|9|si vindemiatores venissent super te non reliquissent racemum si fures in nocte rapuissent quod sufficeret sibi
JER|49|10|ego vero discoperui Esau revelavi abscondita eius et celari non poterit vastatum est semen eius et fratres eius et vicini eius et non erit
JER|49|11|relinque pupillos tuos ego eos faciam vivere et viduae tuae in me sperabunt
JER|49|12|quia haec dicit Dominus ecce quibus non erat iudicium ut biberent calicem bibentes bibent et tu quasi innocens relinqueris non eris innocens sed bibens bibes
JER|49|13|quia per memet ipsum iuravi dicit Dominus quod in solitudinem et in obprobrium et in desertum et in maledictionem erit Bosra et omnes civitates eius erunt in solitudines sempiternas
JER|49|14|auditum audivi a Domino et legatus ad gentes missus est congregamini et venite contra eam et consurgamus in proelium
JER|49|15|ecce enim parvulum dedi te in gentibus contemptibilem inter homines
JER|49|16|arrogantia tua decepit te et superbia cordis tui qui habitas in cavernis petrae et adprehendere niteris altitudinem collis cum exaltaveris quasi aquila nidum tuum inde detraham te dicit Dominus
JER|49|17|et erit Idumea deserta omnis qui transibit per eam stupebit et sibilabit super omnes plagas eius
JER|49|18|sicuti subversa est Sodoma et Gomorra et vicinae eius ait Dominus non habitabit ibi vir et non incolet eam filius hominis
JER|49|19|ecce quasi leo ascendet de superbia Iordanis ad pulchritudinem robustam quia subito currere eum faciam ad illam et quis erit electus quem praeponam ei quis enim similis mei et quis sustinebit me et quis est iste pastor qui resistat vultui meo
JER|49|20|propterea audite consilium Domini quod iniit de Edom et cogitationes eius quas cogitavit de habitatoribus Theman si non deiecerint eos parvuli gregis nisi dissipaverint cum eis habitaculum eorum
JER|49|21|a voce ruinae eorum commota est terra clamor in mari Rubro auditus est vocis eius
JER|49|22|ecce quasi aquila ascendet et evolabit et expandet alas suas super Bosram et erit cor fortium Idumeae in die illa quasi cor mulieris parturientis
JER|49|23|ad Damascum confusa est Emath et Arfad quia auditum pessimum audierunt turbati sunt in mari sollicitudine quiescere non potuit
JER|49|24|dissoluta est Damascus versa in fugam tremor adprehendit eam angustia et dolores tenuerunt eam quasi parturientem
JER|49|25|quomodo dereliquerunt civitatem laudabilem urbem laetitiae
JER|49|26|ideo cadent iuvenes eius in plateis eius et omnes viri proelii conticescent in die illa ait Dominus exercituum
JER|49|27|et succendam ignem in muro Damasci et devorabit moenia Benadad
JER|49|28|ad Cedar et ad regna Asor quae percussit Nabuchodonosor rex Babylonis haec dicit Dominus surgite ascendite ad Cedar et vastate filios orientis
JER|49|29|tabernacula eorum et greges eorum capient pelles eorum et omnia vasa eorum et camelos eorum tollent sibi et vocabunt super eos formidinem in circuitu
JER|49|30|fugite abite vehementer in voraginibus sedete qui habitatis Asor ait Dominus iniit enim contra vos Nabuchodonosor rex Babylonis consilium et cogitavit adversum vos cogitationes
JER|49|31|consurgite et ascendite ad gentem quietam et habitantem confidenter ait Dominus non ostia non vectes ei soli habitant
JER|49|32|et erunt cameli eorum in direptionem et multitudo iumentorum in praedam et dispergam eos in omnem ventum qui sunt adtonsi in comam et ex omni confinio eorum adducam interitum super eos ait Dominus
JER|49|33|et erit Asor in habitaculum draconum deserta usque in aeternum non manebit ibi vir nec incolet eam filius hominis
JER|49|34|quod factum est verbum Domini ad Hieremiam prophetam adversus Aelam in principio regni Sedeciae regis Iuda dicens
JER|49|35|haec dicit Dominus exercituum ecce ego confringam arcum Aelam summam fortitudinem eorum
JER|49|36|et inducam super Aelam quattuor ventos a quattuor plagis caeli et ventilabo eos in omnes ventos istos et non erit gens ad quam non perveniant profugi Aelam
JER|49|37|et pavere faciam Aelam coram inimicis suis et in conspectu quaerentium animam eorum et adducam super eos malum iram furoris mei dicit Dominus et emittam post eos gladium donec consumam eos
JER|49|38|et ponam solium meum in Aelam et perdam inde reges et principes ait Dominus
JER|49|39|in novissimis autem diebus reverti faciam captivos Aelam dicit Dominus
JER|50|1|verbum quod locutus est Dominus de Babylone et de terra Chaldeorum in manu Hieremiae prophetae
JER|50|2|adnuntiate in gentibus et auditum facite levate signum praedicate et nolite celare dicite capta est Babylon confusus est Bel victus est Marodach confusa sunt sculptilia eius superata sunt idola eorum
JER|50|3|quoniam ascendit contra eam gens ab aquilone quae ponet terram eius in solitudinem et non erit qui habitet in ea ab homine usque ad pecus et moti sunt et abierunt
JER|50|4|in diebus illis et in tempore illo ait Dominus venient filii Israhel ipsi et filii Iuda simul ambulantes et flentes properabunt et Dominum Deum suum quaerent
JER|50|5|in Sion interrogabunt viam huc facies eorum venient et adponentur ad Dominum foedere sempiterno quod nulla oblivione delebitur
JER|50|6|grex perditus factus est populus meus pastores eorum seduxerunt eos feceruntque vagari in montibus de monte in collem transierunt obliti sunt cubilis sui
JER|50|7|omnes qui invenerunt comederunt eos et hostes eorum dixerunt non peccavimus pro eo quod peccaverunt Domino decori iustitiae et expectationi patrum eorum Domino
JER|50|8|recedite de medio Babylonis et de terra Chaldeorum egredimini et estote quasi hedi ante greges
JER|50|9|quoniam ecce ego suscito et adducam in Babylonem congregationem gentium magnarum de terra aquilonis et praeparabuntur adversum eam et inde capietur sagitta eius quasi viri fortis interfectoris non revertetur vacua
JER|50|10|et erit Chaldea in praedam omnes vastantes eam replebuntur ait Dominus
JER|50|11|quoniam exultatis et magna loquimini diripientes hereditatem meam quoniam effusi estis sicut vitulus super herbam et mugistis ut tauri
JER|50|12|confusa est mater vestra nimis et adaequata pulveri quae genuit vos ecce novissima erit in gentibus deserta invia et arens
JER|50|13|ab ira Domini non habitabitur sed redigetur tota in solitudinem omnis qui transit per Babylonem stupebit et sibilabit super universis plagis eius
JER|50|14|praeparamini contra Babylonem per circuitum omnes qui intenditis arcum debellate eam non parcatis iaculis quia Domino peccavit
JER|50|15|clamate adversus eam ubique dedit manum ceciderunt fundamenta eius destructi sunt muri eius quoniam ultio Domini est ultionem accipite de ea sicut fecit facite ei
JER|50|16|disperdite satorem de Babylone et tenentem falcem in tempore messis a facie gladii columbae unusquisque ad populum suum convertetur et singuli ad terram suam fugient
JER|50|17|grex dispersus Israhel leones eiecerunt eum primus comedit eum rex Assur iste novissimus exossavit eum Nabuchodonosor rex Babylonis
JER|50|18|propterea haec dicit Dominus exercituum Deus Israhel ecce ego visitabo regem Babylonis et terram eius sicut visitavi regem Assur
JER|50|19|et reducam Israhel ad habitaculum suum et pascetur Carmelum et Basan et in monte Ephraim et Galaad saturabitur anima eius
JER|50|20|in diebus illis et in tempore illo ait Dominus quaeretur iniquitas Israhel et non erit et peccatum Iuda et non invenietur quoniam propitius ero eis quos reliquero
JER|50|21|super terram dominantium ascende et super habitatores eius visita dissipa et interfice quae post eos sunt ait Dominus et fac iuxta omnia quae praecepi tibi
JER|50|22|vox belli in terra et contritio magna
JER|50|23|quomodo confractus est et contritus est malleus universae terrae quomodo versa est in desertum Babylon in gentibus
JER|50|24|inlaqueavi te et capta es Babylon et nesciebas inventa es et adprehensa quoniam Dominum provocasti
JER|50|25|aperuit Dominus thesaurum suum et protulit vasa irae suae quoniam opus est Domino Deo exercituum in terra Chaldeorum
JER|50|26|venite ad eam ab extremis finibus aperite ut exeant qui conculcent eam tollite de via lapides et redigite in acervos et interficite eam nec sit quicquam reliquum
JER|50|27|dissipate universos fortes eius descendant in occisionem vae eis quia venit dies eorum tempus visitationis eorum
JER|50|28|vox fugientium et eorum qui evaserunt de terra Babylonis ut adnuntient in Sion ultionem Domini Dei nostri ultionem templi eius
JER|50|29|adnuntiate in Babylonem plurimis omnibus qui tendunt arcum consistite adversum eam per gyrum et nullus evadat reddite ei secundum opus suum iuxta omnia quae fecit facite illi quia contra Dominum erecta est adversum Sanctum Israhel
JER|50|30|idcirco cadent iuvenes eius in plateis eius et omnes viri bellatores eius conticescent in die illa ait Dominus
JER|50|31|ecce ego ad te superbe dicit Dominus Deus exercituum quia venit dies tuus tempus visitationis tuae
JER|50|32|et cadet superbus et corruet et non erit qui suscitet eum et succendam ignem in urbibus eius et devorabit omnia in circuitu eius
JER|50|33|haec dicit Dominus exercituum calumniam sustinent filii Israhel et filii Iuda simul omnes qui ceperunt eos tenent nolunt dimittere eos
JER|50|34|redemptor eorum Fortis Dominus exercituum nomen eius iudicio defendet causam eorum ut exterreat terram et commoveat habitatores Babylonis
JER|50|35|gladius ad Chaldeos ait Dominus et ad habitatores Babylonis et ad principes et ad sapientes eius
JER|50|36|gladius ad divinos eius qui stulti erunt gladius ad fortes illius qui timebunt
JER|50|37|gladius ad equos eius et ad currus eius et ad omne vulgus quod est in medio eius et erunt quasi mulieres gladius ad thesauros eius qui diripientur
JER|50|38|siccitas super aquas eius erit et arescent quia terra sculptilium est et in portentis gloriantur
JER|50|39|propterea habitabunt dracones cum fatuis ficariis et habitabunt in ea strutiones et non habitabitur ultra usque ad sempiternum nec extruetur usque ad generationem et generationem
JER|50|40|sicut subvertit Deus Sodomam et Gomorram et vicinas eius ait Dominus non habitabit ibi vir nec incolet eam filius hominis
JER|50|41|ecce populus venit ab aquilone et gens magna et reges multi consurgent a finibus terrae
JER|50|42|arcum et scutum adprehendent crudeles sunt et inmisericordes vox eorum quasi mare sonabit et super equos ascendent sicut vir paratus ad proelium contra te filia Babylon
JER|50|43|audivit rex Babylonis famam eorum et dissolutae sunt manus eius angustia adprehendit eum dolor quasi parturientem
JER|50|44|ecce quasi leo ascendet de superbia Iordanis ad pulchritudinem robustam quia subito currere eum faciam ad illam et quis erit electus quem praeponam ei quis enim similis mei et quis sustinebit me et quis est iste pastor qui resistat vultui meo
JER|50|45|propterea audite consilium Domini quod mente concepit adversum Babylonem et cogitationes eius quas cogitavit super terram Chaldeorum nisi detraxerint eos parvuli gregum nisi dissipatum fuerit cum ipsis habitaculum eorum
JER|50|46|a voce captivitatis Babylonis commota est terra et clamor inter gentes auditus est
JER|51|1|haec dicit Dominus ecce ego suscitabo super Babylonem et super habitatores eius qui cor suum levaverunt contra me quasi ventum pestilentem
JER|51|2|et mittam in Babylonem ventilatores et ventilabunt eam et demolientur terram eius quoniam venerunt super eam undique in die adflictionis eius
JER|51|3|non tendat qui tendit arcum suum et non ascendat loricatus nolite parcere iuvenibus eius interficite omnem militiam eius
JER|51|4|et cadent interfecti in terra Chaldeorum et vulnerati in regionibus eius
JER|51|5|quoniam non fuit viduatus Israhel et Iuda a Deo suo Domino exercituum terra autem eorum repleta est delicto a Sancto Israhel
JER|51|6|fugite de medio Babylonis et salvet unusquisque animam suam nolite tacere super iniquitatem eius quoniam tempus ultionis est Domino vicissitudinem ipse retribuet ei
JER|51|7|calix aureus Babylon in manu Domini inebrians omnem terram de vino eius biberunt gentes et ideo commotae sunt
JER|51|8|subito cecidit Babylon et contrita est ululate super eam tollite resinam ad dolorem eius si forte sanetur
JER|51|9|curavimus Babylonem et non est sanata derelinquamus eam et eamus unusquisque in terram suam quoniam pervenit usque ad caelos iudicium eius et elevatum est usque ad nubes
JER|51|10|protulit Dominus iustitias nostras venite et narremus in Sion opus Domini Dei nostri
JER|51|11|acuite sagittas implete faretras suscitavit Dominus spiritum regum Medorum et contra Babylonem mens eius ut perdat eam quoniam ultio Domini est ultio templi sui
JER|51|12|super muros Babylonis levate signum augete custodiam levate custodes praeparate insidias quia cogitavit Dominus et fecit quaecumque locutus est contra habitatores Babylonis
JER|51|13|quae habitas super aquas multas locuples in thesauris venit finis tuus pedalis praecisionis tuae
JER|51|14|iuravit Dominus exercituum per animam suam quoniam replebo te hominibus quasi brucho et super te celeuma cantabitur
JER|51|15|qui fecit terram in fortitudine sua praeparavit orbem in sapientia sua et prudentia sua extendit caelos
JER|51|16|dante eo vocem multiplicantur aquae in caelo qui levat nubes ab extremo terrae fulgura in pluviam fecit et produxit ventum de thesauris suis
JER|51|17|stultus factus est omnis homo ab scientia confusus est omnis conflator in sculptili quia mendax conflatio eius nec est spiritus in eis
JER|51|18|vana sunt opera et risu digna in tempore visitationis suae peribunt
JER|51|19|non sicut haec pars Iacob quia qui fecit omnia ipse est et Israhel sceptrum hereditatis eius Dominus exercituum nomen eius
JER|51|20|conlidis tu mihi vasa belli et ego conlidam in te gentes et disperdam in te regna
JER|51|21|et conlidam in te equum et equitem eius et conlidam in te currum et ascensorem eius
JER|51|22|et conlidam in te virum et mulierem et conlidam in te senem et puerum et conlidam in te iuvenem et virginem
JER|51|23|et conlidam in te pastorem et gregem eius et conlidam in te agricolam et iugales eius et conlidam in te duces et magistratus
JER|51|24|et reddam Babyloni et cunctis habitatoribus Chaldeae omne malum suum quod fecerunt in Sion in oculis vestris ait Dominus
JER|51|25|ecce ego ad te mons pestifer ait Dominus qui corrumpis universam terram et extendam manum meam super te et evolvam te de petris et dabo te in montem conbustionis
JER|51|26|et non tollent de te lapidem in angulum et lapidem in fundamenta sed perditus in aeternum eris ait Dominus
JER|51|27|levate signum in terra clangite bucina in gentibus sanctificate super eam gentes adnuntiate contra illam regibus Ararat Menni et Aschenez numerate contra eam Thapsar adducite equum quasi bruchum aculeatum
JER|51|28|sanctificate contra eam gentes reges Mediae duces eius et universos magistratus eius cunctamque terram potestatis eius
JER|51|29|et commovebitur terra et turbabitur quia evigilavit contra Babylonem cogitatio Domini ut ponat terram Babylonis desertam et inhabitabilem
JER|51|30|cessaverunt fortes Babylonis a proelio habitaverunt in praesidiis devoratum est robur eorum et facti sunt quasi mulieres incensa sunt tabernacula eius contriti sunt vectes eius
JER|51|31|currens obviam currenti veniet et nuntius obvius nuntianti ut adnuntiet regi Babylonis quia capta est civitas eius a summo usque ad summum
JER|51|32|et vada praeoccupata sunt et paludes incensae sunt igni et viri bellatores conturbati sunt
JER|51|33|quia haec dicit Dominus exercituum Deus Israhel filia Babylon quasi area tempus triturae eius adhuc modicum et veniet tempus messionis eius
JER|51|34|comedit me devoravit me Nabuchodonosor rex Babylonis reddidit me quasi vas inane absorbuit me sicut draco replevit ventrem suum teneritudine mea et eiecit me
JER|51|35|iniquitas adversum me et caro mea super Babylonem dicit habitatio Sion et sanguis meus super habitatores Chaldeae dicit Hierusalem
JER|51|36|propterea haec dicit Dominus ecce ego iudicabo causam tuam et ulciscar ultionem tuam et desertum faciam mare eius et siccabo venam eius
JER|51|37|et erit Babylon in tumulos habitatio draconum stupor et sibilus eo quod non sit habitator
JER|51|38|simul ut leones rugient excutient comas velut catuli leonum
JER|51|39|in calore eorum ponam potus eorum et inebriabo eos ut sopiantur et dormiant somnum sempiternum et non consurgant dicit Dominus
JER|51|40|deducam eos quasi agnos ad victimam quasi arietes cum hedis
JER|51|41|quomodo capta est Sesach et conprehensa est inclita universae terrae quomodo facta est in stuporem Babylon inter gentes
JER|51|42|ascendit super Babylonem mare multitudine fluctuum eius operta est
JER|51|43|factae sunt civitates eius in stuporem terra inhabitabilis et deserta terra in qua nullus habitet nec transeat per eam filius hominis
JER|51|44|et visitabo super Bel in Babylone et eiciam quod absorbuerat de ore eius et non confluent ad eum ultra gentes siquidem et murus Babylonis corruit
JER|51|45|egredimini de medio eius populus meus ut salvet unusquisque animam suam ab ira furoris Domini
JER|51|46|et ne forte mollescat cor vestrum et timeatis auditum qui audietur in terra et veniet in anno auditio et post hunc annum auditio et iniquitas in terra et dominator super dominatorem
JER|51|47|propterea ecce dies veniunt et visitabo super sculptilia Babylonis et omnis terra eius confundetur et universi interfecti eius cadent in medio eius
JER|51|48|et laudabunt super Babylonem caeli et terra et omnia quae in eis sunt quia ab aquilone venient ei praedones ait Dominus
JER|51|49|et quomodo fecit Babylon ut caderent occisi in Israhel sic de Babylone cadent occisi in universa terra
JER|51|50|qui fugistis gladium venite nolite stare recordamini procul Domini et Hierusalem ascendat super cor vestrum
JER|51|51|confusi sumus quoniam audivimus obprobrium operuit ignominia facies nostras quia venerunt alieni super sanctificationem domus Domini
JER|51|52|propterea ecce dies veniunt ait Dominus et visitabo super sculptilia eius et in omni terra eius mugiet vulneratus
JER|51|53|si ascenderit Babylon in caelum et firmaverit in excelso robur suum a me venient vastatores eius ait Dominus
JER|51|54|vox clamoris de Babylone et contritio magna de terra Chaldeorum
JER|51|55|quoniam vastavit Dominus Babylonem et perdidit ex ea vocem magnam et sonabunt fluctus eorum quasi aquae multae dedit sonitum vox eorum
JER|51|56|quia venit super eam id est super Babylonem praedo et adprehensi sunt fortes eius et emarcuit arcus eorum quia fortis ultor Dominus reddens retribuet
JER|51|57|et inebriabo principes eius et sapientes eius duces eius et magistratus eius et fortes eius et dormient somnum sempiternum et non expergiscentur ait Rex Dominus exercituum nomen eius
JER|51|58|haec dicit Dominus exercituum murus Babylonis ille latissimus suffossione suffodietur et portae eius excelsae igni conburentur et labores populorum ad nihilum et gentium in igne erunt et disperibunt
JER|51|59|verbum quod praecepit Hieremias prophetes Saraiae filio Neriae filii Maasiae cum pergeret cum Sedecia rege in Babylonem in anno quarto regni eius Saraias autem erat princeps prophetiae
JER|51|60|et scripsit Hieremias omne malum quod venturum erat super Babylonem in libro uno omnia verba haec quae scripta sunt contra Babylonem
JER|51|61|et dixit Hieremias ad Saraiam cum veneris Babylonem et videris et legeris omnia verba haec
JER|51|62|dices Domine tu locutus es contra locum istum ut disperderes eum ne sit qui in eo habitet ab homine usque ad pecus et ut sit perpetua solitudo
JER|51|63|cumque conpleveris legere librum istum ligabis ad eum lapidem et proicies illum in medio Eufraten
JER|51|64|et dices sic submergetur Babylon et non consurget a facie adflictionis quam ego adduco super eam et dissolventur hucusque verba Hieremiae
JER|52|1|filius viginti et unius anni Sedecias cum regnare coepisset et undecim annis regnavit in Hierusalem et nomen matris eius Amithal filia Hieremiae de Lobna
JER|52|2|et fecit malum in oculis Domini iuxta omnia quae fecerat Ioachim
JER|52|3|quoniam furor Domini erat in Hierusalem et in Iuda usquequo proiceret eos a facie sua et recessit Sedecias a rege Babylonis
JER|52|4|factum est autem in anno nono regni eius in mense decimo decima mensis venit Nabuchodonosor rex Babylonis ipse et omnis exercitus eius adversum Hierusalem et obsederunt eam et aedificaverunt contra eam munitiones in circuitu
JER|52|5|et fuit civitas obsessa usque ad undecimum annum regis Sedeciae
JER|52|6|mense autem quarto nona mensis obtinuit fames in civitate et non erant alimenta populo terrae
JER|52|7|et disrupta est civitas et omnes viri bellatores fugerunt et exierunt de civitate nocte per viam portae quae est inter duos muros et ducit ad hortum regis Chaldeis obsidentibus urbem in gyro et abierunt per viam quae ducit in heremum
JER|52|8|persecutus est autem exercitus Chaldeorum regem et adprehenderunt Sedeciam in deserto quod est iuxta Hiericho et omnis comitatus eius diffugit ab eo
JER|52|9|cumque conprehendissent regem adduxerunt eum ad regem Babylonis in Reblatha quae est in terra Emath et locutus est ad eum iudicia
JER|52|10|et iugulavit rex Babylonis filios Sedeciae in oculis eius sed et omnes principes Iudae occidit in Reblatha
JER|52|11|et oculos Sedeciae eruit et vinxit eum conpedibus et adduxit eum rex Babylonis in Babylonem et posuit eum in domo carceris usque ad diem mortis eius
JER|52|12|in mense autem quinto decima mensis ipse est annus nonusdecimus Nabuchodonosor regis Babylonis venit Nabuzardan princeps militiae qui stabat coram rege Babylonis in Hierusalem
JER|52|13|et incendit domum Domini et domum regis et omnes domos Hierusalem et omnem domum magnam igne conbusit
JER|52|14|et totum murum Hierusalem per circuitum destruxit cunctus exercitus Chaldeorum qui erat cum magistro militiae
JER|52|15|de pauperibus autem populi et de reliquo vulgo quod remanserat in civitate et de perfugis qui transfugerant ad regem Babylonis et ceteros de multitudine transtulit Nabuzardan princeps militiae
JER|52|16|de pauperibus vero terrae reliquit Nabuzardan princeps militiae in vinitores et in agricolas
JER|52|17|columnas quoque aereas quae erant in domo Domini et bases et mare aereum quod erat in domo Domini confregerunt Chaldei et tulerunt omne aes eorum in Babylonem
JER|52|18|et lebetas et creagras et psalteria et fialas et mortariola et omnia vasa aerea quae in ministerio fuerant tulerunt
JER|52|19|et hydrias et thymiamateria et urceos et pelves et candelabra et mortaria et cyatos quotquot aurea aurea et quotquot argentea argentea tulit magister militiae
JER|52|20|columnas duas et mare unum vitulos duodecim aereos qui erant sub basibus quas fecerat rex Salomon in domo Domini non erat pondus aeris omnium vasorum horum
JER|52|21|de columnis autem decem et octo cubiti altitudinis erant in columna una et funiculus duodecim cubitorum circuibat eam porro grossitudo eius quattuor digitorum et intrinsecus cava erat
JER|52|22|et capitella super utramque aerea altitudo capitelli unius quinque cubitorum et retiacula et mala granata
JER|52|23|nonaginta sex dependentia omnia mala granata centum retiaculis circumdabantur
JER|52|24|et tulit magister militiae Saraiam sacerdotem primum et Sophoniam sacerdotem secundum et tres custodes vestibuli
JER|52|25|et de civitate tulit eunuchum unum qui erat praepositus super viros bellatores et septem viros de his qui videbant faciem regis qui inventi sunt in civitate et scribam principem militum qui probabat tirones et sexaginta viros de populo terrae qui inventi sunt in medio civitatis
JER|52|26|tulit autem eos Nabuzardan magister militiae et duxit eos ad regem Babylonis in Reblatha
JER|52|27|et percussit eos rex Babylonis et interfecit eos in Reblatha in terra Emath et translatus est Iuda de terra sua
JER|52|28|iste est populus quem transtulit Nabuchodonosor in anno septimo Iudaeos tria milia et viginti tres
JER|52|29|in anno octavodecimo Nabuchodonosor de Hierusalem animas octingentas triginta duas
JER|52|30|in anno vicesimo tertio Nabuchodonosor transtulit Nabuzardan magister militiae Iudaeorum animas septingentas quadraginta quinque omnes ergo animae quattuor milia sescentae
JER|52|31|et factum est in tricesimo septimo anno transmigrationis Ioachim regis Iudae duodecimo mense vicesima quinta mensis elevavit Evilmerodach rex Babylonis ipso anno regni sui caput Ioachim regis Iudae et eduxit eum de domo carceris
JER|52|32|et locutus est cum eo bona et posuit thronum eius super thronos regum qui erant post se in Babylone
JER|52|33|et mutavit vestimenta carceris eius et comedebat panem coram eo semper cunctis diebus vitae suae
JER|52|34|et cibaria eius cibaria perpetua dabantur ei a rege Babylonis statuta per singulos dies usque ad diem mortis suae cunctis diebus vitae eius
