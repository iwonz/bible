JUDE|1|1|Iudas Iesu Christi servus, frater autem Iacobi, his qui sunt vocati, in Deo Patre dilecti et Christo Iesu conservati:
JUDE|1|2|misericordia vobis et pax et caritas adimpleatur.
JUDE|1|3|Carissimi, omnem sollicitudinem faciens scribendi vobis de communi nostra salute, necesse habui scribere vobis, deprecans certare pro semel tradita sanctis fide.
JUDE|1|4|Subintroierunt enim quidam homines, qui olim praescripti sunt in hoc iudicium, impii, Dei nostri gratiam transferentes in luxuriam, et solum Dominatorem et Dominum nostrum Iesum Christum negantes.
JUDE|1|5|Commonere autem vos volo, scientes vos omnia, quoniam Dominus semel populum de terra Aegypti salvans, secundo eos, qui non crediderunt, perdidit;
JUDE|1|6|angelos vero, qui non servaverunt suum principatum, sed dereliquerunt suum domicilium, in iudicium magni diei vinculis aeternis sub caligine reservavit.
JUDE|1|7|Sicut Sodoma et Gomorra et finitimae civitates, simili modo exfornicatae et abeuntes post carnem alteram, factae sunt exemplum, ignis aeterni poenam sustinentes.
JUDE|1|8|Similiter vero et hi somniantes carnem quidem maculant, dominationem autem spernunt, glorias autem blasphemant.
JUDE|1|9|Cum Michael archangelus cum Diabolo disputans altercaretur de Moysis corpore, non est ausus iudicium inferre blasphemiae, sed dixit: " Increpet te Dominus! ".
JUDE|1|10|Hi autem, quaecumque quidem ignorant, blasphemant; quaecumque autem naturaliter tamquam muta animalia norunt, in his corrumpuntur.
JUDE|1|11|Vae illis, quia via Cain abierunt et errore Balaam mercede effusi sunt et contradictione Core perierunt!
JUDE|1|12|Hi sunt in agapis vestris maculae, convivantes sine timore, semetipsos pascentes; nubes sine aqua, quae a ventis circumferuntur; arbores autumnales infructuosae bis mortuae, eradicatae;
JUDE|1|13|fluctus feri maris despumantes suas confusiones; sidera errantia, quibus procella tenebrarum in aeternum servata est.
JUDE|1|14|Prophetavit autem et his septimus ab Adam Henoch dicens: " Ecce venit Dominus in sanctis milibus suis
JUDE|1|15|facere iudicium contra omnes et arguere omnem animam de omnibus operibus impietatis eorum, quibus impie egerunt, et de omnibus duris, quae locuti sunt contra eum peccatores impii ".
JUDE|1|16|Hi sunt murmuratores, querelosi, secundum concupiscentias suas ambulantes, et os illorum loquitur superba, mirantes personas quaestus causa.
JUDE|1|17|Vos autem, carissimi, memores estote verborum, quae praedicta sunt ab apostolis Domini nostri Iesu Christi,
JUDE|1|18|quoniam dicebant vobis: " In novissimo tempore venient illusores, secundum suas concupiscentias ambulantes impietatum".
JUDE|1|19|Hi sunt qui segregant, animales, Spiritum non habentes.
JUDE|1|20|Vos autem, carissimi, superaedificantes vosmetipsos sanctissimae vestrae fidei, in Spiritu Sancto orantes,
JUDE|1|21|ipsos vos in dilectione Dei servate, exspectantes misericordiam Domini nostri Iesu Christi in vitam aeternam.
JUDE|1|22|Et his quidem miseremini disputantibus;
JUDE|1|23|illos vero salvate de igne rapientes; aliis autem miseremini in timore, odientes et eam, quae carnalis est, maculatam tunicam.
JUDE|1|24|Ei autem, qui potest vos conservare sine peccato et constituere ante conspectum gloriae suae immaculatos in exsultatione,
JUDE|1|25|soli Deo salvatori nostro per Iesum Christum Dominum nostrum gloria, magnificentia, imperium et potestas ante omne saeculum et nunc et in omnia saecula. Amen.
