3JOHN|1|1|The elder, To my dear friend Gaius, whom I love in the truth.
3JOHN|1|2|Dear friend, I pray that you may enjoy good health and that all may go well with you, even as your soul is getting along well.
3JOHN|1|3|It gave me great joy to have some brothers come and tell about your faithfulness to the truth and how you continue to walk in the truth.
3JOHN|1|4|I have no greater joy than to hear that my children are walking in the truth.
3JOHN|1|5|Dear friend, you are faithful in what you are doing for the brothers, even though they are strangers to you.
3JOHN|1|6|They have told the church about your love. You will do well to send them on their way in a manner worthy of God.
3JOHN|1|7|It was for the sake of the Name that they went out, receiving no help from the pagans.
3JOHN|1|8|We ought therefore to show hospitality to such men so that we may work together for the truth.
3JOHN|1|9|I wrote to the church, but Diotrephes, who loves to be first, will have nothing to do with us.
3JOHN|1|10|So if I come, I will call attention to what he is doing, gossiping maliciously about us. Not satisfied with that, he refuses to welcome the brothers. He also stops those who want to do so and puts them out of the church.
3JOHN|1|11|Dear friend, do not imitate what is evil but what is good. Anyone who does what is good is from God. Anyone who does what is evil has not seen God.
3JOHN|1|12|Demetrius is well spoken of by everyone--and even by the truth itself. We also speak well of him, and you know that our testimony is true.
3JOHN|1|13|I have much to write you, but I do not want to do so with pen and ink.
3JOHN|1|14|I hope to see you soon, and we will talk face to face. Peace to you. The friends here send their greetings. Greet the friends there by name.
