EPH|1|1|Paulus, apostolus Christi Iesu per voluntatem Dei, sanctis, qui sunt Ephesi, et fidelibus in Christo Iesu:
EPH|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
EPH|1|3|Benedictus Deus et Pater Domini nostri Iesu Christi,qui benedixit nos in omni benedictione spiritali in caelestibus in Christo,
EPH|1|4|sicut elegit nos in ipso ante mundi constitutionem,ut essemus sancti et immaculati in conspectu eius in caritate;
EPH|1|5|qui praedestinavit nos in adoptionem filiorumper Iesum Christum in ipsum,secundum beneplacitum voluntatis suae,
EPH|1|6|in laudem gloriae gratiae suae,in qua gratificavit nos in Dilecto,
EPH|1|7|in quo habemus redemptionem per sanguinem eius,remissionem peccatorum,secundum divitias gratiae eius,
EPH|1|8|quam superabundare fecit in nobisin omni sapientia et prudentia,
EPH|1|9|notum faciens nobis mysterium voluntatis suae,secundum beneplacitum eius, quod proposuit in eo,
EPH|1|10|in dispensationem plenitudinis temporum:recapitulare omnia in Christo,quae in caelis et quae in terra, in ipso;
EPH|1|11|in quo etiam sorte vocati sumus, praedestinati secundum propositum eius, qui omnia operatur secundum consilium voluntatis suae,
EPH|1|12|ut simus in laudem gloriae eius, qui ante speravimus in Christo;
EPH|1|13|in quo et vos cum audissetis verbum veritatis, evangelium salutis vestrae, in quo et credentes signati estis Spiritu promissionis Sancto,
EPH|1|14|qui est arrabo hereditatis nostrae in redemptionem acquisitionis, in laudem gloriae ipsius.
EPH|1|15|Propterea et ego audiens fidem vestram, quae est in Domino Iesu, et dilectionem in omnes sanctos,
EPH|1|16|non cesso gratias agens pro vobis memoriam faciens in orationibus meis,
EPH|1|17|ut Deus Domini nostri Iesu Christi, Pater gloriae, det vobis Spiritum sapientiae et revelationis in agnitione eius,
EPH|1|18|illuminatos oculos cordis vestri, ut sciatis quae sit spes vocationis eius, quae divitiae gloriae hereditatis eius in sanctis,
EPH|1|19|et quae sit supereminens magnitudo virtutis eius in nos, qui credimus, secundum operationem potentiae virtutis eius,
EPH|1|20|quam operatus est in Christo, suscitans illum a mortuis et constituens ad dexteram suam in caelestibus
EPH|1|21|supra omnem principatum et potestatem et virtutem et dominationem et omne nomen, quod nominatur non solum in hoc saeculo sed et in futuro;
EPH|1|22|et omnia subiecit sub pedibus eius et ipsum dedit caput supra omnia ecclesiae,
EPH|1|23|quae est corpus ipsius, plenitudo eius, qui omnia in omnibus adimpletur.
EPH|2|1|Et vos, cum essetis mortui de lictis et peccatis vestris,
EPH|2|2|in qui bus aliquando ambulastis secundum saeculum mundi huius, secundum principem potestatis aeris, spiritus, qui nunc operatur in filios diffidentiae;
EPH|2|3|in quibus et nos omnes aliquando conversati sumus in concupiscentiis carnis nostrae, facientes voluntates carnis et cogitationum, et eramus natura filii irae, sicut et ceteri.
EPH|2|4|Deus autem, qui dives est in misericordia, propter nimiam caritatem suam, qua dilexit nos,
EPH|2|5|et cum essemus mortui peccatis, convivificavit nos Christo - gratia estis salvati -
EPH|2|6|et conresuscitavit et consedere fecit in caelestibus in Christo Iesu,
EPH|2|7|ut ostenderet in saeculis supervenientibus abundantes divitias gratiae suae in bonitate super nos in Christo Iesu.
EPH|2|8|Gratia enim estis salvati per fidem; et hoc non ex vobis, Dei donum est:
EPH|2|9|non ex operibus, ut ne quis glorietur.
EPH|2|10|Ipsius enim sumus factura, creati in Christo Iesu in opera bona, quae praeparavit Deus, ut in illis ambulemus.
EPH|2|11|Propter quod memores estote, quod aliquando vos gentes in carne, qui dicimini praeputium ab ea, quae dicitur circumcisio in carne manufacta,
EPH|2|12|quia eratis illo in tempore sine Christo, alienati a conversatione Israel et extranei testamentorum promissionis, spem non habentes et sine Deo in mundo.
EPH|2|13|Nunc autem in Christo Iesu vos, qui aliquando eratis longe, facti estis prope in sanguine Christi.
EPH|2|14|Ipse est enim pax nostra, qui fecit utraque unum et medium parietem maceriae solvit, inimicitiam, in carne sua,
EPH|2|15|legem mandatorum in decretis evacuans, ut duos condat in semetipso in unum novum hominem, faciens pacem,
EPH|2|16|et reconciliet ambos in uno corpore Deo per crucem, interficiens inimicitiam in semetipso.
EPH|2|17|Et veniens evangelizavit pacem vobis, qui longe fuistis, et pacem his, qui prope;
EPH|2|18|quoniam per ipsum habemus accessum ambo in uno Spiritu ad Patrem.
EPH|2|19|Ergo iam non estis extranei et advenae, sed estis concives sanctorum et domestici Dei,
EPH|2|20|superaedificati super fundamentum apostolorum et prophetarum, ipso summo angulari lapide Christo Iesu,
EPH|2|21|in quo omnis aedificatio compacta crescit in templum sanctum in Domino,
EPH|2|22|in quo et vos coaedificamini in habitaculum Dei in Spiritu.
EPH|3|1|Huius rei gratia, ego Paulus, vinctus Christi Iesu pro vobis gentibus -
EPH|3|2|si tamen audistis dispensationem gratiae Dei, quae data est mihi pro vobis,
EPH|3|3|quoniam secundum revelationem notum mihi factum est mysterium, sicut supra scripsi in brevi,
EPH|3|4|prout potestis legentes intellegere prudentiam meam in mysterio Christi,
EPH|3|5|quod aliis generationibus non innotuit filiis hominum, sicuti nunc revelatum est sanctis apostolis eius et prophetis in Spiritu,
EPH|3|6|esse gentes coheredes et concorporales et comparticipes promissionis in Christo Iesu per evangelium,
EPH|3|7|cuius factus sum minister secundum donum gratiae Dei, quae data est mihi secundum operationem virtutis eius.
EPH|3|8|Mihi omnium sanctorum minimo data est gratia haec: gentibus evangelizare investigabiles divitias Christi
EPH|3|9|et illuminare omnes, quae sit dispensatio mysterii absconditi a saeculis in Deo, qui omnia creavit,
EPH|3|10|ut innotescat nunc principatibus et potestatibus in caelestibus per ecclesiam multiformis sapientia Dei,
EPH|3|11|secundum propositum saeculorum, quod fecit in Christo Iesu Domino nostro,
EPH|3|12|in quo habemus fiduciam et accessum in confidentia per fidem eius.
EPH|3|13|Propter quod peto, ne deficiatis in tribulationibus meis pro vobis, quae est gloria vestra.
EPH|3|14|Huius rei gratia flecto genua mea ad Patrem,
EPH|3|15|ex quo omnis paternitas in caelis et in terra nominatur,
EPH|3|16|ut det vobis secundum divitias gloriae suae virtute corroborari per Spiritum eius in interiorem hominem,
EPH|3|17|habitare Christum per fidem in cordibus vestris, in caritate radicati et fundati,
EPH|3|18|ut valeatis comprehendere cum omnibus sanctis quae sit latitudo et longitudo et sublimitas et profundum,
EPH|3|19|scire etiam supereminentem scientiae caritatem Christi, ut impleamini in omnem plenitudinem Dei.
EPH|3|20|Ei autem, qui potens est supra omnia facere superabundanter quam petimus aut intellegimus, secundum virtutem, quae operatur in nobis,
EPH|3|21|ipsi gloria in ecclesia et in Christo Iesu in omnes generationes saeculi saeculorum. Amen.
EPH|4|1|Obsecro itaque vos ego, vinctus in Domino, ut digne ambuletis vocatione, qua vocati estis,
EPH|4|2|cum omni humilitate et mansuetudine, cum longanimitate, supportantes invicem in caritate,
EPH|4|3|solliciti servare unitatem spiritus in vinculo pacis;
EPH|4|4|unum corpus et unus Spiritus, sicut et vocati estis in una spe vocationis vestrae;
EPH|4|5|unus Dominus, una fides, unum baptisma;
EPH|4|6|unus Deus et Pater omnium, qui super omnes et per omnia et in omnibus.
EPH|4|7|Unicuique autem nostrum data est gratia secundum mensuram donationis Christi.
EPH|4|8|Propter quod dicit: Ascendens in altum captivam duxit captivitatem,dedit dona hominibus ".
EPH|4|9|Illud autem " ascendit " quid est, nisi quia et descendit in inferiores partes terrae?
EPH|4|10|Qui descendit, ipse est et qui ascendit super omnes caelos, ut impleret omnia.
EPH|4|11|Et ipse dedit quosdam quidem apostolos, quosdam autem prophetas, alios vero evangelistas, alios autem pastores et doctores
EPH|4|12|ad instructionem sanctorum in opus ministerii, in aedificationem corporis Christi,
EPH|4|13|donec occurramus omnes in unitatem fidei et agnitionis Filii Dei, in virum perfectum, in mensuram aetatis plenitudinis Christi,
EPH|4|14|ut iam non simus parvuli fluctuantes et circumacti omni vento doctrinae in fallacia hominum, in astutia ad circumventionem erroris;
EPH|4|15|veritatem autem facientes in caritate crescamus in illum per omnia, qui est caput Christus,
EPH|4|16|ex quo totum corpus compactum et conexum per omnem iuncturam subministrationis secundum operationem in mensura uniuscuiusque partis augmentum corporis facit in aedificationem sui in caritate.
EPH|4|17|Hoc igitur dico et testificor in Domino, ut iam non ambuletis, sicut et gentes ambulant in vanitate sensus sui
EPH|4|18|tenebris obscuratum habentes intellectum, alienati a vita Dei propter ignorantiam, quae est in illis propter caecitatem cordis ipsorum;
EPH|4|19|qui indolentes semetipsos tradiderunt impudicitiae in operationem immunditiae omnis in avaritia.
EPH|4|20|Vos autem non ita didicistis Christum,
EPH|4|21|si tamen illum audistis et in ipso edocti estis, sicut est veritas in Iesu:
EPH|4|22|deponere vos secundum pristinam conversationem veterem hominem, qui corrumpitur secundum desideria erroris,
EPH|4|23|renovari autem spiritu mentis vestrae
EPH|4|24|et induere novum hominem, qui secundum Deum creatus est in iustitia et sanctitate veritatis.
EPH|4|25|Propter quod deponentes mendacium loquimini veritatem unusquisque cum proximo suo, quoniam sumus invicem membra.
EPH|4|26|Irascimini et nolite peccare; sol non occidat super iracundiam vestram,
EPH|4|27|et nolite locum dare Diabolo.
EPH|4|28|Qui furabatur, iam non furetur, magis autem laboret operando manibus bonum, ut habeat unde tribuat necessitatem patienti.
EPH|4|29|Omnis sermo malus ex ore vestro non procedat, sed si quis bonus ad aedificationem opportunitatis, ut det gratiam audientibus.
EPH|4|30|Et nolite contristare Spiritum Sanctum Dei, in quo signati estis in diem redemptionis.
EPH|4|31|Omnis amaritudo et ira et indignatio et clamor et blasphemia tollatur a vobis cum omni malitia.
EPH|4|32|Estote autem invicem benigni, misericordes, donantes invicem, sicut et Deus in Christo donavit vobis.
EPH|5|1|Estote ergo imitatores Dei, sicut filii carissimi,
EPH|5|2|et ambulate in dilectione, sicut et Christus dilexit nos et tradidit seipsum pro nobis oblationem et hostiam Deo in odorem suavitatis.
EPH|5|3|Fornicatio autem et omnis immunditia aut avaritia nec nominetur in vobis, sicut decet sanctos,
EPH|5|4|et turpitudo et stultiloquium aut scurrilitas, quae non decent, sed magis gratiarum actio.
EPH|5|5|Hoc enim scitote intellegentes quod omnis fornicator aut immundus aut avarus, id est idolorum cultor, non habet hereditatem in regno Christi et Dei.
EPH|5|6|Nemo vos decipiat inanibus verbis; propter haec enim venit ira Dei in filios diffidentiae.
EPH|5|7|Nolite ergo effici comparticipes eorum;
EPH|5|8|eratis enim aliquando tenebrae, nunc autem lux in Domino. Ut filii lucis ambulate
EPH|5|9|- fructus enim lucis est in omni bonitate et iustitia et veritate -
EPH|5|10|probantes quid sit beneplacitum Domino;
EPH|5|11|et nolite communicare operibus infructuosis tenebrarum, magis autem et redarguite;
EPH|5|12|quae enim in occulto fiunt ab ipsis, turpe est et dicere;
EPH|5|13|omnia autem, quae arguuntur, a lumine manifestantur,
EPH|5|14|omne enim, quod manifestatur, lumen est. Propter quod dicit: " Surge, qui dormis, et exsurge a mortuis, et illuminabit te Christus ".
EPH|5|15|Videte itaque caute quomodo ambuletis, non quasi insipientes sed ut sapientes,
EPH|5|16|redimentes tempus, quoniam dies mali sunt.
EPH|5|17|Propterea nolite fieri imprudentes, sed intellegite, quae sit voluntas Domini.
EPH|5|18|Et nolite inebriari vino, in quo est luxuria, sed implemini Spiritu
EPH|5|19|loquentes vobismetipsis in psalmis et hymnis et canticis spiritalibus, cantantes et psallentes in cordibus vestris Domino.
EPH|5|20|Gratias agentes semper pro omnibus in nomine Domini nostri Iesu Christi Deo et Patri,
EPH|5|21|subiecti invicem in timore Christi.
EPH|5|22|Mulieres viris suis sicut Domino,
EPH|5|23|quoniam vir caput est mulieris, sicut et Christus caput est ecclesiae, ipse salvator corporis.
EPH|5|24|Sed ut ecclesia subiecta est Christo, ita et mulieres viris in omnibus.
EPH|5|25|Viri, diligite uxores, sicut et Christus dilexit ecclesiam et seipsum tradidit pro ea,
EPH|5|26|ut illam sanctificaret mundans lavacro aquae in verbo,
EPH|5|27|ut exhiberet ipse sibi gloriosam ecclesiam non habentem maculam aut rugam aut aliquid eiusmodi, sed ut sit sancta et immaculata.
EPH|5|28|Ita et viri debent diligere uxores suas ut corpora sua. Qui suam uxorem diligit, seipsum diligit;
EPH|5|29|nemo enim umquam carnem suam odio habuit, sed nutrit et fovet eam sicut et Christus ecclesiam,
EPH|5|30|quia membra sumus corporis eius.
EPH|5|31|Propter hoc relinquet homo patrem et matrem et adhaerebit uxori suae, et erunt duo in carne una.
EPH|5|32|Mysterium hoc magnum est; ego autem dico de Christo et ecclesia!
EPH|5|33|Verumtamen et vos singuli unusquisque suam uxorem sicut seipsum diligat; uxor autem timeat virum.
EPH|6|1|Filii, oboedite parentibus vestris in Domino; hoc enim est iu stum.
EPH|6|2|Honora patrem tuum et matrem, quod est mandatum primum cum promissione,
EPH|6|3|ut bene sit tibi, et sis longaevus super terram.
EPH|6|4|Et, patres, nolite ad iracundiam provocare filios vestros, sed educate illos in disciplina et correptione Domini.
EPH|6|5|Servi, oboedite dominis carnalibus cum timore et tremore, in simplicitate cordis vestri, sicut Christo;
EPH|6|6|non ad oculum servientes, quasi hominibus placentes, sed ut servi Christi facientes voluntatem Dei ex animo;
EPH|6|7|cum bona voluntate servientes, sicut Domino et non hominibus,
EPH|6|8|scientes quoniam unusquisque, si quid fecerit bonum, hoc percipiet a Domino, sive servus sive liber.
EPH|6|9|Et, domini, eadem facite illis, remittentes minas, scientes quia et illorum et vester Dominus est in caelis, et personarum acceptio non est apud eum.
EPH|6|10|De cetero confortamini in Domino et in potentia virtutis eius.
EPH|6|11|Induite armaturam Dei, ut possitis stare adversus insidias Diaboli.
EPH|6|12|Quia non est nobis colluctatio adversus sanguinem et carnem sed adversus principatus, adversus potestates, adversus mundi rectores tenebrarum harum, adversus spiritalia nequitiae in caelestibus.
EPH|6|13|Propterea accipite armaturam Dei, ut possitis resistere in die malo et, omnibus perfectis, stare.
EPH|6|14|State ergo succincti lumbos vestros in veritate et induti loricam iustitiae
EPH|6|15|et calceati pedes in praeparatione evangelii pacis,
EPH|6|16|inomnibus sumentes scutum fidei, in quo possitis omnia tela Maligni ignea exstinguere;
EPH|6|17|et galeam salutis assumite et gladium Spiritus, quod est verbum Dei;
EPH|6|18|per omnem orationem et obsecrationem orantes omni tempore in Spiritu, et in ipso vigilantes in omni instantia et obsecratione pro omnibus sanctis
EPH|6|19|et pro me, ut detur mihi sermo in aperitione oris mei cum fiducia notum facere mysterium evangelii,
EPH|6|20|pro quo legatione fungor in catena, ut in ipso audeam, prout oportet me, loqui.
EPH|6|21|Ut autem et vos sciatis, quae circa me sunt, quid agam, omnia nota vobis faciet Tychicus, carissimus frater et fidelis minister in Domino,
EPH|6|22|quem misi ad vos in hoc ipsum, ut cognoscatis, quae circa nos sunt, et consoletur corda vestra.
EPH|6|23|Pax fratribus et caritas cum fide a Deo Patre et Domino Iesu Christo.
EPH|6|24|Gratia cum omnibus, qui diligunt Dominum nostrum Iesum Christum in incorruptione.
