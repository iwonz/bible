JUDG|1|1|І сталося по смерті Ісуса, і питалися Ізраїлеві сини Господа, говорячи: Хто з нас вийде спереду на ханаанеянина, щоб воювати з ним?
JUDG|1|2|І сказав Господь: Юда піде. Оце Я дав Край у його руку.
JUDG|1|3|І сказав Юда до Симеона, свого брата: Іди зо мною на мій жеребок, і будемо воювати з ханаанеянином, то піду й я з тобою на твій жеребок. І пішов із ним Симеон.
JUDG|1|4|І піднявся Юда, а Господь дав ханаанеянина та періззеянина в їхню руку. І вони побили їх у Безеку, десять тисяч чоловіка.
JUDG|1|5|І знайшли вони в Безеку Адоні-Безека, і воювали з ним, і побили ханаанеянина та періззеянина.
JUDG|1|6|І втікав Адоні-Безек, а вони гналися за ним, і зловили його, і повідрубували великі пальці його рук та його ніг.
JUDG|1|7|І сказав Адоні-Безек: Сімдесят царів з відрубаними великими пальцями їхніх рук та їхніх ніг часто збирали поживу під столом моїм. Як робив я, так відплатив мені Бог!
JUDG|1|8|І воювали Юдині сини з Єрусалимом, і здобули його, і побили його вістрям меча, а місто пустили з огнем.
JUDG|1|9|А потому Юдині сини зійшли воювати з ханаанеянином, мешканцем гори, і Неґеву, і Шефелі.
JUDG|1|10|І пішов Юда до ханаанеянина, що сидить у Хевроні, а ім'я Хеврону було колись: Кір'ят-Арба, і побили Шешая, й Ахімана та Талмая.
JUDG|1|11|А звідти пішов він до мешканців Девіру, а ім'я Девіру колись: Кір'ят-Сефер.
JUDG|1|12|І сказав Калев: Хто поб'є Кір'ят-Сефер та здобуде його, то дам йому Ахсу, дочку мою, за жінку.
JUDG|1|13|І здобув його Отніїл, син Кенезів, брат Калевів, молодший від нього. І він дав йому свою дочку Ахсу за жінку.
JUDG|1|14|І сталося, коли вона прийшла, то намовила його жадати поля від її батька. І зійшла вона з осла, а Калев сказав їй: Що тобі?
JUDG|1|15|І вона сказала йому: Дай мені дара благословення! Бо ти дав мені землю суху, то дай мені водні джерела. І Калев дав їй Ґуллот-горішній та Ґуллот-долішній.
JUDG|1|16|А сини Кенея, Мойсеєвого тестя, пішли з міста Пальм з Юдиними синами до Юдиної пустині, що на півдні Араду. І пішов він, і осівся з народом.
JUDG|1|17|І пішов Юда з Симеоном, своїм братом, та й побили ханаанеянина, мешканця Цефату, і вчинили його закляттям. І назвав ім'я того міста: Хорма.
JUDG|1|18|І здобув Юда Аззу та границю її, й Ашкелон та границю його, і Екрон та границю його.
JUDG|1|19|І був Господь з Юдою, і він повиганяв мешканців гори. Та не міг він повиганяти мешканців долини, бо вони мали залізні колесниці.
JUDG|1|20|І дали Калевові Хеврон, як говорив був Мойсей, і він вигнав звідти трьох велетнів.
JUDG|1|21|А євусеянина, мешканця Єрусалиму, не вигнали Веніяминові сини, і осів євусеянин із Веніяминовими синами в Єрусалимі, і сидять тут аж до цього дня.
JUDG|1|22|І пішов також дім Йосипів до Бет-Елу, а Господь був з ними.
JUDG|1|23|І вивідав Йосипів дім у Бет-Елі, а ім'я того міста колись було Луз.
JUDG|1|24|І побачили сторожі чоловіка, що виходив із того міста, та й сказали до нього: Покажи нам вхід до міста, а ми вчинимо тобі милість!
JUDG|1|25|І він показав їм вхід до міста, і вони побили те місто вістрям меча, а того чоловіка та ввесь його рід відпустили.
JUDG|1|26|І пішов той чоловік до краю хіттеян, і збудував місто, та й назвав ім'я йому: Луз, воно ім'я його аж до цього дня.
JUDG|1|27|А Манасія не повиганяв мешканців Бет-Шеану та його залежних міст, і Таанаху та його залежних міст, і мешканців Дору та його залежних міст, і мешканців Ївлеаму та його залежних міст, і мешканців Міґіддо та його залежних міст, і ханаанеянин волів сидіти в тому краї.
JUDG|1|28|І сталося, коли Ізраїль зміцнився, то він наклав на ханаанеянина данину, але вигнати не вигнав його.
JUDG|1|29|І Єфрем не вигнав ханаанеянина, що мешкає в Ґезері, і осівся ханаанеянин серед нього в Ґезері.
JUDG|1|30|Завулон не повиганяв мешканців Кітрону та мешканців Нагалолу, і осівся ханаанеянин серед нього, і став за данину.
JUDG|1|31|Асир не повиганяв мешканців Акко, і мешканців Сидону, і Ахлаву, і Ахзіву, і Хелби, і Афіку, і Рехову.
JUDG|1|32|І осівся асирець серед ханаанеянина, мешканця того Краю, бо він не вигнав його.
JUDG|1|33|Нефталим не повиганяв мешканців Бет-Шемешу, і мешканців Бет-Анату, і він осівся серед ханаанеянина, мешканця того Краю, а мешканці Бет-Шемешу та Бет-Анату стали їм за данину.
JUDG|1|34|І тиснув амореянин Данових синів на гору, бо не давав йому сходити на долину.
JUDG|1|35|І волів амореянин сидіти на горі Херес в Айялоні та в Шаалевімі, та стала сильною рука Йосипового дому, він став за данину.
JUDG|1|36|А границя аморейська від Маале-Акраббім, і від Сели та вище.
JUDG|2|1|І прийшов Ангол Господній з Ґілґалу до Бохіму, та й сказав: Я вивів вас із Єгипту до того Краю, що присягнув був вашим батькам. І сказав Я: не зламаю Свого заповіту з вами повіки!
JUDG|2|2|А ви не складете заповіту з мешканцями цього Краю, їхні жертівники порозбиваєте, та не слухали ви Мого голосу. Що це ви зробили?
JUDG|2|3|І Я теж сказав: Не прожену їх від вас, і вони стануть вам терням у боки, а їхні боги стануть вам пасткою.
JUDG|2|4|І сталося, як Ангол Господній говорив ці слова до всіх Ізраїлевих синів, то народ підніс свій голос, та й заплакав.
JUDG|2|5|І назвали ім'я того місця: Бохім, і приносили там жертви Господеві.
JUDG|2|6|А Ісус відпустив народ, і Ізраїлеві сини розійшлися кожен до свого спадку, щоб посісти той Край.
JUDG|2|7|І служив народ Господеві по всі дні Ісуса та по всі дні старших, які продовжили дні свої по Ісусі, що бачили всякий великий чин Господа, якого зробив Він Ізраїлеві.
JUDG|2|8|І вмер Ісус, син Навинів, раб Господній, віку ста й десяти літ.
JUDG|2|9|І поховали його в межах спадщини його, у Тімнат-Хересі, в Єфремових горах, на північ від гори Ґааш.
JUDG|2|10|І також усе це покоління було прилучене до батьків своїх, а по них настало інше покоління, що не знало Господа, а також тих діл, які чинив Він Ізраїлеві.
JUDG|2|11|І Ізраїлеві сини чинили зло в Господніх очах, і служили Ваалам.
JUDG|2|12|І вони покинули Господа, Бога батьків своїх, що вивів їх із єгипетського краю, та й пішли за іншими богами, за богами тих народів, що були в їхніх околицях, і вклонялися їм, і гнівили Господа.
JUDG|2|13|І покинули вони Господа, та й служили Ваалові та Астартам.
JUDG|2|14|І запалав Господній гнів на Ізраїля, і Він дав їх у руку грабіжників, і вони їх грабували. І Він передав їх у руку навколишніх їхніх ворогів, і вони не могли вже встояти перед своїми ворогами.
JUDG|2|15|У всьому, де вони ходили, Господня рука була проти них на зло, як говорив був Господь, і як заприсягнув їм Господь. І Він дуже їх тиснув.
JUDG|2|16|І поставив Господь суддів, і вони рятували їх від руки їхніх грабіжників.
JUDG|2|17|Та вони не слухалися також своїх суддів, бо блудили за іншими богами, і вклонялися їм. Вони скоро відхилялися з тієї дороги, якою йшли їхні батьки, щоб слухатися Господніх наказів. Вони так не робили!
JUDG|2|18|А коли Господь ставив їм суддів, то Господь був із суддею, і рятував їх із руки їхніх ворогів по всі дні того судді, бо Господь жалував їх через їхній стогін через тих, що їх переслідували та гнобили їх.
JUDG|2|19|І бувало, як умирав той суддя, вони знову псувалися більше від своїх батьків, щоб іти за іншими богами, щоб їм служити та щоб їм вклонятися, і вони не кидали чинів своїх та своєї неслухняної дороги.
JUDG|2|20|І запалився Господній гнів на Ізраїля, і Він сказав: За те, що люд цей переступив Мого заповіта, що Я наказав був їхнім батькам, і не слухалися Мого голосу,
JUDG|2|21|тож Я більше не виганятиму перед ними нікого з тих народів, що Ісус позоставив, умираючи,
JUDG|2|22|щоб випробувати ними Ізраїля, чи держатимуться вони Господньої дороги, щоб нею ходити, як держалися їхні батьки, чи ні.
JUDG|2|23|І Господь позоставив тих людей, щоб їх скоро не виганяти, і не дав їх у руку Ісусову.
JUDG|3|1|А оце ті народи, що Господь позоставив на випробування ними Ізраїля, усі ті, що не знали всіх війн ханаанських,
JUDG|3|2|тільки щоб пізнали покоління Ізраїлевих синів, щоб навчити їх війни, тільки таких, що перед тим не знали їх:
JUDG|3|3|п'ять володарів филистимських, і всі ханаанеяни, і сидоняни, і хіввеяни, мешканці гори Ливану, від гори Баал-Гермон аж до виходу до Гамату.
JUDG|3|4|І були вони залишені на випробування ними Ізраїля, щоб пізнати, чи будуть вони слухатися заповідей Господа, які Він наказав був їхнім батькам через Мойсея.
JUDG|3|5|А Ізраїлеві сини сиділи серед ханаанеянина, хіттеянина, і амореянина, і періззеянина, і хіввеянина, і євусеянина.
JUDG|3|6|І вони брали їхніх дочок собі за жінок, а своїх дочок давали їхнім синам, та служили їхнім богам.
JUDG|3|7|І Ізраїлеві сини робили зло в Господніх очах, і забули Господа, Бога свого, та й служили Ваалам та Астартам.
JUDG|3|8|І запалився Господній гнів на Ізраїля, і Він передав їх у руку Кушан-Ріш'атаїма, царя Араму двох річок. І служили Ізраїлеві сини Кушан-Ріш'атаїмові вісім літ.
JUDG|3|9|І кликали Ізраїлеві сини до Господа, і Господь поставив для Ізраїлевих синів рятівника, і він врятував їх, Отніїла, сина Кеназа, брата Калева, молодшого від нього.
JUDG|3|10|І був на ньому Дух Господній, і судив він Ізраїля. І вийшов він на війну, і Господь дав у його руку Кушан-Ріш'атаїма, царя арамського. І була сильна рука його над Кушан-Ріш'атаїмом.
JUDG|3|11|І мав Край мир сорок літ, і помер Отніїл, син Кеназа.
JUDG|3|12|А Ізраїлеві сини й далі чинили зло в Господніх очах, і Господь зміцнив Еґлона, царя моавського, над Ізраїлем через те, що вони робили зло в Господніх очах.
JUDG|3|13|І зібрав він до себе синів Аммонових та Амаликових, та й пішов і підбив Ізраїля. І вони посіли Місто Пальм.
JUDG|3|14|І служили Ізраїлеві сини Еґлонові, цареві моавському, вісімнадцять літ.
JUDG|3|15|І кликали Ізраїлеві сини до Господа, і Господь поставив їм рятівника, Егуда, сина Ґерового, сина ємінеянина, чоловіка лівшу, з безвладною правою рукою. І послали Ізраїлеві сини через нього дарунка Еґлонові, цареві моавському.
JUDG|3|16|І зробив собі Егуд меча, а в нього два вістря, ґошед довжина його, він прип'яв його під своїм убранням на стегні своєї правиці.
JUDG|3|17|І приніс він того дарунка Еґлонові, цареві моавському. А Еґлон чоловік дуже товстий.
JUDG|3|18|І сталося, коли він скінчив підносити того дарунка, то відпустив тих, що несли того дарунка.
JUDG|3|19|А він вернувся від бовванів, що при Ґілґалі, та й сказав: У мене таємна справа до тебе, о царю! А той сказав: Тихо! І вийшли від нього всі, хто стояв при ньому.
JUDG|3|20|І Егуд увійшов до нього, а він сидить у прохолодній горниці, що була для нього самого. І сказав Егуд: Я маю Боже слово для тебе. І той устав із стільця.
JUDG|3|21|І простяг Егуд свою лівицю, і витяг меча з-над стегна своєї правиці, та й загнав його йому в живіт.
JUDG|3|22|І ввійшла також ручка за вістрям, а сало закрило за вістрям, бо він не витягнув меча з його живота. І ввійшло вістря до міжкроччя.
JUDG|3|23|І вийшов Егуд до сіней, і зачинив за собою двері тієї горниці, та й замкнув.
JUDG|3|24|І він вийшов. А царські раби ввійшли та й побачили, аж ось двері горниці замкнені. І вони сказали: Певне він для потреби своєї в прохолодному покої.
JUDG|3|25|І чекали вони аж допізна, а ото він не відчиняє дверей горниці. І взяли вони ключа, і відчинили, аж ось їхній пан лежить мертвий на землі!
JUDG|3|26|А Егуд утік, поки вони зволікались. І він перейшов ті боввани, і сховався втечею до Сеїру.
JUDG|3|27|І сталося, коли він прийшов, то засурмив у сурму на Єфремових горах. І Ізраїлеві сини зійшли з ним з гори, а він перед ними.
JUDG|3|28|І сказав він до них: Біжіть за мною, бо Господь дав у вашу руку ваших моавських ворогів! І зійшли вони за ним, і захопили йорданські переходи до Моаву, і не дали нікому перейти.
JUDG|3|29|І побили вони Моава того часу, близько десяти тисяч чоловіка, кожного кремезного й кожного сильного чоловіка, і ніхто не втік.
JUDG|3|30|І був того дня приборканий Моав під Ізраїлеву руку, а Край мав мир вісімдесят літ.
JUDG|3|31|А по ньому був Шамґар, син Аната. І побив він филистимлян шістсот чоловіка києм на худобу. І він теж урятував Ізраїля.
JUDG|4|1|А Ізраїлеві сини ще більше чинили зло в Господніх очах, а Егуд умер.
JUDG|4|2|І передав їх Господь у руку Явіна, царя ханаанського, що царював у Гацорі. А зверхником його війська був Сісера, і він сидів у Харошет-Ґаґґоїмі.
JUDG|4|3|І кликали Ізраїлеві сини до Господа, бо той мав дев'ятсот залізних колесниць, і він сильно утискав Ізраїлевих синів двадцять літ.
JUDG|4|4|А Девора пророчиця, жінка Лаппідота, вона судила Ізраїля того часу.
JUDG|4|5|І сиділа вона під Девориною Пальмою, між Рамою та між Бет-Елом в Єфремових горах, а Ізраїлеві сини приходили до неї на суд.
JUDG|4|6|І вона послала й покликала Барака, Авіноамового сина, з Кедешу Нефталимового. І сказала до нього: Ось наказав Господь, Бог Ізраїлів: Іди, зійдеш на гору фавор, і візьмеш з собою десять тисяч чоловіка з синів Нефталимових та з синів Завулонових.
JUDG|4|7|А я приведу до тебе, до Кішонської долини, Сісеру, начальника Явінового війська, і колесниці його, і натовп його, та й дам його в твою руку.
JUDG|4|8|І сказав до неї Барак: Якщо ти підеш зо мною, то піду, а якщо не підеш зо мною, не піду.
JUDG|4|9|А вона відказала: Піти піду з тобою, тільки не буде твоя слава на тій дорозі, якою ти підеш, бо в руку жінки Господь передасть Сісеру. І встала Девора, і пішла з Бараком до Кедешу.
JUDG|4|10|І скликав Барак Завулона та Нефталима до Кедешу, і пішло за ним десять тисяч чоловіка. І пішла з ним Девора.
JUDG|4|11|А кенеянин Хевер відділився від Каїна, з Ховавових синів, Мойсеєвого тестя, і розклав намета свого аж до Елону в Цаананімі, що при Кедеші.
JUDG|4|12|І донесли Сісері, що Барак, син Авіноамів, зійшов на гору Фавор.
JUDG|4|13|І скликав Сісера всі свої колесниці, дев'ятсот залізних колесниць, та ввесь народ, що з ним, з Харошет-Ґаґґоїму до кішонської долини.
JUDG|4|14|І сказала Девора до Барака: Уставай, бо це той день, коли Господь дав Сісеру в твою руку. Ось Господь вийшов перед тобою. І зійшов Барак з гори Фавор, а за ним десять тисяч чоловіка.
JUDG|4|15|І Господь привів у замішання Сісеру, і всі колесниці та ввесь той табір вістрям меча перед Бараком. І зійшов Сісера з колесниці, і побіг пішки.
JUDG|4|16|А Барак гнався за колесницями та за табором аж до Харошет-Ґаґґоїму. І впав увесь табір Сісерин від вістря меча, не позосталось ані одного.
JUDG|4|17|А Сісера втік пішки до намету Яїли, жінки кенеянина Хевера, бо був мир між Явіном, царем Гацору, та між домом кенеянина Хевера.
JUDG|4|18|І вийшла Яїл навпроти Сісери, і сказала до нього: Зайди, пане мій, зайди до мене, не бійся! І він зайшов до неї до намету, і вона накрила його килимом.
JUDG|4|19|І сказав він до неї: Напій мене трохи водою, бо я спрагнений. І відкрила вона молочного бурдюка, і напоїла його, та й накрила його.
JUDG|4|20|І сказав він до неї: Стань при вході намету. І якщо хто ввійде й запитає тебе та скаже: Чи є тут хто? то ти відповіси: Нема.
JUDG|4|21|І взяла Яїл, жінка Хеверона, наметового кілка, і взяла в свою руку молотка, і підійшла тихо до нього, та й всадила того кілка в його скроню, аж у землю. А він спав, змучений, і він помер.
JUDG|4|22|А ось Барак женеться за Сісерою. І вийшла Яїл навпроти нього й сказала йому: Іди, і я покажу тобі того чоловіка, що ти шукаєш. І ввійшов він до неї, а ось Сісера лежить мертвий, а кілок у скроні його!...
JUDG|4|23|Так приборкав Бог того дня Явіна, царя ханаанського, перед Ізраїлевими синами.
JUDG|4|24|А рука Ізраїлевих синів була все тяжча над Явіном, царем ханаанським, аж поки вони вигубили Явіна, царя ханаанського.
JUDG|5|1|І співала Девора й Барак, син Авіноамів, того дня, говорячи:
JUDG|5|2|Що в Ізраїлі закнязювали князі, що народ себе жертвувати став, поблагословіте ви Господа!
JUDG|5|3|Почуйте, царі, уші наставте, князі: я Господеві я буду співати, виспівувати буду Господа, Бога Ізраїля!
JUDG|5|4|Господи, як Ти йшов із Сеїру, як виходив із поля едомського, то тремтіла земля, також капало небо, і хмари дощили водою.
JUDG|5|5|Перед Господнім лицем розпливалися гори, цей Сінай перед Господом, Богом Ізраїля.
JUDG|5|6|За днів Шамґара, сина Анатового, спорожніли дороги, подорожні ж ходили крутими дорогами.
JUDG|5|7|Не стало селянства в Ізраїлі, не стало, аж поки я не повстала, Девора, аж поки я не повстала, мати в Ізраїлі.
JUDG|5|8|Коли вибрав нових він богів, тоді в брамах війна зачалась. Поправді кажу вам, небачений щит був і спис в сорок тисяч Ізраїля!
JUDG|5|9|Серце моє до Ізраїлевих тих начальників, що жертвуються для народу, поблагословіте ви Господа!
JUDG|5|10|Ті, хто їздить на білих ослицях, хто сидить на килимах та дорогою ходить, оповідайте!
JUDG|5|11|Через крик при ділінні здобичі між місцями, де воду беруть, там виспівують правди Господні, правди селянства Його у Ізраїлі. Тоді то зійшов був до брам Господній народ.
JUDG|5|12|Збудися, збудися, Деворо! Збудися, збудися, і пісню співай! Устань, Бараку, і візьми до неволі своїх полонених, сину Авіноамів!
JUDG|5|13|Тоді позосталий зійшов до потужних народу, проти хоробрих Господь був до мене зійшов.
JUDG|5|14|Від Єфрема прийшли були ті, що в Амалику їх корень; Веніямин за тобою, серед народів твоїх; від Махіра зійшли були провідники; а від Завулона оті, хто веде пером писаря.
JUDG|5|15|І князі Іссахарові разом з Деворою, і Іссахар, як Барак, був відпущений пішки в долину. Великі вивідування у Рувимових відділах!
JUDG|5|16|Чого ти усівсь між кошарами, щоб слухати мекання стад? Великі вивідування у Рувимових відділах!
JUDG|5|17|Пробуває Ґілеад на тім боці Йордану, а Дан чому на кораблях буде мешкати він? На березі моря осівся Асир, і при потоках своїх пробуває.
JUDG|5|18|Завулон це народ, що прирік свою душу на смерть, а Нефталим на польових висотах.
JUDG|5|19|Царі прибули, воювали, тоді воювали царі ханаанські в Таанах при воді Меґідда, та здобичі срібла не взяли.
JUDG|5|20|Із неба войовано, зорі з доріг своїх битих воювали з Сісерою.
JUDG|5|21|Кішонський потік позмітав їх, потік стародавній, Кішонський потік. З силою будеш ступати, о душе моя!
JUDG|5|22|Тоді стукотіли копита коня від бігу швидкого, від бігу його скакунів!
JUDG|5|23|Прокляніте Мероза, каже Ангол Господній, проклясти прокляніть його мешканців, бо вони не прийшли Господеві на поміч, Господеві на поміч з хоробрими!
JUDG|5|24|Нехай буде благословенна між жінками Яїл, жінка кенанеянина Хевера, нехай буде благословенна вона між жінками в наметі.
JUDG|5|25|Води він просив подала молока, у царській чаші принесла п'янке молоко.
JUDG|5|26|Ліву руку свою до кілка простягає, а правицю свою до молотка робітничого. І вгатила Сісеру, і розбила вона йому голову, і скроню розбила й пробила йому..
JUDG|5|27|Між ноги її він схилився, упав і лежав, між ноги її він схилився, упав, де схиливсь, там забитий упав.
JUDG|5|28|Через вікно виглядала та голосила Сісерина мати крізь ґрати: Чому колесниця його припізнилась вернутись? Чому припізнились колеса запряжок його?
JUDG|5|29|Мудрі княгині її дають відповідь їй, та й вона сама відповідає собі:
JUDG|5|30|Ось здобич знаходять та ділять вони, бранка, дві бранці на кожного мужа! А здобич із шат кольорових Сісері, здобич із шат кольорових, різнобарвна тканина, на два боки гаптована, жінці на шию.
JUDG|5|31|Нехай отак згинуть усі вороги Твої, Господи! А хто любить Його, той як сонце, що сходить у силі своїй! І Край мав мир сорок літ.
JUDG|6|1|А Ізраїлеві сини чинили зло в очах Господніх, і Господь дав їх у руку мідіянітян на сім літ.
JUDG|6|2|І зміцніла Мідіянова рука над Ізраїлем. Ізраїлеві сини поробили собі зо страху перед мідіянітянами проходи, що в горах, і печери, і твердині.
JUDG|6|3|І бувало, якщо посіяв Ізраїль, то підіймався Мідіян і Амалик та сини Кедему, і йшли на нього.
JUDG|6|4|І вони таборували в них, і нищили врожай землі аж до підходу до Гази. І не лишали вони в Ізраїлі ані поживи, ані штуки дрібної худоби, ані вола, ані осла,
JUDG|6|5|бо вони й їхня худоба та їхні намети ходили, і приходили в такій кількості, як сарана, а їм та їхнім верблюдам не було числа. І вони приходили до Краю, щоб пустошити його.
JUDG|6|6|І через Мідіяна Ізраїль дуже зубожів, і Ізраїлеві сини кликали до Господа.
JUDG|6|7|І сталося, коли Ізраїлеві сини кликали до Господа через Мідіяна,
JUDG|6|8|то Господь послав до Ізраїлевих синів мужа пророка, а він сказав їм: Так сказав Господь, Бог Ізраїлів: Я вивів вас із Єгипту, і випровадив вас із дому рабства.
JUDG|6|9|І Я спас вас з руки Єгипту, і з руки всіх, хто вас тиснув. І Я повиганяв їх перед вами, а їхній Край віддав вам.
JUDG|6|10|І сказав Я до вас: Я Господь, Бог ваш! Не будете боятися аморейських богів, що в їхньому краї сидите ви. Та ви не послухалися Мого голосу!
JUDG|6|11|І прийшов Ангол Господній, і всівся під дубом, що в Офрі, який належить аві-езріянину Йоашеві. А син його Гедеон молотив пшеницю в виноградному чавилі, щоб заховатися перед мідіянітянами.
JUDG|6|12|І явився до нього Ангол Господній, і промовив йому: Господь з тобою, хоробрий мужу!
JUDG|6|13|А Гедеон сказав до нього: О, Пане мій, якщо Господь з нами, то нащо прийшло на нас усе це? І де всі Його чуда, про які оповідали нам наші батьки, говорячи: Ось з Єгипту вивів нас Господь? А тепер Господь покинув нас, і віддав нас у руку Мідіяна.
JUDG|6|14|І обернувся до нього Господь і сказав: Іди з цією своєю силою, і ти спасеш Ізраїля з мідіянської руки. Оце Я послав тебе.
JUDG|6|15|І відказав Йому Гедеон: О, Господи мій, чим я спасу Ізраїля? Ось моя тисяча найнужденніша в Манасії, а я наймолодший у домі батька свого.
JUDG|6|16|І сказав йому Господь: Але Я буду з тобою, і ти поб'єш мідіянітян, як одного чоловіка.
JUDG|6|17|А той до Нього сказав: Якщо знайшов я милість в очах Твоїх, то зроби мені ознаку, що Ти говориш зо мною.
JUDG|6|18|Не відходь же звідси, аж поки я не прийду до Тебе, і не принесу дарунка мого, і не покладу перед лицем Твоїм. А Той відказав: Я буду сидіти аж до твого повернення.
JUDG|6|19|І Гедеон увійшов до хати, і спорядив козеня, і опрісноків з ефи муки, м'ясо поклав до коша, а юшку влив до горщика. І приніс він до Нього під дуб, та й поставив перед Ним.
JUDG|6|20|І сказав до нього Ангол Божий: Візьми це м'ясо й ці опрісноки, та й поклади на оцю скелю, а юшку вилий. І той так зробив.
JUDG|6|21|І витягнув Ангол Господній кінець палиці, що в руці Його, і доторкнувся до м'яса та до опрісноків, і знявся зо скелі огонь, та й поїв те м'ясо та опрісноки, а Ангол Господній зник з його очей.
JUDG|6|22|І побачив Гедеон, що це Ангол Господній. І сказав Гедеон: Ах, Владико, Господи, бож я бачив Господнього Ангола обличчя в обличчя.
JUDG|6|23|І сказав йому Господь: Мир тобі, не бійся, не помреш!
JUDG|6|24|І Гедеон збудував там жертівника для Господа, і назвав ім'я йому: Єгова-Шалом. Він іще є аж до цього дня в Офрі Авіезеровій.
JUDG|6|25|І сталося тієї ночі, і сказав йому Господь: Візьми бичка з волів батька свого, і другого бичка семилітнього, і розбий Ваалового жертівника батька свого, а святе дерево, що при ньому, зрубай.
JUDG|6|26|І збудуєш жертівника Господеві, Богові своєму, на верху цієї твердині, у порядку. І візьмеш другого бичка, і принесеш цілопалення дровами з святого дерева, яке зрубаєш.
JUDG|6|27|І взяв Гедеон десять людей зо своїх рабів, і зробив, як говорив до нього Господь. І сталося, через те, що боявся дому батька свого та людей того міста, щоб робити вдень, то зробив уночі.
JUDG|6|28|І встали люди того міста рано вранці, аж ось жертівник Ваалів розбитий, а святе дерево, що при ньому, порубане, а другого бичка принесено в жертву на збудованому жертівнику.
JUDG|6|29|І говорили вони один одному: Хто зробив оцю річ? І вони вивідували й шукали, та й сказали: Гедеон, син Йоашів, зробив оцю річ.
JUDG|6|30|І сказали люди того міста до Йоаша: Виведи сина свого, і нехай він помре, бо розбив Ваалового жертівника та порубав святе дерево, що при ньому.
JUDG|6|31|І сказав Йоаш до всіх, що стояли при ньому: Чи ви будете обставати за Ваалом? Чи ви допоможете йому? Хто буде обставати за ним, той буде забитий до ранку. Якщо він Бог, то нехай сам заступається за себе, коли той розбив його жертівника.
JUDG|6|32|І він назвав ім'я йому того дня: Єруббаал, говорячи: Нехай змагається з ним Ваал, бо він розбив його жертівника.
JUDG|6|33|А всі мідіяніти й амаликитяни та сини Кедему були зібрані разом, і перейшли Йордан, і таборували в долині Ізреел.
JUDG|6|34|А Дух Господній зійшов на Гедеона, і він засурмив у сурму, і був скликаний Авіезер за ним.
JUDG|6|35|І він послав послів по всьому Манасії, і був скликаний за ним і він. І послав він послів до Асира, і до Завулона, і до Нефталима, і вони вийшли навперейми них.
JUDG|6|36|І сказав Гедеон до Бога: Якщо Ти спасеш Ізраїля моєю рукою, як говорив,
JUDG|6|37|то ось я розстелю на тоці вовняне руно; якщо роса буде на самім руні, а на всій землі сухо, то я буду знати, що Ти спасеш Ізраїля моєю рукою, як говорив!
JUDG|6|38|І сталося так. І встав він рано взавтра, і розстелив руно, і вичавив росу з руна, повне горня води.
JUDG|6|39|І сказав Гедеон до Бога: Нехай не запалиться гнів Твій на мене, нехай я скажу тільки цей раз, нехай но я спробую руном тільки цей раз: нехай буде сухо на самім руні, а на всій землі нехай буде роса.
JUDG|6|40|І Бог зробив так тієї ночі, і було сухо на самім руні, а на всій землі була роса.
JUDG|7|1|І встав рано вранці Єруббаал, це Гедеон, та ввесь народ, що з ним, і таборували над Ен-Хародом. А мідіянітянський табір був із півночі від Ґів'ат-Гамморев долині.
JUDG|7|2|І сказав Господь до Гедеона: Численний той народ, що з тобою, щоб Я дав мідіянітян в його руку, щоб не запишався надо Мною Ізраїль, говорячи: Рука моя спасла мене.
JUDG|7|3|А тепер поклич до ушей люду, говорячи: Хто боїться й тремтить, нехай вернеться й відійде від гори Ґілеад. І вернулося з народу двадцять і дві тисячі, а десять тисяч позосталось.
JUDG|7|4|І сказав Господь до Гедеона: Ще численний цей народ. Зведи їх до води, і Я там переберу його тобі. І буде, як Я скажу тобі: Цей піде з тобою, той піде з тобою, а кожен, що скажу тобі: Цей не піде з тобою, той не піде.
JUDG|7|5|І привів він народ до води. І сказав Господь до Гедеона: Кожен, хто буде хлептати воду язиком своїм, як хлепче пес, поставиш його окремо. А кожен, хто припаде на коліна свої, щоб пити, поставиш його окремо.
JUDG|7|6|І було число тих, що хлептали, носячи рукою своєю до уст своїх, три сотні чоловіка, а вся решта народу припали на коліна свої, щоб пити воду.
JUDG|7|7|І сказав Господь до Гедеона: Трьома сотнями мужів, що хлептали, спасу тебе, і дам мідіянітян у твою руку, а ввесь народ піде кожен на своє місце.
JUDG|7|8|І взяли вони в свою руку поживу народу та свої сурми, а всіх інших ізраїльтян він відпустив, кожного до намету свого, а три сотні мужа затримав. А мідіянітянський табір був під ним у долині.
JUDG|7|9|І сталося тієї ночі, і сказав до нього Господь: Устань, зійди до табору, бо Я дав його в руку твою.
JUDG|7|10|А якщо ти боїшся зійти, зійди ти та Пура, твій слуга, до табору.
JUDG|7|11|І почуєш, що вони говорять, а потім зміцняться твої руки, і ти зійдеш до табору. І зійшов він та Пура, слуга його, до краю озброєних у таборі.
JUDG|7|12|А мідіянітяни й амаликитяни та всі сини Кедему лежали в долині, як сарана, щодо численности. А верблюдам їх нема числа, як пісок на березі моря, щодо численности.
JUDG|7|13|І прийшов Гедеон, аж ось один оповідає другові своєму сон. І він казав: Оце снився мені сон, а ото буханець ячмінного хліба котиться в мідіянітянському таборі. І докотився він аж до намету, та й ударив його, а той упав, і перевернув його догори, і намет той бухнув.
JUDG|7|14|І відповів його друг та й сказав: Це ніщо інше, як меч Гедеона, Йоашового сина, мужа Ізраїльського, Бог дав у його руку мідіянітян та ввесь табір.
JUDG|7|15|І сталося, як Гедеон почув оповідання про той сон та розгадку його, то вклонився, і вернувся до Ізраїлевого табору та й сказав: Уставайте, бо Господь дав у вашу руку мідіянітянський табір!
JUDG|7|16|І поділив він три сотні тих мужів на три відділи, і дав у руку їх усіх сурми, і порожні глеки, та смолоскипи до середини тих глеків.
JUDG|7|17|І сказав він до них: Що будете бачити від мене, то й ви так зробите. А ось я піду до краю табору, і буде, як я зроблю, так зробите й ви.
JUDG|7|18|І засурмлю в сурму я та всі, що зо мною, то засурмите в сурми й ви навколо всього табору, та й скажете: меч за Господа та за Гедеона!
JUDG|7|19|І прийшов Гедеон та сотня мужів, що з ним, до краю табору, на початку середньої сторожі, коли тільки но поставили сторожу. І засурмили вони в сурми, і побили глеки, що в їхніх руках.
JUDG|7|20|І засурмили три відділи в сурми, і поторощили глеки, і тримали рукою своєї лівиці смолоскипа, а рукою своєї правиці сурми, щоб сурмити. І кричали вони: Меч за Господа та за Гедеона!
JUDG|7|21|І стояли кожен на своїм місці навколо табору, а ввесь табір бігав, і вони кричали й утікали.
JUDG|7|22|І засурмили три сотні сурем, а Господь обернув меча одного на одного та на ввесь табір. І табір побіг аж до Бет-Гашшітта до Церери, аж до Сефат-Авел-Мехоли при Таббаті.
JUDG|7|23|І були скликані ізраїльтяни з Нефталиму, і з Асиру, і з усього Манасії, і вони гналися за мідіянітянами.
JUDG|7|24|А по всіх Єфремових горах Гедеон послав послів, говорячи: Зійдіть навперейми мідіянітян, і заступіть їм воду аж до Бет-Бари та Йордан. І скликали всіх Єфремових людей, та й заступили воду аж до Бет-Бари та Йордан.
JUDG|7|25|І вони захопили двох мідіянітянських князів: Орева та Зеева, і вбили Орева в Цур-Ореві, а Зеева вбили в Екев-Зееві. І гналися за мідіянітянами, а голови Орева та Зеева перенесли до Гедеона на той бік Йордану.
JUDG|8|1|І сказали йому мужі Єфремові: Що це за річ зробив ти нам, що не покликав нас, коли йшов воювати з Мідіяном? І вони сильно сперечалися з ним.
JUDG|8|2|І сказав він до них: Що я зробив тепер таке, як ви? Чи не ліпше пізні виноградини Єфремові від авіезерового винобрання?
JUDG|8|3|У вашу руку Бог дав мідіянітянських князів, Орева та Зеева, і що міг я зробити, як ви? Тоді заспокоївся їхній дух проти нього, як він сказав оце слово.
JUDG|8|4|І прийшов Гедеон до Йордану, і перейшов він та три сотні мужів, що з ним, змучені в погоні.
JUDG|8|5|І сказав він до людей Суккоту: Дайте но буханців хліба народові, що за мною, бо вони змучені, а я женуся за Зевахом та Цалмунною, царями мідіянітянськими.
JUDG|8|6|І сказали суккотські князі: Чи рука Зеваха та Цалмунна вже в твоїй руці, щоб давати хліб твоєму війську?
JUDG|8|7|І сказав Гедеон: Тому то, коли Господь дасть у мою руку Зеваха та Цалмунну, то я буду молотити ваше тіло пустинними тернями та колючками!
JUDG|8|8|І пішов він звідти до Пенуїлу, і говорив до них те саме. А люди Пенуїлу відповіли йому, як відповіли люди Суккоту.
JUDG|8|9|І він сказав також до людей Пенуїлу, говорячи: Коли я вертатимусь у мирі, розіб'ю оцю вежу.
JUDG|8|10|А Зевах та Цалмунна були в Каркорі, і з ними їхні табори, близько п'ятнадцяти тисяч, усі позосталі з усього табору синів Кедему. А тих, що впали, було сто й двадцять тисяч чоловіка, що витягали меча.
JUDG|8|11|А Гедеон пішов дорогою Шехуне-Боголіму зо сходу до Коваху й Йоґбеги. І розбив він табора, коли табір був безпечний.
JUDG|8|12|І втікали Зевах та Цалмунна, а він гнався за ними. І він схопив обох мідіянітянських царів, Зеваха та Цалмунну, а на ввесь табір нагнав жаху.
JUDG|8|13|І вернувся Гедеон, син Йоашів, із війни з Маале-Гахересу.
JUDG|8|14|І захопив він юнака з людей Суккоту, та й запитався його. І той написав йому ймення князів Суккоту та старших його, сімдесят і сім чоловіка.
JUDG|8|15|І прийшов він до людей Суккоту та й сказав їм: Ось Зевах та Цалмунна, що ви ображали мене, говорячи: Чи рука Зеваха та Цалмунни тепер у твоїй руці, що дамо хліба твоїм змученим людям?
JUDG|8|16|І схопив він старших того міста, і пустинне терня та колючки, і побив ними суккотських людей.
JUDG|8|17|А пенуїльську вежу розбив, і позабивав людей того міста.
JUDG|8|18|І сказав він до Зеваха та до Цалмунни: Які ті люди, що ви повбивали на Фаворі? А ті сказали: Як ти, так вони одне, мають вигляд царських синів.
JUDG|8|19|А він сказав: То брати мої, сини моєї матері. Як живий Господь, коли б ви були позоставили їх при житті, не повбивав би я вас!
JUDG|8|20|І сказав він до Єтера, свого первенця: Устань, забий їх! Та той юнак не витяг свого меча, бо боявся, бо він був ще малий.
JUDG|8|21|І сказав Зевах та Цалмунна: Устань ти, і кинься на нас, бо по чоловікові сила його. І встав Гедеон, і вбив Зеваха та Цалмунну, і забрав оздобні місяці, що були на шиях їхніх верблюдів.
JUDG|8|22|І сказали Ізраїлеві мужі до Гедеона: Пануй над нами і ти, і син твій, і син твого сина, бо ти спас нас від руки Мідіяна.
JUDG|8|23|І сказав до них Гедеон: Не буду панувати над вами я, і не буде панувати над вами син мій, Господь пануватиме над вами.
JUDG|8|24|І сказав до них Гедеон: Попрошу від вас прохання, і дайте мені кожен носову сережку зо своєї здобичі, бо в них, мідіянітян, були золоті носові сережки, бо ізмаїльтяни вони.
JUDG|8|25|І сказали вони: Дати дамо. І розтягнули одежу, і кидали туди кожен носову сережку зо своєї здобичі.
JUDG|8|26|І була вага золотих носових сережок, що він просив, тисяча й сімсот шеклів золота, крім оздобних місяців, і сережок, і пурпурових шат, що були на мідіянітянських царях, і окрім нашийників, що на шиях їхніх верблюдів.
JUDG|8|27|А Гедеон зробив із того ефода, і поставив його у своєму місті, в Офрі. І за ним чинив там перелюб увесь Ізраїль, і це стало пасткою для Гедеона та для дому його.
JUDG|8|28|І був упокорений Мідіян перед Ізраїлевими синами, і він більш не підіймав своєї голови. І Край мав мир сорок літ за Гедеонових днів.
JUDG|8|29|І пішов Еруббаал, син Йоашів, та й осівся в своїм домі.
JUDG|8|30|А в Гедеона було сімдесят синів, що походили зо стегон його, бо він мав багато жінок.
JUDG|8|31|А наложниця його, що в Сихемі, породила йому сина й вона, а він назвав ім'я йому: Авімелех.
JUDG|8|32|І помер Гедеон, син Йоашів, у добрій сивизні, і був похований у гробі Йоаша, батька свого, в Офрі авіезеровій.
JUDG|8|33|І сталося, як помер Гедеон, то Ізраїлеві сини знову чинили перелюб із Ваалами, і поставили собі Ваал-Берита за бога.
JUDG|8|34|І Ізраїлеві сини не пам'ятали Господа, Бога свого, що спасав їх від руки всіх їхніх навколишніх ворогів.
JUDG|8|35|І не зробили вони милости з домом Єруббаала-Гедеона такої, як усе те добро, яке він зробив для Ізраїля.
JUDG|9|1|І пішов Авімелех, син Єруббаалів, до Сихему, до братів своєї матері, і говорив до них та до всього роду батьківського дому своєї матері, кажучи:
JUDG|9|2|Говоріть голосно до всіх сихемських господарів: Що ліпше для вас: чи панування над вами семидесяти мужів, усіх Єруббаалових синів, чи панування над вами мужа одного? І пам'ятайте, що я кість ваша та тіло ваше.
JUDG|9|3|І говорили брати його матері про нього голосно до сихемських господарів усі ті слова, і їхнє серце схилилося до Авімелеха, бо вони сказали: Він наш брат.
JUDG|9|4|І дали йому сімдесят шеклів срібла з дому Баал-Беріта, а Авімелех найняв за них пустих та легковажних людей, і вони пішли за ним.
JUDG|9|5|А він прийшов до дому свого батька в Офру, і повбивав своїх братів, синів Єруббаалових, сімдесят чоловіка на однім камені. І позостався тільки Йотам, син Єруббаалів, наймолодший, бо сховався.
JUDG|9|6|І були зібрані всі сихемські господарі та ввесь Бет-Мілло, і вони пішли та й настановили Авімелеха за царя при Елон-Муццаві, що в Сихемі.
JUDG|9|7|І повідомили про це Йотама, і він пішов, і став на верхів'ї гори Ґаріззім, і підвищив свій голос, і закликав та й сказав їм: Почуйте мене, сихемські господарі, і хай почує вас Бог!
JUDG|9|8|Пішли були раз дерева, щоб помазати царя над собою, і сказали вони до оливки: Царюй ти над нами!
JUDG|9|9|А оливка сказала до них: Чи я загубила свій товщ, що Бога й людей ним шанують, і сторожити піду над деревами?
JUDG|9|10|І сказали дерева до фіґи: Іди ти, та й над нами царюй!
JUDG|9|11|І сказала їм фіґа: Чи я загубила свої солодощі та свій добрий врожай, і сторожити піду над деревами?
JUDG|9|12|І дерева промовили до винограду: Іди ти, та й над нами царюй!
JUDG|9|13|І промовив до них виноград: Чи я загубив свого сока, що Бога й людей веселити, і сторожити піду над деревами?
JUDG|9|14|Тоді всі дерева сказали тернині: Іди ти, та й над нами царюй!
JUDG|9|15|А тернина сказала деревам: якщо справді мене на царя над собою помазуєте, підійдіть, поховайтеся в тіні моїй! А як ні, то ось вийде огонь із тернини, та кедри ливанські поїсть!
JUDG|9|16|А тепер, якщо направду й у невинності зробили ви, що настановили Авімелеха царем, і якщо ви добре зробили з Єруббаалом та з домом його, і якщо ви зробили йому за заслугою рук його,
JUDG|9|17|бо мій батько воював за вас, і кинув був життя своє на небезпеку, і врятував вас із руки Мідіяна,
JUDG|9|18|а ви сьогодні повстали на дім батька мого, та й повбивали синів його, сімдесят люда, на одному камені, і настановили царем Авімелеха, сина його невільниці, над сихемськими господарями, бо він брат ваш,
JUDG|9|19|і якщо в правді й невинності зробили ви з Єруббаалом та з домом його цього дня, то радійте Авімелехом, і нехай і він радіє вами!
JUDG|9|20|А як ні, вийде огонь з Авімелеха, та й поїсть господарів Сихему й Бет-Мілло, і вийде огонь із господарів Сихему й з Бет-Мілло, та й з'їсть Авімелеха.
JUDG|9|21|І втік Йотам і збіг, і пішов до Бееру, і сидів там перед братом своїм.
JUDG|9|22|І володів Авімелех над Ізраїлем три роки.
JUDG|9|23|І послав Господь злого духа між Авімелехом та між сихемськими господарями, і зрадили сихемські господарі Авімелеха,
JUDG|9|24|щоб прийшла кривда семидесяти Єруббаалових синів, а їхня кров спала на Авімелеха, їхнього брата, що їх повбивав, та на сихемських господарів, що зміцнили його руки забити братів своїх.
JUDG|9|25|І сихемські господарі поставили на верхів'ях гір чатівників на нього, і вони грабували все, що приходило до них на дорозі. І сказано про це Авімелеху.
JUDG|9|26|І прийшов Ґаал, Еведів син, та брати його, і вони прийшли до Сихему, і довірилися йому сихемські господарі.
JUDG|9|27|І виходили вони в поле, і збирали виноград свій, і вичавлювали, і робили празник. І входили вони до дому свого бога, і їли й пили та проклинали Авімелеха.
JUDG|9|28|І говорив Ґаал, син Еведів: Хто Авімелех і хто Сихем, що будемо служити йому? Чи ж він не син Єруббаалів, а Зевул начальник його? Служіть людям Гемора, батька Сихема, а чому ми будемо служити йому?
JUDG|9|29|А хто дав би цього народа в мою руку, то я прогнав би Авімелеха. І він скаже до Авімелеха: Помнож своє військо, та й вийди!
JUDG|9|30|І почув Зевул, голова міста, слова Ґаала, сина Еведового, і запалився його гнів.
JUDG|9|31|І послав він послів до Авімелеха з хитрістю, говорячи: Ось Ґаал, син Еведів, та брати його приходять до Сихему, і ось вони підбурюють місто проти тебе.
JUDG|9|32|А тепер устань уночі ти та той народ, що з тобою, і чатуй на полі.
JUDG|9|33|І буде, встанеш рано вранці, як сходитиме сонце, і нападеш на місто. І ось, він та народ той, що з ним, вийдуть до тебе, а ти зробиш йому, як знайде потрібним рука твоя.
JUDG|9|34|І встав уночі Авімелех та ввесь народ, що з ним, та й чатували над Сихемом чотири відділи.
JUDG|9|35|І вийшов Ґаал, син Еведів, і став при вході міської брами. І встав Авімелех та народ, що з ним, із засідки.
JUDG|9|36|А Ґаал побачив той народ, та й сказав до Зевула: Ось народ сходить із верхів гір. І сказав до нього Зевул: Ти бачиш гірську тінь, немов людей!
JUDG|9|37|А Ґаал далі говорив та казав: Ось народ сходить з верхів'я, а один відділ приходить із дороги Елон-Меоненіму.
JUDG|9|38|І сказав до нього Зевул: Де тоді уста твої, що говорили: Хто Авімелех, що ми будем служити йому? А оце той народ, що ти погорджував ним. Виходь же тепер, та й воюй з ним!
JUDG|9|39|І вийшов Ґаал перед сихемськими господарями, та й воював з Авімелехом.
JUDG|9|40|І Авімелех погнав його, і він побіг перед ним. І нападало багато трупів аж до входу до брами.
JUDG|9|41|І осівся Авімелех в Арумі, а Зевул вигнав Ґаала та братів його, щоб не сиділи в Сихемі.
JUDG|9|42|І сталося другого дня, і вийшов народ на поле, а Авімелеху донесли про це.
JUDG|9|43|І взяв він людей, і поділив їх на три відділи, та й чатував на полі. І побачив він, аж ось народ виходить із міста, і встав він на них, та й побив їх.
JUDG|9|44|А Авімелех та відділи, що з ним, напали й стали при вході міської брами, а два відділи напали на все, що в полі, та й повбивали їх.
JUDG|9|45|І Авімелех воював із містом цілий той день, та й здобув місто, а народ, що був у ньому, позабивав. І зруйнував він те місто, та й обсіяв його сіллю.
JUDG|9|46|І почули про це всі, хто був у сихемській башті, і ввійшли до твердині, до дому бога Беріта.
JUDG|9|47|І було донесено Авімелехові, що зібралися всі господарі сихемської башти.
JUDG|9|48|І вийшов Авімелех на гору Цалмон, він та ввесь народ, що з ним. І взяв Авімелех сокири в свою руку, та й настинав галуззя з дерева, і позносив його, і поклав на своє плече. І сказав він до народу, що з ним: Що ви бачили, що зробив я, поспішно зробіть, як я.
JUDG|9|49|І настинав також увесь народ кожен галуззя собі, і пішли за Авімелехом, і поскладали над печерою, та й підпалили над ними ту печеру огнем. І повмирали всі люди сихемської вежі, близько тисячі чоловіків та жінок.
JUDG|9|50|І пішов Авімелех до Тевецу, і таборував при Тевеці, та й здобув його.
JUDG|9|51|А в середині міста була міцна башта, і повтікали туди всі чоловіки й жінки та всі господарі міста, і замкнули за собою, та й вийшли на дах тієї башти.
JUDG|9|52|І прийшов Авімелех аж до башти, та й воював із нею. І підійшов він аж до входу башти, щоб спалити її огнем.
JUDG|9|53|Тоді одна жінка кинула горішнього каменя від жорен на Авімелехову голову, та й розторощила йому черепа.
JUDG|9|54|І він зараз кликнув до юнака, свого зброєноші, та й сказав йому: Витягни свого меча, та й забий мене, щоб не сказали про мене: Його жінка забила! І його юнак проколов його, і він помер.
JUDG|9|55|І побачили ізраїльтяни, що Авімелех помер, та й порозходилися кожен на своє місце.
JUDG|9|56|І Бог віддав Авімелехові зло, яке він зробив був своєму батькові, що повбивав сімдесят братів своїх.
JUDG|9|57|А все зло сихемських людей Бог повернув на їхню голову, і прийшло на них прокляття Йотама, Єруббаалового сина.
JUDG|10|1|І став по Авімелехові на спасіння Ізраїля Тола, син Пуї, сина Додового, муж Іссахарів. І він сидів у Шамірі в Єфремових горах.
JUDG|10|2|І судив він Ізраїля двадцять і три роки, та й помер, і був похований в Шамірі.
JUDG|10|3|І став по ньому Яір ґілеадеянин, і судив Ізраїля двадцять і два роки.
JUDG|10|4|І було в нього тридцять синів, що їздили на тридцяти молодих ослах, а в них тридцять міст, їх кличуть аж до цього дня: Яірові села, що в ґілеадському краї.
JUDG|10|5|І помер Яір, і був похований в Камоні.
JUDG|10|6|А Ізраїлеві сини й далі чинили зло в Господніх очах, і служили Ваалам та Астартам, і богам арамським, і богам сидонським, і богам моавським, і богам аммонських синів, і богам филистимським. І покинули вони Господа, і не служили Йому.
JUDG|10|7|І запалився Господній гнів на Ізраїля, і Він передав їх в руку филистимлян та в руку синів Аммонових.
JUDG|10|8|І вони били й мучили Ізраїлевих синів від того року, і гнобили вісімнадцять років усіх Ізраїлевих синів, що по той бік Йордану в аморейському краї, що в Ґілеаді.
JUDG|10|9|І перейшли Аммонові сини Йордан, щоб воювати також з Юдою й з Веніямином та з Єфремовим домом. І Ізраїлеві було дуже тісно!
JUDG|10|10|І кликали Ізраїлеві сини до Господа, говорячи: Згрішили ми Тобі, бо ми покинули свого Бога, і служили Ваалам.
JUDG|10|11|І сказав Господь до Ізраїлевих синів: Чи ж не спас Я вас від Єгипту, і від амореянина, і від Аммонових синів, і від филистимлян?
JUDG|10|12|А сидоняни, і Амалик, і Маон гнобили вас, і ви кликали до Мене, і Я спас вас від їхньої руки.
JUDG|10|13|А ви полишили Мене, і служили іншим богам, тому більше не спасатиму вас.
JUDG|10|14|Ідіть, і кличте до тих богів, що ви вибрали їх, вони спасуть вас у часі вашого утиску.
JUDG|10|15|І сказали Ізраїлеві сини до Господа: Згрішили ми! Зроби Ти нам усе, як добре в очах Твоїх. Тільки спаси нас цього дня!
JUDG|10|16|І повикидали вони з-поміж себе чужих богів, та й служили Господеві. І знетерпеливилась душа Його через Ізраїлеве страждання.
JUDG|10|17|А Аммонові сини були скликані, та й таборували в Ґілеаді. І були зібрані Ізраїлеві сини, та й таборували в Міцпі.
JUDG|10|18|І сказали той народ та ґілеадські князі, один до одного: Хто той чоловік, що зачне воювати з Аммоновими синами? Він стане головою для всіх ґілеадських мешканців.
JUDG|11|1|А ґілеадянин Їфтах був хоробрий вояк. А він був син блудливої жінки, і з нею Ґілеад породив Їфтаха.
JUDG|11|2|І породила Ґілеадова жінка йому синів. І повиростали сини тієї жінки, та й вигнали Їфтаха, і сказали йому: Не будеш володіти в домі нашого батька, бо ти син іншої жінки!
JUDG|11|3|І втік Їфтах перед своїми братами, і осівся в краї Тов. І зібралися до Їфтаха гулящі люди, та й виходили з ним.
JUDG|11|4|І сталося по часі, і воювали Аммонові сини з Ізраїлем.
JUDG|11|5|І сталося, як воювали Аммонові сини з Ізраїлем, то пішли ґілеадські старші, щоб забрати Їфтаха з краю Тов.
JUDG|11|6|І сказали вони до Їфтаха: Іди ж, і будеш нам провідником, і будемо воювати з Аммоновими синами.
JUDG|11|7|І сказав Їфтах до ґілеадських старших: Чи ж не ви зненавидили мене, і вигнали мене з дому мого батька? І чого ви прийшли до мене тепер, коли ви в біді?
JUDG|11|8|І сказали ґілеадські старші до Їфтаха: Зате ми тепер вернулися до тебе! І ти піди з нами, і будемо воювати з Аммоновими синами, і станеш нам головою для всіх мешканців ґілеадських.
JUDG|11|9|І сказав Їфтах до ґілеадських старших: Якщо ви мене вернете воювати з Аммоновими синами, і Господь дасть їх, щоб були побиті передо мною, то чи я стану вам головою?
JUDG|11|10|І сказали ґілеадські старші до Їфтаха: Нехай Господь буде свідком поміж нами, що так, як слово твоє, так зробимо.
JUDG|11|11|І пішов Їфтах з ґілеадськими старшими, і народ настановив його собі за голову та провідника, а Їфтах промовляв усі свої слова перед Господнім лицем у Міцпі.
JUDG|11|12|І послав Їфтах послів до царів Аммонових синів, говорячи: Що тобі до мене, що ти прийшов до мене воювати з моїм краєм?
JUDG|11|13|І сказав цар Аммонових синів до Їфтахових послів: Бо Ізраїль забрав мій край, коли він виходив з Єгипту, від Арнону й аж до Яббоку та аж до Йордану. А тепер верни ж їх у мирі.
JUDG|11|14|А Їфтах ще послав послів до царя Аммонових синів,
JUDG|11|15|і сказав йому: Так сказав Їфтах: Не взяв Ізраїль краю Моавого та краю Аммонових синів,
JUDG|11|16|бо коли йшли вони з Єгипту, то Ізраїль ішов по пустині аж до Червоного моря, і прийшов до Кадешу.
JUDG|11|17|І послав Ізраїль послів до едомського царя, говорячи: Нехай я перейду твоїм краєм, та не послухав едомський цар. І послав він також до царя моавського, та й той не хотів. І осівся Ізраїль у Кадешу.
JUDG|11|18|І пішов він пустинею, і обійшов край едомський та край моавський, і прийшов зо сходу сонця до моавського краю, та й таборували по тім боці Арнону, а в моавські границі не входили, бо Арнон границя Моава.
JUDG|11|19|І послав Ізраїль послів до Сихона, царя аморейського, царя хешбонського, і сказав йому Ізраїль: Нехай ми перейдемо твоїм краєм аж до місця свого.
JUDG|11|20|І не вірив Сихон Ізраїлеві, щоб він мирно перейшов його границями. І зібрав Сихон увесь народ свій, та й таборували в Йохці, і воювали з Ізраїлем.
JUDG|11|21|І дав Господь, Бог Ізраїля, Сихона та ввесь народ його в Ізраїлеву руку, вони побили їх. І посів Ізраїль увесь край амореянина, мешканця того краю.
JUDG|11|22|І вони посіли всю аморейську країну від Арнону й аж до Яббоку, і від пустині та аж до Йордану.
JUDG|11|23|А тепер Господь, Бог Ізраїлів, вигнав Амореянина перед народом Своїм, Ізраїлем, а ти посядеш його?
JUDG|11|24|Отож, що дасть тобі на насліддя Кемош, бог твій, те ти посядеш, а все, де вигнав Господь, Бог наш, перед нами, те ми посядемо.
JUDG|11|25|А тепер чи справді ти ліпший від Балака, Ціппорового сина, царя моавського? Чи сваритися сварився він з Ізраїлем? Чи воювати воював із ними?
JUDG|11|26|Коли Ізраїль сидів у Хешбоні та в підлеглих містах його, і в Ар'орі та в підлеглих містах його, і по всіх містах, що над Арноном, три сотні літ, то чому не відібрали ви їх за той час?
JUDG|11|27|А тобі я не згрішив, а ти робиш зо мною зло, щоб воювати зо мною. Нехай розсудить Господь, що судить сьогодні між Ізраїлевими синами та між синами Аммоновими.
JUDG|11|28|Та цар Аммонових синів не послухався слів Їфтаха, що до нього посилав.
JUDG|11|29|І Дух Господній перебував на Їфтахові, і він перейшов Ґілеад та Манасію, і перейшов ґілеадську Міцпе, а з ґілеадської Міцпе перейшов до Аммонових синів.
JUDG|11|30|І обіцяв Їфтах обітницю Господеві й сказав: Якщо справді даси Ти Аммонових синів у мою руку,
JUDG|11|31|то станеться, виходячий, що вийде з дверей мого дому навпроти мене, коли я вертатимусь з миром від Аммонових синів, то буде він для Господа, і я принесу його в цілопалення.
JUDG|11|32|І прийшов Їфтах до Аммонових синів воювати з ними, а Господь дав їх у його руку.
JUDG|11|33|І він побив їх дуже великою поразкою від Ароеру й аж туди, де йти до Мінніту, двадцять міст, і аж до Авел-Кераміму. І впокорилися Аммонові сини перед синами Ізраїлевими.
JUDG|11|34|І прийшов Їфтах до Міцпи до свого дому, аж ось виходить навпроти нього дочка його з бубнами та з танцями! А вона була в нього тільки одна, не було в нього, окрім неї, ані сина, ані дочки.
JUDG|11|35|І сталося, як він побачив її, то роздер одежу свою та й сказав: Ах, дочко моя! Ти справді повалила мене, і ти стала однією з тих, що нещасливлять мене. Бо я дав Господеві обіта, і не можу відмовитися від нього.
JUDG|11|36|А вона відказала йому: Батьку мій, ти дав обітницю Господеві, зроби мені, як вийшло з твоїх уст, коли Господь зробив тобі пімсту на твоїх ворогів, на Аммонових синів.
JUDG|11|37|І сказала вона до свого батька: Нехай буде мені зроблена оця річ: відпусти мене на два місяці, і нехай я піду й зійду на гору, і нехай оплачу дівування своє я та приятельки мої.
JUDG|11|38|А він сказав: Іди! І послав її на два місяці. І пішла вона та її приятельки, і оплакувала дівування своє.
JUDG|11|39|І сталося в кінці двох місяців, і вернулася вона до батька свого, а він учинив над нею свою обітницю, яку обіцяв був, і вона не пізнала мужа. І сталося це звичаєм в Ізраїлі:
JUDG|11|40|рік-річно ходять Ізраїлеві дочки плакати за дочкою ґілеадянина Їфтаха, чотири дні в році.
JUDG|12|1|І були скликані Єфремові люди, і перейшли на північ та й сказали до Їфтаха: Чому перейшов ти Йордан, щоб воювати з Аммоновими синами, а нас не покликав піти з собою? Ми спалимо огнем твій дім із тобою.
JUDG|12|2|І сказав їм Їфтах: Велику боротьбу мав я та народ мій з Аммоновими синами. І кликав я вас, та ви не спасли мене з його руки.
JUDG|12|3|І коли я побачив, що ви не спасете, то поклав я душу свою на небезпеку, і перейшов Йордан до Аммонових синів, а Господь дав їх у мою руку. І чого прийшли ви до мене цього дня, щоб воювати зо мною?
JUDG|12|4|І зібрав Їфтах усіх ґілеадських людей, та й воював з Єфремом. І побили ґілеадські люди Єфрема, бо ті сказали: Ви Єфремові втікачі, Ґілеад поміж Єфремом та поміж Манасією.
JUDG|12|5|І зайняв Ґілеад йорданські переходи до Єфрема. І сталося, коли говорили Єфремові втікачі: Нехай я перейду, то ґілеадські люди йому говорили: Чи ти єфремівець? Той казав: Ні.
JUDG|12|6|І казали йому: Скажи но шібболет. А той казав: Сібболет, бо не міг вимовити так. І хапали його, і різали при йорданськім переході. І впало того часу в Єфрема сорок і дві тисячі.
JUDG|12|7|І судив Їфтах Ізраїля шість років. І помер ґілеадянин Їфтах, і був похований у місті Ґілеаді.
JUDG|12|8|А по ньому Ізраїля судив Івцан з Віфлеєму.
JUDG|12|9|І було в нього тридцять синів, а тридцять дочок він відпустив заміж назовні, і тридцять дочок впровадив для синів своїх з-назовні. І судив він Ізраїля сім літ.
JUDG|12|10|І помер Івцан і був похований в Віфлеємі.
JUDG|12|11|А по ньому Ізраїля судив завулонівець Елон, і судив Ізраїля десять літ.
JUDG|12|12|І помер завулонівець Елон, і був похований в Айялоні, у Завулоновім краї.
JUDG|12|13|А по ньому Ізраїля судив Авдон, син Гіллела, пір'атонянин.
JUDG|12|14|І було в нього сорок синів та тридцять онуків, що їздили на семидесяти молодих ослах. І судив він Ізраїля вісім літ.
JUDG|12|15|І помер Авдон, син Гіллела, пір'атонянин, і був похований в Єфремовім краї, на горі амаликеянина.
JUDG|13|1|А Ізраїлеві сини й далі робили зло в Господніх очах. І Господь віддав їх у руку филистимлян на сорок літ.
JUDG|13|2|І був один чоловік з Цар'ї, данівець з роду, а ім'я йому Маноах. А жінка його була неплідна, і не родила.
JUDG|13|3|І явився Ангол Господній до тієї жінки, та й промовив до неї: Ось ти неплідна, і не роджала, але ти зачнеш і породиш сина.
JUDG|13|4|А тепер стережись, і не пий вина та п'янкого напою, і не їж нічого нечистого,
JUDG|13|5|бо ось ти зачнеш, і сина породиш, і бритва не торкнеться його голови, бо дитя те буде Божим назореєм від утроби, і він зачне спасати Ізраїля з руки филистимлян.
JUDG|13|6|І прийшла та жінка, та й сказала до чоловіка свого, говорячи: Божий чоловік приходив до мене, а вигляд його як вигляд Божого Ангола, дуже грізний. І я не питала його, звідки він, а ймення свого він мені не сказав.
JUDG|13|7|І сказав він мені: Ось ти зачнеш, і породиш сина, а тепер не пий вина та п'янкого напою, і не їж жодної нечистости, бо дитя те буде Божим назореєм від утроби аж до дня смерти своєї.
JUDG|13|8|І благав Маноах Господа, та й сказав: О Господи, Божий чоловік, що його посилав Ти, нехай прийде ще до нас, і нехай нас навчить, що ми зробимо для дитини, що народиться.
JUDG|13|9|І вислухав Бог цей Маноахів голос, і прийшов Божий Ангол ще до тієї жінки. А вона сиділа на полі, і Маноаха, чоловіка її, не було з нею.
JUDG|13|10|І поспішила та жінка, і побігла та й оповіла чоловікові своєму, і сказала до нього: Ось з'явився мені той чоловік, що приходив був того дня до мене.
JUDG|13|11|І встав, і пішов Маноах за своєю жінкою, і прийшов до того чоловіка, та й сказав йому: Чи ти той чоловік, що говорив до цієї жінки? А той сказав: Я.
JUDG|13|12|І сказав Маноах: Тепер нехай сповниться слово твоє. Та як нам виховувати ту дитину, і що чинити з нею?
JUDG|13|13|І сказав Ангол Господній до Маноаха: Усього, що сказав я жінці, нехай вона стережеться.
JUDG|13|14|Усього, що виходить із виноградного куща, не буде вона їсти, а вина та напою п'янкого нехай не п'є, і нічого нечистого нехай не їсть. Нехай додержує всього, що я наказав.
JUDG|13|15|І сказав Маноах до Ангола Господнього: Нехай ми задержимо тебе, і приготовимо для тебе козля.
JUDG|13|16|І сказав Ангол Господній до Маноаха: Якщо ти задержиш мене, я не буду їсти твого хліба. А якщо приготуєш цілопалення для Господа принесеш його. Бо Маноах не знав, що це Ангол Господній.
JUDG|13|17|І сказав Маноах до Господнього Ангола: Яке ім'я твоє? Коли сповниться твоє слово, то ми вшануємо тебе.
JUDG|13|18|І сказав йому Ангол Господній: Чому ти питаєшся про моє ім'я? Воно дивне.
JUDG|13|19|І взяв Маноах козля та жертву хлібну, і на скелі приніс Господеві. І Він учинив чудо, а Маноах та його жінка бачили те.
JUDG|13|20|І сталося, коли полум'я підіймалося з-над жертівника до неба, то Ангол Господній вознісся в полум'ї жертівника. А Маноах та жінка його бачили це, та й попадали обличчям своїм на землю.
JUDG|13|21|І Ангол Господній більш уже не появлявся до Маноаха та до жінки його. Тоді Маноах пізнав, що це Ангол Господній.
JUDG|13|22|І сказав Маноах до своєї жінки: Ми справді помремо, бо ми бачили Бога.
JUDG|13|23|І сказала йому жінка його: Коли б Господь хотів був повбивати нас, не взяв би з нашої руки цілопалення та хлібної жертви, і не дав би нам побачити всього цього, і не об'явив би нам цього часу речі, як це.
JUDG|13|24|І породила та жінка сина, і назвала ім'я йому: Самсон. І виростав той хлопець, і Господь благословляв його.
JUDG|13|25|А Дух Господній почав діяти в ньому в Дановім таборі між Цор'а та між Ештаолом.
JUDG|14|1|І зійшов Самсон до Тімни, і побачив у Тімні жінку з филистимських дочок.
JUDG|14|2|І пішов він, і розповів своєму батькові та своїй матері, та й сказав: Я нагледів у Тімні жінку з филистимських дочок, а тепер візьміть її мені за жінку.
JUDG|14|3|І сказав йому батько його та мати його: Чи ж нема жінки серед дочок братів твоїх та серед усього мого народу, що ти йдеш узяти жінку з необрізаних филистимлян? І сказав Самсон до свого батька: Візьми її мені, бо вона люба очам моїм.
JUDG|14|4|А батько його та мати його не знали, що це від Господа, бо він шукав зачіпки з филистимлянами. А того часу филистимляни панували над Ізраїлем.
JUDG|14|5|І зійшов Самсон і батько його та мати його до Тімни, і прийшли аж до тімненських виноградників, аж ось навпроти нього ричить левчук.
JUDG|14|6|І зійшов на нього Дух Господній, і він розірвав того левчука, як розривають ягня, а в руці його не було нічого. І він не сказав своєму батькові та своїй матері, що зробив.
JUDG|14|7|І він зійшов, і говорив до тієї жінки, і вона стала улюблена в Самсонових очах.
JUDG|14|8|А по часі він вертався забрати її, і звернув із дороги побачити падло лева, аж ось рій бджіл у тілі того лева та мед.
JUDG|14|9|І він вишкріб його на свою долоню, і пішов, і їв та й їв. І він пішов до батька свого й до матері своєї, та й дав їм, і вони їли. І він не сказав їм, що той мед він зішкріб із тіла лева.
JUDG|14|10|І зійшов його батько до тієї жінки, а Самсон справив там прийняття, бо так роблять юнаки.
JUDG|14|11|І сталося, коли вони побачили його, то взяли тридцятеро дружків, і були з ним.
JUDG|14|12|І сказав їм Самсон: Нехай но я загадаю вам загадку. Якщо справді розгадаєте її мені за сім день прийняття, і відгадаєте, то я дам тридцять лляних сорочок та тридцять змін одежі.
JUDG|14|13|А якщо не зможете розгадати мені, то ви мені дасте тридцять лляних сорочок та тридцять змін одежі. І вони сказали йому: Загадуй загадку свою, а ми послухаємо її.
JUDG|14|14|І він сказав їм: З їдячого вийшло їстивне, а з сильного вийшло солодке. І не могли вони розгадати за три дні.
JUDG|14|15|І сталося сьомого дня, і сказали вони до Самсонової жінки: Намов свого чоловіка, і нехай він розгадає нам ту загадку, щоб ми не спалили огнем тебе та дім твого батька. Чи ви нас покликали, щоб посісти маєток наш, чи ні?
JUDG|14|16|І плакала Самсонова жінка при ньому сім день і казала: Ти певне ненавидиш мене й не любиш мене. Ти загадав загадку синам мого народу, а мені не розгадав. А він їй сказав: Таж батькові своєму та матері своїй не розгадав я, а розгадаю тобі?
JUDG|14|17|А вона плакала при ньому сім день, коли в них було прийняття. І сталося сьомого дня, і він розгадав їй, бо вона докучала йому. А вона розгадала ту загадку синам свого народу.
JUDG|14|18|І сказали йому люди того міста сьомого дня, поки зайшло сонце: Що солодше від меду, і що сильніше від лева? А він їм відказав: Якби ви не орали моєю телицею, то ви загадки не відгадали б моєї.
JUDG|14|19|І зійшов на нього Дух Господній, і він пішов до Ашкелону, та й побив з них тридцятеро чоловіка, і пороздягав їх, і віддав ті зміни одежі тим, що розгадали загадку. І запалився гнів його, і він пішов до дому батька свого.
JUDG|14|20|А Самсонова жінка досталася дружкові його, що приятелював із ним.
JUDG|15|1|А по часі сталося в днях жнив пшениці, і відвідав Самсон з козлям свою жінку та й сказав: Нехай увійду я до моєї жінки, до кімнати. Та батько її не дав йому ввійти.
JUDG|15|2|І сказав її батько: Я дійсно подумав був, що ти справді зненавидів її, а тому я дав її твоєму дружкові. Чи молодша сестра її не ліпша від неї? Нехай же вона буде тобі замість неї.
JUDG|15|3|І сказав їм Самсон: Цього разу я не буду винний перед филистимлянами, коли я зроблю їм зло.
JUDG|15|4|І пішов Самсон, та й зловив три сотні лисиць. І взяв він смолоскипи, і обернув хвоста до хвоста, і прив'язав одного смолоскипа всередині поміж два хвости.
JUDG|15|5|І запалив він огонь у тих смолоскипах, і пустив лисиць в филистимські жита. І попалив він стирти та жита, і оливкові сади.
JUDG|15|6|І сказали филистимляни: Хто це зробив? А їм відказали: Самсон, зять тімнеянина, бо він забрав його жінку й віддав її дружкові його. І пішли филистимляни, та й спалили огнем її та батька її.
JUDG|15|7|І сказав їм Самсон: Хоч ви й зробили так, як це, та проте я конче пімщуся на вас, і аж тоді перестану.
JUDG|15|8|І він сильно побив їх дошкульною поразкою. І пішов він, і осівся в щілині скелі Етам.
JUDG|15|9|І посходили филистимляни, і таборували в Юди, і розтяглися до Лехі.
JUDG|15|10|І сказали Юдині люди: Чого ви посходили проти нас? А ті відказали: Ми прийшли зв'язати Самсона, щоб зробити йому, як нам він зробив.
JUDG|15|11|І пішли три тисячі люда від Юди до щілини скелі Етам. І сказали вони Самсонові: Чи ти не знав, що над нами панують филистимляни? І що це ти нам учинив? А він їм сказав: Як вони зробили мені, так я зробив їм.
JUDG|15|12|І сказали йому: Ми зійшли зв'язати тебе, щоб віддати тебе в руку филистимлян. І сказав їм Самсон: Присягніть мені, що ви не заб'єте мене.
JUDG|15|13|А вони сказали йому, говорячи: Ні, а тільки зв'яжемо тебе та дамо тебе в їхню руку, а забити не заб'ємо тебе. І зв'язали його двома новими шнурами, і звели його зо скелі.
JUDG|15|14|Він прийшов аж до Лехі, а филистимляни зняли крик проти нього. І зійшов на нього Дух Господній, і стали ті сукані шнури, що на раменах його, як лляні, що перегоріли в огні, і поспадали з його рук пута його.
JUDG|15|15|І знайшов він свіжу ослячу щелепу, і простяг свою руку й узяв його, та й побив ним тисячу чоловіка.
JUDG|15|16|І сказав Самсон: Ослячою цією щелепою дійсно поклав їх на купу, ослячою цією щелепою тисячу люда побив я.
JUDG|15|17|І сталося, як скінчив він це говорити, то кинув ту щелепу зо своєї руки, і назвав ім'я тому місцю: Рамат-Лехі.
JUDG|15|18|І сильно він спрагнув, і кликнув до Господа та й сказав: Ти дав у руку Свого раба це велике спасіння, а тепер я помру від прагнення, і впаду в руку необрізаних.
JUDG|15|19|І пробив Бог джерело, що в Лехі, і вийшла з нього вода, і він напився, і вернувся його дух, і він ожив. Тому назвав він ім'я йому: Ен-Гаккоре, що в Лехі, і так воно зветься аж до цього дня.
JUDG|15|20|І судив він Ізраїля за днів филистимлян двадцять літ.
JUDG|16|1|І пішов Самсон до Гази, і побачив там жінку блудницю, і ввійшов до неї.
JUDG|16|2|А аззеянам донесли, говорячи: Самсон прийшов сюди! І оточили вони, і чатували на нього всю ніч у міській брамі. І вони тихо поводилися всю ніч, говорячи: Будемо чатувати аж до ранішнього світу, і заб'ємо його.
JUDG|16|3|І лежав Самсон аж до півночі. А опівночі встав, і схопив за двері міської брами та за обидва бічні одвірки, та й вирвав їх разом із засувом, і поклав на свої плечі, і виніс їх на верхів'я гори, що навпроти Хеврону.
JUDG|16|4|І сталося потому, і покохав він жінку в долині Сорек, а ім'я їй Деліла.
JUDG|16|5|І прийшли до неї филистимські володарі, та й сказали їй: Намов його та й побач, у чому його велика сила, і чим переможемо його та зв'яжемо його, щоб упокорити його? А ми кожен дамо тобі тисячу й сто шеклів срібла.
JUDG|16|6|І сказала Деліла до Самсона: Розкажи мені, у чому твоя велика сила, і чим можна зв'язати, щоб упокорити тебе?
JUDG|16|7|І сказав їй Самсон: Якщо зв'яжуть мене сімома мокрими шнурами, що ще не висушені, то ослабну та й стану, як кожен із людей.
JUDG|16|8|І принесли їй филистимські володарі сім мокрих шнурів, що ще не були висушені, а вона зв'язала його ними.
JUDG|16|9|А засідка сиділа в неї в іншій кімнаті. І вона сказала до нього: Филистимляни на тебе, Самсоне! І він розірвав ті шнури, як розривається нитка з клоччя, коли понюхає огню. І не пізнана була його сила.
JUDG|16|10|І сказала Деліла до Самсона: Оце ти обманив мене, і говорив мені лжу. Розкажи ж мені тепер, чим можна зв'язати тебе?
JUDG|16|11|А він їй сказав: Якщо справді зв'яжуть мене новими суканими шнурами, якими не робилася робота, то ослабну й стану, як кожен із людей.
JUDG|16|12|І взяла Деліла нові шнури, та й зв'язала його ними, і сказала до нього: Филистимляни на тебе, Самсоне! А засідка сиділа в іншій кімнаті. І він зірвав їх зо своїх плечей, немов нитку.
JUDG|16|13|І сказала Деліла Самсонові: Досі ти обманював мене, і говорив мені лжу. Розкажи ж мені, чим можна зв'язати тебе? А він їй сказав: Якщо утчеш сім кучерів моєї голови з основою.
JUDG|16|14|І вона прибила їх ткацьким клинком, та й сказала до нього: Филистимляни на тебе, Самсоне! А він обудився зо сну свого, та й вирвав ткацького клинка тканини та основу.
JUDG|16|15|І сказала вона до нього: Як ти говориш: кохаю тебе, а серце твоє не зо мною? Оце тричі обманив ти мене, і не розповів мені, у чому твоя велика сила.
JUDG|16|16|І сталося, коли вона докучала йому своїми словами по всі дні, та напирала на нього, то знетерпеливилася душа його на смерть.
JUDG|16|17|І виложив він їй усе серце своє, та й сказав їй: Бритва не торкалась моєї голови, бо я Божий назорей від утроби своєї матері. Якщо я буду оголений, то відступить від мене сила моя, і я ослабну, та й стану, як кожна людина.
JUDG|16|18|І побачила Деліла, що він розповів їй усе своє серце, і послала й покликала филистимських володарів, говорячи: Прийдіть і цим разом, бо він розповів мені все своє серце. І прийшли до неї филистимські володарі, і знесли срібло в своїй руці.
JUDG|16|19|А вона приспала його на колінах своїх, і покликала чоловіка та й наказала оголити сім кучерів його голови. І став він слабнути, і відступила від нього сила його.
JUDG|16|20|І сказала вона: Филистимляни на тебе, Самсоне! І збудився він зо сну свого та й сказав: Вийду я, як раз-у-раз, і стрясуся. А він не знав, що Господь відступився від нього.
JUDG|16|21|І взяли його филистимляни, та й вибрали очі йому. І вони звели його до Гази, і зв'язали його мідяними ланцюгами, і він молов у домі ув'язнених.
JUDG|16|22|А волос голови його зачав рости по тому, як був він оголений.
JUDG|16|23|А филистимські володарі зібралися, щоб принести велику жертву Даґонові, своєму богові, та повеселитися. І сказали вони: Наш бог передав у нашу руку Самсона, ворога нашого.
JUDG|16|24|І бачив його народ, і хвалили своїх богів, і говорили: Наш бог передав у нашу руку нашого ворога та спустошителя нашого краю, який наші трупи намножив.
JUDG|16|25|І сталося, коли їхнє серце звеселилося, то сказали вони: Покличте Самсона, і нехай він посмішить нас. І покликали Самсона з дому ув'язнених, і він витівав жарти перед ними, а вони поставили його поміж стовпами.
JUDG|16|26|І сказав Самсон юнакові, що держав його за руку: Пусти мене, і дай доторкнутися мені до тих стовпів, що на них цей дім стоїть міцно, і нехай я обіпруся на них.
JUDG|16|27|А той дім був повен чоловіків та жінок, і туди зібралися всі филистимські володарі, а на даху було близько трьох тисяч чоловіків та жінок, що приглядалися до жартів Самсона.
JUDG|16|28|І кликнув Самсон до Господа, та й сказав: Владико Господи, згадай же про мене, та зміцни мене тільки цього разу, Боже, і нехай я пімщу филистимлянам одну пімсту за двоє очей своїх!
JUDG|16|29|І обняв Самсон обидва серединні стовпи, що на них міцно стояв той дім, і обперся на них, на одного правицею своєю, а на одного лівицею своєю.
JUDG|16|30|І сказав Самсон: Нехай помру я разом із филистимлянами! І він з великою силою сперся на стовпи, і впав той дім на володарів та на ввесь той народ, що в ньому... І були ті померлі, що він повбивав їх при своїй смерті, численніші за тих, що повбивав їх за свого життя.
JUDG|16|31|І зійшли його брати та ввесь дім його батька, і понесли його, і винесли та й поховали його між Цор'а та між Ештаолом у гробі Маноаха, батька його. А він судив Ізраїля двадцять літ.
JUDG|17|1|І був чоловік з Єфремових гір, а ім'я йому Миха.
JUDG|17|2|І сказав він до своєї матері: Тисяча й сто шеклів срібла, що в тебе взяті, а ти прокляла за них, і також сказала це, щоб і я чув, ось те срібло зо мною, це я його взяв. І сказала мати його: Благословенний син мій у Господа!
JUDG|17|3|І він вернув ту тисячу й сто шеклів срібла своїй матері. І сказала його мати: Я справді посвятила те срібло Господеві з своєї руки за сина свого, щоб зробити боввана різьбленого та боввана литого. А тепер звертаю його тобі.
JUDG|17|4|Та він вернув те срібло своїй матері. І взяла його мати дві сотні шеклів срібла та й дала його золотареві, а він зробив із нього боввана різьбленого та боввана литого; і було це в домі Михи.
JUDG|17|5|А цей чоловік Миха мав удома божницю. І зробив він ефода та терафи, і висвятив одного з синів своїх, і він був йому за священика.
JUDG|17|6|Того часу не було царя в Ізраїлі, кожен робив, що правдиве було в його очах.
JUDG|17|7|І був юнак із Віфлеєму Юдиного, з Юдиного роду, а він Левит, і він був там приходько.
JUDG|17|8|І пішов той чоловік з того міста, із Віфлеєму Юдиного, щоб часово пожити, де знайде. І прийшов він до Єфремових гір до дому Михи, щоб далі йти своєю дорогою.
JUDG|17|9|І сказав йому Миха: Звідкіля ти приходиш? А той йому відказав: Я Левит із Віфлеєму Юдейського, а я йду, щоб часово пожити, де знайду.
JUDG|17|10|І сказав йому Миха: Зоставайся ж зо мною, і будь мені за отця та за священика, а я дам тобі десять шеклів срібла на рік і потрібну одежу та поживу твою. І пішов той Левит до нього,
JUDG|17|11|і погодився Левит сидіти з тим чоловіком. І був той юнак йому, як один із синів його.
JUDG|17|12|І Миха висвятив того Левита, і був йому той юнак за священика, і був у Михиному домі.
JUDG|17|13|І сказав Миха: Тепер я знаю, що Господь зробить добро мені, бо цей Левит став мені за священика.
JUDG|18|1|Того часу не було царя в Ізраїлі, і того часу Данове плем'я шукало собі наділу на оселю, бо до того дня не випало йому жеребка на наділ серед Ізраїлевих племен.
JUDG|18|2|І Данові сини послали зо свого роду п'ятеро люда з загалу людей військових, щоб вони вивідали Край та дослідили його. І сказали до них: Ідіть, дослідіть цей Край. І вони зійшли на Єфремові гори аж до Михиного дому, і переночували там.
JUDG|18|3|Коли вони були біля Михиного дому, то вони пізнали голос того юнака Левита, та й знайшли туди й сказали йому: Хто тебе привів сюди, і що ти тут робиш? І що ти тут маєш?
JUDG|18|4|І сказав він до них: Так і так зробив мені Миха, і він найняв мене, і я став йому за священика.
JUDG|18|5|А вони сказали йому: Запитай же Бога, і нехай ми пізнаємо, чи пощаститься наша дорога, якою ми йдемо.
JUDG|18|6|І сказав їм священик: Ідіть із миром, перед Господом ваша дорога, якою ви підете.
JUDG|18|7|І пішли ті п'ятеро людей, і прийшли в Лаїш та й побачили той народ, що в ньому, він сидить безпечно, за звичаєм сидонян, спокійний та безпечний. І не було нікого, хто робив би їм щось зле в Краю, посів би владу над ними, і вони далеко від сидонян, і нема їм діла ні до кого.
JUDG|18|8|І прийшли вони до братів своїх у Цор'у та в Ештаол. І сказали їм брати їх: Що ви принесли?
JUDG|18|9|А вони відказали: Устаньте, і підемо на них, бо ми бачили той Край, і ось дуже він добрий. А ви мовчите? Не лініться, щоб піти, щоб прийти та посісти той Край.
JUDG|18|10|Як ви підете, то ввійдете до народу безпечного, а Край той широкий, бо Бог дав його в вашу руку, це місце, що там нема недостачі жодної речі, що на землі.
JUDG|18|11|І рушили звідти з Данового роду з Цор'и та з Ештаолу шістсот чоловіка, оперезаних зброєю.
JUDG|18|12|І пішли вони й таборували в Кір'ят-Єарімі в Юді. Тому вони назвали ім'я тому місцю: Махане-Дан, і так воно зветься аж до цього дня, оце за Кір'ят-Єарімом.
JUDG|18|13|І перейшли вони звідти на Єфремові гори, і прийшли аж до Михиного дому.
JUDG|18|14|І відповіли п'ятеро тих мужів, що ходили вивідати той Край до Лаїшу, і сказали своїм браттям: Чи ви знаєте, що в цих домах є ефод та терафи, і бовван різьблений та бовван литий? А тепер знайте, що зробите.
JUDG|18|15|І вони зайшли туди до дому того юнака Левита, до Михиного дому, і запитали його про мир.
JUDG|18|16|А шість сотень мужа, що з Данових синів, оперезаних своєю зброєю, стояли при вході до брами.
JUDG|18|17|І пішли п'ятеро тих мужів, що ходили вивідати той Край, увійшли туди, узяли різьбленого боввана, і ефода та терафи, і боввана литого. А при вході до брами стояв священик та шістсот мужа, оперезаних зброєю.
JUDG|18|18|І ті ввійшли до Михиного дому, і взяли різьбленого боввана, ефода й терафи та боввана литого. І сказав до них той священик: Що ви робите?
JUDG|18|19|А вони відказали йому: Мовчи! Поклади свою руку на уста свої та й іди з нами, і стань нам за отця та за священика. Чи тобі ліпше бути священиком дому одного чоловіка, чи бути тобі священиком для племени та для роду Ізраїлевого?
JUDG|18|20|І стало добре на серці того священика, і він узяв ефода та терафи й різьбленого боввана, і ввійшов поміж народ.
JUDG|18|21|І повернулися вони та й пішли, а дітей, і худобу, і тягар пустили перед себе.
JUDG|18|22|Коли вони віддалилися від Михиного дому, то люди, що в домах, які разом із домом Михиним, були скликані, та й догнали Данових синів.
JUDG|18|23|І кричали вони до Данових синів, а ті обернули обличчя свої та й сказали до Михи: Що тобі, що ти кричиш?
JUDG|18|24|І він сказав: Ви забрали бога мого, що я зробив, та священика, та й пішли. І що мені ще? І що то ви говорите мені: що тобі?
JUDG|18|25|І сказали до нього Данові сини: Мовчи, щоб не чути нам твого голосу, а то наші люди із злости нападуть на вас, і ти долучиш душу свою до своєї рідні.
JUDG|18|26|І Данові сини пішли на свою дорогу. І побачив Миха, що вони сильніші від нього, і обернувся, та й пішов до свого дому.
JUDG|18|27|А вони взяли, що зробив був Миха, та священика, що був у нього, та й пішли на Лаїш, на народ спокійний та безпечний. І вони побили їх вістрям меча, а місто спалили огнем.
JUDG|18|28|А рятівника не було, бо далеке воно від Сидону, і не було в них діла ні з ким, і воно було в долині, що при Бет-Рехові. А вони збудували місто, та й осілися в ньому.
JUDG|18|29|І вони назвали ім'я тому містові: Дан, іменем Дана, їхнього батька, що був уроджений Ізраїлеві, але напочатку ім'я того міста було Лаїш.
JUDG|18|30|І поставили Данові сини того різьбленого боввана в себе, а Йонатан, син Ґершома, Манасіїного сина, він та сини його були священиками для Данового племени аж до дня виходу на вигнання того краю.
JUDG|18|31|І поклали вони в себе Михиного різьбленого боввана, що зробив він, і він був у них по всі дні буття Божого дому в Шіло.
JUDG|19|1|І сталося тими днями, а царя в Ізраїлі не було і був один Левит приходько на узбіччях Єфремових гір. І взяв він собі жінку наложницю з Юдиного Віфлеєму.
JUDG|19|2|А наложниця його чинила перелюб при ньому, та й пішла від нього до дому свого батька, до Віфлеєму Юдиного, і була там чотири місяці часу.
JUDG|19|3|І встав її муж та й пішов за нею, щоб поговорити до серця її, щоб вернути її, а з ним був слуга його та пара ослів. І вона ввела його до дому батька свого. І побачив його батько тієї молодої жінки, та й радісно вийшов назустріч йому.
JUDG|19|4|І тримав його тесть його, батько тієї молодої жінки, і сидів із ним три дні, і їли й пили вони та ночували там.
JUDG|19|5|І сталося четвертого дня, і повставали вони рано вранці, та й встали, щоб іти. І сказав батько тієї молодої жінки до зятя свого: Підкріпи своє серце кавалком хліба, а потім підете.
JUDG|19|6|І сіли вони, і обоє разом їли та пили. А батько тієї молодої жінки сказав до того чоловіка: Зволь же й переночуй, і нехай буде добре тобі на серці!
JUDG|19|7|Але встав той чоловік, щоб іти, а тесть його сильно просив його. І вернувся він, і переночував там.
JUDG|19|8|І встав він рано вранці п'ятого дня, щоб іти, а батько тієї молодої жінки сказав: Підкріпи ж своє серце! І зволікали вони аж до схилку дня, і їли обоє вони.
JUDG|19|9|І встав той чоловік, щоб іти, він та наложниця його та слуга його. І сказав йому тесть його, батько тієї молодої жінки: Ось день схилився на вечір, переночуй же! Ось день кладеться, ночуй тут, і нехай буде добре тобі на серці! І встанете взавтра рано, у дорогу свою, та й підеш до намету свого.
JUDG|19|10|Та той чоловік не хотів ночувати. І встав він та й пішов, і прийшов навпроти Євусу, це Єрусалим. А з ним пара нав'ючених ослів, і його наложниця з ним.
JUDG|19|11|Вони були при Євусі, а день дуже схилився. І сказав слуга до пана свого: Ходім, і зайдімо до цього євусейського міста, та й переночуємо в ньому.
JUDG|19|12|І сказав до нього пан його: Не заходьмо до міста чужинців, бо вони не з Ізраїлевих синів, а перейдімо до Ґів'и.
JUDG|19|13|І сказав він до слуги свого: Ходім, і прийдемо до одного з тих міст, і переночуємо в Ґів'ї або в Рамі.
JUDG|19|14|І перейшли вони та й пішли. А сонце зайшло їм при Ґів'ї, що була Веніяминова.
JUDG|19|15|І зійшли вони туди, щоб увійти переночувати в Ґів'ї. І він увійшов та й сів на майдані того міста, та ніхто не брав їх до дому переночувати.
JUDG|19|16|Аж ось старий чоловік іде ввечорі з поля з своєї роботи. А цей чоловік був з Єфремових гір, і він був приходько в Ґів'ї. А люди того місця сини Веніяминові.
JUDG|19|17|І звів він очі свої та й побачив того чоловіка мандрівника на міському майдані. І сказав той старий чоловік: Куди ти йдеш та звідки приходиш?
JUDG|19|18|А той до нього сказав: Ми переходимо з Юдиного Віфлеєму аж до узбіччя єфремових гір, звідти я. І ходив я аж до Юдиного Віфлеєму, і йду до Господнього дому, та нема нікого, хто взяв би мене до дому.
JUDG|19|19|Є й солома, і паша для наших ослів, є хліб та вино мені й невільниці твоїй та слузі з твоїми рабами, не бракує жодної речі.
JUDG|19|20|І сказав той старий чоловік: Мир тобі, нехай уся недостача твоя на мені, тільки на майдані не ночуй!
JUDG|19|21|І він увів його до свого дому, і дав ослам корму, а самі вони пообмивали ноги свої та й їли й пили.
JUDG|19|22|Коли вони звеселили серце своє, аж ось люди того міста, люди розпусні, оточили той дім та стукали в двері. І казали вони тому старому чоловікові, власникові того дому, говорячи: Виведи чоловіка, що ввійшов до дому твого, і ми пізнаєм його!
JUDG|19|23|І вийшов до них той чоловік, власник того дому, та й сказав їм: Ні, мої браття, не робіть же ви зла! По тому, як увійшов цей чоловік до мого дому, не зробіть такої гидоти!
JUDG|19|24|Ось дочка моя дівчина, та його наложниця, я їх виведу, а ви візьміть їх, і зробіть їм, що вам до вподоби, а тому чоловікові ви не зробите цієї огидної речі!
JUDG|19|25|Та ті люди не хотіли слухати його. І схопив той чоловік свою наложницю, і вивів до них назовні. І вони познали її, і безчестили її цілу ніч аж до ранку, і відпустили її, як зійшла рання зоря.
JUDG|19|26|І прийшла та жінка, як ранок вертався, та й упала, і лежала при вході дому того чоловіка, що пан її був там, аж до світу.
JUDG|19|27|А пан її встав рано, і відчинив двері дому та й вийшов, щоб іти своєю дорогою, аж ось та жінка, його наложниця, лежить при вході до дому, а руки її на порозі.
JUDG|19|28|І сказав він до неї: Уставай і підемо! Та вона не відповіла, бо вмерла. І взяв він її на осла. І встав той чоловік, і пішов до свого місця.
JUDG|19|29|І ввійшов він до дому свого, і взяв ножа, і схопив свою наложницю та й порізав її за костями її на дванадцять кусків, і порозсилав по всій Ізраїлевій країні.
JUDG|19|30|І сталося, кожен, хто це бачив, то говорив: Не бувало й не бачено такого, як це, від дня виходу Ізраїлевих синів з єгипетського краю аж до цього дня! Зверніть увагу на це, радьте та говоріть!
JUDG|20|1|І повиходили всі Ізраїлеві сини, і була зібрана громада, як один чоловік, від Дану аж до Беер-Шеви, а ґілеадський край до Господа в Міцпу.
JUDG|20|2|І стали проводирі всього того народу, усі Ізраїлеві племена, на зборах Божого народу, чотириста тисяч пішого люду, хто витягує меча.
JUDG|20|3|І почули Веніяминові сини, що Ізраїлеві сини ввійшли до Міцпи. І сказали Ізраїлеві сини: Скажіть, як сталося таке зло?
JUDG|20|4|І відповів той чоловік Левит, чоловік тієї замордованої жінки, та й сказав: До Ґів'и, що Веніяминова, увійшов я та наложниця моя, щоб ночувати.
JUDG|20|5|І встали на мене господарі Ґів'и, і вночі оточили через мене той дім. Мене замишляли забити, а наложницю мою збезчестили, і померла вона.
JUDG|20|6|І схопив я наложницю, і порізав її, та й послав її по всьому полі Ізраїлевого володіння, бо вони вчинили розпусту та гидоту серед Ізраїля.
JUDG|20|7|Ось ви всі Ізраїлеві сини, дайте собі тут слово та раду!
JUDG|20|8|І встав увесь народ, як один муж, говорячи: Не підемо ніхто до намету свого, і не знайдемо ніхто до дому свого!
JUDG|20|9|А тепер оце та річ, що зробимо Ґів'ї: підемо на неї за жеребком!
JUDG|20|10|І візьмемо десятеро людей на сотню, щодо всіх Ізраїлевих племен, і сотню на тисячу, і тисячу на десять тисяч, щоб узяли поживи для народу, щоб вони прийшли зробити Ґів'ї Веніямина, згідно з усією гидотою, що він зробив Ізраїлеві.
JUDG|20|11|І був зібраний кожен ізраїльтянин до того міста разом, як один чоловік.
JUDG|20|12|І послали Ізраїлеві племена людей по всіх Веніяминових родах, говорячи: Що це за зло, що сталось між вами?
JUDG|20|13|А тепер давайте тих людей, розпусних синів, що в Ґів'ї, і ми повбиваємо їх, та й вигубимо зло з Ізраїля. Та не хотіли Веніяминові сини слухати голосу своїх братів, Ізраїлевих синів.
JUDG|20|14|І Веніяминові сини були зібрані з міст до Ґів'ї, щоб піти на війну з Ізраїлевими синами.
JUDG|20|15|І Веніяминові сини з міст були перелічені того дня, двадцять і шість тисяч чоловіка, що витягують меча, окрім мешканців Ґів'и, із них були перелічені сім сотень вибраного чоловіка.
JUDG|20|16|З усього того народу було сім сотень вибраного чоловіка, із нечинною рукою правиці своєї, лівші, кожен той кидав каменем із пращі на волос, і не схибував.
JUDG|20|17|І були перелічені ізраїльтяни, окрім Веніямина, чотириста тисяч чоловіка, що витягують меча, кожен військовий.
JUDG|20|18|І встали вони, і ввійшли до Бет-Елу, і питалися Бога, та й сказали Ізраїлеві сини: Хто піде нам спереду на бій з Веніяминовими синами? І сказав Господь: Юда спереду.
JUDG|20|19|І встали Ізраїлеві сини рано вранці, і таборували при Ґів'ї.
JUDG|20|20|І вийшов Ізраїльтянин на війну з Веніямином, і сточили ізраїльтяни з ними бій при Ґів'ї.
JUDG|20|21|І вийшли Веніяминові сини з Ґів'и, та й повалили між Ізраїлем того дня двадцять і дві тисячі чоловіка на землю.
JUDG|20|22|І зміцнився народ, Ізраїлеві мужі, і точили бій далі в тому місці, де точили бій першого дня.
JUDG|20|23|І ввійшли Ізраїлеві сини до Бет-Елу, та й плакали перед Господнім лицем аж до вечора. І питалися вони Господа, говорячи: Чи далі піду я на бій з синами Веніямина, мого брата? І сказав Господь: Ідіть на нього!
JUDG|20|24|І прийшли Ізраїлеві сини до Веніяминових синів дня другого.
JUDG|20|25|А Веніямин вийшов із Ґів'ї другого дня навпроти них, та й повалив між Ізраїлевими синами на землю ще вісімнадцять тисяч чоловіка, усі ті, що витягають меча.
JUDG|20|26|І прийшли всі Ізраїлеві сини та ввесь народ, і ввійшли до Бет-Елу, та й плакали, і сиділи там перед Господнім лицем, і постили того дня аж до вечора. І принесли вони цілопалення та мирні жертви перед Господнім лицем.
JUDG|20|27|І питалися Ізраїлеві сини Господа (а за тих днів ковчег Божого заповіту був там.
JUDG|20|28|А Пінхас, син Елеазара, Ааронового сина, стояв тими днями перед Його лицем), говорячи: Чи далі піду ще на бій з синами Веніямина, мого брата, чи спинюся? А Господь сказав: Ідіть, бо взавтра Я дам його в твою руку.
JUDG|20|29|І поставив Ізраїль засідку навколо Ґів'ї.
JUDG|20|30|І пішли Ізраїлеві сини на синив Веніяминових третього дня, і сточили бій проти Ґів'ї, як і раніш.
JUDG|20|31|І вийшли Веніяминові сини навпроти народу, одірвалися від міста, і зачали класти трупи з народу, як раз-у-раз, на битих дорогах, що одна йде до Бет-Елу, а одна до Ґів'ї, у полі, коло тридцяти чоловіка між Ізраїлем.
JUDG|20|32|І сказали Веніяминові сини: Биті вони перед нами, як перше! А Ізраїлеві сини сказали: Утікаймо, і відірвемо їх від міста на дороги.
JUDG|20|33|І кожен муж Ізраїля повстав із свого місця, і сточили бій у Баал-Тамарі, а Ізраїлева засідка рушила з свого місця, з Мааре-Ґева.
JUDG|20|34|І прийшли перед Ґів'у десять тисяч чоловіка, вибраного з усього Ізраїля, і бій став тяжкий. А вони не знали, що суне на них те зло.
JUDG|20|35|І вдарив Господь Веніямина перед Ізраїлем, і Ізраїлеві сини повалили того дня між Веніямином двадцять і п'ять тисяч і сто чоловіка, усі ті, що витягають меча.
JUDG|20|36|І побачили Веніяминові сини, що побиті вони, а ізраїльтяни уступили місце Веніяминові, бо вірили засідці, яку поставили на Ґів'у.
JUDG|20|37|А засідка поспішилася, і напала на Ґів'у. І засідка вступилася, і побила все місто вістрям меча.
JUDG|20|38|А Ізраїльтянин мав із засідкою умовленого знака, щоб із міста підняла великий дим.
JUDG|20|39|І відступили ізраїльтяни в бою, а Веніямин зачав класти трупи в Ізраїлі, близько тридцятеро люда, бо казали вони: Дійсно, справді побитий він перед нами, як за першого бою!
JUDG|20|40|А з міста став підійматися стовп диму. І обернувся Веніямин позад себе, аж ось усе місто піднялося димом до неба!
JUDG|20|41|І обернувся Ізраїльтянин, а Веніяминівець перестрашився, бо побачив, що досягло його те зло.
JUDG|20|42|І обернулися вони перед Ізраїльтянином до дороги на пустиню, та бій досягав його, а ті, що з міст, валили його в середині його.
JUDG|20|43|Вони оточили Веніямина, гнали його до Менухи, топтали його аж до Ґів'ї зо сходу сонця.
JUDG|20|44|Полягло тоді з Веніямина вісімнадцять тисяч чоловіка, усе це люди хоробрі.
JUDG|20|45|І повернулися вони, і втікли в пустиню до Села-Ріммону. А ті побили поодиноких утікачів по дорогах, як дозбирюється останній виноград, п'ять тисяч люда. І гналися за ними аж до Ґід'ому, і побили з нього дві тисячі люда.
JUDG|20|46|І було всіх, що впали того дня з Веніямина, двадцять і п'ять тисяч чоловіка, що витягають меча, усе це люди хоробрі.
JUDG|20|47|І обернулися вони, і повтікали в пустиню до Села-Ріммону, шістсот чоловіка. І сиділи вони в Села-Ріммоні чотири місяці.
JUDG|20|48|А ізраїльтяни вернулися до Веніяминових синів, та й повбивали їх вістрям меча, мужчин із міста, і худобу, і все знайдене. А всі міста, що знаходились по дорозі, пустили з огнем.
JUDG|21|1|І присягнув Ізраїльтянин в Міцпі, говорячи: Жоден із нас не дасть своєї дочки Веніяминові за жінку!
JUDG|21|2|І посходився народ до Бет-Елу, та й сидів там аж до вечора перед Божим лицем. І піднесли вони голос свій, та й плакали плачем великим.
JUDG|21|3|І сказали вони: Чому, Господи, Боже Ізраїлів, сталося це між Ізраїлем, щоб сьогодні бракувало з Ізраїля одне плем'я?
JUDG|21|4|І сталося назавтра, і встав рано народ, та й збудували жертівника, і принесли цілопалення та мирні жертви.
JUDG|21|5|І сказали Ізраїлеві сини: Хто зо всіх Ізраїлевих племен не ввійшов до зборів до Господа? Бо та присяга була велика на того, хто не прийшов до Господа, до Міцпи, говорячи: Такий буде конче забитий.
JUDG|21|6|І жалували Ізраїлеві сини за Веніямином, своїм братом, та й сказали: Сьогодні відрубане з Ізраїля одне плем'я!
JUDG|21|7|Що ми зробимо їм, позосталим, щодо жінок? А ми присягнули Господом, що не дамо їм із дочок наших за жінок.
JUDG|21|8|І сказали вони: Яке одне з Ізраїлевих племен не прийшло до Господа до Міцпи? Аж ось виявилось, що з Явешу ґілеадського ніхто не приходив до табору на збори.
JUDG|21|9|І був переглянений народ, а оце не було там нікого з мешканців Явешу ґілеадського!
JUDG|21|10|І послала громада туди дванадцять тисяч чоловіка хоробрих людей, і наказали їм, говорячи: Ідіть, і повбиваєте мешканців ґілеадського Явешу вістрям меча, і жінок і дітей.
JUDG|21|11|А це та річ, що ви зробите: Кожного чоловіка та кожну жінку, що пізнала чоловіка, зробите закляттям.
JUDG|21|12|І знайшли вони з мешканців ґілеадського Явешу чотири сотні дівчат паннів, що не пізнали чоловіка, і спровадили їх до табору в Шіло, що в ханаанському Краї.
JUDG|21|13|І послала вся та громада, а ті говорили до Веніяминових синів, що в Села-Ріммоні, та й кликнули їм: Мир!
JUDG|21|14|І вернувся Веніямин того часу, і дали їм тих жінок, яких позоставили при житті, із жінок ґілеадського Явешу. Та не знайшли їм досить.
JUDG|21|15|А народ той жалував за Веніямином, бо Господь зробив пролома в Ізраїлевих племенах.
JUDG|21|16|І сказали старші громади: Що ми зробимо позосталим щодо жінок? Бо вигублена жінка з Веніямина.
JUDG|21|17|І сказали вони: Останки насліддя для Веніямина, і не буде витерте плем'я з Ізраїля.
JUDG|21|18|А ми не можемо дати їм жінок із наших дочок, бо Ізраїлеві сини присягли, говорячи: Проклятий, хто дає жінку Веніяминові!
JUDG|21|19|І сказали вони: Ось буває рік-у-рік свято Господнє в Шіло, що на північ від Бет-Елу, на схід сонця від дороги, що провадить з Бет-Елу до Сихему, і з півдня від Левони.
JUDG|21|20|І наказали вони Веніяминовим синам, говорячи: Ідіть, і будете чатувати в виноградниках.
JUDG|21|21|І побачите, аж ось дочки Шіла вийдуть танцювати танці, то ви вийдете з виноградників, та й схопите собі кожен свою жінку з дочок Шіла, і підете в Веніяминів край.
JUDG|21|22|І буде, коли їхні батьки або їхні брати прийдуть до нас сваритися, то ми скажемо їм: Змилуйтеся над ними, бо не взяли ми для кожного з них жінку на війні, і ви не дали їж, тому цього часу ви винні.
JUDG|21|23|І зробили так Веніяминові сини, і взяли жінок за числом своїм із тих, що танцювали, що їх вони викрали. І пішли вони, і вернулися до наділу свого, і побудували міста, та й осілися в них.
JUDG|21|24|І порозходилися звідти Ізраїлеві сини того часу кожен до племени свого та до роду свого, і пішли звідти кожен до спадку свого.
JUDG|21|25|Того часу не було царя в Ізраїлі, кожен робив, що здавалося правдивим в його очах!
