JER|1|1|Verba Ieremiae filii Helciae de sacerdotibus, qui fuerunt in Anathoth in terra Beniamin.
JER|1|2|Quod factum est verbum Domini ad eum in diebus Iosiae filii Amon regis Iudae, in tertio decimo anno regni eius.
JER|1|3|Et factum est in diebus Ioachim filii Iosiae regis Iudae, usque ad consummationem undecimi anni Sedeciae filii Iosiae regis Iudae, usque ad transmigrationem Ierusalem in mense quinto.
JER|1|4|Et factum est verbum Domini ad me dicens:
JER|1|5|" Priusquam te formarem in utero, novi teet, antequam exires de vulva, sanctificavi teet prophetam gentibus dedi te ".
JER|1|6|Et dixi: " Heu, Domine Deus! Ecce nescio loqui, quia puer ego sum ".
JER|1|7|Et dixit Dominus ad me: " Noli dicere: "Puer sum",quoniam, ad quoscumque mittam te, ibiset universa, quaecumque mandavero tibi, loqueris.
JER|1|8|Ne timeas a facie eorum,quia tecum ego sum, ut eruam te ",dicit Dominus.
JER|1|9|Et misit Dominus manum suam et tetigit os meum; et dixit Dominus ad me: Ecce dedi verba mea in ore tuo;
JER|1|10|ecce constitui te hodie super gentes et super regna,ut evellas et destruaset disperdas et dissipeset aedifices et plantes ".
JER|1|11|Et factum est verbum Domini ad me dicens: " Quid tu vides, Ieremia? ". Et dixi: " Virgam amygdali vigilantis ego video ".
JER|1|12|Et dixit Dominus ad me: "Bene vidisti, quia vigilo ego super verbo meo, ut faciam illud ".
JER|1|13|Et factum est verbum Domini secundo ad me dicens: " Quid tu vides? ". Et dixi: " Ollam succensam ego video; et facies eius a facie aquilonis ".
JER|1|14|Et dixit Dominus ad me: Ab aquilone pandetur malumsuper omnes habitatores terrae;
JER|1|15|quia ecce ego convocaboomnia regna aquilonis,ait Dominus,et venient et ponent unusquisque solium suumin introitu portarum Ierusalemet contra omnes muros eius in circuituet contra universas urbes Iudae;
JER|1|16|et loquar iudicia mea cum eissuper omnem malitiam eorum,qui dereliquerunt meet incensum obtulerunt diis alieniset adoraverunt opus manuum suarum.
JER|1|17|Tu ergo accinge lumbos tuoset surge et loquere ad eos omnia,quae ego praecipio tibi;ne timeas a facie eorum,alioquin timere te faciam vultum eorum.
JER|1|18|Ego quippe dedi te hodiein civitatem munitamet in columnam ferreamet in murum aereumcontra omnem terramregibus Iudae, principibus eiuset sacerdotibus et populo terrae;
JER|1|19|et bellabunt adversum te et non praevalebunt,quia tecum ego sum,ait Dominus,ut eripiam te ".
JER|2|1|Et factum est verbum Domini ad me dicens:
JER|2|2|" Vade et clama in auribus Ierusalem dicens:Haec dicit Dominus:Recordatus sum tui, caritatis adulescentiae tuaeet amoris desponsationis tuae,quando secuta es me in deserto,in terra, quae non seminatur.
JER|2|3|Sanctus Domino Israel,primitiae frugum eius;omnes, qui devorabant eum, delinquebant;mala veniebant super eos,dicit Dominus.
JER|2|4|Audite verbum Domini, domus Iacobet omnes cognationes domus Israel.
JER|2|5|Haec dicit Dominus:Quid invenerunt patres vestri in me iniquitatis,quia elongaverunt a meet ambulaverunt post vanitatemet vani facti sunt?
JER|2|6|Et non dixerunt: "Ubi est Dominus,qui ascendere nos fecit de terra Aegypti,qui traduxit nos per desertum,per terram inhabitabilem et inviam,per terram sitis et caliginis,per terram, in qua non ambulavit vir,neque habitavit homo?".
JER|2|7|Et induxi vos in terram hortorum,ut comederetis fructum eius et optima illius;et ingressi contaminastis terram meamet hereditatem meam posuistis in abominationem.
JER|2|8|Sacerdotes non dixerunt:Ubi est Dominus?".Et tractantes legem nescierunt me,et pastores praevaricati sunt in me,et prophetae prophetaverunt in Baalet, quae nihil prosunt, secuti sunt.
JER|2|9|Propterea adhuc iudicio contendam vobiscum,ait Dominus,et cum filiis filiorum vestrorum disceptabo.
JER|2|10|En transite ad insulas Cetthim et videteet in Cedar mittite et considerate vehementeret videte, si factum est huiuscemodi:
JER|2|11|si mutavit gens deos,et certe ipsi non sunt dii;populus vero meus mutavit gloriam suamin id, quod nihil prodest.
JER|2|12|Obstupescite, caeli, super hocet inhorrescite supra modum,dicit Dominus.
JER|2|13|Duo enim mala fecit populus meus:me dereliquerunt fontem aquae vivae,ut foderent sibi cisternas,cisternas dissipatas,quae continere non valent aquas.
JER|2|14|Numquid servus est Israelaut vernaculus?Quare ergo factus est in praedam?Super eum rugierunt leones
JER|2|15|et dederunt vocem suam;posuerunt terram eius in solitudinem:civitates eius exustae sunt,et non est qui habitet in eis.
JER|2|16|Filii quoque Mempheos et Taphnesdecalvabunt tibi verticem.
JER|2|17|Numquid non istud factum est tibi,quia dereliquisti Dominum Deum tuumeo tempore, quo ducebat te per viam?
JER|2|18|Et nunc quid tibi vis in via Aegypti,ut bibas aquam Nili?Et quid tibi cum via Assyriorum,ut bibas aquam Fluminis?
JER|2|19|Arguet te malitia tua,et aversio tua increpabit te;scito et vide quia malum et amarum estreliquisse te Dominum Deum tuum et non esse timorem mei apud te,dicit Dominus, Deus exercituum.
JER|2|20|A saeculo confregisti iugum tuum,rupisti vincula tuaet dixisti: "Non serviam".In omni enim colle sublimiet sub omni ligno frondosotu prosternebaris meretrix.
JER|2|21|Ego autem plantavi te vineam electam,omne semen verum;quomodo ergo conversa esin palmites vineae alienae?
JER|2|22|Si laveris te nitroet multiplicaveris tibi herbam fullonum,maculata es in iniquitate tua coram me,dicit Dominus Deus.
JER|2|23|Quomodo dicis: "Non sum polluta,post Baalim non ambulavi"?Vide viam tuam in convalle,scito quid feceris:camelus levis contorquens vias suas.
JER|2|24|Onager assuetus in solitudinein desiderio animae suae attrahit aerem;libidinem eius quis avertet?Omnes, qui quaerunt eam, non deficient,in menstruis eius invenient eam.
JER|2|25|Prohibe pedem tuum a nuditateet guttur tuum a siti.Et dixisti: "Vanum est, nequaquam;adamavi quippe alienoset post eos ambulabo".
JER|2|26|Quomodo confunditur fur, quando deprehenditur,sic confusi sunt domus Israel,ipsi et reges eorum, principeset sacerdotes et prophetae eorum
JER|2|27|dicentes ligno: "Pater meus es tu" et lapidi: "Tu me genuisti".Verterunt ad me tergum et non faciem,sed in tempore afflictionis suae dicent:Surge et libera nos!".
JER|2|28|Ubi sunt dii tui, quos fecisti tibi?Surgant et liberent te in tempore afflictionis tuae;secundum numerum quippe civitatum tuarumfacti sunt dii tui, Iuda.
JER|2|29|Quid vultis mecum iudicio contendere?Omnes praevaricati estis in me,dicit Dominus.
JER|2|30|Frustra percussi filios vestros:disciplinam non receperunt.Devoravit gladius vester prophetas vestros:quasi leo vastator.
JER|2|31|O generatio, vos videte verbum Domini:numquid solitudo factus sum Israeliaut terra tenebrarum?Quare ergo dixit populus meus: "Recessimus,non veniemus ultra ad te"?
JER|2|32|Numquid obliviscitur virgo ornamenti sui,sponsa fasciae pectoralis suae?Populus vero meus oblitus est meidiebus innumeris.
JER|2|33|Quam bene paras viam tuamad quaerendum amorem!Et insuper in malumdocuisti vias tuas,
JER|2|34|et in fimbriis tuis inventus estsanguis animarum pauperum innocentium:non effringentes invenisti eos;sed in omnibus his
JER|2|35|dixisti: "Innocens ego sum,propterea aversus est furor eius a me".Ecce ego iudicio contendam tecum, eo quod dixeris: "Non peccavi".
JER|2|36|Quam leviter mutas vias tuas!Et ab Aegypto confunderis,sicut confusa es ab Assyria.
JER|2|37|Nam et ab ista egredieris,et manus tuae erunt super caput tuum,quoniam obtrivit Dominus illos, quibus confisus es,et nihil habebis prosperum in eis.
JER|3|1|Si dimiserit vir uxorem suam,et recedens ab eoduxerit virum alterum,numquid revertetur ad eam ultra?Numquid non pollutaet contaminata est terra illa?Tu autem fornicata es cum amatoribus multiset reverteris ad me?,dicit Dominus.
JER|3|2|Leva oculos tuos ad colles et vide,ubi non prostrata sis.In viis sedebas exspectans eosquasi Arabs in solitudine;et polluisti terramin fornicationibus tuis et in malitia tua.
JER|3|3|Quam ob rem prohibitae sunt stillae pluviarum,et serotinus imber non fuit.Frons mulieris meretricis facta est tibi;noluisti erubescere.
JER|3|4|Nonne amodo vocas me: "Pater meus,dux adulescentiae meae tu es!
JER|3|5|Numquid irascetur in perpetuumaut perseverabit in finem?".Ecce locuta eset fecisti mala et praevaluisti ".
JER|3|6|Et dixit Dominus ad me in diebus Iosiae regis: " Numquid vidisti, quae fecerit aversatrix Israel? Abiit sibimet super omnem montem excelsum et sub omni ligno frondoso et fornicata est ibi.
JER|3|7|Et dixi: "Cum fecerit haec omnia, ad me revertetur"; et non est reversa. Et vidit praevaricatrix soror eius, Iuda;
JER|3|8|et vidit quia pro eo quod moechata esset aversatrix Israel, dimisissem eam et dedissem ei libellum repudii, et non timuit praevaricatrix Iuda, soror eius, sed abiit et fornicata est etiam ipsa;
JER|3|9|et facilitate fornicationis suae contaminavit terram et moechata est cum lapide et ligno.
JER|3|10|Sed in omnibus his non est reversa ad me praevaricatrix soror eius Iuda in toto corde suo sed in mendacio ", ait Dominus.
JER|3|11|Et dixit Dominus ad me: " Iustificavit animam suam aversatrix Israel comparatione praevaricatricis Iudae.
JER|3|12|Vade et clama sermones istos contra aquilonem et dices:Revertere, aversatrix Israel,ait Dominus,et non avertam faciem meam a vobis,quia pius ego sum,dicit Dominus,et non irascar in perpetuum.
JER|3|13|Verumtamen scito iniquitatem tuam,quia in Dominum Deum tuum praevaricata eset dispersisti vias tuas alienissub omni ligno frondoso;et vocem meam non audistis,ait Dominus.
JER|3|14|Convertimini, filii, qui aversi estis a me, dicit Dominus, quia ego Dominus vester sum; et assumam vos unum de civitate et duos de cognatione et introducam vos in Sion;
JER|3|15|et dabo vobis pastores iuxta cor meum, et pascent vos scientia et doctrina.
JER|3|16|Cumque multiplicati fueritis et creveritis in terra in diebus illis, ait Dominus, non dicent ultra: "Arca testamenti Domini", neque ascendet super cor, neque recordabuntur illius, nec requiretur, nec fiet ultra.
JER|3|17|In tempore illo vocabunt Ierusalem Solium Domini, et congregabuntur ad eam omnes gentes in nomine Domini in Ierusalem; et non ambulabunt ultra post pravitatem cordis sui pessimi.
JER|3|18|In diebus illis ibit domus Iudae ad domum Israel, et venient simul de terra aquilonis ad terram, quam dedi in hereditatem patribus vestris.
JER|3|19|Ego autem dixi:Quomodo ponam te in filiiset tribuam tibi terram desiderabilem,hereditatem praeclarissimam inter gentes?Et dixi: Patrem vocabitis meet post me ingredi non cessabitis.
JER|3|20|Sed, quomodo contemnit mulier amatorem suum,sic contempsistis me, domus Israel ",dicit Dominus.
JER|3|21|Vox in collibus audita est,ploratus et supplicatio filiorum Israel,quoniam iniquam fecerunt viam suam,obliti sunt Domini Dei sui.
JER|3|22|" Convertimini, filii, qui aversi estis a me,et sanabo aversiones vestras ". Ecce nos venimus ad te;tu enim es Dominus Deus noster.
JER|3|23|Vere mendaces erant colleset tumultus montium;vere in Domino Deo nostrosalus Israel.
JER|3|24|Confusio comedit laborem patrum nostrorumab adulescentia nostra,greges eorum et armenta eorum,filios eorum et filias eorum.
JER|3|25|Dormiemus in confusione nostra,et operiet nos ignominia nostra,quoniam Domino Deo nostro peccavimusnos et patres nostriab adulescentia nostra usque ad hanc diemet non audivimus vocem Domini Dei nostri ".
JER|4|1|" Si converteris, Israel,ait Dominus,ad me convertere;si abstuleris abominationes tuas a facie mea,non effugies.
JER|4|2|Et iurabis: "Vivit Dominus!"in veritate et in iudicio et in iustitia,et benedicentur in ipso genteset in ipso gloriabuntur.
JER|4|3|Haec enim dicit Dominusviro Iudae et Ierusalem:Novate vobis novaleet nolite serere super spinas.
JER|4|4|Circumcidimini Dominoet auferte praeputia cordium vestrorum,viri Iudae et habitatores Ierusalem,ne forte egrediatur ut ignis indignatio meaet succendatur, et non sit qui exstinguat,propter malitiam operum vestrorum.
JER|4|5|Annuntiate in Iudaet in Ierusalem auditum facite;et loquimini et canite tuba in terra,clamate fortiter et dicite:Congregamini, et ingrediamur civitates munitas".
JER|4|6|Levate signum in Sion,fugite, nolite stare,quia malum ego adduco ab aquiloneet contritionem magnam.
JER|4|7|Ascendit leo de cubili suo,et praedo gentium se levavit;egressus est de loco suo,ut ponat terram tuam in solitudinem:civitates tuae vastabuntur,remanentes absque habitatore.
JER|4|8|Super hoc accingite vos ciliciis,plangite et ululate,quia non est aversa ira furoris Domini a nobis.
JER|4|9|Et erit in die illa,dicit Dominus,peribit cor regiset cor principum,et obstupescent sacerdotes,et prophetae consternabuntur ".
JER|4|10|Et dixi: " Heu, Domine Deus!Ergo decepisti populum istum et Ierusalemdicens: "Pax erit vobis";et ecce pervenit gladius usque ad animam ".
JER|4|11|In tempore illo dicetur populo huic et Ierusalem: Ventus urens collium, qui sunt in deserto,invadit filiam populi meinon ad ventilandum et ad purgandum.
JER|4|12|Ventus plenior his veniet mihi,nunc et ego loquar iudicia mea cum eis ".
JER|4|13|Ecce quasi nubes ascendet,et quasi tempestas currus eius;velociores aquilis equi illius.Vae nobis, quoniam vastati sumus!
JER|4|14|Lava a malitia cor tuum,Ierusalem, ut salva fias;usquequo morabuntur in tecogitationes iniquae?
JER|4|15|Vox enim annuntiantis a Danet notam facientis calamitatem de monte Ephraim.
JER|4|16|Nuntiate gentibus. Ecce adsunt!Auditum facite hoc super Ierusalem: Custodes venerunt de terra longinquaet dederunt super civitates Iudae vocem suam;
JER|4|17|quasi custodes agrorum facti sunt super eam in gyro,quia adversus me contumax erat ",dicit Dominus.
JER|4|18|Via tua et opera tuafecerunt haec tibi;ista malitia tua, quia amara,quia tetigit cor tuum.
JER|4|19|Viscera mea, viscera mea! Doleo.Parietes cordis mei!Turbatur in me cor meum:non tacebo,quoniam vocem bucinae audivit anima mea,clamorem proelii.
JER|4|20|Contritio super contritionem vocata est,quoniam vastata est omnis terra,repente vastata sunt tabernacula mea,subito tentoria mea.
JER|4|21|Usquequo videbo vexillum,audiam vocem bucinae?
JER|4|22|" Quia stultus populus meus:me non cognoverunt;filii insipientes sunt et vecordes:sapientes sunt, ut faciant mala,bene autem facere nesciunt ".
JER|4|23|Aspexi terram, et ecce vacua erat et deserta;et caelos, et non erat lux in eis.
JER|4|24|Aspexi montes, et ecce movebantur,et omnes colles conturbati sunt.
JER|4|25|Aspexi, et ecce non erat homo,et omne volatile caeli recesserat.
JER|4|26|Aspexi, et ecce hortus desertus,et omnes urbes eius destructae sunta facie Domini et a facie irae furoris eius.
JER|4|27|Haec enim dicit Dominus: Deserta erit omnis terra,sed tamen consummationem non faciam.
JER|4|28|Super hoc lugebit terra,et maerebunt caeli desuper,eo quod locutus sum,statui et non paenitet menec avertar ab eo ".
JER|4|29|A voce equitis et mittentis sagittamfugit omnis civitas;ingressi sunt silvas condensaset ascenderunt rupes;universae urbes derelictae sunt,et non habitat in eis homo.
JER|4|30|Tu autem, vastata, quid facies?Cum vestieris te coccino,cum ornata fueris monili aureo,et pinxeris stibio oculos tuos,frustra componeris;contempserunt te amatores tui,animam tuam quaerent.
JER|4|31|Vocem enim quasi parturientis audivi,angustias ut puerperae;vox filiae Sionintermorientis expandentisque manus suas: Vae mihi, quia defecit anima meapropter interfectores! ".
JER|5|1|Circuite vias Ierusalemet aspicite et considerateet quaerite in plateis eius,an inveniatis virum,an sit qui faciat iudicium et quaerentem fidem,et propitius ero ei.
JER|5|2|Quod si etiam " Vivit Dominus! " dixerint,certe falso iurabunt.
JER|5|3|Domine, nonne oculi tui respiciunt fidem?Percussisti eos, et non doluerunt,attrivisti eos, et renuerunt accipere disciplinam:induraverunt facies suas supra petram,noluerunt reverti.
JER|5|4|Ego autem dixi: " Ecce pauperes illi stulte agunt,quia ignorant viam Domini,iudicium Dei sui.
JER|5|5|Ibo igitur ad optimateset loquar eis;ipsi enim noverunt viam Domini,iudicium Dei sui ".Ecce hi simul confregerunt iugum, ruperunt vincula.
JER|5|6|Idcirco percussit eos leo de silva,lupus deserti vastabit eos,pardus vigilans super civitates eorum:omnis, qui egressus fuerit ex eis, lacerabitur,quia multiplicatae sunt praevaricationes eorum,confortatae sunt aversiones eorum.
JER|5|7|" Super quo propitius tibi esse potero?Filii tui dereliquerunt meet iuraverunt in his, qui non sunt dii;saturavi eos, et moechati suntet in domum meretricis gregatim confluebant.
JER|5|8|Equi impinguati et admissarii facti sunt:unusquisque ad uxorem proximi sui hinniebat.
JER|5|9|Numquid super his non visitabo,dicit Dominus,et in gente tali non ulciscetur anima mea?
JER|5|10|Ascendite muros eius et dissipate,consummationem autem nolite facere;auferte propagines eius,quia non sunt Domini.
JER|5|11|Praevaricatione enim praevaricata est in medomus Israel et domus Iudae ",ait Dominus.
JER|5|12|Negaverunt Dominumet dixerunt: "Non est ipse;neque veniet super nos malum,et gladium et famem non videbimus.
JER|5|13|Prophetae erunt in ventum,et responsum non est in eis.Haec ergo evenient illis ".
JER|5|14|Propterea haec dicit Dominus, Deus exercituum: Quia locuti estis verbum istud,ecce ego do verba mea in ore tuo in ignemet populum istum in ligna,et vorabit eos.
JER|5|15|Ecce ego adducam super vos gentem de longinquo,domus Israel,ait Dominus,gentem robustam,gentem antiquam,gentem, cuius ignorabis linguamnec intelleges quid loquatur.
JER|5|16|Pharetra eius quasi sepulcrum patensuniversi fortes.
JER|5|17|Et comedet segetes tuas et panem tuum,devorabit filios tuos et filias tuas,comedet gregem tuum et armenta tua,comedet vineam tuam et ficum tuam;et conteret urbes munitas tuas,in quibus tu habes fiduciam, gladio.
JER|5|18|Verumtamen et in diebus illis,ait Dominus,non faciam in vobis consummationem ".
JER|5|19|Quod si dixeritis: " Quare fecit nobis Dominus Deus noster haec omnia?, dices ad eos: " Sicut dereliquistis me et servistis diis alienis in terra vestra, sic servietis alienis in terra non vestra ".
JER|5|20|Annuntiate hoc domui Iacobet auditum facite in Iuda dicentes:
JER|5|21|" Audi, popule stulte, qui non habes cor,qui habentes oculos non vident,et aures et non audiunt.
JER|5|22|Numquid me non timebitis,ait Dominus,et a facie mea non trepidabitis?Qui posui arenam terminum mari, praeceptum sempiternum, quod non praeteribit;et commovebuntur et non poterunt,et intumescent fluctus eius, et non transibunt illud ".
JER|5|23|Populo autem huic factum est cor contumax et rebelle;recesserunt et abierunt
JER|5|24|et non dixerunt in corde suo: Metuamus Dominum Deum nostrum,qui dat nobis pluviamtemporaneam et serotinam in tempore suo,hebdomadas statutas messiscustodientem nobis ".
JER|5|25|Iniquitates vestrae declinaverunt haec,et peccata vestra prohibuerunt bonum a vobis,
JER|5|26|quia inventi sunt in populo meo impii,insidiantes quasi incurvati aucupes,laqueos ponentes ad capiendos viros.
JER|5|27|Sicut decipula plena avibus,sic domus eorum plenae dolo;ideo magnificati sunt et ditati,
JER|5|28|incrassati sunt et impinguati:et transgressi sunt terminos mali.Causam non iudicaverunt,causam pupilli, ut ipsi prospere agant,et iudicium pauperum non iudicaverunt.
JER|5|29|Numquid super his non visitabo,dicit Dominus,aut super gentem huiuscemodinon ulciscetur anima mea?
JER|5|30|Stupor et mirabiliafacta sunt in terra:
JER|5|31|prophetae prophetabant mendacium,et sacerdotes applaudebant manibus suis,et populus meus dilexit talia.Quid igitur facietis in novissimo eius?
JER|6|1|Fugite, filii Beniamin,de medio Ierusalem;et in Thecua clangite bucinaet super Bethcharem levate vexillum,quia malum visum est ab aquiloneet contritio magna.
JER|6|2|Speciosam et delicatam silere fecifiliam Sion.
JER|6|3|Ad eam venient pastores et greges eorum,figent in ea tentoria in circuitu;pascet unusquisque partem suam.
JER|6|4|" Sanctificate super eam bellum,consurgite, et ascendamus in meridie;vae nobis, quia declinavit dies,quia longiores factae sunt umbrae vesperi!
JER|6|5|Surgite, et ascendamus in nocteet dissipemus domos eius ".
JER|6|6|Quia haec dicit Dominus exercituum: Caedite lignum eiuset fundite circa Ierusalem aggerem;haec est civitas visitationis,omnis calumnia in medio eius.
JER|6|7|Sicut effluere facit cisterna aquam suam,sic illa effluere facit malitiam suam;violentia et vastitas auditur in ea,coram me semper afflictio et plaga.
JER|6|8|Erudire, Ierusalem,ne forte recedat anima mea a te,ne forte ponam te desertam,terram inhabitabilem ".
JER|6|9|Haec dicit Dominus exercituum: Usque ad racemum colligent quasi in vineareliquias Israel.Converte manum tuamquasi vindemiator ad palmites ".
JER|6|10|Cui loquar et quem contestabor, ut audiat?Ecce incircumcisae aures eorum,et audire non possunt;ecce verbum Domini factum est eis in opprobrium,et non suscipient illud.
JER|6|11|Idcirco furore Domini plenus sum,laboravi sustinens. Effunde super parvulum foriset super concilium iuvenum simul;etiam vir cum muliere capietur,senex cum pleno dierum.
JER|6|12|Et transibunt domus eorum ad alteros,agri et uxores pariter,quia extendam manum meamsuper habitantes terram ",dicit Dominus.
JER|6|13|A minore quippe usque ad maioremomnes avaritiae student,et a propheta usque ad sacerdotemcuncti faciunt dolum.
JER|6|14|Et curant contritionem populi mei in levitatedicentes: " Pax, pax "; et non est pax.
JER|6|15|Confusi sunt, quia abominationem fecerunt;quin potius confusione non sunt confusiet erubescere nescierunt. Quam ob rem cadent inter ruentes;tempore, quo visitavero eos, corruent ",dicit Dominus.
JER|6|16|Haec dicit Dominus: State super vias et videteet interrogate de semitis antiquis,quae sit via bona, et ambulate in eaet invenietis refrigerium animabus vestris ".Et dixerunt: " Non ambulabimus! ".
JER|6|17|Et constitui super vos speculatores: Audite vocem tubae ".Et dixerunt: " Non audiemus! ".
JER|6|18|Ideo audite, gentes,et cognosce, congregatio,quanta ego faciam eis.
JER|6|19|Audi terra: " Ecce ego adducam mala super populum istum,fructum cogitationum eorum,quia verba mea non audieruntet legem meam proiecerunt.
JER|6|20|Ut quid mihi tus, quod de Saba venit,et calamus suave olens de terra longinqua?Holocautomata vestra non sunt accepta,et victimae vestrae non placent mihi ".
JER|6|21|Propterea haec dicit Dominus: Ecce ego dabo in populum istum offendicula,et offendent in eis patres et filii simul,vicinus et proximus peribunt ".
JER|6|22|Haec dicit Dominus: Ecce populus venit de terra aquilonis,et gens magna consurget a finibus terrae;
JER|6|23|arcum et acinacem arripiet,crudelis est et non miserebitur;vox eorum quasi mare sonabit,et super equos ascendent,praeparati quasi vir ad proeliumadversum te, filia Sion ".
JER|6|24|" Audivimus famam eius;dissolutae sunt manus nostrae,tribulatio apprehendit nos,dolores ut parturientem ".
JER|6|25|Nolite exire ad agroset in via ne ambuletis,quoniam gladius inimici,pavor in circuitu.
JER|6|26|Filia populi mei, accingere cilicioet volutare in cinere,luctum unigeniti fac tibi,planctum amarum,quia repente veniet vastator super nos.
JER|6|27|Probatorem dedi te in populo meo;et scies et probabis viam eorum.
JER|6|28|Omnes isti principes rebelles,ambulantes fraudulenter.Aes et ferrum,omnia isti corrumpunt.
JER|6|29|Sufflavit sufflatorium in igne,consumptum est plumbum;frustra conflavit conflator,scoriae enim non sunt separatae.
JER|6|30|Argentum reprobum vocate eos,quia Dominus proiecit illos.
JER|7|1|Verbum, quod factum est ad Ieremiam a Domino dicens:
JER|7|2|" Sta in porta domus Domini et praedica ibi verbum istud et dic: Audite verbum Domini, omnis Iuda, qui ingredimini per portas has, ut adoretis Dominum.
JER|7|3|Haec dicit Dominus exercituum, Deus Israel: Bonas facite vias vestras et opera vestra, et habitare vos faciam in loco isto.
JER|7|4|Nolite confidere in verbis mendacii dicentes: "Templum Domini, templum Domini, templum Domini est".
JER|7|5|Quoniam, si bene direxeritis vias vestras et opera vestra, si feceritis iudicium inter virum et proximum eius,
JER|7|6|advenae et pupillo et viduae non feceritis calumniam nec sanguinem innocentem effuderitis in loco hoc et post deos alienos non ambulaveritis in malum vobismetipsis,
JER|7|7|habitare vos faciam in loco isto, in terra, quam dedi patribus vestris a saeculo usque in saeculum.
JER|7|8|Ecce vos confiditis vobis in sermonibus mendacii, qui non proderunt.
JER|7|9|Quid? Furari, occidere, adulterari, iurare mendaciter, incensum offerre Baal et ire post deos alienos, quos ignoratis;
JER|7|10|et venitis et statis coram me in domo hac, super quam invocatum est nomen meum, et dicitis: "Liberati sumus", eo quod faciatis omnes abominationes istas.
JER|7|11|Numquid spelunca latronum facta est domus ista, super quam invocatum est nomen meum in oculis vestris?Ecce, etiam ego vidi, dicit Dominus.
JER|7|12|Ite ad locum meum in Silo, ubi habitavit nomen meum a principio, et videte, quae fecerim ei propter malitiam populi mei Israel.
JER|7|13|Et nunc, quia fecistis omnia opera haec, dicit Dominus, et locutus sum ad vos mane consurgens et loquens, et non audistis, et vocavi vos, et non respondistis,
JER|7|14|faciam domui huic, super quam invocatum est nomen meum, et in qua vos habetis fiduciam, et loco, quem dedi vobis et patribus vestris, sicut feci Silo;
JER|7|15|et proiciam vos a facie mea, sicut proieci omnes fratres vestros, universum semen Ephraim.
JER|7|16|Tu ergo, noli orare pro populo hoc nec assumas pro eis deprecationem et orationem et non obsistas mihi, quia non exaudiam te.
JER|7|17|Nonne vides, quid isti faciant in civitatibus Iudae et in plateis Ierusalem?
JER|7|18|Filii colligunt ligna, et patres succendunt ignem, et mulieres commiscent farinam, ut faciant placentas reginae caeli et libent diis alienis, ut me ad iracundiam provocent.
JER|7|19|Numquid me ad iracundiam provocant, dicit Dominus, nonne semetipsos in confusionem vultus sui?
JER|7|20|Ideo haec dicit Dominus Deus: Ecce furor meus et indignatio mea effunditur super locum istum, super homines et super iumenta et super lignum regionis et super fruges terrae et succendetur et non exstinguetur.
JER|7|21|Haec dicit Dominus exercituum, Deus Israel: Holocautomata vestra addite victimis vestris et comedite carnes,
JER|7|22|quia non sum locutus cum patribus vestris et non praecepi eis in die, qua eduxi eos de terra Aegypti, de verbo holocautomatum et victimarum.
JER|7|23|Sed hoc verbum praecepi eis dicens: Audite vocem meam, et ero vobis Deus, et vos eritis mihi populus; et ambulate in omni via, quam mandaverim vobis, ut bene sit vobis.
JER|7|24|Et non audierunt nec inclinaverunt aurem suam, sed abierunt in voluntatibus et in pravitate cordis sui mali factique sunt retrorsum et non in ante
JER|7|25|a die, qua egressi sunt patres eorum de terra Aegypti, usque ad diem hanc. Et misi ad vos omnes servos meos prophetas, per diem consurgens diluculo et mittens;
JER|7|26|et non audierunt me nec inclinaverunt aurem suam, sed induraverunt cervicem suam et peius operati sunt quam patres eorum.
JER|7|27|Et loqueris ad eos omnia verba haec, et non audient te; et vocabis eos, et non respondebunt tibi;
JER|7|28|et dices ad eos: Haec est gens, quae non audivit vocem Domini Dei sui nec recepit disciplinam. Periit fides et ablata est de ore eorum.
JER|7|29|Tonde capillum tuum et proiceet sume in collibus planctum,quia sprevit Dominuset proiecit generationem furoris sui.
JER|7|30|Quia fecerunt filii Iudae malum in oculis meis, dicit Dominus; posuerunt abominationes suas in domo, super quam invocatum est nomen meum, ut polluerent eam;
JER|7|31|et aedificaverunt excelsa Topheth, quae est in valle Benennom, ut incenderent filios suos et filias suas igni: quae non praecepi nec cogitavi in corde meo.
JER|7|32|Ideo ecce dies venient, dicit Dominus, et non dicetur amplius Topheth et vallis Benennom sed vallis Interfectionis; et sepelient in Topheth, eo quod non sit locus.
JER|7|33|Et erit morticinum populi huius in cibum volucribus caeli et bestiis terrae, et non erit qui abigat.
JER|7|34|Et quiescere faciam de urbibus Iudae et de plateis Ierusalem vocem gaudii et vocem laetitiae, vocem sponsi et vocem sponsae: in desolationem enim erit terra ".
JER|8|1|" In illo tempore, ait Dominus, eicient ossa regum Iudae et ossa principum eius et ossa sacerdotum et ossa prophetarum et ossa eorum, qui habitaverunt Ierusalem de sepulcris suis;
JER|8|2|et expandent ea ad solem et lunam et omnem militiam caeli, quae dilexerunt et quibus servierunt et post quae ambulaverunt et quae quaesierunt et adoraverunt; non colligentur et non sepelientur: in sterquilinium super faciem terrae erunt.
JER|8|3|Et eligent magis mortem quam vitam omnes, qui residui fuerint de cognatione hac pessima in universis locis, ad quae eiecero eos, dicit Dominus exercituum.
JER|8|4|Et dices ad eos: Haec dicit Dominus:Numquid, qui cadit, non resurget, et, qui aversus est, non revertetur?
JER|8|5|Quare ergo aversus est populus iste,Ierusalem aversione perpetua?Apprehenderunt mendaciumet noluerunt reverti.
JER|8|6|Attendi et auscultavi:nemo, quod bonum est, loquitur,nullus est, qui agat paenitentiamsuper malitia sua dicens:Quid feci?".Omnes conversi sunt ad cursum suum,quasi equus impetu vadens in proelio.
JER|8|7|Etiam ciconia in caelonovit tempus suum;turtur et hirundo et turduscustodierunt tempus adventus sui;populus autem meus non novitiudicium Domini.
JER|8|8|Quomodo dicitis: "Sapientes nos sumus,et lex Domini nobiscum est"?Vere mendacium operatus eststilus mendax scribarum.
JER|8|9|Confusi sunt sapientes,perterriti et capti sunt;verbum enim Domini proiecerunt,et sapientia nulla est in eis.
JER|8|10|Propterea dabo mulieres eorum exteris,agros eorum expugnatoribus,quia a minimo usque ad maximumomnes avaritiam sequuntur,a propheta usque ad sacerdotemcuncti faciunt mendacium.
JER|8|11|Et sanant contritionemfiliae populi mei in levitatedicentes "Pax, pax", cum non sit pax.
JER|8|12|Confusi sunt, quia abominationem fecerunt;quin immo confusione non sunt confusiet erubescere nescierunt,idcirco cadent inter corruentes,in tempore visitationis suae corruent,dicit Dominus.
JER|8|13|Congregans congregabo eos,ait Dominus;non est uva in vitibus,et non sunt ficus in ficulnea,folium defluxit,et dabo eis gradientes super eos.
JER|8|14|"Quare sedemus?Convenite, et ingrediamur civitates munitaset pereamus ibi,quia Dominus Deus noster tradidit nos in interitumet potum dedit nobis aquam fellis;peccavimus enim Domino.
JER|8|15|Exspectavimus pacem, et non est bonum,tempus medelae, et ecce formido".
JER|8|16|A Dan auditus est fremitus equorum eius,a voce hinnituum fortium equorum eiuscommota est omnis terra;et venient et devorabunt terram et plenitudinem eius,urbem et habitatores eius.
JER|8|17|Quia ecce ego mittam vobisserpentes regulos,quibus non est incantatio,et mordebunt vos ",ait Dominus.
JER|8|18|Hilaritas mea facta est dolor in me,cor meum maerens.
JER|8|19|Ecce vox clamoris filiae populi meide terra longinqua: Numquid Dominus non est in Sion?Aut rex eius non est in ea? ". Quare ergo me ad iracundiam concitaverunt in sculptilibus suiset in vanitatibus alienis? ".
JER|8|20|" Transiit messis, finita est aestas,et nos salvati non sumus ".
JER|8|21|Super contritione filiae populi meicontritus sum et contristatus;stupor obtinuit me.
JER|8|22|Numquid resina non est in Galaad?Aut medicus non est ibi?Quare enim non est obductacicatrix filiae populi mei?
JER|8|23|Quis dabit capiti meo aquamet oculis meis fontem lacrimarum,et plorabo die ac nocteinterfectos filiae populi mei?
JER|9|1|Quis dabit mihi in solitudine deversorium viatorum,et de relinquam populum meum et recedam ab eis?Quia omnes adulteri sunt,coetus praevaricatorum.
JER|9|2|" Et tenderunt linguam suam quasi arcum;mendacium, et non veritas, invaluit in terra,quia de malo ad malum egressi suntet me non cognoverunt,dicit Dominus.
JER|9|3|Unusquisque se a proximo suo custodiatet in omni fratre suo non habeat fiduciam,quia omnis frater supplantat,et omnis amicus fraudulenter incedit,
JER|9|4|et vir fratrem suum decipit,et veritatem non loquuntur;docuerunt enim linguam suam loqui mendacium,inique egerunt, noluerunt converti.
JER|9|5|Iniuria super iniuriam,dolus super dolum.Renuerunt scire me ",dicit Dominus.
JER|9|6|Propterea haec dicit Dominus exercituum: Ecce ego conflabo et probabo eos;quid enim aliud faciam filiae populi mei?
JER|9|7|Sagitta vulnerans lingua eorum;dolum locuta est in ore suo:pacem cum amico suo loquituret occulte ponit ei insidias.
JER|9|8|Numquid super his non visitabo eos,dicit Dominus,aut in gente huiusmodinon ulciscetur anima mea? ".
JER|9|9|Super montes assumam fletum ac lamentumet super pascua deserti planctum,quoniam incensa sunt,eo quod non sit vir pertransiens,et non audiunt vocem gregis;a volucre caeli usque ad pecoratransmigraverunt, recesserunt.
JER|9|10|" Et dabo Ierusalem in acervos arenaeet cubilia thoum,et civitates Iudae dabo in desolationem,eo quod non sit habitator ".
JER|9|11|Quis est vir sapiens, qui intellegat hoc,et ad quem verbum oris Domini fiat,ut annuntiet istud:Quare perierit terra,exusta sit quasi desertum,eo quod non sit qui pertranseat?
JER|9|12|Et dixit Dominus: " Quia dereliquerunt legem meam, quam dedi eis, et non audierunt vocem meam et non ambulaverunt in ea;
JER|9|13|et abierunt post pravitatem cordis sui et post Baalim, quos didicerunt a patribus suis ".
JER|9|14|Idcirco haec dicit Dominus exercituum, Deus Israel: " Ecce ego cibabo populum istum absinthio et potum dabo eis aquam fellis;
JER|9|15|et dispergam eos in gentibus, quas non noverunt ipsi et patres eorum, et mittam post eos gladium, donec consumantur.
JER|9|16|Haec dicit Dominus exercituum:Attendite et vocate lamentatrices, et veniant;et ad eas, quae sapientes sunt, mittite, et properent! ".
JER|9|17|Festinentet assumant super nos lamentum:deducant oculi nostri lacrimas,et palpebrae nostrae defluant aquis.
JER|9|18|Quia vox lamentationis audita est de Sion: Quomodo vastati sumus et confusi vehementer,quia dereliquimus terram,quoniam deiecta sunt tabernacula nostra ".
JER|9|19|Audite ergo, mulieres, verbum Domini;et assumant aures vestrae sermonem oris eius,et docete filias vestras lamentum,et unaquaeque proximam suam planctum.
JER|9|20|Quia ascendit mors per fenestras nostras,ingressa est domos nostras,disperdere parvulos deforis,iuvenes de plateis.
JER|9|21|Loquere. Haec dicit Dominus: Et cadet morticinum hominisquasi stercus super faciem regioniset quasi manipulus post tergum metentis,et non est qui colligat ".
JER|9|22|Haec dicit Dominus: Non glorietur sapiens in sapientia sua,et non glorietur fortis in fortitudine sua,et non glorietur dives in divitiis suis;
JER|9|23|sed in hoc glorietur, qui gloriatur:scire et nosse me,quia ego sum Dominus, qui facio misericordiamet iudicium et iustitiam in terra;haec enim placent mihi,ait Dominus.
JER|9|24|Ecce dies veniunt, dicit Dominus, et visitabo super omnem, qui circumcisum habet praeputium,
JER|9|25|super Aegyptum et super Iudam et super Edom et super filios Ammon et super Moab et super omnes, qui attonsi sunt in comam, habitantes in deserto, quia omnes gentes habent praeputium, omnis autem domus Israel incircumcisi sunt corde ".
JER|10|1|Audite verbum, quod locutus est Dominus super vos, domus Israel.
JER|10|2|Haec dicit Dominus: Iuxta vias gentium nolite discereet a signis caeli nolite metuere,quae timent gentes,
JER|10|3|quia leges populorum vanae sunt.Quia lignum de saltu praeciditopus manuum artificis in ascia,
JER|10|4|argento et auro decoravit illud,clavis et malleis firmavit,ut non moveatur;
JER|10|5|sicut formido in cucumerario suntet non loquentur,portantur, quia incedere non valent:nolite ergo timere ea,quia nec male possunt facere nec bene ".
JER|10|6|Non est similis tui, Domine;magnus es tu,et magnum nomen tuum in fortitudine.
JER|10|7|Quis non timebit te, o rex gentium?Te enim decet,quoniam inter cunctos sapientes gentiumet in universis regnis earum nullus est similis tui.
JER|10|8|Pariter insipientes et fatui sunt;doctrina vanitatis eorum lignum est.
JER|10|9|Argentum involutum, quod de Tharsis affertur,et aurum de Ophaz,opus artificis et manuum aurificis,hyacinthus et purpura indumentum eorum;opus artificum universa haec.
JER|10|10|Dominus autem Deus verus est,ipse Deus vivens et rex sempiternus;ab indignatione eius commovebitur terra,et non sustinebunt gentes comminationem eius.
JER|10|11|Sic ergo dicetis eis: " Dii, qui caelos et terram non fecerunt, pereant de terra et de his, quae sub caelis sunt ".
JER|10|12|Qui fecit terram in fortitudine sua,firmavit orbem in sapientia suaet prudentia sua extendit caelos.
JER|10|13|Ad vocem suam dat multitudinem aquarum in caeloet elevat nebulas ab extremitatibus terrae;fulgura in pluviam facitet educit ventum de thesauris suis.
JER|10|14|Stultus factus est omnis homo absque scientia;confusus est omnis artifex in sculptili,quoniam falsum est, quod conflavit,et non est spiritus in eis.
JER|10|15|Vana sunt et opus risu dignum;in tempore visitationis suae peribunt.
JER|10|16|Non est his similis pars Iacob:qui enim formavit omnia, ipse est,et Israel tribus hereditatis eius,Dominus exercituum nomen illi.
JER|10|17|Congrega de terra sarcinam tuam,quae habitas in obsidione,
JER|10|18|quia haec dicit Dominus: Ecce ego longe proiciam habitatores terrae in hac viceet tribulabo eos, ita ut inveniant me ".
JER|10|19|Vae mihi super contritione mea,pessima plaga mea!Ego autem dixi: Plane haec infirmitas mea est,et portabo illam ".
JER|10|20|Tabernaculum meum vastatum est, omnes funiculi mei dirupti sunt;filii mei exierunt a me et non subsistunt,non est qui extendat ultra tentorium meumet erigat pelles meas.
JER|10|21|Quia stulte egerunt pastoreset Dominum non quaesierunt;propterea non prosperati sunt,et omnis grex eorum dispersus est.
JER|10|22|Vox auditionis ecce venitet commotio magna de terra aquilonis,ut ponat civitates Iudae solitudinemet habitaculum thoum.
JER|10|23|" Scio, Domine, quia non est hominis via eius,nec viri est, ut ambulet et dirigat gressus suos.
JER|10|24|Corripe me, Domine,verumtamen in iudicio et non in furore tuo,ne forte ad nihilum redigas me ".
JER|10|25|Effunde indignationem tuam super gentes,quae non cognoverunt te,et super cognationes,quae nomen tuum non invocaverunt;quia comederunt Iacobet devoraverunt eumet consumpserunt illumet pascua eius dissipaverunt.
JER|11|1|Verbum, quod factum est ad Ieremiam a Domino dicens:
JER|11|2|" Audite verba pacti huius et loquimini ad viros Iudae et habitatores Ierusalem.
JER|11|3|Et dices ad eos: Haec dicit Dominus, Deus Israel: Maledictus vir, qui non audierit verba pacti huius,
JER|11|4|quod praecepi patribus vestris in die, qua eduxi eos de terra Aegypti, de fornace ferrea, dicens: Audite vocem meam et facite omnia, quae praecipio vobis, et eritis mihi in populum, et ego ero vobis in Deum;
JER|11|5|ut suscitem iuramentum, quod iuravi patribus vestris, daturum me eis terram fluentem lacte et melle, sicut est dies haec ". Et respondi et dixi: " Amen, Domine ".
JER|11|6|Et dixit Dominus ad me: " Vociferare omnia verba haec in civitatibus Iudae et in foris Ierusalem dicens: Audite verba pacti huius et facite illa.
JER|11|7|Quia contestans contestatus sum patres vestros in die, qua eduxi eos de terra Aegypti, usque ad diem hanc; mane consurgens contestatus sum et dixi: Audite vocem meam.
JER|11|8|Et non audierunt nec inclinaverunt aurem suam, sed abierunt unusquisque in pravitate cordis sui mali; et induxi super eos omnia verba pacti huius, quod praecepi, ut facerent, et non fecerunt ".
JER|11|9|Et dixit Dominus ad me: " Inventa est coniuratio in viris Iudae et in habitatoribus Ierusalem.
JER|11|10|Reversi sunt ad iniquitates patrum suorum priorum, qui noluerunt audire verba mea; et hi ergo abierunt post deos alienos, ut servirent eis: irritum fecerunt domus Israel et domus Iudae pactum meum, quod pepigi cum patribus eorum.
JER|11|11|Quam ob rem haec dicit Dominus: Ecce ego inducam super eos mala, de quibus exire non poterunt; et clamabunt ad me, et non exaudiam eos.
JER|11|12|Et ibunt civitates Iudae et habitatores Ierusalem et clamabunt ad deos, quibus sacrificant, et non salvabunt eos in tempore afflictionis eorum.
JER|11|13|Secundum numerum enim civitatum tuarum erant dii tui, Iuda, et secundum numerum viarum Ierusalem posuistis aras confusioni, aras ad sacrificandum Baal.
JER|11|14|Tu ergo noli orare pro populo hoc et ne assumas pro eis deprecationem et orationem, quia non exaudiam in tempore clamoris eorum ad me, in tempore afflictionis eorum.
JER|11|15|Quid est dilectae meae,ut in domo mea perficiat consilia mala?Numquid vota et carnes sanctaeauferent a te malitias tuas,in quibus glorieris? ".
JER|11|16|Olivam uberem, pulchram, fructibus speciosam,vocabit Dominus nomen tuum;ad vocem strepitus grandissuccendit ignem in ea,et combusti sunt rami eius.
JER|11|17|Et Dominus exercituum, qui plantavit te, locutus est super te malum, pro malis domus Israel et domus Iudae, quae fecerunt sibi ad irritandum me, sacrificantes Baal.
JER|11|18|Tu autem, Domine, demonstrasti mihi, et cognovi;tunc ostendisti mihi opera eorum.
JER|11|19|Et ego quasi agnus mansuetus, qui portatur ad victimam; et non cognovi quia super me cogitaverunt consilia: " Caedamus lignum in vigore eius et eradamus eum de terra viventium, et nomen eius non memoretur amplius ".
JER|11|20|Tu autem, Domine exercituum,qui iudicas iuste et probas renes et corda:videam ultionem tuam ex eis;tibi enim revelavi causam meam.
JER|11|21|Propterea haec dicit Dominus super viros Anathoth, qui quaerunt animam tuam et dicunt: " Non prophetabis in nomine Domini et non morieris in manibus nostris ".
JER|11|22|Propterea haec dicit Dominus exercituum: " Ecce ego visitabo super eos: iuvenes morientur in gladio, filii eorum et filiae eorum morientur in fame,
JER|11|23|et reliquiae non erunt eis; inducam enim malum super viros Anathoth, annum visitationis eorum ".
JER|12|1|Iustus quidem tu es, Domine, si disputem tecum;verumtamen de iudiciis loquar ad te.Quare via impiorum prosperatur?Bene est omnibus, qui praevaricantur et inique agunt.
JER|12|2|Plantasti eos, et radicem miserunt,proficiunt et faciunt fructum;prope es tu ori eorumet longe a renibus eorum.
JER|12|3|Et tu, Domine, nosti me, vidisti meet probasti cor meum tecum;segrega eos quasi gregem ad victimamet sanctifica eos in diem occisionis.
JER|12|4|Usquequo lugebit terra,et herba omnis regionis siccabiturpropter malitiam habitantium in ea?Consumptum est animal et volucre,quoniam dixerunt: "Non videbit novissima nostra".
JER|12|5|" Si cum peditibus currens laborasti,quomodo contendere poteris cum equis?Cum autem in terra pacis securus fueris,quid facies in silva condensa Iordanis?
JER|12|6|Nam et fratres tui et domus patris tui,etiam ipsi fraudulenter egerunt adversum teet clamaverunt post te plena voce;ne credas eis, cum locuti fuerint tibi bona ".
JER|12|7|" Reliqui domum meam,dimisi hereditatem meam;dedi dilectam animae meaein manu inimicorum eius.
JER|12|8|Facta est mihi hereditas meaquasi leo in silva;dedit contra me vocem, ideo odivi eam.
JER|12|9|Numquid avis discolor hereditas mea mihi?Numquid aves in circuitu contra eam?Venite, congregamini, omnes bestiae campi,properate ad devorandum.
JER|12|10|Pastores multi demoliti sunt vineam meam,conculcaverunt partem meam;dederunt portionem meam desiderabilemin desertum solitudinis.
JER|12|11|Posuerunt eam in dissipationem;lugetque coram me desolata,vastata est omnis terra,quia nullus est qui recogitet corde ".
JER|12|12|Super omnes colles in deserto venerunt vastatores,quia gladius Domini devoratab extremo terrae usque ad extremum eius;non est pax universae carni.
JER|12|13|Seminaverunt triticum et spinas messuerunt,laboraverunt, et non eis proderit;confundemini a fructibus vestrispropter iram furoris Domini.
JER|12|14|Haec dicit Dominus adversum omnes vicinos meos pessimos, qui tangunt hereditatem, quam distribui populo meo Israel: "Ecce ego evellam eos de terra sua et domum Iudae evellam de medio eorum.
JER|12|15|Et erit: cum evulsero eos, convertar et miserebor eorum et reducam eos, virum ad hereditatem suam et virum in terram suam.
JER|12|16|Et erit: si eruditi didicerint vias populi mei, ut iurent in nomine meo: "Vivit Dominus!", sicut docuerunt populum meum iurare in Baal, aedificabuntur in medio populi mei.
JER|12|17|Quod si non audierint, evellam gentem illam evulsione et perditione ", ait Dominus.
JER|13|1|Haec dixit Dominus ad me: " Vade et posside tibi lumba re lineum et pones illud super lumbos tuos et in aquam non inferes illud ".
JER|13|2|Et possedi lumbare iuxta verbum Domini et posui circa lumbos meos.
JER|13|3|Et factus est sermo Domini ad me secundo dicens:
JER|13|4|" Tolle lumbare, quod possedisti, quod est circa lumbos tuos, et surgens vade ad Euphraten et absconde ibi illud in foramine petrae ".
JER|13|5|Et abii et abscondi illud ad Euphraten, sicut praeceperat mihi Dominus.
JER|13|6|Et factum est, post dies plurimos dixit Dominus ad me: " Surge, vade ad Euphraten et tolle inde lumbare, quod praecepi tibi, ut absconderes ibi ".
JER|13|7|Et abii ad Euphraten et fodi et tuli lumbare de loco, ubi absconderam illud; et ecce, computruerat lumbare, ita ut nulli usui aptum esset.
JER|13|8|Et factum est verbum Domini ad me dicens:
JER|13|9|" Haec dicit Dominus: Sic putrescere faciam superbiam Iudae et superbiam Ierusalem multam;
JER|13|10|populus iste pessimus - qui nolunt audire verba mea et ambulant in pravitate cordis sui abieruntque post deos alienos, ut servirent eis et adorarent eos - erit sicut lumbare istud, quod nulli usui aptum est.
JER|13|11|Sicut enim adhaeret lumbare ad lumbos viri, sic agglutinavi mihi omnem domum Israel et omnem domum Iudae, dicit Dominus, ut esset mihi in populum et in nomen et in laudem et in gloriam, et non audierunt.
JER|13|12|Dices ergo ad eos sermonem istum: Haec dicit Dominus, Deus Israel: Omnis laguncula implebitur vino. Et dicent ad te: "Numquid ignoramus quia omnis laguncula implebitur vino?".
JER|13|13|Et dices ad eos: Haec dicit Dominus: Ecce ego implebo omnes habitatores terrae huius et reges, qui sedent de stirpe David super thronum eius, et sacerdotes et prophetas et omnes habitatores Ierusalem ebrietate;
JER|13|14|et collidam eos, virum in fratrem suum et patres et filios pariter, ait Dominus; non parcam et non concedam neque miserebor, ut non disperdam eos.
JER|13|15|Audite et auribus percipite; nolite elevari,quia Dominus locutus est.
JER|13|16|Date Domino Deo vestro gloriam,antequam contenebrescat,et antequam offendant pedes vestriad montes caliginosos;exspectabitis lucem,et ponet eam in umbram mortiset in caliginem.
JER|13|17|Quod si hoc non audieritis,in abscondito plorabit anima meaa facie superbiae;plorans plorabitet deducet oculus meus lacrimam,quia captus est grex Domini.
JER|13|18|" Dic regi et dominatrici:In humo sedete,quoniam descendit de capite vestrocorona gloriae vestrae.
JER|13|19|Civitates austri clausae sunt,et non est qui aperiat;translata est omnis Iudatransmigratione perfecta.
JER|13|20|Leva oculos tuos et videvenientes ab aquilone:Ubi est grex, qui datus est tibi,pecus inclitum tuum?
JER|13|21|Quid dices, cum visitaverit te?Tu enim ipsa docuisti eos adversum te,amicos in caput tuum;numquid non dolores apprehendent tequasi mulierem parturientem?
JER|13|22|Quod si dixeris in corde tuo:Quare venerunt mihi haec?".Propter multitudinem iniquitatis tuaerevelatae sunt laciniae tuae,pollutae sunt plantae tuae.
JER|13|23|Numquid mutare potest Aethiops pellem suamaut pardus varietates suas?Tunc et vos poteritis benefacere,cum didiceritis malum.
JER|13|24|Et disseminabo eos quasi stipulam,quae raptatur in vento deserti.
JER|13|25|Haec sors tua parsque mensurae tuae a me,dicit Dominus,quia oblita es meiet confisa es in mendacio.
JER|13|26|Unde et ego sublevabo lacinias tuas super faciem tuam,et apparebit ignominia tua,
JER|13|27|adulteria tua et hinnitus tuus,scelus fornicationis tuae.Super colles in agro vidi abominationes tuas.Vae tibi, Ierusalem! Non mundaberis;usquequo adhuc? ".
JER|14|1|Quod factum est verbum Domini ad Ieremiam de sic citate.
JER|14|2|Luget Iuda,et portae eius languescuntet contristatae iacent in terra,et clamor Ierusalem ascendit.
JER|14|3|Maiores eorum miserunt minores suos ad aquam:venerunt ad cisternas,non invenerunt aquam;reportaverunt vasa sua vacua,confusi sunt et afflictiet operuerunt capita sua.
JER|14|4|Propter terrae vastitatem,quia non venit pluvia in terram,confusi sunt agricolae,operuerunt capita sua.
JER|14|5|Nam et cerva in agro peperit et reliquit,quia non erat herba.
JER|14|6|Et onagri steterunt in collibus,traxerunt aerem quasi thoes;defecerunt oculi eorum,quia non erat herba.
JER|14|7|" Si iniquitates nostrae testificantur adversus nos,Domine, fac propter nomen tuum,quoniam multae sunt aversiones nostrae,tibi peccavimus.
JER|14|8|Exspectatio Israel,salvator eius in tempore tribulationis,quare quasi peregrinus es in terraet quasi viator declinans ad pernoctandum?
JER|14|9|Quare es velut vir attonitus,ut fortis, qui non potest salvare?Tu autem in medio nostri es, Domine,et nomen tuum invocatum est super nos;ne derelinquas nos ".
JER|14|10|Haec dicit Dominus populo huic: " Ita diligunt vagari, pedes suos non prohibent et Domino non placent ". Nunc recordatus est iniquitatum eorum et visitat peccata eorum.
JER|14|11|Et dixit Dominus ad me: " Noli orare pro populo isto in bonum.
JER|14|12|Cum ieiunaverint, non exaudiam preces eorum; et, si obtulerint holocautomata et oblationes, non suscipiam ea; quoniam gladio et fame et peste consumam eos ".
JER|14|13|Et dixi: " Heu, Domine Deus! Ecce prophetae dicunt eis: "Non videbitis gladium, et fames non erit in vobis, sed pacem veram dabit vobis in loco isto" ".
JER|14|14|Et dixit Dominus ad me: " Falso prophetae vaticinantur in nomine meo: non misi eos et non praecepi eis neque locutus sum ad eos; visionem mendacem et divinationem et fraudulentiam et seductionem cordis sui prophetant vobis.
JER|14|15|Idcirco haec dicit Dominus contra prophetas, qui prophetant in nomine meo, quos ego non misi, dicentes: "Gladius et fames non erit in terra hac": In gladio et fame consumentur prophetae illi;
JER|14|16|et homines, quibus prophetant, erunt proiecti in viis Ierusalem prae fame et gladio, et non erit qui sepeliat eos: ipsi et uxores eorum, filii et filiae eorum, et effundam super eos malum suum.
JER|14|17|Et dices ad eos verbum istud:Deducant oculi mei lacrimamper noctem et diem, et non taceant,quoniam contritione magna contrita estvirgo filia populi mei,plaga pessima vehementer.
JER|14|18|Si egressus fuero ad agros,ecce occisi gladio;et, si introiero in civitatem,ecce attenuati fame;propheta quoque et sacerdosabierunt per terram nescientes ".
JER|14|19|Numquid proiciens abiecisti Iudam,aut Sion abominata est anima tua?Quare ergo percussisti nos,ita ut nulla sit sanitas?Exspectavimus pacem, et non est bonum,et tempus curationis, et ecce turbatio.
JER|14|20|Cognovimus, Domine, impietates nostras,iniquitates patrum nostrorum, quia peccavimus tibi.
JER|14|21|Ne des nos in opprobrium propter nomen tuum,ne facias contumeliam solio gloriae tuae;recordare, ne irritum facias foedus tuum nobiscum.
JER|14|22|Numquid sunt in sculptilibus gentium, qui pluant,aut caeli possunt dare imbres?Nonne tu es Dominus Deus noster,quem exspectamus?Tu enim fecisti omnia haec.
JER|15|1|Et dixit Dominus ad me: " Si steterit Moyses et Samuel co ram me, non est anima mea ad populum istum; eice illos a facie mea, et egrediantur.
JER|15|2|Quod si dixerint ad te: "Quo egrediemur?", dices ad eos: Haec dicit Dominus:Qui ad mortem, ad mortem;et qui ad gladium, ad gladium;et qui ad famem, ad famem;et qui ad captivitatem, ad captivitatem.
JER|15|3|Et mandabo super eos quattuor species, dicit Dominus: gladium ad occisionem et canes ad lacerandum et volatilia caeli et bestias terrae ad devorandum et dissipandum.
JER|15|4|Et dabo eos in commotionem universis regnis terrae, propter Manassem filium Ezechiae regem Iudae, super omnibus, quae fecit in Ierusalem.
JER|15|5|Quis enim miserebitur tui, Ierusalem,aut quis contristabitur pro te,aut quis ibit ad rogandum de pace tua?
JER|15|6|Tu reppulisti me,dicit Dominus,retrorsum abiisti;et extendi manum meam super te et interfeci te:laboravi miserans.
JER|15|7|Et ventilavi eos ventilabroin portis terrae;orbavi et disperdidi populum meum:a viis suis non sunt reversi.
JER|15|8|Multiplicatae sunt mihi viduae eiussuper arenam maris,induxi eis super matremmilitem vastatorem meridie,misi super eam repenteperturbationem et terrorem.
JER|15|9|Infirmata est, quae peperit septem,exhalavit animam suam;occidit ei sol, cum adhuc esset dies,confusa est et erubuit,et residuos eorum in gladium daboin conspectu inimicorum eorum ",ait Dominus.
JER|15|10|Vae mihi, mater mea,quoniam genuisti me virum rixaeet virum discordiae in universa terra!Non feneravi, nec feneravit mihi quisquam;omnes maledicunt mihi.
JER|15|11|Amen, Domine, ministravi tibi in bonum,intercessi apud te in tempore afflictioniset in tempore tribulationis pro inimico.
JER|15|12|Numquid frangitur ferroferrum aquilonis et aes?
JER|15|13|" Divitias tuas et thesauros tuosin direptionem dabo gratis,propter omnia peccata tua,in omnibus terminis tuis.
JER|15|14|Et servire te faciam inimicis tuisin terra, quam nescis,quia ignis succensus est in furore meo:super vos ardebit ".
JER|15|15|Tu scis, Domine;recordare mei et visita meet vindica me de his, qui persequuntur me;noli in patientia tua abripere me,scito quoniam sustinui pro te opprobrium.
JER|15|16|Inventi sunt sermones tui, et comedi eos,et factum est mihi verbum tuumin gaudium et in laetitiam cordis mei,quoniam invocatum est nomen tuum super me,Domine, Deus exercituum.
JER|15|17|Non sedi in concilio ludentiumet gloriatus sum;a facie manus tuae solus sedebam,quoniam indignatione replesti me.
JER|15|18|Quare factus est dolor meus perpetuus,et plaga mea desperabilis renuit curari?Factus es mihi quasi rivus mendax,aquae infideles.
JER|15|19|Propter hoc haec dixit Dominus: Si converteris, convertam te,et ante faciem meam stabis;et si separaveris pretiosum a vili,quasi os meum eris;convertentur ipsi ad te,et tu non converteris ad eos.
JER|15|20|Et dabo te populo huicin murum aereum fortem;et bellabunt adversum teet non praevalebunt,quia ego tecum sum,ut salvem te et eruam te,dicit Dominus.
JER|15|21|Et liberabo te de manu pessimorumet redimam te de manu fortium ".
JER|16|1|Et factum est verbum Domi ni ad me dicens:
JER|16|2|" Non acci pies uxorem, et non erunt tibi filii et filiae in loco isto.
JER|16|3|Quia haec dicit Dominus super filios et filias, qui generantur in loco isto, et super matres eorum, quae genuerunt eos, et super patres eorum, de quorum stirpe sunt nati in terra hac:
JER|16|4|Mortibus aegrotationum morientur, non plangentur et non sepelientur; in sterquilinium super faciem terrae erunt et gladio et fame consumentur, et erit cadaver eorum in escam volatilibus caeli et bestiis terrae ".
JER|16|5|Haec enim dixit Dominus: "Ne ingrediaris domum convivii neque vadas ad plangendum neque lugebis eos, quia abstuli pacem meam a populo isto, dicit Dominus, misericordiam et miserationes.
JER|16|6|Et morientur grandes et parvi in terra ista, non sepelientur neque plangentur, et non se incident, neque calvitium fiet pro eis.
JER|16|7|Et non frangent lugenti panem ad consolandum super mortuo et non dabunt ei calicem ad consolandum super patre suo et matre.
JER|16|8|Et domum convivii non ingredieris, ut sedeas cum eis et comedas et bibas.
JER|16|9|Quia haec dicit Dominus exercituum, Deus Israel: Ecce ego auferam de loco isto in oculis vestris et in diebus vestris vocem gaudii et vocem laetitiae, vocem sponsi et vocem sponsae.
JER|16|10|Et cum annuntiaveris populo huic omnia verba haec, et dixerint tibi: Quare locutus est Dominus super nos omne malum grande istud? Quae iniquitas nostra et quod peccatum nostrum, quod peccavimus Domino Deo nostro?",
JER|16|11|dices ad eos: Quia dereliquerunt me patres vestri, ait Dominus, et abierunt post deos alienos et servierunt eis et adoraverunt eos et me dereliquerunt et legem meam non custodierunt.
JER|16|12|Sed et vos peius operati estis quam patres vestri: ecce enim ambulat unusquisque post pravitatem cordis sui mali, ut me non audiat.
JER|16|13|Et eiciam vos de terra hac in terram, quam ignoratis, vos et patres vestri; et servietis ibi diis alienis, die ac nocte, quia non dabo vobis gratiam.
JER|16|14|Propterea ecce dies veniunt, dicit Dominus, et non dicetur ultra: Vivit Dominus, qui eduxit filios Israel de terra Aegypti!",
JER|16|15|sed: "Vivit Dominus, qui eduxit filios Israel de terra aquilonis et de universis terris, ad quas eieci eos!". Et reducam eos in terram suam, quam dedi patribus eorum.
JER|16|16|Ecce ego mittam piscatores multos, dicit Dominus, et piscabuntur eos; et post haec mittam eis multos venatores, et venabuntur eos de omni monte et de omni colle et de cavernis petrarum.
JER|16|17|Quia oculi mei super omnes vias eorum: non sunt absconditae a facie mea, et non est occulta iniquitas eorum ab oculis meis.
JER|16|18|Et reddam primum dupliciter iniquitates et peccata eorum, quia contaminaverunt terram meam in morticinis idolorum suorum et abominationibus suis impleverunt hereditatem meam ".
JER|16|19|Domine, fortitudo mea et praesidium meumet refugium meum in die tribulationis;ad te gentes venient ab extremis terrae et dicent: Vere mendacium possederunt patres nostri,vanitatem, quae nihil prodest ".
JER|16|20|Numquid faciet sibi homo deos,et ipsi non sunt dii?
JER|16|21|" Idcirco ecce ego ostendam eis per vicem hanc,ostendam eis manum meam et virtutem meam,et scient quia nomen mihi Dominus ".
JER|17|1|Peccatum Iudae scriptum est stilo ferreo,in ungue adamantino exaratumsuper tabulam cordis eorumet in cornibus ararum eorum,
JER|17|2|ut recordarentur filii eorum ararum suarumet palorum suorum iuxta ligna frondentiain collibus excelsis,
JER|17|3|montibus in campo. Divitias tuas, omnes thesauros tuosin direptionem dabo,excelsa tua propter peccatain universis finibus tuis.
JER|17|4|Et relinques hereditatem tuam,quam dedi tibi;et servire te faciam inimicis tuisin terra, quam ignoras,quoniam ignem succendistis in naribus meis;usque in aeternum ardebit ".
JER|17|5|Haec dicit Dominus: Maledictus homo, qui confidit in homineet ponit carnem brachium suum,et a Domino recedit cor eius;
JER|17|6|erit enim quasi myricae in desertoet non videbit, cum venerit bonum,sed habitabit in siccitate in deserto,in terra salsuginis et inhabitabili.
JER|17|7|Benedictus vir, qui confidit in Domino,et erit Dominus fiducia eius;
JER|17|8|et erit quasi lignum,quod transplantatur super aquas,quod ad humorem mittit radices suaset non timebit, cum venerit aestus;et erit folium eius viride,et in anno siccitatis non erit sollicitumnec aliquando desinet facere fructum
JER|17|9|Dolosum est cor super omnia et insanabile;quis cognoscet illud?
JER|17|10|Ego Dominus scrutans cor et probans renes,qui do unicuique iuxta viam suamet iuxta fructum operum suorum.
JER|17|11|Perdix fovit, quae non peperit,ita faciens divitias sed non in iudicio.In dimidio dierum suorum derelinquet easet in novissimo suo erit insipiens ".
JER|17|12|Solium gloriae, altitudo a principio,locus sanctificationis nostrae!
JER|17|13|Exspectatio Israel, Domine,omnes, qui te derelinquunt, confundentur;recedentes a te in terra scribentur,quoniam dereliquerunt venamaquarum viventium, Dominum.
JER|17|14|Sana me, Domine, et sanabor;salvum me fac, et salvus ero,quoniam laus mea tu es.
JER|17|15|Ecce ipsi dicunt ad me: Ubi est verbum Domini? Veniat ".
JER|17|16|Et ego non institi pro malo apud teet diem calamitatis non desideravi,tu scis: quod egressum est de labiis meis,rectum in conspectu tuo fuit.
JER|17|17|Non sis mihi tu formidini;refugium meum tu in die afflictionis.
JER|17|18|Confundantur, qui me persequuntur,et non confundar ego;paveant illi, et non paveam ego;induc super eos diem afflictioniset duplici contritione contere eos.
JER|17|19|Haec dixit Dominus ad me: " Vade et sta in porta Filiorum populi, per quam ingrediuntur reges Iudae et egrediuntur, et in cunctis portis Ierusalem;
JER|17|20|et dices ad eos: Audite verbum Domini, reges Iudae et omnis Iuda cunctique habitatores Ierusalem, qui ingredimini per portas istas.
JER|17|21|Haec dicit Dominus: Custodite animas vestras et nolite portare pondera in die sabbati nec inferatis per portas Ierusalem;
JER|17|22|et nolite efferre onera de domibus vestris in die sabbati et omne opus non facietis: sanctificate diem sabbati, sicut praecepi patribus vestris.
JER|17|23|Et non audierunt nec inclinaverunt aurem suam; sed induraverunt cervicem suam, ne audirent me et ne acciperent disciplinam.
JER|17|24|Et erit: si audieritis me, dicit Dominus, ut non inferatis onera per portas civitatis huius in die sabbati, et si sanctificaveritis diem sabbati, ne faciatis in eo omne opus,
JER|17|25|ingredientur per portas civitatis huius reges et principes sedentes super solium David et ascendentes in curribus et equis, ipsi et principes eorum, viri Iudae et habitatores Ierusalem; et habitabitur civitas haec in sempiternum.
JER|17|26|Et venient de civitatibus Iudae et de circuitu Ierusalem et de terra Beniamin et de Sephela et de montuosis et a Nageb, portantes holocaustum et victimam et sacrificium et tus, et inferent oblationem laudis in domum Domini.
JER|17|27|Si autem non audieritis me, ut sanctificetis diem sabbati et ne portetis onus intrantes per portas Ierusalem in die sabbati, succendam ignem in portis eius, et devorabit domos Ierusalem et non exstinguetur ".
JER|18|1|Verbum, quod factum est ad Ieremiam a Domino dicens:
JER|18|2|" Surge et descende in domum figuli et ibi audies verba mea ".
JER|18|3|Et descendi in domum figuli, et ecce ipse faciebat opus super rotam;
JER|18|4|et dissipatum est vas, quod ipse faciebat e luto manibus suis, et rursus fecit illud vas alterum, sicut placuerat in oculis eius, ut faceret.
JER|18|5|Et factum est verbum Domini ad me dicens:
JER|18|6|" Numquid sicut figulus iste non potero vobis facere, domus Israel?, ait Dominus. Ecce, sicut lutum in manu figuli, sic vos in manu mea, domus Israel.
JER|18|7|Repente loquar adversum gentem et adversum regnum, ut eradicem et destruam et disperdam illud;
JER|18|8|si paenitentiam egerit gens illa a malo suo, propter quod locutus sum adversus eam, agam et ego paenitentiam super malo, quod cogitavi ut facerem ei.
JER|18|9|Et subito loquar de gente et de regno, ut aedificem et plantem illud;
JER|18|10|si fecerit malum in oculis meis, ut non audiat vocem meam, paenitentiam agam super bono, quod locutus sum ut facerem ei.
JER|18|11|Nunc ergo, dic viro Iudae et habitatoribus Ierusalem dicens: Haec dicit Dominus: Ecce ego fingo contra vos malum et cogito contra vos cogitationem; revertatur unusquisque a via sua mala, et dirigite vias vestras et opera vestra ".
JER|18|12|Qui dixerunt: " Vanum est; post cogitationes enim nostras ibimus et unusquisque pravitatem cordis sui mali faciemus ".
JER|18|13|Ideo haec dicit Dominus: Interrogate gentes:quis audivit talia horribilia,quae fecit nimis virgo Israel?
JER|18|14|Numquid deficiet de petra agrinix Libani,aut arescent aquae erumpentesfrigidae et defluentes?
JER|18|15|Quia oblitus est mei populus meus,vanitati sacrificanteset impingentes in viis suis,in semitis antiquis,ut ambularent per callesin itinere non trito,
JER|18|16|ut poneret terram eorum in desolationemet in sibilum sempiternum:omnis, qui praeterierit per eam, obstupescetet movebit caput suum.
JER|18|17|Sicut ventus urens dispergam eoscoram inimico;dorsum et non faciem ostendam eis in die perditionis eorum ".
JER|18|18|Et dixerunt: " Venite, et cogitemus contra Ieremiam cogitationes; non enim peribit lex a sacerdote, neque consilium a sapiente, nec sermo a propheta. Venite, et percutiamus eum lingua et non attendamus ad universos sermones eius ".
JER|18|19|Attende, Domine, ad meet audi vocem adversariorum meorum.
JER|18|20|Numquid redditur pro bono malum,quia foderunt foveam animae meae?Recordare quod steterim in conspectu tuo,ut loquerer pro eis bonumet averterem indignationem tuam ab eis.
JER|18|21|Propterea da filios eorum in famemet deduc eos in manus gladii;fiant uxores eorum absque liberis et viduae,et viri eorum interficiantur morte,iuvenes eorum confodiantur gladio in proelio.
JER|18|22|Audiatur clamor de domibus eorum;adduces enim super eos latronem repente,quia foderunt foveam, ut caperent me,et laqueos absconderunt pedibus meis.
JER|18|23|Tu autem, Domine, scis omne consilium eorumadversum me in mortem;ne propitieris iniquitati eorum,et peccatum eorum a facie tua non deleatur.Fiant corruentes in conspectu tuo;in tempore furoris tui abutere eis.
JER|19|1|Haec dicit Dominus: " Vade et eme lagunculam figuli testeam et accipe de senioribus populi et de senioribus sacerdotum
JER|19|2|et egredere ad vallem Benennom, quae est iuxta introitum portae Fictilium, et praedicabis ibi verba, quae ego loquar ad te,
JER|19|3|et dices: Audite verbum Domini, reges Iudae et habitatores Ierusalem: Haec dicit Dominus exercituum, Deus Israel: Ecce ego inducam afflictionem super locum istum, ita ut omnis, qui audierit illam, tinniant aures eius,
JER|19|4|eo quod dereliquerint me et alienum fecerint locum istum et sacrificaverint in eo diis alienis, quos nescierunt ipsi et patres eorum et reges Iudae; et repleverunt locum istum sanguine innocentium;
JER|19|5|et aedificaverunt excelsa Baal ad comburendos filios suos igne in holocaustum Baal: quae non praecepi nec locutus sum, nec ascenderunt in cor meum.
JER|19|6|Propterea ecce dies veniunt, dicit Dominus, et non vocabitur amplius locus iste Topheth et vallis Benennom sed vallis Occisionis.
JER|19|7|Et dissipabo consilium Iudae et Ierusalem in loco isto; et subvertam eos gladio in conspectu inimicorum suorum et in manu quaerentium animas eorum et dabo cadavera eorum escam volatilibus caeli et bestiis terrae.
JER|19|8|Et ponam civitatem hanc in stuporem et in sibilum; omnis, qui praeterierit per eam, obstupescet et sibilabit super universa plaga eius.
JER|19|9|Et cibabo eos carnibus filiorum suorum et carnibus filiarum suarum; et unusquisque carnem amici sui comedet in obsidione et in angustia, in qua concludent eos inimici eorum et qui quaerunt animas eorum.
JER|19|10|Et conteres lagunculam in oculis virorum, qui ibunt tecum,
JER|19|11|et dices ad eos: Haec dicit Dominus exercituum: Sic conteram populum istum et civitatem istam, sicut conteritur vas figuli, quod non potest ultra instaurari; et in Topheth sepelientur, eo quod non sit alius locus ad sepeliendum.
JER|19|12|Sic faciam loco huic, ait Dominus, et habitatoribus eius, ut ponam civitatem istam sicut Topheth;
JER|19|13|et erunt domus Ierusalem et domus regum Iudae sicut locus Topheth, immundae: omnes domus, in quarum domatibus sacrificaverunt omni militiae caeli et libaverunt libamina diis alienis ".
JER|19|14|Venit autem Ieremias de Topheth, quo miserat eum Dominus ad prophetandum, et stetit in atrio domus Domini et dixit ad omnem populum:
JER|19|15|" Haec dicit Dominus exercituum, Deus Israel: Ecce ego inducam super civitatem hanc et super omnes urbes eius universa mala, quae locutus sum adversum eam, quoniam induraverunt cervicem suam, ut non audirent sermones meos ".
JER|20|1|Et audivit Phassur filius Em mer sacerdos, qui constitutus erat princeps in domo Domini, Ieremiam prophetantem sermones istos;
JER|20|2|et percussit Phassur Ieremiam prophetam et misit eum in nervum, quod erat in porta Beniamin superiore in domo Domini.
JER|20|3|Cumque illuxisset in crastinum, eduxit Phassur Ieremiam de nervo; et dixit ad eum Ieremias: " Non Phassur vocavit Dominus nomen tuum sed Pavorem undique.
JER|20|4|Quia haec dicit Dominus: Ecce ego dabo te in pavorem, te et omnes amicos tuos, et corruent gladio inimicorum suorum, et oculi tui videbunt; et omnem Iudam dabo in manu regis Babylonis, et traducet eos in Babylonem et percutiet eos gladio.
JER|20|5|Et dabo universam substantiam civitatis huius et omnem laborem eius omneque pretium et cunctos thesauros regum Iudae dabo in manu inimicorum eorum; et diripient eos et tollent et ducent in Babylonem.
JER|20|6|Tu autem, Phassur et omnes habitatores domus tuae, ibitis in captivitatem; et in Babylonem venies et ibi morieris ibique sepelieris, tu et omnes amici tui, quibus prophetasti mendacium ".
JER|20|7|Seduxisti me, Domine, et seductus sum;fortior me fuisti et invaluisti.Factus sum in derisum tota die,omnes subsannant me.
JER|20|8|Quia quotiescumque loquor, vociferor,iniquitatem et vastitatem clamito;et factus est mihi sermo Dominiin opprobrium et in derisum tota die.
JER|20|9|Et dixi: " Non recordabor eiusneque loquar ultra in nomine illius ".Et factus est in corde meo quasi ignis exaestuansclaususque in ossibus meis:et defeci, ferre non sustinens.
JER|20|10|Audivi enim contumelias multorumet terrorem in circuitu: Denuntiate, et denuntiemus eum ".Omnes pacifici mei observabant lapsum meum: Forte decipietur, et praevalebimus adversus eumet consequemur ultionem ex eo ".
JER|20|11|Dominus autem mecum est quasi bellator fortis;idcirco, qui persequuntur me,cadent et infirmi erunt.Confundentur vehementer, quia non prosperati sunt;opprobrium sempiternum, quod numquam delebitur.
JER|20|12|Et tu, Domine exercituum,probator iusti, qui vides renes et cor,videam, quaeso, ultionem tuam ex eis;tibi enim revelavi causam meam.
JER|20|13|Cantate Domino, laudate Dominum,quia liberavit animam pauperisde manu malorum.
JER|20|14|Maledicta dies, in qua natus sum;dies, in qua peperit me mater mea,non sit benedicta.
JER|20|15|Maledictus vir, qui annuntiavit patri meodicens: " Natus est tibi puer masculus "et gaudio laetificavit eum;
JER|20|16|sit homo ille, ut sunt civitates,quas subvertit Dominuset non paenituit eum:audiat clamorem maneet ululatum in tempore meridiano,
JER|20|17|qui non me interfecit a vulva,ut fieret mihi mater mea sepulcrum,et vulva eius conceptus aeternus.
JER|20|18|Quare de vulva egressus sum,ut viderem laborem et dolorem,et consumerentur in confusione dies mei?
JER|21|1|Verbum, quod factum est ad Ieremiam a Domino, quando misit ad eum rex Sedecias Phassur filium Melchiae et Sophoniam filium Maasiae sacerdotem dicens:
JER|21|2|" Interroga pro nobis Dominum, quia Nabuchodonosor rex Babylonis proeliatur adversum nos; si forte faciat Dominus nobiscum secundum omnia mirabilia sua, et recedat a nobis ".
JER|21|3|Et dixit Ieremias ad eos: " Sic dicetis Sedeciae:
JER|21|4|Haec dicit Dominus, Deus Israel: Ecce ego convertam vasa belli, quae in manibus vestris sunt et quibus vos pugnatis adversum regem Babylonis et Chaldaeos, qui obsident vos in circuitu murorum; et congregabo eos in medio civitatis huius.
JER|21|5|Et debellabo ego vos in manu extenta et in brachio forti et in furore et in indignatione et in ira grandi
JER|21|6|et percutiam habitatores civitatis huius, homines et bestias: pestilentia magna morientur.
JER|21|7|Et post haec, ait Dominus, dabo Sedeciam regem Iudae et servos eius et populum eius, qui derelicti sunt in civitate hac a peste et gladio et fame, in manu Nabuchodonosor regis Babylonis et in manu inimicorum eorum et in manu quaerentium animam eorum; et percutiet eos in ore gladii et non flectetur neque parcet nec miserebitur.
JER|21|8|Et ad populum hunc dices: Haec dicit Dominus: Ecce ego do coram vobis viam vitae et viam mortis:
JER|21|9|qui habitaverit in urbe hac, morietur gladio et fame et peste; qui autem egressus fuerit et transfugerit ad Chaldaeos, qui obsident vos, vivet, et erit ei anima sua quasi spolium.
JER|21|10|Posui enim faciem meam super civitatem hanc in malum et non in bonum, ait Dominus: in manu regis Babylonis dabitur, et exuret eam igni.
JER|21|11|Et domui regis Iudae:Audite verbum Domini,
JER|21|12|domus David. Haec dicit Dominus:Iudicate mane iudiciumet eruite vi oppressum de manu expoliantis,ne forte egrediatur ut ignis indignatio meaet succendatur, et non sit qui exstinguat,propter malitiam operum vestrorum.
JER|21|13|Ecce ego ad te, habitatricem vallis,petram in planitie,ait Dominus;qui dicitis: "Quis invadet nos?Et quis ingredietur domos nostras?".
JER|21|14|Et visitabo super vos iuxta fructum operum vestrorum,dicit Dominus;et succendam ignem in saltu eius,et devorabit omnia in circuitu eius ".
JER|22|1|Haec dicit Dominus: " Descende in domum regis Iudae et loqueris ibi verbum hoc
JER|22|2|et dices: Audi verbum Domini, rex Iudae, qui sedes super solium David, tu et servi tui et populus tuus, qui ingredimini per portas istas.
JER|22|3|Haec dicit Dominus: Facite iudicium et iustitiam et liberate vi oppressum de manu expoliantis et advenam et pupillum et viduam nolite affligere neque opprimatis inique et sanguinem innocentem ne effundatis in loco isto.
JER|22|4|Si enim facientes feceritis verbum istud, ingredientur per portas domus huius reges, sedentes de genere David super thronum eius et ascendentes currus et equos, ipsi et servi et populus eorum.
JER|22|5|Quod si non audieritis verba haec, in memetipso iuravi, dicit Dominus, quia in solitudinem erit domus haec.
JER|22|6|Quia haec dicit Dominus super domum regis Iudae:Galaad tu mihi,caput Libani,verumtamen ponam te solitudinem,urbes inhabitabiles,
JER|22|7|et sanctificabo super teinterficientem virum et arma eius,et succident electas cedros tuaset praecipitabunt in ignem.
JER|22|8|Et pertransibunt gentes multae per civitatem hanc, et dicet unusquisque proximo suo: "Quare fecit Dominus sic civitati huic grandi?".
JER|22|9|Et respondebunt: "Eo quod dereliquerint pactum Domini Dei sui et adoraverint deos alienos et servierint eis" ".
JER|22|10|Nolite flere mortuumneque lugeatis super eum fletu;plangite eum, qui egreditur,quia non revertetur ultranec videbit terram nativitatis suae.
JER|22|11|Quia haec dicit Dominus ad Sellum filium Iosiae regem Iudae, qui regnavit pro Iosia patre suo: " Qui egressus est de loco isto, non revertetur huc amplius,
JER|22|12|sed in loco, ad quem transtulerunt eum, ibi morietur et terram istam non videbit amplius ".
JER|22|13|Vae, qui aedificat domum suam in iniustitiaet cenacula sua non in iudicio,proximum suum servire facit gratiset mercedem eius non reddet ei;
JER|22|14|qui dicit: " Aedificabo mihi domum latamet cenacula spatiosa ";qui aperit sibi fenestraset facit laquearia cedrinapingitque sinopide!
JER|22|15|Numquid regnabis,quoniam gloriaris in cedris?Pater tuus numquid non comedit et bibit?Sed fecit iudicium et iustitiam,tunc bene erat ei.
JER|22|16|Iudicavit causam pauperis et egeni,tunc bene. Numquid non hoc est nosse me? ",dicit Dominus.
JER|22|17|Tui vero oculi et cor tuum nonnisi ad avaritiamet ad sanguinem innocentem fundendumet ad calumniam et ad oppressionem faciendam.
JER|22|18|Propterea haec dicit Dominus ad Ioachim filium Iosiae regem Iudae: Non plangent eum:Vae, frater meus!" et "Vae, soror!".Non concrepabunt ei:Vae, domine!" et "Vae, inclite!".
JER|22|19|Sepultura asini sepelietur,tractus et proiectus longeextra portas Ierusalem ".
JER|22|20|Ascende Libanum et clamaet in Basan da vocem tuamet clama de Abarim,quia contriti sunt omnes amatores tui.
JER|22|21|Locutus sum ad te in securitate tua,et dixisti: " Non audiam! ".Haec est via tua ab adulescentia tua,quia non audisti vocem meam.
JER|22|22|Omnes pastores tuos pascet ventus,et amatores tui in captivitatem ibunt,quia tunc confunderis et erubescesab omni malitia tua.
JER|22|23|Quae sedes in Libanoet nidificas in cedris,quomodo congemisces,cum venerint tibi doloresquasi dolores parturientis!
JER|22|24|" Vivo ego, dicit Dominus, quia si fuerit Iechonias, filius Ioachim rex Iudae, anulus in manu dextera mea, inde evellam eum
JER|22|25|et dabo te in manu quaerentium animam tuam et in manu, quorum tu formidas faciem, in manu Nabuchodonosor, regis Babylonis, et in manu Chaldaeorum;
JER|22|26|et mittam te et matrem tuam, quae genuit te, in terram alienam, in qua nati non estis, ibique moriemini;
JER|22|27|et in terram, ad quam ipsi levant animam suam, ut revertantur, illuc non revertentur ".
JER|22|28|Numquid vas despectum et contritum, vir iste Iechonias? Numquid vas absque omni voluptate? Quare abiecti sunt, ipse et semen eius, et proiecti in terram, quam ignoraverunt?
JER|22|29|Terra, terra, terra, audi sermonem Domini!
JER|22|30|Haec dicit Dominus: " Scribite virum istum sterilem, virum, qui in diebus suis non prosperabitur; nec enim erit de semine eius vir, qui sedeat super solium David et potestatem habeat ultra in Iuda ".
JER|23|1|"Vae pastoribus, qui disper dunt et dissipant gregem pascuae meae!, dicit Dominus.
JER|23|2|Ideo haec dicit Dominus, Deus Israel, ad pastores, qui pascunt populum meum: Vos dissipastis gregem meum et eiecistis eos et non visitastis eos; ecce ego visitabo super vos malitiam operum vestrorum, ait Dominus.
JER|23|3|Et ego congregabo reliquias gregis mei de omnibus terris, ad quas eiecero eos, et convertam eos ad rura sua, et crescent et multiplicabuntur.
JER|23|4|Et suscitabo super eos pastores, et pascent eos; non formidabunt ultra et non pavebunt, et nullus quaeretur ex numero, dicit Dominus.
JER|23|5|Ecce dies veniunt,dicit Dominus,et suscitabo David germen iustum;et regnabit rex et sapiens eritet faciet iudicium et iustitiam in terra.
JER|23|6|In diebus illis salvabitur Iuda,et Israel habitabit confidenter;et hoc est nomen, quod vocabunt eum:Dominus iustitia nostra.
JER|23|7|Propter hoc ecce dies veniunt, dicit Dominus, et non dicent ultra: Vivit Dominus, qui eduxit filios Israel de terra Aegypti!",
JER|23|8|sed: "Vivit Dominus, qui eduxit et adduxit semen domus Israel de terra aquilonis et de cunctis terris!", ad quas eieceram eos; et habitabunt in terra sua ".
JER|23|9|Ad prophetas.Contritum est cor meum in medio mei,contremuerunt omnia ossa mea;factus sum quasi vir ebriuset quasi homo madidus a vino,a facie Dominiet a facie verborum sanctorum eius;
JER|23|10|quia adulteris repleta est terra,quia a facie maledictionis luxit terra,arefacta sunt arva deserti,factus est cursus eorum malus,et fortitudo eorum iniustitia.
JER|23|11|" Propheta namque et sacerdos polluti sunt,et in domo mea inveni malum eorum,ait Dominus.
JER|23|12|Idcirco via eorum erit quasi lubricum;in tenebras proicientur et cadent in eis;afferam enim super eos mala,annum visitationis eorum,ait Dominus.
JER|23|13|Et in prophetis Samariae vidi fatuitatem:prophetabant in Baalet decipiebant populum meum Israel.
JER|23|14|Et in prophetis Ierusalem vidi horribilia:adulterium faciunt et in mendacio ambulant;et confortaverunt manus pessimorum,ut non converteretur unusquisque a malitia sua:facti sunt mihi omnes ut Sodoma,et habitatores eius quasi Gomorra ".
JER|23|15|Propterea haec dicit Dominus exercituum ad prophetas: Ecce ego cibabo eos absinthioet potabo eos felle;a prophetis enim Ierusalemegressa est pollutio super omnem terram.
JER|23|16|Haec dicit Dominus exercituum: Nolite audire verba prophetarum, qui prophetant vobis et decipiunt vos; visionem cordis sui loquuntur, non de ore Domini.
JER|23|17|Dicunt his, qui despiciunt me:Locutus est Dominus: Pax erit vobis";et omni, qui ambulat in pravitate cordis sui,dixerunt: "Non veniet super vos malum".
JER|23|18|Quis enim affuit in consilio Domini et vidit et audivit sermonem eius? Quis consideravit verbum illius et audivit?
JER|23|19|Ecce turbo Domini, indignatio egressa est,et tempestas erumpens super caput impiorum irruet.
JER|23|20|Non cessabit furor Domini, usque dum faciatet usque dum compleat cogitationes cordis sui;in novissimis diebus intellegetis consilium eius.
JER|23|21|Non mittebam prophetas,et ipsi currebant;non loquebar ad eos,et ipsi prophetabant.
JER|23|22|Si stetissent in consilio meo,nota fecissent verba mea populo meoet avertissent utique eos a via sua malaet ab operibus suis pessimis.
JER|23|23|Putasne Deus e vicino ego sum,dicit Dominus,et non Deus de longe?
JER|23|24|Si occultabitur vir in absconditis,ego non videbo eum?,dicit Dominus.Numquid non caelum et terram ego impleo?,dicit Dominus.
JER|23|25|Audivi, quae dixerunt prophetae prophetantes in nomine meo mendacium atque dicentes: "Somniavi, somniavi".
JER|23|26|Usquequo istud est in corde prophetarum vaticinantium mendacium et prophetantium seductionem cordis sui?
JER|23|27|Qui volunt facere, ut obliviscatur populus meus nominis mei, propter somnia eorum, quae narrat unusquisque ad proximum suum, sicut obliti sunt patres eorum nominis mei propter Baal.
JER|23|28|Propheta, qui habet somnium, narret somnium et, qui habet sermonem meum, loquatur sermonem meum vere.Quid paleis ad triticum?,dicit Dominus.
JER|23|29|Numquid non verba mea sunt quasi ignis,dicit Dominus,et quasi malleus conterens petram?
JER|23|30|Propterea ecce ego ad prophetas, ait Dominus, qui furantur verba mea unusquisque a proximo suo.
JER|23|31|Ecce ego ad prophetas, ait Dominus, qui assumunt linguas suas et aiunt: Dicit Dominus".
JER|23|32|Ecce ego ad prophetantes somnia mendacii, ait Dominus, qui narraverunt ea et seduxerunt populum meum in mendaciis suis et in iactantia sua, cum ego non misissem eos nec mandassem eis; qui nihil profuerunt populo huic, dicit Dominus.
JER|23|33|Si interrogaverit te populus iste vel propheta aut sacerdos dicens: Quod est onus Domini", dices ad eos: Vos estis onus; proiciam quippe vos, dicit Dominus.
JER|23|34|Et propheta et sacerdos et populus, qui dicit: "Onus Domini", visitabo super virum illum et super domum eius.
JER|23|35|Haec dicetis unusquisque ad proximum et ad fratrem suum: "Quid respondit Dominus?" et "Quid locutus est Dominus?".
JER|23|36|Sed "Onus Domini" ultra non memorabitis, quia onus erit unicuique sermo suus, et pervertitis verba Dei viventis, Domini exercituum, Dei nostri.
JER|23|37|Haec dices ad prophetam: "Quid respondit tibi Dominus?" et "Quid locutus est Dominus?".
JER|23|38|Si autem "Onus Domini" dixeritis, propter hoc haec dicit Dominus: Quia dixistis sermonem istum: "Onus Domini", et misi ad vos dicens: Nolite dicere: "Onus Domini";
JER|23|39|propterea, ecce ego tollam vos portans et proiciam vos et civitatem, quam dedi vobis et patribus vestris, a facie mea;
JER|23|40|et dabo vos in opprobrium sempiternum et in ignominiam aeternam, quae numquam oblivione delebitur ".
JER|24|1|Ostendit mihi Dominus, et ecce duo calathi pleni ficis positi ante templum Domini, postquam transtulit Nabuchodonosor rex Babylonis Iechoniam filium Ioachim regem Iudae et principes eius et fabrum et inclusorem de Ierusalem et adduxit eos in Babylonem.
JER|24|2|Calathus unus ficus bonas habebat nimis, ut solent ficus esse primi temporis; et calathus unus ficus habebat malas nimis, quae comedi non poterant, eo quod essent malae.
JER|24|3|Et dixit Dominus ad me: " Quid tu vides, Ieremia? ". Et dixi: " Ficus, ficus bonas, bonas valde, et malas, malas valde, quae comedi non possunt, eo quod sint malae ".
JER|24|4|Et factum est verbum Domini ad me dicens:
JER|24|5|" Haec dicit Dominus, Deus Israel: Sicut ficus hae bonae, sic cognoscam transmigrationem Iudae, quam emisi de loco isto in terram Chaldaeorum, in bonum.
JER|24|6|Et ponam oculos meos super eos ad placandum et reducam eos in terram hanc et aedificabo eos et non destruam et plantabo eos et non evellam.
JER|24|7|Et dabo eis cor, ut sciant me quia ego sum Dominus; et erunt mihi in populum, et ego ero eis in Deum, quia revertentur ad me in toto corde suo.
JER|24|8|Et sicut ficus pessimae, quae comedi non possunt, eo quod sint malae, haec dicit Dominus, sic dabo Sedeciam regem Iudae et principes eius et reliquos de Ierusalem, qui remanserunt in terra hac et qui habitant in terra Aegypti.
JER|24|9|Et dabo eos in vexationem afflictionemque omnibus regnis terrae, in opprobrium et in proverbium et in derisum et in maledictionem in universis locis, ad quae eieci eos.
JER|24|10|Et mittam in eis gladium et famem et pestem, donec consumantur de terra, quam dedi eis et patribus eorum ".
JER|25|1|Verbum, quod factum est ad Ieremiam de omni populo Iudae in anno quarto Ioachim filii Iosiae regis Iudae - ipse est annus primus Nabuchodonosor regis Babylonis -
JER|25|2|quod locutus est Ieremias propheta ad omnem populum Iudae et ad universos habitatores Ierusalem dicens:
JER|25|3|" A tertio decimo anno Iosiae filii Amon regis Iudae usque ad diem hanc, iste tertius et vicesimus est annus, factum est verbum Domini ad me, et locutus sum ad vos de nocte consurgens et loquens, et non audistis.
JER|25|4|Et misit Dominus ad vos omnes servos suos prophetas, consurgens diluculo mittensque; et non audistis neque inclinastis aures vestras, ut audiretis,
JER|25|5|cum diceret: "Revertimini unusquisque a via sua mala et a pessimis cogitationibus vestris, et habitabitis in terra, quam dedit Dominus vobis et patribus vestris, a saeculo et usque in saeculum;
JER|25|6|et nolite ire post deos alienos, ut serviatis eis adoretisque eos, neque me ad iracundiam provocetis in operibus manuum vestrarum, et non affligam vos.
JER|25|7|Et non audistis me, dicit Dominus, ut me ad iracundiam provocaretis in operibus manuum vestrarum, in malum vestrum".
JER|25|8|Propterea haec dicit Dominus exercituum: Pro eo quod non audistis verba mea,
JER|25|9|ecce ego mittam et assumam universas cognationes aquilonis, ait Dominus, et Nabuchodonosor regem Babylonis, servum meum, et adducam eos super terram istam et super habitatores eius et super omnes nationes, quae in circuitu illius sunt; et interficiam eos et ponam eos in stuporem et in sibilum et in ruinas sempiternas.
JER|25|10|Perdamque ex eis vocem gaudii et vocem laetitiae, vocem sponsi et vocem sponsae, vocem molae et lumen lucernae,
JER|25|11|et erit universa terra haec in solitudinem et in stuporem, et servient omnes gentes istae regi Babylonis septuaginta annis.
JER|25|12|Cumque impleti fuerint septuaginta anni, visitabo super regem Babylonis et super gentem illam, dicit Dominus, iniquitatem eorum et super terram Chaldaeorum; et ponam illam in solitudines sempiternas.
JER|25|13|Et adducam super terram illam omnia verba mea, quae locutus sum contra eam, omne, quod scriptum est in libro isto, quaecumque prophetavit Ieremias adversum omnes gentes.
JER|25|14|Quia servient eis etiam illi, gentes multae et reges magni, et reddam eis secundum opera eorum et secundum facta manuum suarum ".
JER|25|15|Quia sic dicit Dominus, Deus Israel, ad me: " Sume calicem vini furoris huius de manu mea et propinabis de illo cunctis gentibus, ad quas ego mittam te;
JER|25|16|et bibent et turbabuntur et insanient a facie gladii, quem ego mittam inter eos ".
JER|25|17|Et accepi calicem de manu Domini et propinavi cunctis gentibus, ad quas misit me Dominus,
JER|25|18|Ierusalem et civitatibus Iudae et regibus eius et principibus eius, ut darem eos in solitudinem et in stuporem, in sibilum et in maledictionem, sicut est dies ista;
JER|25|19|pharaoni regi Aegypti et servis eius et principibus eius et omni populo eius;
JER|25|20|et omni vulgo promiscuo et cunctis regibus terrae Us et cunctis regibus terrae Philisthim et Ascaloni et Gazae et Accaroni et reliquiis Azoti,
JER|25|21|Edom et Moab et filiis Ammon;
JER|25|22|et cunctis regibus Tyri et universis regibus Sidonis et regibus terrae insularum, qui sunt trans mare;
JER|25|23|et Dedan et Thema et Buz et universis, qui attonsi sunt in comam;
JER|25|24|et cunctis regibus Arabiae et cunctis regibus vulgi promiscui, qui habitant in deserto,
JER|25|25|et cunctis regibus Zimri et cunctis regibus Elam et cunctis regibus Medorum,
JER|25|26|cunctis quoque regibus aquilonis de prope et de longe, unicuique post fratrem suum et omnibus regnis terrae, quae super faciem eius sunt; et rex Sesach bibet post eos.
JER|25|27|" Et dices ad eos: Haec dicit Dominus exercituum, Deus Israel: Bibite et inebriamini et vomite; et cadite neque surgatis a facie gladii, quem ego mittam inter vos.
JER|25|28|Cumque noluerint accipere calicem de manu tua, ut bibant, dices ad eos: Haec dicit Dominus exercituum: Bibentes bibetis;
JER|25|29|quia ecce in civitate, super quam invocatum est nomen meum, ego incipio affligere, et vos immunes eritis? Non eritis immunes; gladium enim ego voco super omnes habitatores terrae, dicit Dominus exercituum.
JER|25|30|Et tu prophetabis ad eos omnia verba haec et dices ad illos:Dominus de excelso rugietet de habitaculo sancto suo dabit vocem suam;rugiens rugiet super pascua sua,celeuma quasi calcantium concineturadversus omnes habitatores terrae.
JER|25|31|Pervenit sonitus usque ad extrema terrae,quia iudicium Domino cum gentibus;in iudicium venit ipse cum omni carne;impios tradidit gladio,dicit Dominus.
JER|25|32|Haec dicit Dominus exercituum:Ecce afflictio egreditur de gente in gentem,et turbo magnus surgit a summitatibus terrae ".
JER|25|33|Et erunt interfecti Domini in die illa a summo terrae usque ad summum eius; non plangentur et non colligentur neque sepelientur: in sterquilinium super faciem terrae erunt.
JER|25|34|Ululate, pastores, et clamate;et volutamini vos in pulvere, optimates gregis,quia completi sunt dies vestri ad occisionemet ad dispersionem vestram,et cadetis quasi vasa pretiosa.
JER|25|35|Et peribit fuga a pastoribus,et salvatio ab optimatibus gregis.
JER|25|36|Vox clamoris pastorumet ululatus optimatium gregis,quia vastavit Dominus pascua eorum.
JER|25|37|Et conticuerunt arva pacisa facie irae furoris Domini.
JER|25|38|Dereliquit quasi leo umbraculum suum,quia facta est terra eorum in desolationem,a facie irae violentaeet a facie irae furoris Domini.
JER|26|1|In principio regni Ioachim filii Iosiae regis Iudae factum est verbum istud a Domino dicens:
JER|26|2|" Haec dicit Dominus: Sta in atrio domus Domini et loqueris ad omnes civitates Iudae, de quibus veniunt, ut adorent in domo Domini, universos sermones, quos ego mandavi tibi, ut loquaris ad eos: noli subtrahere verbum,
JER|26|3|si forte audiant et convertantur unusquisque a via sua mala, et paeniteat me mali, quod cogito facere eis propter malitiam operum eorum.
JER|26|4|Et dices ad eos: Haec dicit Dominus: Si non audieritis me, ut ambuletis in lege mea, quam dedi vobis,
JER|26|5|ut audiatis sermones servorum meorum prophetarum, quos ego misi ad vos de nocte consurgens et dirigens, et non audistis,
JER|26|6|dabo domum istam sicut Silo et urbem hanc dabo in maledictionem cunctis gentibus terrae ".
JER|26|7|Et audierunt sacerdotes et prophetae et omnis populus Ieremiam loquentem verba haec in domo Domini.
JER|26|8|Cumque complesset Ieremias loquens omnia, quae praeceperat ei Dominus, ut loqueretur ad universum populum, apprehenderunt eum sacerdotes et prophetae et omnis populus dicens: " Morte moriaris!
JER|26|9|Quare prophetasti in nomine Domini dicens: "Sicut Silo erit domus haec, et urbs ista desolabitur, eo quod non sit habitator"? ".Et congregatus est omnis populus adversus Ieremiam in domo Domini.
JER|26|10|Et audierunt principes Iudae verba haec et ascenderunt de domo regis in domum Domini et sederunt in introitu portae domus Domini Novae.
JER|26|11|Et locuti sunt sacerdotes et prophetae ad principes et ad omnem populum dicentes: " Iudicium mortis est viro huic, quia prophetavit adversus civitatem istam, sicut audistis auribus vestris ".
JER|26|12|Et ait Ieremias ad omnes principes et ad universum populum dicens: " Dominus misit me, ut prophetarem ad domum istam et ad civitatem hanc omnia verba, quae audistis.
JER|26|13|Nunc ergo bonas facite vias vestras et opera vestra et audite vocem Domini Dei vestri, et paenitebit Dominum mali, quod locutus est adversum vos.
JER|26|14|Ego autem ecce in manibus vestris sum; facite mihi, quod bonum et rectum est in oculis vestris.
JER|26|15|Verumtamen scitote et cognoscite quod si occideritis me, sanguinem innocentem tradetis contra vosmetipsos et contra civitatem istam et habitatores eius; in veritate enim misit me Dominus ad vos, ut loquerer in auribus vestris omnia verba haec ".
JER|26|16|Et dixerunt principes et omnis populus ad sacerdotes et prophetas: " Non est viro huic iudicium mortis, quia in nomine Domini Dei nostri locutus est ad nos ".
JER|26|17|Surrexerunt ergo viri de senioribus terrae et dixerunt ad omnem coetum populi loquentes:
JER|26|18|" Michaeas Morasthites fuit propheta in diebus Ezechiae regis Iudae et ait ad omnem populum Iudae dicens: "Haec dicit Dominus exercituum:Sion quasi ager arabitur,et Ierusalem in acervum lapidum erit,et mons domus in excelsa silvarum".
JER|26|19|Numquid morte condemnavit eum Ezechias rex Iudae et omnis Iuda? Numquid non timuerunt Dominum et deprecati sunt faciem Domini, et paenituit Dominum mali, quod locutus fuerat adversum eos? Et nos facimus malum grande contra animas nostras! ".
JER|26|20|Fuit quoque vir prophetans in nomine Domini Urias filius Semei de Cariathiarim et prophetavit adversus civitatem istam et adversus terram hanc iuxta omnia verba Ieremiae.
JER|26|21|Et audivit rex Ioachim et omnes potentes et principes eius verba haec, et quaesivit rex interficere eum; et audivit Urias et timuit fugitque et ingressus est Aegyptum.
JER|26|22|Et misit rex Ioachim viros in Aegyptum, Elnathan filium Achobor et viros cum eo in Aegyptum;
JER|26|23|et eduxerunt Uriam de Aegypto et adduxerunt eum ad regem Ioachim, et percussit eum gladio et proiecit cadaver eius in sepulcris filiorum vulgi.
JER|26|24|Igitur manus Ahicam filii Saphan fuit cum Ieremia, ut non traderetur in manus populi, et interficerent eum.
JER|27|1|In principio regni Sedeciae filii Iosiae regis Iudae factum est verbum istud ad Ieremiam a Domino dicens:
JER|27|2|" Haec dicit Dominus ad me: Fac tibi vincula et iuga et pones ea in collo tuo
JER|27|3|et mittes ea ad regem Edom et ad regem Moab et ad regem filiorum Ammon et ad regem Tyri et ad regem Sidonis in manu nuntiorum, qui venerunt Ierusalem ad Sedeciam regem Iudae;
JER|27|4|et praecipies eis, ut ad dominos suos loquantur: Haec dicit Dominus exercituum, Deus Israel: Haec dicetis ad dominos vestros:
JER|27|5|Ego feci terram et hominem et iumenta, quae sunt super faciem terrae, in fortitudine mea magna et in brachio meo extento et dedi eam ei, qui placuit in oculis meis.
JER|27|6|Et nunc itaque ego dedi omnes terras istas in manu Nabuchodonosor regis Babylonis servi mei, insuper et bestias agri dedi ei, ut serviant illi;
JER|27|7|et servient ei omnes gentes et filio eius et filio filii eius, donec veniat tempus terrae eius etiam ipsius; et servient ei gentes multae et reges magni.
JER|27|8|Gens autem et regnum, quod non servierit Nabuchodonosor regi Babylonis, et quicumque non curvaverit collum suum sub iugo regis Babylonis, in gladio et in fame et in peste visitabo super gentem illam, ait Dominus, donec consumam eos in manu eius.
JER|27|9|Vos ergo nolite audire prophetas vestros et divinos et somniatores et augures et maleficos, qui dicunt vobis: "Non servietis regi Babylonis",
JER|27|10|quia mendacium prophetant vobis, ut longe vos faciant de terra vestra, et eiciam vos, et pereatis.
JER|27|11|Porro gens, quae subiecerit cervicem suam sub iugo regis Babylonis et servierit ei, dimittam eam in terra sua, dicit Dominus, et colet eam et habitabit in ea ".
JER|27|12|Et ad Sedeciam regem Iudae locutus sum secundum omnia verba haec dicens: " Subicite colla vestra sub iugo regis Babylonis et servite ei et populo eius, et vivetis.
JER|27|13|Quare moriemini tu et populus tuus gladio, fame et peste, sicut locutus est Dominus ad gentem, quae servire noluerit regi Babylonis?
JER|27|14|Nolite audire verba prophetarum dicentium vobis: "Non servietis regi Babylonis", quia mendacium ipsi loquuntur vobis.
JER|27|15|Quia non misi eos, ait Dominus, et ipsi prophetant in nomine meo mendaciter, ut eiciam vos et pereatis, tam vos quam prophetae, qui vaticinantur vobis ".
JER|27|16|Et ad sacerdotes et ad populum istum locutus sum dicens: " Haec dicit Dominus: Nolite audire verba prophetarum vestrorum, qui prophetant vobis dicentes: "Ecce vasa domus Domini revertentur de Babylone nunc cito". Mendacium enim prophetant vobis.
JER|27|17|Nolite ergo audire eos, sed servite regi Babylonis, ut vivatis. Quare datur haec civitas in solitudinem?
JER|27|18|Et si prophetae sunt, et est verbum Domini in eis, occurrant Domino exercituum, ut non veniant vasa, quae derelicta fuerant in domo Domini et in domo regis Iudae et in Ierusalem, in Babylonem ".
JER|27|19|Quia haec dicit Dominus exercituum ad columnas et ad mare et ad bases et ad reliqua vasorum, quae remanserunt in civitate hac,
JER|27|20|quae non tulit Nabuchodonosor rex Babylonis, cum transferret Iechoniam filium Ioachim regem Iudae de Ierusalem in Babylonem et omnes optimates Iudae et Ierusalem;
JER|27|21|quia haec dicit Dominus exercituum, Deus Israel, ad vasa, quae derelicta sunt in domo Domini et in domo regis Iudae et Ierusalem:
JER|27|22|"In Babylonem transferentur et ibi erunt usque ad diem visitationis eorum, dicit Dominus; et afferri faciam ea et restitui in loco isto ".
JER|28|1|Et factum est in anno illo, in principio regni Sedeciae regis Iudae, in anno quarto in mense quinto, dixit ad me Hananias filius Azur propheta de Gabaon in domo Domini coram sacerdotibus et omni populo dicens:
JER|28|2|" Haec dicit Domi nus exercituum, Deus Israel: Contrivi iugum regis Babylonis.
JER|28|3|Adhuc duo anni dierum, et ego referri faciam ad locum istum omnia vasa domus Domini, quae tulit Nabuchodonosor rex Babylonis de loco isto et transtulit ea in Babylonem.
JER|28|4|Et Iechoniam filium Ioachim regem Iudae et omnem transmigrationem Iudae, qui ingressi sunt in Babylonem, ego convertam ad locum istum, ait Dominus; conteram enim iugum regis Babylonis ".
JER|28|5|Et dixit Ieremias propheta ad Hananiam prophetam in oculis sacerdotum et in oculis omnis populi, qui stabat in domo Domini,
JER|28|6|et ait Ieremias propheta: " Amen, sic faciat Dominus! Suscitet Dominus verba tua, quae prophetasti, ut referantur vasa in domum Domini et omnis transmigratio de Babylone ad locum istum.
JER|28|7|Verumtamen audi verbum hoc, quod ego loquor in auribus tuis et in auribus universi populi:
JER|28|8|Prophetae, qui fuerunt ante me et ante te ab initio et prophetaverunt super terras multas et super regna magna de proelio et de afflictione et de peste;
JER|28|9|propheta, qui vaticinatur pacem, cum venerit verbum eius, scietur propheta, quem misit Dominus in veritate ".
JER|28|10|Et tulit Hananias propheta iugum de collo Ieremiae prophetae et confregit illud;
JER|28|11|et ait Hananias in conspectu omnis populi dicens: " Haec dicit Dominus: Sic confringam iugum Nabuchodonosor regis Babylonis post duos annos dierum de collo omnium gentium ". Et abiit Ieremias propheta in viam suam.
JER|28|12|Et factum est verbum Domini ad Ieremiam, postquam confregit Hananias propheta iugum de collo Ieremiae prophetae, dicens:
JER|28|13|"Vade et dices Hananiae: Haec dicit Dominus: Iuga lignea contrivisti et facies pro eis iuga ferrea.
JER|28|14|Quia haec dicit Dominus exercituum, Deus Israel: Iugum ferreum posui super collum cunctarum gentium istarum, ut serviant Nabuchodonosor regi Babylonis, et servient ei; insuper et bestias terrae dedi ei ".
JER|28|15|Et dixit Ieremias propheta ad Hananiam prophetam: "Audi, Hanania! Non misit te Dominus, et tu confidere fecisti populum istum in mendacio.
JER|28|16|Idcirco haec dicit Dominus: Ecce emittam te a facie terrae; hoc anno morieris, adversum enim Dominum praevaricationem locutus es ".
JER|28|17|Et mortuus est Hananias propheta in anno illo, mense septimo.
JER|29|1|Et haec sunt verba epistulae, quam misit Ieremias propheta de Ierusalem ad reliquias seniorum transmigrationis et ad sacerdotes et ad prophetas et ad omnem populum, quem traduxerat Nabuchodonosor de Ierusalem in Babylonem,
JER|29|2|postquam egressus est Iechonias rex et domina et eunuchi et principes Iudae et Ierusalem et faber et inclusor de Ierusalem,
JER|29|3|in manu Elasa filii Saphan et Gamariae filii Helciae, quos misit Sedecias rex Iudae ad Nabuchodonosor regem Babylonis in Babylonem dicens:
JER|29|4|" Haec dicit Dominus exercituum, Deus Israel, omni transmigrationi, quam transtuli de Ierusalem in Babylonem:
JER|29|5|Aedificate domos et habitate et plantate hortos et comedite fructum eorum,
JER|29|6|accipite uxores et generate filios et filias et date filiis vestris uxores et filias vestras date viris, et pariant filios et filias, et multiplicamini ibi et nolite esse pauci numero.
JER|29|7|Et quaerite pacem civitatis, ad quam transmigrare vos feci, et orate pro ea ad Dominum, quia in pace illius erit pax vobis.
JER|29|8|Haec enim dicit Dominus exercituum, Deus Israel: Non vos seducant prophetae vestri, qui sunt in medio vestrum, et divini vestri, et ne attendatis ad somnia vestra, quae vos somniatis,
JER|29|9|quia falso ipsi prophetant vobis in nomine meo, et non misi eos, dicit Dominus.
JER|29|10|Quia haec dicit Dominus: Cum impleti fuerint in Babylone septuaginta anni, visitabo vos et suscitabo super vos verbum meum bonum, ut reducam vos ad locum istum.
JER|29|11|Ego enim scio cogitationes, quas ego cogito super vos, ait Dominus, cogitationes pacis et non afflictionis, ut dem vobis posteritatem et spem.
JER|29|12|Et invocabitis me et ibitis; et orabitis me, et ego exaudiam vos.
JER|29|13|Quaeretis me et invenietis, cum quaesieritis me in toto corde vestro.
JER|29|14|Et inveniar a vobis, ait Dominus, et reducam captivitatem vestram et congregabo vos de universis gentibus et de cunctis locis, ad quae expuli vos, dicit Dominus; et reverti vos faciam ad locum, de quo transmigrare vos feci.
JER|29|15|Quia dixistis: "Suscitavit nobis Dominus prophetas in Babylone".
JER|29|16|Quia haec dicit Dominus ad regem, qui sedet super solium David, et ad omnem populum habitatorem urbis huius, ad fratres vestros, qui non sunt egressi vobiscum in transmigrationem,
JER|29|17|haec dicit Dominus exercituum: Ecce mittam in eis gladium et famem et pestem et ponam eos quasi ficus malas, quae comedi non possunt, eo quod pessimae sint;
JER|29|18|et persequar eos in gladio et in fame et in pestilentia et dabo eos in vexationem universis regnis terrae, in maledictionem et in stuporem et in sibilum et in opprobrium cunctis gentibus, ad quas ego eieci eos,
JER|29|19|eo quod non audierint verba mea, dicit Dominus, quae misi ad eos per servos meos prophetas, de nocte consurgens et mittens, et non audistis, dicit Dominus.
JER|29|20|Vos ergo audite verbum Domini, omnis transmigratio, quam emisi de Ierusalem in Babylonem.
JER|29|21|Haec dicit Dominus exercituum, Deus Israel, ad Achab filium Colaiae et ad Sedeciam filium Maasiae, qui prophetant vobis in nomine meo mendaciter: Ecce ego tradam eos in manu Nabuchodonosor regis Babylonis, et percutiet eos in oculis vestris;
JER|29|22|et assumetur ex eis maledictio omni transmigrationi Iudae, quae est in Babylone, dicentium: "Ponat te Dominus sicut Sedeciam et sicut Achab, quos frixit rex Babylonis in igne!";
JER|29|23|pro eo quod fecerint stultitiam in Israel et moechati sunt in uxores amicorum suorum et locuti sunt verbum in nomine meo mendaciter, quod non mandavi eis. Ego enim scio et sum testis, dicit Dominus.
JER|29|24|Et ad Semeiam Nehelamiten dices:
JER|29|25|Haec dicit Dominus exercituum, Deus Israel, pro eo quod misisti in nomine tuo epistulas ad omnem populum, qui est in Ierusalem, et ad Sophoniam filium Maasiae sacerdotem et ad universos sacerdotes dicens:
JER|29|26|"Dominus dedit te sacerdotem pro Ioiada sacerdote, ut sis praefectus in domo Domini super omnem virum arrepticium et prophetantem, ut mittas eum in nervum et in vincula.
JER|29|27|Et nunc quare non increpasti Ieremiam Anathothiten, qui prophetat vobis?
JER|29|28|Quia super hoc misit ad nos in Babylonem dicens: Longum est; aedificate domos et habitate et plantate hortos et comedite fructum eorum" ".
JER|29|29|Legit ergo Sophonias sacerdos epistulam istam in auribus Ieremiae prophetae.
JER|29|30|Et factum est verbum Domini ad Ieremiam dicens:
JER|29|31|" Mitte ad omnem transmigrationem dicens: Haec dicit Dominus ad Semeiam Nehelamiten: Pro eo quod prophetavit vobis Semeias, et ego non misi eum, et fecit vos confidere in mendacio,
JER|29|32|idcirco haec dicit Dominus: Ecce ego visitabo super Semeiam Nehelamiten et super semen eius; non erit ei vir sedens in medio populi huius, et non videbit bonum, quod ego faciam populo meo, ait Dominus, quia praevaricationem locutus est adversus Dominum ".
JER|30|1|Verbum, quod factum est ad Ieremiam a Domino dicens:
JER|30|2|" Haec dicit Dominus, Deus Israel, dicens: Scribe tibi omnia verba, quae locutus sum ad te, in libro;
JER|30|3|ecce enim dies veniunt, dicit Dominus, et convertam sortem populi mei Israel et Iudae, ait Dominus, et convertam eos ad terram, quam dedi patribus eorum, et possidebunt eam ".
JER|30|4|Et haec verba, quae locutus est Dominus ad Israel et ad Iudam:
JER|30|5|" Quoniam haec dicit Dominus:Vocem terroris audivimus,formido et non est pax.
JER|30|6|Interrogate et videte, si generat masculus;quare ergo vidi omnis viri manumsuper lumbum suum quasi parturientis,et conversae sunt universae facies in auruginem?
JER|30|7|Vae, quia magna dies illa,nec est similis eius,tempusque tribulationis est Iacob,et ex ipso salvabitur.
JER|30|8|Et erit: in die illa, ait Dominus exercituum, conteram iugum eius de collo tuo et vincula tua dirumpam; et non dominabuntur ei amplius alieni,
JER|30|9|sed servient Domino Deo suo et David regi suo, quem suscitabo eis.
JER|30|10|Tu ergo ne timeas, serve meus Iacob,ait Dominus,neque paveas, Israel,quia ecce ego salvabo te de terra longinquaet semen tuum de terra captivitatis eorum;et revertetur Iacob et quiescetet securus erit, et non erit quem formidet;
JER|30|11|quoniam tecum ego sum,ait Dominus,ut salvem te.Faciam enim consummationem in cunctis gentibus,in quibus dispersi te;te autem non faciam in consummationem,sed castigabo te in iudicionec quasi innocenti parcam tibi.
JER|30|12|Quia haec dicit Dominus:Insanabilis fractura tua,pessima plaga tua;
JER|30|13|non est qui iudicet iudicium tuum;sunt ulceri medicamina,tibi vero cicatrix non obducitur.
JER|30|14|Omnes amatores tui obliti sunt tui,te non quaerunt;plaga enim inimici percussi tecastigatione crudeli:propter multitudinem iniquitatis tuaedura facta sunt peccata tua.
JER|30|15|Quid clamas super contritione tua?Insanabilis est dolor tuus.Propter multitudinem iniquitatis tuaeet propter dura peccata tua feci haec tibi.
JER|30|16|Propterea omnes, qui comedunt te, devorabuntur,et universi hostes tui in captivitatem ducentur,et, qui te vastant, vastabuntur,cunctosque praedatores tuos dabo in praedam.
JER|30|17|Obducam enim cicatricem tibiet a vulneribus tuis sanabo te,dicit Dominus,quia Eiectam vocaverunt te,Sion haec, quae non habebat requirentem.
JER|30|18|Haec dicit Dominus:Ecce ego convertam sortem tabernaculorum Iacobet tectis eius miserebor,et aedificabitur civitas in ruinis suis,et arx in loco suo fundabitur;
JER|30|19|et egredietur de eis laus voxque ludentium.Et multiplicabo eos, et non imminuentur,et glorificabo eos, et non attenuabuntur.
JER|30|20|Et erunt filii eius sicut a principio,et coetus eius coram me permanebit,et visitabo adversum omnes, qui tribulant eum.
JER|30|21|Et erit dux eius ex eo,et princeps de medio eius procedet; et applicabo eum, et accedet ad me.Quis enim iste est, qui pignori dabit cor suum,ut appropinquet mihi?,ait Dominus.
JER|30|22|Et eritis mihi in populum,et ego ero vobis in Deum.
JER|30|23|Ecce turbo Domini, furor egrediens,procella ruens;in capite impiorum conquiescet.
JER|30|24|Non cessabit ab ira indignationis Dominus,donec faciat et compleatcogitationes cordis sui;in novissimo dierum intellegetis ea.
JER|31|1|In tempore illo,dicit Dominus,ero Deus universis cognationibus Israel,et ipsi erunt mihi in populum.
JER|31|2|Haec dicit Dominus:Invenit gratiam in desertopopulus, qui remanserat a gladio;vadet ad requiem suam Israel ".
JER|31|3|De longe Dominus apparuit mihi: In caritate perpetua dilexi te;ideo attraxi te in misericordia.
JER|31|4|Rursumque aedificabo te, et aedificaberis,virgo Israel;adhuc ornaberis tympanis tuiset egredieris in choro ludentium.
JER|31|5|Adhuc plantabis vineas in montibus Samariae;plantabunt plantanteset vindemiabunt.
JER|31|6|Quia erit dies, in qua clamabunt custodesin monte Ephraim:Surgite, et ascendamus in Sionad Dominum Deum nostrum".
JER|31|7|Quia haec dicit Dominus:Exsultate in laetitia propter Iacobet hinnite capiti gentium;personate, canite et dicite:Salva, Domine, populum tuum,reliquias Israel".
JER|31|8|Ecce ego adducam eos de terra aquiloniset congregabo eos ab extremis terrae;inter quos erunt caecus et claudus, praegnans et pariens simul:coetus magnus revertentium huc.
JER|31|9|In fletu venient,et in deprecatione reducam eoset adducam eos per torrentes aquarumin via recta, et non impingent in ea, quia factus sum Israeli pater,et Ephraim primogenitus meus est ".
JER|31|10|Audite verbum Domini, gentes,et annuntiate in insulis, quae procul sunt, et dicite: Qui dispersit Israel, congregabit eumet custodiet eum sicut pastor gregem suum ".
JER|31|11|Redemit enim Dominus Iacobet liberavit eum de manu potentioris.
JER|31|12|Et venient et laudabunt in monte Sionet confluent ad bona Dominisuper frumento et vino et oleoet fetu pecorum et armentorum;eritque anima eorum quasi hortus irriguus,et ultra non esurient.
JER|31|13|Tunc laetabitur virgo in choro,iuvenes et senes simul. Et convertam luctum eorum in gaudiumet consolabor eos et laetificabo a dolore suo.
JER|31|14|Et inebriabo animam sacerdotum pinguedine,et populus meus bonis meis adimplebitur ",ait Dominus.
JER|31|15|Haec dicit Dominus: Vox in Rama audita estlamentationis, luctus et fletusRachel plorantis filios suoset nolentis consolari super eis, quia non sunt ".
JER|31|16|Haec dicit Dominus: Quiescat vox tua a ploratu,et oculi tui a lacrimis,quia est merces operi tuo,ait Dominus,et revertentur de terra inimici.
JER|31|17|Et est spes novissimis tuis,ait Dominus,et revertentur filii ad terminos suos.
JER|31|18|Audiens audivi Ephraim transmigrantem:Castigasti me, et eruditus sumquasi iuvenculus indomitus;converte me, et convertar,quia tu Dominus Deus meus.
JER|31|19|Postquam enim convertisti me,egi paenitentiam;et postquam ostendisti mihi,percussi femur meum;confusus sum et erubui,quoniam sustinui opprobrium adulescentiae meae".
JER|31|20|Estne filius honorabilis mihi Ephraimaut puer delectabilis,quia ex quo locutus sum de eo,adhuc recordabor eius?Idcirco conturbata sunt viscera mea super eum:miserans miserebor eius ",ait Dominus.
JER|31|21|Statue tibi lapides,pone tibi signa,dirige cor tuum in iter,viam, in qua ambulasti;revertere, virgo Israel,revertere ad civitates tuas istas.
JER|31|22|Usquequo vagaberis,filia rebellis?Quia creavit Dominus novum super terram:femina circumdabit virum.
JER|31|23|Haec dicit Dominus exercituum, Deus Israel: " Adhuc dicent verbum istud in terra Iudae et in urbibus eius, cum convertero sortem eorum: "Benedicat tibi Dominus, habitaculum iustitiae, mons sanctus".
JER|31|24|Et habitabunt in eo Iudas et omnes civitates eius simul, agricolae et minantes greges.
JER|31|25|Quia inebriavi animam lassam et omnem animam esurientem saturavi ".
JER|31|26|Ideo quasi de somno suscitatus sum et vidi, et somnus meus dulcis mihi.
JER|31|27|" Ecce dies veniunt, dicit Dominus, et seminabo domum Israel et domum Iudae semine hominum et semine iumentorum.
JER|31|28|Et sicut vigilavi super eos, ut evellerem et demolirer et dissiparem et disperderem et affligerem, sic vigilabo super eos, ut aedificem et plantem, ait Dominus.
JER|31|29|In diebus illis non dicent ultra:Patres comederunt uvam acerbam, et dentes filiorum obstupuerunt",
JER|31|30|sed unusquisque in iniquitate sua morietur; omnis homo, qui comederit uvam acerbam, obstupescent dentes eius.
JER|31|31|Ecce dies veniunt, dicit Dominus, et feriam domui Israel et domui Iudae pactum novum;
JER|31|32|non secundum pactum, quod pepigi cum patribus eorum in die qua apprehendi manum eorum, ut educerem eos de terra Aegypti, pactum, quod irritum fecerunt, et ego dominatus sum eorum, dicit Dominus.
JER|31|33|Sed hoc erit pactum, quod feriam cum domo Israel post dies illos, dicit Dominus: Dabo legem meam in visceribus eorum et in corde eorum scribam eam; et ero eis in Deum, et ipsi erunt mihi in populum.
JER|31|34|Et non docebit ultra vir proximum suum, et vir fratrem suum dicens: Cognosce Dominum"; omnes enim cognoscent me, a minimo eorum usque ad maximum, ait Dominus, quia propitiabor iniquitati eorum et peccati eorum non memorabor amplius ".
JER|31|35|Haec dicit Dominus,qui dat solem in lumine diei,ordinem lunae et stellarum in lumine noctis,qui turbat mare, et fremunt fluctus eius,Dominus exercituum nomen illi:
JER|31|36|" Si defecerint leges istae coram me,dicit Dominus,tunc et semen Israel deficiet,ut non sit gens coram me cunctis diebus ".
JER|31|37|Haec dicit Dominus: Si mensurari potuerint caeli sursum,et investigari fundamenta terrae deorsum,et ego abiciam universum semen Israelpropter omnia, quae fecerunt,dicit Dominus.
JER|31|38|Ecce dies veniunt, dicit Dominus, et aedificabitur civitas Domino a turre Hananeel usque ad portam Anguli,
JER|31|39|et exibit ultra norma mensurae in conspectu eius super collem Gareb et vertetur in Goa,
JER|31|40|et omnis vallis cadaverum et cineris et universa regio usque ad torrentem Cedron et usque ad angulum portae Equorum orientalis sanctum Domini; non evelletur et non destruetur ultra in perpetuum ".
JER|32|1|Verbum, quod factum est ad Ieremiam a Domino in anno decimo Sedeciae regis Iudae; ipse est annus decimus octavus Nabuchodonosor.
JER|32|2|Tunc exercitus regis Babylonis obsidebat Ierusalem, et Ieremias propheta erat clausus in atrio custodiae, qui erat in domo regis Iudae.
JER|32|3|Clauserat enim eum Sedecias rex Iudae dicens: " Quare vaticinaris dicens: "Haec dicit Dominus: Ecce ego dabo civitatem istam in manu regis Babylonis, et capiet eam;
JER|32|4|et Sedecias rex Iudae non effugiet de manu Chaldaeorum, sed tradetur in manus regis Babylonis, et loquetur os eius cum ore illius, et oculi eius oculos illius videbunt;
JER|32|5|et in Babylonem ducet Sedeciam, et ibi erit, donec visitem eum, ait Dominus; si autem dimicaveritis adversum Chaldaeos, nihil prosperum habebitis"? ".
JER|32|6|Et dixit Ieremias: " Factum est verbum Domini ad me dicens:
JER|32|7|Ecce Hanameel filius Sellum patruelis tuus veniet ad te dicens: "Eme tibi agrum meum, qui est in Anathoth; tibi enim competit ex propinquitate, ut emas".
JER|32|8|Et venit ad me Hanameel filius patrui mei secundum verbum Domini ad vestibulum custodiae et ait ad me: "Posside agrum meum, qui est in Anathoth in terra Beniamin, quia tibi competit hereditas, et tu propinquus es, ut possideas". Intellexi autem quod verbum Domini esset
JER|32|9|et emi agrum ab Hanameel filio patrui mei, qui est in Anathoth, et appendi ei argentum: septem et decem siclos argenteos.
JER|32|10|Et scripsi in libro et signavi et adhibui testes et appendi argentum in statera.
JER|32|11|Et accepi librum possessionis signatum, continentem stipulationes et rata, et apertum;
JER|32|12|et dedi librum possessionis Baruch filio Neriae filii Maasiae in oculis Hanameel patruelis mei et in oculis testium, qui obsignaverant in libro emptionis, et in oculis omnium Iudaeorum, qui sedebant in atrio custodiae.
JER|32|13|Et praecepi Baruch coram eis dicens:
JER|32|14|Haec dicit Dominus exercituum, Deus Israel: Sume libros istos, librum emptionis hunc signatum et librum hunc, qui apertus est; et pones illos in vase fictili, ut permanere possint diebus multis.
JER|32|15|Haec enim dicit Dominus exercituum, Deus Israel: Adhuc possidebuntur domus et agri et vineae in terra ista.
JER|32|16|Et oravi ad Dominum, postquam tradidi librum possessionis Baruch filio Neriae, dicens:
JER|32|17|Heu, Domine Deus, ecce tu fecisti caelum et terram in fortitudine tua magna et in brachio tuo extento; non erit tibi difficile omne verbum,
JER|32|18|qui facis misericordiam in milibus et reddis iniquitatem patrum in sinum filiorum eorum post eos; Deus magne, potens, Dominus exercituum nomen eius:
JER|32|19|magnus consilio et potens in operibus, cuius oculi aperti sunt super omnes vias filiorum Adam, ut reddas unicuique secundum vias suas et secundum fructum operum eius.
JER|32|20|Qui posuisti signa et portenta in terra Aegypti usque ad diem hanc et in Israel et in hominibus; et fecisti tibi nomen, sicut est dies haec.
JER|32|21|Et eduxisti populum tuum Israel de terra Aegypti in signis et in portentis et in manu robusta et in brachio extento et in terrore magno.
JER|32|22|Et dedisti eis terram hanc, quam iurasti patribus eorum, ut dares eis, terram fluentem lacte et melle.
JER|32|23|Et ingressi sunt et possederunt eam; et non oboedierunt voci tuae et in lege tua non ambulaverunt: omnia, quae mandasti eis, ut facerent, non fecerunt; et occurrere fecisti eis omnia mala haec.
JER|32|24|Ecce munitiones exstructae sunt adversum civitatem, ut capiatur, et urbs data est in manu Chaldaeorum, qui proeliantur adversus eam, in gladio et fame et pestilentia; et quaecumque locutus es, acciderunt, ut tu ipse cernis.
JER|32|25|Et tu dicis mihi, Domine Deus: Eme agrum argento et adhibe testes, cum urbs data sit in manu Chaldaeorum ".
JER|32|26|Et factum est verbum Domini ad Ieremiam dicens:
JER|32|27|" Ecce ego Dominus, Deus universae carnis; numquid mihi difficile erit omne verbum?
JER|32|28|Propterea haec dicit Dominus: Ecce ego tradam civitatem istam in manus Chaldaeorum et in manus regis Babylonis, et capiet eam.
JER|32|29|Et venient Chaldaei proeliantes adversum urbem hanc et succendent eam igni et comburent eam et domos, in quarum domatibus sacrificabant Baal et libabant diis alienis libamina ad irritandum me.
JER|32|30|Erant enim filii Israel et filii Iudae iugiter facientes malum in oculis meis ab adulescentia sua, filii Israel, qui usque nunc exacerbant me in opere manuum suarum, dicit Dominus.
JER|32|31|Quia in furorem et in indignationem meam facta est mihi civitas haec a die, qua aedificaverunt eam, usque ad diem istam, qua auferetur de conspectu meo
JER|32|32|propter omnem malitiam filiorum Israel et filiorum Iudae, quam fecerunt, ad iracundiam me provocantes, ipsi et reges eorum, principes eorum et sacerdotes eorum et prophetae eorum, viri Iudae et habitatores Ierusalem.
JER|32|33|Et verterunt ad me terga et non facies, cum docerem eos diluculo consurgens et erudiens, et nollent audire, ut acciperent disciplinam.
JER|32|34|Et posuerunt idola sua in domo, super quam invocatum est nomen meum, ut polluerent eam;
JER|32|35|et aedificaverunt excelsa Baal, quae sunt in valle Benennom, ut initiarent filios suos et filias suas Moloch; quod non mandavi eis, nec ascendit in cor meum, ut facerent abominationem hanc et in peccatum deducerent Iudam ".
JER|32|36|Et nunc propter ista, haec dicit Dominus, Deus Israel, ad civitatem hanc, de qua vos dicitis quod tradatur in manus regis Babylonis in gladio et in fame et in peste:
JER|32|37|" Ecce ego congregabo eos de universis terris, ad quas eieci eos in furore meo et in ira mea et in indignatione grandi; et reducam eos ad locum istum et habitare eos faciam confidenter.
JER|32|38|Et erunt mihi in populum, et ego ero eis in Deum.
JER|32|39|Et dabo eis cor unum et viam unam, ut timeant me universis diebus, et bene sit eis et filiis eorum post eos.
JER|32|40|Et feriam eis pactum sempiternum et non desinam eis benefacere et timorem meum dabo in corde eorum, ut non recedant a me.
JER|32|41|Et laetabor super eis, cum bene eis fecero, et plantabo eos in terra ista in veritate, in toto corde meo et in tota anima mea.
JER|32|42|Quia haec dicit Dominus: Sicut adduxi super populum istum omne malum hoc grande, sic adducam super eos omne bonum, quod ego loquor ad eos,
JER|32|43|et possidebuntur agri in terra ista, de qua vos dicitis quod deserta sit, eo quod non remanserit homo et iumentum, et data sit in manu Chaldaeorum.
JER|32|44|Agri ementur pecunia et scribentur in libro, et imprimetur signum, et testes adhibebuntur in terra Beniamin et in circuitu Ierusalem, in civitatibus Iudae et in civitatibus montanis et in civitatibus Sephelae et in civitatibus, quae ad austrum sunt, quia convertam sortem eorum ", ait Dominus.
JER|33|1|Et factum est verbum Domi ni ad Ieremiam secundo, cum adhuc clausus esset in atrio custodiae, dicens:
JER|33|2|" Haec dicit Dominus, qui facturus est id, Dominus, qui formaturus est illud et paraturus, Dominus nomen eius:
JER|33|3|Clama ad me, et exaudiam te et annuntiabo tibi grandia et inaccessibilia, quae nescis.
JER|33|4|Quia haec dicit Dominus, Deus Israel, super domos urbis huius et ad domos regis Iudae, quae destructae sunt, pro munitionibus et pro gladio
JER|33|5|venientium, ut dimicent cum Chaldaeis et impleant eas cadaveribus hominum, quos percussi in furore meo et in indignatione mea, abscondens faciem meam a civitate hac propter omnem malitiam eorum.
JER|33|6|Ecce ego obducam ei cicatricem et sanitatem et curabo eos et revelabo illis abundantiam pacis et veritatis
JER|33|7|et convertam sortem Iudae et sortem Israel et aedificabo eos sicut a principio.
JER|33|8|Et emundabo illos ab omni iniquitate sua, in qua peccaverunt mihi, et propitius ero cunctis iniquitatibus eorum, in quibus deliquerunt mihi et spreverunt me;
JER|33|9|et erit mihi in nomen et in gaudium et in laudem et in exsultationem cunctis gentibus terrae, quae audierint omnia bona, quae ego facturus sum eis; et pavebunt et turbabuntur in universis bonis et in omni pace, quam ego faciam eis.
JER|33|10|Haec dicit Dominus: Adhuc audietur in loco isto, quem vos dicitis esse desertum, eo quod non sit homo et iumentum in civitatibus Iudae et foris Ierusalem, quae desolatae sunt absque homine et absque habitatore et absque pecore,
JER|33|11|vox gaudii et vox laetitiae, vox sponsi et vox sponsae, vox dicentium:Confitemini Domino exercituum, quoniam bonus Dominus,quoniam in aeternum misericordia eius";et portantium vota in domum Domini; reducam enim sortem terrae sicut a principio, dicit Dominus.
JER|33|12|Haec dicit Dominus exercituum: Adhuc erit in loco isto deserto, absque homine et absque iumento, et in cunctis civitatibus eius habitaculum pastorum accubantium gregum.
JER|33|13|In civitatibus montuosis et in civitatibus Sephelae et in civitatibus, quae ad austrum sunt, et in terra Beniamin et in circuitu Ierusalem et in civitatibus Iudae adhuc transibunt greges ad manum numerantis, ait Dominus.
JER|33|14|Ecce dies veniunt, dicit Dominus, et suscitabo verbum bonum, quod locutus sum ad domum Israel et ad domum Iudae.
JER|33|15|In diebus illis et in tempore illo germinare faciam David germen iustitiae, et faciet iudicium et iustitiam in terra.
JER|33|16|In diebus illis salvabitur Iuda, et Ierusalem habitabit confidenter; et hoc est nomen, quod vocabit eam: Dominus iustitia nostra.
JER|33|17|Quia haec dicit Dominus: Non interibit de David vir, qui sedeat super thronum domus Israel;
JER|33|18|et de sacerdotibus Levitis non interibit vir a facie mea, qui offerat holocautomata et incendat sacrificium et caedat victimas omnibus diebus ".
JER|33|19|Et factum est verbum Domini ad Ieremiam dicens:
JER|33|20|" Haec dicit Dominus: Si irritum potest fieri pactum meum cum die et pactum meum cum nocte, ut non sit dies et nox in tempore suo,
JER|33|21|et pactum meum irritum esse poterit cum David servo meo, ut non sit ex eo filius, qui regnet in throno eius, et cum Levitis sacerdotibus ministris meis.
JER|33|22|Sicuti enumerari non possunt stellae caeli et metiri arena maris, sic multiplicabo semen David servi mei et Levitas ministros meos ".
JER|33|23|Et factum est verbum Domini ad Ieremiam dicens:
JER|33|24|" Numquid non vidisti quid populus hic locutus sit dicens: "Duae cognationes, quas elegerat Dominus, abiectae sunt", et populum meum despexerunt, eo quod non sit ultra gens coram eis?
JER|33|25|Haec dicit Dominus: Si pactum meum inter diem et noctem et leges caelo et terrae non posui,
JER|33|26|equidem et semen Iacob et David servi mei proiciam, ut non assumam de semine eius principes seminis Abraham et Isaac et Iacob; reducam enim sortem eorum et miserebor eis ".
JER|34|1|Verbum, quod factum est ad Ieremiam a Domino, quando Nabuchodonosor rex Babylonis et omnis exercitus eius universaque regna terrae, quae erant sub potestate manus eius, et omnes populi bellabant contra Ierusalem et contra omnes urbes eius, dicens:
JER|34|2|" Haec dicit Dominus, Deus Israel: Vade et loquere ad Sedeciam regem Iudae et dices ad eum: Haec dicit Dominus: Ecce ego tradam civitatem hanc in manus regis Babylonis, et succendet eam igni;
JER|34|3|et tu non effugies de manu eius, sed comprehensione capieris et in manu eius traderis, et oculi tui oculos regis Babylonis videbunt, et os eius cum ore tuo loquetur, et Babylonem introibis.
JER|34|4|Attamen audi verbum Domini, Sedecia rex Iudae. Haec dicit Dominus ad te: Non morieris in gladio,
JER|34|5|sed in pace morieris et secundum combustiones patrum tuorum regum priorum, qui fuerunt ante te, sic comburent tibi et "Vae, domine!" plangent te, quia verbum ego locutus sum ", dicit Dominus.
JER|34|6|Et locutus est Ieremias propheta ad Sedeciam regem Iudae universa verba haec in Ierusalem;
JER|34|7|et exercitus regis Babylonis pugnabat contra Ierusalem et contra omnes civitates Iudae, quae reliquae erant, contra Lachis et contra Azeca: hae enim supererant de civitatibus Iudae urbes munitae.
JER|34|8|Verbum, quod factum est ad Ieremiam a Domino, postquam percussit rex Sedecias foedus cum omni populo in Ierusalem praedicans eis libertatem,
JER|34|9|ut dimitteret unusquisque servum suum et unusquisque ancillam suam, Hebraeum et Hebraeam, liberos et nequaquam dominarentur eis, id est in Iudaeo et fratre suo.
JER|34|10|Audierunt ergo omnes principes et universus populus, qui inierant pactum, ut dimitteret unusquisque servum suum et unusquisque ancillam suam liberos et ultra non dominarentur eis; audierunt igitur et dimiserunt.
JER|34|11|Et conversi sunt deinceps et retraxerunt servos et ancillas suas, quos dimiserant liberos, et subiugaverunt in famulos et in famulas.
JER|34|12|Et factum est verbum Domini ad Ieremiam a Domino dicens:
JER|34|13|" Haec dicit Dominus, Deus Israel: Ego percussi foedus cum patribus vestris in die, qua eduxi eos de terra Aegypti de domo servitutis, dicens:
JER|34|14|Cum completi fuerint septem anni, dimittat unusquisque fratrem suum Hebraeum, qui venditus est ei, et serviet tibi sex annis, et dimittes eum a te liberum, et non audierunt patres vestri me nec inclinaverunt aurem suam.
JER|34|15|Et conversi estis vos hodie et fecistis, quod rectum est in oculis meis, ut praedicaretis libertatem unusquisque ad proximum suum; et inistis pactum in conspectu meo in domo, super quam invocatum est nomen meum.
JER|34|16|Et reversi estis et commaculastis nomen meum et reduxistis unusquisque servum suum et unusquisque ancillam suam, quos dimiseratis, ut essent liberi et suae potestatis, et subiugastis eos, ut sint vobis servi et ancillae.
JER|34|17|Propterea haec dicit Dominus: Vos non audistis me, ut praedicaretis libertatem unusquisque fratri suo et unusquisque amico suo; ecce ego praedico vobis libertatem, ait Dominus, ad gladium et pestem et famem et dabo vos in commotionem cunctis regnis terrae.
JER|34|18|Et dabo viros, qui praevaricantur foedus meum et non observaverunt verba foederis, quibus assensi sunt in conspectu meo, sicut vitulum, quem conciderunt in duas partes et transierunt inter divisiones eius,
JER|34|19|principes Iudae et principes Ierusalem, eunuchi et sacerdotes et omnis populus terrae, qui transierunt inter divisiones vituli;
JER|34|20|et dabo eos in manu inimicorum suorum et in manu quaerentium animam eorum, et erit morticinum eorum in escam volatilibus caeli et bestiis terrae.
JER|34|21|Et Sedeciam regem Iudae et principes eius dabo in manus inimicorum suorum et in manus quaerentium animas eorum et in manus exercituum regis Babylonis, qui recesserunt a vobis.
JER|34|22|Ecce ego praecipio, dicit Dominus, et reducam eos in civitatem hanc; et proeliabuntur adversus eam et capient eam et incendent igni; et civitates Iudae dabo in solitudinem, eo quod non sit habitator ".
JER|35|1|Verbum, quod factum est ad Ieremiam a Domino in die bus Ioachim filii Iosiae regis Iudae dicens:
JER|35|2|" Vade ad domum Rechabitarum et loquere eis; et introduces eos in domum Domini in unam exedram et dabis eis bibere vinum ".
JER|35|3|Et assumpsi Iezoniam filium Ieremiae filii Habsaniae et fratres eius et omnes filios eius et universam domum Rechabitarum;
JER|35|4|et introduxi eos in domum Domini ad exedram filiorum Hanan filii Iegdaliae hominis Dei, quod erat iuxta exedram principum super exedram Maasiae filii Sellum, qui erat custos vestibuli.
JER|35|5|Et posui coram filiis domus Rechabitarum scyphos plenos vino et calices et dixi ad eos: " Bibite vinum ".
JER|35|6|Qui responderunt: " Non bibemus vinum, quia Ionadab filius Rechab pater noster praecepit nobis dicens: "Non bibetis vinum, vos et filii vestri, usque in sempiternum
JER|35|7|et domum non aedificabitis et sementem non seretis et vineas non plantabitis, nec habebitis, sed in tabernaculis habitabitis cunctis diebus vestris, ut vivatis diebus multis super faciem terrae, in qua vos peregrinamini".
JER|35|8|Oboedivimus ergo voci Ionadab filii Rechab patris nostri in omnibus, quae praecepit nobis, ita ut non biberemus vinum cunctis diebus nostris, nos et mulieres nostrae, filii et filiae nostrae,
JER|35|9|et non aedificaremus domos ad habitandum et vineam et agrum et sementem non habuimus,
JER|35|10|sed habitavimus in tabernaculis; et oboedientes fecimus iuxta omnia, quae praecepit nobis Ionadab pater noster.
JER|35|11|Cum autem ascendisset Nabuchodonosor rex Babylonis ad terram, diximus: Venite, et ingrediamur Ierusalem a facie exercitus Chaldaeorum et a facie exercitus Syriae. Et mansimus in Ierusalem ".
JER|35|12|Et factum est verbum Domini ad Ieremiam dicens:
JER|35|13|" Haec dicit Dominus exercituum, Deus Israel: Vade et dic viris Iudae et habitatoribus Ierusalem: Numquid non recipietis disciplinam, ut oboediatis verbis meis?, dicit Dominus.
JER|35|14|Praevaluerunt sermones Ionadab filii Rechab, quos praecepit filiis suis, ut non biberent vinum, et non biberunt usque ad diem hanc, quia oboedierunt praecepto patris sui; ego autem locutus sum ad vos de mane consurgens et loquens, et non oboedistis mihi.
JER|35|15|Misique ad vos omnes servos meos prophetas, consurgens diluculo mittensque et dicens: Convertimini unusquisque a via sua pessima et bona facite opera vestra et nolite sequi deos alienos neque colatis eos, et habitabitis in terra, quam dedi vobis et patribus vestris, et non inclinastis aurem vestram neque audistis me.
JER|35|16|Firmaverunt igitur filii Ionadab filii Rechab praeceptum patris sui, quod praeceperat eis; populus autem iste non oboedivit mihi.
JER|35|17|Idcirco haec dicit Dominus exercituum, Deus Israel: Ecce ego adducam super Iudam et super omnes habitatores Ierusalem universam afflictionem, quam locutus sum adversum illos, eo quod locutus sum ad illos, et non audierunt, vocavi illos, et non responderunt mihi ".
JER|35|18|Domui autem Rechabitarum dixit Ieremias: " Haec dicit Dominus exercituum, Deus Israel: Pro eo quod oboedistis praecepto Ionadab patris vestri et custodistis omnia mandata eius et fecistis universa, quae praecepit vobis,
JER|35|19|propterea haec dicit Dominus exercituum, Deus Israel: Non deficiet vir de stirpe Ionadab filii Rechab stans in conspectu meo cunctis diebus ".
JER|36|1|Et factum est in anno quarto Ioachim filii Iosiae regis Iudae, factum est verbum hoc ad Ieremiam a Domino dicens:
JER|36|2|" Tolle volumen libri et scribes in eo omnia verba, quae locutus sum tibi adversum Israel et Iudam et adversum omnes gentes a die qua locutus sum ad te ex diebus Iosiae usque ad diem hanc,
JER|36|3|si forte, audiente domo Iudae universa mala, quae ego cogito facere eis, revertatur unusquisque a via sua pessima, et propitius ero iniquitati et peccato eorum ".
JER|36|4|Vocavit ergo Ieremias Baruch filium Neriae; et scripsit Baruch ex ore Ieremiae omnes sermones Domini, quos locutus est ad eum, in volumine libri.
JER|36|5|Et praecepit Ieremias Baruch dicens: " Ego impeditus sum nec valeo ingredi domum Domini.
JER|36|6|Ingredere ergo tu et lege de volumine, in quo scripsisti ex ore meo verba Domini, audiente populo in domo Domini, in die ieiunii; insuper et audiente universo Iuda, qui veniunt de civitatibus suis, leges eis,
JER|36|7|si forte cadat oratio eorum in conspectu Domini, et revertatur unusquisque a via sua pessima, quoniam magnus furor et indignatio est, quam locutus est Dominus adversus populum hunc ".
JER|36|8|Et fecit Baruch filius Neriae iuxta omnia, quae praeceperat ei Ieremias propheta, legens ex volumine sermones Domini in domo Domini.
JER|36|9|Factum est autem in anno quinto Ioachim filii Iosiae regis Iudae, in mense nono, praedicaverunt ieiunium in conspectu Domini omni populo in Ierusalem et universae multitudini, quae confluxerat de civitatibus Iudae in Ierusalem.
JER|36|10|Legitque Baruch ex volumine sermones Ieremiae in domo Domini, in exedra Gamariae filii Saphan scribae in vestibulo superiore, in introitu portae Novae domus Domini, audiente omni populo.
JER|36|11|Cumque audisset Michaeas filius Gamariae filii Saphan omnes sermones Domini ex libro,
JER|36|12|descendit in domum regis ad exedram scribae; et ecce ibi omnes principes sedebant: Elisama scriba et Dalaias filius Semiae et Elnathan filius Achobor et Gamarias filius Saphan et Sedecias filius Hananiae et universi principes.
JER|36|13|Et nuntiavit eis Michaeas omnia verba, quae audivit, legente Baruch ex volumine in auribus populi.
JER|36|14|Miserunt itaque omnes principes ad Baruch Iudi filium Nathaniae filii Selemiae filii Chusi dicentes: " Volumen, ex quo legisti audiente populo, sume in manu tua et veni ". Tulit ergo Baruch filius Neriae volumen in manu sua et venit ad eos.
JER|36|15|Et dixerunt ad eum: " Sede et lege haec in auribus nostris "; et legit Baruch in auribus eorum.
JER|36|16|Igitur cum audissent omnia verba, obstupuerunt unusquisque ad proximum suum; et dixerunt ad Baruch: "Nuntiare debemus regi omnes sermones istos".
JER|36|17|Et interrogaverunt Baruch dicentes: " Indica nobis, quomodo scripsisti omnes sermones istos ex ore eius ".
JER|36|18|Dixit autem eis Baruch: " Ex ore suo loquebatur ad me omnes sermones istos, et ego scribebam in volumine atramento ".
JER|36|19|Et dixerunt principes ad Baruch: " Vade et abscondere, tu et Ieremias, et nemo sciat, ubi sitis ".
JER|36|20|Et ingressi sunt ad regem in atrium, porro volumen deposuerunt in exedra Elisamae scribae; et nuntiaverunt audiente rege omnes sermones.
JER|36|21|Misitque rex Iudi, ut sumeret volumen; qui, tollens illud de exedra Elisamae scribae, legit audiente rege et universis principibus, qui stabant circa regem.
JER|36|22|Rex autem sedebat in domo hiemali in mense nono, et posita erat arula coram eo plena prunis;
JER|36|23|cumque legisset Iudi tres pagellas vel quattuor, scidit eas scalpello scribae et proiecit in ignem, qui erat super arulam, donec consumeretur omne volumen igni, qui erat in arula.
JER|36|24|Et non timuerunt neque sciderunt vestimenta sua rex et omnes servi eius, qui audierunt universos sermones istos.
JER|36|25|Verumtamen Elnathan et Dalaias et Gamarias instanter rogaverunt regem, ne combureret librum, et non audivit eos.
JER|36|26|Et praecepit rex Ierameel filio regis et Saraiae filio Azriel et Selemiae filio Abdeel, ut comprehenderent Baruch scribam et Ieremiam prophetam; abscondit autem eos Dominus.
JER|36|27|Et factum est verbum Domini ad Ieremiam, postquam combusserat rex volumen et sermones, quos scripserat Baruch ex ore Ieremiae, dicens:
JER|36|28|"Rursum tolle volumen aliud et scribe in eo omnes sermones priores, qui erant in primo volumine, quod combussit Ioachim rex Iudae.
JER|36|29|Et super Ioachim regem Iudae dices: Haec dicit Dominus: Tu combussisti volumen illud dicens: "Quare scripsisti in eo annuntians: Certe veniet rex Babylonis et vastabit terram hanc et cessare faciet ex illa hominem et iumentum?".
JER|36|30|Propterea haec dicit Dominus contra Ioachim regem Iudae: Non erit ex eo, qui sedeat super solium David, et cadaver eius proicietur ad aestum per diem et ad gelu per noctem;
JER|36|31|et visitabo contra eum et contra semen eius et contra servos eius iniquitates suas; et adducam super eos et super habitatores Ierusalem et super viros Iudae omne malum, quod locutus sum ad eos, et non audierunt ".
JER|36|32|Ieremias autem tulit volumen aliud et dedit illud Baruch filio Neriae scribae; qui scripsit in eo ex ore Ieremiae omnes sermones libri, quem combusserat Ioachim rex Iudae igni; et insuper additi sunt multi sermones similes illis.
JER|37|1|Et regnavit rex Sedecias filius Iosiae pro Iechonia filio Ioachim; quem constituit regem Nabuchodonosor rex Babylonis in terra Iudae.
JER|37|2|Et non oboedivit, ipse et servi eius et populus terrae, verbis Domini, quae locutus est in manu Ieremiae prophetae.
JER|37|3|Et misit rex Sedecias Iuchal filium Selemiae et Sophoniam filium Maasiae sacerdotem ad Ieremiam prophetam dicens: " Ora pro nobis Dominum Deum nostrum ".
JER|37|4|Ieremias autem libere ambulabat in medio populi; non enim miserant eum in custodiam carceris.
JER|37|5|Igitur exercitus pharaonis egressus est de Aegypto, et audientes Chaldaei, qui obsidebant Ierusalem, huiuscemodi nuntium recesserunt ab Ierusalem.
JER|37|6|Et factum est verbum Domini ad Ieremiam prophetam dicens:
JER|37|7|" Haec dicit Dominus, Deus Israel: Sic dicetis regi Iudae, qui misit vos ad me interrogandum: Ecce exercitus pharaonis, qui egressus est vobis in auxilium, revertetur in terram suam in Aegyptum;
JER|37|8|et redient Chaldaei et bellabunt contra civitatem hanc et capient eam et succendent eam igni.
JER|37|9|Haec dicit Dominus: Nolite decipere animas vestras dicentes: "Euntes abibunt et recedent a nobis Chaldaei", quia non abibunt.
JER|37|10|Sed et si percusseritis omnem exercitum Chaldaeorum, qui proeliantur adversum vos, et derelicti fuerint ex eis aliqui vulnerati, singuli de tentorio suo consurgent et incendent civitatem hanc igni ".
JER|37|11|Ergo cum recessisset exercitus Chaldaeorum ab Ierusalem propter exercitum pharaonis,
JER|37|12|egressus est Ieremias de Ierusalem, ut iret in terram Beniamin et divideret ibi possessionem in conspectu populi.
JER|37|13|Cumque pervenisset ad portam Beniamin, erat ibi custos portae nomine Ierias filius Selemiae filii Hananiae; et apprehendit Ieremiam prophetam dicens: " Ad Chaldaeos profugis ".
JER|37|14|Et respondit Ieremias: " Falsum est! Non fugio ad Chaldaeos ". Et non audivit eum; sed comprehendit Ierias Ieremiam et adduxit eum ad principes.
JER|37|15|Et irati sunt principes contra Ieremiam, quem caesum miserunt in carcerem, qui erat in domo Ionathan scribae; eam enim in carcerem fecerant.
JER|37|16|Itaque ingressus est Ieremias in domum laci fornice tectam; et sedit ibi Ieremias diebus multis.
JER|37|17|Mittens autem Sedecias rex tulit eum et interrogavit eum in domo sua abscondite et dixit: " Putasne est sermo a Domino? ". Et dixit Ieremias: " Est "; et ait: "In manus regis Babylonis traderis ".
JER|37|18|Et dixit Ieremias ad regem Sedeciam: " Quid peccavi tibi et servis tuis et populo isti, quia misistis me in domum carceris?
JER|37|19|Ubi sunt prophetae vestri, qui prophetabant vobis et dicebant: "Non veniet rex Babylonis super vos et super terram hanc"?
JER|37|20|Nunc ergo audi, obsecro, domine mi rex; valeat deprecatio mea in conspectu tuo, et ne me remittas in domum Ionathan scribae, ne moriar ibi.
JER|37|21|Praecepit ergo rex Sedecias, ut traderetur Ieremias in vestibulo custodiae, et daretur ei torta panis cotidie ex vico Pistorum, donec consumerentur omnes panes de civitate. Et mansit Ieremias in vestibulo custodiae.
JER|38|1|Audivit autem Saphatias fi lius Matthan et Godolias fi lius Phassur et Iuchal filius Selemiae et Phassur filius Melchiae sermones, quos Ieremias loquebatur ad omnem populum dicens:
JER|38|2|" Haec dicit Dominus: Quicumque manserit in civitate hac, morietur gladio et fame et peste; qui autem profugerit ad Chaldaeos, vivet, et erit anima eius quasi spolium et vivet.
JER|38|3|Haec dicit Dominus: Certe tradetur civitas haec in manu exercitus regis Babylonis, et capiet eam ".
JER|38|4|Et dixerunt principes regi: " Rogamus, ut occidatur homo iste; de industria enim dissolvit manus virorum bellantium, qui remanserunt in civitate hac, et manus universi populi loquens ad eos iuxta verba haec; siquidem homo iste non quaerit pacem populo huic sed malum ".
JER|38|5|Et dixit rex Sedecias: " Ecce ipse in manibus vestris est; nequit enim rex vobis quidquam negare ".
JER|38|6|Tulerunt ergo Ieremiam et proiecerunt eum in lacum Melchiae filii regis, qui erat in vestibulo custodiae. Et submiserunt Ieremiam funibus. Et in lacu non erat aqua sed lutum; descendit itaque Ieremias in caenum.
JER|38|7|Audivit autem Abdemelech Aethiops, vir eunuchus, qui erat in domo regis, quod misissent Ieremiam in lacum; porro rex sedebat in porta Beniamin.
JER|38|8|Et egressus est Abdemelech de domo regis et locutus est ad regem dicens:
JER|38|9|" Domine mi rex, malefecerunt viri isti omnia, quaecumque perpetrarunt contra Ieremiam prophetam, mittentes eum in lacum, ut moriatur ibi fame; non sunt enim panes ultra in civitate ".
JER|38|10|Praecepit itaque rex Abdemelech Aethiopi dicens: " Tolle tecum hinc triginta viros et leva Ieremiam prophetam de lacu, antequam moriatur ".
JER|38|11|Assumptis ergo Abdemelech secum viris, ingressus est domum regis, in conclave, quod erat sub thesauro, et tulit inde pannos ex vestibus veteribus et scissis et submisit eos ad Ieremiam in lacum per funiculos.
JER|38|12|Dixitque Abdemelech Aethiops ad Ieremiam: " Pone veteres pannos et haec scissa sub scapuli et postea funes ". Fecit ergo Ieremias sic;
JER|38|13|et extraxerunt Ieremiam funibus et eduxerunt eum de lacu. Mansit autem Ieremias in vestibulo custodiae.
JER|38|14|Et misit rex Sedecias et tulit ad se Ieremiam prophetam ad ostium tertium, quod erat in domo Domini; et dixit rex ad Ieremiam: "Interrogo ego te sermonem, ne abscondas a me aliquid ".
JER|38|15|Dixit autem Ieremias ad Sedeciam: " Si annuntiavero tibi, numquid non interficies me? Et si consilium dedero tibi, non me audies ".
JER|38|16|Iuravit ergo rex Sedecias Ieremiae clam dicens: " Vivit Dominus, qui fecit nobis animam hanc, non occidam te et non tradam te in manu virorum istorum, qui quaerunt animam tuam ".
JER|38|17|Et dixit Ieremias ad Sedeciam: " Haec dicit Dominus exercituum, Deus Israel: Si profectus exieris ad principes regis Babylonis, vivet anima tua, et civitas haec non succendetur igni, et salvus eris tu et domus tua;
JER|38|18|si autem non exieris ad principes regis Babylonis, tradetur civitas haec in manu Chaldaeorum, et succendent eam igni, et tu non effugies de manu eorum ".
JER|38|19|Et dixit rex Sedecias ad Ieremiam: " Sollicitus sum propter Iudaeos, qui transfugerunt ad Chaldaeos, ne forte tradar in manus eorum, et illudant mihi ".
JER|38|20|Respondit autem Ieremias: " Non te tradent; audi, quaeso, vocem Domini, quam ego loquor ad te, et bene tibi erit, et vivet anima tua.
JER|38|21|Quod si nolueris egredi, iste est sermo, quem ostendit mihi Dominus:
JER|38|22|Ecce omnes mulieres, quae remanserunt in domo regis Iudae, educentur ad principes regis Babylonis et ipsae dicent:Seduxerunt te et praevaluerunt adversum teviri pacifici tui;demersi sunt in caeno pedes tui,illi autem recesserunt a te".
JER|38|23|Et omnes uxores tuae et filii tui educentur ad Chaldaeos, et non effugies manus eorum, sed in manu regis Babylonis capieris; et civitatem hanc comburet igni ".
JER|38|24|Dixit ergo Sedecias ad Ieremiam: " Nullus sciat verba haec, et non morieris.
JER|38|25|Si autem audierint principes quia locutus sum tecum, et venerint ad te et dixerint tibi: "Indica nobis, quid locutus sis cum rege, ne celes nos, et non te interficiemus, et quid locutus est tecum rex",
JER|38|26|dices ad eos: "Prostravi ego preces meas coram rege, ne me reduci iuberet in domum Ionathan, et ibi morerer" ".
JER|38|27|Venerunt ergo omnes principes ad Ieremiam et interrogaverunt eum, et locutus est eis iuxta omnia verba, quae praeceperat ei rex; et cessaverunt ab eo: nihil enim fuerat auditum.
JER|38|28|Mansit vero Ieremias in vestibulo custodiae usque ad diem, quo capta est Ierusalem.Et factum est ut caperetur Ierusalem.
JER|39|1|Anno nono Sedeciae regis Iudae, mense decimo, venit Nabuchodonosor rex Babylonis et omnis exercitus eius ad Ierusalem et obsidebant eam.
JER|39|2|Undecimo autem anno Sedeciae, mense quarto, nona mensis, aperta est civitas;
JER|39|3|et ingressi sunt omnes principes regis Babylonis et sederunt in porta Media: Nergelsereser Samegarnabu, Sarsachim princeps eunuchorum, Nergelsereser princeps magorum et omnes reliqui principes regis Babylonis.
JER|39|4|Cumque vidisset eos Sedecias rex Iudae et omnes viri bellatores, fugerunt et egressi sunt nocte de civitate per viam horti regis et per portam, quae erat inter duos muros, et egressi sunt ad viam Arabae.
JER|39|5|Persecutus est autem eos exercitus Chaldaeorum; et comprehenderunt Sedeciam in campestribus Iericho et captum adduxerunt ad Nabuchodonosor regem Babylonis in Rebla, quae est in terra Emath; et locutus est ad eum iudicia.
JER|39|6|Et occidit rex Babylonis filios Sedeciae in Rebla in oculis eius, et omnes nobiles Iudae occidit rex Babylonis;
JER|39|7|oculos quoque Sedeciae eruit et vinxit eum compedibus, ut duceretur in Babylonem.
JER|39|8|Domum quoque regis et domum vulgi succenderunt Chaldaei igni; et murum Ierusalem subverterunt.
JER|39|9|Et reliquias populi, quae remanserant in civitate, et perfugas, qui transfugerant ad eum, et superfluos artificum, qui remanserant, transtulit Nabuzardan magister satellitum in Babylonem.
JER|39|10|Et de plebe pauperum, qui nihil penitus habebant, dimisit Nabuzardan magister satellitum in terra Iudae; et dedit eis vineas et agros in die illa.
JER|39|11|Praeceperat autem Nabuchodonosor rex Babylonis de Ieremia Nabuzardan magistro satellitum dicens:
JER|39|12|" Tolle illum et pone super eum oculos tuos nihilque ei mali facias, sed, ut voluerit, sic facies ei ".
JER|39|13|Misit ergo Nabuzardan princeps satellitum et Nabusezban princeps eunuchorum et Nergelsereser princeps magorum et omnes optimates regis Babylonis
JER|39|14|miserunt et tulerunt Ieremiam de vestibulo custodiae et tradiderunt eum Godoliae filio Ahicam filii Saphan, ut duceret domum. Et habitavit in populo.
JER|39|15|Ad Ieremiam autem factus fuerat sermo Domini, cum clausus esset in vestibulo custodiae, dicens:
JER|39|16|" Vade et dic Abdemelech Aethiopi dicens: Haec dicit Dominus exercituum, Deus Israel: Ecce ego inducam sermones meos super civitatem hanc in malum et non in bonum; et erunt in conspectu tuo in die illa.
JER|39|17|Et liberabo te in die illa, ait Dominus, et non traderis in manus virorum, quos tu formidas;
JER|39|18|sed eruens liberabo te, et gladio non cades, sed erit tibi anima tua quasi spolium, quia in me habuisti fiduciam ", ait Dominus.
JER|40|1|Sermo, qui factus est ad Ieremiam a Domino, postquam dimissus est a Nabuzardan magistro satellitum de Rama, quando tulit eum vinctum catenis in medio omnium, qui migrabant de Ierusalem et Iuda et ducebantur in Babylonem.
JER|40|2|Tollens ergo princeps satellitum Ieremiam, dixit ad eum: " Dominus Deus tuus locutus est malum hoc super locum istum
JER|40|3|et adduxit; et fecit Dominus, sicut locutus est, quia peccastis Domino et non audistis vocem eius, et factus est vobis sermo hic.
JER|40|4|Nunc ergo ecce solvi te hodie de catenis, quae sunt in manibus tuis. Si placet tibi, ut venias mecum in Babylonem, veni, et ponam oculos meos super te; si autem displicet tibi venire mecum in Babylonem, reside; ecce omnis terra in conspectu tuo est: quod elegeris et quo placuerit tibi ut vadas, illuc perge ".
JER|40|5|Cum nondum reverteretur, dixit: " Revertere ad Godoliam filium Ahicam filii Saphan, quem praeposuit rex Babylonis civitatibus Iudae; habita ergo cum eo in medio populi vel quocumque placuerit tibi ut vadas, vade ". Dedit quoque ei magister satellitum cibaria et munuscula et dimisit eum.
JER|40|6|Venit autem Ieremias ad Godoliam filium Ahicam in Maspha et habitavit cum eo in medio populi, qui relictus fuerat in terra.
JER|40|7|Cumque audissent omnes principes exercitus, qui dispersi fuerant per regiones, ipsi et viri eorum, quod praefecisset rex Babylonis Godoliam filium Ahicam terrae et quod commendasset ei viros et mulieres et parvulos et de pauperibus terrae, qui non fuerant translati in Babylonem,
JER|40|8|venerunt ad Godoliam in Maspha; Ismael, inquam, filius Nathaniae et Iohanan et Ionathan filii Caree et Saraia filius Thanehumeth et filii Ophi, qui erant de Netopha, et Iezonias filius Maachathi, ipsi et viri eorum.
JER|40|9|Et iuravit eis Godolias filius Ahicam filii Saphan et comitibus eorum dicens: "Nolite timere servire Chaldaeis; habitate in terra et servite regi Babylonis, et bene erit vobis.
JER|40|10|Ecce ego habito in Maspha, ut stem coram Chaldaeis, qui veniunt ad nos; vos autem colligite vindemiam et messem et oleum et condite in vasis vestris et manete in urbibus vestris, quas tenetis ".
JER|40|11|Sed et omnes Iudaei, qui erant in Moab et in filiis Ammon et in Edom et in universis regionibus, audito quod dedisset rex Babylonis reliquias in Iudaea et quod praeposuisset super eos Godoliam filium Ahicam filii Saphan,
JER|40|12|reversi sunt, inquam, omnes Iudaei de universis locis, ad quae profugerant, et venerunt in terram Iudae ad Godoliam in Maspha et collegerunt vinum et messem multam nimis.
JER|40|13|Iohanan autem filius Caree et omnes principes exercitus, qui dispersi fuerant in regionibus, venerunt ad Godoliam in Maspha
JER|40|14|et dixerunt ei: " Scito quod Baalis rex filiorum Ammon misit Ismael filium Nathaniae percutere animam tuam "; et non credidit eis Godolias filius Ahicam.
JER|40|15|Iohanan vero filius Caree dixit ad Godoliam seorsum in Maspha loquens: Ibo et percutiam Ismael filium Nathaniae, nullo sciente, ne interficiat animam tuam, et dissipentur omnes Iudaei, qui congregati sunt ad te, et peribunt reliquiae Iudae ".
JER|40|16|Et ait Godolias filius Ahicam ad Iohanan filium Caree: " Noli facere verbum hoc; falsum enim tu loqueris de Ismael ".
JER|41|1|Et factum est in mense septi mo, venit Ismael filius Nathaniae filii Elisama de semine regali et optimates regis et decem viri cum eo ad Godoliam filium Ahicam in Maspha; et comederunt ibi panes simul in Maspha.
JER|41|2|Surrexit autem Ismael filius Nathaniae et decem viri, qui cum eo erant, et percusserunt Godoliam filium Ahicam filii Saphan gladio; et interfecerunt eum, quem praefecerat rex Babylonis terrae.
JER|41|3|Omnes quoque Iudaeos, qui erant cum Godolia in Maspha, et Chaldaeos, qui reperti sunt ibi, et viros bellatores percussit Ismael.
JER|41|4|Secundo autem die postquam occiderat Godoliam, nullo adhuc sciente,
JER|41|5|venerunt viri de Sichem et de Silo et de Samaria, octoginta viri, rasi barba et scissis vestibus et incisi in cute, et munera et tus habebant in manu, ut offerrent in domo Domini.
JER|41|6|Egressus ergo Ismael filius Nathaniae in occursum eorum de Maspha, incedens et plorans ibat. Cum autem occurrisset eis, dixit ad eos: " Venite ad Godoliam filium Ahicam ".
JER|41|7|Qui cum venissent ad medium civitatis, interfecit eos Ismael filius Nathaniae et proiecit in medium laci, ipse et viri, qui erant cum eo.
JER|41|8|Decem autem viri reperti sunt inter eos, qui dixerunt ad Ismael: " Noli occidere nos, quia habemus thesauros in agro, frumenti et hordei et olei et mellis "; et cessavit et non interfecit eos cum fratribus suis.
JER|41|9|Lacus autem, in quem proiecerat Ismael omnia cadavera virorum, quos percussit, est lacus magnus, quem fecit rex Asa propter Baasa regem Israel; ipsum replevit Ismael filius Nathaniae occisis.
JER|41|10|Et captivas duxit Ismael omnes reliquias populi, qui erant in Maspha, filias regis et universum populum, qui remanserat in Maspha, quos commendaverat Nabuzardan princeps satellitum Godoliae filio Ahicam; et cepit eos Ismael filius Nathaniae et abiit, ut transiret ad filios Ammon.
JER|41|11|Audivit autem Iohanan filius Caree et omnes principes bellatorum, qui erant cum eo, omne malum, quod fecerat Ismael filius Nathaniae,
JER|41|12|et, assumptis universis viris, profecti sunt, ut bellarent adversum Ismael filium Nathaniae; et invenerunt eum ad aquas multas, quae sunt in Gabaon.
JER|41|13|Cumque vidisset omnis populus, qui erat cum Ismael, Iohanan filium Caree et universos principes bellatorum, qui erant cum eo, laetati sunt.
JER|41|14|Et omnis populus, quem ceperat Ismael in Maspha, reversus est et abiit ad Iohanan filium Caree;
JER|41|15|Ismael autem filius Nathaniae fugit cum octo viris a facie Iohanan et abiit ad filios Ammon.
JER|41|16|Tulit ergo Iohanan filius Caree et omnes principes bellatorum, qui erant cum eo, universas reliquias vulgi, quas reduxerat ab Ismael filio Nathaniae venientes de Maspha, postquam percussit Godoliam filium Ahicam, viros fortes ad proelium et mulieres et pueros et eunuchos, quos reduxerat de Gabaon.
JER|41|17|Et abierunt et sederunt in Gherutchamaam, quae est iuxta Bethlehem, ut pergerent et introirent Aegyptum
JER|41|18|a facie Chaldaeorum; timebant enim eos, quia percusserat Ismael filius Nathaniae Godoliam filium Ahicam, quem praeposuerat rex Babylonis in regione.
JER|42|1|Et accesserunt omnes princi pes bellatorum, scilicet Iohanan filius Caree et Iezonias filius Osaiae et universum vulgus, a parvo usque ad magnum,
JER|42|2|dixeruntque ad Ieremiam prophetam: " Cadat oratio nostra in conspectu tuo, et ora pro nobis ad Dominum Deum tuum pro universis reliquiis istis, quia derelicti sumus pauci de pluribus, sicut oculi tui nos intuentur;
JER|42|3|et annuntiet nobis Dominus Deus tuus viam, per quam pergamus, et verbum, quod faciamus ".
JER|42|4|Dixit autem ad eos Ieremias propheta: " Audivi. Ecce ego oro ad Dominum Deum vestrum secundum verba vestra; omne verbum, quodcumque responderit pro vobis, indicabo vobis nec celabo vos quidquam ".
JER|42|5|Et illi dixerunt ad Ieremiam: " Sit Dominus inter nos testis verax et fidelis, si non iuxta omne verbum, in quo miserit te Dominus Deus tuus ad nos, sic faciemus.
JER|42|6|Sive bonum est sive malum, voci Domini Dei nostri, ad quem mittimus te, oboediemus, ut bene sit nobis, cum audierimus vocem Domini Dei nostri ".
JER|42|7|Cum autem completi essent decem dies, factum est verbum Domini ad Ieremiam;
JER|42|8|vocavitque Iohanan filium Caree et omnes principes bellatorum, qui erant cum eo, et universum populum a minimo usque ad magnum
JER|42|9|et dixit ad eos: " Haec dicit Dominus, Deus Israel, ad quem misistis me, ut prosternerem preces vestras in conspectu eius:
JER|42|10|Si quiescentes manseritis in terra hac, aedificabo vos et non destruam, plantabo et non evellam; iam enim placatus sum super malo, quod feci vobis.
JER|42|11|Nolite timere a facie regis Babylonis, quem vos pavidi formidatis; nolite metuere eum, dicit Dominus, quia vobiscum sum ego, ut salvos vos faciam et eruam de manu eius;
JER|42|12|et dabo vobis, ut misericordiam inveniatis, et ipse miserebitur vestri et habitare vos faciet in terra vestra.
JER|42|13|Si autem dixeritis vos: "Non habitabimus in terra ista", nec audieritis vocem Domini Dei vestri
JER|42|14|dicentes: "Nequaquam, sed ad terram Aegypti pergemus, ubi non videbimus bellum et clangorem tubae non audiemus et famem non sustinebimus et ibi habitabimus",
JER|42|15|propter hoc nunc audite verbum Domini, reliquiae Iudae: Haec dicit Dominus exercituum, Deus Israel: Si posueritis faciem vestram, ut ingrediamini Aegyptum, et intraveritis, ut ibi peregrinemini,
JER|42|16|gladius, quem vos formidatis, ibi comprehendet vos in terra Aegypti, et fames, pro qua estis solliciti, adhaerebit vobis in Aegypto, et ibi moriemini.
JER|42|17|Omnesque viri, qui posuerunt faciem suam, ut ingrediantur Aegyptum et peregrinentur ibi, morientur gladio et fame et peste: nullus de eis remanebit nec effugiet a facie mali, quod ego afferam super eos.
JER|42|18|Quia haec dicit Dominus exercituum, Deus Israel: Sicut effusus est furor meus et indignatio mea super habitatores Ierusalem, sic effundetur indignatio mea super vos, cum ingressi fueritis Aegyptum, et eritis in exsecrationem et in stuporem et in maledictum et in opprobrium et nequaquam ultra videbitis locum istum ".
JER|42|19|Verbum Domini super vos, reliquiae Iudae: " Nolite intrare Aegyptum; scientes scietis quia obtestatus sum vos hodie,
JER|42|20|quia decepistis animas vestras. Vos enim misistis me ad Dominum Deum nostrum dicentes: "Ora pro nobis ad Dominum Deum nostrum et iuxta omnia, quaecumque dixerit tibi Dominus Deus noster, sic annuntia nobis, et faciemus".
JER|42|21|Et annuntiavi vobis hodie, et non audistis vocem Domini Dei vestri super universis, pro quibus misit me ad vos.
JER|42|22|Nunc ergo scientes scietis quia gladio et fame et peste moriemini in loco, ad quem voluistis intrare et ibi peregrinari ".
JER|43|1|Factum est autem, cum complesset Ieremias loquens ad populum universos sermones Domini Dei eorum, pro quibus miserat eum Dominus Deus eorum ad illos omnia verba haec,
JER|43|2|dixit Azarias filius Osaiae et Iohanan filius Caree et omnes viri superbi dicentes ad Ieremiam: " Mendacium tu loqueris; non misit te Dominus Deus noster dicens: "Ne ingrediamini Aegyptum, ut illic peregrinemini",
JER|43|3|sed Baruch filius Neriae incitat te adversum nos, ut tradat nos in manu Chaldaeorum, ut interficiant nos et traducant in Babylonem ".
JER|43|4|Et non audivit Iohanan filius Caree et omnes principes bellatorum et universus populus vocem Domini, ut manerent in terra Iudae.
JER|43|5|Sed tollens Iohanan filius Caree et universi principes bellatorum universos reliquiarum Iudae, qui reversi fuerant de cunctis gentibus, ad quas fuerant ante dispersi, ut peregrinarentur in terra Iudae,
JER|43|6|viros et mulieres et parvulos et filias regis et omnem animam, quam reliquerat Nabuzardan princeps satellitum cum Godolia filio Ahicam filii Saphan, et Ieremiam prophetam et Baruch filium Neriae,
JER|43|7|et ingressi sunt terram Aegypti, quia non oboedierunt voci Domini; et venerunt usque ad Taphnas.
JER|43|8|Et factus est sermo Domini ad Ieremiam in Taphnis dicens:
JER|43|9|" Sume lapides grandes in manu tua et absconde eos in caemento, sub pavimento, quod est ad portam domus pharaonis in Taphnis, cernentibus viris Iudaeis;
JER|43|10|et dices ad eos: Haec dicit Dominus exercituum, Deus Israel: Ecce ego mittam et assumam Nabuchodonosor regem Babylonis servum meum et ponam thronum eius super lapides istos, quos abscondi, et statuet solium suum super eos;
JER|43|11|veniensque percutiet terram Aegypti, quos in mortem, in mortem et, quos in captivitatem, in captivitatem et, quos in gladium, in gladium;
JER|43|12|et succendet ignem in delubris deorum Aegypti et comburet ea et captivos ducet illos et excutiet terram Aegypti, sicut pastor pediculis excutit pallium suum, et egredietur inde in pace;
JER|43|13|et conteret statuas domus Solis, quae sunt in terra Aegypti, et delubra deorum Aegypti comburet igni ".
JER|44|1|Verbum, quod factum est per Ieremiam ad omnes Iudaeos, qui habitabant in terra Aegypti, habitantes in Magdolo et in Taphnis et in Memphi et in terra Phatures, dicens:
JER|44|2|" Haec dicit Dominus exercituum, Deus Israel: Vos vidistis omne malum istud, quod adduxi super Ierusalem et super omnes urbes Iudae; et ecce desertae sunt hodie, et non est in eis habitator
JER|44|3|propter malitiam, quam fecerunt, ut me ad iracundiam provocarent et irent, ut sacrificarent et colerent deos alienos, quos nesciebant et illi et vos et patres vestri.
JER|44|4|Et misi ad vos omnes servos meos prophetas, de nocte consurgens mittensque et dicens: Nolite facere verbum abominationis huiuscemodi, quam odivi.
JER|44|5|Et non audierunt nec inclinaverunt aurem suam, ut converterentur a malis suis et non sacrificarent diis alienis;
JER|44|6|et effusa est indignatio mea et furor meus et succensa est in civitatibus Iudae et in plateis Ierusalem, et versae sunt in solitudinem et vastitatem secundum diem hanc.
JER|44|7|Et nunc haec dicit Dominus exercituum, Deus Israel: Quare vos facitis malum grande contra animas vestras, ut intereat ex vobis vir et mulier, parvulus et lactans de medio Iudae, nec relinquatur vobis quidquam residuum,
JER|44|8|provocantes me in operibus manuum vestrarum, sacrificando diis alienis in terra Aegypti, in quam ingressi estis, ut ibi peregrinemini, et dissipet vos, et sitis in maledictionem et in opprobrium cunctis gentibus terrae?
JER|44|9|Numquid obliti estis mala patrum vestrorum et mala regum Iudae et mala uxorum eius et mala vestra et mala uxorum vestrarum, quae fecerunt in terra Iudae et in plateis Ierusalem?
JER|44|10|Non sunt contriti usque ad diem hanc et non timuerunt et non ambulaverunt in lege mea et in praeceptis meis, quae dedi coram vobis et coram patribus vestris.
JER|44|11|Ideo haec dicit Dominus exercituum, Deus Israel: Ecce ego ponam faciem meam in vobis in malum et disperdam omnem Iudam.
JER|44|12|Et assumam reliquias Iudae, qui posuerunt facies suas, ut ingrederentur terram Aegypti et peregrinarentur ibi, et consumentur omnes in terra Aegypti: cadent in gladio et in fame et consumentur a minimo usque ad maximum, in gladio et in fame morientur; et erunt in exsecrationem et in stuporem et in maledictionem et in opprobrium.
JER|44|13|Et visitabo super habitatores terrae Aegypti, sicut visitavi super Ierusalem, in gladio et in fame et in peste:
JER|44|14|et non erit qui effugiat et sit residuus de reliquiis Iudaeorum, qui venerunt, ut peregrinarentur in terra Aegypti et reverterentur in terram Iudae, ad quam ipsi elevant animas suas, ut revertantur et habitent ibi; non revertentur, nisi qui fugerint ".
JER|44|15|Responderunt autem Ieremiae omnes viri, scientes quod sacrificarent uxores eorum diis alienis, et universae mulieres, quarum stabat multitudo grandis, et omnis populus habitantium in terra Aegypti in Phatures, dicentes:
JER|44|16|" Sermonem, quem locutus es ad nos in nomine Domini, non audiemus ex te,
JER|44|17|sed facientes faciemus omne verbum, quod egressum est de ore nostro, ut sacrificemus reginae caeli et libemus ei libamina, sicut fecimus nos et patres nostri, reges nostri et principes nostri in urbibus Iudae et in plateis Ierusalem, et saturati sumus panibus et bene nobis erat malumque non vidimus.
JER|44|18|Ex eo autem tempore, quo cessavimus sacrificare reginae caeli et libare ei libamina, indigemus omnibus et gladio et fame consumpti sumus.
JER|44|19|Quod si nos sacrificamus reginae caeli et libamus ei libamina, numquid sine viris nostris fecimus ei placentas ad effingendum eam et libandum ei libamina? ".
JER|44|20|Et dixit Ieremias ad omnem populum, adversum viros et adversum mulieres et adversum universam plebem, qui responderant ei verbum, dicens:
JER|44|21|" Numquid non sacrificium, quod sacrificastis in civitatibus Iudae et in plateis Ierusalem, vos et patres vestri, reges vestri et principes vestri et populus terrae, horum recordatus est Dominus, et ascendit super cor eius?
JER|44|22|Et non poterat Dominus ultra portare propter malitiam operum vestrorum et propter abominationes, quas fecistis; et facta est terra vestra in desolationem et in stuporem et in maledictum, eo quod non sit habitator, sicut est dies haec.
JER|44|23|Propterea quod sacrificaveritis et peccaveritis Domino et non audieritis vocem Domini et in lege et in praeceptis et in testimoniis eius non ambulaveritis, idcirco evenerunt vobis mala haec, sicut est dies haec.
JER|44|24|Dixit autem Ieremias ad omnem populum et ad universas mulieres: " Audite verbum Domini, omnis Iuda, qui estis in terra Aegypti.
JER|44|25|Haec dicit Dominus exercituum, Deus Israel, dicens: Vos et uxores vestrae locuti estis ore vestro et manibus vestris implestis dicentes: Faciamus vota nostra, quae vovimus, ut sacrificemus reginae caeli et libemus ei libamina". Implete vota vestra et opere perpetrate ea.
JER|44|26|Ideo audite verbum Domini, omnis Iuda, qui habitatis in terra Aegypti: Ecce ego iuravi in nomine meo magno, ait Dominus, quia nequaquam ultra vocabitur nomen meum ex ore omnis viri Iudae dicentis: "Vivit Dominus Deus", in omni terra Aegypti.
JER|44|27|Ecce ego vigilabo super eos in malum et non in bonum, et consumentur omnes viri Iudae, qui sunt in terra Aegypti, gladio et fame, donec penitus consumantur.
JER|44|28|Et, qui fugerint gladium, revertentur de terra Aegypti in terram Iudae, viri pauci, et scient omnes reliquiae Iudae, quae ingressae sunt terram Aegypti, ut peregrinarentur ibi, cuius sermo compleatur, meus an illorum.
JER|44|29|Et hoc vobis signum, ait Dominus, quod visitem ego super vos in loco isto, ut sciatis quia vere complebuntur sermones mei contra vos in malum.
JER|44|30|Haec dicit Dominus: Ecce ego tradam pharaonem Ophree, regem Aegypti, in manu inimicorum eius et in manu quaerentium animam illius, sicut tradidi Sedeciam regem Iudae in manu Nabuchodonosor regis Babylonis inimici sui et quaerentis animam eius ".
JER|45|1|Verbum, quod locutus est Ieremias propheta ad Baruch filium Neriae, cum scriberet verba haec in libro ex ore Ieremiae, anno quarto Ioachim filii Iosiae regis Iudae, dicens:
JER|45|2|" Haec dicit Dominus, Deus Israel, super te, Baruch.
JER|45|3|Dixisti: "Vae misero mihi, quoniam addidit Dominus dolorem maerori meo; laboravi in gemitu meo et requiem non inveni".
JER|45|4|Haec dices ad eum: Sic dicit Dominus: Ecce, quod aedificavi, ego destruo et, quod plantavi, ego evello, universam terram hanc;
JER|45|5|et tu quaeris tibi grandia? Noli quaerere, quia ecce ego adducam malum super omnem carnem, ait Dominus, et dabo tibi animam tuam quasi spolium in omnibus locis, ad quaecumque perrexeris ".
JER|46|1|Quod factum est verbum Domini ad Ieremiam prophetam contra gentes.
JER|46|2|Ad Aegyptum.Adversum exercitum pharaonis Nechao regis Aegypti, qui erat iuxta fluvium Euphraten in Charchamis, quem percussit Nabuchodonosor rex Babylonis in quarto anno Ioachim filii Iosiae regis Iudae.
JER|46|3|" Praeparate scutum et clipeumet procedite ad bellum.
JER|46|4|Iungite equos et ascendite, equites;state in galeis, polite lanceas, induite vos loricis.
JER|46|5|Quid igitur? Vidi ipsos pavidos et terga vertentes,fortes eorum caesos;fugerunt conciti nec respexerunt:terror undique,ait Dominus.
JER|46|6|Non fugiat velox,nec salvari se putet fortis;ad aquilonem iuxta flumen Euphratenvicti sunt et ruerunt.
JER|46|7|Quis est iste, qui quasi Nilus ascendit,et veluti fluviorum intumescunt gurgites eius?
JER|46|8|Aegyptus Nili instar ascendit,et velut flumina moventur fluctus eius,et dixit: "Ascendens operiam terram,perdam civitatem et habitatores eius".
JER|46|9|Ascendite, equi, et irruite, currus;et procedant fortes,Aethiopia et Phut tenentes scutum et Ludii arripientes et iacientes sagittas.
JER|46|10|Dies autem ille Domini, Dei exercituum, dies ultionis,ut sumat vindictam de inimicis suis: devorat gladius, et saturatur,et inebriatur sanguine eorum;victima enim Domini, Dei exercituum,in terra aquilonis iuxta flumen Euphraten.
JER|46|11|Ascende in Galaad et tolle resinam,virgo filia Aegypti;frustra multiplicas medicamina,tibi vero cicatrix non obducitur.
JER|46|12|Audierunt gentes ignominiam tuam, et ululatus tuus replevit terram,quia fortis impegit in fortem,et ambo pariter conciderunt ".
JER|46|13|Verbum, quod locutus est Dominus ad Ieremiam prophetam super eo quod veniret Nabuchodonosor rex Babylonis percussurus terram Aegypti.
JER|46|14|" Annuntiate Aegyptoet auditum facite in Magdolo,et resonet in Memphi et in Taphnis,dicite: "Sta et praepara te,quia devoravit gladius ea,quae per circuitum tuum sunt".
JER|46|15|Quare deiectus est fortis tuus?Non stetit, quoniam Dominus subvertit eum.
JER|46|16|Multiplicavit ruentes,ceciditque vir ad proximum suum, et dixerunt: "Surge,et revertamur ad populum nostrumet ad terram nativitatis nostrae,a facie gladii saevientis".
JER|46|17|Vocate nomen pharaonis regis Aegypti:Tumultum, qui praetermisit tempus opportunum.
JER|46|18|Vivo ego, inquit rex,Dominus exercituum nomen eius,quoniam sicut Thabor in montibuset sicut Carmelus ad mare veniet.
JER|46|19|Vasa transmigrationis fac tibi,habitatrix filia Aegypti,quia Memphis in solitudinem eritet destruetur et inhabitabilis erit.
JER|46|20|Vitula elegans atque formosa Aegyptus,stimulus ab aquilone venit ei.
JER|46|21|Mercennarii quoque eius,qui versabantur in medio eius quasi vituli saginati,versi sunt et fugerunt simulnec stare potuerunt,quia dies interfectionis eorum venit super eos,tempus visitationis eorum.
JER|46|22|Vox eius quasi serpentis sibilantis,quoniam cum exercitu properabunt et cum securibus venient ei,quasi caedentes ligna.
JER|46|23|Succiderunt saltum eius,ait Dominus,qui supputari non potest;multiplicati sunt enim super locustas,et non est eis numerus.
JER|46|24|Confusa est filia Aegyptiet tradita in manu populi aquilonis ".
JER|46|25|Dixit Dominus exercituum, Deus Israel: " Ecce ego visitabo super Amon de No et super pharaonem et super Aegyptum et super deos eius et super reges eius et super pharaonem et super eos, qui confidunt in eo;
JER|46|26|et dabo eos in manu quaerentium animam eorum et in manu Nabuchodonosor regis Babylonis et in manu servorum eius; et post haec habitabitur sicut diebus pristinis, ait Dominus.
JER|46|27|Et tu ne timeas, serve meus Iacob,et ne paveas, Israel,quia ecce ego salvum te faciam de longinquoet semen tuum de terra captivitatis eorum;et revertetur Iacob et requiescet,securus erit, et non erit qui exterreat eum.
JER|46|28|Et tu noli timere, serve meus Iacob,ait Dominus,quia tecum ego sum,quia ego consumam cunctas gentes, ad quas eieci te;te vero non consumam,sed castigabo te in iudicionec quasi innocenti parcam tibi ".
JER|47|1|Quod factum est verbum Domini ad Ieremiam prophe tam contra Philisthim, antequam percuteret pharao Gazam.
JER|47|2|Haec dicit Dominus: Ecce, aquae ascendunt ab aquiloneet erunt quasi torrens inundanset operient terram et plenitudinem eius,urbem et habitatores eius.Clamabunt homines,et ululabunt omnes habitatores terrae
JER|47|3|a strepitu ungularum fortium equorum eius,a commotione quadrigarum eiuset tumultu rotarum illius;non respexerunt patres filios, manibus dissolutis,
JER|47|4|pro adventu diei, in quo vastabuntur omnes Philisthim,et dissipabitur Tyro et Sidoni omnis superstes auxiliator:depopulatus est enim Dominus Philisthim,reliquias insulae Caphtor.
JER|47|5|Venit calvitium super Gazam,conticuit Ascalon;reliquiae Enacim,usquequo incidetis vos?
JER|47|6|O mucro Domini,usquequo non quiesces?Ingredere in vaginam tuam,refrigerare et sile.
JER|47|7|Quomodo quiescet,cum Dominus praeceperit ei adversus Ascalonemet adversus maritimas regionesibique condixerit illi? ".
JER|48|1|Ad Moab.Haec dicit Dominus exercituum, Deus Israel: Vae super Nabo, quoniam vastata est et confusa!Capta est Cariathaim, confusa est arx et tremuit.
JER|48|2|Non est ultra exsultatio in Moab;in Hesebon cogitaverunt malum contra eam:Venite et disperdamus eam de gente".Tu quoque, Madmen, conticesces, sequeturque te gladius.
JER|48|3|Vox clamoris de Oronaim:Vastitas et contritio magna".
JER|48|4|Contrita est Moab,auditum fecerunt clamorem usque ad Segor.
JER|48|5|Per ascensum enim Luithplorans ascendit in fletu,quoniam in descensu Oronaimhostes ululatum contritionis audierunt:
JER|48|6|"Fugite, salvate animas vestraset eritis quasi myricae in deserto".
JER|48|7|Pro eo enim quod habuisti fiduciamin operibus tuis et in thesauris tuis,tu quoque capieris;et ibit Chamos in transmigrationem,sacerdotes eius et principes eius simul.
JER|48|8|Et veniet praedo ad omnem urbem, et urbs nulla salvabitur;et peribit vallis, et dissipabuntur campestria,quoniam dixit Dominus.
JER|48|9|Date pennas ad volandum;et civitates eius desertae erunt et inhabitabiles.
JER|48|10|Maledictus, qui facit opus Domini neglegenter,et maledictus, qui prohibet gladium suum a sanguine.
JER|48|11|Securus fuit Moab ab adulescentia suaet requievit in faecibus suisnec transfusus est de vase in vaset in transmigrationem non abiit;idcirco permansit gustus eius in eo,et odor eius non est immutatus.
JER|48|12|Propterea, ecce, dies veniunt,dicit Dominus,et mittam ei stratores laguncularum;et sternent eumet vasa eius exhaurientet lagunculas eorum collident.
JER|48|13|Et confundetur Moab a Chamos, sicut confusa est domus Israel a Bethel, in qua habebat fiduciam.
JER|48|14|Quomodo dicitis: "Fortes sumuset viri robusti ad proeliandum"?
JER|48|15|Vastata est Moab,et ascenderunt civitates illius,et electi iuvenes eius descenderunt in occisionem,ait rex, Dominus exercituum nomen eius.
JER|48|16|Prope est interitus Moab ut veniat,et malum eius velociter accurret nimis.
JER|48|17|Lugete super eum,omnes, qui estis in circuitu eius;et universi, qui scitis nomen eius,dicite: "Quomodo confracta est virga fortis,baculus gloriosus?".
JER|48|18|Descende de gloria et sede in siti,habitatrix filia Dibon,quoniam vastator Moab ascendit ad te,dissipavit munitiones tuas.
JER|48|19|Ad viam sta et prospice,habitatrix Aroer;interroga fugientemet eam, quae evasit.Dic: "Quid accidit?".
JER|48|20|Confusus est Moab, quoniam victus est.Ululate et clamate;annuntiate in Arnon,quoniam vastatus est Moab.
JER|48|21|Et iudicium venit ad terram campestrem super Helon et super Iasa et super Mephaath
JER|48|22|et super Dibon et super Nabo et super Bethdeblathaim,
JER|48|23|et super Cariathaim et super Bethgamul et super Bethmaon
JER|48|24|et super Carioth et super Bosra et super omnes civitates terrae Moab, quae longe et quae prope sunt.
JER|48|25|Abscissum est cornu Moab,et brachium eius contritum est,ait Dominus.
JER|48|26|Inebriate eum, quoniam contra Dominum erectus est; et allidet manum Moab in vomitu suo, et erit in derisum etiam ipse.
JER|48|27|Nonne in derisum tibi fuit Israel? Num inter fures repertus est? Quotiescumque enim adversum illum loquebaris, caput movebas.
JER|48|28|Relinquite civitates et habitate in petra,habitatores Moab,et estote quasi columba nidificansin parietibus apertae voraginis.
JER|48|29|Audivimus superbiam Moab,superbus est valde;sublimitatem eius et arrogantiamet superbiam et altitudinem cordis eius.
JER|48|30|Ego scio, ait Dominus, iactantiam eius, et quod non sint rectae fabulationes, nec recta fecerint.
JER|48|31|Ideo super Moab eiulabo et super Moab universam clamabo, super viros Cirhareseth plorabitur.
JER|48|32|Plus quam in planctu Iazer plorabo tibi,vinea Sabama;propagines tuae transierunt mare,usque ad Iazer pervenerunt.Super messem tuam et vindemiam tuampraedo irruit.
JER|48|33|Ablata est laetitia et exsultatiode horto et de terra Moab,et vinum de torcularibus sustuli;nequaquam calcator uvaesolitum celeuma cantabit.
JER|48|34|De clamore Hesebon usque Eleale et Iasa dederunt vocem suam, a Segor usque ad Oronaim, ad Eglatselisiam; aquae quoque Nemrim pessimae erunt.
JER|48|35|Et auferam de Moab, ait Dominus, offerentem in excelsis et sacrificantem diis eius.
JER|48|36|Propterea cor meum ad Moab quasi tibia resonabit, et cor meum ad viros Cirhareseth dabit sonitum tibiarum; quia depositum, quod acquisierunt, periit.
JER|48|37|Omne enim caput calvitium et omnis barba rasa erit, in cunctis manibus incisiones et super lumbos cilicium.
JER|48|38|Super omnia tecta Moab et in plateis eius omnis planctus, quoniam contrivi Moab sicut vas, quod nemini placet, ait Dominus.
JER|48|39|Quomodo victa est, et ululaverunt? Quomodo vertit dorsum Moab et confusus est? Eritque Moab in derisum et in terrorem omnibus in circuitu suo.
JER|48|40|Haec dicit Dominus:Ecce quasi aquila volabitet extendet alas suas ad Moab.
JER|48|41|Capta sunt oppida,et munitiones comprehensae sunt,et erit cor fortium Moab in die illasicut cor mulieris parturientis.
JER|48|42|Et cessabit Moab esse populus,quoniam contra Dominum gloriatus est.
JER|48|43|Pavor et fovea et laqueus super te,o habitator Moab,dicit Dominus.
JER|48|44|Qui fugerit a facie pavoris, cadet in foveam,et, qui conscenderit de fovea, capietur laqueo;adducam enim super Moabannum visitationis eorum,ait Dominus.
JER|48|45|In umbra Hesebon steterunt sine viribus fugientes,sed ignis egressus est de Hesebon,et flamma de medio Sehon,et devoravit tempora Moabet verticem filiorum tumultus.
JER|48|46|Vae tibi, Moab!Periit populus Chamos,quia comprehensi sunt filii tuiet filiae tuae in captivitatem.
JER|48|47|Et convertam sortem Moab in novissimis diebus ",ait Dominus.Hucusque iudicia Moab.
JER|49|1|Ad filios Ammon.Haec dicit Dominus: Numquid filii non sunt Israel,aut heres non est ei?Cur igitur hereditate possedit Melchom Gad,et populus eius in urbibus eius habitavit?
JER|49|2|Ideo ecce dies veniunt,dicit Dominus,et auditum faciam super Rabba filiorum Ammonfremitum proelii;et erit in tumulum dissipata,filiaeque eius igni succendentur,et possidebit Israel possessores suos, ait Dominus.
JER|49|3|Ulula, Hesebon, quoniam vastata es, ut sis in acervum lapidum;clamate, filiae Rabba,accingite vos ciliciis, plangiteet circuite per muros,quoniam Melchom in transmigrationem ducetur,sacerdotes eius et principes eius simul.
JER|49|4|Quid gloriaris in vallibus?Copiose fluxit vallis tua, filia rebellis,quae confidebas in thesauris tuiset dicebas: "Quis veniet ad me?".
JER|49|5|Ecce ego inducam super te terrorem,ait Dominus, Deus exercituum,ab omnibus, qui sunt in circuitu tuo;et dispergemini singuli in viam suam,nec erit qui congreget fugientes.
JER|49|6|Et post haec convertamsortem filiorum Ammon ",ait Dominus.
JER|49|7|Ad Edom.Haec dicit Dominus exercituum: Numquid non ultra est sapientia in Theman?Periit consilium a prudentibus,inutilis facta est sapientia eorum.
JER|49|8|Fugite, terga vertite, descendite in voraginem,habitatores Dedan,quoniam perditionem Esau adduxi super eum,tempore quo visitavi eum.
JER|49|9|Si vindemiatores veniunt super te,non relinquent racemum;si fures in nocte,diripiunt, quod placet sibi.
JER|49|10|Ego vero discooperui Esau,revelavi abscondita eius,et celari non poterit;vastatum est semen eiuset fratres eius et vicini eius, et non erit.
JER|49|11|Relinque pupillos tuos, ego faciam eos vivere;et viduae tuae in me sperabunt.
JER|49|12|Quia haec dicit Dominus: Ecce quibus non erat iudicium, ut biberent calicem, bibentes bibent; et tu quasi innocens relinqueris? Non eris innocens, sed bibens bibes.
JER|49|13|Quia per memetipsum iuravi, dicit Dominus, quod in solitudinem et in opprobrium et in desertum et in maledictionem erit Bosra; et omnes civitates eius erunt in solitudines sempiternas ".
JER|49|14|Auditum audivi a Domino,et legatus ad gentes missus est: Congregamini et venite contra eamet consurgite in proelium ".
JER|49|15|" Ecce enim parvulum dedi te in gentibus,contemptibilem inter homines.
JER|49|16|Arrogantia tua decepit te,et superbia cordis tui,qui habitas in cavernis petraeet tenes altitudinem collis;cum exaltaveris quasi aquila nidum tuum,inde detraham te,dicit Dominus.
JER|49|17|Et erit Edom in desolationem: omnis, qui transibit per eam, stupebit et sibilabit super omnes plagas eius.
JER|49|18|Sicut subversa est Sodoma et Gomorra et vicinae eius, ait Dominus, non habitabit ibi vir, et non peregrinabitur in ea filius hominis.
JER|49|19|Ecce quasi leo ascendet de silva condensa Iordanis ad prata semper virentia, quia subito currere faciam eos ex illa; et, qui erit electus, illum praeponam ei. Quis enim similis mei? Et quis vocabit me in iudicium? Et quis est iste pastor, qui resistat vultui meo?
JER|49|20|Propterea audite consilium Domini, quod iniit de Edom, et cogitationes eius, quas cogitavit de habitatoribus Theman:Certe abstrahent parvulos gregis,certe desolabuntur super eos pascua eorum.
JER|49|21|A voce ruinae eorum commota est terra,clamor in mari Rubro auditus est ocis eius.
JER|49|22|Ecce quasi aquila ascendet et volabitet expandet alas suas super Bosram;et erit cor fortium Edom in die illaquasi cor mulieris parturientis ".
JER|49|23|Ad Damascum. Confusa est Emath et Arphad,quia auditum pessimum audierunt;turbati sunt in mari sollicitudinis,quod quiescere non potuit.
JER|49|24|Dissoluta est Damascus, versa in fugam;tremor apprehendit eam,angustia et dolores tenuerunt eamquasi parturientem.
JER|49|25|Quomodo non erit derelicta civitas laudabilis,urbs laetitiae?
JER|49|26|Ideo cadent iuvenes eius in plateis eius,et omnes viri proelii conticescent in die illa,ait Dominus exercituum.
JER|49|27|Et succendam ignem in muro Damasci,et devorabit moenia Benadad ".
JER|49|28|Ad Cedar et ad regna Asor, quae percussit Nabuchodonosor rex Babylonis.Haec dicit Dominus: Surgite, ascendite ad Cedaret vastate filios orientis.
JER|49|29|Tabernacula eorum et greges eorum capient;tentoria eorum et omnia vasa eorumet camelos eorum tollent sibi;et vocabunt super eos formidinem in circuitu.
JER|49|30|Fugite, abite vehementer,in voraginibus sedete,qui habitatis Asor,ait Dominus;iniit enim contra vosNabuchodonosor rex Babylonis consiliumet cogitavit adversum vos cogitationes.
JER|49|31|Consurgite, et ascenditead gentem quietam et habitantem confidenter,ait Dominus;non ostia nec vectes eis:soli habitant.
JER|49|32|Et erunt cameli eorum in direptionem,et multitudo iumentorum in praedam;et dispergam eos in omnem ventum, qui sunt attonsi in comam,et ex omni confinio eorumadducam interitum super eos,ait Dominus.
JER|49|33|Et erit Asor in habitaculum thoum,deserta usque in aeternum;non manebit ibi vir,nec peregrinabitur in ea filius hominis ".
JER|49|34|Quod factum est verbum Domini ad Ieremiam prophetam super Elam, in principio regni Sedeciae regis Iudae, dicens:
JER|49|35|" Haec dicit Dominus exercituum:Ecce ego confringam arcum Elam, summam fortitudinem eorum;
JER|49|36|et inducam super Elamquattuor ventos a quattuor plagis caeli,et ventilabo eos in omnes ventos istos,et non erit gens,ad quam non perveniant profugi Elam.
JER|49|37|Et pavere faciam Elam coram inimicis suiset in conspectu quaerentium animam eorum;et adducam super eos malumiram furoris mei,dicit Dominus,et mittam post eos gladium,donec consumam eos.
JER|49|38|Et ponam solium meum in Elamet perdam inde regem et principes, ait Dominus.
JER|49|39|In novissimis autem diebusconvertam sortem Elam ",dicit Dominus.
JER|50|1|Verbum, quod locutus est Dominus de Babylone et de terra Chaldaeorum in manu Ieremiae prophetae:
JER|50|2|" Annuntiate in gentibus et auditum facite,levate signum;praedicate et nolite celare, dicite:Capta est Babylon,confusus est Bel,victus est Merodach.Confusa sunt sculptilia eius,superata sunt idola eorum".
JER|50|3|Quoniam ascendit contra eam gens ab aquilone, quae ponet terram eius in solitudinem, et non erit qui habitet in ea ab homine usque ad pecus: et moti sunt et abierunt.
JER|50|4|In diebus illis et in tempore illo, ait Dominus, venient filii Israel ipsi et filii Iudae simul; ambulantes et flentes properabunt et Dominum Deum suum quaerent.
JER|50|5|De Sion interrogabunt, ad cuius viam facies eorum: "Venite, et apponamur ad Dominum foedere sempiterno, quod nulla oblivione delebitur".
JER|50|6|Grex perditus factus est populus meus, pastores eorum seduxerunt eos feceruntque vagari in montibus; de monte in collem transierunt, obliti sunt cubilis sui.
JER|50|7|Omnes, qui invenerunt, comederunt eos, et hostes eorum dixerunt: "Non delinquimus, pro eo quod peccaverunt Domino, habitaculo iustitiae et exspectationi patrum eorum Domino".
JER|50|8|Recedite de medio Babyloniset de terra Chaldaeorum egredimini;et estote quasi haedi ante gregem.
JER|50|9|Quoniam ecce ego suscito et adducam in Babylonemcongregationem gentium magnarumde terra aquilonis;et praeparabuntur adversus eam,et inde capietur:sagitta eorum quasi bellatoris electinon revertetur vacua.
JER|50|10|Et erit Chaldaea in praedam;omnes vastantes eam replebuntur ",ait Dominus.
JER|50|11|Dum exsultatis et magna loquiminidiripientes hereditatem meamdum effusi estis sicut vituli super herbamet hinnitis sicut equi fortes,
JER|50|12|confusa est mater vestra nimis,et in opprobrium facta est, quae genuit vos;ecce novissima erit in gentibus,deserta, invia et arens.
JER|50|13|Ab ira Domini non habitabitur,sed redigetur tota in solitudinem;omnis, qui transibit per Babylonem, stupebitet sibilabit super universis plagis eius.
JER|50|14|Praeparamini contra Babylonem per circuitumomnes, qui tenditis arcum;debellate eam, non parcatis iaculis,quia Domino peccavit.
JER|50|15|Clamate adversus eam;ubique dedit manum,ceciderunt fundamenta eius,destructi sunt muri eius,quoniam ultio Domini est;ultionem accipite de ea:sicut fecit, facite ei.
JER|50|16|Disperdite satorem de Babyloneet tenentem falcem in tempore messis;a facie gladii saevientisunusquisque ad populum suum convertetur,et singuli ad terram suam fugient.
JER|50|17|Ovis dispersa Israel;leones eiecerunt eum.Primus comedit eum rex Assyriae;iste novissimus exossavit eumNabuchodonosor rex Babylonis.
JER|50|18|Propterea haec dicit Dominus exercituum, Deus Israel: " Ecce ego visitabo regem Babylonis et terram eius, sicut visitavi regem Assyriae;
JER|50|19|et reducam Israel ad pascua sua, et pascetur Carmelum et Basan, et in monte Ephraim et Galaad saturabitur anima eius.
JER|50|20|In diebus illis et in tempore illo, ait Dominus, quaeretur iniquitas Israel et non erit, et peccatum Iudae et non invenietur, quoniam propitius ero eis, quos reliquero.
JER|50|21|Super terram Merataim ascendeet super habitatores Phacud.Dissipa et interfice persequens eos,ait Dominus,et fac iuxta omnia, quae praecepi tibi ".
JER|50|22|Vox belli in terraet contritio magna.
JER|50|23|Quomodo confractus est et contritusmalleus universae terrae?Quomodo versa est in desolationem Babylon in gentibus?
JER|50|24|Illaqueavi te, et capta es, Babylon,et nesciebas;inventa es et apprehensa,quoniam Dominum provocasti.
JER|50|25|Aperuit Dominus thesaurum suumet protulit vasa irae suae,quoniam opus est Domino Deo exercituumin terra Chaldaeorum.
JER|50|26|Venite ad eam ab extremis finibus,aperite horrea eius;redigite eam in acervos lapidum quasi manipuloset interficite eam,nec sit quidquam reliquum.
JER|50|27|Dissipate universos tauros eius,descendant in occisionem.Vae eis, quia venit dies eorum,tempus visitationis eorum!
JER|50|28|Vox fugientiumet eorum, qui evaserunt de terra Babylonis,ut annuntient in Sionultionem Domini Dei nostri,ultionem templi eius.
JER|50|29|Convocate in Babylonem sagittarios,omnes, qui tendunt arcum;consistite adversus eam per gyrum, et nullus evadat:reddite ei secundum opus suum,iuxta omnia, quae fecit, facite illi,quia contra Dominum erecta est,adversum Sanctum Israel.
JER|50|30|" Idcirco cadent iuvenes eius in plateis eius,et omnes viri bellatores eius conticescent in die illa,ait Dominus.
JER|50|31|Ecce ego ad te, Superbia,dicit Dominus, Deus exercituum,quia venit dies tuus,tempus visitationis tuae.
JER|50|32|Et cadet Superbia et corruet,et non erit qui suscitet eam;et succendam ignem in urbibus eius,et devorabit omnia in circuitu eius ".
JER|50|33|Haec dicit Dominus exercituum: " Calumniam sustinent filii Israel et filii Iudae simul; omnes, qui ceperunt eos, tenent, nolunt dimittere eos.
JER|50|34|Redemptor eorum fortis, Dominus exercituum nomen eius, iudicio defendet causam eorum, ut quietem det terrae et conturbet habitatores Babylonis.
JER|50|35|Gladius ad Chaldaeos,ait Dominus,et ad habitatores Babyloniset ad principes et ad sapientes eius!
JER|50|36|Gladius ad divinos eius, qui stulti erunt!Gladius ad fortes illius, qui timebunt!
JER|50|37|Gladius ad equos eius et ad currus eiuset ad omne vulgus, quod est in medio eius;et erunt quasi mulieres!Gladius ad thesauros eius, qui diripientur!
JER|50|38|Siccitas super aquas eius erit, et arescent,quia terra sculptilium est,et in portentis insaniunt.
JER|50|39|Propterea habitabunt dracones cum thoibus, et habitabunt in ea struthiones; et non inhabitabitur ultra usque in sempiternum nec exstruetur usque ad generationem et generationem.
JER|50|40|Sicut subvertit Deus Sodomam et Gomorram et vicinas eius, ait Dominus, non habitabit ibi vir, et non peregrinabitur in ea filius hominis.
JER|50|41|Ecce populus venit ab aquilone, et gens magna et reges multi consurgent a finibus terrae.
JER|50|42|Arcum et acinacem apprehendent, crudeles sunt et immisericordes; vox eorum quasi mare sonabit, et super equos ascendent sicut vir paratus ad proelium contra te, filia Babylon.
JER|50|43|Audivit rex Babylonis famam eorum, et dissolutae sunt manus eius; angustia apprehendit eum, dolor quasi parturientem.
JER|50|44|Ecce quasi leo ascendet de silva condensa Iordanis ad prata semper virentia, quia subito currere faciam eos ex illa et, qui erit electus, illum praeponam ei. Quis enim similis mei? Et quis vocabit me in iudicium? Et quis est iste pastor, qui resistat vultui meo? ".
JER|50|45|Propterea audite consilium Domini, quod mente concepit adversum Babylonem, et cogitationes eius, quas cogitavit super terram Chaldaeorum: certe abstrahent parvulos gregis, certe desolabuntur super eos pascua eorum.
JER|50|46|A voce captivitatis Babylonis commota est terra, et clamor inter gentes auditus est.
JER|51|1|Haec dicit Dominus: Ecce ego suscitabo super Babylonemet super habitatores Chaldaeaequasi ventum pestilentem;
JER|51|2|et mittam in Babylonem ventilatores,et ventilabunt eamet demolientur terram eius,quoniam venerunt super eam undiquein die afflictionis.
JER|51|3|Non tendat, qui tendit arcum suum,et non ascendat loricatus;nolite parcere iuvenibus eius,interficite omnem militiam eius ".
JER|51|4|Et cadent interfecti in terra Chaldaeorumet vulnerati in plateis eius,
JER|51|5|quoniam non est viduatus Israel et Iudaa Deo suo, Domino exercituum;terra autem eorum repleta est delictoin conspectu Sancti Israel.
JER|51|6|Fugite de medio Babylonis,et salvet unusquisque animam suam;nolite perire in poena eius,quoniam tempus ultionis est Domino:vicissitudinem ipse retribuet ei.
JER|51|7|Calix aureus Babylon in manu Dominiinebrians omnem terram;de vino eius biberunt genteset ideo insaniunt.
JER|51|8|Subito cecidit Babylon et contrita est.Ululate super eam;tollite resinam ad dolorem eius,si forte sanetur.
JER|51|9|" Curavimus Babylonem,et non est sanata.Derelinquite eam,et eamus unusquisque in terram suam,quoniam pervenit usque ad caelos iudicium eiuset elevatum est usque ad nubes.
JER|51|10|Protulit Dominus iustitias nostras;venite, et narremus in Sionopus Domini Dei nostri ".
JER|51|11|Acuite sagittas, implete pharetras;suscitavit Dominus spiritum regum Medorum,et contra Babylonem mens eius est, ut perdat eam,quoniam ultio Dominiest ultio templi sui.
JER|51|12|Super muros Babylonis levate signum,augete custodiam,ponite custodes, praeparate insidias,quia cogitavit Dominus,et facit quaecumque locutus estcontra habitatores Babylonis.
JER|51|13|Quae habitas super aquas multas,locuples in thesauris,venit finis tuus,pedalis praecisionis tuae.
JER|51|14|Iuravit Dominus exercituum per animam suam: Quoniam, etsi replevero te hominibus quasi brucho,super te celeuma cantabitur ".
JER|51|15|Qui fecit terram in fortitudine sua,praeparavit orbem in sapientia sua et prudentia sua extendit caelos;
JER|51|16|dante eo vocem, multiplicantur aquae in caelo;qui levat nubes ab extremo terrae,fulgura in pluviam facitet producit ventum de thesauris suis.
JER|51|17|Stultus factus est omnis homo, absque scientia;confusus est omnis conflator in sculptili,quia mendax conflatio eius,nec est spiritus in eis.
JER|51|18|Vana sunt opera et risu digna,in tempore visitationis suae peribunt.
JER|51|19|Non sicut haec pars Iacob,quia, qui fecit omnia, ipse est,et Israel tribus hereditatis eius:Dominus exercituum nomen eius.
JER|51|20|" Malleus tu mihi, vas belli:et ego collisi in te genteset dispersi in te regna
JER|51|21|et collisi in te equum et equitem eiuset collisi in te currum et ascensorem eius
JER|51|22|et collisi in te virum et mulieremet collisi in te senem et puerumet collisi in te iuvenem et virginem
JER|51|23|et collisi in te pastorem et gregem eiuset collisi in te agricolam et iugales eiuset collisi in te duces et magistratus.
JER|51|24|Et reddam Babyloni et cunctis habitatoribus Chaldaeae omne malum suum, quod fecerunt in Sion in oculis vestris, ait Dominus.
JER|51|25|Ecce ego ad te, mons pestifer,ait Dominus,qui corrumpis universam terram;et extendam manum meam super teet evolvam te de petriset dabo te in montem combustionis.
JER|51|26|Et non tollent de te lapidem in angulumet lapidem in fundamenta,sed perditus in aeternum eris ",ait Dominus.
JER|51|27|Levate signum in terra,clangite bucina in gentibus,sanctificate super eam gentes,vocate contra illam regnaArarat, Menni et Aschenez.Constituite super eam scribas,adducite equos quasi bruchum aculeatum.
JER|51|28|Sanctificate contra eam gentes, reges Mediae, duces eius et universos magistratus eius cunctamque terram potestatis eius.
JER|51|29|Et commovebitur terra et conturbabitur,quia impletur contra Babylonem cogitatio Domini,ut ponat terram Babylonisdesertam et inhabitabilem.
JER|51|30|Cessaverunt fortes Babylonis a proelio,habitaverunt in praesidiis;devoratum est robur eorum,et facti sunt quasi mulieres;incensa sunt tabernacula eius,contriti sunt vectes eius.
JER|51|31|Currens obviam currenti veniet,et nuntius obvius nuntianti,ut annuntiet regi Babylonisquia capta est civitas eiusa summo usque ad summum.
JER|51|32|Et vada praeoccupata sunt,et paludes incensae sunt igni;et viri bellatores conturbati sunt.
JER|51|33|Quia haec dicit Dominus exercituum, Deus Israel: Filia Babylonis quasi area tempore triturae eius;adhuc modicum, et veniet tempus messionis eius ".
JER|51|34|" Comedit me, devoravit me Nabuchodonosor;rex Babylonis reddidit me quasi vas inane,absorbuit me quasi draco,replevit ventrem suum deliciis meis et eiecit me ".
JER|51|35|" Iniquitas adversum me et caro mea super Babylonem! ",dicit habitatio Sion. Et sanguis meus super habitatores Chaldaeae! ",dicit Ierusalem.
JER|51|36|Propterea haec dicit Dominus: Ecce ego iudicabo causam tuamet ulciscar ultionem tuamet desertum faciam mare eiuset siccabo venam eius;
JER|51|37|et erit Babylon in tumulos,habitatio thoum,stupor et sibilus,eo quod non sit habitator.
JER|51|38|Simul ut leones rugient,frement veluti catuli leonum.
JER|51|39|In calore eorum ponam potus eorumet inebriabo eos, ut sopianturet dormiant somnum sempiternum et non consurgant,dicit Dominus.
JER|51|40|Deducam eos quasi agnos ad victimam,quasi arietes cum haedis ".
JER|51|41|Quomodo capta est Babel,et comprehensa est gloria universae terrae?Quomodo facta est in stuporemBabylon inter gentes?
JER|51|42|Ascendit super Babylonem mare,multitudine fluctuum eius operta est.
JER|51|43|Factae sunt civitates eius in stuporem,terra inhabitabilis et deserta,terra, in qua nullus habitet,nec transeat per eam filius hominis.
JER|51|44|" Et visitabo super Bel in Babyloneet eiciam, quod absorbuerat, de ore eius;et non confluent ad eum ultra gentes,siquidem et murus Babylonis corruet.
JER|51|45|Egredimini de medio eius, populus meus,ut salvet unusquisque animam suamab ira furoris Domini.
JER|51|46|Et ne forte mollescat cor vestrum, et timeatis auditum, qui audietur in terra; et veniet in anno auditio, et post hunc annum auditio, et iniquitas in terra, et dominator super dominatorem.
JER|51|47|Propterea ecce dies veniunt, et visitabo super sculptilia Babylonis, et omnis terra eius confundetur, et universi interfecti eius cadent in medio eius.
JER|51|48|Et laudabunt super Babylonem caeli et terra et omnia, quae in eis sunt, quia ab aquilone venient ei praedones, ait Dominus.
JER|51|49|Et Babylon cadet, occisi in Israel, sicut pro Babylone ceciderunt occisi universae terrae.
JER|51|50|Qui fugistis gladium, ite, nolite stare; recordamini procul Domini, et Ierusalem ascendat super cor vestrum.
JER|51|51|"Confusi sumus, quoniam audivimus opprobrium; operuit ignominia facies nostras, quia venerunt alieni super sanctificationem domus Domini".
JER|51|52|Propterea ecce dies veniunt, ait Dominus, et visitabo super sculptilia eius, et in omni terra eius gemet vulneratus.
JER|51|53|Si ascenderit Babylon in caelum et firmaverit in excelso robur suum, a me venient vastatores eius ", ait Dominus.
JER|51|54|Vox clamoris de Babylone et contritio magna de terra Chaldaeorum,
JER|51|55|quoniam vastavit Dominus Babylonem et perdidit ex ea vocem magnam; et sonabunt fluctus eorum quasi aquae multae, dedit sonitum vox eorum.
JER|51|56|Quia venit super eam, id est super Babylonem, praedo; et apprehensi sunt fortes eius, et fractus est arcus eorum, quia Deus ultor Dominus reddens retribuet.
JER|51|57|" Et inebriabo principes eius et sapientes eius et duces eius et magistratus eius et fortes eius; et dormient somnum sempiternum et non expergiscentur ", ait rex, Dominus exercituum nomen eius.
JER|51|58|Haec dicit Dominus exercituum: Murus Babylonis ille latissimus funditus suffodietur,et portae eius excelsae igni comburentur;et laboraverunt populi pro nihilo,et gentes pro igni lassatae sunt ".
JER|51|59|Verbum, quod praecepit Ieremias propheta Saraiae filio Neriae filii Maasiae, cum pergeret cum Sedecia rege Iudae in Babylonem in anno quarto regni eius; Saraias autem erat princeps, qui mansionibus praeerat.
JER|51|60|Et scripsit Ieremias omne malum, quod venturum erat super Babylonem, in libro uno, omnia verba haec, quae scripta sunt contra Babylonem.
JER|51|61|Et dixit Ieremias ad Saraiam: " Cum veneris in Babylonem et videris et legeris omnia verba haec,
JER|51|62|dices: "Domine, tu locutus es contra locum istum, ut disperderes eum, ne sit qui in eo habitet ab homine usque ad pecus, et ut sit perpetua solitudo".
JER|51|63|Cumque compleveris legere librum istum, ligabis ad eum lapidem et proicies illum in medium Euphraten
JER|51|64|et dices: "Sic submergetur Babylon et non consurget a facie afflictionis, quam ego adduco super eam, et dissolvetur" ".Hucusque verba Ieremiae.
JER|52|1|Filius viginti et unius anni erat Sedecias, cum regnare coepisset, et undecim annis regnavit in Ierusalem; et nomen matris eius Amital filia Ieremiae de Lobna.
JER|52|2|Et fecit malum in oculis Domini iuxta omnia, quae fecerat Ioachim,
JER|52|3|quoniam furor Domini erat in Ierusalem et in Iuda, usquequo proiceret eos a facie sua.Et recessit Sedecias a rege Babylonis.
JER|52|4|Factum est autem in anno nono regni eius, in mense decimo decima mensis, venit Nabuchodonosor rex Babylonis, ipse et omnis exercitus eius, adversus Ierusalem; et obsederunt eam et aedificaverunt contra eam munitiones in circuitu.
JER|52|5|Et fuit civitas obsessa usque ad undecimum annum regis Sedeciae.
JER|52|6|Mense autem quarto, nona mensis, obtinuit fames in civitate, et non erant alimenta populo terrae.
JER|52|7|Et dirupta est civitas, et omnes viri bellatores fugerunt exieruntque de civitate nocte per viam portae, quae est inter duos muros et ducit ad hortum regis, Chaldaeis obsidentibus urbem in gyro, et abierunt per viam, quae ducit in Arabam.
JER|52|8|Persecutus est autem Chaldaeorum exercitus regem, et apprehenderunt Sedeciam in campestribus Iericho, et omnis comitatus eius diffugit ab eo.
JER|52|9|Cumque comprehendissent regem, adduxerunt eum ad regem Babylonis in Rebla, quae est in terra Emath; et locutus est ad eum iudicia.
JER|52|10|Et iugulavit rex Babylonis filios Sedeciae in oculis eius, sed et omnes principes Iudae occidit in Rebla;
JER|52|11|et oculos Sedeciae eruit et vinxit eum compedibus et adduxit eum rex Babylonis in Babylonem et posuit eum in domo carceris usque ad diem mortis eius.
JER|52|12|In mense autem quinto, decima mensis, ipse est annus nonus decimus Nabuchodonosor regis Babylonis, venit Nabuzardan princeps satellitum, qui stabat coram rege Babylonis, in Ierusalem.
JER|52|13|Et incendit domum Domini et domum regis; et omnes domos Ierusalem et omnem domum magnam igni combussit;
JER|52|14|et totum murum Ierusalem per circuitum destruxit cunctus exercitus Chaldaeorum, qui erat cum magistro satellitum.
JER|52|15|De pauperibus autem populi et de reliquo vulgo, quod remanserat in civitate, et de perfugis, qui transfugerant ad regem Babylonis, et superfluos artificum transtulit Nabuzardan princeps satellitum.
JER|52|16|De pauperibus vero terrae reliquit Nabuzardan princeps satellitum in vinitores et in agricolas.
JER|52|17|Columnas quoque aereas, quae erant in domo Domini, et bases et mare aereum, quod erat in domo Domini, confregerunt Chaldaei et tulerunt omne aes eorum in Babylonem.
JER|52|18|Et lebetes et vatilla et cultros et phialas et mortariola et omnia vasa aerea, quae in ministerio fuerant, tulerunt;
JER|52|19|et pelves et thymiamateria et phialas et lebetes et candelabra et mortaria et cyathos, quotquot aurea aurea, et quotquot argentea argentea, tulit magister satellitum;
JER|52|20|columnas duas et mare unum et vitulos duodecim aereos, qui erant subtus basi, quam fecerat rex Salomon domui Domini. Non erat pondus aeris omnium horum vasorum.
JER|52|21|De columnis autem, decem et octo cubiti altitudinis erant in columna una, et funiculus duodecim cubitorum circuibat eam; porro grossitudo eius quattuor digitorum, et intrinsecus cava erat.
JER|52|22|Et capitella super utramque aerea: altitudo capitelli unius quinque cubitorum, et retiacula et malogranata super capitellum in circuitu omnia aerea; similiter columnae secundae.
JER|52|23|Et malogranata nonaginta sex dependentia; omnia malogranata centum super retiacula in circuitu.
JER|52|24|Et tulit magister satellitum Saraiam sacerdotem primum et Sophoniam sacerdotem secundum et tres custodes vestibuli.
JER|52|25|Et de civitate tulit eunuchum unum, qui erat praepositus super viros bellatores, et septem viros de his, qui videbant faciem regis, qui inventi sunt in civitate, et scribam principis militum, qui ex populo terrae probabat tirones, et sexaginta viros de populo terrae, qui inventi sunt in medio civitatis.
JER|52|26|Tulit autem eos Nabuzardan magister satellitum et duxit eos ad regem Babylonis in Rebla;
JER|52|27|et percussit eos rex Babylonis et interfecit eos in Rebla in terra Emath. Et translatus est Iuda de terra sua.
JER|52|28|Iste est populus, quem transtulit Nabuchodonosor: in anno septimo, Iudaeos tria millia et viginti tres;
JER|52|29|in anno octavo decimo Nabuchodonosor de Ierusalem animas octingentas triginta duas;
JER|52|30|in anno vicesimo tertio Nabuchodonosor transtulit Nabuzardan magister satellitum animas Iudaeorum septingentas quadraginta quinque; omnes ergo animae quattuor milia sescentae.
JER|52|31|Et factum est in tricesimo septimo anno transmigrationis Ioachin regis Iudae, duodecimo mense vicesima quinta mensis, elevavit Evilmerodach rex Babylonis, ipso anno regni sui, caput Ioachin regis Iudae; et eduxit eum de domo carceris.
JER|52|32|Et locutus est cum eo bona et posuit thronum eius super thronos regum, qui erant secum in Babylone.
JER|52|33|Et mutavit vestimenta carceris eius, et comedebat panem coram eo semper cunctis diebus vitae suae.
JER|52|34|Et cibaria eius, cibaria perpetua dabantur ei a rege Babylonis statuta per singulos dies, usque ad diem mortis suae, cunctis diebus vitae eius.
