LUKE|1|1|Quoniam quidem multi conati sunt ordinare narrationem, quae in nobis completae sunt, rerum,
LUKE|1|2|sicut tradiderunt nobis, qui ab initio ipsi viderunt et ministri fuerunt verbi,
LUKE|1|3|visum est et mihi, adsecuto a principio omnia, diligenter ex ordine tibi scribere, optime Theophile,
LUKE|1|4|ut cognoscas eorum verborum, de quibus eruditus es, firmitatem.
LUKE|1|5|Fuit in diebus Herodis regis Iudaeae sacerdos quidam nomine Zacharias de vice Abiae, et uxor illi de filiabus Aaron, et nomen eius Elisabeth.
LUKE|1|6|Erant autem iusti ambo ante Deum, incedentes in omnibus mandatis et iustificationibus Domini, irreprehensibiles.
LUKE|1|7|Et non erat illis filius, eo quod esset Elisabeth sterilis, et ambo processissent in diebus suis.
LUKE|1|8|Factum est autem, cum sacerdotio fungeretur in ordine vicis suae ante Deum,
LUKE|1|9|secundum consuetudinem sacerdotii sorte exiit, ut incensum poneret ingressus in templum Domini;
LUKE|1|10|et omnis multitudo erat populi orans foris hora incensi.
LUKE|1|11|Apparuit autem illi angelus Domini stans a dextris altaris incensi;
LUKE|1|12|et Zacharias turbatus est videns, et timor irruit super eum.
LUKE|1|13|Ait autem ad illum angelus: " Ne timeas, Zacharia, quoniam exaudita est deprecatio tua, et uxor tua Elisabeth pariet tibi filium, et vocabis nomen eius Ioannem.
LUKE|1|14|Et erit gaudium tibi et exsultatio, et multi in nativitate eius gaudebunt:
LUKE|1|15|erit enim magnus coram Domino et vinum et siceram non bibet et Spiritu Sancto replebitur adhuc ex utero matris suae
LUKE|1|16|et multos filiorum Israel convertet ad Dominum Deum ipsorum.
LUKE|1|17|Et ipse praecedet ante illum in spiritu et virtute Eliae, ut convertat corda patrum in filios et incredibiles ad prudentiam iustorum, parare Domino plebem perfectam ".
LUKE|1|18|Et dixit Zacharias ad angelum: " Unde hoc sciam? Ego enim sum senex, et uxor mea processit in diebus suis ".
LUKE|1|19|Et respondens angelus dixit ei: " Ego sum Gabriel, qui adsto ante Deum, et missus sum loqui ad te et haec tibi evangelizare.
LUKE|1|20|Et ecce: eris tacens et non poteris loqui usque in diem, quo haec fiant, pro eo quod non credidisti verbis meis, quae implebuntur in tempore suo ".
LUKE|1|21|Et erat plebs exspectans Zachariam, et mirabantur quod tardaret ipse in templo.
LUKE|1|22|Egressus autem non poterat loqui ad illos, et cognoverunt quod visionem vidisset in templo; et ipse erat innuens illis et permansit mutus.
LUKE|1|23|Et factum est, ut impleti sunt dies officii eius, abiit in domum suam.
LUKE|1|24|Post hos autem dies concepit Elisabeth uxor eius et occultabat se mensibus quinque dicens:
LUKE|1|25|" Sic mihi fecit Dominus in diebus, quibus respexit auferre opprobrium meum inter homines ".
LUKE|1|26|In mense autem sexto missus est angelus Gabriel a Deo in civitatem Galilaeae, cui nomen Nazareth,
LUKE|1|27|ad virginem desponsatam viro, cui nomen erat Ioseph de domo David, et nomen virginis Maria.
LUKE|1|28|Et ingressus ad eam dixit: " Ave, gratia plena, Dominus tecum ".
LUKE|1|29|Ipsa autem turbata est in sermone eius et cogitabat qualis esset ista salutatio.
LUKE|1|30|Et ait angelus ei: " Ne timeas, Maria; invenisti enim gratiam apud Deum.
LUKE|1|31|Et ecce concipies in utero et paries filium et vocabis nomen eius Iesum.
LUKE|1|32|Hic erit magnus et Filius Altissimi vocabitur, et dabit illi Dominus Deus sedem David patris eius,
LUKE|1|33|et regnabit super domum Iacob in aeternum, et regni eius non erit finis.
LUKE|1|34|Dixit autem Maria ad angelum: " Quomodo fiet istud, quoniam virum non cognosco? ".
LUKE|1|35|Et respondens angelus dixit ei: " Spiritus Sanctus superveniet in te, et virtus Altissimi obumbrabit tibi: ideoque et quod nascetur sanctum, vocabitur Filius Dei.
LUKE|1|36|Et ecce Elisabeth cognata tua et ipsa concepit filium in senecta sua, et hic mensis est sextus illi, quae vocatur sterilis,
LUKE|1|37|quia non erit impossibile apud Deum omne verbum ".
LUKE|1|38|Dixit autem Maria: " Ecce ancilla Domini; fiat mihi secundum verbum tuum ". Et discessit ab illa angelus.
LUKE|1|39|Exsurgens autem Maria in diebus illis abiit in montana cum festinatione in civitatem Iudae
LUKE|1|40|et intravit in domum Zachariae et salutavit Elisabeth.
LUKE|1|41|Et factum est, ut audivit salutationem Mariae Elisabeth, exsultavit infans in utero eius, et repleta est Spiritu Sancto Elisabeth
LUKE|1|42|et exclamavit voce magna et dixit: " Benedicta tu inter mulieres, et benedictus fructus ventris tui.
LUKE|1|43|Et unde hoc mihi, ut veniat mater Domini mei ad me?
LUKE|1|44|Ecce enim ut facta est vox salutationis tuae in auribus meis, exsultavit in gaudio infans in utero meo.
LUKE|1|45|Et beata, quae credidit, quoniam perficientur ea, quae dicta sunt ei a Domino ".
LUKE|1|46|Et ait Maria: Magnificat anima mea Dominum,
LUKE|1|47|et exsultavit spiritus meus in Deo salvatore meo,
LUKE|1|48|quia respexit humilitatem ancillae suae.Ecce enim ex hoc beatam me dicent omnes generationes,
LUKE|1|49|quia fecit mihi magna, qui potens est,et sanctum nomen eius,
LUKE|1|50|et misericordia eius in progenies et progeniestimentibus eum.
LUKE|1|51|Fecit potentiam in brachio suo,dispersit superbos mente cordis sui;
LUKE|1|52|deposuit potentes de sedeet exaltavit humiles;
LUKE|1|53|esurientes implevit boniset divites dimisit inanes.
LUKE|1|54|Suscepit Israel puerum suum,recordatus misericordiae,
LUKE|1|55|sicut locutus est ad patres nostros,Abraham et semini eius in saecula ".
LUKE|1|56|Mansit autem Maria cum illa quasi mensibus tribus et reversa est in domum suam.
LUKE|1|57|Elisabeth autem impletum est tempus pariendi, et peperit filium.
LUKE|1|58|Et audierunt vicini et cognati eius quia magnificavit Dominus misericordiam suam cum illa, et congratulabantur ei.
LUKE|1|59|Et factum est, in die octavo venerunt circumcidere puerum et vocabant eum nomine patris eius, Zachariam.
LUKE|1|60|Et respondens mater eius dixit: " Nequaquam, sed vocabitur Ioannes ".
LUKE|1|61|Et dixerunt ad illam: " Nemo est in cognatione tua, qui vocetur hoc nomine ".
LUKE|1|62|Innuebant autem patri eius quem vellet vocari eum.
LUKE|1|63|Et postulans pugillarem scripsit dicens: " Ioannes est nomen eius ". Et mirati sunt universi.
LUKE|1|64|Apertum est autem ilico os eius et lingua eius, et loquebatur benedicens Deum.
LUKE|1|65|Et factus est timor super omnes vicinos eorum, et super omnia montana Iudaeae divulgabantur omnia verba haec.
LUKE|1|66|Et posuerunt omnes, qui audierant, in corde suo dicentes: " Quid putas puer iste erit? ". Etenim manus Domini erat cum illo.
LUKE|1|67|Et Zacharias pater eius impletus est Spiritu Sancto et prophetavit dicens:
LUKE|1|68|" Benedictus Dominus, Deus Israel,quia visitavit et fecit redemptionem plebi suae
LUKE|1|69|et erexit cornu salutis nobisin domo David pueri sui,
LUKE|1|70|sicut locutus est per os sanctorum,qui a saeculo sunt, prophetarum eius,
LUKE|1|71|salutem ex inimicis nostriset de manu omnium, qui oderunt nos;
LUKE|1|72|ad faciendam misericordiam cum patribus nostriset memorari testamenti sui sancti,
LUKE|1|73|iusiurandum, quod iuravit ad Abraham patrem nostrum,daturum se nobis,
LUKE|1|74|ut sine timore, de manu inimicorum liberati,serviamus illi
LUKE|1|75|in sanctitate et iustitia coram ipsoomnibus diebus nostris.
LUKE|1|76|Et tu, puer, propheta Altissimi vocaberis:praeibis enim ante faciem Domini parare vias eius,
LUKE|1|77|ad dandam scientiam salutis plebi eiusin remissionem peccatorum eorum,
LUKE|1|78|per viscera misericordiae Dei nostri,in quibus visitabit nos oriens ex alto,
LUKE|1|79|illuminare his, qui in tenebris et in umbra mortis sedent,ad dirigendos pedes nostros in viam pacis ".
LUKE|1|80|Puer autem crescebat et confortabatur spiritu et erat in deserto usque in diem ostensionis suae ad Israel.
LUKE|2|1|Factum est autem, in diebus il lis exiit edictum a Caesare Au gusto, ut describeretur universus orbis.
LUKE|2|2|Haec descriptio prima facta est praeside Syriae Quirino.
LUKE|2|3|Et ibant omnes, ut profiterentur, singuli in suam civitatem.
LUKE|2|4|Ascendit autem et Ioseph a Galilaea de civitate Nazareth in Iudaeam in civitatem David, quae vocatur Bethlehem, eo quod esset de domo et familia David,
LUKE|2|5|ut profiteretur cum Maria desponsata sibi, uxore praegnante.
LUKE|2|6|Factum est autem, cum essent ibi, impleti sunt dies, ut pareret,
LUKE|2|7|et peperit filium suum primogenitum; et pannis eum involvit et reclinavit eum in praesepio, quia non erat eis locus in deversorio.
LUKE|2|8|Et pastores erant in regione eadem vigilantes et custodientes vigilias noctis supra gregem suum.
LUKE|2|9|Et angelus Domini stetit iuxta illos, et claritas Domini circumfulsit illos, et timuerunt timore magno.
LUKE|2|10|Et dixit illis angelus: " Nolite timere; ecce enim evangelizo vobis gaudium magnum, quod erit omni populo,
LUKE|2|11|quia natus est vobis hodie Salvator, qui est Christus Dominus, in civitate David.
LUKE|2|12|Et hoc vobis signum: invenietis infantem pannis involutum et positum in praesepio ".
LUKE|2|13|Et subito facta est cum angelo multitudo militiae caelestis laudantium Deum et dicentium:
LUKE|2|14|" Gloria in altissimis Deo,et super terram pax in hominibus bonae voluntatis ".
LUKE|2|15|Et factum est, ut discesserunt ab eis angeli in caelum, pastores loquebantur ad invicem: " Transeamus usque Bethlehem et videamus hoc verbum, quod factum est, quod Dominus ostendit nobis ".
LUKE|2|16|Et venerunt festinantes et invenerunt Mariam et Ioseph et infantem positum in praesepio.
LUKE|2|17|Videntes autem notum fecerunt verbum, quod dictum erat illis de puero hoc.
LUKE|2|18|Et omnes, qui audierunt, mirati sunt de his, quae dicta erant a pastoribus ad ipsos.
LUKE|2|19|Maria autem conservabat omnia verba haec conferens in corde suo.
LUKE|2|20|Et reversi sunt pastores glorificantes et laudantes Deum in omnibus, quae audierant et viderant, sicut dictum est ad illos.
LUKE|2|21|Et postquam consummati sunt dies octo, ut circumcideretur, vocatum est nomen eius Iesus, quod vocatum est ab angelo, priusquam in utero conciperetur.
LUKE|2|22|Et postquam impleti sunt dies purgationis eorum secundum legem Moysis, tulerunt illum in Hierosolymam, ut sisterent Domino,
LUKE|2|23|sicut scriptum est in lege Domini: " Omne masculinum adaperiens vulvam sanctum Domino vocabitur ",
LUKE|2|24|et ut darent hostiam secundum quod dictum est in lege Domini: par turturum aut duos pullos columbarum.
LUKE|2|25|Et ecce homo erat in Ierusalem, cui nomen Simeon, et homo iste iustus et timoratus, exspectans consolationem Israel, et Spiritus Sanctus erat super eum;
LUKE|2|26|et responsum acceperat ab Spiritu Sancto non visurum se mortem nisi prius videret Christum Domini.
LUKE|2|27|Et venit in Spiritu in templum. Et cum inducerent puerum Iesum parentes eius, ut facerent secundum consuetudinem legis pro eo,
LUKE|2|28|et ipse accepit eum in ulnas suas et benedixit Deum et dixit:
LUKE|2|29|" Nunc dimittis servum tuum, Domine,secundum verbum tuum in pace,
LUKE|2|30|quia viderunt oculi meisalutare tuum,
LUKE|2|31|quod parastiante faciem omnium populorum,
LUKE|2|32|lumen ad revelationem gentiumet gloriam plebis tuae Israel ".
LUKE|2|33|Et erat pater eius et mater mirantes super his, quae dicebantur de illo.
LUKE|2|34|Et benedixit illis Simeon et dixit ad Mariam matrem eius: " Ecce positus est hic in ruinam et resurrectionem multorum in Israel et in signum, cui contradicetur
LUKE|2|35|- et tuam ipsius animam pertransiet gladius - ut revelentur ex multis cordibus cogitationes ".
LUKE|2|36|Et erat Anna prophetissa, filia Phanuel, de tribu Aser. Haec processerat in diebus multis et vixerat cum viro annis septem a virginitate sua;
LUKE|2|37|et haec vidua usque ad annos octoginta quattuor, quae non discedebat de templo, ieiuniis et obsecrationibus serviens nocte ac die.
LUKE|2|38|Et haec ipsa hora superveniens confitebatur Deo et loquebatur de illo omnibus, qui exspectabant redemptionem Ierusalem.
LUKE|2|39|Et ut perfecerunt omnia secundum legem Domini, reversi sunt in Galilaeam in civitatem suam Nazareth.
LUKE|2|40|Puer autem crescebat et confortabatur plenus sapientia; et gratia Dei erat super illum.
LUKE|2|41|Et ibant parentes eius per omnes annos in Ierusalem in die festo Paschae.
LUKE|2|42|Et cum factus esset annorum duodecim, ascendentibus illis secundum consuetudinem diei festi,
LUKE|2|43|consummatisque diebus, cum redirent, remansit puer Iesus in Ierusalem, et non cognoverunt parentes eius.
LUKE|2|44|Existimantes autem illum esse in comitatu, venerunt iter diei et requirebant eum inter cognatos et notos;
LUKE|2|45|et non invenientes regressi sunt in Ierusalem requirentes eum.
LUKE|2|46|Et factum est, post triduum invenerunt illum in templo sedentem in medio doctorum, audientem illos et interrogantem eos;
LUKE|2|47|stupebant autem omnes, qui eum audiebant, super prudentia et responsis eius.
LUKE|2|48|Et videntes eum admirati sunt, et dixit Mater cius ad illum: " Fili, quid fecisti nobis sic? Ecce pater tuus et ego dolentes quaerebamus te ".
LUKE|2|49|Et ait ad illos: " Quid est quod me quaerebatis? Nesciebatis quia in his, quae Patris mei sunt, oportet me esse? ".
LUKE|2|50|Et ipsi non intellexerunt verbum, quod locutus est ad illos.
LUKE|2|51|Et descendit cum eis et venit Nazareth et erat subditus illis. Et mater eius conservabat omnia verba in corde suo.
LUKE|2|52|Et Iesus proficiebat sapientia et aetate et gratia apud Deum et homines.
LUKE|3|1|Anno autem quinto decimo im perii Tiberii Caesaris, procu rante Pontio Pilato Iudaeam, tetrarcha autem Galilaeae Herode, Philippo autem fratre eius tetrarcha Ituraeae et Trachonitidis regionis, et Lysania Abilinae tetrarcha,
LUKE|3|2|sub principe sacerdotum Anna et Caipha, factum est verbum Dei super Ioannem Zachariae filium in deserto.
LUKE|3|3|Et venit in omnem regionem circa Iordanem praedicans baptismum paenitentiae in remissionem peccatorum,
LUKE|3|4|sicut scriptum est in libro sermonum Isaiae prophetae: Vox clamantis in deserto:Parate viam Domini,rectas facite semitas eius.
LUKE|3|5|Omnis vallis implebitur,et omnis mons et collis humiliabitur;et erunt prava in directa,et aspera in vias planas:
LUKE|3|6|et videbit omnis caro salutare Dei" ".
LUKE|3|7|Dicebat ergo ad turbas, quae exibant, ut baptizarentur ab ipso: " Genimina viperarum, quis ostendit vobis fugere a ventura ira?
LUKE|3|8|Facite ergo fructus dignos paenitentiae et ne coeperitis dicere in vobis ipsis: "Patrem habemus Abraham"; dico enim vobis quia potest Deus de lapidibus istis suscitare Abrahae filios.
LUKE|3|9|Iam enim et securis ad radicem arborum posita est; omnis ergo arbor non faciens fructum bonum exciditur et in ignem mittitur ".
LUKE|3|10|Et interrogabant eum turbae dicentes: " Quid ergo faciemus? ".
LUKE|3|11|Respondens autem dicebat illis: " Qui habet duas tunicas, det non habenti; et, qui habet escas, similiter faciat ".
LUKE|3|12|Venerunt autem et publicani, ut baptizarentur, et dixerunt ad illum: " Magister, quid faciemus? ".
LUKE|3|13|At ille dixit ad eos: " Nihil amplius quam constitutum est vobis, faciatis ".
LUKE|3|14|Interrogabant autem eum et milites dicentes: " Quid faciemus et nos? ". Et ait illis: " Neminem concutiatis neque calumniam faciatis et contenti estote stipendiis vestris ".
LUKE|3|15|Existimante autem populo et cogitantibus omnibus in cordibus suis de Ioanne, ne forte ipse esset Christus,
LUKE|3|16|respondit Ioannes dicens omnibus: " Ego quidem aqua baptizo vos. Venit autem fortior me, cuius non sum dignus solvere corrigiam calceamentorum eius: ipse vos baptizabit in Spiritu Sancto et igni;
LUKE|3|17|cuius ventilabrum in manu eius ad purgandam aream suam et ad congregandum triticum in horreum suum, paleas autem comburet igni inexstinguibili ".
LUKE|3|18|Multa quidem et alia exhortans evangelizabat populum.
LUKE|3|19|Herodes autem tetrarcha, cum corriperetur ab illo de Herodiade uxore fratris sui et de omnibus malis, quae fecit Herodes,
LUKE|3|20|adiecit et hoc supra omnia et inclusit Ioannem in carcere.
LUKE|3|21|Factum est autem, cum baptizaretur omnis populus, et Iesu baptizato et orante, apertum est caelum,
LUKE|3|22|et descendit Spiritus Sanctus corporali specie sicut columba super ipsum; et vox de caelo facta est: " Tu es Filius meus dilectus; in te complacui mihi ".
LUKE|3|23|Et ipse Iesus erat incipiens quasi annorum triginta, ut putabatur, filius Ioseph, qui fuit Heli,
LUKE|3|24|qui fuit Matthat, qui fuit Levi, qui fuit Melchi, qui fuit Iannae, qui fuit Ioseph,
LUKE|3|25|qui fuit Matthathiae, qui fuit Amos, qui fuit Nahum, qui fuit Esli, qui fuit Naggae,
LUKE|3|26|qui fuit Maath, qui fuit Matthathiae, qui fuit Semei, qui fuit Iosech, qui fuit Ioda,
LUKE|3|27|qui fuit Ioanna, qui fuit Resa, qui fuit Zorobabel, qui fuit Salathiel, qui fuit Neri,
LUKE|3|28|qui fuit Melchi, qui fuit Addi, qui fuit Cosam, qui fuit Elmadam, qui fuit Her,
LUKE|3|29|qui fuit Iesu, qui fuit Eliezer, qui fuit Iorim, qui fuit Matthat, qui fuit Levi,
LUKE|3|30|qui fuit Simeon, qui fuit Iudae, qui fuit Ioseph, qui fuit Iona, qui fuit Eliachim,
LUKE|3|31|qui fuit Melea, qui fuit Menna, qui fuit Matthatha, qui fuit Nathan, qui fuit David,
LUKE|3|32|qui fuit Iesse, qui fuit Obed, qui fuit Booz, qui fuit Salmon, qui fuit Naasson,
LUKE|3|33|qui fuit Aminadab, qui fuit Admin, qui fuit Arni, qui fuit Esrom, qui fuit Phares, qui fuit Iudae,
LUKE|3|34|qui fuit Iacob, qui fuit Isaac, qui fuit Abrahae, qui fuit Thare, qui fuit Nachor,
LUKE|3|35|qui fuit Seruch, qui fuit Ragau, qui fuit Phaleg, qui fuit Heber, qui fuit Sala,
LUKE|3|36|qui fuit Cainan, qui fuit Arphaxad, qui fuit Sem, qui fuit Noe, qui fuit Lamech,
LUKE|3|37|qui fuit Mathusala, qui fuit Henoch, qui fuit Iared, qui fuit Malaleel, qui fuit Cainan,
LUKE|3|38|qui fuit Enos, qui fuit Seth, qui fuit Adam, qui fuit Dei.
LUKE|4|1|Iesus autem plenus Spiritu Sancto regressus est ab Iordane et agebatur in Spiritu in deserto
LUKE|4|2|diebus quadraginta et tentabatur a Diabolo. Et nihil manducavit in diebus illis et, consummatis illis, esuriit.
LUKE|4|3|Dixit autem illi Diabolus: " Si Filius Dei es, dic lapidi huic, ut panis fiat ".
LUKE|4|4|Et respondit ad illum Iesus: " Scriptum est: "Non in pane solo vivet homo" ".
LUKE|4|5|Et sustulit illum et ostendit illi omnia regna orbis terrae in momento temporis;
LUKE|4|6|et ait ei Diabolus: " Tibi dabo potestatem hanc universam et gloriam illorum, quia mihi tradita est, et, cui volo, do illam:
LUKE|4|7|tu ergo, si adoraveris coram me, erit tua omnis ".
LUKE|4|8|Et respondens Iesus dixit illi: " Scriptum est: "Dominum Deum tuum adorabis et illi soli servies" ".
LUKE|4|9|Duxit autem illum in Ierusalem et statuit eum supra pinnam templi et dixit illi: " Si Filius Dei es, mitte te hinc deorsum.
LUKE|4|10|Scriptum est enim:Angelis suis mandabit de te,ut conservent te"
LUKE|4|11|et: "In manibus tollent te,ne forte offendas ad lapidem pedem tuum" ".
LUKE|4|12|Et respondens Iesus ait illi: " Dictum est: "Non tentabis Dominum Deum tuum" ".
LUKE|4|13|Et consummata omni tentatione, Diabolus recessit ab illo usque ad tempus.
LUKE|4|14|Et regressus est Iesus in virtute Spiritus in Galilaeam. Et fama exiit per universam regionem de illo.
LUKE|4|15|Et ipse docebat in synagogis eorum et magnificabatur ab omnibus.
LUKE|4|16|Et venit Nazareth, ubi erat nutritus, et intravit secundum consuetudinem suam die sabbati in synagogam et surrexit legere.
LUKE|4|17|Et tradi tus est illi liber prophetae Isaiae; etut revolvit librum, invenit locum, ubi scriptum erat:
LUKE|4|18|" Spiritus Domini super me;propter quod unxit meevangelizare pauperibus,misit me praedicare captivis remissionemet caecis visum,dimittere confractos in remissione,
LUKE|4|19|praedicare annum Domini acceptum ".
LUKE|4|20|Et cum plicuisset librum, reddidit ministro et sedit; et omnium in synagoga oculi erant intendentes in eum.
LUKE|4|21|Coepit autem dicere ad illos: " Hodie impleta est haec Scriptura in auribus vestris ".
LUKE|4|22|Et omnes testimonium illi dabant et mirabantur in verbis gratiae, quae procedebant de ore ipsius, et dicebant: " Nonne hic filius est Ioseph? ".
LUKE|4|23|Et ait illis: " Utique dicetis mihi hanc similitudinem: "Medice, cura teipsum; quanta audivimus facta in Capharnaum, fac et hic in patria tua".
LUKE|4|24|Ait autem: " Amen dico vobis: Nemo propheta acceptus est in patria sua.
LUKE|4|25|In veritate autem dico vobis: Multae viduae erant in diebus Eliae in Israel, quando clausum est caelum annis tribus et mensibus sex, cum facta est fames magna in omni terra;
LUKE|4|26|et ad nullam illarum missus est Elias nisi in Sarepta Sidoniae ad mulierem viduam.
LUKE|4|27|Et multi leprosi erant in Israel sub Eliseo propheta; et nemo eorum mundatus est nisi Naaman Syrus ".
LUKE|4|28|Et repleti sunt omnes in synagoga ira haec audientes;
LUKE|4|29|et surrexerunt et eiecerunt illum extra civitatem et duxerunt illum usque ad supercilium montis, supra quem civitas illorum erat aedificata, ut praecipitarent eum.
LUKE|4|30|Ipse autem transiens per medium illorum ibat.
LUKE|4|31|Et descendit in Capharnaum civitatem Galilaeae. Et docebat illos sabbatis;
LUKE|4|32|et stupebant in doctrina eius, quia in potestate erat sermo ipsius.
LUKE|4|33|Et in synagoga erat homo habens spiritum daemonii immundi; et exclamavit voce magna:
LUKE|4|34|" Sine; quid nobis et tibi, Iesu Nazarene? Venisti perdere nos? Scio te qui sis: Sanctus Dei ".
LUKE|4|35|Et increpavit illi Iesus dicens: " Obmutesce et exi ab illo! ". Et cum proiecisset illum daemonium in medium, exiit ab illo nihilque illum nocuit.
LUKE|4|36|Et factus est pavor in omnibus; et colloquebantur ad invicem dicentes: Quod est hoc verbum, quia in potestate et virtute imperat immundis spiritibus, et exeunt? ".
LUKE|4|37|Et divulgabatur fama de illo in omnem locum regionis.
LUKE|4|38|Surgens autem de synagoga introivit in domum Simonis. Socrus autem Simonis tenebatur magna febri; et rogaverunt illum pro ea.
LUKE|4|39|Et stans super illam imperavit febri, et dimisit illam; et continuo surgens ministrabat illis.
LUKE|4|40|Cum sol autem occidisset, omnes, qui habebant infirmos variis languoribus, ducebant illos ad eum; at ille singulis manus imponens curabat eos.
LUKE|4|41|Exibant autem daemonia a multis clamantia et dicentia: " Tu es Filius Dei ". Et increpans non sinebat ea loqui, quia sciebant ipsum esse Christum.
LUKE|4|42|Facta autem die, egressus ibat in desertum locum; et turbae requirebant eum et venerunt usque ad ipsum et detinebant illum, ne discederet ab eis.
LUKE|4|43|Quibus ille ait: " Et aliis civitatibus oportet me evangelizare regnum Dei, quia ideo missus sum ".
LUKE|4|44|Et erat praedicans in synagogis Iudaeae.
LUKE|5|1|Factum est autem, cum turba urgeret illum et audiret verbum Dei, et ipse stabat secus stagnum Genesareth
LUKE|5|2|et vidit duas naves stantes secus stagnum; piscatores autem descenderant de illis et lavabant retia.
LUKE|5|3|Ascendens autem in unam navem, quae erat Simonis, rogavit eum a terra reducere pusillum; et sedens docebat de navicula turbas.
LUKE|5|4|Ut cessavit autem loqui, dixit ad Simonem: " Duc in altum et laxate retia vestra in capturam ".
LUKE|5|5|Et respondens Simon dixit: " Praeceptor, per totam noctem laborantes nihil cepimus; in verbo autem tuo laxabo retia ".
LUKE|5|6|Et cum hoc fecissent, concluserunt piscium multitudinem copiosam; rumpebantur autem retia eorum.
LUKE|5|7|Et annuerunt sociis, qui erant in alia navi, ut venirent et adiuvarent eos; et venerunt et impleverunt ambas naviculas, ita ut mergerentur.
LUKE|5|8|Quod cum videret Simon Petrus, procidit ad genua Iesu dicens: " Exi a me, quia homo peccator sum, Domine ".
LUKE|5|9|Stupor enim circumdederat eum et omnes, qui cum illo erant, in captura piscium, quos ceperant;
LUKE|5|10|similiter autem et Iacobum et Ioannem, filios Zebedaei, qui erant socii Simonis. Et ait ad Simonem Iesus: " Noli timere; ex hoc iam homines eris capiens ".
LUKE|5|11|Et subductis ad terram navibus, relictis omnibus, secuti sunt illum.
LUKE|5|12|Et factum est, cum esset in una civitatum, et ecce vir plenus lepra; et videns Iesum et procidens in faciem rogavit eum dicens: " Domine, si vis, potes me mundare ".
LUKE|5|13|Et extendens manum tetigit illum dicens: " Volo, mundare! "; et confestim lepra discessit ab illo.
LUKE|5|14|Et ipse praecepit illi, ut nemini diceret, sed: " Vade, ostende te sacerdoti et offer pro emundatione tua, sicut praecepit Moyses, in testimonium illis ".
LUKE|5|15|Perambulabat autem magis sermo de illo, et conveniebant turbae multae, ut audirent et curarentur ab infirmitatibus suis;
LUKE|5|16|ipse autem secedebat in desertis et orabat.
LUKE|5|17|Et factum est, in una dierum, et ipse erat docens, et erant pharisaei sedentes et legis doctores, qui venerant ex omni castello Galilaeae et Iudaeae et Ierusalem; et virtus Domini erat ei ad sanandum.
LUKE|5|18|Et ecce viri portantes in lecto hominem, qui erat paralyticus, et quaerebant eum inferre et ponere ante eum.
LUKE|5|19|Et non invenientes qua parte illum inferrent prae turba, ascenderunt supra tectum et per tegulas summiserunt illum cum lectulo in medium ante Iesum.
LUKE|5|20|Quorum fidem ut vidit, dixit: " Homo, remittuntur tibi peccata tua ".
LUKE|5|21|Et coeperunt cogitare scribae et pharisaei dicentes: " Quis est hic, qui loquitur blasphemias? Quis potest dimittere peccata nisi solus Deus?.
LUKE|5|22|Ut cognovit autem Iesus cogitationes eorum, respondens dixit ad illos: Quid cogitatis in cordibus vestris?
LUKE|5|23|Quid est facilius, dicere: "Dimittuntur tibi peccata tua", an dicere: Surge et ambula"?
LUKE|5|24|Ut autem sciatis quia Filius hominis potestatem habet in terra dimittere peccata - ait paralytico -: Tibi dico: Surge, tolle lectulum tuum et vade in domum tuam ".
LUKE|5|25|Et confestim surgens coram illis tulit, in quo iacebat, et abiit in domum suam magnificans Deum.
LUKE|5|26|Et stupor apprehendit omnes, et magnificabant Deum; et repleti sunt timore dicentes: " Vidimus mirabilia hodie ".
LUKE|5|27|Et post haec exiit et vidit publicanum nomine Levi sedentem ad teloneum et ait illi: " Sequere me ".
LUKE|5|28|Et relictis omnibus, surgens secutus est eum.
LUKE|5|29|Et fecit ei convivium magnum Levi in domo sua; et erat turba multa publicanorum et aliorum, qui cum illis erant discumbentes.
LUKE|5|30|Et murmurabant pharisaei et scribae eorum adversus discipulos eius dicentes: " Quare cum publicanis et peccatoribus manducatis et bibitis? ".
LUKE|5|31|Et respondens Iesus dixit ad illos: " Non egent, qui sani sunt, medico, sed qui male habent.
LUKE|5|32|Non veni vocare iustos sed peccatores in paenitentiam ".
LUKE|5|33|At illi dixerunt ad eum: " Discipuli Ioannis ieiunant frequenter et obsecrationes faciunt, similiter et pharisaeorum; tui autem edunt et bibunt ".
LUKE|5|34|Quibus Iesus ait: " Numquid potestis convivas nuptiarum, dum cum illis est sponsus, facere ieiunare?
LUKE|5|35|Venient autem dies; et cum ablatus fuerit ab illis sponsus, tunc ieiunabunt in illis diebus ".
LUKE|5|36|Dicebat autem et similitudinem ad illos: " Nemo abscindit commissuram a vestimento novo et immittit in vestimentum vetus; alioquin et novum rumpet, et veteri non conveniet commissura a novo.
LUKE|5|37|Et nemo mittit vinum novum in utres veteres; alioquin rumpet vinum novum utres et ipsum effundetur, et utres peribunt;
LUKE|5|38|sed vinum novum in utres novos mittendum est.
LUKE|5|39|Et nemo bibens vetus vult novum; dicit enim: "Vetus melius est!" ".
LUKE|6|1|Factum est autem in sabbato, cum transiret per sata, et velle bant discipuli eius spicas et manducabant confricantes manibus.
LUKE|6|2|Quidam autem pharisaeorum dixerunt: " Quid facitis, quod non licet in sabbatis? ".
LUKE|6|3|Et respondens Iesus ad eos dixit: " Nec hoc legistis, quod fecit David, cum esurisset ipse et qui cum eo erant?
LUKE|6|4|Quomodo intravit in domum Dei et panes propositionis sumpsit et manducavit et dedit his, qui cum ipso erant, quos non licet manducare nisi tantum sacerdotibus? ".
LUKE|6|5|Et dicebat illis: " Dominus est sabbati Filius hominis ".
LUKE|6|6|Factum est autem in alio sabbato, ut intraret in synagogam et doceret; et erat ibi homo, et manus eius dextra erat arida.
LUKE|6|7|Observabant autem illum scribae et pharisaei, si sabbato curaret, ut invenirent accusare illum.
LUKE|6|8|Ipse vero sciebat cogitationes eorum et ait homini, qui habebat manum aridam: " Surge et sta in medium ". Et surgens stetit.
LUKE|6|9|Ait autem ad illos Iesus: " Interrogo vos, si licet sabbato bene facere an male; animam salvam facere an perdere? ".
LUKE|6|10|Et circumspectis omnibus illis, dixit illi: " Extende manum tuam ". Et fecit; et restituta est manus eius.
LUKE|6|11|Ipsi autem repleti sunt insipientia et colloquebantur ad invicem quidnam facerent Iesu.
LUKE|6|12|Factum est autem in illis diebus, exiit in montem orare et erat pernoctans in oratione Dei.
LUKE|6|13|Et cum dies factus esset, vocavit discipulos suos et elegit Duodecim ex ipsis, quos et apostolos nominavit:
LUKE|6|14|Simonem, quem et cognominavit Petrum, et Andream fratrem eius et Iacobum et Ioannem et Philippum et Bartholomaeum
LUKE|6|15|et Matthaeum et Thomam et Iacobum Alphaei et Simonem, qui vocatur Zelotes,
LUKE|6|16|et Iudam Iacobi et Iudam Iscarioth, qui fuit proditor.
LUKE|6|17|Et descendens cum illis stetit in loco campestri, et turba multa discipulorum eius, et multitudo copiosa plebis ab omni Iudaea et Ierusalem et maritima Tyri et Sidonis,
LUKE|6|18|qui venerunt, ut audirent eum et sanarentur a languoribus suis; et, qui vexabantur a spiritibus immundis, curabantur.
LUKE|6|19|Et omnis turba quaerebant eum tangere, quia virtus de illo exibat et sanabat omnes.
LUKE|6|20|Et ipse, elevatis oculis suis in discipulos suos, dicebat: Beati pauperes, quia vestrum est regnum Dei.
LUKE|6|21|Beati, qui nunc esuritis, quia saturabimini.Beati, qui nunc fletis, quia ridebitis.
LUKE|6|22|Beati eritis, cum vos oderint homines et cum separaverint vos et exprobraverint et eiecerint nomen vestrum tamquam malum propter Filium hominis.
LUKE|6|23|Gaudete in illa die et exsultate, ecce enim merces vestra multa in caelo; secundum haec enim faciebant prophetis patres eorum.
LUKE|6|24|Verumtamen vae vobis divitibus, quia habetis consolationem vestram!
LUKE|6|25|Vae vobis, qui saturati estis nunc, quia esurietis!Vae vobis, qui ridetis nunc, quia lugebitis et flebitis!
LUKE|6|26|Vae, cum bene vobis dixerint omnes homines! Secundum haec enim faciebant pseudoprophetis patres eorum.
LUKE|6|27|Sed vobis dico, qui auditis: Diligite inimicos vestros, bene facite his, qui vos oderunt;
LUKE|6|28|benedicite male dicentibus vobis, orate pro calumniantibus vos.
LUKE|6|29|Ei, qui te percutit in maxillam, praebe et alteram; et ab eo, qui aufert tibi vestimentum, etiam tunicam noli prohibere.
LUKE|6|30|Omni petenti te tribue; et ab eo, qui aufert, quae tua sunt, ne repetas.
LUKE|6|31|Et prout vultis, ut faciant vobis homines, facite illis similiter.
LUKE|6|32|Et si diligitis eos, qui vos diligunt, quae vobis est gratia? Nam et peccatores diligentes se diligunt.
LUKE|6|33|Et si bene feceritis his, qui vobis bene faciunt, quae vobis est gratia? Si quidem et peccatores idem faciunt.
LUKE|6|34|Et si mutuum dederitis his, a quibus speratis recipere, quae vobis gratia est? Nam et peccatores peccatoribus fenerantur, ut recipiant aequalia.
LUKE|6|35|Verumtamen diligite inimicos vestros et bene facite et mutuum date nihil desperantes; et erit merces vestra multa, et eritis filii Altissimi, quia ipse benignus est super ingratos et malos.
LUKE|6|36|Estote misericordes, sicut et Pater vester misericors est.
LUKE|6|37|Et nolite iudicare et non iudicabimini; et nolite condemnare et non condemnabimini. Dimittite et dimittemini;
LUKE|6|38|date, et dabitur vobis: mensuram bonam, confertam, coagitatam, supereffluentem dabunt in sinum vestrum; eadem quippe mensura, qua mensi fueritis, remetietur vobis ".
LUKE|6|39|Dixit autem illis et similitudinem: " Numquid potest caecus caecum ducere? Nonne ambo in foveam cadent?
LUKE|6|40|Non est discipulus super magistrum; perfectus autem omnis erit sicut magister eius.
LUKE|6|41|Quid autem vides festucam in oculo fratris tui, trabem autem, quae in oculo tuo est, non consideras?
LUKE|6|42|Quomodo potes dicere fratri tuo: "Frater, sine eiciam festucam, quae est in oculo tuo", ipse in oculo tuo trabem non videns? Hypocrita, eice primum trabem de oculo tuo et tunc perspicies, ut educas festucam, quae est in oculo fratris tui.
LUKE|6|43|Non est enim arbor bona faciens fructum malum, neque iterum arbor mala faciens fructum bonum.
LUKE|6|44|Unaquaeque enim arbor de fructu suo cognoscitur; neque enim de spinis colligunt ficus, neque de rubo vindemiant uvam.
LUKE|6|45|Bonus homo de bono thesauro cordis profert bonum, et malus homo de malo profert malum: ex abundantia enim cordis os eius loquitur.
LUKE|6|46|Quid autem vocatis me: "Domine, Domine", et non facitis, quae dico?
LUKE|6|47|Omnis, qui venit ad me et audit sermones meos et facit eos, ostendam vobis cui similis sit:
LUKE|6|48|similis est homini aedificanti domum, qui fodit in altum et posuit fundamentum supra petram; inundatione autem facta, illisum est flumen domui illi et non potuit eam movere; bene enim aedificata erat.
LUKE|6|49|Qui autem audivit et non fecit, similis est homini aedificanti domum suam supra terram sine fundamento; in quam illisus est fluvius, et continuo cecidit, et facta est ruina domus illius magna ".
LUKE|7|1|Cum autem implesset omnia verba sua in aures plebis, intra vit Capharnaum.
LUKE|7|2|Centurionis autem cuiusdam servus male habens erat moriturus, qui illi erat pretiosus.
LUKE|7|3|Et cum audisset de Iesu, misit ad eum seniores Iudaeorum rogans eum, ut veniret et salvaret servum eius.
LUKE|7|4|At illi cum venissent ad Iesum, rogabant eum sollicite dicentes: " Dignus est, ut hoc illi praestes:
LUKE|7|5|diligit enim gentem nostram et synagogam ipse aedificavit nobis ".
LUKE|7|6|Iesus autem ibat cum illis. At cum iam non longe esset a domo, misit centurio amicos dicens ei: " Domine, noli vexari; non enim dignus sum, ut sub tectum meum intres,
LUKE|7|7|propter quod et meipsum non sum dignum arbitratus, ut venirem ad te; sed dic verbo, et sanetur puer meus.
LUKE|7|8|Nam et ego homo sum sub potestate constitutus, habens sub me milites, et dico huic: "Vade", et vadit; et alii: "Veni", et venit; et servo meo: "Fac hoc", et facit ".
LUKE|7|9|Quo audito, Iesus miratus est eum et conversus sequentibus se turbis dixit: " Dico vobis, nec in Israel tantam fidem inveni! ".
LUKE|7|10|Et reversi, qui missi fuerant, domum, invenerunt servum sanum.
LUKE|7|11|Et factum est, deinceps ivit in civitatem, quae vocatur Naim, et ibant cum illo discipuli eius et turba copiosa.
LUKE|7|12|Cum autem appropinquaret portae civitatis, et ecce defunctus efferebatur filius unicus matri suae; et haec vidua erat, et turba civitatis multa cum illa.
LUKE|7|13|Quam cum vidisset Dominus, misericordia motus super ea dixit illi: " Noli flere! ".
LUKE|7|14|Et accessit et tetigit loculum; hi autem, qui portabant, steterunt. Et ait: " Adulescens, tibi dico: Surge! ".
LUKE|7|15|Et resedit, qui erat mortuus, et coepit loqui; et dedit illum matri suae.
LUKE|7|16|Accepit autem omnes timor, et magnificabant Deum dicentes: " Propheta magnus surrexit in nobis " et: " Deus visitavit plebem suam ".
LUKE|7|17|Et exiit hic sermo in universam Iudaeam de eo et omnem circa regionem.
LUKE|7|18|Et nuntiaverunt Ioanni discipuli eius de omnibus his.
LUKE|7|19|Et convocavit duos de discipulis suis Ioannes et misit ad Dominum dicens: " Tu es qui venturus es, an alium exspectamus? ".
LUKE|7|20|Cum autem venissent ad eum viri, dixerunt: " Ioannes Baptista misit nos ad te dicens: "Tu es qui venturus es, an alium exspectamus?" ".
LUKE|7|21|In ipsa hora curavit multos a languoribus et plagis et spiritibus malis et caecis multis donavit visum.
LUKE|7|22|Et respondens dixit illis: " Euntes nuntiate Ioanni, quae vidistis et audistis: caeci vident, claudi ambulant, leprosi mundantur et surdi audiunt, mortui resurgunt, pauperes evangelizantur;
LUKE|7|23|et beatus est, quicumque non fuerit scandalizatus in me ".
LUKE|7|24|Et cum discessissent nuntii Ioannis, coepit dicere de Ioanne ad turbas: Quid existis in desertum videre? Arundinem vento moveri?
LUKE|7|25|Sed quid existis videre? Hominem mollibus vestimentis indutum? Ecce, qui in veste pretiosa sunt et deliciis, in domibus regum sunt.
LUKE|7|26|Sed quid existis videre? Prophetam? Utique, dico vobis, et plus quam prophetam.
LUKE|7|27|Hic est, de quo scriptum est:Ecce mitto angelum meum ante faciem tuam,qui praeparabit viam tuam ante te".
LUKE|7|28|Dico vobis: Maior inter natos mulierum Ioanne nemo est; qui autem minor est in regno Dei, maior est illo.
LUKE|7|29|Et omnis populus audiens et publicani iustificaverunt Deum, baptizati baptismo Ioannis;
LUKE|7|30|pharisaei autem et legis periti consilium Dei spreverunt in semetipsos, non baptizati ab eo.
LUKE|7|31|Cui ergo similes dicam homines generationis huius, et cui similes sunt?
LUKE|7|32|Similes sunt pueris sedentibus in foro et loquentibus ad invicem, quod dicit:Cantavimus vobis tibiis, et non saltastis;lamentavimus, et non plorastis!".
LUKE|7|33|Venit enim Ioannes Baptista neque manducans panem neque bibens vinum, et dicitis: "Daemonium habet!";
LUKE|7|34|venit Filius hominis manducans et bibens, et dicitis: "Ecce homo devorator et bibens vinum, amicus publicanorum et peccatorum!".
LUKE|7|35|Et iustificata est sapientia ab omnibus filiis suis ".
LUKE|7|36|Rogabat autem illum quidam de pharisaeis, ut manducaret cum illo; et ingressus domum pharisaei discubuit.
LUKE|7|37|Et ecce mulier, quae erat in civitate peccatrix, ut cognovit quod accubuit in domo pharisaei, attulit alabastrum unguenti;
LUKE|7|38|et stans retro secus pedes eius flens lacrimis coepit rigare pedes eius et capillis capitis sui tergebat, et osculabatur pedes eius et unguento ungebat.
LUKE|7|39|Videns autem pharisaeus, qui vocaverat eum, ait intra se dicens: " Hic si esset propheta, sciret utique quae et qualis mulier, quae tangit eum, quia peccatrix est ".
LUKE|7|40|Et respondens Iesus dixit ad illum: " Simon, habeo tibi aliquid dicere. At ille ait: " Magister, dic ".
LUKE|7|41|" Duo debitores erant cuidam feneratori: unus debebat denarios quingentos, alius quinquaginta.
LUKE|7|42|Non habentibus illis, unde redderent, donavit utrisque. Quis ergo eorum plus diliget eum? ".
LUKE|7|43|Respondens Simon dixit: " Aestimo quia is, cui plus donavit ". At ille dixit ei: " Recte iudicasti ".
LUKE|7|44|Et conversus ad mulierem, dixit Simoni: " Vides hanc mulierem? Intravi in domum tuam: aquam pedibus meis non dedisti; haec autem lacrimis rigavit pedes meos et capillis suis tersit.
LUKE|7|45|Osculum mihi non dedisti; haec autem, ex quo intravi, non cessavit osculari pedes meos.
LUKE|7|46|Oleo caput meum non unxisti; haec autem unguento unxit pedes meos.
LUKE|7|47|Propter quod dico tibi: Remissa sunt peccata eius multa, quoniam dilexit multum; cui autem minus dimittitur, minus diligit ".
LUKE|7|48|Dixit autem ad illam: " Remissa sunt peccata tua ".
LUKE|7|49|Et coeperunt, qui simul accumbebant, dicere intra se: " Quis est hic, qui etiam peccata dimittit?".
LUKE|7|50|Dixit autem ad mulierem: " Fides tua te salvam fecit; vade in pace! ".
LUKE|8|1|Et factum est deinceps, et ipse iter faciebat per civitatem et ca stellum praedicans et evangelizans regnum Dei; et Duodecim cum illo
LUKE|8|2|et mulieres aliquae, quae erant curatae ab spiritibus malignis et infirmitatibus: Maria, quae vocatur Magdalene, de qua daemonia septem exierant,
LUKE|8|3|et Ioanna uxor Chuza, procuratoris Herodis, et Susanna et aliae multae, quae ministrabant eis de facultatibus suis.
LUKE|8|4|Cum autem turba plurima conveniret, et de singulis civitatibus properarent ad eum, dixit per similitudinem:
LUKE|8|5|" Exiit, qui seminat, seminare semen suum. Et dum seminat ipse, aliud cecidit secus viam et conculcatum est, et volucres caeli comederunt illud.
LUKE|8|6|Et aliud cecidit super petram et natum aruit, quia non habebat umorem.
LUKE|8|7|Et aliud cecidit inter spinas, et simul exortae spinae suffocaverunt illud.
LUKE|8|8|Et aliud cecidit in terram bonam et ortum fecit fructum centuplum ". Haec dicens clamabat: " Qui habet aures audiendi, audiat ".
LUKE|8|9|Interrogabant autem eum discipuli eius, quae esset haec parabola.
LUKE|8|10|Quibus ipse dixit: " Vobis datum est nosse mysteria regni Dei, ceteris autem in parabolis, ut videntes non videant et audientes non intellegant.
LUKE|8|11|Est autem haec parabola: Semen est verbum Dei.
LUKE|8|12|Qui autem secus viam, sunt qui audiunt; deinde venit Diabolus et tollit verbum de corde eorum, ne credentes salvi fiant.
LUKE|8|13|Qui autem supra petram: qui cum audierint, cum gaudio suscipiunt verbum; et hi radices non habent, qui ad tempus credunt, et in tempore tentationis recedunt.
LUKE|8|14|Quod autem in spinis cecidit: hi sunt, qui audierunt et a sollicitudinibus et divitiis et voluptatibus vitae euntes suffocantur et non referunt fructum.
LUKE|8|15|Quod autem in bonam terram: hi sunt, qui in corde bono et optimo audientes verbum retinent et fructum afferunt in patientia.
LUKE|8|16|Nemo autem lucernam accendens operit eam vaso aut subtus lectum ponit, sed supra candelabrum ponit, ut intrantes videant lumen.
LUKE|8|17|Non enim est occultum, quod non manifestetur, nec absconditum, quod non cognoscatur et in palam veniat.
LUKE|8|18|Videte ergo quomodo audiatis: qui enim habet, dabitur illi; et, quicumque non habet, etiam quod putat se habere, auferetur ab illo ".
LUKE|8|19|Venerunt autem ad illum mater et fratres eius, et non poterant adire ad eum prae turba.
LUKE|8|20|Et nuntiatum est illi: " Mater tua et fratres tui stant foris volentes te videre ".
LUKE|8|21|Qui respondens dixit ad eos: " Mater mea et fratres mei hi sunt, qui verbum Dei audiunt et faciunt ".
LUKE|8|22|Factum est autem in una dierum, et ipse ascendit in navem et discipuli eius, et ait ad illos: " Transfretemus trans stagnum ". Et ascenderunt.
LUKE|8|23|Navigantibus autem illis, obdormivit. Et descendit procella venti in stagnum, et complebantur et periclitabantur.
LUKE|8|24|Accedentes autem suscitaverunt eum dicentes: " Praeceptor, praeceptor, perimus! ". At ille surgens increpavit ventum et tempestatem aquae, et cessaverunt, et facta est tranquillitas.
LUKE|8|25|Dixit autem illis: " Ubi est fides vestra? ". Qui timentes mirati sunt dicentes ad invicem: " Quis putas hic est, quia et ventis imperat et aquae, et oboediunt ei? ".
LUKE|8|26|Enavigaverunt autem ad regionem Gergesenorum, quae est contra Galilaeam.
LUKE|8|27|Et cum egressus esset ad terram, occurrit illi vir quidam de civitate, qui habebat daemonia et iam tempore multo vestimento non induebatur neque in domo manebat sed in monumentis.
LUKE|8|28|Is ut vidit Iesum, exclamans procidit ante illum et voce magna dixit: " Quid mihi et tibi est, Iesu, Fili Dei Altissimi? Obsecro te, ne me torqueas ".
LUKE|8|29|Praecipiebat enim spiritui immundo, ut exiret ab homine. Multis enim temporibus arripiebat illum, vinciebatur catenis et compedibus custoditus; et ruptis vinculis, agebatur a daemonio in deserta.
LUKE|8|30|Interrogavit autem illum Iesus dicens: " Quod tibi nomen est? ". At ille dixit: " Legio ", quia intraverunt daemonia multa in eum.
LUKE|8|31|Et rogabant eum, ne imperaret illis, ut in abyssum irent.
LUKE|8|32|Erat autem ibi grex porcorum multorum pascentium in monte; et rogaverunt eum, ut permitteret eis in illos ingredi. Et permisit illis.
LUKE|8|33|Exierunt ergo daemonia ab homine et intraverunt in porcos, et impetu abiit grex per praeceps in stagnum et suffocatus est.
LUKE|8|34|Quod ut viderunt factum, qui pascebant, fugerunt et nuntiaverunt in civitatem et in villas.
LUKE|8|35|Exierunt autem videre, quod factum est, et venerunt ad Iesum et invenerunt hominem sedentem, a quo daemonia exierant, vestitum ac sana mente ad pedes Iesu et timuerunt.
LUKE|8|36|Nuntiaverunt autem illis hi, qui viderant, quomodo sanus factus esset, qui a daemonio vexabatur.
LUKE|8|37|Et rogaverunt illum omnis multitudo regionis Gergesenorum, ut discederet ab ipsis, quia timore magno tenebantur. Ipse autem ascendens navem reversus est.
LUKE|8|38|Et rogabat illum vir, a quo daemonia exierant, ut cum eo esset. Dimisit autem eum dicens:
LUKE|8|39|" Redi domum tuam et narra quanta tibi fecit Deus ". Et abiit per universam civitatem praedicans quanta illi fecisset Iesus.
LUKE|8|40|Cum autem rediret Iesus, excepit illum turba; erant enim omnes exspectantes eum.
LUKE|8|41|Et ecce venit vir, cui nomen Iairus, et ipse princeps synagogae erat, et cecidit ad pedes Iesu rogans eum, ut intraret in domum eius,
LUKE|8|42|quia filia unica erat illi fere annorum duodecim, et haec moriebatur. Et dum iret, a turbis comprimebatur.
LUKE|8|43|Et mulier quaedam erat in fluxu sanguinis ab annis duodecim, quae in medicos erogaverat omnem substantiam suam nec ab ullo potuit curari;
LUKE|8|44|accessit retro et tetigit fimbriam vestimenti eius, et confestim stetit fluxus sanguinis eius.
LUKE|8|45|Et ait Iesus: " Quis est, qui me tetigit? ". Negantibus autem omnibus, dixit Petrus: " Praeceptor, turbae te comprimunt et affligunt ".
LUKE|8|46|At dixit Iesus: " Tetigit me aliquis; nam et ego novi virtutem de me exisse ".
LUKE|8|47|Videns autem mulier quia non latuit, tremens venit et procidit ante eum et ob quam causam tetigerit eum indicavit coram omni populo et quemadmodum confestim sanata sit.
LUKE|8|48|At ipse dixit illi: " Filia, fides tua te salvam fecit. Vade in pace ".
LUKE|8|49|Adhuc illo loquente, venit quidam e domo principis synagogae dicens: " Mortua est filia tua; noli amplius vexare magistrum ".
LUKE|8|50|Iesus autem, audito hoc verbo, respondit ei: " Noli timere; crede tantum, et salva erit ".
LUKE|8|51|Et cum venisset domum, non permisit intrare secum quemquam nisi Petrum et Ioannem et Iacobum et patrem puellae et matrem.
LUKE|8|52|Flebant autem omnes et plangebant illam. At ille dixit: " Nolite flere; non est enim mortua, sed dormit ".
LUKE|8|53|Et deridebant eum scientes quia mortua esset.
LUKE|8|54|Ipse autem tenens manum eius clamavit dicens: " Puella, surge! ".
LUKE|8|55|Et reversus est spiritus eius, et surrexit continuo; et iussit illi dari manducare.
LUKE|8|56|Et stupuerunt parentes eius, quibus praecepit, ne alicui dicerent, quod factum erat.
LUKE|9|1|Convocatis autem Duodecim, dedit illis virtutem et potesta tem super omnia daemonia, et ut languores curarent,
LUKE|9|2|et misit illos praedicare regnum Dei et sanare infirmos;
LUKE|9|3|et ait ad illos: " Nihil tuleritis in via, neque virgam neque peram neque panem neque pecuniam, neque duas tunicas habeatis.
LUKE|9|4|Et in quamcumque domum intraveritis, ibi manete et inde exite.
LUKE|9|5|Et quicumque non receperint vos, exeuntes de civitate illa pulverem pedum vestrorum excutite in testimonium supra illos ".
LUKE|9|6|Egressi autem circumibant per castella evangelizantes et curantes ubique.
LUKE|9|7|Audivit autem Herodes tetrarcha omnia, quae fiebant, et haesitabat, eo quod diceretur a quibusdam: " Ioannes surrexit a mortuis ";
LUKE|9|8|a quibusdam vero: " Elias apparuit "; ab aliis autem: " Propheta unus de antiquis surrexit ".
LUKE|9|9|Et ait Herodes: " Ioannem ego decollavi; quis autem est iste, de quo audio ego talia? ". Et quaerebat videre eum.
LUKE|9|10|Et reversi apostoli narraverunt illi, quaecumque fecerunt. Et assumptis illis, secessit seorsum ad civitatem, quae vocatur Bethsaida.
LUKE|9|11|Quod cum cognovissent turbae, secutae sunt illum. Et excepit illos et loquebatur illis de regno Dei et eos, qui cura indigebant, sanabat.
LUKE|9|12|Dies autem coeperat declinare; et accedentes Duodecim dixerunt illi: " Dimitte turbam, ut euntes in castella villasque, quae circa sunt, divertant et inveniant escas, quia hic in loco deserto sumus ".
LUKE|9|13|Ait autem ad illos: " Vos date illis manducare ". At illi dixerunt: " Non sunt nobis plus quam quinque panes et duo pisces, nisi forte nos eamus et emamus in omnem hanc turbam escas ".
LUKE|9|14|Erant enim fere viri quinque milia. Ait autem ad discipulos suos: " Facite illos discumbere per convivia ad quinquagenos ".
LUKE|9|15|Et ita fecerunt et discumbere fecerunt omnes.
LUKE|9|16|Acceptis autem quinque panibus et duobus piscibus, respexit in caelum et benedixit illis et fregit et dabat discipulis suis, ut ponerent ante turbam.
LUKE|9|17|Et manducaverunt et saturati sunt omnes; et sublatum est, quod superfuit illis, fragmentorum cophini duodecim.
LUKE|9|18|Et factum est, cum solus esset orans, erant cum illo discipuli, et interrogavit illos dicens: " Quem me dicunt esse turbae? ".
LUKE|9|19|At illi responderunt et dixerunt: " Ioannem Baptistam, alii autem Eliam, alii vero: Propheta unus de prioribus surrexit ".
LUKE|9|20|Dixit autem illis: " Vos autem quem me esse dicitis? ". Respondens Petrus dixit: " Christum Dei ".
LUKE|9|21|At ille increpans illos praecepit, ne cui dicerent hoc,
LUKE|9|22|dicens: " Oportet Filium hominis multa pati et reprobari a senioribus et principibus sacerdotum et scribis et occidi et tertia die resurgere ".
LUKE|9|23|Dicebat autem ad omnes: " Si quis vult post me venire, abneget semetipsum et tollat crucem suam cotidie et sequatur me.
LUKE|9|24|Qui enim voluerit animam suam salvam facere, perdet illam; qui autem perdiderit animam suam propter me, hic salvam faciet illam.
LUKE|9|25|Quid enim proficit homo, si lucretur universum mundum, se autem ipsum perdat vel detrimentum sui faciat?
LUKE|9|26|Nam qui me erubuerit et meos sermones, hunc Filius hominis erubescet, cum venerit in gloria sua et Patris et sanctorum angelorum.
LUKE|9|27|Dico autem vobis vere: Sunt aliqui hic stantes, qui non gustabunt mortem, donec videant regnum Dei ".
LUKE|9|28|Factum est autem post haec verba fere dies octo, et assumpsit Petrum et Ioannem et Iacobum et ascendit in montem, ut oraret.
LUKE|9|29|Et facta est, dum oraret, species vultus eius altera, et vestitus eius albus, refulgens.
LUKE|9|30|Et ecce duo viri loquebantur cum illo, et erant Moyses et Elias,
LUKE|9|31|qui visi in gloria dicebant exodum eius, quam completurus erat in Ierusalem.
LUKE|9|32|Petrus vero et qui cum illo gravati erant somno; et evigilantes viderunt gloriam eius et duos viros, qui stabant cum illo.
LUKE|9|33|Et factum est, cum discederent ab illo, ait Petrus ad Iesum: " Praeceptor, bonum est nos hic esse; et faciamus tria tabernacula: unum tibi et unum Moysi et unum Eliae ", nesciens quid diceret.
LUKE|9|34|Haec autem illo loquente, facta est nubes et obumbravit eos; et timuerunt intrantibus illis in nubem.
LUKE|9|35|Et vox facta est de nube dicens: " Hic est Filius meus electus; ipsum audite ".
LUKE|9|36|Et dum fieret vox, inventus est Iesus solus. Et ipsi tacuerunt et nemini dixerunt in illis diebus quidquam ex his, quae viderant.
LUKE|9|37|Factum est autem in sequenti die, descendentibus illis de monte, occurrit illi turba multa.
LUKE|9|38|Et ecce vir de turba exclamavit dicens: " Magister, obsecro te, respice in filium meum, quia unicus est mihi;
LUKE|9|39|et ecce spiritus apprehendit illum, et subito clamat, et dissipat eum cum spuma et vix discedit ab eo dilanians eum;
LUKE|9|40|et rogavi discipulos tuos, ut eicerent illum, et non potuerunt ".
LUKE|9|41|Respondens autem Iesus dixit: " O generatio infidelis et perversa, usquequo ero apud vos et patiar vos? Adduc huc filium tuum ".
LUKE|9|42|Et cum accederet, elisit illum daemonium et dissipavit. Et increpavit Iesus spiritum immundum et sanavit puerum et reddidit illum patri eius.
LUKE|9|43|Stupebant autem omnes in magnitudine Dei.Omnibusque mirantibus in omnibus, quae faciebat, dixit ad discipulos suos:
LUKE|9|44|" Ponite vos in auribus vestris sermones istos: Filius enim hominis futurum est ut tradatur in manus hominum ".
LUKE|9|45|At illi ignorabant verbum istud, et erat velatum ante eos, ut non sentirent illud, et time bant interrogare eum de hoc verbo.
LUKE|9|46|Intravit autem cogitatio in eos, quis eorum maior esset.
LUKE|9|47|At Iesus sciens cogitationem cordis illorum, apprehendens puerum statuit eum secus se
LUKE|9|48|et ait illis: " Quicumque susceperit puerum istum in nomine meo, me recipit; et, quicumque me receperit, recipit eum, qui me misit; nam qui minor est inter omnes vos, hic maior est ".
LUKE|9|49|Respondens autem Ioannes dixit: " Praeceptor, vidimus quendam in nomine tuo eicientem daemonia et prohibuimus eum, quia non sequitur nobiscum ".
LUKE|9|50|Et ait ad illum Iesus: " Nolite prohibere; qui enim non est adversus vos, pro vobis est ".
LUKE|9|51|Factum est autem, dum complerentur dies assumptionis eius, et ipse faciem suam firmavit, ut iret Ierusalem,
LUKE|9|52|et misit nuntios ante conspectum suum. Et euntes intraverunt in castellum Samaritanorum, ut pararent illi.
LUKE|9|53|Et non receperunt eum, quia facies eius erat euntis Ierusalem.
LUKE|9|54|Cum vidissent autem discipuli Iacobus et Ioannes, dixerunt: " Domine, vis dicamus, ut ignis descendat de caelo et consumat illos? ".
LUKE|9|55|Et conversus increpavit illos.
LUKE|9|56|Et ierunt in aliud castellum.
LUKE|9|57|Et euntibus illis in via, dixit quidam ad illum: " Sequar te, quocumque ieris ".
LUKE|9|58|Et ait illi Iesus: " Vulpes foveas habent, et volucres caeli nidos, Filius autem hominis non habet, ubi caput reclinet ".
LUKE|9|59|Ait autem ad alterum: " Sequere me ". Ille autem dixit: " Domine, permitte mihi primum ire et sepelire patrem meum ".
LUKE|9|60|Dixitque ei Iesus: " Sine, ut mortui sepeliant mortuos suos; tu autem vade, annuntia regnum Dei ".
LUKE|9|61|Et ait alter: " Sequar te, Domine, sed primum permitte mihi renuntiare his, qui domi sunt ".
LUKE|9|62|Ait ad illum Iesus: " Nemo mittens manum suam in aratrum et aspiciens retro, aptus est regno Dei ".
LUKE|10|1|Post haec autem designavit Dominus alios septuaginta duos et misit illos binos ante faciem suam in omnem civitatem et locum, quo erat ipse venturus.
LUKE|10|2|Et dicebat illis: " Messis quidem multa, operarii autem pauci; rogate ergo Dominum messis, ut mittat operarios in messem suam.
LUKE|10|3|Ite; ecce ego mitto vos sicut agnos inter lupos.
LUKE|10|4|Nolite portare sacculum neque peram neque calceamenta et neminem per viam salutaveritis.
LUKE|10|5|In quamcumque domum intraveritis, primum dicite: "Pax huic domui".
LUKE|10|6|Et si ibi fuerit filius pacis, requiescet super illam pax vestra; sin autem, ad vos revertetur.
LUKE|10|7|In eadem autem domo manete edentes et bibentes, quae apud illos sunt: dignus enim est operarius mercede sua. Nolite transire de domo in domum.
LUKE|10|8|Et in quamcumque civitatem intraveritis, et susceperint vos, manducate, quae apponuntur vobis,
LUKE|10|9|et curate infirmos, qui in illa sunt, et dicite illis: "Appropinquavit in vos regnum Dei".
LUKE|10|10|In quamcumque civitatem intraveritis, et non receperint vos, exeuntes in plateas eius dicite:
LUKE|10|11|"Etiam pulverem, qui adhaesit nobis ad pedes de civitate vestra, extergimus in vos; tamen hoc scitote, quia appropinquavit regnum Dei".
LUKE|10|12|Dico vobis quia Sodomis in die illa remissius erit quam illi civitati.
LUKE|10|13|Vae tibi, Chorazin! Vae tibi, Bethsaida! Quia si in Tyro et Sidone factae fuissent virtutes, quae in vobis factae sunt, olim in cilicio et cinere sedentes paeniterent.
LUKE|10|14|Verumtamen Tyro et Sidoni remissius erit in iudicio quam vobis.
LUKE|10|15|Et tu, Capharnaum, numquid usque in caelum exaltaberis? Usque ad infernum demergeris!
LUKE|10|16|Qui vos audit, me audit; et, qui vos spernit, me spernit; qui autem me spernit, spernit eum, qui me misit ".
LUKE|10|17|Reversi sunt autem septuaginta duo cum gaudio dicentes: " Domine, etiam daemonia subiciuntur nobis in nomine tuo! ".
LUKE|10|18|Et ait illis: " Videbam Satanam sicut fulgur de caelo cadentem.
LUKE|10|19|Ecce dedi vobis potestatem calcandi supra serpentes et scorpiones et supra omnem virtutem inimici; et nihil vobis nocebit.
LUKE|10|20|Verumtamen in hoc nolite gaudere, quia spiritus vobis subiciuntur; gaudete autem quod nomina vestra scripta sunt in caelis ".
LUKE|10|21|In ipsa hora exsultavit Spiritu Sancto et dixit: " Confiteor tibi, Pater, Domine caeli et terrae, quod abscondisti haec a sapientibus et prudentibus et revelasti ea parvulis; etiam, Pater, quia sic placuit ante te.
LUKE|10|22|Omnia mihi tradita sunt a Patre meo; et nemo scit qui sit Filius, nisi Pater, et qui sit Pater, nisi Filius et cui voluerit Filius revelare ".
LUKE|10|23|Et conversus ad discipulos seorsum dixit: " Beati oculi, qui vident, quae videtis.
LUKE|10|24|Dico enim vobis: Multi prophetae et reges voluerunt videre, quae vos videtis, et non viderunt, et audire, quae auditis, et non audierunt ".
LUKE|10|25|Et ecce quidam legis peritus surrexit tentans illum dicens: " Magister, quid faciendo vitam aeternam possidebo? ".
LUKE|10|26|At ille dixit ad eum: " In Lege quid scriptum est? Quomodo legis? ".
LUKE|10|27|Ille autem respondens dixit: " Diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex omnibus viribus tuis et ex omni mente tua et proximum tuum sicut teipsum ".
LUKE|10|28|Dixitque illi: " Recte respondisti; hoc fac et vives ".
LUKE|10|29|Ille autem, volens iustificare seipsum, dixit ad Iesum: " Et quis est meus proximus? ".
LUKE|10|30|Suscipiens autem Iesus dixit: " Homo quidam descendebat ab Ierusalem in Iericho et incidit in latrones, qui etiam despoliaverunt eum et, plagis impositis, abierunt, semivivo relicto.
LUKE|10|31|Accidit autem, ut sacerdos quidam descenderet eadem via et, viso illo, praeterivit;
LUKE|10|32|similiter et Levita, cum esset secus locum et videret eum, pertransiit.
LUKE|10|33|Samaritanus autem quidam iter faciens, venit secus eum et videns eum misericordia motus est,
LUKE|10|34|et appropians alligavit vulnera eius infundens oleum et vinum; et imponens illum in iumentum suum duxit in stabulum et curam eius egit.
LUKE|10|35|Et altera die protulit duos denarios et dedit stabulario et ait: "Curam illius habe, et, quodcumque supererogaveris, ego, cum rediero, reddam tibi".
LUKE|10|36|Quis horum trium videtur tibi proximus fuisse illi, qui incidit in latrones? ".
LUKE|10|37|At ille dixit: " Qui fecit misericordiam in illum ". Et ait illi Iesus: Vade et tu fac similiter ".
LUKE|10|38|Cum autem irent, ipse intravit in quoddam castellum, et mulier quaedam Martha nomine excepit illum.
LUKE|10|39|Et huic erat soror nomine Maria, quae etiam sedens secus pedes Domini audiebat verbum illius.
LUKE|10|40|Martha autem satagebat circa frequens ministerium; quae stetit et ait: Domine, non est tibi curae quod soror mea reliquit me solam ministrare? Dic ergo illi, ut me adiuvet ".
LUKE|10|41|Et respondens dixit illi Dominus: " Martha, Martha, sollicita es et turbaris erga plurima,
LUKE|10|42|porro unum est necessarium; Maria enim optimam partem elegit, quae non auferetur ab ea ".
LUKE|11|1|Et factum est cum esset in loco quodam orans, ut cessa vit, dixit unus ex discipulis eius ad eum: " Domine, doce nos orare, sicut et Ioannes docuit discipulos suos ".
LUKE|11|2|Et ait illis: " Cum oratis, dicite:Pater, sanctificetur nomen tuum,adveniat regnum tuum;
LUKE|11|3|panem nostrum cotidianum da nobis cotidie,
LUKE|11|4|et dimitte nobis peccata nostra,si quidem et ipsi dimittimus omni debenti nobis,et ne nos inducas in tentationem ".
LUKE|11|5|Et ait ad illos: " Quis vestrum habebit amicum et ibit ad illum media nocte et dicet illi: "Amice, commoda mihi tres panes,
LUKE|11|6|quoniam amicus meus venit de via ad me, et non habeo, quod ponam ante illum";
LUKE|11|7|et ille de intus respondens dicat: "Noli mihi molestus esse; iam ostium clausum est, et pueri mei mecum sunt in cubili; non possum surgere et dare tibi".
LUKE|11|8|Dico vobis: Et si non dabit illi surgens, eo quod amicus eius sit, propter improbitatem tamen eius surget et dabit illi, quotquot habet necessarios.
LUKE|11|9|Et ego vobis dico: Petite, et dabitur vobis; quaerite, et invenietis; pulsate, et aperietur vobis.
LUKE|11|10|Omnis enim qui petit, accipit; et, qui quaerit, invenit; et pulsanti aperietur.
LUKE|11|11|Quem autem ex vobis patrem filius petierit piscem, numquid pro pisce serpentem dabit illi?
LUKE|11|12|Aut si petierit ovum, numquid porriget illi scorpionem?
LUKE|11|13|Si ergo vos, cum sitis mali, nostis dona bona dare filiis vestris, quanto magis Pater de caelo dabit Spiritum Sanctum petentibus se ".
LUKE|11|14|Et erat eiciens daemonium, et illud erat mutum; et factum est, cum daemonium exisset, locutus est mutus. Et admiratae sunt turbae;
LUKE|11|15|quidam autem ex eis dixerunt: " In Beelzebul principe daemoniorum eicit daemonia ".
LUKE|11|16|Et alii tentantes signum de caelo quaerebant ab eo.
LUKE|11|17|Ipse autem sciens cogitationes eorum dixit eis: " Omne regnum in seipsum divisum desolatur, et domus supra domum cadit.
LUKE|11|18|Si autem et Satanas in seipsum divisus est, quomodo stabit regnum ipsius? Quia dicitis in Beelzebul eicere me daemonia.
LUKE|11|19|Si autem ego in Beelzebul eicio daemonia, filii vestri in quo eiciunt? Ideo ipsi iudices vestri erunt.
LUKE|11|20|Porro si in digito Dei eicio daemonia, profecto pervenit in vos regnum Dei.
LUKE|11|21|Cum fortis armatus custodit atrium suum, in pace sunt ea, quae possidet;
LUKE|11|22|si autem fortior illo superveniens vicerit eum, universa arma eius auferet, in quibus confidebat, et spolia eius distribuet.
LUKE|11|23|Qui non est mecum, adversum me est; et, qui non colligit mecum, dispergit.
LUKE|11|24|Cum immundus spiritus exierit de homine, perambulat per loca inaquosa quaerens requiem; et non inveniens dicit: "Revertar in domum meam unde exivi".
LUKE|11|25|Et cum venerit, invenit scopis mundatam et exornatam.
LUKE|11|26|Et tunc vadit et assumit septem alios spiritus nequiores se, et ingressi habitant ibi; et sunt novissima hominis illius peiora prioribus.
LUKE|11|27|Factum est autem, cum haec diceret, extollens vocem quaedam mulier de turba dixit illi: " Beatus venter, qui te portavit, et ubera, quae suxisti! ".
LUKE|11|28|At ille dixit: " Quinimmo beati, qui audiunt verbum Dei et custodiunt!.
LUKE|11|29|Turbis autem concurrentibus, coepit dicere: " Generatio haec generatio nequam est; signum quaerit, et signum non dabitur illi, nisi signum Ionae.
LUKE|11|30|Nam sicut Ionas fuit signum Ninevitis, ita erit et Filius hominis generationi isti.
LUKE|11|31|Regina austri surget in iudicio cum viris generationis huius et condemnabit illos, quia venit a finibus terrae audire sapientiam Salomonis, et ecce plus Salomone hic.
LUKE|11|32|Viri Ninevitae surgent in iudicio cum generatione hac et condemnabunt illam, quia paenitentiam egerunt ad praedicationem Ionae, et ecce plus Iona hic.
LUKE|11|33|Nemo lucernam accendit et in abscondito ponit neque sub modio sed supra candelabrum, ut, qui ingrediuntur, lumen videant.
LUKE|11|34|Lucerna corporis est oculus tuus. Si oculus tuus fuerit simplex, totum corpus tuum lucidum erit; si autem nequam fuerit, etiam corpus tuum tenebrosum erit.
LUKE|11|35|Vide ergo, ne lumen, quod in te est, tenebrae sint.
LUKE|11|36|Si ergo corpus tuum totum lucidum fuerit non habens aliquam partem tenebrarum, erit lucidum totum, sicut quando lucerna in fulgore suo illuminat te ".
LUKE|11|37|Et cum loqueretur, rogavit illum quidam pharisaeus, ut pranderet apud se; et ingressus recubuit.
LUKE|11|38|Pharisaeus autem videns miratus est quod non baptizatus esset ante prandium.
LUKE|11|39|Et ait Dominus ad illum: " Nunc vos pharisaei, quod de foris est calicis et catini, mundatis; quod autem intus est vestrum, plenum est rapina et iniquitate.
LUKE|11|40|Stulti! Nonne, qui fecit, quod de foris est, etiam id, quod de intus est, fecit?
LUKE|11|41|Verumtamen, quae insunt, date eleemosynam; et ecce omnia munda sunt vobis.
LUKE|11|42|Sed vae vobis pharisaeis, quia decimatis mentam et rutam et omne holus et praeteritis iudicium et caritatem Dei! Haec autem oportuit facere et illa non omittere.
LUKE|11|43|Vae vobis pharisaeis, quia diligitis primam cathedram in synagogis et salutationes in foro!
LUKE|11|44|Vae vobis, quia estis ut monumenta, quae non parent, et homines ambulantes supra nesciunt! ".
LUKE|11|45|Respondens autem quidam ex legis peritis ait illi: " Magister, haec dicens etiam nobis contumeliam facis ".
LUKE|11|46|At ille ait: " Et vobis legis peritis: Vae, quia oneratis homines oneribus, quae portari non possunt, et ipsi uno digito vestro non tangitis sarcinas!
LUKE|11|47|Vae vobis, quia aedificatis monumenta prophetarum, patres autem vestri occiderunt illos!
LUKE|11|48|Profecto testificamini et consentitis operibus patrum vestrorum, quoniam ipsi quidem eos occiderunt, vos autem aedificatis.
LUKE|11|49|Propterea et sapientia Dei dixit: Mittam ad illos prophetas et apostolos, et ex illis occident et persequentur,
LUKE|11|50|ut requiratur sanguis omnium prophetarum, qui effusus est a constitutione mundi, a generatione ista,
LUKE|11|51|a sanguine Abel usque ad sanguinem Zachariae, qui periit inter altare et aedem. Ita dico vobis: Requiretur ab hac generatione.
LUKE|11|52|Vae vobis legis peritis, quia tulistis clavem scientiae! Ipsi non introistis et eos, qui introibant, prohibuistis ".
LUKE|11|53|Cum autem inde exisset, coeperunt scribae et pharisaei graviter insistere et eum allicere in sermone de multis
LUKE|11|54|insidiantes ei, ut caperent aliquid ex ore eius.
LUKE|12|1|Interea multis turbis cir cumstantibus, ita ut se invi cem conculcarent, coepit dicere ad discipulos suos primum: " Attendite a fermento pharisaeorum, quod est hypocrisis.
LUKE|12|2|Nihil autem opertum est, quod non reveletur, neque absconditum, quod non sciatur.
LUKE|12|3|Quoniam, quae in tenebris dixistis, in lumine audientur; et, quod in aurem locuti estis in cubiculis, praedicabitur in tectis.
LUKE|12|4|Dico autem vobis amicis meis: Ne terreamini ab his, qui occidunt corpus et post haec non habent amplius, quod faciant.
LUKE|12|5|Ostendam autem vobis quem timeatis: Timete eum, qui postquam occiderit, habet potestatem mittere in gehennam. Ita dico vobis: Hunc timete.
LUKE|12|6|Nonne quinque passeres veneunt dipundio? Et unus ex illis non est in oblivione coram Deo.
LUKE|12|7|Sed et capilli capitis vestri omnes numerati sunt. Nolite timere; multis passeribus pluris estis.
LUKE|12|8|Dico autem vobis: Omnis, quicumque confessus fuerit in me coram hominibus, et Filius hominis confitebitur in illo coram angelis Dei;
LUKE|12|9|qui autem negaverit me coram hominibus, denegabitur coram angelis Dei.
LUKE|12|10|Et omnis, qui dicet verbum in Filium hominis, remittetur illi; ei autem, qui in Spiritum Sanctum blasphemaverit, non remittetur.
LUKE|12|11|Cum autem inducent vos in synagogas et ad magistratus et potestates, nolite solliciti esse qualiter aut quid respondeatis aut quid dicatis:
LUKE|12|12|Spiritus enim Sanctus docebit vos in ipsa hora, quae oporteat dicere ".
LUKE|12|13|Ait autem quidam ei de turba: " Magister, dic fratri meo, ut dividat mecum hereditatem ".
LUKE|12|14|At ille dixit ei: " Homo, quis me constituit iudicem aut divisorem super vos? ".
LUKE|12|15|Dixitque ad illos: " Videte et cavete ab omni avaritia, quia si cui res abundant, vita eius non est ex his, quae possidet ".
LUKE|12|16|Dixit autem similitudinem ad illos dicens: " Hominis cuiusdam divitis uberes fructus ager attulit.
LUKE|12|17|Et cogitabat intra se dicens: "Quid faciam, quod non habeo, quo congregem fructus meos?".
LUKE|12|18|Et dixit: "Hoc faciam: destruam horrea mea et maiora aedificabo et illuc congregabo omne triticum et bona mea;
LUKE|12|19|et dicam animae meae: Anima, habes multa bona posita in annos plurimos; requiesce, comede, bibe, epulare".
LUKE|12|20|Dixit autem illi Deus: "Stulte! Hac nocte animam tuam repetunt a te; quae autem parasti, cuius erunt?".
LUKE|12|21|Sic est qui sibi thesaurizat et non fit in Deum dives ".
LUKE|12|22|Dixitque ad discipulos suos: " Ideo dico vobis: nolite solliciti esse animae quid manducetis, neque corpori quid vestiamini.
LUKE|12|23|Anima enim plus est quam esca, et corpus quam vestimentum.
LUKE|12|24|Considerate corvos, quia non seminant neque metunt, quibus non est cellarium neque horreum, et Deus pascit illos; quanto magis vos pluris estis volucribus.
LUKE|12|25|Quis autem vestrum cogitando potest adicere ad aetatem suam cubitum?
LUKE|12|26|Si ergo neque, quod minimum est, potestis, quid de ceteris solliciti estis?
LUKE|12|27|Considerate lilia quomodo crescunt: non laborant neque nent; dico autem vobis: Nec Salomon in omni gloria sua vestiebatur sicut unum ex istis.
LUKE|12|28|Si autem fenum, quod hodie in agro est et cras in clibanum mittitur, Deus sic vestit, quanto magis vos, pusillae fidei.
LUKE|12|29|Et vos nolite quaerere quid manducetis aut quid bibatis et nolite solliciti esse.
LUKE|12|30|Haec enim omnia gentes mundi quaerunt; Pater autem vester scit quoniam his indigetis.
LUKE|12|31|Verumtamen quaerite regnum eius; et haec adicientur vobis.
LUKE|12|32|Noli timere, pusillus grex, quia complacuit Patri vestro dare vobis regnum.
LUKE|12|33|Vendite, quae possidetis, et date eleemosynam. Facite vobis sacculos, qui non veterescunt, thesaurum non deficientem in caelis, quo fur non appropiat, neque tinea corrumpit;
LUKE|12|34|ubi enim thesaurus vester est, ibi et cor vestrum erit.
LUKE|12|35|Sint lumbi vestri praecincti et lucernae ardentes,
LUKE|12|36|et vos similes hominibus exspectantibus dominum suum, quando revertatur a nuptiis, ut, cum venerit et pulsaverit, confestim aperiant ei.
LUKE|12|37|Beati, servi illi, quos, cum venerit dominus, invenerit vigilantes. Amen dico vobis, quod praecinget se et faciet illos discumbere et transiens ministrabit illis.
LUKE|12|38|Et si venerit in secunda vigilia, et si in tertia vigilia venerit, et ita invenerit, beati sunt illi.
LUKE|12|39|Hoc autem scitote, quia, si sciret pater familias, qua hora fur veniret, non sineret perfodi domum suam.
LUKE|12|40|Et vos estote parati, quia, qua hora non putatis, Filius hominis venit.
LUKE|12|41|Ait autem Petrus: " Domine, ad nos dicis hanc parabolam an et ad omnes?.
LUKE|12|42|Et dixit Dominus: " Quis putas est fidelis dispensator et prudens, quem constituet dominus super familiam suam, ut det illis in tempore tritici mensuram?
LUKE|12|43|Beatus ille servus, quem, cum venerit dominus eius, invenerit ita facientem.
LUKE|12|44|Vere dico vobis: Supra omnia, quae possidet, constituet illum.
LUKE|12|45|Quod si dixerit servus ille in corde suo: "Moram facit dominus meus venire", et coeperit percutere pueros et ancillas et edere et bibere et inebriari,
LUKE|12|46|veniet dominus servi illius in die, qua non sperat, et hora, qua nescit, et dividet eum partemque eius cum infidelibus ponet.
LUKE|12|47|Ille autem servus, qui cognovit voluntatem domini sui et non praeparavit vel non fecit secundum voluntatem eius, vapulabit multis;
LUKE|12|48|qui autem non cognovit et fecit digna plagis, vapulabit paucis. Omni autem, cui multum datum est, multum quaeretur ab eo; et cui commendaverunt multum, plus petent ab eo.
LUKE|12|49|Ignem veni mittere in terram et quid volo? Si iam accensus esset!
LUKE|12|50|Baptisma autem habeo baptizari et quomodo coartor, usque dum perficiatur!
LUKE|12|51|Putatis quia pacem veni dare in terram? Non, dico vobis, sed separationem.
LUKE|12|52|Erunt enim ex hoc quinque in domo una divisi: tres in duo, et duo in tres;
LUKE|12|53|dividentur pater in filium et filius in patrem, mater in filiam et filia in matrem, socrus in nurum suam et nurus in socrum ".
LUKE|12|54|Dicebat autem et ad turbas: " Cum videritis nubem orientem ab occasu, statim dicitis: "Nimbus venit", et ita fit;
LUKE|12|55|et cum austrum flantem, dicitis: "Aestus erit", et fit.
LUKE|12|56|Hypocritae, faciem terrae et caeli nostis probare, hoc autem tempus quomodo nescitis probare?
LUKE|12|57|Quid autem et a vobis ipsis non iudicatis, quod iustum est?
LUKE|12|58|Cum autem vadis cum adversario tuo ad principem, in via da operam liberari ab illo, ne forte trahat te apud iudicem, et iudex tradat te exactori, et exactor mittat te in carcerem.
LUKE|12|59|Dico tibi: Non exies inde, donec etiam novissimum minutum reddas ".
LUKE|13|1|Aderant autem quidam ipso in tempore nuntiantes illi de Galilaeis, quorum sanguinem Pilatus miscuit cum sacrificiis eorum.
LUKE|13|2|Et respondens dixit illis: " Putatis quod hi Galilaei prae omnibus Galilaeis peccatores fuerunt, quia talia passi sunt?
LUKE|13|3|Non, dico vobis, sed, nisi paenitentiam egeritis, omnes similiter peribitis.
LUKE|13|4|Vel illi decem et octo, supra quos cecidit turris in Siloam et occidit eos, putatis quia et ipsi debitores fuerunt praeter omnes homines habitantes in Ierusalem?
LUKE|13|5|Non, dico vobis, sed, si non paenitentiam egeritis, omnes similiter peribitis ".
LUKE|13|6|Dicebat autem hanc similitudinem: " Arborem fici habebat quidam plantatam in vinea sua et venit quaerens fructum in illa et non invenit.
LUKE|13|7|Dixit autem ad cultorem vineae: "Ecce anni tres sunt, ex quo venio quaerens fructum in ficulnea hac et non invenio. Succide ergo illam. Ut quid etiam terram evacuat?".
LUKE|13|8|At ille respondens dicit illi: "Domine, dimitte illam et hoc anno, usque dum fodiam circa illam et mittam stercora,
LUKE|13|9|et si quidem fecerit fructum in futurum; sin autem succides eam" ".
LUKE|13|10|Erat autem docens in una synagogarum sabbatis.
LUKE|13|11|Et ecce mulier, quae habebat spiritum infirmitatis annis decem et octo et erat inclinata nec omnino poterat sursum respicere.
LUKE|13|12|Quam cum vidisset Iesus, vocavit et ait illi: " Mulier, dimissa es ab infirmitate tua ",
LUKE|13|13|et imposuit illi manus; et confestim erecta est et glorificabat Deum.
LUKE|13|14|Respondens autem archisynagogus, indignans quia sabbato curasset Iesus, dicebat turbae: " Sex dies sunt, in quibus oportet operari; in his ergo venite et curamini et non in die sabbati ".
LUKE|13|15|Respondit autem ad illum Dominus et dixit: " Hypocritae, unusquisque vestrum sabbato non solvit bovem suum aut asinum a praesepio et ducit adaquare?
LUKE|13|16|Hanc autem filiam Abrahae, quam alligavit Satanas ecce decem et octo annis, non oportuit solvi a vinculo isto die sabbati? ".
LUKE|13|17|Et cum haec diceret, erubescebant omnes adversarii eius, et omnis populus gaudebat in universis, quae gloriose fiebant ab eo.
LUKE|13|18|Dicebat ergo: " Cui simile est regnum Dei, et cui simile existimabo illud?
LUKE|13|19|Simile est grano sinapis, quod acceptum homo misit in hortum suum, et crevit et factum est in arborem, et volucres caeli requieverunt in ramis eius ".
LUKE|13|20|Et iterum dixit: " Cui simile aestimabo regnum Dei?
LUKE|13|21|Simile est fermento, quod acceptum mulier abscondit in farinae sata tria, donec fermentaretur totum ".
LUKE|13|22|Et ibat per civitates et castella docens et iter faciens in Hierosolymam.
LUKE|13|23|Ait autem illi quidam: " Domine, pauci sunt, qui salvantur? ". Ipse autem dixit ad illos:
LUKE|13|24|" Contendite intrare per angustam portam, quia multi, dico vobis, quaerent intrare et non poterunt.
LUKE|13|25|Cum autem surrexerit pater familias et clauserit ostium, et incipietis foris stare et pulsare ostium dicentes: "Domine, aperi nobis"; et respondens dicet vobis: "Nescio vos unde sitis".
LUKE|13|26|Tunc incipietis dicere: "Manducavimus coram te et bibimus, et in plateis nostris docuisti";
LUKE|13|27|et dicet loquens vobis: "Nescio vos unde sitis; discedite a me, omnes operarii iniquitatis".
LUKE|13|28|Ibi erit fletus et stridor dentium, cum videritis Abraham et Isaac et Iacob et omnes prophetas in regno Dei, vos autem expelli foras.
LUKE|13|29|Et venient ab oriente et occidente et aquilone et austro et accumbent in regno Dei.
LUKE|13|30|Et ecce sunt novissimi, qui erunt primi, et sunt primi, qui erunt novissimi ".
LUKE|13|31|In ipsa hora accesserunt quidam pharisaeorum dicentes illi: " Exi et vade hinc, quia Herodes vult te occidere ".
LUKE|13|32|Et ait illis: " Ite, dicite vulpi illi: "Ecce eicio daemonia et sanitates perficio hodie et cras et tertia consummor.
LUKE|13|33|Verumtamen oportet me hodie et cras et sequenti ambulare, quia non capit prophetam perire extra Ierusalem".
LUKE|13|34|Ierusalem, Ierusalem, quae occidis prophetas et lapidas eos, qui missi sunt ad te, quotiens volui congregare filios tuos, quemadmodum avis nidum suum sub pinnis, et noluistis.
LUKE|13|35|Ecce relinquitur vobis domus vestra. Dico autem vobis: Non videbitis me, donec veniat cum dicetis: "Benedictus, qui venit in nomine Domini" ".
LUKE|14|1|Et factum est, cum intraret in domum cuiusdam princi pis pharisaeorum sabbato manducare panem, et ipsi observabant eum.
LUKE|14|2|Et ecce homo quidam hydropicus erat ante illum.
LUKE|14|3|Et respondens Iesus dixit ad legis peritos et pharisaeos dicens: " Licet sabbato curare an non? ".
LUKE|14|4|At illi tacuerunt. Ipse vero apprehensum sanavit eum ac dimisit.
LUKE|14|5|Et ad illos dixit: " Cuius vestrum filius aut bos in puteum cadet, et non continuo extrahet illum die sabbati? ".
LUKE|14|6|Et non poterant ad haec respondere illi.
LUKE|14|7|Dicebat autem ad invitatos parabolam, intendens quomodo primos accubitus eligerent, dicens ad illos:
LUKE|14|8|" Cum invitatus fueris ab aliquo ad nuptias, non discumbas in primo loco, ne forte honoratior te sit invitatus ab eo,
LUKE|14|9|et veniens is qui te et illum vocavit, dicat tibi: "Da huic locum"; et tunc incipias cum rubore novissimum locum tenere.
LUKE|14|10|Sed cum vocatus fueris, vade, recumbe in novissimo loco, ut, cum venerit qui te invitavit, dicat tibi: "Amice, ascende superius"; tunc erit tibi gloria coram omnibus simul discumbentibus.
LUKE|14|11|Quia omnis, qui se exaltat, humiliabitur; et, qui se humiliat, exaltabitur ".
LUKE|14|12|Dicebat autem et ei, qui se invitaverat: " Cum facis prandium aut cenam, noli vocare amicos tuos neque fratres tuos neque cognatos neque vicinos divites, ne forte et ipsi te reinvitent, et fiat tibi retributio.
LUKE|14|13|Sed cum facis convivium, voca pauperes, debiles, claudos, caecos;
LUKE|14|14|et beatus eris, quia non habent retribuere tibi. Retribuetur enim tibi in resurrectione iustorum ".
LUKE|14|15|Haec cum audisset quidam de simul discumbentibus, dixit illi: " Beatus, qui manducabit panem in regno Dei ".
LUKE|14|16|At ipse dixit ei: " Homo quidam fecit cenam magnam et vocavit multos;
LUKE|14|17|et misit servum suum hora cenae dicere invitatis: "Venite, quia iam paratum est".
LUKE|14|18|Et coeperunt simul omnes excusare. Primus dixit ei: "Villam emi et necesse habeo exire et videre illam; rogo te, habe me excusatum".
LUKE|14|19|Et alter dixit: "Iuga boum emi quinque et eo probare illa; rogo te, habe me excusatum".
LUKE|14|20|Et alius dixit: "Uxorem duxi et ideo non possum venire".
LUKE|14|21|Et reversus servus nuntiavit haec domino suo. Tunc iratus pater familias dixit servo suo: "Exi cito in plateas et vicos civitatis et pauperes ac debiles et caecos et claudos introduc huc".
LUKE|14|22|Et ait servus: "Domine, factum est, ut imperasti, et adhuc locus est".
LUKE|14|23|Et ait dominus servo: "Exi in vias et saepes, et compelle intrare, ut impleatur domus mea.
LUKE|14|24|Dico autem vobis, quod nemo virorum illorum, qui vocati sunt, gustabit cenam meam" ".
LUKE|14|25|Ibant autem turbae multae cum eo; et conversus dixit ad illos:
LUKE|14|26|" Si quis venit ad me et non odit patrem suum et matrem et uxorem et filios et fratres et sorores, adhuc et animam suam, non potest esse meus discipulus.
LUKE|14|27|Et, qui non baiulat crucem suam et venit post me, non potest esse meus discipulus.
LUKE|14|28|Quis enim ex vobis volens turrem aedificare, non prius sedens computat sumptus, si habet ad perficiendum?
LUKE|14|29|Ne, posteaquam posuerit fundamentum et non potuerit perficere, omnes, qui vident, incipiant illudere ei
LUKE|14|30|dicentes: "Hic homo coepit aedificare et non potuit consummare".
LUKE|14|31|Aut quis rex, iturus committere bellum adversus alium regem, non sedens prius cogitat, si possit cum decem milibus occurrere ei, qui cum viginti milibus venit ad se?
LUKE|14|32|Alioquin, adhuc illo longe agente, legationem mittens rogat ea, quae pacis sunt.
LUKE|14|33|Sic ergo omnis ex vobis, qui non renuntiat omnibus, quae possidet, non potest meus esse discipulus.
LUKE|14|34|Bonum est sal; si autem sal quoque evanuerit, in quo condietur?
LUKE|14|35|Neque in terram neque in sterquilinium utile est, sed foras proiciunt illud. Qui habet aures audiendi, audiat ".
LUKE|15|1|Erant autem appropinquan tes ei omnes publicani et pec catores, ut audirent illum.
LUKE|15|2|Et murmurabant pharisaei et scribae dicentes: " Hic peccatores recipit et manducat cum illis ".
LUKE|15|3|Et ait ad illos parabolam istam dicens:
LUKE|15|4|" Quis ex vobis homo, qui habet centum oves et si perdiderit unam ex illis, nonne dimittit nonaginta novem in deserto et vadit ad illam, quae perierat, donec inveniat illam?
LUKE|15|5|Et cum invenerit eam, imponit in umeros suos gaudens
LUKE|15|6|et veniens domum convocat amicos et vicinos dicens illis: Congratulamini mihi, quia inveni ovem meam, quae perierat".
LUKE|15|7|Dico vobis: Ita gaudium erit in caelo super uno peccatore paenitentiam agente quam super nonaginta novem iustis, qui non indigent paenitentia.
LUKE|15|8|Aut quae mulier habens drachmas decem, si perdiderit drachmam unam, nonne accendit lucernam et everrit domum et quaerit diligenter, donec inveniat?
LUKE|15|9|Et cum invenerit, convocat amicas et vicinas dicens: "Congratulamini mihi, quia inveni drachmam, quam perdideram".
LUKE|15|10|Ita dico vobis: Gaudium fit coram angelis Dei super uno peccatore paenitentiam agente ".
LUKE|15|11|Ait autem: " Homo quidam habebat duos filios.
LUKE|15|12|Et dixit adulescentior ex illis patri: "Pater, da mihi portionem substantiae, quae me contingit". Et divisit illis substantiam.
LUKE|15|13|Et non post multos dies, congregatis omnibus, adulescentior filius peregre profectus est in regionem longinquam et ibi dissipavit substantiam suam vivendo luxuriose.
LUKE|15|14|Et postquam omnia consummasset, facta est fames valida in regione illa, et ipse coepit egere.
LUKE|15|15|Et abiit et adhaesit uni civium regionis illius, et misit illum in villam suam, ut pasceret porcos;
LUKE|15|16|et cupiebat saturari de siliquis, quas porci manducabant, et nemo illi dabat.
LUKE|15|17|In se autem reversus dixit: "Quanti mercennarii patris mei abundant panibus, ego autem hic fame pereo.
LUKE|15|18|Surgam et ibo ad patrem meum et dicam illi: Pater, peccavi in caelum et coram te
LUKE|15|19|et iam non sum dignus vocari filius tuus; fac me sicut unum de mercennariis tuis".
LUKE|15|20|Et surgens venit ad patrem suum.Cum autem adhuc longe esset, vidit illum pater ipsius et misericordia motus est et accurrens cecidit supra collum eius et osculatus est illum.
LUKE|15|21|Dixitque ei filius: "Pater, peccavi in caelum et coram te; iam non sum dignus vocari filius tuus".
LUKE|15|22|Dixit autem pater ad servos suos: "Cito proferte stolam primam et induite illum et date anulum in manum eius et calceamenta in pedes
LUKE|15|23|et adducite vitulum saginatum, occidite et manducemus et epulemur,
LUKE|15|24|quia hic filius meus mortuus erat et revixit, perierat et inventus est". Et coeperunt epulari.
LUKE|15|25|Erat autem filius eius senior in agro et, cum veniret et appropinquaret domui, audivit symphoniam et choros
LUKE|15|26|et vocavit unum de servis et interrogavit quae haec essent.
LUKE|15|27|Isque dixit illi: "Frater tuus venit, et occidit pater tuus vitulum saginatum, quia salvum illum recepit".
LUKE|15|28|Indignatus est autem et nolebat introire. Pater ergo illius egressus coepit rogare illum.
LUKE|15|29|At ille respondens dixit patri suo: "Ecce tot annis servio tibi et numquam mandatum tuum praeterii, et numquam dedisti mihi haedum, ut cum amicis meis epularer;
LUKE|15|30|sed postquam filius tuus hic, qui devoravit substantiam tuam cum meretricibus, venit, occidisti illi vitulum saginatum".
LUKE|15|31|At ipse dixit illi: "Fili, tu semper mecum es, et omnia mea tua sunt;
LUKE|15|32|epulari autem et gaudere oportebat, quia frater tuus hic mortuus erat et revixit, perierat et inventus est" ".
LUKE|16|1|Dicebat autem et ad disci pulos: " Homo quidam erat dives, qui habebat vilicum, et hic diffamatus est apud illum quasi dissipasset bona ipsius.
LUKE|16|2|Et vocavit illum et ait illi: "Quid hoc audio de te? Redde rationem vilicationis tuae; iam enim non poteris vilicare".
LUKE|16|3|Ait autem vilicus intra se: "Quid faciam, quia dominus meus aufert a me vilicationem? Fodere non valeo, mendicare erubesco.
LUKE|16|4|Scio quid faciam, ut, cum amotus fuero a vilicatione, recipiant me in domos suas".
LUKE|16|5|Convocatis itaque singulis debitoribus domini sui, dicebat primo: Quantum debes domino meo?".
LUKE|16|6|At ille dixit: "Centum cados olei". Dixitque illi: "Accipe cautionem tuam et sede cito, scribe quinquaginta".
LUKE|16|7|Deinde alii dixit: "Tu vero quantum debes?". Qui ait: "Centum coros tritici". Ait illi: "Accipe litteras tuas et scribe octoginta".
LUKE|16|8|Et laudavit dominus vilicum iniquitatis, quia prudenter fecisset, quia filii huius saeculi prudentiores filiis lucis in generatione sua sunt.
LUKE|16|9|Et ego vobis dico: Facite vobis amicos de mammona iniquitatis, ut, cum defecerit, recipiant vos in aeterna tabernacula.
LUKE|16|10|Qui fidelis est in minimo, et in maiori fidelis est; et, qui in modico iniquus est, et in maiori iniquus est.
LUKE|16|11|Si ergo in iniquo mammona fideles non fuistis, quod verum est, quis credet vobis?
LUKE|16|12|Et si in alieno fideles non fuistis, quod vestrum est, quis dabit vobis?
LUKE|16|13|Nemo servus potest duobus dominis servire: aut enim unum odiet et alterum diliget, aut uni adhaerebit et alterum contemnet. Non potestis Deo servire et mammonae ".
LUKE|16|14|Audiebant autem omnia haec pharisaei, qui erant avari, et deridebant illum.
LUKE|16|15|Et ait illis: " Vos estis, qui iustificatis vos coram hominibus; Deus autem novit corda vestra, quia, quod hominibus altum est, abominatio est ante Deum.
LUKE|16|16|Lex et Prophetae usque ad Ioannem; ex tunc regnum Dei evangelizatur, et omnis in illud vim facit.
LUKE|16|17|Facilius est autem caelum et terram praeterire, quam de Lege unum apicem cadere.
LUKE|16|18|Omnis, qui dimittit uxorem suam et ducit alteram, moechatur; et, qui dimissam a viro ducit, moechatur.
LUKE|16|19|Homo quidam erat dives et induebatur purpura et bysso et epulabatur cotidie splendide.
LUKE|16|20|Quidam autem pauper nomine Lazarus iacebat ad ianuam eius ulceribus plenus
LUKE|16|21|et cupiens saturari de his, quae cadebant de mensa divitis; sed et canes veniebant et lingebant ulcera eius.
LUKE|16|22|Factum est autem ut moreretur pauper et portaretur ab angelis in sinum Abrahae; mortuus est autem et dives et sepultus est.
LUKE|16|23|Et in inferno elevans oculos suos, cum esset in tormentis, videbat Abraham a longe et Lazarum in sinu eius.
LUKE|16|24|Et ipse clamans dixit: "Pater Abraham, miserere mei et mitte Lazarum, ut intingat extremum digiti sui in aquam, ut refrigeret linguam meam, quia crucior in hac flamma".
LUKE|16|25|At dixit Abraham: "Fili, recordare quia recepisti bona tua in vita tua, et Lazarus similiter mala; nunc autem hic consolatur, tu vero cruciaris.
LUKE|16|26|Et in his omnibus inter nos et vos chaos magnum firmatum est, ut hi, qui volunt hinc transire ad vos, non possint, neque inde ad nos transmeare".
LUKE|16|27|Et ait: "Rogo ergo te, Pater, ut mittas eum in domum patris mei
LUKE|16|28|- habeo enim quinque fratres - ut testetur illis, ne et ipsi veniant in locum hunc tormentorum".
LUKE|16|29|Ait autem Abraham: "Habent Moysen et Prophetas; audiant illos".
LUKE|16|30|At ille dixit: "Non, pater Abraham, sed si quis ex mortuis ierit ad eos, paenitentiam agent".
LUKE|16|31|Ait autem illi: "Si Moysen et Prophetas non audiunt, neque si quis ex mortuis resurrexerit, credent" ".
LUKE|17|1|Et ad discipulos suos ait: " Impossibile est ut non ve niant scandala; vae autem illi, per quem veniunt!
LUKE|17|2|Utilius est illi, si lapis molaris imponatur circa collum eius et proiciatur in mare, quam ut scandalizet unum de pusillis istis.
LUKE|17|3|Attendite vobis!Si peccaverit frater tuus, increpa illum et, si paenitentiam egerit, dimitte illi;
LUKE|17|4|et si septies in die peccaverit in te et septies conversus fuerit ad te dicens: "Paenitet me", dimittes illi ".
LUKE|17|5|Et dixerunt apostoli Domino: " Adauge nobis fidem! ".
LUKE|17|6|Dixit autem Dominus: " Si haberetis fidem sicut granum sinapis, diceretis huic arbori moro: "Eradicare et transplantare in mare", et oboediret vobis.
LUKE|17|7|Quis autem vestrum habens servum arantem aut pascentem, qui regresso de agro dicet illi: "Statim transi, recumbe",
LUKE|17|8|et non dicet ei: "Para, quod cenem, et praecinge te et ministra mihi, donec manducem et bibam, et post haec tu manducabis et bibes"?
LUKE|17|9|Numquid gratiam habet servo illi, quia fecit, quae praecepta sunt?
LUKE|17|10|Sic et vos, cum feceritis omnia, quae praecepta sunt vobis, dicite: Servi inutiles sumus; quod debuimus facere, fecimus" ".
LUKE|17|11|Et factum est, dum iret in Ierusalem, et ipse transibat per mediam Samariam et Galilaeam.
LUKE|17|12|Et cum ingrederetur quoddam castellum, occurrerunt ei decem viri leprosi, qui steterunt a longe
LUKE|17|13|et levaverunt vocem dicentes: " Iesu praeceptor, miserere nostri! ".
LUKE|17|14|Quos ut vidit, dixit: " Ite, ostendite vos sacerdotibus ". Et factum est, dum irent, mundati sunt.
LUKE|17|15|Unus autem ex illis, ut vidit quia sanatus est, regressus est cum magna voce magnificans Deum
LUKE|17|16|et cecidit in faciem ante pedes eius gratias agens ei; et hic erat Samaritanus.
LUKE|17|17|Respondens autem Iesus dixit: " Nonne decem mundati sunt? Et novem ubi sunt?
LUKE|17|18|Non sunt inventi qui redirent, ut darent gloriam Deo, nisi hic alienigena? ".
LUKE|17|19|Et ait illi: " Surge, vade; fides tua te salvum fecit ".
LUKE|17|20|Interrogatus autem a pharisaeis: " Quando venit regnum Dei? ", respondit eis et dixit: " Non venit regnum Dei cum observatione,
LUKE|17|21|neque dicent: "Ecce hic" aut: "Illic"; ecce enim regnum Dei intra vos est ".
LUKE|17|22|Et ait ad discipulos: " Venient dies, quando desideretis videre unum diem Filii hominis et non videbitis.
LUKE|17|23|Et dicent vobis: "Ecce hic", "Ecce illic"; nolite ire neque sectemini.
LUKE|17|24|Nam sicut fulgur coruscans de sub caelo in ea, quae sub caelo sunt, fulget, ita erit Filius hominis in die sua.
LUKE|17|25|Primum autem oportet illum multa pati et reprobari a generatione hac.
LUKE|17|26|Et sicut factum est in diebus Noe, ita erit et in diebus Filii hominis:
LUKE|17|27|edebant, bibebant, uxores ducebant, dabantur ad nuptias, usque in diem, qua intravit Noe in arcam, et venit diluvium et perdidit omnes.
LUKE|17|28|Similiter sicut factum est in diebus Lot: edebant, bibebant, emebant, vendebant, plantabant, aedificabant;
LUKE|17|29|qua die autem exiit Lot a Sodomis, pluit ignem et sulphur de caelo et omnes perdidit.
LUKE|17|30|Secundum haec erit, qua die Filius hominis revelabitur.
LUKE|17|31|In illa die, qui fuerit in tecto, et vasa eius in domo, ne descendat tollere illa; et, qui in agro, similiter non redeat retro.
LUKE|17|32|Memores estote uxoris Lot.
LUKE|17|33|Quicumque quaesierit animam suam salvam facere, perdet illam; et, quicumque perdiderit illam, vivificabit eam.
LUKE|17|34|Dico vobis: Illa nocte erunt duo in lecto uno:unus assumetur, et alter relinquetur;
LUKE|17|35|duae erunt molentes in unum: una assumetur, et altera relinquetur ". 36) 37 Respondentes dicunt illi: " Ubi, Domine? ". Qui dixit eis: " Ubicumque fuerit corpus, illuc congregabuntur et aquilae ".
LUKE|18|1|Dicebat autem parabolam ad illos, quoniam oportet semper orare et non deficere,
LUKE|18|2|dicens: " Iudex quidam erat in quadam civitate, qui Deum non timebat et hominem non reverebatur.
LUKE|18|3|Vidua autem erat in civitate illa et veniebat ad eum dicens: "Vindica me de adversario meo".
LUKE|18|4|Et nolebat per multum tempus; post haec autem dixit intra se: "Etsi Deum non timeo nec hominem revereor,
LUKE|18|5|tamen quia molesta est mihi haec vidua, vindicabo illam, ne in novissimo veniens suggillet me" ".
LUKE|18|6|Ait autem Dominus: " Audite quid iudex iniquitatis dicit;
LUKE|18|7|Deus autem non faciet vindictam electorum suorum clamantium ad se die ac nocte, et patientiam habebit in illis?
LUKE|18|8|Dico vobis: Cito faciet vindictam illorum. Verumtamen Filius hominis veniens, putas, inveniet fidem in terra? ".
LUKE|18|9|Dixit autem et ad quosdam, qui in se confidebant tamquam iusti et aspernabantur ceteros, parabolam istam:
LUKE|18|10|" Duo homines ascenderunt in templum, ut orarent: unus pharisaeus et alter publicanus.
LUKE|18|11|Pharisaeus stans haec apud se orabat: "Deus, gratias ago tibi, quia non sum sicut ceteri hominum, raptores, iniusti, adulteri, velut etiam hic publicanus;
LUKE|18|12|ieiuno bis in sabbato, decimas do omnium, quae possideo".
LUKE|18|13|Et publicanus a longe stans nolebat nec oculos ad caelum levare, sed percutiebat pectus suum dicens: "Deus, propitius esto mihi peccatori".
LUKE|18|14|Dico vobis: Descendit hic iustificatus in domum suam ab illo. Quia omnis, qui se exaltat, humiliabitur; et, qui se humiliat, exaltabitur ".
LUKE|18|15|Afferebant autem ad illum et infantes, ut eos tangeret; quod cum viderent, discipuli increpabant illos.
LUKE|18|16|Iesus autem convocans illos dixit: " Sinite pueros venire ad me et nolite eos vetare; talium est enim regnum Dei.
LUKE|18|17|Amen dico vobis: Quicumque non acceperit regnum Dei sicut puer, non intrabit in illud ".
LUKE|18|18|Et interrogavit eum quidam princeps dicens: " Magister bone, quid faciens vitam aeternam possidebo? ".
LUKE|18|19|Dixit autem ei Iesus: " Quid me dicis bonum? Nemo bonus nisi solus Deus.
LUKE|18|20|Mandata nosti: non moechaberis, non occides, non furtum facies, non falsum testimonium dices, honora patrem tuum et matrem ".
LUKE|18|21|Qui ait: " Haec omnia custodivi a iuventute ".
LUKE|18|22|Quo audito, Iesus ait ei: " Adhuc unum tibi deest: omnia, quaecumque habes, vende et da pauperibus et habebis thesaurum in caelo: et veni, sequere me ".
LUKE|18|23|His ille auditis, contristatus est, quia dives erat valde.
LUKE|18|24|Videns autem illum Iesus tristem factum dixit: " Quam difficile, qui pecunias habent, in regnum Dei intrant.
LUKE|18|25|Facilius est enim camelum per foramen acus transire, quam divitem intrare in regnum Dei ".
LUKE|18|26|Et dixerunt, qui audiebant: " Et quis potest salvus fieri? ".
LUKE|18|27|Ait autem illis: " Quae impossibilia sunt apud homi nes, possibilia sunt apud Deum ".
LUKE|18|28|Ait autem Petrus: " Ecce nos dimisimus nostra et secuti sumus te ".
LUKE|18|29|Qui dixit eis: " Amen dico vobis: Nemo est, qui reliquit domum aut uxorem aut fratres aut parentes aut filios propter regnum Dei,
LUKE|18|30|et non recipiat multo plura in hoc tempore et in saeculo venturo vitam aeternam ".
LUKE|18|31|Assumpsit autem Duodecim et ait illis: " Ecce ascendimus Ierusalem, et consummabuntur omnia, quae scripta sunt per Prophetas de Filio hominis:
LUKE|18|32|tradetur enim gentibus et illudetur et contumeliis afficietur et conspuetur;
LUKE|18|33|et, postquam flagellaverint, occident eum, et die tertia resurget ".
LUKE|18|34|Et ipsi nihil horum intellexerunt; et erat verbum istud absconditum ab eis, et non intellegebant, quae dicebantur.
LUKE|18|35|Factum est autem, cum appropinquaret Iericho, caecus quidam sedebat secus viam mendicans.
LUKE|18|36|Et cum audiret turbam praetereuntem, interrogabat quid hoc esset.
LUKE|18|37|Dixerunt autem ei: " Iesus Nazarenus transit ".
LUKE|18|38|Et clamavit dicens: " Iesu, fili David, miserere mei! ".
LUKE|18|39|Et qui praeibant, increpabant eum, ut taceret; ipse vero multo magis clamabat: " Fili David, miserere mei! ".
LUKE|18|40|Stans autem Iesus iussit illum adduci ad se. Et cum appropinquasset, interrogavit illum:
LUKE|18|41|" Quid tibi vis faciam? ". At ille dixit: " Domine, ut videam ".
LUKE|18|42|Et Iesus dixit illi: " Respice! Fides tua te salvum fecit ". 43 Et confestim vidit et sequebatur illum magnificans Deum. Et omnis plebs, ut vidit, dedit laudem Deo.
LUKE|19|1|Et ingressus perambulabat Iericho.
LUKE|19|2|Et ecce vir nomine Zacchaeus, et hic erat princeps publicanorum et ipse dives.
LUKE|19|3|Et quaerebat videre Iesum, quis esset, et non poterat prae turba, quia statura pusillus erat.
LUKE|19|4|Et praecurrens ascendit in arborem sycomorum, ut videret illum, quia inde erat transiturus.
LUKE|19|5|Et cum venisset ad locum, suspiciens Iesus dixit ad eum: " Zacchaee, festinans descende, nam hodie in domo tua oportet me manere ".
LUKE|19|6|Et festinans descendit et excepit illum gaudens.
LUKE|19|7|Et cum viderent, omnes murmurabant dicentes: " Ad hominem peccatorem divertit! ".
LUKE|19|8|Stans autem Zacchaeus dixit ad Dominum: " Ecce dimidium bonorum meorum, Domine, do pauperibus et, si quid aliquem defraudavi, reddo quadruplum ".
LUKE|19|9|Ait autem Iesus ad eum: " Hodie salus domui huic facta est, eo quod et ipse filius sit Abrahae;
LUKE|19|10|venit enim Filius hominis quaerere et salvum facere, quod perierat ".
LUKE|19|11|Haec autem illis audientibus, adiciens dixit parabolam, eo quod esset prope Ierusalem, et illi existimarent quod confestim regnum Dei manifestaretur.
LUKE|19|12|Dixit ergo: " Homo quidam nobilis abiit in regionem longinquam accipere sibi regnum et reverti.
LUKE|19|13|Vocatis autem decem servis suis, dedit illis decem minas et ait ad illos: "Negotiamini, dum venio".
LUKE|19|14|Cives autem eius oderant illum et miserunt legationem post illum dicentes: "Nolumus hunc regnare super nos!".
LUKE|19|15|Et factum est ut rediret, accepto regno, et iussit ad se vocari servos illos, quibus dedit pecuniam, ut sciret quantum negotiati essent.
LUKE|19|16|Venit autem primus dicens: "Domine, mina tua decem minas acquisivit".
LUKE|19|17|Et ait illi: "Euge, bone serve; quia in modico fidelis fuisti, esto potestatem habens supra decem civitates".
LUKE|19|18|Et alter venit dicens: "Mina tua, domine, fecit quinque minas".
LUKE|19|19|Et huic ait: "Et tu esto supra quinque civitates".
LUKE|19|20|Et alter venit dicens: "Domine, ecce mina tua, quam habui repositam in sudario;
LUKE|19|21|timui enim te, quia homo austerus es: tollis, quod non posuisti, et metis, quod non seminasti".
LUKE|19|22|Dicit ei: "De ore tuo te iudico, serve nequam! Sciebas quod ego austerus homo sum, tollens quod non posui et metens quod non seminavi?
LUKE|19|23|Et quare non dedisti pecuniam meam ad mensam? Et ego veniens cum usuris utique exegissem illud".
LUKE|19|24|Et adstantibus dixit: "Auferte ab illo minam et date illi, qui decem minas habet".
LUKE|19|25|Et dixerunt ei: "Domine, habet decem minas!".
LUKE|19|26|Dico vobis: "Omni habenti dabitur; ab eo autem, qui non habet, et, quod habet, auferetur.
LUKE|19|27|Verumtamen inimicos meos illos, qui noluerunt me regnare super se, adducite huc et interficite ante me! ".
LUKE|19|28|Et his dictis, praecedebat ascendens Hierosolymam.
LUKE|19|29|Et factum est, cum appropinquasset ad Bethfage et Bethaniam, ad montem, qui vocatur Oliveti, misit duos discipulos
LUKE|19|30|dicens: " Ite in castellum, quod contra est, in quod introeuntes invenietis pullum asinae alligatum, cui nemo umquam hominum sedit; solvite illum et adducite.
LUKE|19|31|Et si quis vos interrogaverit: "Quare solvitis?", sic dicetis: "Dominus eum necessarium habet" ".
LUKE|19|32|Abierunt autem, qui missi erant, et invenerunt, sicut dixit illis.
LUKE|19|33|Solventibus autem illis pullum, dixerunt domini eius ad illos: " Quid solvitis pullum? ".
LUKE|19|34|At illi dixerunt: " Dominus eum necessarium habet ".
LUKE|19|35|Et duxerunt illum ad Iesum; et iactantes vestimenta sua supra pullum, imposuerunt Iesum.
LUKE|19|36|Eunte autem illo, substernebant vestimenta sua in via.
LUKE|19|37|Et cum appropinquaret iam ad descensum montis Oliveti, coeperunt omnis multitudo discipulorum gaudentes laudare Deum voce magna super omnibus, quas viderant, virtutibus
LUKE|19|38|dicentes: Benedictus, qui venit rex in nomine Domini!Pax in caelo, et gloria in excelsis! ".
LUKE|19|39|Et quidam pharisaeorum de turbis dixerunt ad illum: " Magister, increpa discipulos tuos! ".
LUKE|19|40|Et respondens dixit: " Dico vobis: Si hi tacuerint, lapides clamabunt!.
LUKE|19|41|Et ut appropinquavit, videns civitatem flevit super illam
LUKE|19|42|dicens: " Si cognovisses et tu in hac die, quae ad pacem tibi! Nunc autem abscondita sunt ab oculis tuis.
LUKE|19|43|Quia venient dies in te, et circumdabunt te inimici tui vallo et obsidebunt te et coangustabunt te undique
LUKE|19|44|et ad terram prosternent te et filios tuos, qui in te sunt, et non relinquent in te lapidem super lapidem, eo quod non cognoveris tempus visitationis tuae ".
LUKE|19|45|Et ingressus in templum, coepit eicere vendentes
LUKE|19|46|dicens illis: " Scriptum est: "Et erit domus mea domus orationis". Vos autem fecistis illam speluncam latronum ".
LUKE|19|47|Et erat docens cotidie in templo. Principes autem sacerdotum et scribae et principes plebis quaerebant illum perdere
LUKE|19|48|et non inveniebant quid facerent; omnis enim populus suspensus erat audiens illum.
LUKE|20|1|Et factum est in una dierum, docente illo populum in tem plo et evangelizante, supervenerunt principes sacerdotum et scribae cum senioribus
LUKE|20|2|et aiunt dicentes ad illum: " Dic nobis: In qua potestate haec facis, aut quis est qui dedit tibi hanc potestatem? ".
LUKE|20|3|Respondens autem dixit ad illos: " Interrogabo vos et ego verbum; et dicite mihi:
LUKE|20|4|Baptismum Ioannis de caelo erat an ex hominibus? ".
LUKE|20|5|At illi cogitabant inter se dicentes: " Si dixerimus: "De caelo", dicet: Quare non credidistis illi?;
LUKE|20|6|si autem dixerimus: "Ex hominibus", plebs universa lapidabit nos; certi sunt enim Ioannem prophetam esse ".
LUKE|20|7|Et responderunt se nescire unde esset.
LUKE|20|8|Et Iesus ait illis: " Neque ego dico vobis in qua potestate haec facio.
LUKE|20|9|Coepit autem dicere ad plebem parabolam hanc: " Homo plantavit vineam et locavit eam colonis et ipse peregre fuit multis temporibus.
LUKE|20|10|Et in tempore misit ad cultores servum, ut de fructu vineae darent illi; cultores autem caesum dimiserunt eum inanem.
LUKE|20|11|Et addidit alterum servum mittere; illi autem hunc quoque caedentes et afficientes contumelia dimiserunt inanem.
LUKE|20|12|Et addidit tertium mittere; qui et illum vulnerantes eiecerunt.
LUKE|20|13|Dixit autem dominus vineae: "Quid faciam? Mittam filium meum dilectum; forsitan hunc verebuntur".
LUKE|20|14|Quem cum vidissent coloni, cogitaverunt inter se dicentes: "Hic est heres. Occidamus illum, ut nostra fiat hereditas".
LUKE|20|15|Et eiectum illum extra vineam occiderunt. Quid ergo faciet illis dominus vineae?
LUKE|20|16|Veniet et perdet colonos istos et dabit vineam aliis ".Quo audito, dixerunt: " Absit! ".
LUKE|20|17|Ille autem aspiciens eos ait: " Quid est ergo hoc, quod scriptum est:Lapidem quem reprobaverunt aedificantes,hic factus est in caput anguli"?
LUKE|20|18|Omnis, qui ceciderit supra illum lapidem, conquassabitur; supra quem autem ceciderit, comminuet illum ".
LUKE|20|19|Et quaerebant scribae et principes sacerdotum mittere in illum manus in illa hora et timuerunt populum; cognoverunt enim quod ad ipsos dixerit similitudinem istam.
LUKE|20|20|Et observantes miserunt insidiatores, qui se iustos simularent, ut caperent eum in sermone, et sic traderent illum principatui et potestati praesidis.
LUKE|20|21|Et interrogaverunt illum dicentes: " Magister, scimus quia recte dicis et doces et non accipis personam, sed in veritate viam Dei doces.
LUKE|20|22|Licet nobis dare tributum Caesari an non? ".
LUKE|20|23|Considerans autem dolum illorum dixit ad eos:
LUKE|20|24|" Ostendite mihi denarium. Cuius habet imaginem et inscriptionem? ".
LUKE|20|25|At illi dixerunt: " Caesaris ". Et ait illis: " Reddite ergo, quae Caesaris sunt, Caesari et, quae Dei sunt, Deo ".
LUKE|20|26|Et non potuerunt verbum eius reprehendere coram plebe et mirati in responso eius tacuerunt.
LUKE|20|27|Accesserunt autem quidam sadducaeorum, qui negant esse resurrectionem, et interrogaverunt eum
LUKE|20|28|dicentes: " Magister, Moyses scripsit nobis, si frater alicuius mortuus fuerit habens uxorem et hic sine filiis fuerit, ut accipiat eam frater eius uxorem et suscitet semen fratri suo.
LUKE|20|29|Septem ergo fratres erant: et primus accepit uxorem et mortuus est sine filiis;
LUKE|20|30|et sequens
LUKE|20|31|et tertius accepit illam, similiter autem et septem non reliquerunt filios et mortui sunt.
LUKE|20|32|Novissima mortua est et mulier.
LUKE|20|33|Mulier ergo in resurrectione cuius eorum erit uxor? Si quidem septem habuerunt eam uxorem ".
LUKE|20|34|Et ait illis Iesus: " Filii saeculi huius nubunt et traduntur ad nuptias;
LUKE|20|35|illi autem, qui digni habentur saeculo illo et resurrectione ex mortuis, neque nubunt neque ducunt uxores.
LUKE|20|36|Neque enim ultra mori possunt: aequales enim angelis sunt et filii sunt Dei, cum sint filii resurrectionis.
LUKE|20|37|Quia vero resurgant mortui, et Moyses ostendit secus rubum, sicut dicit: "Dominum Deum Abraham et Deum Isaac et Deum Iacob".
LUKE|20|38|Deus autem non est mortuorum sed vivorum: omnes enim vivunt ei ".
LUKE|20|39|Respondentes autem quidam scribarum dixerunt: " Magister, bene dixisti.
LUKE|20|40|Et amplius non audebant eum quidquam interrogare.
LUKE|20|41|Dixit autem ad illos: " Quomodo dicunt Christum filium David esse?
LUKE|20|42|Ipse enim David dicit in libro Psalmorum:Dixit Dominus Domino meo: Sede a dextris meis,
LUKE|20|43|donec ponam inimicos tuos scabellum pedum tuorum".
LUKE|20|44|David ergo Dominum illum vocat; et quomodo filius eius est? ".
LUKE|20|45|Audiente autem omni populo, dixit discipulis suis:
LUKE|20|46|" Attendite a scribis, qui volunt ambulare in stolis et amant salutationes in foro et primas cathedras in synagogis et primos discubitus in conviviis,
LUKE|20|47|qui devorant domos viduarum et simulant longam orationem. Hi accipient damnationem maiorem ".
LUKE|21|1|Respiciens autem vidit eos, qui mittebant munera sua in gazophylacium, divites.
LUKE|21|2|Vidit autem quandam viduam pauperculam mittentem illuc minuta duo
LUKE|21|3|et dixit: " Vere dico vobis: Vidua haec pauper plus quam omnes misit.
LUKE|21|4|Nam omnes hi ex abundantia sua miserunt in munera; haec autem ex inopia sua omnem victum suum, quem habebat, misit ".
LUKE|21|5|Et quibusdam dicentibus de templo, quod lapidibus bonis et donis ornatum, esset dixit:
LUKE|21|6|" Haec quae videtis, venient dies, in quibus non relinquetur lapis super lapidem, qui non destruatur ".
LUKE|21|7|Interrogaverunt autem illum dicentes: " Praeceptor, quando ergo haec erunt, et quod signum, cum fieri incipient? ".
LUKE|21|8|Qui dixit: " Videte, ne seducamini. Multi enim venient in nomine meo dicentes: "Ego sum" et: "Tempus appropinquavit". Nolite ergo ire post illos.
LUKE|21|9|Cum autem audieritis proelia et seditiones, nolite terreri; oportet enim primum haec fieri, sed non statim finis ".
LUKE|21|10|Tunc dicebat illis: " Surget gens contra gentem, et regnum adversus regnum;
LUKE|21|11|et terrae motus magni et per loca fames et pestilentiae erunt, terroresque et de caelo signa magna erunt.
LUKE|21|12|Sed ante haec omnia inicient vobis manus suas et persequentur tradentes in synagogas et custodias, et trahemini ad reges et praesides propter nomen meum;
LUKE|21|13|continget autem vobis in testimonium.
LUKE|21|14|Ponite ergo in cordibus vestris non praemeditari quemadmodum respondeatis;
LUKE|21|15|ego enim dabo vobis os et sapientiam, cui non poterunt resistere vel contradicere omnes adversarii vestri.
LUKE|21|16|Trademini autem et a parentibus et fratribus et cognatis et amicis, et morte afficient ex vobis,
LUKE|21|17|et eritis odio omnibus propter nomen meum.
LUKE|21|18|Et capillus de capite vestro non peribit.
LUKE|21|19|In patientia vestra possidebitis animas vestras.
LUKE|21|20|Cum autem videritis circumdari ab exercitu Ierusalem, tunc scitote quia appropinquavit desolatio eius.
LUKE|21|21|Tunc, qui in Iudaea sunt, fugiant in montes; et, qui in medio eius, discedant; et, qui in regionibus, non intrent in eam.
LUKE|21|22|Quia dies ultionis hi sunt, ut impleantur omnia, quae scripta sunt.
LUKE|21|23|Vae autem praegnantibus et nutrientibus in illis diebus! Erit enim pressura magna super terram et ira populo huic,
LUKE|21|24|et cadent in ore gladii et captivi ducentur in omnes gentes, et Ierusalem calcabitur a gentibus, donec impleantur tempora nationum.
LUKE|21|25|Et erunt signa in sole et luna et stellis, et super terram pressura gentium prae confusione sonitus maris et fluctuum,
LUKE|21|26|arescentibus hominibus prae timore et exspectatione eorum, quae supervenient orbi, nam virtutes caelorum movebuntur.
LUKE|21|27|Et tunc videbunt Filium hominis venientem in nube cum potestate et gloria magna.
LUKE|21|28|His autem fieri incipientibus, respicite et levate capita vestra, quoniam appropinquat redemptio vestra ".
LUKE|21|29|Et dixit illis similitudinem: " Videte ficulneam et omnes arbores:
LUKE|21|30|cum iam germinaverint, videntes vosmetipsi scitis quia iam prope est aestas.
LUKE|21|31|Ita et vos, cum videritis haec fieri, scitote quoniam prope est regnum Dei.
LUKE|21|32|Amen dico vobis: Non praeteribit generatio haec, donec omnia fiant.
LUKE|21|33|Caelum et terra transibunt, verba autem mea non transibunt.
LUKE|21|34|Attendite autem vobis, ne forte graventur corda vestra in crapula et ebrietate et curis huius vitae, et superveniat in vos repentina dies illa;
LUKE|21|35|tamquam laqueus enim superveniet in omnes, qui sedent super faciem omnis terrae.
LUKE|21|36|Vigilate itaque omni tempore orantes, ut possitis fugere ista omnia, quae futura sunt, et stare ante Filium hominis ".
LUKE|21|37|Erat autem diebus docens in templo, noctibus vero exiens morabatur in monte, qui vocatur Oliveti.
LUKE|21|38|Et omnis populus manicabat ad eum in templo audire eum.
LUKE|22|1|Appropinquabat autem dies festus Azymorum, qui dici tur Pascha.
LUKE|22|2|Et quaerebant principes sacerdotum et scribae quomodo eum interficerent; timebant vero plebem.
LUKE|22|3|Intravit autem Satanas in Iudam, qui cognominabatur Iscarioth, unum de Duodecim;
LUKE|22|4|et abiit et locutus est cum principibus sacerdotum et magistratibus, quemadmodum illum traderet eis.
LUKE|22|5|Et gavisi sunt et pacti sunt pecuniam illi dare.
LUKE|22|6|Et spopondit et quaerebat opportunitatem, ut eis traderet illum sine turba.
LUKE|22|7|Venit autem dies Azymorum, in qua necesse erat occidi Pascha.
LUKE|22|8|Et misit Petrum et Ioannem dicens: " Euntes parate nobis Pascha, ut manducemus ".
LUKE|22|9|At illi dixerunt ei: "Ubi vis paremus? ".
LUKE|22|10|Et dixit ad eos: " Ecce, introeuntibus vobis in civitatem, occurret vobis homo amphoram aquae portans; sequimini eum in domum, in quam intrat.
LUKE|22|11|Et dicetis patri familias domus: "Dicit tibi Magister: Ubi est deversorium, ubi Pascha cum discipulis meis manducem?".
LUKE|22|12|Ipse vobis ostendet cenaculum magnum stratum; ibi parate ".
LUKE|22|13|Euntes autem invenerunt, sicut dixit illis, et paraverunt Pascha.
LUKE|22|14|Et cum facta esset hora, discubuit, et apostoli cum eo.
LUKE|22|15|Et ait illis: " Desiderio desideravi hoc Pascha manducare vobiscum, antequam patiar.
LUKE|22|16|Dico enim vobis: Non manducabo illud, donec impleatur in regno Dei ".
LUKE|22|17|Et accepto calice, gratias egit et dixit: " Accipite hoc et dividite inter vos.
LUKE|22|18|Dico enim vobis: Non bibam amodo de generatione vitis, donec regnum Dei veniat ".
LUKE|22|19|Et accepto pane, gratias egit et fregit et dedit eis dicens: " Hoc est corpus meum, quod pro vobis datur. Hoc facite in meam commemorationem ".
LUKE|22|20|Similiter et calicem, postquam cenavit, dicens: " Hic calix novum testamentum est in sanguine meo, qui pro vobis funditur.
LUKE|22|21|Verumtamen ecce manus tradentis me mecum est in mensa;
LUKE|22|22|et quidem Filius hominis, secundum quod definitum est, vadit; verumtamen vae illi homini, per quem traditur! ".
LUKE|22|23|Et ipsi coeperunt quaerere inter se, quis esset ex eis, qui hoc facturus esset.
LUKE|22|24|Facta est autem et contentio inter eos, quis eorum videretur esse maior.
LUKE|22|25|Dixit autem eis: " Reges gentium dominantur eorum; et, qui potestatem habent super eos, benefici vocantur.
LUKE|22|26|Vos autem non sic, sed qui maior est in vobis, fiat sicut iunior; et, qui praecessor est, sicut ministrator.
LUKE|22|27|Nam quis maior est: qui recumbit, an qui ministrat? Nonne qui recumbit? Ego autem in medio vestrum sum, sicut qui ministrat.
LUKE|22|28|Vos autem estis, qui permansistis mecum in tentationibus meis;
LUKE|22|29|et ego dispono vobis, sicut disposuit mihi Pater meus regnum,
LUKE|22|30|ut edatis et bibatis super mensam meam in regno meo et sedeatis super thronos iudicantes duodecim tribus Israel.
LUKE|22|31|Simon, Simon, ecce Satanas expetivit vos, ut cribraret sicut triticum;
LUKE|22|32|ego autem rogavi pro te, ut non deficiat fides tua. Et tu, aliquando conversus, confirma fratres tuos ".
LUKE|22|33|Qui dixit ei: " Domine, tecum paratus sum et in carcerem et in mortem ire ".
LUKE|22|34|Et ille dixit: " Dico tibi, Petre, non cantabit hodie gallus, donec ter abneges nosse me ".
LUKE|22|35|Et dixit eis: " Quando misi vos sine sacculo et pera et calceamentis, numquid aliquid defuit vobis? ". At illi dixerunt: " Nihil ".
LUKE|22|36|Dixit ergo eis: " Sed nunc, qui habet sacculum, tollat, similiter et peram; et, qui non habet, vendat tunicam suam et emat gladium.
LUKE|22|37|Dico enim vobis: Hoc, quod scriptum est, oportet impleri in me, illud: Cum iniustis deputatus est". Etenim ea, quae sunt de me, adimpletionem habent ".
LUKE|22|38|At illi dixerunt: " Domine, ecce gladii duo hic ". At ille dixit eis: " Satis est ".
LUKE|22|39|Et egressus ibat secundum consuetudinem in montem Olivarum; secuti sunt autem illum et discipuli.
LUKE|22|40|Et cum pervenisset ad locum, dixit illis: " Orate, ne intretis in tentationem ".
LUKE|22|41|Et ipse avulsus est ab eis, quantum iactus est lapidis, et, positis genibus, orabat
LUKE|22|42|dicens: " Pater, si vis, transfer calicem istum a me; verumtamen non mea voluntas sed tua fiat ".
LUKE|22|43|Apparuit autem illi angelus de caelo confortans eum. Et factus in agonia prolixius orabat.
LUKE|22|44|Et factus est sudor eius sicut guttae sanguinis decurrentis in terram.
LUKE|22|45|Et cum surrexisset ab oratione et venisset ad discipulos, invenit eos dormientes prae tristitia
LUKE|22|46|et ait illis: " Quid dormitis? Surgite; orate, ne intretis in tentationem ".
LUKE|22|47|Adhuc eo loquente, ecce turba; et, qui vocabatur Iudas, unus de Duodecim, antecedebat eos et appropinquavit Iesu, ut oscularetur eum.
LUKE|22|48|Iesus autem dixit ei: " Iuda, osculo Filium hominis tradis? ".
LUKE|22|49|Videntes autem hi, qui circa ipsum erant, quod futurum erat, dixerunt: Domine, si percutimus in gladio? ".
LUKE|22|50|Et percussit unus ex illis servum principis sacerdotum et amputavit auriculam eius dextram.
LUKE|22|51|Respondens autem Iesus ait: " Sinite usque huc! ". Et cum tetigisset auriculam eius, sanavit eum.
LUKE|22|52|Dixit autem Iesus ad eos, qui venerant ad se principes sacerdotum et magistratus templi et seniores: " Quasi ad latronem existis cum gladiis et fustibus?
LUKE|22|53|Cum cotidie vobiscum fuerim in templo, non extendistis manus in me; sed haec est hora vestra et potestas tenebrarum ".
LUKE|22|54|Comprehendentes autem eum, duxerunt et introduxerunt in domum principis sacerdotum. Petrus vero sequebatur a longe.
LUKE|22|55|Accenso autem igni in medio atrio et circumsedentibus illis, sedebat Petrus in medio eorum.
LUKE|22|56|Quem cum vidisset ancilla quaedam sedentem ad lumen et eum fuisset intuita, dixit:
LUKE|22|57|" Et hic cum illo erat! ". At ille negavit eum dicens:
LUKE|22|58|" Mulier, non novi illum! ". Et post pusillum alius videns eum dixit: " Et tu de illis es! ". Petrus vero ait: " O homo, non sum! ".
LUKE|22|59|Et intervallo facto quasi horae unius, alius quidam affirmabat dicens: Vere et hic cum illo erat, nam et Galilaeus est! ".
LUKE|22|60|Et ait Petrus: " Homo, nescio quid dicis! ". Et continuo adhuc illo loquente cantavit gallus.
LUKE|22|61|Et conversus Dominus respexit Petrum; et recordatus est Petrus verbi Domini, sicut dixit ei: " Priusquam gallus cantet hodie, ter me negabis ".
LUKE|22|62|Et egressus foras flevit amare.
LUKE|22|63|Et viri, qui tenebant illum, illudebant ei caedentes;
LUKE|22|64|et velaverunt eum et interrogabant eum dicentes: " Prophetiza: Quis est, qui te percussit? ".
LUKE|22|65|Et alia multa blasphemantes dicebant in eum.
LUKE|22|66|Et ut factus est dies, convenerunt seniores plebis et principes sacerdotum et scribae et duxerunt illum in concilium suum
LUKE|22|67|dicentes: " Si tu es Christus, dic nobis ". Et ait illis: " Si vobis dixero, non credetis;
LUKE|22|68|si autem interrogavero, non respondebitis mihi.
LUKE|22|69|Ex hoc autem erit Filius hominis sedens a dextris virtutis Dei ".
LUKE|22|70|Dixerunt autem omnes: " Tu ergo es Filius Dei? ". Qui ait ad illos: " Vos dicitis quia ego sum ".
LUKE|22|71|At illi dixerunt: " Quid adhuc desideramus testimonium? Ipsi enim audivimus de ore eius! ".
LUKE|23|1|Et surgens omnis multitudo eorum duxerunt illum ad Pi latum.
LUKE|23|2|Coeperunt autem accusare illum dicentes: " Hunc invenimus subvertentem gentem nostram et prohibentem tributa dare Caesari et dicentem se Christum regem esse ".
LUKE|23|3|Pilatus autem interrogavit eum dicens: " Tu es rex Iudaeorum? ". At ille respondens ait: " Tu dicis ".
LUKE|23|4|Ait autem Pilatus ad principes sacerdotum et turbas: " Nihil invenio causae in hoc homine ".
LUKE|23|5|At illi invalescebant dicentes: " Commovet populum docens per universam Iudaeam et in cipiens a Galilaea usque huc! ".
LUKE|23|6|Pilatus autem audiens interrogavit si homo Galilaeus esset;
LUKE|23|7|et ut cognovit quod de Herodis potestate esset, remisit eum ad Herodem, qui et ipse Hierosolymis erat illis diebus.
LUKE|23|8|Herodes autem, viso Iesu, gavisus est valde; erat enim cupiens ex multo tempore videre eum, eo quod audiret de illo et sperabat signum aliquod videre ab eo fieri.
LUKE|23|9|Interrogabat autem illum multis sermonibus; at ipse nihil illi respondebat.
LUKE|23|10|Stabant etiam principes sacerdotum et scribae constanter accusantes eum.
LUKE|23|11|Sprevit autem illum Herodes cum exercitu suo et illusit indutum veste alba et remisit ad Pilatum.
LUKE|23|12|Facti sunt autem amici inter se Herodes et Pilatus in ipsa die; nam antea inimici erant ad invicem.
LUKE|23|13|Pilatus autem, convocatis principibus sacerdotum et magistratibus et plebe,
LUKE|23|14|dixit ad illos: " Obtulistis mihi hunc hominem quasi avertentem populum, et ecce ego coram vobis interrogans nullam causam inveni in homine isto ex his, in quibus eum accusatis,
LUKE|23|15|sedneque Herodes; remisit enim illum ad nos. Et ecce nihil dignum morte actum est ei.
LUKE|23|16|Emendatum ergo illum dimittam ".
LUKE|23|17|()
LUKE|23|18|Exclamavit autem universa turba dicens: " Tolle hunc et dimitte nobis Barabbam! ",
LUKE|23|19|qui erat propter seditionem quandam factam in civitate et homicidium missus in carcerem.
LUKE|23|20|Iterum autem Pilatus locutus est ad illos volens dimittere Iesum,
LUKE|23|21|at illi succlamabant dicentes: " Crucifige, crucifige illum! ".
LUKE|23|22|Ille autem tertio dixit ad illos: " Quid enim mali fecit iste? Nullam causam mortis invenio in eo; corripiam ergo illum et dimittam ".
LUKE|23|23|At illi instabant vocibus magnis postulantes, ut crucifigeretur, et invalescebant voces eorum.
LUKE|23|24|Et Pilatus adiudicavit fieri petitionem eorum:
LUKE|23|25|dimisit autem eum, qui propter seditionem et homicidium missus fuerat in carcerem, quem petebant; Iesum vero tradidit voluntati eorum.
LUKE|23|26|Et cum abducerent eum, apprehenderunt Simonem quendam Cyrenensem venientem de villa et imposuerunt illi crucem portare post Iesum.
LUKE|23|27|Sequebatur autem illum multa turba populi et mulierum, quae plangebant et lamentabant eum.
LUKE|23|28|Conversus autem ad illas Iesus dixit: " Filiae Ierusalem, nolite flere super me, sed super vos ipsas flete et super filios vestros,
LUKE|23|29|quoniam ecce venient dies, in quibus dicent: "Beatae steriles et ventres, qui non genuerunt, et ubera, quae non lactaverunt!".
LUKE|23|30|Tunc incipient dicere montibus: "Cadite super nos!", et collibus: Operite nos!",
LUKE|23|31|quia si in viridi ligno haec faciunt, in arido quid fiet? ".
LUKE|23|32|Ducebantur autem et alii duo nequam cum eo, ut interficerentur.
LUKE|23|33|Et postquam venerunt in locum, qui vocatur Calvariae, ibi crucifixerunt eum et latrones, unum a dextris et alterum a sinistris.
LUKE|23|34|Iesus autem dicebat: " Pater, dimitte illis, non enim sciunt quid faciunt ".Dividentes vero vestimenta eius miserunt sortes.
LUKE|23|35|Et stabat populus exspectans. Et deridebant illum et principes dicentes: " Alios salvos fecit; se salvum faciat, si hic est Christus Dei electus! ".
LUKE|23|36|Illudebant autem ei et milites accedentes, acetum offerentes illi
LUKE|23|37|et dicentes: " Si tu es rex Iudaeorum, salvum te fac! ".
LUKE|23|38|Erat autem et superscriptio super illum: " Hic est rex Iudaeorum ".
LUKE|23|39|Unus autem de his, qui pendebant, latronibus blasphemabat eum dicens: " Nonne tu es Christus? Salvum fac temetipsum et nos! ".
LUKE|23|40|Respondens autem alter increpabat illum dicens: " Neque tu times Deum, quod in eadem damnatione es?
LUKE|23|41|Et nos quidem iuste, nam digna factis recipimus! Hic vero nihil mali gessit ".
LUKE|23|42|Et dicebat: " Iesu, memento mei, cum veneris in regnum tuum ".
LUKE|23|43|Et dixit illi: " Amen dico tibi: Hodie mecum eris in paradiso ".
LUKE|23|44|Et erat iam fere hora sexta, et tenebrae factae sunt in universa terra usque in horam nonam,
LUKE|23|45|et obscuratus est sol, et velum templi scissum est medium.
LUKE|23|46|Et clamans voce magna Iesus ait: " Pater, in manus tuas commendo spiritum meum "; et haec dicens exspiravit.
LUKE|23|47|Videns autem centurio, quod factum fuerat, glorificavit Deum dicens: " Vere hic homo iustus erat! ".
LUKE|23|48|Et omnis turba eorum, qui simul aderant ad spectaculum istud et videbant, quae fiebant, percutientes pectora sua revertebantur.
LUKE|23|49|Stabant autem omnes noti eius a longe et mulieres, quae secutae erant eum a Galilaea, haec videntes.
LUKE|23|50|Et ecce vir nomine Ioseph, qui erat decurio, vir bonus et iustus
LUKE|23|51|Chic non consenserat consilio et actibus eorum - ab Arimathaea civitate Iudaeorum, qui exspectabat regnum Dei,
LUKE|23|52|hic accessit ad Pilatum et petiit corpus Iesu
LUKE|23|53|et depositum involvit sindone et posuit eum in monumento exciso, in quo nondum quisquam positus fuerat.
LUKE|23|54|Et dies erat Parasceves, et sabbatum illucescebat.
LUKE|23|55|Subsecutae autem mulieres, quae cum ipso venerant de Galilaea, viderunt monumentum et quemadmodum positum erat corpus eius;
LUKE|23|56|et revertentes paraverunt aromata et unguenta et sabbato quidem siluerunt secundum mandatum.
LUKE|24|1|Prima autem sabbatorum, valde diluculo venerunt ad monumentum portantes, quae paraverant, aromata.
LUKE|24|2|Et invenerunt lapidem revolutum a monumento;
LUKE|24|3|et ingressae non invenerunt corpus Domini Iesu.
LUKE|24|4|Et factum est, dum mente haesitarent de isto, ecce duo viri steterunt secus illas in veste fulgenti.
LUKE|24|5|Cum timerent autem et declinarent vultum in terram, dixerunt ad illas: " Quid quaeritis viventem cum mortuis?
LUKE|24|6|Non est hic, sed surrexit. Recordamini qualiter locutus est vobis, cum adhuc in Galilaea esset,
LUKE|24|7|dicens: "Oportet Filium hominis tradi in manus hominum peccatorum et crucifigi et die tertia resurgere" ".
LUKE|24|8|Et recordatae sunt verborum eius
LUKE|24|9|et regressae a monumento nuntiaverunt haec omnia illis Undecim et ceteris omnibus.
LUKE|24|10|Erat autem Maria Magdalene et Ioanna et Maria Iacobi; et ceterae cum eis dicebant ad apostolos haec.
LUKE|24|11|Et visa sunt ante illos sicut deliramentum verba ista, et non credebant illis.
LUKE|24|12|Petrus autem surgens cucurrit ad monumentum et procumbens videt linteamina sola; et rediit ad sua mirans, quod factum fuerat.
LUKE|24|13|Et ecce duo ex illis ibant ipsa die in castellum, quod erat in spatio stadiorum sexaginta ab Ierusalem nomine Emmaus;
LUKE|24|14|et ipsi loquebantur ad invicem de his omnibus, quae acciderant.
LUKE|24|15|Et factum est, dum fabularentur et secum quaererent, et ipse Iesus appropinquans ibat cum illis;
LUKE|24|16|oculi autem illorum tenebantur, ne eum agnoscerent.
LUKE|24|17|Et ait ad illos: " Qui sunt hi sermones, quos confertis ad invicem ambulantes? ". Et steterunt tristes.
LUKE|24|18|Et respondens unus, cui nomen Cleopas, dixit ei: " Tu solus peregrinus es in Ierusalem et non cognovisti, quae facta sunt in illa his diebus? ".
LUKE|24|19|Quibus ille dixit: " Quae? ". Et illi dixerunt ei: " De Iesu Nazareno, qui fuit vir propheta, potens in opere et sermone coram Deo et omni populo;
LUKE|24|20|et quomodo eum tradiderunt summi sacerdotes et principes nostri in damnationem mortis et crucifixerunt eum.
LUKE|24|21|Nos autem sperabamus, quia ipse esset redempturus Israel; at nunc super haec omnia tertia dies hodie quod haec facta sunt.
LUKE|24|22|Sed et mulieres quaedam ex nostris terruerunt nos, quae ante lucem fuerunt ad monumentum
LUKE|24|23|et, non invento corpore eius, venerunt dicentes se etiam visionem angelorum vidisse, qui dicunt eum vivere.
LUKE|24|24|Et abierunt quidam ex nostris ad monumentum et ita invenerunt, sicut mulieres dixerunt, ipsum vero non viderunt ".
LUKE|24|25|Et ipse dixit ad eos: " O stulti et tardi corde ad credendum in omnibus, quae locuti sunt Prophetae!
LUKE|24|26|Nonne haec oportuit pati Christum et intrare in gloriam suam? ".
LUKE|24|27|Et incipiens a Moyse et omnibus Prophetis interpretabatur illis in omnibus Scripturis, quae de ipso erant.
LUKE|24|28|Et appropinquaverunt castello, quo ibant, et ipse se finxit longius ire.
LUKE|24|29|Et coegerunt illum dicentes: " Mane nobiscum, quoniam advesperascit, et inclinata est iam dies ". Et intravit, ut maneret cum illis.
LUKE|24|30|Et factum est, dum recumberet cum illis, accepit panem et benedixit ac fregit et porrigebat illis.
LUKE|24|31|Et aperti sunt oculi eorum, et cognoverunt eum; et ipse evanuit ab eis.
LUKE|24|32|Et dixerunt ad invicem: " Nonne cor nostrum ardens erat in nobis, dum loqueretur nobis in via et aperiret nobis Scripturas? ".
LUKE|24|33|Et surgentes eadem hora regressi sunt in Ierusalem et invenerunt congregatos Undecim et eos, qui cum ipsis erant,
LUKE|24|34|dicentes: " Surrexit Dominus vere et apparuit Simoni ".
LUKE|24|35|Et ipsi narrabant, quae gesta erant in via, et quomodo cognoverunt eum in fractione panis.
LUKE|24|36|Dum haec autem loquuntur, ipse stetit in medio eorum et dicit eis: " Pax vobis! ".
LUKE|24|37|Conturbati vero et conterriti existimabant se spiritum videre.
LUKE|24|38|Et dixit eis: " Quid turbati estis, et quare cogitationes ascendunt in corda vestra?
LUKE|24|39|Videte manus meas et pedes meos, quia ipse ego sum! Palpate me et videte, quia spiritus carnem et ossa non habet, sicut me videtis habere ".
LUKE|24|40|Et cum hoc dixisset, ostendit eis manus et pedes.
LUKE|24|41|Adhuc autem illis non credentibus prae gaudio et mirantibus, dixit eis: Habetis hic aliquid, quod manducetur? ".
LUKE|24|42|At illi obtulerunt ei partem piscis assi.
LUKE|24|43|Et sumens, coram eis manducavit.
LUKE|24|44|Et dixit ad eos: " Haec sunt verba, quae locutus sum ad vos, cum adhuc essem vobiscum, quoniam necesse est impleri omnia, quae scripta sunt in Lege Moysis et Prophetis et Psalmis de me ".
LUKE|24|45|Tunc aperuit illis sensum, ut intellegerent Scripturas.
LUKE|24|46|Et dixit eis: " Sic scriptum est, Christum pati et resurgere a mortuis die tertia,
LUKE|24|47|et praedicari in nomine eius paenitentiam in remissionem peccatorum in omnes gentes, incipientibus ab Ierusalem.
LUKE|24|48|Vos estis testes horum.
LUKE|24|49|Et ecce ego mitto promissum Patris mei in vos; vos autem sedete in civitate, quoadusque induamini virtutem ex alto ".
LUKE|24|50|Eduxit autem eos foras usque in Bethaniam et, elevatis manibus suis, benedixit eis.
LUKE|24|51|Et factum est, dum benediceret illis, recessit ab eis et ferebatur in caelum.
LUKE|24|52|Et ipsi adoraverunt eum et regressi sunt in Ierusalem cum gaudio magno
LUKE|24|53|et erant semper in templo benedicentes Deum.
