ACTS|1|1|Першу книгу я був написав, о Теофіле, про все те, що Ісус від початку чинив та навчав,
ACTS|1|2|аж до дня, коли через Духа Святого подав Він накази апостолам, що їх вибрав, і вознісся.
ACTS|1|3|А по муці Своїй Він ставав перед ними живий із засвідченнями багатьма, і сорок день їм з'являвся та про Божеє Царство казав.
ACTS|1|4|А зібравшися з ними, Він звелів, щоб вони не відходили з Єрусалиму, а чекали обітниці Отчої, що про неї казав ви чули від Мене.
ACTS|1|5|Іван бо водою христив, ви ж охрищені будете Духом Святим через кілька тих днів!
ACTS|1|6|А вони, зійшовшись, питали Його й говорили: Чи не часу цього відбудуєш Ти, Господи, царство Ізраїлеві?
ACTS|1|7|А Він їм відказав: То не ваша справа знати час та добу, що Отець поклав у владі Своїй.
ACTS|1|8|Та ви приймете силу, як Дух Святий злине на вас, і Моїми ви свідками будете в Єрусалимі, і в усій Юдеї та в Самарії, та аж до останнього краю землі.
ACTS|1|9|І, прорікши оце, як дивились вони, Він угору возноситись став, а хмара забрала Його сперед їхніх очей...
ACTS|1|10|А коли вони пильно дивились на небо, як Він віддалявся, то два мужі у білій одежі ось стали при них,
ACTS|1|11|та й сказали: Галілейські мужі, чого стоїте й задивляєтесь на небо? Той Ісус, що вознісся на небо від вас, прийде так, як бачили ви, як ішов Він на небо!
ACTS|1|12|Тоді вони повернулись до Єрусалиму з гори, що Оливною зветься, і що знаходиться поблизько Єрусалиму, на віддаль дороги суботнього дня.
ACTS|1|13|А прийшовши, увійшли вони в горницю, де й перебували: Петро та Іван, та Яків та Андрій, Пилип та Фома, Варфоломій та Матвій, Яків Алфеїв та Симон Зилот, та Юда Яковів.
ACTS|1|14|Вони всі однодушно були на невпинній молитві, із жінками, і з Марією, матір'ю Ісусовою, та з братами Його.
ACTS|1|15|Тими ж днями Петро став посеред братів а народу було поіменно до ста двадцяти та й промовив:
ACTS|1|16|Мужі-браття! Належало збутись Писанню тому, що устами Давидовими Дух Святий був прорік про Юду, який показав дорогу для тих, хто Ісуса схопив,
ACTS|1|17|бо він був зарахований з нами, і жереб служіння оцього прийняв.
ACTS|1|18|І він поле набув за заплату злочинства, а впавши сторчма, він тріснув надвоє, і все нутро його вилилось...
ACTS|1|19|І стало відоме це всім, хто замешкує в Єрусалимі, тому й поле те назване їхньою мовою Акелдама, що є: Поле крови.
ACTS|1|20|Бо написано в книзі Псалмів: Нехай пусткою стане мешкання його, і нехай пожильця в нім не буде, а також: А служіння його забере нехай інший.
ACTS|1|21|Отже треба, щоб один із тих мужів, що сходились з нами повсякчас, як Господь Ісус входив і виходив між нами,
ACTS|1|22|зачавши від хрищення Іванового аж до дня, коли Він вознісся від нас, щоб той разом із нами був свідком Його воскресення.
ACTS|1|23|І поставили двох: Йосипа, що Варсавою зветься, і що Юстом був названий, та Маттія.
ACTS|1|24|А молившись, казали: Ти, Господи, знавче всіх сердець, покажи з двох одного, котрого Ти вибрав,
ACTS|1|25|щоб він зайняв місце тієї служби й апостольства, що Юда від нього відпав, щоб іти в своє місце.
ACTS|1|26|І дали жеребки їм, і впав жеребок на Маттія, і він зарахований був до одинадцятьох апостолів.
ACTS|2|1|Коли ж почався день П'ятдесятниці, всі вони однодушно знаходилися вкупі.
ACTS|2|2|І нагло зчинився шум із неба, ніби буря раптова зірвалася, і переповнила ввесь той дім, де сиділи вони.
ACTS|2|3|І з'явилися їм язики поділені, немов би огненні, та й на кожному з них по одному осів.
ACTS|2|4|Усі ж вони сповнились Духом Святим, і почали говорити іншими мовами, як їм Дух промовляти давав.
ACTS|2|5|Перебували ж в Єрусалимі юдеї, люди побожні, від усякого народу під небом.
ACTS|2|6|А коли оцей гомін зчинився, зібралася безліч народу, та й диву далися, бо кожен із них тут почув, що вони розмовляли їхньою власною мовою!...
ACTS|2|7|Усі ж побентежилися та дивувалися, та й казали один до одного: Хіба ж не галілеяни всі ці, що говорять?
ACTS|2|8|Як же кожен із нас чує свою власну мову, що ми в ній народились?
ACTS|2|9|Парфяни та мідяни та еламіти, також мешканці Месопотамії, Юдеї та Каппадокії, Понту та Азії,
ACTS|2|10|і Фріґії та Памфілії, Єгипту й лівійських земель край Кірени, і захожі римляни,
ACTS|2|11|юдеї й нововірці, крітяни й араби, усі чуємо ми, що говорять вони про великі діла Божі мовами нашими!
ACTS|2|12|І всі не виходили з дива, і безрадні були, і говорили один до одного: Що ж то статися має?
ACTS|2|13|А інші казали глузуючи: Вони повпивались вином молодим!
ACTS|2|14|Ставши ж Петро із Одинадцятьма, свій голос підніс та й промовив до них: Мужі юдейські та мешканці Єрусалиму! Нехай вам оце стане відоме, і послухайте слів моїх!
ACTS|2|15|Бо не п'яні вони, як ви думаєте, бо третя година дня,
ACTS|2|16|а це те, що пророк Йоіл передрік:
ACTS|2|17|І буде останніми днями, говорить Господь: Я виллю від Духа Свого на всяке тіло, і будуть пророкувати сини ваші та ваші доньки, юнаки ж ваші бачити будуть видіння, а старим вашим сни будуть снитися.
ACTS|2|18|І на рабів Моїх і на рабинь Моїх за тих днів Я також виллю від Духа Свого, і пророкувати вони будуть!
ACTS|2|19|І дам чуда на небі вгорі, а внизу на землі ці знамена: кров, і огонь, і куряву диму.
ACTS|2|20|Переміниться сонце на темряву, а місяць на кров, перше ніж день Господній настане, великий та славний!
ACTS|2|21|І станеться, що кожен, хто покличе Господнє Ім'я, той спасеться.
ACTS|2|22|Мужі ізраїльські, послухайте ви оцих слів: Ісуса Назарянина, Мужа, що Його Бог прославив вам силою, і чудами, і тими знаменами, що Бог через Нього вчинив серед вас, як самі ви те знаєте,
ACTS|2|23|Того, що був виданий певною волею та передбаченням Божим, ви руками беззаконників розп'яли та забили.
ACTS|2|24|Та Бог воскресив Його, пута смерти усунувши, вона бо тримати Його не могла.
ACTS|2|25|Бо каже про Нього Давид: Мав я Господа завсіди перед очима своїми, бо Він по правиці моїй, щоб я не захитався.
ACTS|2|26|Тому серце моє звеселилось, і зрадів мій язик, і тіло моє відпочине в надії.
ACTS|2|27|Бо не позоставиш Ти в аду моєї душі, і не даси Ти Своєму Святому побачити тління!
ACTS|2|28|Ти дороги життя об'явив мені, Ти мене переповниш утіхою перед обличчям Своїм!
ACTS|2|29|Мужі-браття! Нехай буде вільно мені сміло сказати вам про патріярха Давида, що помер і похований, і знаходиться гріб його в нас аж до цього дня.
ACTS|2|30|А бувши ж пророком, та відаючи, що Бог клятвою клявся йому посадити на престолі його від плоду його стегон,
ACTS|2|31|у передбаченні він говорив про Христове воскресення, що не буде зоставлений в аду, ані тіло Його не зазнає зотління.
ACTS|2|32|Бог Ісуса Цього воскресив, чого свідки всі ми!
ACTS|2|33|А отож, як правицею Божою був Він вознесений, і обітницю Духа Святого прийняв від Отця, то й злив Він оте, що ви бачите й чуєте.
ACTS|2|34|Не зійшов бо на небо Давид, але сам він говорить: Промовив Господь Господеві моєму: Сядь праворуч Мене,
ACTS|2|35|доки не покладу Я Твоїх ворогів підніжком ногам Твоїм!
ACTS|2|36|Ото ж, нехай ввесь Ізраїлів дім твердо знає, що і Господом, і Христом учинив Бог Його, Того Ісуса, що Його розп'яли ви!
ACTS|2|37|Як почули ж оце, вони серцем розжалобились, та й сказали Петрові та іншим апостолам: Що ж ми маємо робити, мужі-браття?
ACTS|2|38|А Петро до них каже: Покайтеся, і нехай же охриститься кожен із вас у Ім'я Ісуса Христа на відпущення ваших гріхів, і дара Духа Святого ви приймете!
ACTS|2|39|Бо для вас ця обітниця, і для ваших дітей, і для всіх, що далеко знаходяться, кого б тільки покликав Господь, Бог наш.
ACTS|2|40|І іншими багатьома словами він засвідчував та вмовляв їх, говорячи: Рятуйтесь від цього лукавого роду!
ACTS|2|41|Отож ті, хто прийняв його слово, охристилися. І пристало до них того дня душ тисяч зо три!
ACTS|2|42|І вони перебували в науці апостольській, та в спільноті братерській, і в ламанні хліба, та в молитвах.
ACTS|2|43|І був острах у кожній душі, бо багато чинили апостоли чуд та знамен.
ACTS|2|44|А всі віруючі були вкупі, і мали все спільним.
ACTS|2|45|І вони продавали маєтки та добра, і всім їх ділили, як кому чого треба було.
ACTS|2|46|І кожного дня перебували вони однодушно у храмі, і, ломлячи хліб по домах, поживу приймали із радістю та в сердечній простоті,
ACTS|2|47|вихваляючи Бога та маючи ласку в усього народу. І щоденно до Церкви Господь додавав тих, що спасалися.
ACTS|3|1|А Петро та Іван на дев'яту годину молитви йшли разом у храм.
ACTS|3|2|І несено там чоловіка одного, що кривий був з утроби своєї матері. Його садовили щоденно в воротях храму, що Красними звалися, просити милостині від тих, хто до храму йшов.
ACTS|3|3|Як побачив же він, що Петро та Іван хочуть у храм увійти, став просити в них милостині.
ACTS|3|4|Петро ж із Іваном поглянув на нього й сказав: Подивися на нас!
ACTS|3|5|І той подивився на них, сподіваючися щось дістати від них.
ACTS|3|6|Та промовив Петро: Срібла й золота в мене нема, але що я маю, даю тобі: У Ім'я Ісуса Христа Назарянина устань та й ходи!
ACTS|3|7|І, узявши його за правицю, він підвів його. І хвилі тієї зміцнилися ноги й суглобці його!...
ACTS|3|8|І, зірвавшись, він устав та й ходив, і з ними у храм увійшов, ходячи та підскакуючи, і хвалячи Бога!
ACTS|3|9|Народ же ввесь бачив, як ходив він та Бога хвалив.
ACTS|3|10|І пізнали його, що це той, що при Красних воротях храму сидів ради милостині. І вони переповнились жахом та подивом із того, що сталось йому!
ACTS|3|11|А тому, що тримався він Петра та Івана, увесь народ зачудований збігся до них на той ґанок, який Соломоновим зветься.
ACTS|3|12|І, побачивши це, промовив Петро до народу: Мужі ізраїльські! Чого ви дивуєтесь цим, та чого ви на нас позираєте так, ніби те, що він ходить, ми зробили своєю силою чи благочестям?
ACTS|3|13|Бог Авраамів, та Ісаків, та Яковів, Бог наших батьків, Сина Свого прославив, Ісуса, Якого ви видали, і відцуралися перед Пилатом, як він присудив був пустити Його.
ACTS|3|14|Але ви відцурались Святого та Праведного, і домагалися видати вам душогубця.
ACTS|3|15|Начальника ж життя ви забили, та Його воскресив Бог із мертвих, чого свідками ми!
ACTS|3|16|І через віру в Ім'я Його вздоровило Ім'я Його того, кого бачите й знаєте. І віра, що від Нього, принесла йому вздоровлення це перед вами всіма.
ACTS|3|17|А тепер, браття, знаю, що вчинили ви це з несвідомости, як і ваші начальники.
ACTS|3|18|А Бог учинив так, як Він провіщав був устами Своїх усіх пророків, щоб терпіти Христові.
ACTS|3|19|Покайтеся ж та наверніться, щоб Він змилувався над вашими гріхами,
ACTS|3|20|щоб часи відпочинку прийшли від обличчя Господнього, і щоб послав заповідженого вам Ісуса Христа,
ACTS|3|21|що Його небо мусить прийняти аж до часу відновлення всього, про що провіщав Бог від віку устами всіх святих пророків Своїх!
ACTS|3|22|Бо Мойсей провіщав: Господь Бог вам Пророка підійме від ваших братів, як мене; у всім Його слухайтеся, про що тільки Він вам говоритиме!
ACTS|3|23|І станеться, що кожна душа, яка не послухала б того Пророка, знищена буде з народу.
ACTS|3|24|Так само всі пророки від Самуїла й наступних, скільки їх говорило, також провіщали ці дні.
ACTS|3|25|Сини ви пророків і того заповіту, що Бог вашим батькам заповів, промовляючи до Авраама: І в насінні твоїм усі народи землі благословлені будуть!
ACTS|3|26|Воскресивши Свого Отрока, Бог послав Його перше до вас, щоб вас поблагословити, щоб кожен із вас відвернувся від злих своїх учинків!
ACTS|4|1|А коли промовляли вони до народу оце, до них приступили священики, і влада сторожі храму й саддукеї,
ACTS|4|2|обурюючись, що навчають народ та звіщають в Ісусі воскресіння з мертвих.
ACTS|4|3|І руки наклали на них, і до в'язниці всадили до ранку, бо вже вечір настав був.
ACTS|4|4|І багато-хто з тих, хто слухав слово, увірували; число ж мужів таких було тисяч із п'ять.
ACTS|4|5|І сталось, що ранком зібралися в Єрусалимі начальники їхні, і старші та книжники,
ACTS|4|6|і Анна первосвященик, і Кайяфа, і Іван, і Олександер, і скільки було їх із роду первосвященичого.
ACTS|4|7|І, поставивши їх посередині, запиталися: Якою ви силою чи яким ви ім'ям те робили?
ACTS|4|8|Тоді Петро, переповнений Духом Святим, промовив до них: Начальники люду та старшини Ізраїлеві!
ACTS|4|9|Як сьогодні беруть нас на допит про те добродійство недужій людині, як вона вздоровлена,
ACTS|4|10|нехай буде відомо всім вам, і всім людям Ізраїлевим, що Ім'ям Ісуса Христа Назарянина, що Його розп'яли ви, то Його воскресив Бог із мертвих, Ним поставлений він перед вами здоровий!
ACTS|4|11|Він камінь, що ви, будівничі, відкинули, але каменем став Він наріжним!
ACTS|4|12|І нема ні в кім іншім спасіння. Бо під небом нема іншого Ймення, даного людям, що ним би спастися ми мали.
ACTS|4|13|А бачивши сміливість Петра та Івана, і спостерігши, що то люди обидва невчені та прості, дивувалися, і пізнали їх, що вони з Ісусом були.
ACTS|4|14|Та бачивши, що вздоровлений чоловік стоїть з ними, нічого навпроти сказати не могли.
ACTS|4|15|І, звелівши їм вийти із синедріону, зачали радитися між собою,
ACTS|4|16|говорячи: Що робити нам із цими людьми? Бож усім мешканцям Єрусалиму відомо, що вчинили вони явне чудо, і не можемо того заперечити.
ACTS|4|17|Та щоб більш не поширювалось це в народі, то з погрозою заборонімо їм, щоб нікому з людей вони не говорили про Це Ім'я.
ACTS|4|18|І, закликавши їх, наказали їм не говорити, і взагалі не навчати про Ісусове Ймення.
ACTS|4|19|І відповіли їм Петро та Іван, та й сказали: Розсудіть, чи це справедливе було б перед Богом, щоб слухатись вас більш, як Бога?
ACTS|4|20|Бо не можемо ми не казати про те, що ми бачили й чули!
ACTS|4|21|А вони пригрозили їм ще, і відпустили їх, не знайшовши нічого, щоб їх покарати, через людей, бо всі славили Бога за теє, що сталось.
ACTS|4|22|Бо років більш сорока мав той чоловік, що на нім відбулося це чудо вздоровлення.
ACTS|4|23|Коли ж їх відпустили, вони до своїх прибули й сповістили, про що первосвященики й старші до них говорили.
ACTS|4|24|Вони ж, вислухавши, однодушно свій голос до Бога піднесли й промовили: Владико, що небо, і землю, і море, і все, що в них є, Ти створив!
ACTS|4|25|Ти устами Давида, Свого слуги, отця нашого, сказав Духом Святим: Чого люди бунтуються, а народи задумують марне?
ACTS|4|26|Повстають царі земні, і збираються старші докупи на Господа та на Христа Його.
ACTS|4|27|Бо справді зібралися в місці оцім проти Отрока Святого Твого Ісуса, що Його намастив Ти, Ірод та Понтій Пилат із поганами та з народом Ізраїлевим,
ACTS|4|28|учинити оте, що рука Твоя й воля Твоя наперед встановили були, щоб збулося.
ACTS|4|29|І тепер споглянь, Господи, на їхні погрози, і дай Своїм рабам із повною сміливістю слово Твоє повідати,
ACTS|4|30|коли руку Свою простягатимеш Ти на вздоровлення, і щоб знамена та чуда чинились Ім'ям Твого Святого Отрока Ісуса.
ACTS|4|31|Як вони ж помолились, затряслося те місце, де зібрались були, і переповнилися всі Святим Духом, і зачали говорити Слово Боже з сміливістю!
ACTS|4|32|А люди, що ввірували, мали серце одне й одну душу, і жаден із них не вважав що з маєтку свого за своє, але в них усе спільним було.
ACTS|4|33|І апостоли з великою силою свідчили про воскресення Ісуса Господа, і благодать велика на всіх них була!
ACTS|4|34|Бо жаден із них не терпів недостачі: бо, хто мав поле чи дім, продавали, і заплату за продаж приносили,
ACTS|4|35|та й клали в ногах у апостолів, і роздавалося кожному, хто потребу в чім мав.
ACTS|4|36|Так, Йосип, що Варнавою що в перекладі є син потіхи був прозваний від апостолів, Левит, родом кіпрянин,
ACTS|4|37|мавши поле, продав, а гроші приніс, та й поклав у ногах у апостолів.
ACTS|5|1|А один чоловік, на ймення Ананій, із своєю дружиною Сапфірою, продав був маєтка,
ACTS|5|2|та й з відома дружини своєї присвоїв частину з заплати, а якусь там частину приніс та й поклав у ногах у апостолів.
ACTS|5|3|І промовив Петро: Ананію, чого сатана твоє серце наповнив, щоб ти Духу Святому неправду сказав та присвоїв із заплати за землю?
ACTS|5|4|Хіба те, що ти мав, не твоє все було, а продане не в твоїй владі було? Чого ж в серце своє ти цю справу поклав? Ти не людям неправду сказав, але Богові!
ACTS|5|5|Як Ананій зачув ці слова, то впав та й умер... І обгорнув жах великий усіх, що це чули!
ACTS|5|6|Юнаки ж повставали, обгорнули його, і винесли та й поховали.
ACTS|5|7|І сталось, годин через три прийшла й дружина його, про випадок нічого не знавши.
ACTS|5|8|І промовив до неї Петро: Скажи мені, чи за стільки ви землю оту продали? Вона ж відказала: Так, за стільки.
ACTS|5|9|До неї ж Петро: Чому це ви змовилися спокушувати Господнього Духа? Он ті входять у двері, що чоловіка твого поховали, і тебе вони винесуть...
ACTS|5|10|І вона зараз упала до ніг його, та й умерла. Як ввійшли ж юнаки, то знайшли її мертвою, і, винісши, біля мужа її поховали.
ACTS|5|11|І обгорнув страх великий всю Церкву та всіх, що чули про це...
ACTS|5|12|А руками апостолів стались знамена та чуда великі в народі. І були однодушно всі в Соломоновім ґанку.
ACTS|5|13|А з сторонніх ніхто приставати не важивсь до них, але люд прославляв їх.
ACTS|5|14|І все збільшувалось тих, хто вірує в Господа, безліч чоловіків і жінок,
ACTS|5|15|так що хворих стали виносити на вулиці, та й клали на ложа та ноші, щоб, як ітиме Петро, то хоч тінь його впала б на кого із них.
ACTS|5|16|І безліч люду збиралась до Єрусалиму з довколишніх міст, і несли недужих та хворих від духів нечистих, і були вони всі вздоровлювані!
ACTS|5|17|А первосвященик, уставши, та й усі, хто був із ним, хто належав до саддукейської єресі, переповнились заздрощами,
ACTS|5|18|і руки наклали вони на апостолів, і до в'язниці громадської вкинули їх.
ACTS|5|19|Але Ангол Господній вночі відчинив для них двері в'язничні, і, вивівши їх, проказав:
ACTS|5|20|Ідіть, і, ставши, говоріть до народу у храмі всі слова цього життя.
ACTS|5|21|Як це вчули вони, то в храм рано ввійшли і навчали. А первосвященик і ті, хто був із ним, прийшовши, скликали синедріон і всіх старших з Ізраїлевих синів. І послали в в'язницю, щоб їх привели.
ACTS|5|22|А служба, прийшовши, не знайшла їх у в'язниці, а вернувшись, сповістила,
ACTS|5|23|говорячи: В'язницю знайшли ми з великою пильністю замкнену, і сторожу, що при дверях стояла; а коли відчинили, то нікого всередині ми не знайшли!
ACTS|5|24|Як почули слова ці начальник сторожі храму та первосвященики, не могли зрозуміти вони, що б то сталося.
ACTS|5|25|Та прийшовши один, сповістив їх, говорячи: Ось ті мужі, що ви їх до в'язниці всадили були, у храмі стоять та й навчають народ.
ACTS|5|26|Пішов тоді старший сторожі зо службою, та й привів їх без насильства, бо боялись народу, щоб їх не побили камінням.
ACTS|5|27|Припровадивши ж їх, поставили перед синедріоном. І спитався їх первосвященик, говорячи:
ACTS|5|28|Чи ми не заборонили з погрозою вам, щоб про Те Ім'я не навчати? І ото, ви своєю наукою переповнили Єрусалим, і хочете кров Чоловіка Того припровадити на нас...
ACTS|5|29|Відповів же Петро та сказали апостоли: Бога повинно слухатися більш, як людей!
ACTS|5|30|Бог наших отців воскресив нам Ісуса, Якому ви смерть були заподіяли, повісивши на дереві.
ACTS|5|31|Його Бог підвищив Своєю правицею на Начальника й Спаса, щоб дати Ізраїлеві покаяння і прощення гріхів.
ACTS|5|32|А тих справ Йому свідками ми й Святий Дух, що Його Бог дав тим, хто слухняний Йому.
ACTS|5|33|Як зачули ж оце, запалилися гнівом вони, та й радилися, як їм смерть заподіяти?...
ACTS|5|34|І встав у синедріоні один фарисей, Гамаліїл на ймення, учитель Закону, поважаний від усього народу, та й звелів на часинку апостолів вивести.
ACTS|5|35|І промовив до них: Мужі ізраїльські! Поміркуйте собі про людей цих, що з ними робити ви маєте.
ACTS|5|36|Бо перед цими днями повстав був Тевда та й казав, що великий він хтось, і до нього пристало з чотириста люда. Він забитий, а всі ті, хто слухав його, розпорошились та обернулись в ніщо.
ACTS|5|37|Після нього повстав, під час перепису, Галілеянин Юда, та й багато людей потягнув за собою. Загинув і він, а всі ті, хто слухав його, розпорошились.
ACTS|5|38|І тепер кажу вам: Відступіться від цих людей, і занехайте їх! Бо коли від людей оця рада чи справа ця буде, розпадеться вона.
ACTS|5|39|А коли те від Бога, то того зруйнувати не зможете, щоб випадком не стати і вам богоборцями! І послухались ради його.
ACTS|5|40|І, покликавши знов апостолів, вибили їх, наказали їм не говорити про Ісусове Ймення, та й їх відпустили.
ACTS|5|41|А вони поверталися з синедріону, радіючи, що сподобились прийняти зневагу за Ймення Господа Ісуса.
ACTS|5|42|І щоденно у храмі й домах безупинно навчали, і звіщали Євангелію Ісуса Христа.
ACTS|6|1|Тими ж днями, як учнів намножилось, зачали нарікати на євреїв огречені, що в щоденному служінні їхні вдовиці занедбані.
ACTS|6|2|Тоді ті Дванадцять покликали багатьох учнів та й сказали: Нам не личить покинути Боже Слово, і служити при столах.
ACTS|6|3|Отож, браття, виглядіть ізпоміж себе сімох мужів доброї слави, повних Духа Святого та мудрости, їх поставимо на службу оцю.
ACTS|6|4|А ми перебуватимемо завжди в молитві та в служінні слову.
ACTS|6|5|І всім людям сподобалося оце слово, і обрали Степана, мужа повного віри та Духа Святого, і Пилипа, і Прохора та Никанора, і Тимона та Пармена, і нововірця Миколу з Антіохії,
ACTS|6|6|їх поставили перед апостолів, і, помолившись, вони руки поклали на них.
ACTS|6|7|І росло Слово Боже, і дуже множилося число учнів у Єрусалимі, і дуже багато священиків були слухняні вірі.
ACTS|6|8|А Степан, повний віри та сили, чинив між народом великі знамена та чуда.
ACTS|6|9|Тому дехто повстав із синагоги, що зветься лібертинська, і кірінейська, і олександрійська, та з тих, хто походить із Кілікії та з Азії, і зачали сперечатись із Степаном.
ACTS|6|10|Але встояти вони не могли проти мудрости й Духа, що він Ним говорив.
ACTS|6|11|Тоді вони підмовили людей, що казали, ніби чули, як він богозневажні слова говорив на Мойсея та Бога.
ACTS|6|12|І людей попідбурювали, і старших та книжників, і, напавши, схопили його, і припровадили в синедріон.
ACTS|6|13|Також свідків фальшивих поставили, які говорили: Чоловік оцей богозневажні слова безперестань говорить на це святе місце та проти Закону.
ACTS|6|14|Бо ми чули, як він говорив, що Ісус Назарянин зруйнує це місце та змінить звичаї, які передав нам Мойсей.
ACTS|6|15|Коли всі, хто в синедріоні сидів, на нього споглянули, то бачили лице його, як лице Ангола!
ACTS|7|1|Запитав тоді первосвященик: Чи це так?
ACTS|7|2|Степан же промовив: Послухайте, мужі-браття й отці! Бог слави з'явивсь Авраамові, отцеві нашому, як він у Месопотамії був, перше ніж оселився в Харані,
ACTS|7|3|і промовив до нього: Вийди із своєї землі та від роду свого, та й піди до землі, що тобі покажу.
ACTS|7|4|Тоді він вийшов із землі халдейської, та й оселився в Харані. А звідти, як умер йому батько, Він переселив його в землю оцю, що на ній ви живете тепер.
ACTS|7|5|Та спадщини на ній Він не дав йому навіть на крок, але обіцяв дати її на володіння йому й його родові по нім, хоч дитини не мав він.
ACTS|7|6|І сказав Бог отак, що насіння його буде приходьком у краї чужому, і поневолять його, і будуть гнобити чотириста років.
ACTS|7|7|Але Я сказав Бог буду судити народ, що його поневолить. Опісля ж вони вийдуть, і будуть служити Мені на цім місці.
ACTS|7|8|І дав Він йому заповіта обрізання. І породив так Ісака, і восьмого дня він обрізав його. А Ісак породив Якова, а Яків дванадцятьох патріярхів.
ACTS|7|9|А ті патріярхи позаздрили Йосипові, і продали його до Єгипту. Але Бог був із ним,
ACTS|7|10|і його визволив від усіх його утисків, і дав йому благодать та мудрість перед фараоном, царем єгипетським, а він настановив його за правителя над Єгиптом та всім своїм домом.
ACTS|7|11|А як голод прийшов на всю землю єгипетську та ханаанську, та велика біда, то поживи тоді не знаходили наші батьки.
ACTS|7|12|Коли ж Яків зачув, що в Єгипті є збіжжя, то послав батьків наших уперше.
ACTS|7|13|А як удруге послав, то був пізнаний Йосип братами своїми, і фараонові знаний став Йосипів рід.
ACTS|7|14|Тоді Йосип послав, щоб покликати Якова, батька свого, та всю родину свою сімдесят і п'ять душ.
ACTS|7|15|І подався Яків в Єгипет, та й умер там він сам та наші батьки.
ACTS|7|16|І їх перенесли в Сихем, і поклали до гробу, що Авраам був купив за ціну срібла від синів Еммора Сихемового.
ACTS|7|17|А коли наближавсь час обітниці, що нею Бог клявсь Авраамові, розрісся народ і намножився в Єгипті,
ACTS|7|18|аж поки настав інший цар ув Єгипті, що не знав уже Йосипа.
ACTS|7|19|Він хитро наш люд обманив, і силою змушував наших отців викидати дітей своїх, щоб вони не лишались живі.
ACTS|7|20|Того часу родився Мойсей, і гарний він був перед Богом. Він годований був у домі батька свойого три місяці.
ACTS|7|21|А коли він був викинений, то дочка фараона забрала його, та й за сина собі його викохала.
ACTS|7|22|І Мойсей був навчений всієї премудрости єгипетської, і був міцний у словах та в ділах своїх.
ACTS|7|23|А коли йому сповнилося сорок років, йому спало на серце відвідати братів своїх, синів Ізраїлевих.
ACTS|7|24|Як угледів же він, що одному з них діється кривда, заступився, і відомстив за окривдженого, убивши єгиптянина.
ACTS|7|25|Він же думав, що брати розуміють, що рукою його Бог дає їм визволення, та не зрозуміли вони.
ACTS|7|26|А наступного дня, як сварились вони, він з'явився й хотів погодити їх, кажучи: Люди, ви браття, чого один одного кривдите?
ACTS|7|27|А той, що ближнього кривдив, його відіпхнув та сказав: Хто наставив над нами тебе за старшого й суддю?
ACTS|7|28|Чи хочеш убити й мене, як учора вбив ти єгиптянина?
ACTS|7|29|І втік Мойсей через слово оце, і стався приходьком у землі мадіямській, де зродив двох синів.
ACTS|7|30|А коли сорок років проминуло, то з'явивсь йому Ангол Господній у полум'ї куща огняного в пустині Сінайської гори.
ACTS|7|31|А Мойсей, як побачив, дивувався з видіння. А коли підійшов, щоб розглянути, був голос Господній до нього:
ACTS|7|32|Я Бог отців твоїх, Бог Авраамів, і Бог Ісаків, і Бог Яковів! І затрусився Мойсей, і не відваживсь поглянути...
ACTS|7|33|І промовив до нього Господь: Скинь взуття з своїх ніг, бо те місце, на якому стоїш, то святая земля!
ACTS|7|34|Добре бачив Я утиск народу Свого, що в Єгипті, і стогін його Я почув, і зійшов, щоб їх визволити. Тепер ось іди, Я пошлю до Єгипту тебе.
ACTS|7|35|Цього Мойсея, що його відцурались вони, сказавши: Хто наставив тебе за старшого й суддю, цього Бог через Ангола, якому з'явився в кущі, послав за старшого й визвольника.
ACTS|7|36|Він їх вивів, чуда й знамена вчинивши в землі єгипетській, і на Червоному морі, і сорок років у пустині.
ACTS|7|37|Це той Мойсей, що прорік Ізраїлевим синам: Господь Бог вам підійме Пророка від ваших братів, як мене, Його слухайте!
ACTS|7|38|Це той, що в пустині на зборах був з Анголом, який промовляв йому на Сінайській горі, та з отцями нашими, і що прийняв він живі слова, щоб їх нам передати;
ACTS|7|39|що його не хотіли отці наші слухати, але відіпхнули, і звернулися серцем своїм до Єгипту,
ACTS|7|40|промовивши до Аарона: Зроби нам богів, які йшли б перед нами, бо не знаємо, що сталося з тим Мойсеєм, який вивів нас із краю єгипетського...
ACTS|7|41|І зробили вони тими днями теля, і бовванові жертви приносили та веселилися з діл своїх рук.
ACTS|7|42|Але Бог відвернувся від них, і попустив їх вклонятися силі небесній, як написано в книзі Пророків: Чи заколення й жертви Мені ви приносили сорок років у пустині, о доме Ізраїлів?
ACTS|7|43|Ви ж носили намета Молохового, і зорю вашого бога Ромфана, зображення, що їх ви зробили, щоб вклонятися їм... Через те запроваджу вас аж за Вавилон!
ACTS|7|44|У наших отців на пустині була скинія свідоцтва, як Той ізвелів, Хто Мойсею казав, щоб зробив її за зразком, якого він бачив.
ACTS|7|45|Її наші отці й узяли, і внесли з Ісусом у землю народів, яких вигнав Бог з-перед обличчя наших отців, аж до часу Давида.
ACTS|7|46|Він у Бога знайшов благодать, і просив, щоб оселю знайти для Бога Якова.
ACTS|7|47|І Соломон збудував Йому дім.
ACTS|7|48|Але не в рукотворнім Всевишній живе, як говорить пророк:
ACTS|7|49|Мені небо престол, а земля то підніжок ногам Моїм! Який Мені дім ви збудуєте, говорить Господь, або місце яке для Мого відпочинку?
ACTS|7|50|Хіба не рука Моя все це створила?...
ACTS|7|51|О ви, твердошиї, люди серця й вух необрізаних! Ви завжди противитесь Духові Святому, як ваші батьки, так і ви!
ACTS|7|52|Котрого з пророків батьки ваші не переслідували? Вони ж тих повбивали, хто звіщав прихід Праведного, Якому тепер ви сталися зрадниками та убійниками,
ACTS|7|53|ви, що Закона одержали через зарядження Анголів, та не зберігали його!...
ACTS|7|54|Як зачули ж оце, вони запалилися гнівом у серцях своїх, і скреготали зубами на нього...
ACTS|7|55|А Степан, повний Духа Святого, на небо споглянув, і побачив Божу славу й Ісуса, що по Божій правиці стояв,
ACTS|7|56|і промовив: Ось я бачу відчинене небо, і Сина Людського, що по Божій правиці стоїть!...
ACTS|7|57|Та вони гучним голосом стали кричати та вуха собі затуляти, та й кинулися однодушно на нього!...
ACTS|7|58|І за місто вони його вивели, і зачали побивати камінням його. А свідки плащі свої склали в ногах юнака, який звався Савлом.
ACTS|7|59|І побивали камінням Степана, що молився й казав: Господи Ісусе, прийми духа мого!...
ACTS|7|60|Упавши ж навколішки, скрикнув голосом гучним: Не залічи їм, о Господи, цього гріха! І, промовивши це, він спочив...
ACTS|8|1|А Савл похваляв його вбивство. І утиск великий постав того дня проти єрусалимської Церкви, і всі, крім апостолів, розпорошилися по краях юдейських та самарійських.
ACTS|8|2|І поховали Степана мужі побожні, і плакали ревно за ним.
ACTS|8|3|А Савл нищив Церкву, вдирався в доми, витягав чоловіків і жінок та давав до в'язниці...
ACTS|8|4|Ходили тоді розпорошенці, та Боже Слово благовістили.
ACTS|8|5|Ось Пилип прийшов до самарійського міста, і проповідував їм про Христа.
ACTS|8|6|А люди вважали на те, що Пилип говорив, і згідно слухали й бачили чуда, які він чинив.
ACTS|8|7|Із багатьох бо, що мали їх, духи нечисті виходили з криком великим, і багато розслаблених та кривих уздоровилися.
ACTS|8|8|І радість велика в тім місті була!
ACTS|8|9|Був один чоловік, на ім'я йому Симон, що до того в цім місті займавсь ворожбитством та дурив самарійський народ, видаючи себе за якогось великого.
ACTS|8|10|Його слухали всі, від найменшого аж до найбільшого, кажучи: Він сила Божа, що зветься велика!
ACTS|8|11|Його ж слухалися, бо він їх довший час дивував ворожбитством.
ACTS|8|12|Та коли йняли віри Пилипові, що благовістив про Боже Царство й Ім'я Ісуса Христа, чоловіки й жінки охристилися.
ACTS|8|13|Увірував навіть сам Симон, і, охристившись, тримався Пилипа; а бачивши чуда й знамена великі, він дуже дивувався.
ACTS|8|14|Як зачули ж апостоли, які в Єрусалимі були, що Боже Слово прийняла Самарія, то послали до них Петра та Івана.
ACTS|8|15|А вони, як прийшли, помолились за них, щоб Духа Святого вони прийняли,
ACTS|8|16|бо ще ні на одного з них Він не сходив, а були вони тільки охрищені в Ім'я Господа Ісуса.
ACTS|8|17|Тоді на них руки поклали, і прийняли вони Духа Святого!
ACTS|8|18|Як побачив же Симон, що через накладання апостольських рук Святий Дух подається, то приніс він їм гроші,
ACTS|8|19|і сказав: Дайте й мені таку владу, щоб той, на кого покладу свої руки, одержав би Духа Святого!
ACTS|8|20|Та промовив до нього Петро: Нехай згине з тобою те срібло твоє, бо ти думав набути дар Божий за гроші!
ACTS|8|21|У цім ділі нема тобі частки ні уділу, бо серце твоє перед Богом не слушне.
ACTS|8|22|Тож покайся за це лихе діло своє, і проси Господа, може прощений буде тобі замір серця твого!
ACTS|8|23|Бо я бачу, що ти пробуваєш у жовчі гіркій та в путах неправди.
ACTS|8|24|А Симон озвався й сказав: Помоліться за мене до Господа, щоб мене не спіткало нічого з того, про що ви говорили...
ACTS|8|25|А вони ж, засвідчивши, і Слово Господнє звістивши, повернулись до Єрусалиму, і звіщали Євангелію в багатьох самарійських оселях.
ACTS|8|26|А Ангол Господній промовив Пилипові, кажучи: Устань та на південь іди, на дорогу, що від Єрусалиму до Гази спускається, порожня вона.
ACTS|8|27|І, вставши, пішов він. І ось муж етіопський, скопець, вельможа Кандаки, цариці етіопської, що був над усіма її скарбами, що до Єрусалиму прибув поклонитись,
ACTS|8|28|вертався, і, сидючи на повозі своїм, читав пророка Ісаю.
ACTS|8|29|А Дух до Пилипа промовив: Підійди, та й пристань до цього повозу.
ACTS|8|30|Пилип же підбіг і почув, що той читає пророка Ісаю, та й спитав: Чи розумієш, що ти читаєш?
ACTS|8|31|А той відказав: Як же можу, як ніхто не напутить мене? І впросив він Пилипа піднятись та сісти з ним.
ACTS|8|32|А слово Писання, що його він читав, було це: Як вівцю на заріз Його ведено, і як ягня супроти стрижія безголосе, так Він не відкрив Своїх уст!
ACTS|8|33|У приниженні суд Йому віднятий був, а про рід Його хто розповість? Бо життя Його із землі забирається...
ACTS|8|34|Відізвався ж скопець до Пилипа й сказав: Благаю тебе, це про кого говорить пророк? Чи про себе, чи про іншого кого?
ACTS|8|35|А Пилип відкрив уста свої, і, зачавши від цього Писання, благовістив про Ісуса йому.
ACTS|8|36|І, як шляхом вони їхали, прибули до якоїсь води. І озвався скопець: Ось вода. Що мені заважає христитись?
ACTS|8|37|А Пилип відказав: Якщо віруєш із повного серця свого, то можна. А той відповів і сказав: Я вірую, що Ісус Христос то Син Божий!
ACTS|8|38|І звелів, щоб повіз спинився. І обидва Пилип та скопець увійшли до води, і охристив він його.
ACTS|8|39|А коли вони вийшли з води, Дух Господній Пилипа забрав, і скопець уже більше не бачив його. І він їхав, радіючи, шляхом своїм.
ACTS|8|40|А Пилип опинився в Азоті, і, переходячи, звіщав Євангелію всім містам, аж поки прийшов у Кесарію.
ACTS|9|1|А Савл, іще дишучи грізьбою й убивством на учнів Господніх, приступивши до первосвященика,
ACTS|9|2|попросив від нього листи у Дамаск синагогам, щоб, коли знайде яких чоловіків та жінок, що тієї дороги вони, то зв'язати й привести до Єрусалиму.
ACTS|9|3|А коли він ішов й наближався до Дамаску, то ось нагло осяяло світло із неба його,
ACTS|9|4|а він повалився на землю, і голос почув, що йому говорив: Савле, Савле, чому ти Мене переслідуєш?
ACTS|9|5|А він запитав: Хто Ти, Пане? А Той: Я Ісус, що Його переслідуєш ти. Трудно тобі бити ногою колючку!
ACTS|9|6|А він, затрусившися та налякавшися, каже: Чого, Господи, хочеш, щоб я вчинив? А до нього Господь: Уставай, та до міста подайся, а там тобі скажуть, що маєш робити!
ACTS|9|7|А люди, що йшли з ним, онімілі стояли, бо вони чули голос, та нікого не бачили.
ACTS|9|8|Тоді Савл підвівся з землі, і хоч очі розплющені мав, нікого не бачив... І за руку його повели й привели до Дамаску.
ACTS|9|9|І три дні невидющий він був, і не їв, і не пив.
ACTS|9|10|А в Дамаску був учень один, на ймення Ананій. І Господь у видінні промовив до нього: Ананію! А він відказав: Ось я, Господи!
ACTS|9|11|Господь же до нього: Устань, і піди на вулицю, що Простою зветься, і пошукай в домі Юдовім Савла на ймення, тарсянина, ось бо він молиться,
ACTS|9|12|і мужа в видінні він бачив, на ймення Ананія, що до нього прийшов і руку на нього поклав, щоб став він видющий...
ACTS|9|13|Відповів же Ананій: Чув я, Господи, від багатьох про цього чоловіка, скільки зла він учинив в Єрусалимі святим Твоїм!
ACTS|9|14|І тут має владу від первосвящеників, щоб в'язати усіх, хто кличе Ім'я Твоє.
ACTS|9|15|І промовив до нього Господь: Іди, бо для Мене посудина вибрана він, щоб носити Ім'я Моє перед народами, і царями, і синами Ізраїля.
ACTS|9|16|Бо Я покажу йому, скільки має він витерпіти за Ім'я Моє.
ACTS|9|17|І Ананій пішов, і до дому ввійшов, і руки поклавши на нього, промовив: Савле брате, Господь Ісус, що з'явився тобі на дорозі, якою ти йшов, послав ось мене, щоб став ти видющий, і наповнився Духа Святого!
ACTS|9|18|І хвилі тієї відпала з очей йому ніби луска, і зараз видющий він став... І, вставши, охристився,
ACTS|9|19|і, прийнявши поживу, на силах зміцнів.
ACTS|9|20|І він зараз зачав у синагогах звіщати про Ісуса, що Він Божий Син,
ACTS|9|21|І дивом усі дивувалися, хто чув, і говорили: Хіба це не той, що переслідував в Єрусалимі визнавців оцього Ім'я, та й сюди не на те він прибув, щоб отих пов'язати й привести до первосвящеників?
ACTS|9|22|А Савл іще більше зміцнявся, і непокоїв юдеїв, що в Дамаску жили, удоводнюючи, що Той то Христос.
ACTS|9|23|А як часу минуло доволі, юдеї змовилися його вбити,
ACTS|9|24|та Савлові стала відома їхня змова. А вони день і ніч чатували в воротях, щоб убити його.
ACTS|9|25|Тому учні забрали його вночі, та й із муру спустили в коші.
ACTS|9|26|А коли він до Єрусалиму прибув, то силкувався пристати до учнів, та його всі лякалися, не вірячи, що він учень.
ACTS|9|27|Варнава тоді взяв його та й привів до апостолів, і їм розповів, як дорогою той бачив Господа, і як Він йому промовляв, і як сміливо навчав у Дамаску в Ісусове Ймення.
ACTS|9|28|І він із ними входив і виходив до Єрусалиму, і відважно звіщав в Ім'я Господа.
ACTS|9|29|Він також розмовляв й сперечався з огреченими, а вони намагалися вбити його.
ACTS|9|30|Тому браття, довідавшися, відвели його до Кесарії, і до Тарсу його відіслали.
ACTS|9|31|А Церква по всій Юдеї, і Галілеї, і Самарії мала мир, будуючись і ходячи в страсі Господньому, і сповнялася втіхою Духа Святого.
ACTS|9|32|І сталося, як Петро всіх обходив, то прибув і до святих, що мешкали в Лідді.
ACTS|9|33|Знайшов же він там чоловіка одного, на ймення Еней, що на ліжку лежав вісім років, він розслаблений був.
ACTS|9|34|І промовив до нього Петро: Енею, тебе вздоровляє Ісус Христос. Уставай, і постели собі сам! І той зараз устав...
ACTS|9|35|І його оглядали усі, хто мешкав у Лідді й Сароні, які навернулися до Господа.
ACTS|9|36|А в Йоппії була одна учениця, на ймення Тавіта, що в перекладі Сарною зветься. Вона повна була добрих вчинків та милостині, що чинила.
ACTS|9|37|І трапилося тими днями, що вона занедужала й умерла. Обмили ж її й поклали в горниці.
ACTS|9|38|А що Лідда лежить недалеко Йоппії, то учні, прочувши, що в ній пробуває Петро, послали до нього двох мужів, що благали: Не гайся прибути до нас!
ACTS|9|39|І, вставши Петро, пішов із ними. А коли він прибув, то ввели його в горницю. І обступили його всі вдовиці, плачучи та показуючи йому сукні й плащі, що їх Сарна робила, як із ними була.
ACTS|9|40|Петро ж із кімнати всіх випровадив, і, ставши навколішки, помолився, і, звернувшись до тіла, промовив: Тавіто, вставай! А вона свої очі розплющила, і сіла, уздрівши Петра...
ACTS|9|41|Він же руку подав їй, і підвів її, і закликав святих і вдовиць, та й поставив живою її.
ACTS|9|42|А це стало відоме по цілій Йоппії, і багато-хто в Господа ввірували.
ACTS|9|43|І сталось, що він багато днів пробув у Йоппії, в одного гарбарника Симона.
ACTS|10|1|Проживав же один чоловік у Кесарії, на ймення Корнилій, сотник полку, що звавсь Італійським.
ACTS|10|2|З усім домом своїм він побожний був та богобійний, подавав людям щедру милостиню, і завжди Богові молився.
ACTS|10|3|Явно він у видінні, десь коло години дев'ятої дня, бачив Ангола Божого, що до нього зійшов і промовив йому: Корнилію!
ACTS|10|4|Він поглянув на нього й жахнувся, й сказав: Що, Господи? Той же йому відказав: Молитви твої й твоя милостиня перед Богом згадалися.
ACTS|10|5|Тепер же пошли до Йоппії людей, та й приклич Симона, що зветься Петром.
ACTS|10|6|Він гостює в одного гарбарника Симона, що дім має при морі. Він скаже тобі, що ти маєш робити.
ACTS|10|7|Коли ж Ангол, що йому говорив, відійшов, той закликав двох із своїх слуг домових, і вояка богобійного з тих, що служили при ньому,
ACTS|10|8|і розповів їм усе та й послав їх в Йоппію.
ACTS|10|9|А наступного дня, як у дорозі були вони та наближались до міста, Петро вийшов на горницю, щоб помолитись, о годині десь шостій.
ACTS|10|10|І став він голодний, і їсти схотів. Як йому ж готували, захоплення на нього найшло,
ACTS|10|11|і бачить він небо відкрите, і якуюсь посудину, що сходила, немов простирало велике, яка, за чотири кінці прив'язана, спускалась додолу.
ACTS|10|12|У ній же знаходились чотириногі всілякі, і земне гаддя, і небесні пташки.
ACTS|10|13|І голос почувся до нього: Устань, заколи, Петре, і їж!
ACTS|10|14|А Петро відказав: Жадним способом, Господи, бо ніколи не їв я нічого огидного чи то нечистого!
ACTS|10|15|І знов голос удруге до нього: Що від Бога очищене, не вважай за огидне того!
ACTS|10|16|І це сталося тричі, і посудина знов була взята на небо.
ACTS|10|17|Як Петро ж у собі бентежився, що б то значило те видіння, що бачив, то ось посланці від Корнилія, розпитавши про Симонів дім, спинилися перед ворітьми,
ACTS|10|18|і спиталися, крикнувши: Чи то тут сидить Симон, що зветься Петро?
ACTS|10|19|Як Петро ж над видінням роздумував, Дух промовив до нього: Онде три чоловіки шукають тебе.
ACTS|10|20|Але встань і зійди, і піди з ними без жадного сумніву, бо то Я їх послав!
ACTS|10|21|І зійшовши Петро до тих мужів, промовив: Ось я той, що його ви шукаєте. З якої причини прийшли ви?
ACTS|10|22|А вони відказали: Сотник Корнилій, муж праведний та богобійний, слави доброї в усього люду юдейського, святим Анголом був у видінні наставлений, щоб до дому свого покликати тебе та послухати слів твоїх.
ACTS|10|23|Тоді він покликав й гостинно прийняв їх. А другого дня він устав та й із ними пішов; також дехто з братів із Йоппії пішли з ним.
ACTS|10|24|І назавтра прийшли вони до Кесарії. А Корнилій чекав їх, рідню й близьких друзів покликавши.
ACTS|10|25|А як увіходив Петро, Корнилій зустрінув його, і до ніг йому впав і вклонився.
ACTS|10|26|Та Петро його підвів, промовляючи: Устань, бо й сам я людина!
ACTS|10|27|І, розмовляючи з ним, увійшов, і знайшов багатьох, що зібралися,
ACTS|10|28|і промовив до них: Ви знаєте, що невільно юдеєві приставати й приходити до чужаниці. Та відкрив мені Бог, щоб я жадну людину не мав за огидну чи то за нечисту.
ACTS|10|29|Тому я без вагання прибув, як покликано. Тож питаю я вас: З якої причини ви слали по мене?
ACTS|10|30|А Корнилій сказав: Четвертого дня аж до цієї години я постив, а о дев'ятій годині молився я в домі своїм. І ото, перед мене став муж у блискучій одежі
ACTS|10|31|й сказав: Корнилію, почута молитва твоя, і твої милостині перед Богом згадалися.
ACTS|10|32|Тож пошли до Йоппії, і приклич Симона, що зветься Петром. Він гостює в гарбарника Симона, у господі край моря, він прийде й розповість тобі.
ACTS|10|33|Я зараз по тебе послав, ти добре зробив, що прийшов. Тож тепер перед Богом ми всі стоїмо, щоб почути все те, що Господь наказав був тобі.
ACTS|10|34|А Петро відкрив уста свої та й промовив: Пізнаю я поправді, що не дивиться Бог на обличчя,
ACTS|10|35|але в кожнім народі приємний Йому, хто боїться Його й чинить правду.
ACTS|10|36|Він слово послав для Ізраїлевих синів, благовістячи мир через Ісуса Христа, що Господь Він усім.
ACTS|10|37|Ви знаєте справу, що по всій Юдеї була й зачалась з Галілеї, після хрищення, що Іван проповідував,
ACTS|10|38|Ісуса, що був із Назарету, як помазав Його Святим Духом і силою Бог. І ходив Він, добро чинячи й усіх уздоровлюючи, кого поневолив диявол, бо Бог був із Ним.
ACTS|10|39|І ми свідки всьому, що Він учинив у Юдейському краї та в Єрусалимі, та вбили Його, на дереві повісивши...
ACTS|10|40|Але Бог воскресив Його третього дня, і дав Йому, щоб з'явився,
ACTS|10|41|не всьому народові, але наперед Богом вибраним свідкам, нам, що з Ним їли й пили, як воскрес Він із мертвих.
ACTS|10|42|І Він нам звелів, щоб народові ми проповідували та засвідчили, що то Він є призначений Богом Суддя для живих і для мертвих.
ACTS|10|43|Усі пророки свідкують про Нього, що кожен, хто вірує в Нього, одержить прощення гріхів Його Йменням.
ACTS|10|44|Як Петро говорив ще слова ці, злинув Святий Дух на всіх, хто слухав слова.
ACTS|10|45|А обрізані віруючі, що з Петром прибули, здивувалися дивом, що дар Духа Святого пролився також на поган!
ACTS|10|46|Бо чули вони, що мовами різними ті розмовляли та Бога звеличували... Петро тоді відповів:
ACTS|10|47|Чи хто може заборонити христитись водою оцим, що одержали Духа Святого, як і ми?
ACTS|10|48|І звелів охриститися їм у Ймення Ісуса Христа. Тоді просили його позостатися в них кілька днів.
ACTS|11|1|Почули ж апостоли й браття, що в Юдеї були, що й погани прийняли Слово Боже.
ACTS|11|2|І, як Петро повернувся до Єрусалиму, з ним стали змагатися ті, хто з обрізання,
ACTS|11|3|кажучи: Чого ти ходив до людей необрізаних та споживав із ними?
ACTS|11|4|Петро ж розпочав і їм розповів за порядком, говорячи:
ACTS|11|5|Був я в місті йоппійськім і молився, і бачив в захопленні видіння: якась посудина сходила, немов простирало велике, яка, за чотири кінці прив'язана, спускалася з неба й підійшла аж до мене.
ACTS|11|6|Зазирнувши до неї, я поглянув, і побачив там чотириногих землі, і звірів, і гаддя, і небесних пташок.
ACTS|11|7|І голос почув я, що мені промовляв: Устань, Петре, заколи та й їж!
ACTS|11|8|А я відказав: Жадним способом, Господи, бо ніколи нічого огидного чи то нечистого в уста мої не ввіходило!
ACTS|11|9|І відповів мені голос із неба вдруге: Що від Бога очищене, не вважай за огидне того!
ACTS|11|10|І це сталося тричі, і все знов було взяте на небо.
ACTS|11|11|І ось три чоловіки, посланці з Кесарії до мене, перед домом, де був я, спинилися зараз.
ACTS|11|12|І сказав мені Дух іти з ними без жадного сумніву. Зо мною ж пішли й оці шестеро браття, і ввійшли ми до дому того чоловіка.
ACTS|11|13|І він нам розповів, як у домі своїм бачив Ангола, який став і сказав: Пошли до Йоппії, та приклич того Симона, що зветься Петром,
ACTS|11|14|він слова тобі скаже, якими спасешся і ти, і ввесь дім твій.
ACTS|11|15|А як я промовляв, злинув на них Святий Дух, як спочатку й на нас.
ACTS|11|16|І я згадав слово Господнє, як Він говорив: Іван ось водою христив, ви ж охрищені будете Духом Святим.
ACTS|11|17|Отож, коли Бог дав однаковий дар їм, як і нам, що ввірували в Господа Ісуса Христа, то хто ж я такий, щоб міг заперечити Богові?
ACTS|11|18|І, почувши таке, замовкли вони, і Бога хвалили, говорячи: Отож, і поганам Бог дав покаяння в життя!
ACTS|11|19|А ті, хто розпорошився від переслідування, що знялося було через Степана, перейшли навіть до Фінікії, і Кіпру, і Антіохії, не звістуючи слова нікому, крім юдеїв.
ACTS|11|20|А між ними були мужі деякі з Кіпру та з Кірінеї, що до Антіохії прийшли, і промовляли й до греків, благовістячи про Господа Ісуса.
ACTS|11|21|І Господня рука була з ними; і велике число їх увірувало, і навернулось до Господа!
ACTS|11|22|І вістка про них досягла до вух єрусалимської Церкви, і до Антіохії послали Варнаву.
ACTS|11|23|А він, як прийшов і благодать Божу побачив, звеселився, і всіх став просити, щоб серцем рішучим трималися Господа.
ACTS|11|24|Бо він добрий був муж, повний Духа Святого та віри. І прилучилось багато народу до Господа!
ACTS|11|25|Після того подався Варнава до Тарсу, щоб Савла шукати.
ACTS|11|26|А знайшовши, привів в Антіохію. І збирались у Церкві вони цілий рік, і навчали багато народу, і в Антіохії найперш християнами названо учнів.
ACTS|11|27|Прибули ж тими днями пророки від Єрусалиму до Антіохії.
ACTS|11|28|І встав один з них, на ймення Агав, і Духом прорік, що голод великий у цілому світі настане, як за Клавдія був.
ACTS|11|29|Тоді учні, усякий із своєї спроможности, постановили послати допомогу братам, що в Юдеї жили.
ACTS|11|30|Що й зробили, через руки Варнави та Савла, пославши до старших.
ACTS|12|1|А Цар Ірод тоді підніс руки, щоб декого з Церкви гнобити.
ACTS|12|2|І мечем він стяв Якова, брата Іванового.
ACTS|12|3|А бачивши, що подобалося це юдеям, він задумав схопити й Петра. Були ж дні Опрісноків.
ACTS|12|4|І, схопивши його, посадив до в'язниці, і передав чотирьом чвіркам вояків, щоб його стерегли, бажаючи вивести людям його по Пасці.
ACTS|12|5|Отож, у в'язниці Петра стерегли, а Церква ревно молилася Богові за нього.
ACTS|12|6|А як Ірод хотів його вивести, Петро спав тієї ночі між двома вояками, закутий у два ланцюги, і сторожа пильнувала в'язницю при дверях.
ACTS|12|7|І ось Ангол Господній з'явився, і в в'язниці засяяло світло. І, доторкнувшись до боку Петрового, він збудив його, кажучи: Мерщій вставай! І ланцюги йому з рук поспадали.
ACTS|12|8|А Ангол до нього промовив: Підпережися, і взуй сандалі свої. І він так учинив. І каже йому: Зодягнися в плаща свого, та й за мною йди.
ACTS|12|9|І, вийшовши, він ішов услід за ним, і не знав, чи то правда, що робилось від Ангола, бо думав, що видіння він бачить.
ACTS|12|10|Як сторожу минули вони першу й другу, то прийшли до залізної брами, що до міста веде, і вона відчинилась сама їм. І, вийшовши, пройшли одну вулицю, і відступив Ангол зараз від нього.
ACTS|12|11|Сказав же Петро, опритомнівши: Тепер знаю правдиво, що Господь послав Свого Ангола, і видер мене із рук Іродових та від усього чекання народу юдейського.
ACTS|12|12|А зміркувавши, він прийшов до садиби Марії, матері Івана, званого Марком, де багато зібралося й молилося.
ACTS|12|13|І як Петро в фіртку брами постукав, то вийшла послухати служниця, що звалася Рода,
ACTS|12|14|та голос Петрів розпізнавши, вона з радощів не відчинила воріт, а прибігши, сказала, що Петро при воротях стоїть!...
ACTS|12|15|А вони їй сказали: Чи ти навісна? Та вона запевняла своє, що є так. Вони ж говорили: То Ангол його!
ACTS|12|16|А Петро й далі стукав. Коли ж відчинили, вони його вгледіли та й дивувалися.
ACTS|12|17|Махнувши ж рукою до них, щоб мовчали, він їм розповів, як Господь його вивів із в'язниці. І сказав: Сповістіть про це Якова й браттю. І, вийшовши, він до іншого місця пішов.
ACTS|12|18|Коли ж настав день, поміж вояками зчинилась велика тривога, що то сталось з Петром.
ACTS|12|19|А Ірод, пошукавши його й не знайшовши, віддав варту під суд, і звелів їх стратити. А сам із Юдеї відбув в Кесарію, і там перебував.
ACTS|12|20|А Ірод розгніваний був на тирян та сидонян. І вони однодушно до нього прийшли, і вблагали царського постельника Власта, та й миру просили, бо їхня земля годувалась з царської.
ACTS|12|21|Дня ж призначеного Ірод убрався в одежу царську, і на підвищенні сів та й до них говорив.
ACTS|12|22|А натовп кричав: Голос Божий, а не людський!
ACTS|12|23|І Ангол Господній уразив зненацька його, бо він не віддав слави Богові. І черва його з'їла, і він умер...
ACTS|12|24|Слово ж Боже росло та помножувалось.
ACTS|12|25|А Варнава та Савл, службу виконавши, повернулись із Єрусалиму, узявши з собою Івана, що прозваний Марком.
ACTS|13|1|А в Антіохії, у тамошній Церкві були ці пророки та вчителі: Варнава й Семен, званий Ніґер, і кірінеянин Луцій, і Манаїл, що був вигодуваний із тетрархом Іродом, та ще Савл.
ACTS|13|2|Як служили ж вони Господеві та постили, прорік Святий Дух: Відділіть Варнаву та Савла для Мене на справу, до якої покликав Я їх!
ACTS|13|3|Тоді, попостивши та помолившись, вони руки поклали на них, і відпустили.
ACTS|13|4|Вони ж, послані бувши від Духа Святого, прийшли в Селевкію, а звідти до Кіпру відплинули.
ACTS|13|5|Як були ж в Саламіні, то звіщали вони Слово Боже по синагогах юдейських; до послуг же мали й Івана.
ACTS|13|6|А коли перейшли аж до Пафи ввесь острів, то знайшли ворожбита одного, лжепророка юдеянина, йому на ім'я Варісус.
ACTS|13|7|Він був при проконсулі Сергії Павлі, чоловіку розумнім. Той закликав Варнаву та Савла, і прагнув послухати Божого Слова.
ACTS|13|8|Але їм опирався Еліма ворожбит той, бо ім'я його перекладається так, і намагавсь відвернути від віри проконсула.
ACTS|13|9|Але Савл, що й Павло він, переповнився Духом Святим і на нього споглянув,
ACTS|13|10|і промовив: О сину дияволів, повний всякого підступу та всілякої злости, ти ворогу всякої правди! Чи не перестанеш ти плутати простих Господніх доріг?
ACTS|13|11|І тепер ось на тебе Господня рука, ти станеш сліпий, і сонця бачити не будеш до часу! І миттю обняв того морок та темрява, і став він ходити навпомацки та шукати поводатора...
ACTS|13|12|Тоді той проконсул, як побачив, що сталося, увірував, і дивувався науці Господній!
ACTS|13|13|І, як від Пафа Павло й ті, хто з ним був, відпливли, то вони прибули в Памфілійську Пергію. А Іван, відлучившись від них, повернувся до Єрусалиму.
ACTS|13|14|А вони, пішовши з Пергії, прийшли до Пісідійської Антіохії, і дня суботнього до синагоги ввійшли й посідали.
ACTS|13|15|А по відчитанні Закону й Пророків, старші синагоги послали до них, переказуючи: Мужі-браття, якщо маєте слово потіхи для люду, промовте!
ACTS|13|16|Тоді Павло встав, і давши знака рукою, промовив: Послухайте, мужі ізраїльтяни, та ви, богобійні!
ACTS|13|17|Бог цих Ізраїлевих людей вибрав Собі отців наших, і підвищив народ, як він перебував у єгипетськім краї, і рукою потужною вивів їх із нього,
ACTS|13|18|і літ із сорок Він їх годував у пустині,
ACTS|13|19|а вигубивши сім народів в землі ханаанській, поділив жеребком їхню землю між ними,
ACTS|13|20|майже що по чотириста й п'ятидесяти роках. Після того аж до Самуїла пророка Він їм суддів давав.
ACTS|13|21|А потім забажали царя, і Бог дав їм Саула, сина Кісового, мужа з Веніяминового племени, на чотири десятки років.
ACTS|13|22|А його віддаливши, поставив царем їм Давида, про якого й сказав, засвідчуючи: Знайшов Я Давида, сина Єссеєвого, чоловіка за серцем Своїм, що всю волю Мою він виконувати буде.
ACTS|13|23|За обітницею, із його насіння підняв Бог Ісуса, як спасіння Ізраїлеві,
ACTS|13|24|як Іван перед самим приходом Його усьому народові Ізраїлевому проповідував хрищення на покаяння.
ACTS|13|25|А коли свою путь Іван виконав, то він промовляв: Я не Той, за Кого ви мене вважаєте, але йде он за мною, що Йому розв'язати ремінця від узуття Його я недостойний.
ACTS|13|26|Мужі-браття, сини роду Авраамового, та хто богобоязний із вас! Для вас було послане слово спасіння цього.
ACTS|13|27|Бо мешканці Єрусалиму та їхня старшина Його не пізнали, а пророчі слова які щосуботи читаються вони сповнили присудом,
ACTS|13|28|і хоч жадної провини смертельної в Ісусі вони не знайшли, все ж просили Пилата вбити Його.
ACTS|13|29|Коли ж усе виповнилось, що про Нього написане, то зняли Його з дерева, та й до гробу поклали.
ACTS|13|30|Але Бог воскресив Його з мертвих!
ACTS|13|31|Він з'являвся багато днів тим, що були поприходили з Ним із Галілеї до Єрусалиму, і що тепер вони свідки Його перед людьми.
ACTS|13|32|І ми благовістимо вам ту обітницю, що дана була нашим отцям,
ACTS|13|33|що її нам, їхнім дітям, Бог виконав, воскресивши Ісуса, як написано в другім псалмі: Ти Мій Син, Я сьогодні Тебе породив!
ACTS|13|34|А що Він воскресив Його з мертвих, щоб більш не вернувся в зотління, те так заповів: Я дам вам ті милості, що обіцяні вірно Давиду були!
ACTS|13|35|Тому то й деінде говорить: Не даси Ти Своєму Святому побачити тління!
ACTS|13|36|Бо Давид, що часу свого послужив волі Божій, спочив, і злучився з отцями своїми, і тління побачив.
ACTS|13|37|Але Той, що Бог воскресив Його з мертвих, тління не побачив.
ACTS|13|38|Отже, мужі-браття, хай відомо вам буде, що прощення гріхів через Нього звіщається вам.
ACTS|13|39|І в усім, у чому ви не могли виправдатись Законом Мойсеєвим, через Нього виправдується кожен віруючий.
ACTS|13|40|Отож, стережіться, щоб на вас не прийшло, що в Пророків провіщене:
ACTS|13|41|Дивіться, погордющі, і дивуйтеся та пощезайте, бо Я діло роблю за днів ваших, те діло, що йому не повірите ви, якби хто розповів вам!
ACTS|13|42|А як стали виходити вони, то їх прошено, щоб на другу суботу до них говорили ті самі слова.
ACTS|13|43|А коли розійшлась синагога, то багато з юдеїв та й із нововірців побожних пішли за Павлом та Варнавою, а вони промовляли до них і намовляли їх перебувати в благодаті Божій.
ACTS|13|44|А в наступну суботу зібралося майже все місто послухати Божого Слова.
ACTS|13|45|Як юдеї ж побачили натовп, то наповнились заздрощів, і стали перечити мові Павла та богозневажати.
ACTS|13|46|Тоді Павло та Варнава мужньо промовили: До вас перших потрібно було говорить Слово Боже; та коли ви його відкидаєте, а себе вважаєте за недостойних вічного життя, то ось до поган ми звертаємось.
ACTS|13|47|Бо так заповів нам Господь: Я світлом поставив Тебе для поган, щоб спасінням Ти був аж до краю землі!
ACTS|13|48|А погани, почувши таке, раділи та Слово Господнє хвалили. І всі ті, хто призначений був в життя вічне, увірували.
ACTS|13|49|І ширилось Слово Господнє по цілій країні.
ACTS|13|50|Юдеї ж підбили побожних впливових жінок та значніших у місті, і зняли переслідування на Павла та Варнаву, та й вигнали їх із своєї землі.
ACTS|13|51|Вони ж, обтрусивши із ніг своїх порох на них, подалися в Іконію.
ACTS|13|52|А учні сповнялися радощів і Духа Святого.
ACTS|14|1|І трапилось, що в Іконії вкупі ввійшли вони до синагоги юдейської, і промовили так, що безліч юдеїв й огречених увірували.
ACTS|14|2|Невірні ж юдеї підбурили та роз'ятрили душі поган на братів.
ACTS|14|3|Та проте довгий час пробули вони там, промовляючи мужньо про Господа, що свідоцтво давав слову благодаті Своєї, і робив, щоб знамена та чуда чинились їхніми руками.
ACTS|14|4|А в місті народ поділився, і пристали одні до юдеїв, а інші тримались апостолів.
ACTS|14|5|Коли ж кинулися ті погани й юдеї з своїми старшими, щоб зневажити їх та камінням побити,
ACTS|14|6|то, дізнавшись про це, вони повтікали до міст лікаонських, до Лістри та Дервії, та в околиці їхні,
ACTS|14|7|і Євангелію там звіщали.
ACTS|14|8|А в Лістрі сидів один чоловік, безвладний на ноги, що кривий був з утроби своєї матері, і ніколи ходити не міг.
ACTS|14|9|Він слухав, як Павло говорив, який пильно на нього споглянув, і побачив, що має він віру вздоровленим бути,
ACTS|14|10|то голосом гучним промовив: Устань просто на ноги свої! А той скочив, і ходити почав...
ACTS|14|11|А люди, побачивши, що Павло вчинив, піднесли свій голос, говорячи по-лікаонському: Боги людям вподібнились, та до нас ось зійшли!...
ACTS|14|12|І Варнаву вони звали Зевсом, а Гермесом Павла, бо він провід мав у слові.
ACTS|14|13|А жрець Зевса, що святиня його перед містом була, припровадив бики та вінки до воріт, та й з народом приносити жертву хотів.
ACTS|14|14|Та коли про це почули апостоли Варнава й Павло, то роздерли одежі свої, та й кинулися між народ, кричачи
ACTS|14|15|та говорячи: Що це робите, люди? Таж і ми такі самі смертельні, подібні вам люди, і благовістимо вам, від оцих ось марнот навернутись до Бога Живого, що створив небо й землю, і море, і все, що в них є.
ACTS|14|16|За минулих родів попустив Він усім народам, щоб ходили стежками своїми,
ACTS|14|17|але не зоставив Себе Він без свідчення, добро чинячи: подавав нам із неба дощі та врожайні часи, та наповнював їжею й радощами серця наші.
ACTS|14|18|І, говорячи це, заледве спинили народ не приносити їм жертов.
ACTS|14|19|А з Антіохії та з Іконії посходились юдеї, і, підбуривши натовп, камінням побили Павла, та й за місто геть виволікли, мавши думку, що вмер він...
ACTS|14|20|Коли ж учні його оточили, то він устав, та й вернувся до міста. А наступного дня він відбув із Варнавою в Дервію.
ACTS|14|21|І, як звістили Євангелію тому містові, і учнів багато придбали, вони повернулися в Лістру, та в Іконію, та в Антіохію,
ACTS|14|22|душі учнів зміцняючи, просячи перебувати в вірі, та навчаючи, що через великі утиски треба нам входити у Боже Царство.
ACTS|14|23|І рукопоклали їм пресвітерів по Церквах, і помолилися з постом та й їх передали Господеві, в Якого ввірували.
ACTS|14|24|Як вони ж перейшли Пісідію, прибули в Памфілію;
ACTS|14|25|і, звістивши Господнє Слово в Пергії, вони в Атталію ввійшли,
ACTS|14|26|а звідти поплинули в Антіохію, звідки були благодаті Божій віддані на діло, що його й закінчили.
ACTS|14|27|А прибувши та скликавши Церкву, вони розповіли, як багато вчинив Бог із ними, і що відкрив двері і віри поганам.
ACTS|14|28|І перебували вони немалий час із учнями.
ACTS|15|1|А дехто, що з Юдеї прийшли, навчали братів: Якщо ви не обріжетеся за звичаєм Мойсеєвим, то спастися не можете.
ACTS|15|2|Коли ж суперечка повстала й чимале змагання в Павла та в Варнави з ними, то постановили, щоб Павло та Варнава, та дехто ще інший із них, пішли в справі цій до апостолів й старших у Єрусалим.
ACTS|15|3|Тож вони, відпроваджені Церквою, ішли через Фінікію та Самарію, розповідуючи про поганське навернення, і радість велику чинили всім браттям.
ACTS|15|4|Коли ж в Єрусалим прибули вони, були прийняті Церквою, та апостолами, та старшими, і вони розповіли, як багато вчинив Бог із ними.
ACTS|15|5|Але дехто, що ввірували з фарисейської партії, устали й сказали, що потрібно поганів обрізувати й наказати, щоб Закона Мойсеєвого берегли.
ACTS|15|6|І зібрались апостоли й старші, щоб розглянути справу оцю.
ACTS|15|7|Як велике ж змагання повстало, Петро встав і промовив до них: Мужі-браття, ви знаєте, що з давнішніх днів вибрав Бог поміж нами мене, щоб погани почули слово Євангелії через уста мої, та й увірували.
ACTS|15|8|І засвідчив їм Бог Серцезнавець, давши їм Духа Святого, як і нам,
ACTS|15|9|і між нами та ними різниці Він жадної не вчинив, очистивши вірою їхні серця.
ACTS|15|10|Отож, чого Бога тепер спокушуєте, щоб учням на шию покласти ярмо, якого ані наші отці, ані ми не здолали понести?
ACTS|15|11|Та ми віруємо, що спасемося благодаттю Господа Ісуса так само, як і вони.
ACTS|15|12|І вся громада замовкла, і слухали пильно Варнаву й Павла, що розповідали, які то знамена та чуда вчинив через них Бог між поганами!
ACTS|15|13|Як замовкли ж вони, то Яків озвався й промовив: Мужі-браття, послухайте також мене.
ACTS|15|14|Симон ось розповів, як зглянувся Бог від початку, щоб вибрати люд із поганів для Ймення Свого.
ACTS|15|15|І пророчі слова з цим погоджуються, як написано:
ACTS|15|16|Потому вернуся, і відбудую Давидову скинію занепалу, і відбудую руїни її, і наново поставлю її,
ACTS|15|17|щоб шукали Господа люди зосталі та всі народи, над якими Ім'я Моє кликано, говорить Господь, що чинить це все!
ACTS|15|18|Господеві відвіку відомі всі вчинки Його.
ACTS|15|19|Тому думаю я, щоб не турбувати поган, що до Бога навертаються,
ACTS|15|20|але написати до них, щоб стримувались від занечищення ідольського, та від блуду, і задушенини, і від крови.
ACTS|15|21|Бо своїх проповідників має Мойсей по містах здавендавна, і щосуботи читають його в синагогах.
ACTS|15|22|Тоді постановили апостоли й старші з цілою Церквою вибрати мужів із них, і послати до Антіохії з Павлом та Варнавою Юду, що зветься Варсавва, і Силу, мужів проводирів між братами,
ACTS|15|23|написавши своїми руками оце: Апостоли й старші брати до братів, що з поган в Антіохії, і Сирії, і Кілікії: Вітаємо вас!
ACTS|15|24|Через те, що ми чули, що деякі з вас, яким ми того не доручували, стурбували наукою вас, і захитали вам душі,
ACTS|15|25|то ми постановили однодушно, зібравшися, щоб обраних мужів послати до вас із коханими нашими Варнавою та Павлом,
ACTS|15|26|людьми тими, що душі свої віддали за Ім'я Господа нашого Ісуса Христа.
ACTS|15|27|Тож ми Юду та Силу послали, що вияснять усно те саме.
ACTS|15|28|Бо зволилось Духові Святому і нам, тягару вже ніякого не накладати на вас, окрім цього необхідного:
ACTS|15|29|стримуватися від ідольських жертов та крови, і задушенини, та від блуду. Оберегаючися від того, ви зробите добре. Бувайте здорові!...
ACTS|15|30|Посланці ж прийшли в Антіохію, і, зібравши народ, доручили листа.
ACTS|15|31|А перечитавши, раділи з потішення того.
ACTS|15|32|А Юда та Сила, самі бувши пророками, частим словом підбадьорували та зміцняли братів.
ACTS|15|33|А як перебули вони там якийсь час, то брати їх відпустили з миром до тих, хто їх вислав.
ACTS|15|34|Але Сила схотів лишитися там, а Юда вернувся до Єрусалиму.
ACTS|15|35|А Павло з Варнавою в Антіохії жили, навчаючи та благовістячи разом із іншими багатьома Слово Господнє.
ACTS|15|36|А по декількох днях промовив Павло до Варнави: Ходімо знов, і відвідаймо наших братів у кожному місті, де ми провіщали Слово Господнє, як вони пробувають.
ACTS|15|37|А Варнава хотів був узяти з собою Івана, що званий був Марком.
ACTS|15|38|Та Павло вважав за потрібне не брати з собою того, хто від них відлучився з Памфілії, та з ними на працю не йшов.
ACTS|15|39|І повстала незгода, і розлучились вони між собою. Тож Варнава взяв Марка, і поплинув до Кіпру.
ACTS|15|40|А Павло вибрав Силу й пішов, Божій благодаті братами доручений.
ACTS|15|41|І проходив він Сирію та Кілікію, Церкви зміцнюючи.
ACTS|16|1|І прибув він у Дервію й Лістру. І ото був там один учень, на ім'я Тимофій, син наверненої однієї юдеянки, а батько був геллен.
ACTS|16|2|Добре свідоцтво про нього давали брати, що були в Лістрі та в Іконії.
ACTS|16|3|Павло захотів його взяти з собою, і, взявши, обрізав його через юдеїв, що були в тих місцях, бо всі знали про батька його, що був геллен.
ACTS|16|4|Як міста ж переходили, то їм передавали, щоб вони берегли оті постанови, які видали в Єрусалимі апостоли та старші.
ACTS|16|5|А Церкви зміцнювалися в вірі, і щоденно зростали кількістю.
ACTS|16|6|А що Дух Святий їм не звелів провіщати слово в Азії, то вони перейшли через Фрігію та через країну галатську.
ACTS|16|7|Дійшовши ж до Мізії, хотіли піти до Вітінії, та їм не дозволив Дух Ісусів.
ACTS|16|8|Обминувши ж Мізію, прибули до Троади.
ACTS|16|9|І Павлові з'явилось видіння вночі: якийсь македонянин став перед ним і благав його, кажучи: Прийди в Македонію, і нам поможи!
ACTS|16|10|Як побачив він це видіння, то ми зараз хотіли піти в Македонію, зрозумівши, що Господь нас покликав звіщати їм Євангелію.
ACTS|16|11|Тож відпливши з Троади, прибули ми навпрост у Самотракію, а другого дня до Неаполя,
ACTS|16|12|звідтіля ж у Филипи, що є перше місто-осада в тій частині Македонії. І пробули ми в цім місті днів кілька.
ACTS|16|13|Дня ж суботнього вийшли ми з міста над річку, де, за звичаєм, було місце молитви, і, посідавши, розмовляли з жінками, що посходились.
ACTS|16|14|Прислухалася й жінка одна, що звалася Лідія, купчиха кармазином з міста Тіятір, що Бога вона шанувала. Господь же їй серце відкрив, щоб уважати на те, що Павло говорив.
ACTS|16|15|А коли охристилась вона й її дім, то благала нас, кажучи: Якщо ви признали, що вірна я Господеві, то прийдіть до господи моєї й живіть. І змусила нас.
ACTS|16|16|І сталось, як ми йшли на молитву, то нас перестріла служниця одна, що мала віщунського духа, яка ворожбитством давала великий прибуток панам своїм.
ACTS|16|17|Вона йшла слідкома за Павлом та за нами, і кричала, говорячи: Оці люди це раби Всевишнього Бога, що вам провіщають дорогу спасіння!
ACTS|16|18|І багато днів вона це робила. І обуривсь Павло, і, обернувшись, промовив до духа: У Ім'я Ісуса Христа велю я тобі вийди з неї! І того часу той вийшов.
ACTS|16|19|А пани її, бачивши, що пропала надія на їхній прибуток, схопили Павла й Силу, і потягли їх на ринок до старших.
ACTS|16|20|Коли ж їх привели до начальників, то сказали: Ці люди, юдеї, наше місто бунтують,
ACTS|16|21|і навчають звичаїв, яких нам, римлянам, не годиться приймати, ані виконувати.
ACTS|16|22|І натовп піднявся на них. А начальники здерли одежу із них, та звеліли їх різками сікти.
ACTS|16|23|І, завдавши багато їм ран, посадили в в'язницю, наказавши в'язничному дозорцеві, щоб їх пильно стеріг.
ACTS|16|24|Одержавши такого наказа, той їх повкидав до внутрішньої в'язниці, а їхні ноги забив у колоди.
ACTS|16|25|А північної пори Павло й Сила молилися, і Богові співали, а ув'язнені слухали їх.
ACTS|16|26|І ось нагло повстало велике трясіння землі, аж основи в'язничні були захиталися! І повідчинялися зараз усі двері, а кайдани з усіх поспадали...
ACTS|16|27|Як прокинувся ж сторож в'язничний, і побачив відчинені двері в'язниці, то витяг меча та й хотів себе вбити, мавши думку, що повтікали ув'язнені.
ACTS|16|28|А Павло скрикнув голосом гучним, говорячи: Не чини собі жодного зла, бо всі ми ось тут!
ACTS|16|29|Зажадавши ж той світла, ускочив, і тремтячий припав до Павла та до Сили.
ACTS|16|30|І вивів їх звідти й спитав: Добродії! Що треба робити мені, щоб спастися?
ACTS|16|31|А вони відказали: Віруй в Господа Ісуса, і будеш спасений ти сам та твій дім.
ACTS|16|32|І Слово Господнє звіщали йому та й усім, хто був у домі його.
ACTS|16|33|І сторож забрав їх того ж часу вночі, їхні рани обмив, і охристився негайно він сам та його всі домашні.
ACTS|16|34|І він їх запровадив до дому свого, і поживу поставив, і радів із усім домом своїм, що ввірував у Бога.
ACTS|16|35|А коли настав день, то прислали начальники слуг поліційних, наказуючи: Відпусти тих людей!
ACTS|16|36|І сказав той в'язничний дозорець слова ці Павлові: що прислали начальники, щоб вас відпустити. Отож, вийдіть тепер та й з миром ідіть!
ACTS|16|37|А Павло відказав їм: Нас, римлян, незасуджених, різками сікли прилюдно, і до в'язниці всадили, а тепер нас таємно виводять? Але ні! Хай вони самі прийдуть, та й виведуть нас!
ACTS|16|38|Ці ж слова поліційні слуги донесли начальникам. А ті налякались, почувши, що римляни вони.
ACTS|16|39|І прийшли, та їх перепросили, а вивівши, благали, щоб із міста пішли.
ACTS|16|40|І, вийшовши з в'язниці, прибули вони до Лідії, а з братами побачившись, потішили їх та й пішли.
ACTS|17|1|Як вони перейшли Амфіполь й Аполлонію, то прийшли до Солуня, де була синагога юдейська.
ACTS|17|2|І Павло, за звичаєм своїм, до них увійшов, і з ними змагавсь три суботі з Писання,
ACTS|17|3|виказуючи та доводячи, що мусів Христос постраждати й воскреснути з мертвих, і що Христос Той Ісус, про Якого я вам проповідую.
ACTS|17|4|І ввірували дехто з них і до Павла та до Сили пристали, безліч побожних із гелленів та немало з шляхетних жінок.
ACTS|17|5|А невірні юдеї були запалилися заздрістю, і якихсь негідних людей назбирали на вулицях, учинили збіговисько та й бунтували те місто, а набігши на хату Ясонову, шукали апостолів, щоб до натовпу вивести їх.
ACTS|17|6|А як їх не знайшли, потягли до начальників міста Ясона та декого з братті, кричачи: Ті, що світ сколотили, і сюди ось вони поприходили!
ACTS|17|7|А Ясон їх до себе прийняв. Вони всі проти наказів кесаря чинять, говорячи, ніби інший є цар Ісус...
ACTS|17|8|І вони зворохобили народ та начальників міста, що слухали це.
ACTS|17|9|Але, узявши поруку з Ясона та з інших, вони їх відпустили.
ACTS|17|10|А брати відіслали негайно вночі Павла й Силу до Верії. І, прибувши вони, пішли в синагогу юдейську.
ACTS|17|11|Ці були шляхетніші за солунян, і слова прийняли з повним запалом, і Писання досліджували день-у-день, чи так воно є.
ACTS|17|12|Тож багато із них тоді ввірували, і з почесних гелленських жінок та немало із мужів.
ACTS|17|13|Як солунські ж юдеї довідалися, що Павло проповідує Боже Слово й у Верії, прибули вони, і там баламутили та бунтували народ.
ACTS|17|14|Тоді браття негайно Павла відпустили, щоб до моря йшов; а Сила та Тимофій позосталися там.
ACTS|17|15|А ті, що Павла відпроваджували, провели його аж до Атен, а прийнявши наказа про Силу та Тимофія, щоб до нього вернулися якнайшвидше, відбули.
ACTS|17|16|Як Павло ж їх чекав ув Атенах, у ньому кипів його дух, як бачив це місто, повне ідолів.
ACTS|17|17|Тож він розмовляв у синагозі з юдеями та з богобійними, і на ринку щоденно зо стрічними.
ACTS|17|18|А дехто з філософів епікуреїв та стоїків сперечалися з ним. Одні говорили: Що то хоче сказати оцей пустомов? А інші: Здається, він проповідник чужих богів, бо він їм звіщав Євангелію про Ісуса й воскресення.
ACTS|17|19|І, взявши його, повели в ареопаг та й казали: Чи можемо знати, що то є ця наука нова, яку проповідуєш ти?
ACTS|17|20|Бо чудне щось вкладаєш до наших вух. Отже хочемо знати, що то значити має?
ACTS|17|21|А всі атеняни та захожі чужинці нічим іншим радніш не займалися, як аби щось нове говорити чи слухати.
ACTS|17|22|Тоді Павло став посередині ареопагу й промовив: Мужі атенські! Із усього я бачу, що ви дуже побожні.
ACTS|17|23|Бо, проходячи та оглядаючи святощі ваші, я знайшов також жертівника, що на ньому написано: Незнаному Богові. Ось Того, Кого навмання ви шануєте, Того я проповідую вам.
ACTS|17|24|Бог, що створив світ і все, що в ньому, бувши Господом неба й землі, проживає не в храмах, рукою збудованих,
ACTS|17|25|і Він не вимагає служіння рук людських, ніби в чомусь Він мав би потребу, бо Сам дає всім і життя, і дихання, і все.
ACTS|17|26|І ввесь людський рід Він з одного створив, щоб замешкати всю поверхню землі, і призначив окреслені доби й границі замешкання їх,
ACTS|17|27|щоб Бога шукали вони, чи Його не відчують і не знайдуть, хоч Він недалеко від кожного з нас.
ACTS|17|28|Бо ми в Нім живемо, і рухаємось, і існуємо, як і деякі з ваших поетів казали: Навіть рід ми Його!
ACTS|17|29|Отож, бувши Божим тим родом, не повинні ми думати, що Божество подібне до золота, або срібла, чи до каменю, твору мистецтва чи людської вигадки.
ACTS|17|30|Не зважаючи ж Бог на часи невідомости, ось тепер усім людям наказує, щоб скрізь каялися,
ACTS|17|31|бо Він визначив день, коли хоче судити поправді ввесь світ через Мужа, що Його наперед Він поставив, і Він подав доказа всім, із мертвих Його воскресивши.
ACTS|17|32|Як почули ж вони про воскресення мертвих, то одні насміхатися стали, а інші казали: Про це будемо слухати тебе іншим разом...
ACTS|17|33|Так вийшов Павло з-поміж них.
ACTS|17|34|А деякі мужі пристали до нього й увірували, серед них і Діонисій Ареопагіт, і жінка, Дамара ім'ям, та інші із ними.
ACTS|18|1|Після цього він вийшов з Атен і прибув до Коринту.
ACTS|18|2|І знайшов він одного юдея, на ймення Акилу, родом із Понту, що недавно прибув із Італії, та Прискиллу, його дружину, бо Клавдій звелів усім юдеям, щоб покинули Рим. І до них він прийшов,
ACTS|18|3|а що був він того ж ремесла, то в них позостався та працював; ремесло ж їхнє було виробляти намети.
ACTS|18|4|І він щосуботи розмову точив у синагозі, переконуючи юдеїв та гелленів.
ACTS|18|5|А коли прибули Сила та Тимофій з Македонії, Павло слову віддався, і він свідчив юдеям, що Ісус то Христос.
ACTS|18|6|Як вони ж спротивлялися та богозневажали, то він обтрусив одежу свою та промовив до них: Ваша кров на голову вашу! Я чистий. Відтепер я піду до поган.
ACTS|18|7|І, вийшовши звідти, він прибув до господи одного, на ім'я Тита Юста, що був богобійний, його ж дім межував із синагогою.
ACTS|18|8|А Крисп, старший синагоги, увірував в Господа з усім домом своїм; і багато з коринтян, почувши, увірували й охристились.
ACTS|18|9|Сказав же Павлові Господь у видінні вночі: Не бійся, але говори й не мовчи,
ACTS|18|10|бо з тобою ось Я, і на тебе ніхто не накинеться, щоб тобі заподіяти зло, бо Я маю в цім місті багато людей.
ACTS|18|11|І позостався він рік і шість місяців, навчаючи в них Слова Божого.
ACTS|18|12|А коли Галліон був в Ахаї проконсулом, то проти Павла однодушно повстали юдеї, і на суд привели його,
ACTS|18|13|кажучи: Цей людей намовляє, щоб Богові честь віддавали незгідно з Законом!
ACTS|18|14|Як Павло ж хотів уста відкрити, сказав Галліон до юдеїв: О юдеї, якби сталася кривда яка, або злий учинок, то я б справедливо вас вислухав.
ACTS|18|15|Та коли спір іде про слово та ймення й Закон ваш, то самі доглядайте, я суддею цього бути не хочу.
ACTS|18|16|І прогнав їх від суду.
ACTS|18|17|Тоді всі схопили Состена, начальника над синагогою, та й перед судом його били. Галліон же на те зовсім не зважав.
ACTS|18|18|А Павло, перебувши доволі ще днів, попрощався з братами, і поплинув у Сирію, і з ним Прискилла й Акила; він у Кенхреях обстриг собі голову, бо обітницю дав був.
ACTS|18|19|І прибув він в Ефес, і там їх позоставив, а сам у синагогу ввійшов і розмовляв із юдеями.
ACTS|18|20|Як просили ж його довший час позостатися в них, то він не згодився,
ACTS|18|21|але попрощався й сказав: Знов вернуся до вас, коли буде на те воля Божа! І відплив із Ефесу.
ACTS|18|22|І, побувши в Кесарії, він піднявся, і, привіт славши Церкві, відбув в Антіохію.
ACTS|18|23|І, пробувши там деякий час, він вибрався в подорож знову, за порядком проходячи через країну галатську та Фріґію, та всіх учнів зміцняючи.
ACTS|18|24|Один же юдей, на ім'я Аполлос, родом з Олександрії, красномовець та сильний в Писанні, прибув до Ефесу.
ACTS|18|25|Він був навчений дороги Господньої, і, палаючи духом, промовляв і про Господа пильно навчав, знаючи тільки Іванове хрищення.
ACTS|18|26|І він сміливо став промовляти в синагозі. Як Акила й Прискилла почули його, то його прийняли, і докладніш розповіли йому про дорогу Господню.
ACTS|18|27|А коли він схотів перейти до Ахаї, брати написали до учнів, нагадуючи, щоб його прийняли. А прибувши, помагав він багато тим, хто ввірував благодаттю,
ACTS|18|28|бо він переконував пильно юдеїв, Писанням прилюдно доводячи, що Ісус то Христос.
ACTS|19|1|І сталося, що коли Аполлос перебував у Коринті, то Павло, перейшовши горішні країни, прибув до Ефесу, і деяких учнів знайшов,
ACTS|19|2|та й спитав їх: Чи ви Духа Святого одержали, як увірували? А вони відказали йому: Та ми навіть не чули, чи є Дух Святий!
ACTS|19|3|І він запитав: Тож у що ви христились? Вони ж відказали: В Іванове хрищення.
ACTS|19|4|І промовив Павло: Таж Іван христив хрищенням на покаяння, говорячи людям, щоб вірили в Того, Хто прийде по ньому, цебто в Ісуса.
ACTS|19|5|Як почули ж оце, то христились вони в Ім'я Господа Ісуса.
ACTS|19|6|А коли Павло руки на них поклав, то зійшов на них Дух Святий, і різними мовами стали вони промовляти та пророкувати!
ACTS|19|7|А всіх їх було чоловіка з дванадцять.
ACTS|19|8|А до синагоги ввійшовши, промовляв він відважно, три місяці про Боже Царство навчаючи та переконуючи.
ACTS|19|9|А коли опиралися дехто й не вірували, і дорогу Господню лихословили перед народом, то він їх покинув і виділив учнів, і щодня проповідував у школі одного Тирана.
ACTS|19|10|Це ж два роки продовжувалось, так що всі, хто замешкував в Азії, юдеї та геллени, слухали слово про Господа.
ACTS|19|11|І Бог чуда чинив надзвичайні руками Павловими,
ACTS|19|12|так що навіть хустки й пояси з його тіла приносили хворим, і хвороби їх кидали, і духи лукаві виходили з них.
ACTS|19|13|Дехто ж із мандрівних ворожбитів юдейських зачали закликати Ім'я Господа Ісуса над тими, хто мав злих духів, проказуючи: Заклинаємо вас Ісусом, Якого Павло проповідує!
ACTS|19|14|Це ж робили якісь сім синів юдейського первосвященика Скеви.
ACTS|19|15|Відповів же злий дух і сказав їм: Я знаю Ісуса, і знаю Павла, а ви хто такі?
ACTS|19|16|І скочив на них чоловік, що в ньому злий дух був, і, перемігши обох, подужав їх так, що втекли вони з дому нагі та поранені.
ACTS|19|17|І це стало відоме юдеям та гелленам, усім, що в Ефесі замешкують, і острах напав на всіх їх, і славилося Ім'я Господа Ісуса.
ACTS|19|18|І багато-хто з тих, що ввірували, приходили, визнаваючи та відкриваючи вчинки свої.
ACTS|19|19|І багато-хто з тих, що займалися чарами, позносили книги свої та й перед усіма попалили. І злічили ціну їх, і вийшло на срібло п'ятдесят тисяч драхм.
ACTS|19|20|Так могуче росло та зміцнялося Божеє Слово!
ACTS|19|21|А як сповнилось це, Павло в Дусі задумав перейти Македонію та Ахаю, та й удатись у Єрусалим, говорячи: Як побуду я там, то треба мені й Рим побачити.
ACTS|19|22|Тож він послав у Македонію двох із тих, що служили йому, Тимофія й Ераста, а сам позостався якийсь час ув Азії.
ACTS|19|23|І розрух чималий був стався там часу того за Господню дорогу.
ACTS|19|24|Бо один золотар, Дмитро на ім'я, що робив срібляні Артемідині храмки, та ремісникам заробіток чималий давав,
ACTS|19|25|згромадив він їх і ще інших подібних робітників, та й промовив: Ви знаєте, мужі, що з цього ремесла заробіток ми маємо.
ACTS|19|26|І ви бачите й чуєте, що не тільки в Ефесі, але мало не в усій Азії цей Павло збаламутив і відвернув багатенно народу, говорячи, ніби то не боги, що руками пороблені.
ACTS|19|27|І не тільки оце нам загрожує, що прийде зайняття в упадок, а й храм богині великої Артеміди в ніщо зарахується, і буде зруйнована й велич тієї, що шанує її ціла Азія та цілий світ.
ACTS|19|28|Почувши ж оце, вони переповнились гнівом, та й стали кричати, говорячи: Артеміда ефеська велика!
ACTS|19|29|І місто наповнилось заколотом. І кинулися однодушно до видовища, схопивши Павлових супутників Гая та Аристарха, македонян.
ACTS|19|30|Як Павло ж хотів у народ увійти, то учні його не пустили.
ACTS|19|31|Також дехто з азійських начальників, що були йому приятелі, послали до нього й просили, щоб він не вдававсь на видовище.
ACTS|19|32|І кожен що інше кричав, бо збори бурхливі були, і багатенно з них навіть не знали, чого ради зібралися.
ACTS|19|33|А з народу взяли Олександра, бо юдеї його висували. І Олександер дав знака рукою, і хотів виправдатися перед народом.
ACTS|19|34|А коли розпізнали, що юдеянин він, то злилися всі в один голос, і годин зо дві гукали: Артеміда ефеська велика!
ACTS|19|35|А як писар міський заспокоїв народ, то промовив: Мужі ефеські, яка ж то людина не знає, що місто Ефес то храмовий доглядач Артеміди великої й її образу, упалого з неба?
ACTS|19|36|Коли ж цьому перечити не можна, то потрібно вам бути спокійними, і не робити необачно нічого.
ACTS|19|37|А ви ж привели цих людей, що ані святокрадці, ані вашої богині не зневажили.
ACTS|19|38|Отож, як Дмитро та його ремісники мають справу на кого, то суди є на ринку й проконсули, один одного хай позивають.
ACTS|19|39|А коли чогось іншого допоминаєтеся, то те вирішиться на законнім зібранні.
ACTS|19|40|Бо ось є небезпека, що нас за сьогоднішній розрух оскаржити можуть, і немає жадної причини, якою могли б виправдати це зборище.
ACTS|19|41|(19-40) І, промовивши це, розпустив він громаду.
ACTS|20|1|А як заколот стих, то Павло скликав учнів, і, потішивши та попрощавшись із ними, вибрався йти в Македонію.
ACTS|20|2|Перейшовши ж ті сторони та підбадьоривши їх довгим словом, прибув до Геллади,
ACTS|20|3|і прожив там три місяці. А як він захотів був відплинути в Сирію, то змову на нього вчинили юдеї, тому він узяв думку вертатись через Македонію.
ACTS|20|4|Разом із ним пішов Сопатер Піррів із Верії, Аристарх та Секунд із Солуня, і Гай дерв'янин, і Тимофій, а з азійців Тихик та Трохим.
ACTS|20|5|Вони відбули наперед, і нас дожидали в Троаді.
ACTS|20|6|А ми відпливли із Филипів по святах Опрісноків, і прибули днів за п'ять у Троаду до них, де сім день прожили.
ACTS|20|7|А дня першого в тижні, як учні зібралися на ламання хліба, Павло мав промову до них, бо вранці збирався відбути, і затягнув своє слово до півночі.
ACTS|20|8|А в горниці, де зібралися ми, було багато світел.
ACTS|20|9|Юнак же один, Євтих на ім'я, сидів на вікні. Його обгорнув міцний сон, бо задовго Павло промовляв, і він сонний хитнувся, і додолу упав із третього поверху, і підняли його мертвого...
ACTS|20|10|Зійшов же Павло та до нього припав, і, обнявши його, проказав: Заспокойтесь, бо душа його в ньому!
ACTS|20|11|А вернувшись, він хліб переломив і спожив, і бесіду довго точив, аж до досвітку, потім відбув.
ACTS|20|12|А хлопця живим привели, і зраділи немало.
ACTS|20|13|А ми наперед пішли до корабля, та в Асс попливли, щоб звідти забрати Павла, бо він так ізвелів, сам бажаючи пішки піти.
ACTS|20|14|А коли він із нами зійшовся в Ассі, ми взяли його та прибули в Мітілену.
ACTS|20|15|І, відплинувши звідти, ми назавтра пристали навпроти Хіосу, а другого дня припливли до Самосу, наступного ж ми прибули до Мілету.
ACTS|20|16|Бо Павло захотів поминути Ефес, щоб йому не баритися в Азії, бо він квапився, коли буде можливе, бути в Єрусалимі на день П'ятдесятниці.
ACTS|20|17|А з Мілету послав до Ефесу, і прикликав пресвітерів Церкви.
ACTS|20|18|І, як до нього вони прибули, він промовив до них: Ви знаєте, як із першого дня, відколи прибув в Азію, я з вами ввесь час перебував,
ACTS|20|19|і служив Господеві з усією покорою, і з рясними слізьми та напастями, що спіткали мене від юдейської змови,
ACTS|20|20|як нічого корисного я не минув, щоб його вам звістити й навчити вас прилюдно і в домах.
ACTS|20|21|І я свідчив юдеям та гелленам, щоб вони перед Богом покаялись, та ввірували в Господа нашого Ісуса Христа.
ACTS|20|22|І ось тепер, побуджений Духом, подаюсь я в Єрусалим, не відаючи, що там трапитись має мені,
ACTS|20|23|тільки Дух Святий в кожному місті засвідчує, кажучи, що кайдани та муки чекають мене...
ACTS|20|24|Але я ні про що не турбуюсь, і свого життя не вважаю для себе цінним, аби но скінчити дорогу свою та служіння, яке я одержав від Господа Ісуса, щоб засвідчити Євангелію благодаті Божої.
ACTS|20|25|І ось я знаю тепер, що обличчя мого більш не будете бачити всі ви, між якими ходив я, проповідуючи Царство Боже...
ACTS|20|26|Тому дня сьогоднішнього вам свідкую, що я чистий від крови всіх,
ACTS|20|27|бо я не вхилявсь об'являти вам усю волю Божу!
ACTS|20|28|Пильнуйте себе та всієї отари, в якій Святий Дух вас поставив єпископами, щоб пасти Церкву Божу, яку власною кров'ю набув Він.
ACTS|20|29|Бо я знаю, що як я відійду, то ввійдуть між вас вовки люті, що отари щадити не будуть...
ACTS|20|30|Із вас самих навіть мужі постануть, що будуть казати перекручене, аби тільки учнів тягнути за собою...
ACTS|20|31|Тому то пильнуйте, пам'ятаючи, що я кожного з вас день і ніч безперестань навчав зо слізьми ось три роки.
ACTS|20|32|А тепер доручаю вас Богові та слову благодаті Його, Який має силу будувати та дати спадщину, серед усіх освячених.
ACTS|20|33|Ні срібла, ані золота, ні одежі чиєїсь я не побажав...
ACTS|20|34|Самі знаєте, що ці руки мої послужили потребам моїм та отих, хто був зо мною.
ACTS|20|35|Я вам усе показав, що, працюючи так, треба поміч давати слабим, та пам'ятати слова Господа Ісуса, бо Він Сам проказав: Блаженніше давати, ніж брати!
ACTS|20|36|Проказавши ж оце, він навколішки впав, та й із ними всіма помолився.
ACTS|20|37|І знявсь між усіма плач великий, і вони припадали на Павлову шию, і його цілували...
ACTS|20|38|А найтяжче вони сумували з-за слова, яке він прорік, що не бачитимуть більш обличчя його. І вони провели його до корабля.
ACTS|21|1|А як ми розлучилися з ними й відплинули, то дорогою простою в Кос прибули, а другого дня до Родосу, а звідти в Патару.
ACTS|21|2|І знайшли корабля, що плив у Фінікію, увійшли та й поплинули.
ACTS|21|3|А коли показався нам Кіпр, ми лишили ліворуч його та й поплинули в Сирію. І пристали ми в Тирі, бо там корабель вантажа мав скласти.
ACTS|21|4|І, учнів знайшовши, перебули тут сім день. Вони через Духа казали Павлові, щоб до Єрусалиму не йшов.
ACTS|21|5|І, як дні побуту скінчилися, то ми вийшли й пішли, а всі нас проводили з дружинами й дітьми аж за місто. І, ставши навколішки, помолились на березі.
ACTS|21|6|І, попрощавшись один із одним, ми ввійшли в корабель, а вони повернулись додому.
ACTS|21|7|А ми, закінчивши від Тиру плавбу, пристали до Птолемаїди, і, братів привітавши, один день перебули в них.
ACTS|21|8|А назавтра в дорогу ми вибрались, і прийшли в Кесарію. І ввійшли до господи благовісника Пилипа, одного з семи, і позосталися в нього.
ACTS|21|9|Він мав чотири панні дочки, що пророкували.
ACTS|21|10|І коли ми багато днів у них зоставались, то прибув із Юдеї якийсь пророк, Агав на ім'я.
ACTS|21|11|І прийшов він до нас, і взяв пояса Павлового, та й зв'язав свої руки та ноги й сказав: Дух Святий так звіщає: Отак зв'яжуть в Єрусалимі юдеї того мужа, що цей пояс його, і видадуть в руки поган...
ACTS|21|12|Як почули ж оце, то благали ми та тамтешні Павла, щоб до Єрусалиму не йшов.
ACTS|21|13|А Павло відповів: Що робите ви, плачучи та серце мені розриваючи? Бо за Ім'я Господа Ісуса я готовий не тільки зв'язаним бути, а й померти в Єрусалимі!
ACTS|21|14|І не могли ми його вмовити, і замовкли, сказавши: Нехай діється Божая воля!
ACTS|21|15|А після оцих днів приготувались ми, та до Єрусалиму вирушили.
ACTS|21|16|А з нами пішли й деякі учні із Кесарії, ведучи якогось кіпрянина Мнасона, давнього учня, що ми в нього спинитися мали.
ACTS|21|17|А коли ми прийшли в Єрусалим, то брати прийняли нас гостинно.
ACTS|21|18|А другого дня Павло з нами подався до Якова. І всі старші посходились.
ACTS|21|19|Поздоровивши ж їх, розповів він докладно, що Бог через служіння його вчинив між поганами.
ACTS|21|20|Як вони ж це почули, то славили Бога, а до нього промовили: Бачиш, брате, скільки тисяч серед юдеїв увірувало, і всі вони ревні оборонці Закону!
ACTS|21|21|Вони ж чули про тебе, ніби ти всіх юдеїв, що живуть між поганами, навчаєш відступлення від Мойсея, говорячи, щоб дітей не обрізували й не тримались звичаїв.
ACTS|21|22|Що ж почати? Люд збереться напевно, бо почують, що прибув ти.
ACTS|21|23|Отже, зроби це, що порадимо тобі. Ми маємо чотирьох мужів, що обітницю склали на себе.
ACTS|21|24|Візьми їх, та й із ними очисться, і видатки за них заплати, щоб постригли їм голови. І пізнають усі, що неправда про тебе їм сказане, та й що сам ти Закона пильнуєш.
ACTS|21|25|А про тих із поган, що ввірували, ми писали, розсудивши, щоб вони береглися від ідольських жертов та крови й задушенини, та від блуду.
ACTS|21|26|Тоді взяв Павло мужів отих, і назавтра очистився з ними, і ввійшов у храм, і звістив про виконання днів очищення, так, аж за кожного з них була жертва принесена.
ACTS|21|27|А коли ті сім день закінчитися мали, то азійські юдеї, як побачили в храмі його, підбурили ввесь народ, та руки на нього наклали,
ACTS|21|28|кричачи: Ізраїльські мужі, рятуйте! Це людина ота, що проти народу й Закону та місця цього всіх усюди навчає!... А до того у храм упровадив і гелленів, і занечистив це місце святе!
ACTS|21|29|Бо перед тим вони бачили в місті з ним разом Трохима ефесянина, і гадали про нього, що Павло то його ввів у храм.
ACTS|21|30|І порушилося ціле місто, і повстало збіговисько люду. І, схопивши Павла, потягли його поза храм, а двері негайно зачинено...
ACTS|21|31|Як хотіли ж забити його, то вістка досталась до полкового тисяцього, що ввесь Єрусалим збунтувався!
ACTS|21|32|І він зараз узяв вояків та сотників, і подався до них. А вони, як угледіли тисяцького й вояків, то бити Павла перестали.
ACTS|21|33|Приступив тоді тисяцький, та й ухопив його, і двома ланцюгами зв'язати звелів, і допитувати став: хто такий він і що він зробив?
ACTS|21|34|Але кожен що інше викрикував у натовпі. І, не мігши довідатись певного через заколот, він звелів відпровадити його до фортеці.
ACTS|21|35|А коли він до сходів прийшов, то трапилося, що мусіли нести його вояки із-за натовпу людського,
ACTS|21|36|бо безліч народу йшла слідкома та кричала: Геть із ним!
ACTS|21|37|А коли Павло входив до фортеці, то тисяцького поспитався: Чи можна мені щось сказати тобі? А той відказав: То ти вмієш по-грецькому?
ACTS|21|38|Чи не той ти єгиптянин, що перед цими днями призвів був до бунту, і випровадив до пустині чотири тисячі потаємних убійників?
ACTS|21|39|А Павло відказав: Я юдеянин із Тарсу, громадянин відомого міста в Кілікії. Благаю тебе, дозволь мені до народу промовити!
ACTS|21|40|А коли той дозволив, то Павло став на сходах, і дав знака рукою народові. А як тиша велика настала, промовив єврейською мовою, кажучи:
ACTS|22|1|Мужі-браття й батьки! Послухайте ось тепер виправдання мого перед вами!
ACTS|22|2|Як зачули ж вони, що до них він говорить єврейською мовою, то тиша ще більша настала. А він промовляв:
ACTS|22|3|Я юдеянин, що родився в кілікійському Тарсі, а вихований у цім місті, у ніг Гамаліїла докладно навчений Закону отців; горливець я Божий, як і всі ви сьогодні.
ACTS|22|4|Переслідував я аж до смерти цю путь, і в'язав, і до в'язниці вкидав чоловіків і жінок,
ACTS|22|5|як засвідчить про мене первосвященик та вся старшина. Я від них був узяв навіть листи на братів, і пішов до Дамаску, щоб тамтешніх зв'язати й привести до Єрусалиму на кару.
ACTS|22|6|І сталося, як у дорозі я був, і наближавсь до Дамаску опівдня, то ось мене нагло осяяло світло велике з неба!
ACTS|22|7|І я повалився на землю, і голос почув, що мені говорив: Савле, Савле, чому ти Мене переслідуєш?
ACTS|22|8|А я запитав: Хто Ти, Господи? А Він мені відказав: Я Ісус Назарянин, що Його переслідуєш ти...
ACTS|22|9|А ті, що зо мною були, правда, бачили світло, але не почули вони того голосу, що мені говорив.
ACTS|22|10|А я запитав: Що я, Господи, маю робити? Господь же до мене промовив: Уставай та й іди до Дамаску, а там тобі скажуть про все, що тобі призначено робити.
ACTS|22|11|А від ясности світла того невидющим я став... І присутні зо мною за руку мене повели, і до Дамаску прибув я.
ACTS|22|12|А один муж Ананій, у Законі побожний, що добре свідоцтво про нього дають усі юдеї в Дамаску,
ACTS|22|13|до мене прибув, і, ставши, промовив мені: Савле брате, стань видющий! І я хвилі тієї побачив його...
ACTS|22|14|І озвавсь він до мене: Бог отців наших вибрав тебе, щоб ти волю Його зрозумів, і щоб бачив ти Праведника, і почув голос із уст Його.
ACTS|22|15|Бо будеш ти свідком Йому перед усіма людьми про оте, що ти бачив та чув!
ACTS|22|16|А тепер чого гаєшся? Уставай й охристися, і обмий гріхи свої, прикликавши Ймення Його!
ACTS|22|17|І сталось, як вернувся я в Єрусалим, і молився у храмі, то в захоплення впав я,
ACTS|22|18|і побачив Його, що до мене сказав: Поспіши, і піди хутчій з Єрусалиму, бо не приймуть свідоцтва твого про Мене...
ACTS|22|19|А я відказав: Самі вони, Господи, знають, що я до в'язниць садовив та бив по синагогах отих, хто вірував у Тебе.
ACTS|22|20|А коли лилась кров Твого свідка Степана, то сам я стояв та вбивство його похваляв, і одежу вбивців його сторожив...
ACTS|22|21|Але Він до мене промовив: Іди, бо пошлю Я далеко тебе, до поган!
ACTS|22|22|І аж до слова цього його слухали. Аж ось піднесли вони голос свій, гукаючи: Геть такого з землі, бо жити йому не годиться!...
ACTS|22|23|І як вони верещали, і одежу шпурляли, і кидали порох у повітря,
ACTS|22|24|то звелів тисяцький у фортецю його відвести, і звелів бичуванням його допитати, щоб довідатися, з якої причини на нього вони так кричали.
ACTS|22|25|І як його розтягли для ремінних бичів, то Павло сказав сотникові, що стояв: Хіба бичувати дозволено вам громадянина римського та ще й незасудженого?
ACTS|22|26|Якже сотник це почув, то подався до тисяцького, і завідомив, говорячи: Що хочеш робити? Бож римлянин цей чоловік!
ACTS|22|27|Підійшов тоді тисяцький, та й поспитався його: Скажи мені, чи ти римлянин? А він: Так! відказав.
ACTS|22|28|Відповів на те тисяцький: За великі гроші громадянство оце я набув... А Павло відказав: А я в нім і родився!
ACTS|22|29|І відступили негайно від нього оті, що хотіли допитувати його. І злякався тисяцький, довідавшись, що той римлянин, і що він ізв'язав був його.
ACTS|22|30|А другого дня, бажавши довідатись правди, у чому юдеї його оскаржають, він звільнив його та звелів, щоб зібралися первосвященики та ввесь синедріон. І він вивів Павла, і поставив його перед ними.
ACTS|23|1|І вп'явся очима Павло на той синедріон і промовив: Мужі-браття, я аж по сьогоднішній день жив для Бога всім добрим сумлінням!
ACTS|23|2|Але первосвященик Ананій звелів тим, що стояли при ньому, щоб били його по устах.
ACTS|23|3|Тоді промовив до нього Павло: Тебе битиме Бог, ти стіно побілена... Ти ж сидиш, щоб судити мене за Законом, наказуєш бити мене проти Закону?
ACTS|23|4|А присутні сказали: То ти Божому первосвященикові лихословиш?
ACTS|23|5|І промовив Павло: Не знав я, брати, що то первосвященик. Бо написано: На начальника люду твого не лихослов.
ACTS|23|6|І Павло, спостерігши, що частина одна саддукеї, а друга фарисеї, покликнув у синедріоні: Мужі-браття, я фарисей, і син фарисея. За надію на воскресення мертвих мене судять!
ACTS|23|7|Якже він це промовив, колотнеча постала поміж саддукеями та фарисеями, і розділилась юрба.
ACTS|23|8|Саддукеї бо твердять, що немає воскресення, ані Ангола, ані духа, фарисеї ж оце визнають.
ACTS|23|9|І галас великий зчинився. А деякі книжники, із фарисейської групи, уставши, почали сперечатися, кажучи: У чоловікові цьому ми жадного лиха не знаходимо! А коли промовляв Дух до нього, чи Ангол, не противмося Богові.
ACTS|23|10|А коли колотнеча велика зчинилась, то тисяцький, боячись, щоб Павла не роздерли, звелів воякам увійти та забрати його з-поміж них, і відвести в фортецю.
ACTS|23|11|А наступної ночі став Господь перед ним і промовив: Будь бадьорий! Бо як в Єрусалимі про Мене ти свідчив, так треба тобі свідкувати й у Римі!
ACTS|23|12|А коли настав день, то дехто з юдеїв зібрались, та клятву склали, говорячи, що ні їсти, ні пити не будуть, аж доки Павла не заб'ють!
ACTS|23|13|А тих, що закляття таке поклали, було більш сорока.
ACTS|23|14|І вони приступили до первосвящеників та старших і сказали: Ми клятву склали нічого не їсти, аж поки заб'ємо Павла!
ACTS|23|15|Отож разом із синедріоном передайте тисяцькому, щоб до вас він привів його, ніби хочете ви докладніш розізнати про нього. А ми, перше ніж він наблизиться, готові забити його...
ACTS|23|16|Як зачув же сестрінець Павлів про цю змову, то прибув, і ввійшов у фортецю, і Павла завідомив.
ACTS|23|17|Павло ж зараз покликав одного з сотників, та й сказав: Цього юнака запровадь до тисяцького, бо він має йому щось сказати.
ACTS|23|18|Той же взяв його, та й запровадив до тисяцького та сказав: Павло в'язень покликав мене, і просив запровадити до тебе цього юнака, що має тобі щось сказати.
ACTS|23|19|І взяв тисяцький того за руку, і набік відвів і спитав: Що ти маєш звістити мені?
ACTS|23|20|А той розповів: Змову склали юдеї, просити тебе, щоб ти взавтра до синедріону Павла припровадив, ніби хочуть вони докладніш розпізнати про нього.
ACTS|23|21|Отож, не послухайся їх, бо чигає на нього їх більш сорока чоловіка, що клятву склали ні їсти, ні пити, аж доки його не заб'ють... І тепер он готові вони, і чекають твого приречення.
ACTS|23|22|Тоді тисяцький відпустив юнака, наказавши йому не розповідати ані одному, що мені ти це виявив.
ACTS|23|23|І він закликав котрихсь двох із сотників, і наказа: Пришикуйте на третю годину вночі дві сотні вояків, щоб іти до Кесарії, і кіннотчиків сімдесят, та дві сотні стрільців.
ACTS|23|24|Приготуйте також в'ючаків і Павла посадіть, і здоровим його проведіть до намісника Фелікса.
ACTS|23|25|І листа написав він такого ось змісту:
ACTS|23|26|Клавдій Лісій намісникові вседостойному Феліксові поздоровлення!
ACTS|23|27|Цього мужа, що його юдеї схопили були та хотіли забити, урятувава я, із вояками прийшовши, довідавшися, що він римлянин.
ACTS|23|28|І хотів я довідатися про причину, що за неї його оскаржали, та й привів був його до їхнього синедріону.
ACTS|23|29|Я знайшов, що його винуватять у спірних речах їхнього Закону, і що провини не має він жадної, вартої смерти або ланцюгів.
ACTS|23|30|Як донесли ж мені про ту змову, що юдеї вчинили на мужа цього, я зараз до тебе його відіслав, наказавши також позивальникам, щоб перед тобою сказали, що мають на нього. Будь здоровий!
ACTS|23|31|Отож вояки, як наказано їм, забрали Павла, і вночі попровадили в Антипатриду.
ACTS|23|32|А другого дня, полишивши кіннотчиків, щоб ішли з ним, у фортецю вони повернулись.
ACTS|23|33|А ті прибули в Кесарію, і, листа передавши намісникові, поставили також Павла перед ним.
ACTS|23|34|Намісник листа прочитав і спитав, із якого він краю. А довідавшись, що з Кілікії, промовив:
ACTS|23|35|Я тебе переслухаю, як прийдуть і твої позивальники. І звелів стерегти його в Іродовому преторії.
ACTS|24|1|А по п'яти днях прибув первосвященик Ананій з якимись старшими, та з промовцем якимсь Тертилом, що перед намісником скаржилися на Павла.
ACTS|24|2|Коли ж він був покликаний, то Тертил оскаржати зачав, промовляючи: Через тебе великий мир маємо ми, і для народу цього добрі речі впроваджено через дбайливість твою,
ACTS|24|3|це ми завжди і скрізь визнаємо з подякою щирою, вседостойний наш Феліксе!
ACTS|24|4|Та щоб довго тебе не турбувати, то благаю тебе, щоб ти коротко вислухав нас зо своєї ласкавости.
ACTS|24|5|Ми переконались, що цей чоловік то зараза, і що він колотнечу викликує між усіма юдеями в цілому світі, і що він провідник Назорейської єресі.
ACTS|24|6|Він відважився навіть збезчестити храм, і його ми схопили були, і судити хотіли за нашим Законом.
ACTS|24|7|Але тисяцький Лісій прибув, і з великим насильством видер його з наших рук,
ACTS|24|8|а його винувальникам звелів йти до тебе. Ти сам зможеш від нього, розпитавши, дізнатись про все, у чому його ми винуємо.
ACTS|24|9|Юдеї також прилучились до того, говорячи, що то так.
ACTS|24|10|І як намісник дав знака йому говорити, то Павло відповів: Я знаю, що від літ багатьох ти суддя для народу цього, тому буду сміліш боронитись.
ACTS|24|11|Ти можеш довідатися, що нема більш дванадцяти день, як прийшов я до Єрусалиму вклонитися.
ACTS|24|12|І вони ані в храмі, ані в синагогах, ні в місті мене не здибали, щоб я з ким сперечався, або колотнечу в народі здіймав.
ACTS|24|13|І не можуть вони довести тобі того, у чому тепер оскаржають мене.
ACTS|24|14|Але признаюсь тобі, що в дорозі оцій, яку звуть вони єрессю, я Богові отців служу так, що вірую всьому, що в Законі й у Пророків написане.
ACTS|24|15|І маю надію я в Бозі, чого й самі вони сподіваються, що настане воскресення праведних і неправедних.
ACTS|24|16|І я пильно дбаю про те, щоб завсіди мати сумління невинне, щодо Бога й людей.
ACTS|24|17|А по довгих роках я прибув, щоб подати моєму народові милостиню та приноси.
ACTS|24|18|Ось при цьому знайшли мене дехто з юдеїв азійських очищеного в храмі, а не з натовпом чи з колотнечею.
ACTS|24|19|Їм належало б ось перед тебе прибути й казати, коли мають вони що на мене.
ACTS|24|20|Або самі ці нехай скажуть, чи якусь неправду знайшли на мені, як я в синедріоні стояв,
ACTS|24|21|крім отого єдиного виразу, що я його крикнув, стоячи серед них: За воскресення мертвих приймаю від вас суд сьогодні!
ACTS|24|22|Але Фелікс, дуже добре дорогу цю знавши, відрочив їм справу, говорячи: Розсуджу вашу справу, коли тисяцький Лісій прибуде.
ACTS|24|23|І він сотникові наказав сторожити Павла, але мати полегшу, і не боронити нікому з близьких його, щоб служили йому.
ACTS|24|24|А по декількох днях прийшов Фелікс із дружиною своєю Друзіллою, що була юдеянка, і покликав Павла, та слухав від нього про віру в Ісуса Христа.
ACTS|24|25|І як розповідав він про праведність, і про здержливість, та про майбутній суд, то Фелікса страх обгорнув, і він відповів: Тепер іди собі, відповідного ж часу покличу тебе!
ACTS|24|26|Разом із тим і сподівався він, що дасть Павло грошей йому, тому й часто його прикликав і розмову з ним вів.
ACTS|24|27|Як минуло ж два роки, то Фелікс одержав наступника, Порція Феста. А Фелікс бажав догодити юдеям, і в в'язниці Павла залишив.
ACTS|25|1|А коли прибув Фест до свого намісництва, то він по трьох днях відійшов із Кесарії до Єрусалиму.
ACTS|25|2|І поскаржилися йому на Павла первосвященики та головніші з юдеїв, і благали його,
ACTS|25|3|і ніби милости просили для нього, щоб до Єрусалиму його припровадив, вони змову вчинили, щоб смерть заподіяти йому по дорозі.
ACTS|25|4|А Фест відповів, що Павла стережуть у Кесарії, і він сам незабаром туди подається.
ACTS|25|5|Отже, сказав він, хто спроможен із вас, нехай ті вирушають разом зо мною, і коли є неправда яка в чоловікові цьому, нехай оскаржають його.
ACTS|25|6|І, пробувши в них днів не більше як вісім чи десять, він повернувся до Кесарії. А другого дня він засів на суддевім сидінні, і звелів, щоб привести Павла.
ACTS|25|7|Як його ж привели, то стали навколо юдеї, що поприходили з Єрусалиму, і Павлу закидали багато тяжких винувачень, що їх не могли довести,
ACTS|25|8|бо Павло боронився: Я не провинився ні в чім ані проти Закону юдейського, ані проти храму, ані супроти кесаря.
ACTS|25|9|Тоді Фест, що бажав догодити юдеям, промовив Павлові на відповідь: Чи ти хочеш до Єрусалиму піти, і там суд прийняти від мене про це?
ACTS|25|10|Та Павло відказав: Я стою перед судом кесаревим, де належить мені суд прийняти. Юдеїв нічим я не скривдив, як і ти дуже добре те знаєш.
ACTS|25|11|Бо коли допустився я кривди, або гідне смерти вчинив що, то не відмовляюся вмерти. Як нема ж нічого того, у чім вони винуватять мене, то не може ніхто мене видати їм. Відкликаюсь до кесаря!
ACTS|25|12|Тоді Фест, побалакавши з радою, відповідь дав: Ти відкликавсь до кесаря, до кесаря підеш!
ACTS|25|13|Як минуло ж днів кілька, цар Агріппа й Верніка приїхали до Кесарії, щоб Феста вітати.
ACTS|25|14|А що там багато днів вони пробули, то Фест виклав справу Павлову цареві й промовив: Є один чоловік від Фелікса лишений в'язень,
ACTS|25|15|на якого, як в Єрусалимі я був, первосвященики й старші юдейські принесли скаргу, домагаючись його осуду.
ACTS|25|16|Я їм відповів, що римляни не мають звичаю людину якусь видавати на згубу, поки пізваний перед собою не матиме обвинувачів, і не буде йому дано можности для оборони від закидів.
ACTS|25|17|І як зійшлись вони тут, то я, зволікання не роблячи жадного, сів наступного дня на сидіння суддеве, і звелів привести цього мужа.
ACTS|25|18|І винувальники стали круг нього, проте не вказали вини ані жадної з тих, яких я сподівався.
ACTS|25|19|Та мали вони проти нього якісь суперечки про власне своє марновірство, і про якогось Ісуса померлого, про Якого Павло твердив, що живий Він.
ACTS|25|20|І я був непевний у цьому змаганні й спитав, чи не хоче піти він до Єрусалиму, і там суд прийняти про це?
ACTS|25|21|Через те ж, що Павло заявив, щоб залишений був він на кесарів розсуд, я звелів сторожити його, аж поки його не відправлю до кесаря.
ACTS|25|22|А Агріппа промовив до Феста: Хотів би і я цього мужа послухати! Узавтра сказав той почуєш його.
ACTS|25|23|А назавтра Агріппа й Верніка прийшли з превеликою пишнотою, і на залю судову ввійшли разом з тисяцькими та значнішими мужами міста. І як Фест наказав, то Павло був приведений.
ACTS|25|24|І сказав до них Фест: О царю Агріппо, та з нами присутні всі мужі! Ви бачите того, що за нього ввесь люд юдейський мені докучав в Єрусалимі та тут, кричачи, що йому не повинно більш жити.
ACTS|25|25|Я ж дізнавсь, що нічого, вартого смерти, він не вчинив; а що сам він відкликавсь до Августа, розсудив я послати його.
ACTS|25|26|Нічого не маю я певного, що міг би про нього писати до пана. Тому я припровадив його перед вас, а найбільш перед тебе, царю Агріппо, щоб після переслухання мав що писати.
ACTS|25|27|Бо здається мені нерозважливим ув'язненого посилати, і не означити обвинувачень на нього.
ACTS|26|1|А Агріппа сказав до Павла: Дозволяємо тобі говорити про себе самого. Павло тоді простягнув руку, і промовив у своїй обороні:
ACTS|26|2|О царю Агріппо! Уважаю себе за щасливого, що сьогодні я перед тобою боронитися маю з усього, у чім мене винуватять юдеї,
ACTS|26|3|особливо ж тому, що ти знаєш усі юдейські звичаї та суперечки. Тому я прошу мене вислухати терпляче.
ACTS|26|4|А життя моє змалку, що спочатку точилося в Єрусалимі серед народу мого, знають усі юдеї,
ACTS|26|5|які відають здавна мене, аби тільки схотіли засвідчити, що я жив фарисеєм за найдокладнішою сектою нашої віри.
ACTS|26|6|І тепер я стою отут суджений за надію обітниці, що Бог дав її нашим отцям,
ACTS|26|7|а її виконання чекають побачити наші дванадцять племен, служачи Богові безперестанно вдень та вночі. За цю надію, о царю, мене винуватять юдеї!
ACTS|26|8|Чому ви вважаєте за неймовірне, що Бог воскрешає померлих?
ACTS|26|9|Правда, думав був я, що мені належить чинити багато ворожого проти Ймення Ісуса Назарянина,
ACTS|26|10|що я в Єрусалимі й робив, і багато кого зо святих до в'язниць я замкнув, як отримав був владу від первосвящеників; а як їх убивали, я голос давав проти них.
ACTS|26|11|І часто по всіх синагогах караючи їх, до богозневаги примушував я, а лютуючи вельми на них, переслідував їх навіть по закордонних містах.
ACTS|26|12|Коли в цих справах я йшов до Дамаску зо владою та припорученням первосвящеників,
ACTS|26|13|то опівдні, о царю, на дорозі побачив я світло із неба, ясніше від світлости сонця, що осяяло мене та тих, хто разом зо мною йшов!...
ACTS|26|14|І як ми всі повалились на землю, я голос почув, що мені говорив єврейською мовою: Савле, Савле, чому ти Мене переслідуєш? Трудно тобі бити ногою колючку!
ACTS|26|15|А я запитав: Хто Ти, Господи? А Він відказав: Я Ісус, що Його переслідуєш ти.
ACTS|26|16|Але підведися, і стань на ноги свої. Бо на те Я з'явився тобі, щоб тебе вчинити слугою та свідком того, що ти бачив та що Я відкрию тобі.
ACTS|26|17|Визволяю тебе від твого народу та від поган, до яких Я тебе посилаю,
ACTS|26|18|відкрити їм очі, щоб вони навернулись від темряви в світло та від сатаниної влади до Бога, щоб вірою в Мене отримати їм дарування гріхів і долю з освяченими.
ACTS|26|19|Через це я, о царю Агріппо, не був супротивний видінню небесному,
ACTS|26|20|але мешканцям перше Дамаску, потім Єрусалиму й усякого краю юдейського та поганам я проповідував, щоб покаялися й навернулись до Бога, і чинили діла, гідні покаяння.
ACTS|26|21|Через це юдеї в святині схопили мене та й хотіли роздерти.
ACTS|26|22|Але, поміч від Бога одержавши, я стою аж до дня сьогоднішнього та свідкую малому й великому, нічого не розповідаючи, окрім того, що сказали Пророки й Мойсей, що статися має,
ACTS|26|23|що має Христос постраждати, що Він, як перший воскреснувши з мертвих, проповідувати буде світло народові й поганам!
ACTS|26|24|Коли ж він боронився отак, то Фест проказав гучним голосом: Дурієш ти, Павле! Велика наука доводить тебе до нерозуму!
ACTS|26|25|А Павло: Не дурію сказав, о Фесте достойний, але провіщаю слова правди та щирого розуму.
ACTS|26|26|Цар бо знає про це, до нього з відвагою я й промовляю. Бо не гадаю я, щоб із цього щобудь сховалось від нього, бо не в закутку діялось це.
ACTS|26|27|Чи віруєш, царю Агріппо, Пророкам? Я знаю, що віруєш.
ACTS|26|28|Агріппа ж Павлові: Ти малощо не намовляєш мене, щоб я став християнином...
ACTS|26|29|А Павло: Благав би я Бога, щоб чи мало, чи багато, не тільки но ти, але й усі, хто чує сьогодні мене, зробились такими, як і я, крім оцих ланцюгів...
ACTS|26|30|І встав цар та намісник, і Верніка та ті, хто з ними сидів.
ACTS|26|31|І набік вони відійшли, і розмовляли один до одного й казали: Нічого, вартого смерти або ланцюгів, чоловік цей не робить!
ACTS|26|32|Агріппа ж до Феста сказав: Міг би бути відпущений цей чоловік, якби не відкликавсь був до кесаря.
ACTS|27|1|А коли постановлено, щоб відплинули ми до Італії, то віддано Павла та ще деяких інших ув'язнених сотникові, Юлієві на ім'я, з полку Августа.
ACTS|27|2|І посідали ми на корабля адрамітського, що пливсти мав біля місць азійських, та й відчалили. Із нами був Арістарх македонець із Солуня.
ACTS|27|3|А другого дня ми пристали в Сидоні. До Павла ж Юлій ставивсь по-людському, і дозволив до друзів піти, та їхньої опіки зазнати.
ACTS|27|4|А вирушивши звідти, припливли ми до Кіпру, бо вітри супротивні були.
ACTS|27|5|Коли ж переплинули море, що біля Кілікії й Памфілії, то ми прибули до Лікійської Міри.
ACTS|27|6|І там сотник знайшов корабля олександрійського, що плинув в Італію, і всадив нас на нього.
ACTS|27|7|І днів багато помалу пливли ми, і насилу насупроти Кніду приплинули, а що вітер нас не допускав, попливли ми додолу на Кріт при Салмоні.
ACTS|27|8|І коли ми насилу минули його, то припливли до одного місця, що зветься Доброю Пристанню, недалеко якого знаходиться місто Ласея.
ACTS|27|9|А як часу минуло багато, і була вже плавба небезпечна, бо минув уже й піст, то зачав Павло радити,
ACTS|27|10|говорячи їм: О мужі! Я бачу, що буде плавба з перешкодами та з великим ущербком не лиш для вантажу й корабля, але й для наших душ.
ACTS|27|11|Та сотник довіряв більше стерничому та власникові корабля, ніж тому, що Павло говорив.
ACTS|27|12|А що пристань була на зимівлю невигідна, то більшість давала пораду відплинути звідти, щоб, як можна, дістатись до Фініка, і перезимувати в пристані крітській, неприступній західнім вітрам із півдня та з півночі.
ACTS|27|13|А як вітер південний повіяв, то подумали, що бажання вони досягли, тому витягли кітви й попливли покрай Кріту.
ACTS|27|14|Але незабаром ударив на них рвачкий вітер, що зветься евроклідон.
ACTS|27|15|А коли корабель був підхоплений, і не міг противитись вітрові, то йому віддались ми й понеслися.
ACTS|27|16|І наїхали ми на один острівець, що Клавдою зветься, і човна насилу затримати змогли.
ACTS|27|17|Коли ж його витягли, то засобів допомічних добирали й корабля підв'язали. А боявшись, щоб не впасти на Сірт, поспускали вітрила, і носилися так.
ACTS|27|18|А коли зачала буря міцно нас кидати, то другого дня стали ми розвантажуватись,
ACTS|27|19|а третього дня корабельне знаряддя ми повикидали власноруч.
ACTS|27|20|А коли довгі дні не з'являлось ні сонце, ні зорі, і буря чимала на нас напирала, то останню надію ми втратили, щоб нам урятуватись...
ACTS|27|21|А як довго не їли вони, то Павло став тоді серед них і промовив: О мужі, тож треба було мене слухатися та не відпливати від Кріту, і обминули б були ці терпіння та шкоди.
ACTS|27|22|А тепер вас благаю триматись на дусі, бо ні одна душа з вас не згине, окрім корабля.
ACTS|27|23|Бо ночі цієї з'явився мені Ангол Бога, Якому належу й Якому служу,
ACTS|27|24|та і прорік: Не бійся, Павле, бо треба тобі перед кесарем стати, і ось Бог дарував тобі всіх, хто з тобою пливе.
ACTS|27|25|Тому то тримайтесь на дусі, о мужі, бо я вірую Богові, що станеться так, як було мені сказано.
ACTS|27|26|І ми мусимо наткнутись на острів якійсь.
ACTS|27|27|А коли надійшла чотирнадцята ніч, і ми носились по Адріятицькому морю, то десь коло півночі стали домислюватись моряки, що наближуються до якоїсь землі.
ACTS|27|28|І, запустивши оливницю, двадцять сяжнів знайшли. А від'їхавши трохи, запустити оливницю знову, і знайшли сяжнів п'ятнадцять.
ACTS|27|29|І боявшись, щоб не натрапити нам на скелясті місця, ми закинули чотири кітві з корми, і благали, щоб настав день.
ACTS|27|30|А коли моряки намагались утекти з корабля, і човна спускали до моря, вдаючи, ніби кітви закинути з носа хочуть,
ACTS|27|31|то сказав Павло сотникові й воякам: Як вони в кораблі не зостануться, то спастись ви не зможете!
ACTS|27|32|Тоді вояки перерізали мотузи в човна, і дали йому впасти.
ACTS|27|33|А коли розвиднятися стало, то благав Павло всіх, щоб поживу прийняти, і казав: Чотирнадцятий день ось сьогодні без їжі ви перебуваєте, очікуючи та нічого не ївши.
ACTS|27|34|Тому то благаю вас їжу прийняти, бо це на рятунок вам буде, бо жадному з вас не спаде з голови й волосина!
ACTS|27|35|А промовивши це, узяв хліб та подякував Богові перед усіма, і, поламавши, став їсти.
ACTS|27|36|Тоді всі піднеслись на дусі, і, стали поживу приймати.
ACTS|27|37|А всіх душ нас було в кораблі двісті сімдесят шість.
ACTS|27|38|І як наїлись вони, то стали полегшувати корабля, викидаючи збіжжя до моря.
ACTS|27|39|А коли настав день, то вони не могли розпізнати землі, одначе затоку якусь там угледіли, що берега плаского мала, до якого й вирішили, як можна, приплисти з кораблем.
ACTS|27|40|Підняли тоді кітви, і повкидали до моря, і порозв'язували поворозки в стерна, і вітрило мале за вітром поставили, та й покерували до берега.
ACTS|27|41|Та ось ми натрапили на місце, що мало з обох сторін море, і корабель опинивсь на мілкому: ніс загруз й позоставсь нерухомий, а корма розбивалася силою хвиль...
ACTS|27|42|Вояки ж були змовилися повбивати в'язнів, щоб котрийсь не поплив і не втік.
ACTS|27|43|Але сотник хотів урятувати Павла, і заборонив їхній намір, і звелів усім тим, хто пливати вміє, щоб скакали та перші на берег виходили,
ACTS|27|44|а інші хто на дошках, а хто на чімбудь з корабля. І таким чином сталось, що всі врятувались на землю!
ACTS|28|1|А коли врятувалися ми, то довідалися, що острів той зветься Меліта.
ACTS|28|2|Тубільці ж нам виявили надзвичайну людяність, бо вони запалили огонь, ішов бо дощ і був холод, і прийняли нас усіх.
ACTS|28|3|Як Павло ж назбирав купу хмизу та й поклав на огонь, змія вискочила через жар, і почепилась на руку йому...
ACTS|28|4|Як тубільці ж угледіли, що змія почепилась на руку йому, зачали говорити один одному: Либонь цей чоловік душогуб, що йому, від моря врятованому, Помста жити не дозволила!
ACTS|28|5|Він струснув ту звірюку в огонь, і ніякої шкоди не зазнав!
ACTS|28|6|А вони сподівалися, що він спухне або впаде мертвий умить. Коли ж довго чекали того та побачили, що ніякого лиха не сталося з ним, думку змінили й казали, що він бог...
ACTS|28|7|Навкруги ж того місця знаходились, добра начальника острова, на ім'я Публія, він прийняв нас, і три дні ласкаво гостив.
ACTS|28|8|І сталось, що Публіїв батько лежав, слабий на пропасницю та на червінку. До нього Павло ввійшов і помолився, і, руки на нього поклавши, уздоровив його.
ACTS|28|9|Якже трапилось це, то й інші на острові, що мали хвороби, приходили та вздоровлялись.
ACTS|28|10|Вони нас вшанували й великими почестями, а як ми від'їжджали, понакладали, чого було треба.
ACTS|28|11|А по трьох місяцях ми відпливли на олександрійському кораблі, що мав знака братів Діоскурів, і що на острові він перезимував.
ACTS|28|12|І, як ми допливли в Сіракузи, пробули там три дні.
ACTS|28|13|А звідти, пливучи понад берегом, прибули ми до Реґії, а що вітер південний повіяв за день, то другого дня прибули в Путеолі,
ACTS|28|14|де знайшли ми братів, вони ж нас ублагали сім день позостатися в них. І ось так прибули ми до Риму.
ACTS|28|15|А звідти брати, прочувши про нас, назустріч нам вийшли аж до Аппіфору та до Тритаверни. Побачивши їх, Павло дякував Богові та посмілішав.
ACTS|28|16|А коли прибули ми до Риму, Павлові дозволено жити осібно, ураз із вояком, що його сторожив.
ACTS|28|17|І сталось, по трьох днях Павло скликав знатніших з юдеїв. Як зійшлися ж вони, він промовив до них: Мужі-браття! Не вчинив я нічого проти люду чи звичаїв отцівських, та проте мене видано з Єрусалиму ув'язненого в руки римлян.
ACTS|28|18|Вони мене вислухали та й хотіли пустити, бож провини смертельної ні однієї в мені не було.
ACTS|28|19|Та юдеї противилися, тому змушений був я відкликатися на суд кесарів, але не для того, щоб народ свій у чомусь оскаржити.
ACTS|28|20|Тож із цієї причини покликав я вас, щоб побачити й порозмовляти, бо то за надію Ізраїлеву я обкутий цими кайданами...
ACTS|28|21|А вони відказали йому: Не одержали ми ні листів із Юдеї про тебе, ані жоден із братів не прийшов, і не звістив, і не казав чого злого про тебе.
ACTS|28|22|Але прагнемо ми, щоб почути від тебе, яку думку ти маєш, бо відомо про секту цю нам, що їй скрізь спротивляються.
ACTS|28|23|А коли вони визначили йому день, то дуже багато прийшло їх до нього в господу. А він їм від ранку до вечора розповідав, та про Божеє Царство свідоцтва давав, і переконував їх про Ісуса Законом Мойсея й Пророками.
ACTS|28|24|І одні вірили в те, про що він говорив, а інші не вірили.
ACTS|28|25|Вони між собою незгідні були й повиходили, як промовив Павло одне слово, що добре прорік Дух Святий отцям нашим через пророка Ісаю,
ACTS|28|26|промовляючи: Піди до народу цього та й скажи: Ви вухом почуєте, та розуміти не будете, дивитися будете оком, але не побачите!
ACTS|28|27|Затовстіло бо серце людей цих, тяжко чують на вуха вони, і зажмурили очі свої, щоб якось не побачити очима, і не почути вухами, і не зрозуміти їм серцем, і не навернутись, щоб Я їх уздоровив!
ACTS|28|28|Тож нехай для вас буде відоме, що послано Боже спасіння оце до поган, і почують вони!
ACTS|28|29|Як промовив він це, розійшлися юдеї, велику суперечку провадивши поміж собою.
ACTS|28|30|І цілих два роки Павло пробув у найнятім домі своїм, і приймав усіх, хто приходив до нього,
ACTS|28|31|і проповідував він Боже Царство, та з відвагою повною беззаборонно навчав про Господа Ісуса Христа!
