ACTS|1|1|primum quidem sermonem feci de omnibus o Theophile quae coepit Iesus facere et docere
ACTS|1|2|usque in diem qua praecipiens apostolis per Spiritum Sanctum quos elegit adsumptus est
ACTS|1|3|quibus et praebuit se ipsum vivum post passionem suam in multis argumentis per dies quadraginta apparens eis et loquens de regno Dei
ACTS|1|4|et convescens praecepit eis ab Hierosolymis ne discederent sed expectarent promissionem Patris quam audistis per os meum
ACTS|1|5|quia Iohannes quidem baptizavit aqua vos autem baptizabimini Spiritu Sancto non post multos hos dies
ACTS|1|6|igitur qui convenerant interrogabant eum dicentes Domine si in tempore hoc restitues regnum Israhel
ACTS|1|7|dixit autem eis non est vestrum nosse tempora vel momenta quae Pater posuit in sua potestate
ACTS|1|8|sed accipietis virtutem supervenientis Spiritus Sancti in vos et eritis mihi testes in Hierusalem et in omni Iudaea et Samaria et usque ad ultimum terrae
ACTS|1|9|et cum haec dixisset videntibus illis elevatus est et nubes suscepit eum ab oculis eorum
ACTS|1|10|cumque intuerentur in caelum eunte illo ecce duo viri adstiterunt iuxta illos in vestibus albis
ACTS|1|11|qui et dixerunt viri galilaei quid statis aspicientes in caelum hic Iesus qui adsumptus est a vobis in caelum sic veniet quemadmodum vidistis eum euntem in caelum
ACTS|1|12|tunc reversi sunt Hierosolymam a monte qui vocatur Oliveti qui est iuxta Hierusalem sabbati habens iter
ACTS|1|13|et cum introissent in cenaculum ascenderunt ubi manebant Petrus et Iohannes Iacobus et Andreas Philippus et Thomas Bartholomeus et Mattheus Iacobus Alphei et Simon Zelotes et Iudas Iacobi
ACTS|1|14|hii omnes erant perseverantes unianimiter in oratione cum mulieribus et Maria matre Iesu et fratribus eius
ACTS|1|15|et in diebus illis exsurgens Petrus in medio fratrum dixit erat autem turba nominum simul fere centum viginti
ACTS|1|16|viri fratres oportet impleri scripturam quam praedixit Spiritus Sanctus per os David de Iuda qui fuit dux eorum qui conprehenderunt Iesum
ACTS|1|17|quia connumeratus erat in nobis et sortitus est sortem ministerii huius
ACTS|1|18|et hic quidem possedit agrum de mercede iniquitatis et suspensus crepuit medius et diffusa sunt omnia viscera eius
ACTS|1|19|et notum factum est omnibus habitantibus Hierusalem ita ut appellaretur ager ille lingua eorum Acheldemach hoc est ager Sanguinis
ACTS|1|20|scriptum est enim in libro Psalmorum fiat commoratio eius deserta et non sit qui inhabitet in ea et episcopatum eius accipiat alius
ACTS|1|21|oportet ergo ex his viris qui nobiscum congregati sunt in omni tempore quo intravit et exivit inter nos Dominus Iesus
ACTS|1|22|incipiens a baptismate Iohannis usque in diem qua adsumptus est a nobis testem resurrectionis eius nobiscum fieri unum ex istis
ACTS|1|23|et statuerunt duos Ioseph qui vocabatur Barsabban qui cognominatus est Iustus et Matthiam
ACTS|1|24|et orantes dixerunt tu Domine qui corda nosti omnium ostende quem elegeris ex his duobus unum
ACTS|1|25|accipere locum ministerii huius et apostolatus de quo praevaricatus est Iudas ut abiret in locum suum
ACTS|1|26|et dederunt sortes eis et cecidit sors super Matthiam et adnumeratus est cum undecim apostolis
ACTS|2|1|et cum conplerentur dies pentecostes erant omnes pariter in eodem loco
ACTS|2|2|et factus est repente de caelo sonus tamquam advenientis spiritus vehementis et replevit totam domum ubi erant sedentes
ACTS|2|3|et apparuerunt illis dispertitae linguae tamquam ignis seditque supra singulos eorum
ACTS|2|4|et repleti sunt omnes Spiritu Sancto et coeperunt loqui aliis linguis prout Spiritus Sanctus dabat eloqui illis
ACTS|2|5|erant autem in Hierusalem habitantes Iudaei viri religiosi ex omni natione quae sub caelo sunt
ACTS|2|6|facta autem hac voce convenit multitudo et mente confusa est quoniam audiebat unusquisque lingua sua illos loquentes
ACTS|2|7|stupebant autem omnes et mirabantur dicentes nonne omnes ecce isti qui loquuntur Galilaei sunt
ACTS|2|8|et quomodo nos audivimus unusquisque lingua nostra in qua nati sumus
ACTS|2|9|Parthi et Medi et Elamitae et qui habitant Mesopotamiam et Iudaeam et Cappadociam Pontum et Asiam
ACTS|2|10|Frygiam et Pamphiliam Aegyptum et partes Lybiae quae est circa Cyrenen et advenae romani
ACTS|2|11|Iudaei quoque et proselyti Cretes et Arabes audivimus loquentes eos nostris linguis magnalia Dei
ACTS|2|12|stupebant autem omnes et mirabantur ad invicem dicentes quidnam hoc vult esse
ACTS|2|13|alii autem inridentes dicebant quia musto pleni sunt isti
ACTS|2|14|stans autem Petrus cum undecim levavit vocem suam et locutus est eis viri iudaei et qui habitatis Hierusalem universi hoc vobis notum sit et auribus percipite verba mea
ACTS|2|15|non enim sicut vos aestimatis hii ebrii sunt cum sit hora diei tertia
ACTS|2|16|sed hoc est quod dictum est per prophetam Iohel
ACTS|2|17|et erit in novissimis diebus dicit Dominus effundam de Spiritu meo super omnem carnem et prophetabunt filii vestri et filiae vestrae et iuvenes vestri visiones videbunt et seniores vestri somnia somniabunt
ACTS|2|18|et quidem super servos meos et super ancillas meas in diebus illis effundam de Spiritu meo et prophetabunt
ACTS|2|19|et dabo prodigia in caelo sursum et signa in terra deorsum sanguinem et ignem et vaporem fumi
ACTS|2|20|sol convertetur in tenebras et luna in sanguinem antequam veniat dies Domini magnus et manifestus
ACTS|2|21|et erit omnis quicumque invocaverit nomen Domini salvus erit
ACTS|2|22|viri israhelitae audite verba haec Iesum Nazarenum virum adprobatum a Deo in vobis virtutibus et prodigiis et signis quae fecit per illum Deus in medio vestri sicut vos scitis
ACTS|2|23|hunc definito consilio et praescientia Dei traditum per manus iniquorum adfigentes interemistis
ACTS|2|24|quem Deus suscitavit solutis doloribus inferni iuxta quod inpossibile erat teneri illum ab eo
ACTS|2|25|David enim dicit in eum providebam Dominum coram me semper quoniam a dextris meis est ne commovear
ACTS|2|26|propter hoc laetatum est cor meum et exultavit lingua mea insuper et caro mea requiescet in spe
ACTS|2|27|quoniam non derelinques animam meam in inferno neque dabis Sanctum tuum videre corruptionem
ACTS|2|28|notas fecisti mihi vias vitae replebis me iucunditate cum facie tua
ACTS|2|29|viri fratres liceat audenter dicere ad vos de patriarcha David quoniam et defunctus est et sepultus est et sepulchrum eius est apud nos usque in hodiernum diem
ACTS|2|30|propheta igitur cum esset et sciret quia iureiurando iurasset illi Deus de fructu lumbi eius sedere super sedem eius
ACTS|2|31|providens locutus est de resurrectione Christi quia neque derelictus est in inferno neque caro eius vidit corruptionem
ACTS|2|32|hunc Iesum resuscitavit Deus cui omnes nos testes sumus
ACTS|2|33|dextera igitur Dei exaltatus et promissione Spiritus Sancti accepta a Patre effudit hunc quem vos videtis et audistis
ACTS|2|34|non enim David ascendit in caelos dicit autem ipse dixit Dominus Domino meo sede a dextris meis
ACTS|2|35|donec ponam inimicos tuos scabillum pedum tuorum
ACTS|2|36|certissime ergo sciat omnis domus Israhel quia et Dominum eum et Christum Deus fecit hunc Iesum quem vos crucifixistis
ACTS|2|37|his auditis conpuncti sunt corde et dixerunt ad Petrum et ad reliquos apostolos quid faciemus viri fratres
ACTS|2|38|Petrus vero ad illos paenitentiam inquit agite et baptizetur unusquisque vestrum in nomine Iesu Christi in remissionem peccatorum vestrorum et accipietis donum Sancti Spiritus
ACTS|2|39|vobis enim est repromissio et filiis vestris et omnibus qui longe sunt quoscumque advocaverit Dominus Deus noster
ACTS|2|40|aliis etiam verbis pluribus testificatus est et exhortabatur eos dicens salvamini a generatione ista prava
ACTS|2|41|qui ergo receperunt sermonem eius baptizati sunt et adpositae sunt in illa die animae circiter tria milia
ACTS|2|42|erant autem perseverantes in doctrina apostolorum et communicatione fractionis panis et orationibus
ACTS|2|43|fiebat autem omni animae timor multa quoque prodigia et signa per apostolos fiebant in Hierusalem et metus erat magnus in universis
ACTS|2|44|omnes etiam qui credebant erant pariter et habebant omnia communia
ACTS|2|45|possessiones et substantias vendebant et dividebant illa omnibus prout cuique opus erat
ACTS|2|46|cotidie quoque perdurantes unianimiter in templo et frangentes circa domos panem sumebant cibum cum exultatione et simplicitate cordis
ACTS|2|47|conlaudantes Deum et habentes gratiam ad omnem plebem Dominus autem augebat qui salvi fierent cotidie in id ipsum
ACTS|3|1|Petrus autem et Iohannes ascendebant in templum ad horam orationis nonam
ACTS|3|2|et quidam vir qui erat claudus ex utero matris suae baiulabatur quem ponebant cotidie ad portam templi quae dicitur Speciosa ut peteret elemosynam ab introeuntibus in templum
ACTS|3|3|is cum vidisset Petrum et Iohannem incipientes introire in templum rogabat ut elemosynam acciperet
ACTS|3|4|intuens autem in eum Petrus cum Iohanne dixit respice in nos
ACTS|3|5|at ille intendebat in eos sperans se aliquid accepturum ab eis
ACTS|3|6|Petrus autem dixit argentum et aurum non est mihi quod autem habeo hoc tibi do in nomine Iesu Christi Nazareni surge et ambula
ACTS|3|7|et adprehensa ei manu dextera adlevavit eum et protinus consolidatae sunt bases eius et plantae
ACTS|3|8|et exiliens stetit et ambulabat et intravit cum illis in templum ambulans et exiliens et laudans Dominum
ACTS|3|9|et vidit omnis populus eum ambulantem et laudantem Deum
ACTS|3|10|cognoscebant autem illum quoniam ipse erat qui ad elemosynam sedebat ad Speciosam portam templi et impleti sunt stupore et extasi in eo quod contigerat illi
ACTS|3|11|cum teneret autem Petrum et Iohannem concurrit omnis populus ad eos ad porticum qui appellatur Salomonis stupentes
ACTS|3|12|videns autem Petrus respondit ad populum viri israhelitae quid miramini in hoc aut nos quid intuemini quasi nostra virtute aut pietate fecerimus hunc ambulare
ACTS|3|13|Deus Abraham et Deus Isaac et Deus Iacob Deus patrum nostrorum glorificavit Filium suum Iesum quem vos quidem tradidistis et negastis ante faciem Pilati iudicante illo dimitti
ACTS|3|14|vos autem sanctum et iustum negastis et petistis virum homicidam donari vobis
ACTS|3|15|auctorem vero vitae interfecistis quem Deus suscitavit a mortuis cuius nos testes sumus
ACTS|3|16|et in fide nominis eius hunc quem videtis et nostis confirmavit nomen eius et fides quae per eum est dedit integram sanitatem istam in conspectu omnium vestrum
ACTS|3|17|et nunc fratres scio quia per ignorantiam fecistis sicut et principes vestri
ACTS|3|18|Deus autem quae praenuntiavit per os omnium prophetarum pati Christum suum implevit sic
ACTS|3|19|paenitemini igitur et convertimini ut deleantur vestra peccata
ACTS|3|20|ut cum venerint tempora refrigerii a conspectu Domini et miserit eum qui praedicatus est vobis Iesum Christum
ACTS|3|21|quem oportet caelum quidem suscipere usque in tempora restitutionis omnium quae locutus est Deus per os sanctorum suorum a saeculo prophetarum
ACTS|3|22|Moses quidem dixit quia prophetam vobis suscitabit Dominus Deus vester de fratribus vestris tamquam me ipsum audietis iuxta omnia quaecumque locutus fuerit vobis
ACTS|3|23|erit autem omnis anima quae non audierit prophetam illum exterminabitur de plebe
ACTS|3|24|et omnes prophetae a Samuhel et deinceps qui locuti sunt et adnuntiaverunt dies istos
ACTS|3|25|vos estis filii prophetarum et testamenti quod disposuit Deus ad patres vestros dicens ad Abraham et in semine tuo benedicentur omnes familiae terrae
ACTS|3|26|vobis primum Deus suscitans Filium suum misit eum benedicentem vobis ut convertat se unusquisque a nequitia sua
ACTS|4|1|loquentibus autem illis ad populum supervenerunt sacerdotes et magistratus templi et Sadducaei
ACTS|4|2|dolentes quod docerent populum et adnuntiarent in Iesu resurrectionem ex mortuis
ACTS|4|3|et iniecerunt in eis manus et posuerunt eos in custodiam in crastinum erat enim iam vespera
ACTS|4|4|multi autem eorum qui audierant verbum crediderunt et factus est numerus virorum quinque milia
ACTS|4|5|factum est autem in crastinum ut congregarentur principes eorum et seniores et scribae in Hierusalem
ACTS|4|6|et Annas princeps sacerdotum et Caiphas et Iohannes et Alexander et quotquot erant de genere sacerdotali
ACTS|4|7|et statuentes eos in medio interrogabant in qua virtute aut in quo nomine fecistis hoc vos
ACTS|4|8|tunc Petrus repletus Spiritu Sancto dixit ad eos principes populi et seniores
ACTS|4|9|si nos hodie diiudicamur in benefacto hominis infirmi in quo iste salvus factus est
ACTS|4|10|notum sit omnibus vobis et omni plebi Israhel quia in nomine Iesu Christi Nazareni quem vos crucifixistis quem Deus suscitavit a mortuis in hoc iste adstat coram vobis sanus
ACTS|4|11|hic est lapis qui reprobatus est a vobis aedificantibus qui factus est in caput anguli
ACTS|4|12|et non est in alio aliquo salus nec enim nomen aliud est sub caelo datum hominibus in quo oportet nos salvos fieri
ACTS|4|13|videntes autem Petri constantiam et Iohannis conperto quod homines essent sine litteris et idiotae admirabantur et cognoscebant eos quoniam cum Iesu fuerant
ACTS|4|14|hominem quoque videntes stantem cum eis qui curatus fuerat nihil poterant contradicere
ACTS|4|15|iusserunt autem eos foras extra concilium secedere et conferebant ad invicem
ACTS|4|16|dicentes quid faciemus hominibus istis quoniam quidem notum signum factum est per eos omnibus habitantibus in Hierusalem manifestum et non possumus negare
ACTS|4|17|sed ne amplius divulgetur in populum comminemur eis ne ultra loquantur in nomine hoc ulli hominum
ACTS|4|18|et vocantes eos denuntiaverunt ne omnino loquerentur neque docerent in nomine Iesu
ACTS|4|19|Petrus vero et Iohannes respondentes dixerunt ad eos si iustum est in conspectu Dei vos potius audire quam Deum iudicate
ACTS|4|20|non enim possumus quae vidimus et audivimus non loqui
ACTS|4|21|at illi comminantes dimiserunt eos non invenientes quomodo punirent eos propter populum quia omnes clarificabant Deum in eo quod acciderat
ACTS|4|22|annorum enim erat amplius quadraginta homo in quo factum erat signum istud sanitatis
ACTS|4|23|dimissi autem venerunt ad suos et adnuntiaverunt eis quanta ad eos principes sacerdotum et seniores dixissent
ACTS|4|24|qui cum audissent unianimiter levaverunt vocem ad Deum et dixerunt Domine tu qui fecisti caelum et terram et mare et omnia quae in eis sunt
ACTS|4|25|qui Spiritu Sancto per os patris nostri David pueri tui dixisti quare fremuerunt gentes et populi meditati sunt inania
ACTS|4|26|adstiterunt reges terrae et principes convenerunt in unum adversus Dominum et adversus Christum eius
ACTS|4|27|convenerunt enim vere in civitate ista adversus sanctum puerum tuum Iesum quem unxisti Herodes et Pontius Pilatus cum gentibus et populis Israhel
ACTS|4|28|facere quae manus tua et consilium decreverunt fieri
ACTS|4|29|et nunc Domine respice in minas eorum et da servis tuis cum omni fiducia loqui verbum tuum
ACTS|4|30|in eo cum manum tuam extendas sanitates et signa et prodigia fieri per nomen sancti Filii tui Iesu
ACTS|4|31|et cum orassent motus est locus in quo erant congregati et repleti sunt omnes Spiritu Sancto et loquebantur verbum Dei cum fiducia
ACTS|4|32|multitudinis autem credentium erat cor et anima una nec quisquam eorum quae possidebant aliquid suum esse dicebat sed erant illis omnia communia
ACTS|4|33|et virtute magna reddebant apostoli testimonium resurrectionis Iesu Christi Domini et gratia magna erat in omnibus illis
ACTS|4|34|neque enim quisquam egens erat inter illos quotquot enim possessores agrorum aut domorum erant vendentes adferebant pretia eorum quae vendebant
ACTS|4|35|et ponebant ante pedes apostolorum dividebantur autem singulis prout cuique opus erat
ACTS|4|36|Ioseph autem qui cognominatus est Barnabas ab apostolis quod est interpretatum Filius consolationis Levites Cyprius genere
ACTS|4|37|cum haberet agrum vendidit illum et adtulit pretium et posuit ante pedes apostolorum
ACTS|5|1|vir autem quidam nomine Ananias cum Saffira uxore sua vendidit agrum
ACTS|5|2|et fraudavit de pretio agri conscia uxore sua et adferens partem quandam ad pedes apostolorum posuit
ACTS|5|3|dixit autem Petrus Anania cur temptavit Satanas cor tuum mentiri te Spiritui Sancto et fraudare de pretio agri
ACTS|5|4|nonne manens tibi manebat et venundatum in tua erat potestate quare posuisti in corde tuo hanc rem non es mentitus hominibus sed Deo
ACTS|5|5|audiens autem Ananias haec verba cecidit et exspiravit et factus est timor magnus in omnes qui audierant
ACTS|5|6|surgentes autem iuvenes amoverunt eum et efferentes sepelierunt
ACTS|5|7|factum est autem quasi horarum trium spatium et uxor ipsius nesciens quod factum fuerat introiit
ACTS|5|8|respondit autem ei Petrus dic mihi si tanti agrum vendidistis at illa dixit etiam tanti
ACTS|5|9|Petrus autem ad eam quid utique convenit vobis temptare Spiritum Domini ecce pedes eorum qui sepelierunt virum tuum ad ostium et efferent te
ACTS|5|10|confestim cecidit ante pedes eius et exspiravit intrantes autem iuvenes invenerunt illam mortuam et extulerunt et sepelierunt ad virum suum
ACTS|5|11|et factus est timor magnus in universa ecclesia et in omnes qui audierunt haec
ACTS|5|12|per manus autem apostolorum fiebant signa et prodigia multa in plebe et erant unianimiter omnes in porticu Salomonis
ACTS|5|13|ceterorum autem nemo audebat coniungere se illis sed magnificabat eos populus
ACTS|5|14|magis autem augebatur credentium in Domino multitudo virorum ac mulierum
ACTS|5|15|ita ut in plateas eicerent infirmos et ponerent in lectulis et grabattis ut veniente Petro saltim umbra illius obumbraret quemquam eorum
ACTS|5|16|concurrebat autem et multitudo vicinarum civitatum Hierusalem adferentes aegros et vexatos ab spiritibus inmundis qui curabantur omnes
ACTS|5|17|exsurgens autem princeps sacerdotum et omnes qui cum illo erant quae est heresis Sadducaeorum repleti sunt zelo
ACTS|5|18|et iniecerunt manus in apostolos et posuerunt illos in custodia publica
ACTS|5|19|angelus autem Domini per noctem aperiens ianuas carceris et educens eos dixit
ACTS|5|20|ite et stantes loquimini in templo plebi omnia verba vitae huius
ACTS|5|21|qui cum audissent intraverunt diluculo in templum et docebant adveniens autem princeps sacerdotum et qui cum eo erant convocaverunt concilium et omnes seniores filiorum Israhel et miserunt in carcerem ut adducerentur
ACTS|5|22|cum venissent autem ministri et aperto carcere non invenissent illos reversi nuntiaverunt
ACTS|5|23|dicentes carcerem quidem invenimus clausum cum omni diligentia et custodes stantes ad ianuas aperientes autem neminem intus invenimus
ACTS|5|24|ut audierunt autem hos sermones magistratus templi et principes sacerdotum ambigebant de illis quidnam fieret
ACTS|5|25|adveniens autem quidam nuntiavit eis quia ecce viri quos posuistis in carcere sunt in templo stantes et docentes populum
ACTS|5|26|tunc abiit magistratus cum ministris et adduxit illos sine vi timebant enim populum ne lapidarentur
ACTS|5|27|et cum adduxissent illos statuerunt in concilio et interrogavit eos princeps sacerdotum
ACTS|5|28|dicens praecipiendo praecepimus vobis ne doceretis in nomine isto et ecce replestis Hierusalem doctrina vestra et vultis inducere super nos sanguinem hominis istius
ACTS|5|29|respondens autem Petrus et apostoli dixerunt oboedire oportet Deo magis quam hominibus
ACTS|5|30|Deus patrum nostrorum suscitavit Iesum quem vos interemistis suspendentes in ligno
ACTS|5|31|hunc Deus principem et salvatorem exaltavit dextera sua ad dandam paenitentiam Israhel et remissionem peccatorum
ACTS|5|32|et nos sumus testes horum verborum et Spiritus Sanctus quem dedit Deus omnibus oboedientibus sibi
ACTS|5|33|haec cum audissent dissecabantur et cogitabant interficere illos
ACTS|5|34|surgens autem quidam in concilio Pharisaeus nomine Gamalihel legis doctor honorabilis universae plebi iussit foras ad breve homines fieri
ACTS|5|35|dixitque ad illos viri israhelitae adtendite vobis super hominibus istis quid acturi sitis
ACTS|5|36|ante hos enim dies extitit Theodas dicens esse se aliquem cui consensit virorum numerus circiter quadringentorum qui occisus est et omnes quicumque credebant ei dissipati sunt et redactus est ad nihilum
ACTS|5|37|post hunc extitit Iudas Galilaeus in diebus professionis et avertit populum post se et ipse periit et omnes quotquot consenserunt ei dispersi sunt
ACTS|5|38|et nunc itaque dico vobis discedite ab hominibus istis et sinite illos quoniam si est ex hominibus consilium hoc aut opus dissolvetur
ACTS|5|39|si vero ex Deo est non poteritis dissolvere eos ne forte et Deo repugnare inveniamini consenserunt autem illi
ACTS|5|40|et convocantes apostolos caesis denuntiaverunt ne loquerentur in nomine Iesu et dimiserunt eos
ACTS|5|41|et illi quidem ibant gaudentes a conspectu concilii quoniam digni habiti sunt pro nomine Iesu contumeliam pati
ACTS|5|42|omni autem die in templo et circa domos non cessabant docentes et evangelizantes Christum Iesum
ACTS|6|1|in diebus autem illis crescente numero discipulorum factus est murmur Graecorum adversus Hebraeos eo quod dispicerentur in ministerio cotidiano viduae eorum
ACTS|6|2|convocantes autem duodecim multitudinem discipulorum dixerunt non est aequum nos derelinquere verbum Dei et ministrare mensis
ACTS|6|3|considerate ergo fratres viros ex vobis boni testimonii septem plenos Spiritu et sapientia quos constituamus super hoc opus
ACTS|6|4|nos vero orationi et ministerio verbi instantes erimus
ACTS|6|5|et placuit sermo coram omni multitudine et elegerunt Stephanum virum plenum fide et Spiritu Sancto et Philippum et Prochorum et Nicanorem et Timonem et Parmenam et Nicolaum advenam Antiochenum
ACTS|6|6|hos statuerunt ante conspectum apostolorum et orantes inposuerunt eis manus
ACTS|6|7|et verbum Dei crescebat et multiplicabatur numerus discipulorum in Hierusalem valde multa etiam turba sacerdotum oboediebat fidei
ACTS|6|8|Stephanus autem plenus gratia et fortitudine faciebat prodigia et signa magna in populo
ACTS|6|9|surrexerunt autem quidam de synagoga quae appellatur Libertinorum et Cyrenensium et Alexandrinorum et eorum qui erant a Cilicia et Asia disputantes cum Stephano
ACTS|6|10|et non poterant resistere sapientiae et Spiritui quo loquebatur
ACTS|6|11|tunc submiserunt viros qui dicerent se audisse eum dicentem verba blasphemiae in Mosen et Deum
ACTS|6|12|commoverunt itaque plebem et seniores et scribas et concurrentes rapuerunt eum et adduxerunt in concilium
ACTS|6|13|et statuerunt testes falsos dicentes homo iste non cessat loqui verba adversus locum sanctum et legem
ACTS|6|14|audivimus enim eum dicentem quoniam Iesus Nazarenus hic destruet locum istum et mutabit traditiones quas tradidit nobis Moses
ACTS|6|15|et intuentes eum omnes qui sedebant in concilio viderunt faciem eius tamquam faciem angeli
ACTS|7|1|dixit autem princeps sacerdotum si haec ita se habent
ACTS|7|2|qui ait viri fratres et patres audite Deus gloriae apparuit patri nostro Abraham cum esset in Mesopotamiam priusquam moraretur in Charram
ACTS|7|3|et dixit ad illum exi de terra tua et de cognatione tua et veni in terram quam tibi monstravero
ACTS|7|4|tunc exiit de terra Chaldeorum et habitavit in Charram et inde postquam mortuus est pater eius transtulit illum in terram istam in qua nunc vos habitatis
ACTS|7|5|et non dedit illi hereditatem in ea nec passum pedis et repromisit dare illi eam in possessionem et semini eius post ipsum cum non haberet filium
ACTS|7|6|locutus est autem Deus quia erit semen eius accola in terra aliena et servituti eos subicient et male tractabunt eos annis quadringentis
ACTS|7|7|et gentem cui servierint iudicabo ego dixit Deus et post haec exibunt et deservient mihi in loco isto
ACTS|7|8|et dedit illi testamentum circumcisionis et sic genuit Isaac et circumcidit eum die octava et Isaac Iacob et Iacob duodecim patriarchas
ACTS|7|9|et patriarchae aemulantes Ioseph vendiderunt in Aegyptum et erat Deus cum eo
ACTS|7|10|et eripuit eum ex omnibus tribulationibus eius et dedit ei gratiam et sapientiam in conspectu Pharaonis regis Aegypti et constituit eum praepositum super Aegyptum et super omnem domum suam
ACTS|7|11|venit autem fames in universam Aegyptum et Chanaan et tribulatio magna et non inveniebant cibos patres nostri
ACTS|7|12|cum audisset autem Iacob esse frumentum in Aegypto misit patres nostros primum
ACTS|7|13|et in secundo cognitus est Ioseph a fratribus suis et manifestatum est Pharaoni genus eius
ACTS|7|14|mittens autem Ioseph accersivit Iacob patrem suum et omnem cognationem in animabus septuaginta quinque
ACTS|7|15|et descendit Iacob in Aegyptum et defunctus est ipse et patres nostri
ACTS|7|16|et translati sunt in Sychem et positi sunt in sepulchro quod emit Abraham pretio argenti a filiis Emmor filii Sychem
ACTS|7|17|cum adpropinquaret autem tempus repromissionis quam confessus erat Deus Abrahae crevit populus et multiplicatus est in Aegypto
ACTS|7|18|quoadusque surrexit rex alius in Aegypto qui non sciebat Ioseph
ACTS|7|19|hic circumveniens genus nostrum adflixit patres ut exponerent infantes suos ne vivificarentur
ACTS|7|20|eodem tempore natus est Moses et fuit gratus Deo qui nutritus est tribus mensibus in domo patris sui
ACTS|7|21|exposito autem illo sustulit eum filia Pharaonis et enutrivit eum sibi in filium
ACTS|7|22|et eruditus est Moses omni sapientia Aegyptiorum et erat potens in verbis et in operibus suis
ACTS|7|23|cum autem impleretur ei quadraginta annorum tempus ascendit in cor eius ut visitaret fratres suos filios Israhel
ACTS|7|24|et cum vidisset quendam iniuriam patientem vindicavit illum et fecit ultionem ei qui iniuriam sustinebat percusso Aegyptio
ACTS|7|25|existimabat autem intellegere fratres quoniam Deus per manum ipsius daret salutem illis at illi non intellexerunt
ACTS|7|26|sequenti vero die apparuit illis litigantibus et reconciliabat eos in pacem dicens viri fratres estis ut quid nocetis alterutrum
ACTS|7|27|qui autem iniuriam faciebat proximo reppulit eum dicens quis te constituit principem et iudicem super nos
ACTS|7|28|numquid interficere me tu vis quemadmodum interfecisti heri Aegyptium
ACTS|7|29|fugit autem Moses in verbo isto et factus est advena in terra Madiam ubi generavit filios duos
ACTS|7|30|et expletis annis quadraginta apparuit illi in deserto montis Sina angelus in igne flammae rubi
ACTS|7|31|Moses autem videns admiratus est visum et accedente illo ut consideraret facta est vox Domini
ACTS|7|32|ego Deus patrum tuorum Deus Abraham et Deus Isaac et Deus Iacob tremefactus autem Moses non audebat considerare
ACTS|7|33|dixit autem illi Dominus solve calciamentum pedum tuorum locus enim in quo stas terra sancta est
ACTS|7|34|videns vidi adflictionem populi mei qui est in Aegypto et gemitum eorum audivi et descendi liberare eos et nunc veni et mittam te in Aegyptum
ACTS|7|35|hunc Mosen quem negaverunt dicentes quis te constituit principem et iudicem hunc Deus principem et redemptorem misit cum manu angeli qui apparuit illi in rubo
ACTS|7|36|hic eduxit illos faciens prodigia et signa in terra Aegypti et in Rubro mari et in deserto annis quadraginta
ACTS|7|37|hic est Moses qui dixit filiis Israhel prophetam vobis suscitabit Deus de fratribus vestris tamquam me
ACTS|7|38|hic est qui fuit in ecclesia in solitudine cum angelo qui loquebatur ei in monte Sina et cum patribus nostris qui accepit verba vitae dare nobis
ACTS|7|39|cui noluerunt oboedire patres nostri sed reppulerunt et aversi sunt cordibus suis in Aegyptum
ACTS|7|40|dicentes ad Aaron fac nobis deos qui praecedant nos Moses enim hic qui eduxit nos de terra Aegypti nescimus quid factum sit ei
ACTS|7|41|et vitulum fecerunt in illis diebus et obtulerunt hostiam simulacro et laetabantur in operibus manuum suarum
ACTS|7|42|convertit autem Deus et tradidit eos servire militiae caeli sicut scriptum est in libro Prophetarum numquid victimas aut hostias obtulistis mihi annis quadraginta in deserto domus Israhel
ACTS|7|43|et suscepistis tabernaculum Moloch et sidus dei vestri Rempham figuras quas fecistis adorare eas et transferam vos trans Babylonem
ACTS|7|44|tabernaculum testimonii fuit patribus nostris in deserto sicut disposuit loquens ad Mosen ut faceret illud secundum formam quam viderat
ACTS|7|45|quod et induxerunt suscipientes patres nostri cum Iesu in possessionem gentium quas expulit Deus a facie patrum nostrorum usque in diebus David
ACTS|7|46|qui invenit gratiam ante Deum et petiit ut inveniret tabernaculum Deo Iacob
ACTS|7|47|Salomon autem aedificavit illi domum
ACTS|7|48|sed non Excelsus in manufactis habitat sicut propheta dicit
ACTS|7|49|caelum mihi sedis est terra autem scabillum pedum meorum quam domum aedificabitis mihi dicit Dominus aut quis locus requietionis meae est
ACTS|7|50|nonne manus mea fecit haec omnia
ACTS|7|51|dura cervice et incircumcisi cordibus et auribus vos semper Spiritui Sancto resistitis sicut patres vestri et vos
ACTS|7|52|quem prophetarum non sunt persecuti patres vestri et occiderunt eos qui praenuntiabant de adventu Iusti cuius vos nunc proditores et homicidae fuistis
ACTS|7|53|qui accepistis legem in dispositionem angelorum et non custodistis
ACTS|7|54|audientes autem haec dissecabantur cordibus suis et stridebant dentibus in eum
ACTS|7|55|cum autem esset plenus Spiritu Sancto intendens in caelum vidit gloriam Dei et Iesum stantem a dextris Dei et ait ecce video caelos apertos et Filium hominis a dextris stantem Dei
ACTS|7|56|exclamantes autem voce magna continuerunt aures suas et impetum fecerunt unianimiter in eum
ACTS|7|57|et eicientes eum extra civitatem lapidabant et testes deposuerunt vestimenta sua secus pedes adulescentis qui vocabatur Saulus
ACTS|7|58|et lapidabant Stephanum invocantem et dicentem Domine Iesu suscipe spiritum meum
ACTS|7|59|positis autem genibus clamavit voce magna Domine ne statuas illis hoc peccatum et cum hoc dixisset obdormivit Saulus autem erat consentiens neci eius
ACTS|8|1|facta est autem in illa die persecutio magna in ecclesia quae erat Hierosolymis et omnes dispersi sunt per regiones Iudaeae et Samariae praeter apostolos
ACTS|8|2|curaverunt autem Stephanum viri timorati et fecerunt planctum magnum super illum
ACTS|8|3|Saulus vero devastabat ecclesiam per domos intrans et trahens viros ac mulieres tradebat in custodiam
ACTS|8|4|igitur qui dispersi erant pertransiebant evangelizantes verbum
ACTS|8|5|Philippus autem descendens in civitatem Samariae praedicabat illis Christum
ACTS|8|6|intendebant autem turbae his quae a Philippo dicebantur unianimiter audientes et videntes signa quae faciebat
ACTS|8|7|multi enim eorum qui habebant spiritus inmundos clamantes voce magna exiebant multi autem paralytici et claudi curati sunt
ACTS|8|8|factum est ergo magnum gaudium in illa civitate
ACTS|8|9|vir autem quidam nomine Simon qui ante fuerat in civitate magus seducens gentem Samariae dicens esse se aliquem magnum
ACTS|8|10|cui auscultabant omnes a minimo usque ad maximum dicentes hic est virtus Dei quae vocatur Magna
ACTS|8|11|adtendebant autem eum propter quod multo tempore magicis suis dementasset eos
ACTS|8|12|cum vero credidissent Philippo evangelizanti de regno Dei et nomine Iesu Christi baptizabantur viri ac mulieres
ACTS|8|13|tunc Simon et ipse credidit et cum baptizatus esset adherebat Philippo videns etiam signa et virtutes maximas fieri stupens admirabatur
ACTS|8|14|cum autem audissent apostoli qui erant Hierosolymis quia recepit Samaria verbum Dei miserunt ad illos Petrum et Iohannem
ACTS|8|15|qui cum venissent oraverunt pro ipsis ut acciperent Spiritum Sanctum
ACTS|8|16|nondum enim in quemquam illorum venerat sed baptizati tantum erant in nomine Domini Iesu
ACTS|8|17|tunc inponebant manus super illos et accipiebant Spiritum Sanctum
ACTS|8|18|cum vidisset autem Simon quia per inpositionem manus apostolorum daretur Spiritus Sanctus obtulit eis pecuniam
ACTS|8|19|dicens date et mihi hanc potestatem ut cuicumque inposuero manus accipiat Spiritum Sanctum Petrus autem dixit ad eum
ACTS|8|20|pecunia tua tecum sit in perditionem quoniam donum Dei existimasti pecunia possideri
ACTS|8|21|non est tibi pars neque sors in sermone isto cor enim tuum non est rectum coram Deo
ACTS|8|22|paenitentiam itaque age ab hac nequitia tua et roga Deum si forte remittatur tibi haec cogitatio cordis tui
ACTS|8|23|in felle enim amaritudinis et obligatione iniquitatis video te esse
ACTS|8|24|respondens autem Simon dixit precamini vos pro me ad Dominum ut nihil veniat super me horum quae dixistis
ACTS|8|25|et illi quidem testificati et locuti verbum Domini rediebant Hierosolymam et multis regionibus Samaritanorum evangelizabant
ACTS|8|26|angelus autem Domini locutus est ad Philippum dicens surge et vade contra meridianum ad viam quae descendit ab Hierusalem in Gazam haec est deserta
ACTS|8|27|et surgens abiit et ecce vir aethiops eunuchus potens Candacis reginae Aethiopum qui erat super omnes gazas eius venerat adorare in Hierusalem
ACTS|8|28|et revertebatur sedens super currum suum legensque prophetam Esaiam
ACTS|8|29|dixit autem Spiritus Philippo accede et adiunge te ad currum istum
ACTS|8|30|adcurrens autem Philippus audivit illum legentem Esaiam prophetam et dixit putasne intellegis quae legis
ACTS|8|31|qui ait et quomodo possum si non aliquis ostenderit mihi rogavitque Philippum ut ascenderet et sederet secum
ACTS|8|32|locus autem scripturae quam legebat erat hic tamquam ovis ad occisionem ductus est et sicut agnus coram tondente se sine voce sic non aperuit os suum
ACTS|8|33|in humilitate iudicium eius sublatum est generationem illius quis enarrabit quoniam tollitur de terra vita eius
ACTS|8|34|respondens autem eunuchus Philippo dixit obsecro te de quo propheta dicit hoc de se an de alio aliquo
ACTS|8|35|aperiens autem Philippus os suum et incipiens ab scriptura ista evangelizavit illi Iesum
ACTS|8|36|et dum irent per viam venerunt ad quandam aquam et ait eunuchus ecce aqua quid prohibet me baptizari
ACTS|8|37|
ACTS|8|38|et iussit stare currum et descenderunt uterque in aquam Philippus et eunuchus et baptizavit eum
ACTS|8|39|cum autem ascendissent de aqua Spiritus Domini rapuit Philippum et amplius non vidit eum eunuchus ibat enim per viam suam gaudens
ACTS|8|40|Philippus autem inventus est in Azoto et pertransiens evangelizabat civitatibus cunctis donec veniret Caesaream
ACTS|9|1|Saulus autem adhuc inspirans minarum et caedis in discipulos Domini accessit ad principem sacerdotum
ACTS|9|2|et petiit ab eo epistulas in Damascum ad synagogas ut si quos invenisset huius viae viros ac mulieres vinctos perduceret in Hierusalem
ACTS|9|3|et cum iter faceret contigit ut adpropinquaret Damasco et subito circumfulsit eum lux de caelo
ACTS|9|4|et cadens in terram audivit vocem dicentem sibi Saule Saule quid me persequeris
ACTS|9|5|qui dixit quis es Domine et ille ego sum Iesus quem tu persequeris
ACTS|9|6|
ACTS|9|7|sed surge et ingredere civitatem et dicetur tibi quid te oporteat facere viri autem illi qui comitabantur cum eo stabant stupefacti audientes quidem vocem neminem autem videntes
ACTS|9|8|surrexit autem Saulus de terra apertisque oculis nihil videbat ad manus autem illum trahentes introduxerunt Damascum
ACTS|9|9|et erat tribus diebus non videns et non manducavit neque bibit
ACTS|9|10|erat autem quidam discipulus Damasci nomine Ananias et dixit ad illum in visu Dominus Anania at ille ait ecce ego Domine
ACTS|9|11|et Dominus ad illum surgens vade in vicum qui vocatur Rectus et quaere in domo Iudae Saulum nomine Tarsensem ecce enim orat
ACTS|9|12|et vidit virum Ananiam nomine introeuntem et inponentem sibi manus ut visum recipiat
ACTS|9|13|respondit autem Ananias Domine audivi a multis de viro hoc quanta mala sanctis tuis fecerit in Hierusalem
ACTS|9|14|et hic habet potestatem a principibus sacerdotum alligandi omnes qui invocant nomen tuum
ACTS|9|15|dixit autem ad eum Dominus vade quoniam vas electionis est mihi iste ut portet nomen meum coram gentibus et regibus et filiis Israhel
ACTS|9|16|ego enim ostendam illi quanta oporteat eum pro nomine meo pati
ACTS|9|17|et abiit Ananias et introivit in domum et inponens ei manus dixit Saule frater Dominus misit me Iesus qui apparuit tibi in via qua veniebas ut videas et implearis Spiritu Sancto
ACTS|9|18|et confestim ceciderunt ab oculis eius tamquam squamae et visum recepit et surgens baptizatus est
ACTS|9|19|et cum accepisset cibum confortatus est fuit autem cum discipulis qui erant Damasci per dies aliquot
ACTS|9|20|et continuo in synagogis praedicabat Iesum quoniam hic est Filius Dei
ACTS|9|21|stupebant autem omnes qui audiebant et dicebant nonne hic est qui expugnabat in Hierusalem eos qui invocabant nomen istud et huc ad hoc venit ut vinctos illos duceret ad principes sacerdotum
ACTS|9|22|Saulus autem magis convalescebat et confundebat Iudaeos qui habitabant Damasci adfirmans quoniam hic est Christus
ACTS|9|23|cum implerentur autem dies multi consilium fecerunt Iudaei ut eum interficerent
ACTS|9|24|notae autem factae sunt Saulo insidiae eorum custodiebant autem et portas die ac nocte ut eum interficerent
ACTS|9|25|accipientes autem discipuli eius nocte per murum dimiserunt eum submittentes in sporta
ACTS|9|26|cum autem venisset in Hierusalem temptabat iungere se discipulis et omnes timebant eum non credentes quia esset discipulus
ACTS|9|27|Barnabas autem adprehensum illum duxit ad apostolos et narravit illis quomodo in via vidisset Dominum et quia locutus est ei et quomodo in Damasco fiducialiter egerit in nomine Iesu
ACTS|9|28|et erat cum illis intrans et exiens in Hierusalem et fiducialiter agens in nomine Domini
ACTS|9|29|loquebatur quoque et disputabat cum Graecis illi autem quaerebant occidere eum
ACTS|9|30|quod cum cognovissent fratres deduxerunt eum Caesaream et dimiserunt Tarsum
ACTS|9|31|ecclesia quidem per totam Iudaeam et Galilaeam et Samariam habebat pacem et aedificabatur ambulans in timore Domini et consolatione Sancti Spiritus replebatur
ACTS|9|32|factum est autem Petrum dum pertransiret universos devenire et ad sanctos qui habitabant Lyddae
ACTS|9|33|invenit autem ibi hominem quendam nomine Aeneam ab annis octo iacentem in grabatto qui erat paralyticus
ACTS|9|34|et ait illi Petrus Aeneas sanat te Iesus Christus surge et sterne tibi et continuo surrexit
ACTS|9|35|et viderunt illum omnes qui habitabant Lyddae et Saronae qui conversi sunt ad Dominum
ACTS|9|36|in Ioppe autem fuit quaedam discipula nomine Tabitas quae interpretata dicitur Dorcas haec erat plena operibus bonis et elemosynis quas faciebat
ACTS|9|37|factum est autem in diebus illis ut infirmata moreretur quam cum lavissent posuerunt eam in cenaculo
ACTS|9|38|cum autem prope esset Lydda ab Ioppe discipuli audientes quia Petrus esset in ea miserunt duos viros ad eum rogantes ne pigriteris venire usque ad nos
ACTS|9|39|exsurgens autem Petrus venit cum illis et cum advenisset duxerunt illum in cenaculum et circumsteterunt illum omnes viduae flentes et ostendentes tunicas et vestes quas faciebat illis Dorcas
ACTS|9|40|eiectis autem omnibus foras Petrus ponens genua oravit et conversus ad corpus dixit Tabita surge at illa aperuit oculos suos et viso Petro resedit
ACTS|9|41|dans autem illi manum erexit eam et cum vocasset sanctos et viduas adsignavit eam vivam
ACTS|9|42|notum autem factum est per universam Ioppen et crediderunt multi in Domino
ACTS|9|43|factum est autem ut dies multos moraretur in Ioppe apud quendam Simonem coriarium
ACTS|10|1|vir autem quidam erat in Caesarea nomine Cornelius centurio cohortis quae dicitur Italica
ACTS|10|2|religiosus et timens Deum cum omni domo sua faciens elemosynas multas plebi et deprecans Deum semper
ACTS|10|3|vidit in visu manifeste quasi hora nona diei angelum Dei introeuntem ad se et dicentem sibi Corneli
ACTS|10|4|at ille intuens eum timore correptus dixit quid est domine dixit autem illi orationes tuae et elemosynae tuae ascenderunt in memoriam in conspectu Dei
ACTS|10|5|et nunc mitte viros in Ioppen et accersi Simonem quendam qui cognominatur Petrus
ACTS|10|6|hic hospitatur apud Simonem quendam coriarium cuius est domus iuxta mare
ACTS|10|7|et cum discessisset angelus qui loquebatur illi vocavit duos domesticos suos et militem metuentem Dominum ex his qui illi parebant
ACTS|10|8|quibus cum narrasset omnia misit illos in Ioppen
ACTS|10|9|postera autem die iter illis facientibus et adpropinquantibus civitati ascendit Petrus in superiora ut oraret circa horam sextam
ACTS|10|10|et cum esuriret voluit gustare parantibus autem eis cecidit super eum mentis excessus
ACTS|10|11|et videt caelum apertum et descendens vas quoddam velut linteum magnum quattuor initiis submitti de caelo in terram
ACTS|10|12|in quo erant omnia quadrupedia et serpentia terrae et volatilia caeli
ACTS|10|13|et facta est vox ad eum surge Petre et occide et manduca
ACTS|10|14|ait autem Petrus absit Domine quia numquam manducavi omne commune et inmundum
ACTS|10|15|et vox iterum secundo ad eum quae Deus purificavit ne tu commune dixeris
ACTS|10|16|hoc autem factum est per ter et statim receptum est vas in caelum
ACTS|10|17|et dum intra se haesitaret Petrus quidnam esset visio quam vidisset ecce viri qui missi erant a Cornelio inquirentes domum Simonis adstiterunt ad ianuam
ACTS|10|18|et cum vocassent interrogabant si Simon qui cognominatur Petrus illic haberet hospitium
ACTS|10|19|Petro autem cogitante de visione dixit Spiritus ei ecce viri tres quaerunt te
ACTS|10|20|surge itaque et descende et vade cum eis nihil dubitans quia ego misi illos
ACTS|10|21|descendens autem Petrus ad viros dixit ecce ego sum quem quaeritis quae causa est propter quam venistis
ACTS|10|22|qui dixerunt Cornelius centurio vir iustus et timens Deum et testimonium habens ab universa gente Iudaeorum responsum accepit ab angelo sancto accersire te in domum suam et audire verba abs te
ACTS|10|23|introducens igitur eos recepit hospitio sequenti autem die surgens profectus est cum eis et quidam ex fratribus ab Ioppe comitati sunt eum
ACTS|10|24|altera autem die introivit Caesaream Cornelius vero expectabat illos convocatis cognatis suis et necessariis amicis
ACTS|10|25|et factum est cum introisset Petrus obvius ei Cornelius et procidens ad pedes adoravit
ACTS|10|26|Petrus vero levavit eum dicens surge et ego ipse homo sum
ACTS|10|27|et loquens cum illo intravit et invenit multos qui convenerant
ACTS|10|28|dixitque ad illos vos scitis quomodo abominatum sit viro iudaeo coniungi aut accedere ad alienigenam et mihi ostendit Deus neminem communem aut inmundum dicere hominem
ACTS|10|29|propter quod sine dubitatione veni accersitus interrogo ergo quam ob causam accersistis me
ACTS|10|30|et Cornelius ait a nudius quartana die usque in hanc horam orans eram hora nona in domo mea et ecce vir stetit ante me in veste candida et ait
ACTS|10|31|Corneli exaudita est oratio tua et elemosynae tuae commemoratae sunt in conspectu Dei
ACTS|10|32|mitte ergo in Ioppen et accersi Simonem qui cognominatur Petrus hic hospitatur in domo Simonis coriarii iuxta mare
ACTS|10|33|confestim igitur misi ad te et tu bene fecisti veniendo nunc ergo omnes nos in conspectu tuo adsumus audire omnia quaecumque tibi praecepta sunt a Domino
ACTS|10|34|aperiens autem Petrus os dixit in veritate conperi quoniam non est personarum acceptor Deus
ACTS|10|35|sed in omni gente qui timet eum et operatur iustitiam acceptus est illi
ACTS|10|36|verbum misit filiis Israhel adnuntians pacem per Iesum Christum hic est omnium Dominus
ACTS|10|37|vos scitis quod factum est verbum per universam Iudaeam incipiens enim a Galilaea post baptismum quod praedicavit Iohannes
ACTS|10|38|Iesum a Nazareth quomodo unxit eum Deus Spiritu Sancto et virtute qui pertransivit benefaciendo et sanando omnes oppressos a diabolo quoniam Deus erat cum illo
ACTS|10|39|et nos testes sumus omnium quae fecit in regione Iudaeorum et Hierusalem quem et occiderunt suspendentes in ligno
ACTS|10|40|hunc Deus suscitavit tertia die et dedit eum manifestum fieri
ACTS|10|41|non omni populo sed testibus praeordinatis a Deo nobis qui manducavimus et bibimus cum illo postquam resurrexit a mortuis
ACTS|10|42|et praecepit nobis praedicare populo et testificari quia ipse est qui constitutus est a Deo iudex vivorum et mortuorum
ACTS|10|43|huic omnes prophetae testimonium perhibent remissionem peccatorum accipere per nomen eius omnes qui credunt in eum
ACTS|10|44|adhuc loquente Petro verba haec cecidit Spiritus Sanctus super omnes qui audiebant verbum
ACTS|10|45|et obstipuerunt ex circumcisione fideles qui venerant cum Petro quia et in nationes gratia Spiritus Sancti effusa est
ACTS|10|46|audiebant enim illos loquentes linguis et magnificantes Deum
ACTS|10|47|tunc respondit Petrus numquid aquam quis prohibere potest ut non baptizentur hii qui Spiritum Sanctum acceperunt sicut et nos
ACTS|10|48|et iussit eos in nomine Iesu Christi baptizari tunc rogaverunt eum ut maneret aliquot diebus
ACTS|11|1|audierunt autem apostoli et fratres qui erant in Iudaea quoniam et gentes receperunt verbum Dei
ACTS|11|2|cum ascendisset autem Petrus in Hierosolymam disceptabant adversus illum qui erant ex circumcisione
ACTS|11|3|dicentes quare introisti ad viros praeputium habentes et manducasti cum illis
ACTS|11|4|incipiens autem Petrus exponebat illis ordinem dicens
ACTS|11|5|ego eram in civitate Ioppe orans et vidi in excessu mentis visionem descendens vas quoddam velut linteum magnum quattuor initiis submitti de caelo et venit usque ad me
ACTS|11|6|in quod intuens considerabam et vidi quadrupedia terrae et bestias et reptilia et volatilia caeli
ACTS|11|7|audivi autem et vocem dicentem mihi surgens Petre occide et manduca
ACTS|11|8|dixi autem nequaquam Domine quia commune aut inmundum numquam introivit in os meum
ACTS|11|9|respondit autem vox secundo de caelo quae Deus mundavit tu ne commune dixeris
ACTS|11|10|hoc autem factum est per ter et recepta sunt rursum omnia in caelum
ACTS|11|11|et ecce confestim tres viri adstiterunt in domo in qua eram missi a Caesarea ad me
ACTS|11|12|dixit autem Spiritus mihi ut irem cum illis nihil haesitans venerunt autem mecum et sex fratres isti et ingressi sumus in domum viri
ACTS|11|13|narravit autem nobis quomodo vidisset angelum in domo sua stantem et dicentem sibi mitte in Ioppen et accersi Simonem qui cognominatur Petrus
ACTS|11|14|qui loquetur tibi verba in quibus salvus eris tu et universa domus tua
ACTS|11|15|cum autem coepissem loqui decidit Spiritus Sanctus super eos sicut et in nos in initio
ACTS|11|16|recordatus sum autem verbi Domini sicut dicebat Iohannes quidem baptizavit aqua vos autem baptizabimini Spiritu Sancto
ACTS|11|17|si ergo eandem gratiam dedit illis Deus sicut et nobis qui credidimus in Dominum Iesum Christum ego quis eram qui possem prohibere Deum
ACTS|11|18|his auditis tacuerunt et glorificaverunt Deum dicentes ergo et gentibus Deus paenitentiam ad vitam dedit
ACTS|11|19|et illi quidem qui dispersi fuerant a tribulatione quae facta fuerat sub Stephano perambulaverunt usque Foenicen et Cyprum et Antiochiam nemini loquentes verbum nisi solis Iudaeis
ACTS|11|20|erant autem quidam ex eis viri cyprii et cyrenei qui cum introissent Antiochiam loquebantur et ad Graecos adnuntiantes Dominum Iesum
ACTS|11|21|et erat manus Domini cum eis multusque numerus credentium conversus est ad Dominum
ACTS|11|22|pervenit autem sermo ad aures ecclesiae quae erat Hierosolymis super istis et miserunt Barnaban usque Antiochiam
ACTS|11|23|qui cum pervenisset et vidisset gratiam Dei gavisus est et hortabatur omnes proposito cordis permanere in Domino
ACTS|11|24|quia erat vir bonus et plenus Spiritu Sancto et fide et adposita est turba multa Domino
ACTS|11|25|profectus est autem Tarsum ut quaereret Saulum quem cum invenisset perduxit Antiochiam
ACTS|11|26|et annum totum conversati sunt in ecclesia et docuerunt turbam multam ita ut cognominarentur primum Antiochiae discipuli Christiani
ACTS|11|27|in his autem diebus supervenerunt ab Hierosolymis prophetae Antiochiam
ACTS|11|28|et surgens unus ex eis nomine Agabus significabat per Spiritum famem magnam futuram in universo orbe terrarum quae facta est sub Claudio
ACTS|11|29|discipuli autem prout quis habebat proposuerunt singuli eorum in ministerium mittere habitantibus in Iudaea fratribus
ACTS|11|30|quod et fecerunt mittentes ad seniores per manus Barnabae et Sauli
ACTS|12|1|eodem autem tempore misit Herodes rex manus ut adfligeret quosdam de ecclesia
ACTS|12|2|occidit autem Iacobum fratrem Iohannis gladio
ACTS|12|3|videns autem quia placeret Iudaeis adposuit adprehendere et Petrum erant autem dies azymorum
ACTS|12|4|quem cum adprehendisset misit in carcerem tradens quattuor quaternionibus militum custodire eum volens post pascha producere eum populo
ACTS|12|5|et Petrus quidem servabatur in carcere oratio autem fiebat sine intermissione ab ecclesia ad Deum pro eo
ACTS|12|6|cum autem producturus eum esset Herodes in ipsa nocte erat Petrus dormiens inter duos milites vinctus catenis duabus et custodes ante ostium custodiebant carcerem
ACTS|12|7|et ecce angelus Domini adstitit et lumen refulsit in habitaculo percussoque latere Petri suscitavit eum dicens surge velociter et ceciderunt catenae de manibus eius
ACTS|12|8|dixit autem angelus ad eum praecingere et calcia te gallicas tuas et fecit sic et dixit illi circumda tibi vestimentum tuum et sequere me
ACTS|12|9|et exiens sequebatur et nesciebat quia verum est quod fiebat per angelum aestimabat autem se visum videre
ACTS|12|10|transeuntes autem primam et secundam custodiam venerunt ad portam ferream quae ducit ad civitatem quae ultro aperta est eis et exeuntes processerunt vicum unum et continuo discessit angelus ab eo
ACTS|12|11|et Petrus ad se reversus dixit nunc scio vere quia misit Dominus angelum suum et eripuit me de manu Herodis et de omni expectatione plebis Iudaeorum
ACTS|12|12|consideransque venit ad domum Mariae matris Iohannis qui cognominatus est Marcus ubi erant multi congregati et orantes
ACTS|12|13|pulsante autem eo ostium ianuae processit puella ad audiendum nomine Rhode
ACTS|12|14|et ut cognovit vocem Petri prae gaudio non aperuit ianuam sed intro currens nuntiavit stare Petrum ante ianuam
ACTS|12|15|at illi dixerunt ad eam insanis illa autem adfirmabat sic se habere illi autem dicebant angelus eius est
ACTS|12|16|Petrus autem perseverabat pulsans cum autem aperuissent viderunt eum et obstipuerunt
ACTS|12|17|annuens autem eis manu ut tacerent enarravit quomodo Dominus eduxisset eum de carcere dixitque nuntiate Iacobo et fratribus haec et egressus abiit in alium locum
ACTS|12|18|facta autem die erat non parva turbatio inter milites quidnam de Petro factum esset
ACTS|12|19|Herodes autem cum requisisset eum et non invenisset inquisitione facta de custodibus iussit eos duci descendensque a Iudaea in Caesaream ibi commoratus est
ACTS|12|20|erat autem iratus Tyriis et Sidoniis at illi unianimes venerunt ad eum et persuaso Blasto qui erat super cubiculum regis postulabant pacem eo quod alerentur regiones eorum ab illo
ACTS|12|21|statuto autem die Herodes vestitus veste regia sedit pro tribunali et contionabatur ad eos
ACTS|12|22|populus autem adclamabat dei voces et non hominis
ACTS|12|23|confestim autem percussit eum angelus Domini eo quod non dedisset honorem Deo et consumptus a vermibus exspiravit
ACTS|12|24|verbum autem Domini crescebat et multiplicabatur
ACTS|12|25|Barnabas autem et Saulus reversi sunt ab Hierosolymis expleto ministerio adsumpto Iohanne qui cognominatus est Marcus
ACTS|13|1|erant autem in ecclesia quae erat Antiochiae prophetae et doctores in quibus Barnabas et Symeon qui vocabatur Niger et Lucius Cyrenensis et Manaen qui erat Herodis tetrarchae conlactaneus et Saulus
ACTS|13|2|ministrantibus autem illis Domino et ieiunantibus dixit Spiritus Sanctus separate mihi Barnaban et Saulum in opus quod adsumpsi eos
ACTS|13|3|tunc ieiunantes et orantes inponentesque eis manus dimiserunt illos
ACTS|13|4|et ipsi quidem missi ab Spiritu Sancto abierunt Seleuciam et inde navigaverunt Cyprum
ACTS|13|5|et cum venissent Salamina praedicabant verbum Dei in synagogis Iudaeorum habebant autem et Iohannem in ministerio
ACTS|13|6|et cum perambulassent universam insulam usque Paphum invenerunt quendam virum magum pseudoprophetam Iudaeum cui nomen erat Bariesu
ACTS|13|7|qui erat cum proconsule Sergio Paulo viro prudente hic accitis Barnaba et Saulo desiderabat audire verbum Dei
ACTS|13|8|resistebat autem illis Elymas magus sic enim interpretatur nomen eius quaerens avertere proconsulem a fide
ACTS|13|9|Saulus autem qui et Paulus repletus Spiritu Sancto intuens in eum
ACTS|13|10|dixit o plene omni dolo et omni fallacia fili diaboli inimice omnis iustitiae non desinis subvertere vias Domini rectas
ACTS|13|11|et nunc ecce manus Domini super te et eris caecus non videns solem usque ad tempus et confestim cecidit in eum caligo et tenebrae et circumiens quaerebat qui ei manum daret
ACTS|13|12|tunc proconsul cum vidisset factum credidit admirans super doctrinam Domini
ACTS|13|13|et cum a Papho navigassent Paulus et qui cum eo venerunt Pergen Pamphiliae Iohannes autem discedens ab eis reversus est Hierosolymam
ACTS|13|14|illi vero pertranseuntes Pergen venerunt Antiochiam Pisidiae et ingressi synagogam die sabbatorum sederunt
ACTS|13|15|post lectionem autem legis et prophetarum miserunt principes synagogae ad eos dicentes viri fratres si quis est in vobis sermo exhortationis ad plebem dicite
ACTS|13|16|surgens autem Paulus et manu silentium indicens ait viri israhelitae et qui timetis Deum audite
ACTS|13|17|Deus plebis Israhel elegit patres nostros et plebem exaltavit cum essent incolae in terra Aegypti et in brachio excelso eduxit eos ex ea
ACTS|13|18|et per quadraginta annorum tempus mores eorum sustinuit in deserto
ACTS|13|19|et destruens gentes septem in terra Chanaan sorte distribuit eis terram eorum
ACTS|13|20|quasi post quadringentos et quinquaginta annos et post haec dedit iudices usque ad Samuhel prophetam
ACTS|13|21|et exinde postulaverunt regem et dedit illis Deus Saul filium Cis virum de tribu Beniamin annis quadraginta
ACTS|13|22|et amoto illo suscitavit illis David regem cui et testimonium perhibens dixit inveni David filium Iesse virum secundum cor meum qui faciet omnes voluntates meas
ACTS|13|23|huius Deus ex semine secundum promissionem eduxit Israhel salvatorem Iesum
ACTS|13|24|praedicante Iohanne ante faciem adventus eius baptismum paenitentiae omni populo Israhel
ACTS|13|25|cum impleret autem Iohannes cursum suum dicebat quem me arbitramini esse non sum ego sed ecce venit post me cuius non sum dignus calciamenta pedum solvere
ACTS|13|26|viri fratres filii generis Abraham et qui in vobis timent Deum vobis verbum salutis huius missum est
ACTS|13|27|qui enim habitabant Hierusalem et principes eius hunc ignorantes et voces prophetarum quae per omne sabbatum leguntur iudicantes impleverunt
ACTS|13|28|et nullam causam mortis invenientes in eum petierunt a Pilato ut interficerent eum
ACTS|13|29|cumque consummassent omnia quae de eo scripta erant deponentes eum de ligno posuerunt in monumento
ACTS|13|30|Deus vero suscitavit eum a mortuis qui visus est per dies multos his
ACTS|13|31|qui simul ascenderant cum eo de Galilaea in Hierusalem qui usque nunc sunt testes eius ad plebem
ACTS|13|32|et nos vobis adnuntiamus ea quae ad patres nostros repromissio facta est
ACTS|13|33|quoniam hanc Deus adimplevit filiis nostris resuscitans Iesum sicut et in psalmo secundo scriptum est Filius meus es tu ego hodie genui te
ACTS|13|34|quod autem suscitaverit eum a mortuis amplius iam non reversurum in corruptionem ita dixit quia dabo vobis sancta David fidelia
ACTS|13|35|ideoque et alias dicit non dabis Sanctum tuum videre corruptionem
ACTS|13|36|David enim sua generatione cum administrasset voluntati Dei dormivit et adpositus est ad patres suos et vidit corruptionem
ACTS|13|37|quem vero Deus suscitavit non vidit corruptionem
ACTS|13|38|notum igitur sit vobis viri fratres quia per hunc vobis remissio peccatorum adnuntiatur ab omnibus quibus non potuistis in lege Mosi iustificari
ACTS|13|39|in hoc omnis qui credit iustificatur
ACTS|13|40|videte ergo ne superveniat quod dictum est in prophetis
ACTS|13|41|videte contemptores et admiramini et disperdimini quia opus operor ego in diebus vestris opus quod non credetis si quis enarraverit vobis
ACTS|13|42|exeuntibus autem illis rogabant ut sequenti sabbato loquerentur sibi verba haec
ACTS|13|43|cumque dimissa esset synagoga secuti sunt multi Iudaeorum et colentium advenarum Paulum et Barnaban qui loquentes suadebant eis ut permanerent in gratia Dei
ACTS|13|44|sequenti vero sabbato paene universa civitas convenit audire verbum Domini
ACTS|13|45|videntes autem turbas Iudaei repleti sunt zelo et contradicebant his quae a Paulo dicebantur blasphemantes
ACTS|13|46|tunc constanter Paulus et Barnabas dixerunt vobis oportebat primum loqui verbum Dei sed quoniam repellitis illud et indignos vos iudicastis aeternae vitae ecce convertimur ad gentes
ACTS|13|47|sic enim praecepit nobis Dominus posui te in lumen gentibus ut sis in salutem usque ad extremum terrae
ACTS|13|48|audientes autem gentes gavisae sunt et glorificabant verbum Domini et crediderunt quotquot erant praeordinati ad vitam aeternam
ACTS|13|49|disseminabatur autem verbum Domini per universam regionem
ACTS|13|50|Iudaei autem concitaverunt religiosas mulieres et honestas et primos civitatis et excitaverunt persecutionem in Paulum et Barnaban et eiecerunt eos de finibus suis
ACTS|13|51|at illi excusso pulvere pedum in eos venerunt Iconium
ACTS|13|52|discipuli quoque replebantur gaudio et Spiritu Sancto
ACTS|14|1|factum est autem Iconii ut simul introirent synagogam Iudaeorum et loquerentur ita ut crederet Iudaeorum et Graecorum copiosa multitudo
ACTS|14|2|qui vero increduli fuerunt Iudaei suscitaverunt et ad iracundiam concitaverunt animas gentium adversus fratres
ACTS|14|3|multo igitur tempore demorati sunt fiducialiter agentes in Domino testimonium perhibente verbo gratiae suae dante signa et prodigia fieri per manus eorum
ACTS|14|4|divisa est autem multitudo civitatis et quidam quidem erant cum Iudaeis quidam vero cum apostolis
ACTS|14|5|cum autem factus esset impetus gentilium et Iudaeorum cum principibus suis ut contumeliis adficerent et lapidarent eos
ACTS|14|6|intellegentes confugerunt ad civitates Lycaoniae Lystram et Derben et universam in circuitu regionem et ibi evangelizantes erant
ACTS|14|7|et quidam vir in Lystris infirmus pedibus sedebat claudus ex utero matris suae qui numquam ambulaverat
ACTS|14|8|hic audivit Paulum loquentem qui intuitus eum et videns quia haberet fidem ut salvus fieret
ACTS|14|9|dixit magna voce surge super pedes tuos rectus et exilivit et ambulabat
ACTS|14|10|turbae autem cum vidissent quod fecerat Paulus levaverunt vocem suam lycaonice dicentes dii similes facti hominibus descenderunt ad nos
ACTS|14|11|et vocabant Barnaban Iovem Paulum vero Mercurium quoniam ipse erat dux verbi
ACTS|14|12|sacerdos quoque Iovis qui erat ante civitatem tauros et coronas ante ianuas adferens cum populis volebat sacrificare
ACTS|14|13|quod ubi audierunt apostoli Barnabas et Paulus conscissis tunicis suis exilierunt in turbas clamantes
ACTS|14|14|et dicentes viri quid haec facitis et nos mortales sumus similes vobis homines adnuntiantes vobis ab his vanis converti ad Deum vivum qui fecit caelum et terram et mare et omnia quae in eis sunt
ACTS|14|15|qui in praeteritis generationibus dimisit omnes gentes ingredi in vias suas
ACTS|14|16|et quidem non sine testimonio semet ipsum reliquit benefaciens de caelo dans pluvias et tempora fructifera implens cibo et laetitia corda vestra
ACTS|14|17|et haec dicentes vix sedaverunt turbas ne sibi immolarent
ACTS|14|18|supervenerunt autem quidam ab Antiochia et Iconio Iudaei et persuasis turbis lapidantesque Paulum traxerunt extra civitatem aestimantes eum mortuum esse
ACTS|14|19|circumdantibus autem eum discipulis surgens intravit civitatem et postera die profectus est cum Barnaba in Derben
ACTS|14|20|cumque evangelizassent civitati illi et docuissent multos reversi sunt Lystram et Iconium et Antiochiam
ACTS|14|21|confirmantes animas discipulorum exhortantes ut permanerent in fide et quoniam per multas tribulationes oportet nos intrare in regnum Dei
ACTS|14|22|et cum constituissent illis per singulas ecclesias presbyteros et orassent cum ieiunationibus commendaverunt eos Domino in quem crediderunt
ACTS|14|23|transeuntesque Pisidiam venerunt Pamphiliam
ACTS|14|24|et loquentes in Pergen verbum Domini descenderunt in Attaliam
ACTS|14|25|et inde navigaverunt Antiochiam unde erant traditi gratiae Dei in opus quod conpleverunt
ACTS|14|26|cum autem venissent et congregassent ecclesiam rettulerunt quanta fecisset Deus cum illis quia aperuisset gentibus ostium fidei
ACTS|14|27|morati sunt autem tempus non modicum cum discipulis
ACTS|15|1|et quidam descendentes de Iudaea docebant fratres quia nisi circumcidamini secundum morem Mosi non potestis salvi fieri
ACTS|15|2|facta ergo seditione non minima Paulo et Barnabae adversum illos statuerunt ut ascenderent Paulus et Barnabas et quidam alii ex illis ad apostolos et presbyteros in Hierusalem super hac quaestione
ACTS|15|3|illi igitur deducti ab ecclesia pertransiebant Foenicen et Samariam narrantes conversionem gentium et faciebant gaudium magnum omnibus fratribus
ACTS|15|4|cum autem venissent Hierosolymam suscepti sunt ab ecclesia et ab apostolis et senioribus adnuntiantes quanta Deus fecisset cum illis
ACTS|15|5|surrexerunt autem quidam de heresi Pharisaeorum qui crediderant dicentes quia oportet circumcidi eos praecipere quoque servare legem Mosi
ACTS|15|6|conveneruntque apostoli et seniores videre de verbo hoc
ACTS|15|7|cum autem magna conquisitio fieret surgens Petrus dixit ad eos viri fratres vos scitis quoniam ab antiquis diebus in nobis elegit Deus per os meum audire gentes verbum evangelii et credere
ACTS|15|8|et qui novit corda Deus testimonium perhibuit dans illis Spiritum Sanctum sicut et nobis
ACTS|15|9|et nihil discrevit inter nos et illos fide purificans corda eorum
ACTS|15|10|nunc ergo quid temptatis Deum inponere iugum super cervicem discipulorum quod neque patres nostri neque nos portare potuimus
ACTS|15|11|sed per gratiam Domini Iesu credimus salvari quemadmodum et illi
ACTS|15|12|tacuit autem omnis multitudo et audiebant Barnaban et Paulum narrantes quanta fecisset Deus signa et prodigia in gentibus per eos
ACTS|15|13|et postquam tacuerunt respondit Iacobus dicens viri fratres audite me
ACTS|15|14|Simeon narravit quemadmodum primum Deus visitavit sumere ex gentibus populum nomini suo
ACTS|15|15|et huic concordant verba prophetarum sicut scriptum est
ACTS|15|16|post haec revertar et aedificabo tabernaculum David quod decidit et diruta eius reaedificabo et erigam illud
ACTS|15|17|ut requirant ceteri hominum Dominum et omnes gentes super quas invocatum est nomen meum dicit Dominus faciens haec
ACTS|15|18|notum a saeculo est Domino opus suum
ACTS|15|19|propter quod ego iudico non inquietari eos qui ex gentibus convertuntur ad Deum
ACTS|15|20|sed scribere ad eos ut abstineant se a contaminationibus simulacrorum et fornicatione et suffocatis et sanguine
ACTS|15|21|Moses enim a temporibus antiquis habet in singulis civitatibus qui eum praedicent in synagogis ubi per omne sabbatum legitur
ACTS|15|22|tunc placuit apostolis et senioribus cum omni ecclesia eligere viros ex eis et mittere Antiochiam cum Paulo et Barnaba Iudam qui cognominatur Barsabban et Silam viros primos in fratribus
ACTS|15|23|scribentes per manus eorum apostoli et seniores fratres his qui sunt Antiochiae et Syriae et Ciliciae fratribus ex gentibus salutem
ACTS|15|24|quoniam audivimus quia quidam ex nobis exeuntes turbaverunt vos verbis evertentes animas vestras quibus non mandavimus
ACTS|15|25|placuit nobis collectis in unum eligere viros et mittere ad vos cum carissimis nostris Barnaba et Paulo
ACTS|15|26|hominibus qui tradiderunt animas suas pro nomine Domini nostri Iesu Christi
ACTS|15|27|misimus ergo Iudam et Silam qui et ipsi vobis verbis referent eadem
ACTS|15|28|visum est enim Spiritui Sancto et nobis nihil ultra inponere vobis oneris quam haec necessario
ACTS|15|29|ut abstineatis vos ab immolatis simulacrorum et sanguine suffocato et fornicatione a quibus custodientes vos bene agetis valete
ACTS|15|30|illi igitur dimissi descenderunt Antiochiam et congregata multitudine tradiderunt epistulam
ACTS|15|31|quam cum legissent gavisi sunt super consolatione
ACTS|15|32|Iudas autem et Silas et ipsi cum essent prophetae verbo plurimo consolati sunt fratres et confirmaverunt
ACTS|15|33|facto autem ibi tempore dimissi sunt cum pace a fratribus ad eos qui miserant illos
ACTS|15|34|
ACTS|15|35|Paulus autem et Barnabas demorabantur Antiochiae docentes et evangelizantes cum aliis pluribus verbum Domini
ACTS|15|36|post aliquot autem dies dixit ad Barnaban Paulus revertentes visitemus fratres per universas civitates in quibus praedicavimus verbum Domini quomodo se habeant
ACTS|15|37|Barnabas autem volebat secum adsumere et Iohannem qui cognominatur Marcus
ACTS|15|38|Paulus autem rogabat eum qui discessisset ab eis a Pamphilia et non isset cum eis in opus non debere recipi eum
ACTS|15|39|facta est autem dissensio ita ut discederent ab invicem et Barnabas adsumpto Marco navigaret Cyprum
ACTS|15|40|Paulus vero electo Sila profectus est traditus gratiae Domini a fratribus
ACTS|15|41|perambulabat autem Syriam et Ciliciam confirmans ecclesias
ACTS|16|1|pervenit autem in Derben et Lystram et ecce discipulus quidam erat ibi nomine Timotheus filius mulieris iudaeae fidelis patre gentili
ACTS|16|2|huic testimonium reddebant qui in Lystris erant et Iconii fratres
ACTS|16|3|hunc voluit Paulus secum proficisci et adsumens circumcidit eum propter Iudaeos qui erant in illis locis sciebant enim omnes quod pater eius gentilis esset
ACTS|16|4|cum autem pertransirent civitates tradebant eis custodire dogmata quae erant decreta ab apostolis et senioribus qui essent Hierosolymis
ACTS|16|5|et ecclesiae quidem confirmabantur fide et abundabant numero cotidie
ACTS|16|6|transeuntes autem Frygiam et Galatiae regionem vetati sunt a Sancto Spiritu loqui verbum in Asia
ACTS|16|7|cum venissent autem in Mysiam temptabant ire Bithyniam et non permisit eos Spiritus Iesu
ACTS|16|8|cum autem pertransissent Mysiam descenderunt Troadem
ACTS|16|9|et visio per noctem Paulo ostensa est vir macedo quidam erat stans et deprecans eum et dicens transiens in Macedoniam adiuva nos
ACTS|16|10|ut autem visum vidit statim quaesivimus proficisci in Macedoniam certi facti quia vocasset nos Deus evangelizare eis
ACTS|16|11|navigantes autem a Troade recto cursu venimus Samothraciam et sequenti die Neapolim
ACTS|16|12|et inde Philippis quae est prima partis Macedoniae civitas colonia eramus autem in hac urbe diebus aliquot conferentes
ACTS|16|13|die autem sabbatorum egressi sumus foras portam iuxta flumen ubi videbatur oratio esse et sedentes loquebamur mulieribus quae convenerant
ACTS|16|14|et quaedam mulier nomine Lydia purpuraria civitatis Thyatirenorum colens Deum audivit cuius Dominus aperuit cor intendere his quae dicebantur a Paulo
ACTS|16|15|cum autem baptizata esset et domus eius deprecata est dicens si iudicastis me fidelem Domino esse introite in domum meam et manete et coegit nos
ACTS|16|16|factum est autem euntibus nobis ad orationem puellam quandam habentem spiritum pythonem obviare nobis quae quaestum magnum praestabat dominis suis divinando
ACTS|16|17|haec subsecuta Paulum et nos clamabat dicens isti homines servi Dei excelsi sunt qui adnuntiant vobis viam salutis
ACTS|16|18|hoc autem faciebat multis diebus dolens autem Paulus et conversus spiritui dixit praecipio tibi in nomine Iesu Christi exire ab ea et exiit eadem hora
ACTS|16|19|videntes autem domini eius quia exivit spes quaestus eorum adprehendentes Paulum et Silam perduxerunt in forum ad principes
ACTS|16|20|et offerentes eos magistratibus dixerunt hii homines conturbant civitatem nostram cum sint Iudaei
ACTS|16|21|et adnuntiant morem quem non licet nobis suscipere neque facere cum simus Romani
ACTS|16|22|et concurrit plebs adversus eos et magistratus scissis tunicis eorum iusserunt virgis caedi
ACTS|16|23|et cum multas plagas eis inposuissent miserunt eos in carcerem praecipientes custodi ut diligenter custodiret eos
ACTS|16|24|qui cum tale praeceptum accepisset misit eos in interiorem carcerem et pedes eorum strinxit in ligno
ACTS|16|25|media autem nocte Paulus et Silas adorantes laudabant Deum et audiebant eos qui in custodia erant
ACTS|16|26|subito vero terraemotus factus est magnus ita ut moverentur fundamenta carceris et aperta sunt statim ostia omnia et universorum vincula soluta sunt
ACTS|16|27|expergefactus autem custos carceris et videns apertas ianuas carceris evaginato gladio volebat se interficere aestimans fugisse vinctos
ACTS|16|28|clamavit autem Paulus magna voce dicens nihil feceris tibi mali universi enim hic sumus
ACTS|16|29|petitoque lumine introgressus est et tremefactus procidit Paulo et Silae
ACTS|16|30|et producens eos foras ait domini quid me oportet facere ut salvus fiam
ACTS|16|31|at illi dixerunt crede in Domino Iesu et salvus eris tu et domus tua
ACTS|16|32|et locuti sunt ei verbum Domini cum omnibus qui erant in domo eius
ACTS|16|33|et tollens eos in illa hora noctis lavit plagas eorum et baptizatus est ipse et omnes eius continuo
ACTS|16|34|cumque perduxisset eos in domum suam adposuit eis mensam et laetatus est cum omni domo sua credens Deo
ACTS|16|35|et cum dies factus esset miserunt magistratus lictores dicentes dimitte homines illos
ACTS|16|36|nuntiavit autem custos carceris verba haec Paulo quia miserunt magistratus ut dimittamini nunc igitur exeuntes ite in pace
ACTS|16|37|Paulus autem dixit eis caesos nos publice indemnatos homines romanos miserunt in carcerem et nunc occulte nos eiciunt non ita sed veniant
ACTS|16|38|et ipsi nos eiciant nuntiaverunt autem magistratibus lictores verba haec timueruntque audito quod Romani essent
ACTS|16|39|et venientes deprecati sunt eos et educentes rogabant ut egrederentur urbem
ACTS|16|40|exeuntes autem de carcere introierunt ad Lydiam et visis fratribus consolati sunt eos et profecti sunt
ACTS|17|1|cum autem perambulassent Amphipolim et Apolloniam venerunt Thessalonicam ubi erat synagoga Iudaeorum
ACTS|17|2|secundum consuetudinem autem Paulus introivit ad eos et per sabbata tria disserebat eis de scripturis
ACTS|17|3|adaperiens et insinuans quia Christum oportuit pati et resurgere a mortuis et quia hic est Christus Iesus quem ego adnuntio vobis
ACTS|17|4|et quidam ex eis crediderunt et adiuncti sunt Paulo et Silae et de colentibus gentilibusque multitudo magna et mulieres nobiles non paucae
ACTS|17|5|zelantes autem Iudaei adsumentesque de vulgo viros quosdam malos et turba facta concitaverunt civitatem et adsistentes domui Iasonis quaerebant eos producere in populum
ACTS|17|6|et cum non invenissent eos trahebant Iasonem et quosdam fratres ad principes civitatis clamantes quoniam hii qui orbem concitant et huc venerunt
ACTS|17|7|quos suscepit Iason et hii omnes contra decreta Caesaris faciunt regem alium dicentes esse Iesum
ACTS|17|8|concitaverunt autem plebem et principes civitatis audientes haec
ACTS|17|9|et accepto satis ab Iasone et a ceteris dimiserunt eos
ACTS|17|10|fratres vero confestim per noctem dimiserunt Paulum et Silam in Beroeam qui cum advenissent in synagogam Iudaeorum introierunt
ACTS|17|11|hii autem erant nobiliores eorum qui sunt Thessalonicae qui susceperunt verbum cum omni aviditate cotidie scrutantes scripturas si haec ita se haberent
ACTS|17|12|et multi quidem crediderunt ex eis et gentilium mulierum honestarum et viri non pauci
ACTS|17|13|cum autem cognovissent in Thessalonica Iudaei quia et Beroeae praedicatum est a Paulo verbum Dei venerunt et illuc commoventes et turbantes multitudinem
ACTS|17|14|statimque tunc Paulum dimiserunt fratres ut iret usque ad mare Silas autem et Timotheus remanserunt ibi
ACTS|17|15|qui autem deducebant Paulum perduxerunt usque Athenas et accepto mandato ab eo ad Silam et Timotheum ut quam celeriter venirent ad illum profecti sunt
ACTS|17|16|Paulus autem cum Athenis eos expectaret incitabatur spiritus eius in ipso videns idolatriae deditam civitatem
ACTS|17|17|disputabat igitur in synagoga cum Iudaeis et colentibus et in foro per omnes dies ad eos qui aderant
ACTS|17|18|quidam autem epicurei et stoici philosophi disserebant cum eo et quidam dicebant quid vult seminiverbius hic dicere alii vero novorum daemoniorum videtur adnuntiator esse quia Iesum et resurrectionem adnuntiabat eis
ACTS|17|19|et adprehensum eum ad Ariopagum duxerunt dicentes possumus scire quae est haec nova quae a te dicitur doctrina
ACTS|17|20|nova enim quaedam infers auribus nostris volumus ergo scire quidnam velint haec esse
ACTS|17|21|Athenienses autem omnes et advenae hospites ad nihil aliud vacabant nisi aut dicere aut audire aliquid novi
ACTS|17|22|stans autem Paulus in medio Ariopagi ait viri athenienses per omnia quasi superstitiosiores vos video
ACTS|17|23|praeteriens enim et videns simulacra vestra inveni et aram in qua scriptum erat ignoto deo quod ergo ignorantes colitis hoc ego adnuntio vobis
ACTS|17|24|Deus qui fecit mundum et omnia quae in eo sunt hic caeli et terrae cum sit Dominus non in manufactis templis inhabitat
ACTS|17|25|nec manibus humanis colitur indigens aliquo cum ipse det omnibus vitam et inspirationem et omnia
ACTS|17|26|fecitque ex uno omne genus hominum inhabitare super universam faciem terrae definiens statuta tempora et terminos habitationis eorum
ACTS|17|27|quaerere Deum si forte adtractent eum aut inveniant quamvis non longe sit ab unoquoque nostrum
ACTS|17|28|in ipso enim vivimus et movemur et sumus sicut et quidam vestrum poetarum dixerunt ipsius enim et genus sumus
ACTS|17|29|genus ergo cum simus Dei non debemus aestimare auro aut argento aut lapidi sculpturae artis et cogitationis hominis divinum esse simile
ACTS|17|30|et tempora quidem huius ignorantiae despiciens Deus nunc adnuntiat hominibus ut omnes ubique paenitentiam agant
ACTS|17|31|eo quod statuit diem in qua iudicaturus est orbem in aequitate in viro in quo statuit fidem praebens omnibus suscitans eum a mortuis
ACTS|17|32|cum audissent autem resurrectionem mortuorum quidam quidem inridebant quidam vero dixerunt audiemus te de hoc iterum
ACTS|17|33|sic Paulus exivit de medio eorum
ACTS|17|34|quidam vero viri adherentes ei crediderunt in quibus et Dionisius Ariopagita et mulier nomine Damaris et alii cum eis
ACTS|18|1|post haec egressus ab Athenis venit Corinthum
ACTS|18|2|et inveniens quendam Iudaeum nomine Aquilam Ponticum genere qui nuper venerat ab Italia et Priscillam uxorem eius eo quod praecepisset Claudius discedere omnes Iudaeos a Roma accessit ad eos
ACTS|18|3|et quia eiusdem erat artis manebat apud eos et operabatur erat autem scenofactoriae artis
ACTS|18|4|
ACTS|18|5|cum venissent autem de Macedonia Silas et Timotheus instabat verbo Paulus testificans Iudaeis esse Christum Iesum
ACTS|18|6|contradicentibus autem eis et blasphemantibus excutiens vestimenta dixit ad eos sanguis vester super caput vestrum mundus ego ex hoc ad gentes vadam
ACTS|18|7|et migrans inde intravit in domum cuiusdam nomine Titi Iusti colentis Deum cuius domus erat coniuncta synagogae
ACTS|18|8|Crispus autem archisynagogus credidit Domino cum omni domo sua et multi Corinthiorum audientes credebant et baptizabantur
ACTS|18|9|dixit autem Dominus nocte per visionem Paulo noli timere sed loquere et ne taceas
ACTS|18|10|propter quod ego sum tecum et nemo adponetur tibi ut noceat te quoniam populus est mihi multus in hac civitate
ACTS|18|11|sedit autem annum et sex menses docens apud eos verbum Dei
ACTS|18|12|Gallione autem proconsule Achaiae insurrexerunt uno animo Iudaei in Paulum et adduxerunt eum ad tribunal
ACTS|18|13|dicentes quia contra legem hic persuadet hominibus colere Deum
ACTS|18|14|incipiente autem Paulo aperire os dixit Gallio ad Iudaeos si quidem esset iniquum aliquid aut facinus pessimum o viri iudaei recte vos sustinerem
ACTS|18|15|si vero quaestiones sunt de verbo et nominibus et legis vestrae vos ipsi videritis iudex ego horum nolo esse
ACTS|18|16|et minavit eos a tribunali
ACTS|18|17|adprehendentes autem omnes Sosthenen principem synagogae percutiebant ante tribunal et nihil eorum Gallioni curae erat
ACTS|18|18|Paulus vero cum adhuc sustinuisset dies multos fratribus valefaciens navigavit Syriam et cum eo Priscilla et Aquila qui sibi totonderat in Cencris caput habebat enim votum
ACTS|18|19|devenitque Ephesum et illos ibi reliquit ipse vero ingressus synagogam disputavit cum Iudaeis
ACTS|18|20|rogantibus autem eis ut ampliori tempore maneret non consensit
ACTS|18|21|sed valefaciens et dicens iterum revertar ad vos Deo volente profectus est ab Epheso
ACTS|18|22|et descendens Caesaream ascendit et salutavit ecclesiam et descendit Antiochiam
ACTS|18|23|et facto ibi aliquanto tempore profectus est perambulans ex ordine galaticam regionem et Frygiam confirmans omnes discipulos
ACTS|18|24|Iudaeus autem quidam Apollo nomine Alexandrinus natione vir eloquens devenit Ephesum potens in scripturis
ACTS|18|25|hic erat edoctus viam Domini et fervens spiritu loquebatur et docebat diligenter ea quae sunt Iesu sciens tantum baptisma Iohannis
ACTS|18|26|hic ergo coepit fiducialiter agere in synagoga quem cum audissent Priscilla et Aquila adsumpserunt eum et diligentius exposuerunt ei viam Dei
ACTS|18|27|cum autem vellet ire Achaiam exhortati fratres scripserunt discipulis ut susciperent eum qui cum venisset contulit multum his qui crediderant
ACTS|18|28|vehementer enim Iudaeos revincebat publice ostendens per scripturas esse Christum Iesum
ACTS|19|1|factum est autem cum Apollo esset Corinthi ut Paulus peragratis superioribus partibus veniret Ephesum et inveniret quosdam discipulos
ACTS|19|2|dixitque ad eos si Spiritum Sanctum accepistis credentes at illi ad eum sed neque si Spiritus Sanctus est audivimus
ACTS|19|3|ille vero ait in quo ergo baptizati estis qui dixerunt in Iohannis baptismate
ACTS|19|4|dixit autem Paulus Iohannes baptizavit baptisma paenitentiae populum dicens in eum qui venturus esset post ipsum ut crederent hoc est in Iesum
ACTS|19|5|his auditis baptizati sunt in nomine Domini Iesu
ACTS|19|6|et cum inposuisset illis manum Paulus venit Spiritus Sanctus super eos et loquebantur linguis et prophetabant
ACTS|19|7|erant autem omnes viri fere duodecim
ACTS|19|8|introgressus autem synagogam cum fiducia loquebatur per tres menses disputans et suadens de regno Dei
ACTS|19|9|cum autem quidam indurarentur et non crederent maledicentes viam coram multitudine discedens ab eis segregavit discipulos cotidie disputans in scola Tyranni
ACTS|19|10|hoc autem factum est per biennium ita ut omnes qui habitabant in Asia audirent verbum Domini Iudaei atque gentiles
ACTS|19|11|virtutesque non quaslibet Deus faciebat per manus Pauli
ACTS|19|12|ita ut etiam super languidos deferrentur a corpore eius sudaria vel semicintia et recedebant ab eis languores et spiritus nequam egrediebantur
ACTS|19|13|temptaverunt autem quidam et de circumeuntibus iudaeis exorcistis invocare super eos qui habebant spiritus malos nomen Domini Iesu dicentes adiuro vos per Iesum quem Paulus praedicat
ACTS|19|14|erant autem quidam Scevae Iudaei principis sacerdotum septem filii qui hoc faciebant
ACTS|19|15|respondens autem spiritus nequam dixit eis Iesum novi et Paulum scio vos autem qui estis
ACTS|19|16|et insiliens homo in eos in quo erat daemonium pessimum et dominatus amborum invaluit contra eos ita ut nudi et vulnerati effugerent de domo illa
ACTS|19|17|hoc autem notum factum est omnibus Iudaeis atque gentilibus qui habitabant Ephesi et cecidit timor super omnes illos et magnificabatur nomen Domini Iesu
ACTS|19|18|multique credentium veniebant confitentes et adnuntiantes actus suos
ACTS|19|19|multi autem ex his qui fuerant curiosa sectati contulerunt libros et conbuserunt coram omnibus et conputatis pretiis illorum invenerunt pecuniam denariorum quinquaginta milium
ACTS|19|20|ita fortiter verbum Dei crescebat et confirmabatur
ACTS|19|21|his autem expletis posuit Paulus in Spiritu transita Macedonia et Achaia ire Hierosolymam dicens quoniam postquam fuero ibi oportet me et Romam videre
ACTS|19|22|mittens autem in Macedoniam duos ex ministrantibus sibi Timotheum et Erastum ipse remansit ad tempus in Asia
ACTS|19|23|facta est autem in illo tempore turbatio non minima de via
ACTS|19|24|Demetrius enim quidam nomine argentarius faciens aedes argenteas Dianae praestabat artificibus non modicum quaestum
ACTS|19|25|quos convocans et eos qui eiusmodi erant opifices dixit viri scitis quia de hoc artificio adquisitio est nobis
ACTS|19|26|et videtis et auditis quia non solum Ephesi sed paene totius Asiae Paulus hic suadens avertit multam turbam dicens quoniam non sunt dii qui manibus fiunt
ACTS|19|27|non solum autem haec periclitabitur nobis pars in redargutionem venire sed et magnae deae Dianae templum in nihilum reputabitur sed et destrui incipiet maiestas eius quam tota Asia et orbis colit
ACTS|19|28|his auditis repleti sunt ira et exclamaverunt dicentes magna Diana Ephesiorum
ACTS|19|29|et impleta est civitas confusione et impetum fecerunt uno animo in theatrum rapto Gaio et Aristarcho Macedonibus comitibus Pauli
ACTS|19|30|Paulo autem volente intrare in populum non permiserunt discipuli
ACTS|19|31|quidam autem et de Asiae principibus qui erant amici eius miserunt ad eum rogantes ne se daret in theatrum
ACTS|19|32|alii autem aliud clamabant erat enim ecclesia confusa et plures nesciebant qua ex causa convenissent
ACTS|19|33|de turba autem detraxerunt Alexandrum propellentibus eum Iudaeis Alexander ergo manu silentio postulato volebat rationem reddere populo
ACTS|19|34|quem ut cognoverunt Iudaeum esse vox facta est una omnium quasi per horas duas clamantium magna Diana Ephesiorum
ACTS|19|35|et cum sedasset scriba turbas dixit viri ephesii quis enim est hominum qui nesciat Ephesiorum civitatem cultricem esse magnae Dianae Iovisque prolis
ACTS|19|36|cum ergo his contradici non possit oportet vos sedatos esse et nihil temere agere
ACTS|19|37|adduxistis enim homines istos neque sacrilegos neque blasphemantes deam vestram
ACTS|19|38|quod si Demetrius et qui cum eo sunt artifices habent adversus aliquem causam conventus forenses aguntur et pro consulibus sunt accusent invicem
ACTS|19|39|si quid autem alterius rei quaeritis in legitima ecclesia poterit absolvi
ACTS|19|40|nam et periclitamur argui seditionis hodiernae cum nullus obnoxius sit de quo non possimus reddere rationem concursus istius et cum haec dixisset dimisit ecclesiam
ACTS|20|1|postquam autem cessavit tumultus vocatis Paulus discipulis et exhortatus eos valedixit et profectus est ut iret in Macedoniam
ACTS|20|2|cum autem perambulasset partes illas et exhortatus eos fuisset multo sermone venit ad Graeciam
ACTS|20|3|ubi cum fecisset menses tres factae sunt illi insidiae a Iudaeis navigaturo in Syriam habuitque consilium ut reverteretur per Macedoniam
ACTS|20|4|comitatus est autem eum Sopater Pyrri Beroensis Thessalonicensium vero Aristarchus et Secundus et Gaius Derbeus et Timotheus Asiani vero Tychicus et Trophimus
ACTS|20|5|hii cum praecessissent sustinebant nos Troade
ACTS|20|6|nos vero navigavimus post dies azymorum a Philippis et venimus ad eos Troadem in diebus quinque ubi demorati sumus diebus septem
ACTS|20|7|in una autem sabbati cum convenissemus ad frangendum panem Paulus disputabat eis profecturus in crastinum protraxitque sermonem usque in mediam noctem
ACTS|20|8|erant autem lampades copiosae in cenaculo ubi eramus congregati
ACTS|20|9|sedens autem quidam adulescens nomine Eutychus super fenestram cum mergeretur somno gravi disputante diu Paulo eductus somno cecidit de tertio cenaculo deorsum et sublatus est mortuus
ACTS|20|10|ad quem cum descendisset Paulus incubuit super eum et conplexus dixit nolite turbari anima enim ipsius in eo est
ACTS|20|11|ascendens autem frangensque panem et gustans satisque adlocutus usque in lucem sic profectus est
ACTS|20|12|adduxerunt autem puerum viventem et consolati sunt non minime
ACTS|20|13|nos autem ascendentes navem enavigavimus in Asson inde suscepturi Paulum sic enim disposuerat ipse per terram iter facturus
ACTS|20|14|cum autem convenisset nos in Asson adsumpto eo venimus Mytilenen
ACTS|20|15|et inde navigantes sequenti die venimus contra Chium et alia adplicuimus Samum et sequenti venimus Miletum
ACTS|20|16|proposuerat enim Paulus transnavigare Ephesum ne qua mora illi fieret in Asia festinabat enim si possibile sibi esset ut diem pentecosten faceret Hierosolymis
ACTS|20|17|a Mileto autem mittens Ephesum vocavit maiores natu ecclesiae
ACTS|20|18|qui cum venissent ad eum et simul essent dixit eis vos scitis a prima die qua ingressus sum in Asiam qualiter vobiscum per omne tempus fuerim
ACTS|20|19|serviens Domino cum omni humilitate et lacrimis et temptationibus quae mihi acciderunt ex insidiis Iudaeorum
ACTS|20|20|quomodo nihil subtraxerim utilium quo minus adnuntiarem vobis et docerem vos publice et per domos
ACTS|20|21|testificans Iudaeis atque gentilibus in Deum paenitentiam et fidem in Dominum nostrum Iesum Christum
ACTS|20|22|et nunc ecce alligatus ego Spiritu vado in Hierusalem quae in ea eventura sint mihi ignorans
ACTS|20|23|nisi quod Spiritus Sanctus per omnes civitates protestatur mihi dicens quoniam vincula et tribulationes me manent
ACTS|20|24|sed nihil horum vereor nec facio animam pretiosiorem quam me dummodo consummem cursum meum et ministerium quod accepi a Domino Iesu testificari evangelium gratiae Dei
ACTS|20|25|et nunc ecce ego scio quia amplius non videbitis faciem meam vos omnes per quos transivi praedicans regnum Dei
ACTS|20|26|quapropter contestor vos hodierna die quia mundus sum a sanguine omnium
ACTS|20|27|non enim subterfugi quo minus adnuntiarem omne consilium Dei vobis
ACTS|20|28|adtendite vobis et universo gregi in quo vos Spiritus Sanctus posuit episcopos regere ecclesiam Dei quam adquisivit sanguine suo
ACTS|20|29|ego scio quoniam intrabunt post discessionem meam lupi graves in vos non parcentes gregi
ACTS|20|30|et ex vobis ipsis exsurgent viri loquentes perversa ut abducant discipulos post se
ACTS|20|31|propter quod vigilate memoria retinentes quoniam per triennium nocte et die non cessavi cum lacrimis monens unumquemque vestrum
ACTS|20|32|et nunc commendo vos Deo et verbo gratiae ipsius qui potens est aedificare et dare hereditatem in sanctificatis omnibus
ACTS|20|33|argentum aut aurum aut vestem nullius concupivi
ACTS|20|34|ipsi scitis quoniam ad ea quae mihi opus erant et his qui mecum sunt ministraverunt manus istae
ACTS|20|35|omnia ostendi vobis quoniam sic laborantes oportet suscipere infirmos ac meminisse verbi Domini Iesu quoniam ipse dixit beatius est magis dare quam accipere
ACTS|20|36|et cum haec dixisset positis genibus suis cum omnibus illis oravit
ACTS|20|37|magnus autem fletus factus est omnium et procumbentes super collum Pauli osculabantur eum
ACTS|20|38|dolentes maxime in verbo quo dixerat quoniam amplius faciem eius non essent visuri et deducebant eum ad navem
ACTS|21|1|cum autem factum esset ut navigaremus abstracti ab eis recto cursu venimus Cho et sequenti die Rhodum et inde Patara
ACTS|21|2|et cum invenissemus navem transfretantem in Foenicen ascendentes navigavimus
ACTS|21|3|cum paruissemus autem Cypro et relinquentes eam ad sinistram navigabamus in Syriam et venimus Tyrum ibi enim navis erat expositura onus
ACTS|21|4|inventis autem discipulis mansimus ibi diebus septem qui Paulo dicebant per Spiritum ne ascenderet Hierosolymam
ACTS|21|5|et explicitis diebus profecti ibamus deducentibus nos omnibus cum uxoribus et filiis usque foras civitatem et positis genibus in litore oravimus
ACTS|21|6|et cum valefecissemus invicem ascendimus in navem illi autem redierunt in sua
ACTS|21|7|nos vero navigatione explicita a Tyro descendimus Ptolomaida et salutatis fratribus mansimus die una apud illos
ACTS|21|8|alia autem die profecti venimus Caesaream et intrantes in domum Philippi evangelistae qui erat de septem mansimus apud eum
ACTS|21|9|huic autem erant filiae quattuor virgines prophetantes
ACTS|21|10|et cum moraremur per dies aliquot supervenit quidam a Iudaea propheta nomine Agabus
ACTS|21|11|is cum venisset ad nos tulit zonam Pauli et alligans sibi pedes et manus dixit haec dicit Spiritus Sanctus virum cuius est zona haec sic alligabunt in Hierusalem Iudaei et tradent in manus gentium
ACTS|21|12|quod cum audissemus rogabamus nos et qui loci illius erant ne ascenderet Hierosolymam
ACTS|21|13|tunc respondit Paulus et dixit quid facitis flentes et adfligentes cor meum ego enim non solum alligari sed et mori in Hierusalem paratus sum propter nomen Domini Iesu
ACTS|21|14|et cum ei suadere non possemus quievimus dicentes Domini voluntas fiat
ACTS|21|15|post dies autem istos praeparati ascendebamus Hierusalem
ACTS|21|16|venerunt autem et ex discipulis a Caesarea nobiscum adducentes apud quem hospitaremur Mnasonem quendam Cyprium antiquum discipulum
ACTS|21|17|et cum venissemus Hierosolymam libenter exceperunt nos fratres
ACTS|21|18|sequenti autem die introibat Paulus nobiscum ad Iacobum omnesque collecti sunt seniores
ACTS|21|19|quos cum salutasset narrabat per singula quae fecisset Deus in gentibus per ministerium ipsius
ACTS|21|20|at illi cum audissent magnificabant Deum dixeruntque ei vides frater quot milia sint in Iudaeis qui crediderunt et omnes aemulatores sunt legis
ACTS|21|21|audierunt autem de te quia discessionem doceas a Mose eorum qui per gentes sunt Iudaeorum dicens non debere circumcidere eos filios suos neque secundum consuetudinem ingredi
ACTS|21|22|quid ergo est utique oportet convenire multitudinem audient enim te supervenisse
ACTS|21|23|hoc ergo fac quod tibi dicimus sunt nobis viri quattuor votum habentes super se
ACTS|21|24|his adsumptis sanctifica te cum illis et inpende in illis ut radant capita et scient omnes quia quae de te audierunt falsa sunt sed ambulas et ipse custodiens legem
ACTS|21|25|de his autem qui crediderunt ex gentibus nos scripsimus iudicantes ut abstineant se ab idolis immolato et sanguine et suffocato et fornicatione
ACTS|21|26|tunc Paulus adsumptis viris postera die purificatus cum illis intravit in templum adnuntians expletionem dierum purificationis donec offerretur pro unoquoque eorum oblatio
ACTS|21|27|dum autem septem dies consummarentur hii qui de Asia erant Iudaei cum vidissent eum in templo concitaverunt omnem populum et iniecerunt ei manus clamantes
ACTS|21|28|viri israhelitae adiuvate hic est homo qui adversus populum et legem et locum hunc omnes ubique docens insuper et gentiles induxit in templum et violavit sanctum locum istum
ACTS|21|29|viderant enim Trophimum Ephesium in civitate cum ipso quem aestimaverunt quoniam in templum induxisset Paulus
ACTS|21|30|commotaque est civitas tota et facta est concursio populi et adprehendentes Paulum trahebant eum extra templum et statim clausae sunt ianuae
ACTS|21|31|quaerentibus autem eum occidere nuntiatum est tribuno cohortis quia tota confunditur Hierusalem
ACTS|21|32|qui statim adsumptis militibus et centurionibus decucurrit ad illos qui cum vidissent tribunum et milites cessaverunt percutere Paulum
ACTS|21|33|tunc accedens tribunus adprehendit eum et iussit alligari catenis duabus et interrogabat quis esset et quid fecisset
ACTS|21|34|alii autem aliud clamabant in turba et cum non posset certum cognoscere prae tumultu iussit duci eum in castra
ACTS|21|35|et cum venisset ad gradus contigit ut portaretur a militibus propter vim populi
ACTS|21|36|sequebatur enim multitudo populi clamans tolle eum
ACTS|21|37|et cum coepisset induci in castra Paulus dicit tribuno si licet mihi loqui aliquid ad te qui dixit graece nosti
ACTS|21|38|nonne tu es Aegyptius qui ante hos dies tumultum concitasti et eduxisti in desertum quattuor milia virorum sicariorum
ACTS|21|39|et dixit ad eum Paulus ego homo sum quidem iudaeus a Tarso Ciliciae non ignotae civitatis municeps rogo autem te permitte mihi loqui ad populum
ACTS|21|40|et cum ille permisisset Paulus stans in gradibus annuit manu ad plebem et magno silentio facto adlocutus est hebraea lingua dicens
ACTS|22|1|viri fratres et patres audite quam ad vos nunc reddo rationem
ACTS|22|2|cum audissent autem quia hebraea lingua loquitur ad illos magis praestiterunt silentium
ACTS|22|3|et dixit ego sum vir iudaeus natus Tarso Ciliciae nutritus autem in ista civitate secus pedes Gamalihel eruditus iuxta veritatem paternae legis aemulator legis sicut et vos omnes estis hodie
ACTS|22|4|qui hanc viam persecutus sum usque ad mortem alligans et tradens in custodias viros ac mulieres
ACTS|22|5|sicut princeps sacerdotum testimonium mihi reddit et omnes maiores natu a quibus et epistulas accipiens ad fratres Damascum pergebam ut adducerem inde vinctos in Hierusalem uti punirentur
ACTS|22|6|factum est autem eunte me et adpropinquante Damasco media die subito de caelo circumfulsit me lux copiosa
ACTS|22|7|et decidens in terram audivi vocem dicentem mihi Saule Saule quid me persequeris
ACTS|22|8|ego autem respondi quis es Domine dixitque ad me ego sum Iesus Nazarenus quem tu persequeris
ACTS|22|9|et qui mecum erant lumen quidem viderunt vocem autem non audierunt eius qui loquebatur mecum
ACTS|22|10|et dixi quid faciam Domine Dominus autem dixit ad me surgens vade Damascum et ibi tibi dicetur de omnibus quae te oporteat facere
ACTS|22|11|et cum non viderem prae claritate luminis illius ad manum deductus a comitibus veni Damascum
ACTS|22|12|Ananias autem quidam vir secundum legem testimonium habens ab omnibus habitantibus Iudaeis
ACTS|22|13|veniens ad me et adstans dixit mihi Saule frater respice et ego eadem hora respexi in eum
ACTS|22|14|at ille dixit Deus patrum nostrorum praeordinavit te ut cognosceres voluntatem eius et videres Iustum et audires vocem ex ore eius
ACTS|22|15|quia eris testis illius ad omnes homines eorum quae vidisti et audisti
ACTS|22|16|et nunc quid moraris exsurge baptizare et ablue peccata tua invocato nomine ipsius
ACTS|22|17|factum est autem revertenti mihi in Hierusalem et oranti in templo fieri me in stupore mentis
ACTS|22|18|et videre illum dicentem mihi festina et exi velociter ex Hierusalem quoniam non recipient testimonium tuum de me
ACTS|22|19|et ego dixi Domine ipsi sciunt quia ego eram concludens in carcerem et caedens per synagogas eos qui credebant in te
ACTS|22|20|et cum funderetur sanguis Stephani testis tui ego adstabam et consentiebam et custodiebam vestimenta interficientium illum
ACTS|22|21|et dixit ad me vade quoniam ego in nationes longe mittam te
ACTS|22|22|audiebant autem eum usque ad hoc verbum et levaverunt vocem suam dicentes tolle de terra eiusmodi non enim fas est eum vivere
ACTS|22|23|vociferantibus autem eis et proicientibus vestimenta sua et pulverem iactantibus in aerem
ACTS|22|24|iussit tribunus induci eum in castra et flagellis caedi et torqueri eum ut sciret propter quam causam sic adclamarent ei
ACTS|22|25|et cum adstrinxissent eum loris dixit adstanti sibi centurioni Paulus si hominem romanum et indemnatum licet vobis flagellare
ACTS|22|26|quo audito centurio accessit ad tribunum et nuntiavit dicens quid acturus es hic enim homo civis romanus est
ACTS|22|27|accedens autem tribunus dixit illi dic mihi tu Romanus es at ille dixit etiam
ACTS|22|28|et respondit tribunus ego multa summa civitatem hanc consecutus sum et Paulus ait ego autem et natus sum
ACTS|22|29|protinus ergo discesserunt ab illo qui eum torturi erant tribunus quoque timuit postquam rescivit quia civis romanus esset et quia alligasset eum
ACTS|22|30|postera autem die volens scire diligentius qua ex causa accusaretur a Iudaeis solvit eum et iussit sacerdotes convenire et omne concilium et producens Paulum statuit inter illos
ACTS|23|1|intendens autem concilium Paulus ait viri fratres ego omni conscientia bona conversatus sum ante Deum usque in hodiernum diem
ACTS|23|2|princeps autem sacerdotum Ananias praecepit adstantibus sibi percutere os eius
ACTS|23|3|tunc Paulus ad eum dixit percutiet te Deus paries dealbate et tu sedens iudicas me secundum legem et contra legem iubes me percuti
ACTS|23|4|et qui adstabant dixerunt summum sacerdotem Dei maledicis
ACTS|23|5|dixit autem Paulus nesciebam fratres quia princeps est sacerdotum scriptum est enim principem populi tui non maledices
ACTS|23|6|sciens autem Paulus quia una pars esset Sadducaeorum et altera Pharisaeorum exclamavit in concilio viri fratres ego Pharisaeus sum filius Pharisaeorum de spe et resurrectione mortuorum ego iudicor
ACTS|23|7|et cum haec dixisset facta est dissensio inter Pharisaeos et Sadducaeos et soluta est multitudo
ACTS|23|8|Sadducaei enim dicunt non esse resurrectionem neque angelum neque spiritum Pharisaei autem utrumque confitentur
ACTS|23|9|factus est autem clamor magnus et surgentes quidam Pharisaeorum pugnabant dicentes nihil mali invenimus in homine isto quod si spiritus locutus est ei aut angelus
ACTS|23|10|et cum magna dissensio facta esset timens tribunus ne discerperetur Paulus ab ipsis iussit milites descendere et rapere eum de medio eorum ac deducere eum in castra
ACTS|23|11|sequenti autem nocte adsistens ei Dominus ait constans esto sicut enim testificatus es de me Hierusalem sic te oportet et Romae testificari
ACTS|23|12|facta autem die collegerunt se quidam ex Iudaeis et devoverunt se dicentes neque manducaturos neque bibituros donec occiderent Paulum
ACTS|23|13|erant autem plus quam quadraginta qui hanc coniurationem fecerant
ACTS|23|14|qui accesserunt ad principes sacerdotum et seniores et dixerunt devotione devovimus nos nihil gustaturos donec occidamus Paulum
ACTS|23|15|nunc ergo vos notum facite tribuno cum concilio ut producat illum ad vos tamquam aliquid certius cognituri de eo nos vero priusquam adpropiet parati sumus interficere illum
ACTS|23|16|quod cum audisset filius sororis Pauli insidias venit et intravit in castra nuntiavitque Paulo
ACTS|23|17|vocans autem Paulus ad se unum ex centurionibus ait adulescentem hunc perduc ad tribunum habet enim aliquid indicare illi
ACTS|23|18|et ille quidem adsumens eum duxit ad tribunum et ait vinctus Paulus vocans rogavit me hunc adulescentem perducere ad te habentem aliquid loqui tibi
ACTS|23|19|adprehendens autem tribunus manum illius secessit cum eo seorsum et interrogavit illum quid est quod habes indicare mihi
ACTS|23|20|ille autem dixit Iudaeis convenit rogare te ut crastina die Paulum producas in concilium quasi aliquid certius inquisituri sint de illo
ACTS|23|21|tu vero ne credideris illis insidiantur enim ei ex eis viri amplius quadraginta qui se devoverunt non manducare neque bibere donec interficiant eum et nunc parati sunt expectantes promissum tuum
ACTS|23|22|tribunus igitur dimisit adulescentem praecipiens ne cui loqueretur quoniam haec nota sibi fecisset
ACTS|23|23|et vocatis duobus centurionibus dixit illis parate milites ducentos ut eant usque Caesaream et equites septuaginta et lancearios ducentos a tertia hora noctis
ACTS|23|24|et iumenta praeparate ut inponentes Paulum salvum perducerent ad Felicem praesidem
ACTS|23|25|
ACTS|23|26|scribens epistulam continentem haec Claudius Lysias optimo praesidi Felici salutem
ACTS|23|27|virum hunc conprehensum a Iudaeis et incipientem interfici ab eis superveniens cum exercitu eripui cognito quia Romanus est
ACTS|23|28|volensque scire causam quam obiciebant illi deduxi eum in concilium eorum
ACTS|23|29|quem inveni accusari de quaestionibus legis ipsorum nihil vero dignum morte aut vinculis habentem crimen
ACTS|23|30|et cum mihi perlatum esset de insidiis quas paraverunt ei misi ad te denuntians et accusatoribus ut dicant apud te
ACTS|23|31|milites ergo secundum praeceptum sibi adsumentes Paulum duxerunt per noctem in Antipatridem
ACTS|23|32|et postera die dimissis equitibus ut irent cum eo reversi sunt ad castra
ACTS|23|33|qui cum venissent Caesaream et tradidissent epistulam praesidi statuerunt ante illum et Paulum
ACTS|23|34|cum legisset autem et interrogasset de qua provincia esset et cognoscens quia de Cilicia
ACTS|23|35|audiam te inquit cum et accusatores tui venerint iussitque in praetorio Herodis custodiri eum
ACTS|24|1|post quinque autem dies descendit princeps sacerdotum Ananias cum senioribus quibusdam et Tertullo quodam oratore qui adierunt praesidem adversus Paulum
ACTS|24|2|et citato Paulo coepit accusare Tertullus dicens cum in multa pace agamus per te et multa corrigantur per tuam providentiam
ACTS|24|3|semper et ubique suscipimus optime Felix cum omni gratiarum actione
ACTS|24|4|ne diutius autem te protraham oro breviter audias nos pro tua clementia
ACTS|24|5|invenimus hunc hominem pestiferum et concitantem seditiones omnibus Iudaeis in universo orbe et auctorem seditionis sectae Nazarenorum
ACTS|24|6|qui etiam templum violare conatus est quem et adprehendimus
ACTS|24|7|
ACTS|24|8|a quo poteris ipse iudicans de omnibus istis cognoscere de quibus nos accusamus eum
ACTS|24|9|adiecerunt autem et Iudaei dicentes haec ita se habere
ACTS|24|10|respondit autem Paulus annuente sibi praeside dicere ex multis annis esse te iudicem genti huic sciens bono animo pro me satisfaciam
ACTS|24|11|potes enim cognoscere quia non plus sunt dies mihi quam duodecim ex quo ascendi adorare in Hierusalem
ACTS|24|12|et neque in templo invenerunt me cum aliquo disputantem aut concursum facientem turbae neque in synagogis neque in civitate
ACTS|24|13|neque probare possunt tibi de quibus nunc accusant me
ACTS|24|14|confiteor autem hoc tibi quod secundum sectam quam dicunt heresim sic deservio patrio Deo meo credens omnibus quae in lege et prophetis scripta sunt
ACTS|24|15|spem habens in Deum quam et hii ipsi expectant resurrectionem futuram iustorum et iniquorum
ACTS|24|16|in hoc et ipse studeo sine offendiculo conscientiam habere ad Deum et ad homines semper
ACTS|24|17|post annos autem plures elemosynas facturus in gentem meam veni et oblationes et vota
ACTS|24|18|in quibus invenerunt me purificatum in templo non cum turba neque cum tumultu
ACTS|24|19|quidam autem ex Asia Iudaei quos oportebat apud te praesto esse et accusare si quid haberent adversum me
ACTS|24|20|aut hii ipsi dicant si quid invenerunt in me iniquitatis cum stem in concilio
ACTS|24|21|nisi de una hac solummodo voce qua clamavi inter eos stans quoniam de resurrectione mortuorum ego iudicor hodie a vobis
ACTS|24|22|distulit autem illos Felix certissime sciens de via dicens cum tribunus Lysias descenderit audiam vos
ACTS|24|23|iussitque centurioni custodiri eum et habere requiem nec quemquam prohibere de suis ministrare ei
ACTS|24|24|post aliquot autem dies veniens Felix cum Drusilla uxore sua quae erat Iudaea vocavit Paulum et audivit ab eo fidem quae est in Iesum Christum
ACTS|24|25|disputante autem illo de iustitia et castitate et de iudicio futuro timefactus Felix respondit quod nunc adtinet vade tempore autem oportuno accersiam te
ACTS|24|26|simul et sperans quia pecunia daretur a Paulo propter quod et frequenter accersiens eum loquebatur cum eo
ACTS|24|27|biennio autem expleto accepit successorem Felix Porcium Festum volens autem gratiam praestare Iudaeis Felix reliquit Paulum vinctum
ACTS|25|1|Festus ergo cum venisset in provinciam post triduum ascendit Hierosolymam a Caesarea
ACTS|25|2|adieruntque eum principes sacerdotum et primi Iudaeorum adversus Paulum et rogabant eum
ACTS|25|3|postulantes gratiam adversum eum ut iuberet perduci eum Hierusalem insidias tendentes ut eum interficerent in via
ACTS|25|4|Festus autem respondit servari Paulum in Caesarea se autem maturius profecturum
ACTS|25|5|qui ergo in vobis ait potentes sunt descendentes simul si quod est in viro crimen accusent eum
ACTS|25|6|demoratus autem inter eos dies non amplius quam octo aut decem descendit Caesaream et altera die sedit pro tribunali et iussit Paulum adduci
ACTS|25|7|qui cum perductus esset circumsteterunt eum qui ab Hierosolyma descenderant Iudaei multas et graves causas obicientes quas non poterant probare
ACTS|25|8|Paulo autem rationem reddente quoniam neque in legem Iudaeorum neque in templum neque in Caesarem quicquam peccavi
ACTS|25|9|Festus autem volens Iudaeis gratiam praestare respondens Paulo dixit vis Hierosolymam ascendere et ibi de his iudicari apud me
ACTS|25|10|dixit autem Paulus ad tribunal Caesaris sto ubi me oportet iudicari Iudaeis non nocui sicut tu melius nosti
ACTS|25|11|si enim nocui aut dignum morte aliquid feci non recuso mori si vero nihil est eorum quae hii accusant me nemo potest me illis donare Caesarem appello
ACTS|25|12|tunc Festus cum consilio locutus respondit Caesarem appellasti ad Caesarem ibis
ACTS|25|13|et cum dies aliquot transacti essent Agrippa rex et Bernice descenderunt Caesaream ad salutandum Festum
ACTS|25|14|et cum dies plures ibi demorarentur Festus regi indicavit de Paulo dicens vir quidam est derelictus a Felice vinctus
ACTS|25|15|de quo cum essem Hierosolymis adierunt me principes sacerdotum et seniores Iudaeorum postulantes adversus illum damnationem
ACTS|25|16|ad quos respondi quia non est consuetudo Romanis donare aliquem hominem priusquam is qui accusatur praesentes habeat accusatores locumque defendendi accipiat ad abluenda crimina
ACTS|25|17|cum ergo huc convenissent sine ulla dilatione sequenti die sedens pro tribunali iussi adduci virum
ACTS|25|18|de quo cum stetissent accusatores nullam causam deferebant de quibus ego suspicabar malum
ACTS|25|19|quaestiones vero quasdam de sua superstitione habebant adversus eum et de quodam Iesu defuncto quem adfirmabat Paulus vivere
ACTS|25|20|haesitans autem ego de huiusmodi quaestione dicebam si vellet ire Hierosolymam et ibi iudicari de istis
ACTS|25|21|Paulo autem appellante ut servaretur ad Augusti cognitionem iussi servari eum donec mittam eum ad Caesarem
ACTS|25|22|Agrippa autem ad Festum volebam et ipse hominem audire cras inquit audies eum
ACTS|25|23|altera autem die cum venisset Agrippa et Bernice cum multa ambitione et introissent in auditorium cum tribunis et viris principalibus civitatis et iubente Festo adductus est Paulus
ACTS|25|24|et dixit Festus Agrippa rex et omnes qui simul adestis nobiscum viri videtis hunc de quo omnis multitudo Iudaeorum interpellavit me Hierosolymis petens et hic clamantes non oportere eum vivere amplius
ACTS|25|25|ego vero conperi nihil dignum eum morte admisisse ipso autem hoc appellante Augustum iudicavi mittere
ACTS|25|26|de quo quid certum scribam domino non habeo propter quod produxi eum ad vos et maxime ad te rex Agrippa ut interrogatione facta habeam quid scribam
ACTS|25|27|sine ratione enim mihi videtur mittere vinctum et causas eius non significare
ACTS|26|1|Agrippa vero ad Paulum ait permittitur tibi loqui pro temet ipso tunc Paulus extenta manu coepit rationem reddere
ACTS|26|2|de omnibus quibus accusor a Iudaeis rex Agrippa aestimo me beatum apud te cum sim defensurus me hodie
ACTS|26|3|maxime te sciente omnia quae apud Iudaeos sunt consuetudines et quaestiones propter quod obsecro patienter me audias
ACTS|26|4|et quidem vitam meam a iuventute quae ab initio fuit in gente mea in Hierosolymis noverunt omnes Iudaei
ACTS|26|5|praescientes me ab initio si velint testimonium perhibere quoniam secundum certissimam sectam nostrae religionis vixi Pharisaeus
ACTS|26|6|et nunc in spe quae ad patres nostros repromissionis facta est a Deo sto iudicio subiectus
ACTS|26|7|in quam duodecim tribus nostrae nocte ac die deservientes sperant devenire de qua spe accusor a Iudaeis rex
ACTS|26|8|quid incredibile iudicatur apud vos si Deus mortuos suscitat
ACTS|26|9|et ego quidem existimaveram me adversus nomen Iesu Nazareni debere multa contraria agere
ACTS|26|10|quod et feci Hierosolymis et multos sanctorum ego in carceribus inclusi a principibus sacerdotum potestate accepta et cum occiderentur detuli sententiam
ACTS|26|11|et per omnes synagogas frequenter puniens eos conpellebam blasphemare et amplius insaniens in eos persequebar usque in exteras civitates
ACTS|26|12|in quibus dum irem Damascum cum potestate et permissu principum sacerdotum
ACTS|26|13|die media in via vidi rex de caelo supra splendorem solis circumfulsisse me lumen et eos qui mecum simul erant
ACTS|26|14|omnesque nos cum decidissemus in terram audivi vocem loquentem mihi hebraica lingua Saule Saule quid me persequeris durum est tibi contra stimulum calcitrare
ACTS|26|15|ego autem dixi quis es Domine Dominus autem dixit ego sum Iesus quem tu persequeris
ACTS|26|16|sed exsurge et sta super pedes tuos ad hoc enim apparui tibi ut constituam te ministrum et testem eorum quae vidisti et eorum quibus apparebo tibi
ACTS|26|17|eripiens te de populo et gentibus in quas nunc ego mitto te
ACTS|26|18|aperire oculos eorum ut convertantur a tenebris ad lucem et de potestate Satanae ad Deum ut accipiant remissionem peccatorum et sortem inter sanctos per fidem quae est in me
ACTS|26|19|unde rex Agrippa non fui incredulus caelestis visionis
ACTS|26|20|sed his qui sunt Damasci primum et Hierosolymis et in omnem regionem Iudaeae et gentibus adnuntiabam ut paenitentiam agerent et converterentur ad Deum digna paenitentiae opera facientes
ACTS|26|21|hac ex causa me Iudaei cum essem in templo conprehensum temptabant interficere
ACTS|26|22|auxilio autem adiutus Dei usque in hodiernum diem sto testificans minori atque maiori nihil extra dicens quam ea quae prophetae sunt locuti futura esse et Moses
ACTS|26|23|si passibilis Christus si primus ex resurrectione mortuorum lumen adnuntiaturus est populo et gentibus
ACTS|26|24|haec loquente eo et rationem reddente Festus magna voce dixit insanis Paule multae te litterae ad insaniam convertunt
ACTS|26|25|at Paulus non insanio inquit optime Feste sed veritatis et sobrietatis verba eloquor
ACTS|26|26|scit enim de his rex ad quem et constanter loquor latere enim eum nihil horum arbitror neque enim in angulo quicquam horum gestum est
ACTS|26|27|credis rex Agrippa prophetis scio quia credis
ACTS|26|28|Agrippa autem ad Paulum in modico suades me Christianum fieri
ACTS|26|29|et Paulus opto apud Deum et in modico et in magno non tantum te sed et omnes hos qui audiunt hodie fieri tales qualis et ego sum exceptis vinculis his
ACTS|26|30|et exsurrexit rex et praeses et Bernice et qui adsidebant eis
ACTS|26|31|et cum secessissent loquebantur ad invicem dicentes quia nihil morte aut vinculorum dignum quid facit homo iste
ACTS|26|32|Agrippa autem Festo dixit dimitti poterat homo hic si non appellasset Caesarem
ACTS|27|1|ut autem iudicatum est eum navigare in Italiam et tradi Paulum cum reliquis custodiis centurioni nomine Iulio cohortis Augustae
ACTS|27|2|ascendentes autem navem hadrumetinam incipientem navigare circa Asiae loca sustulimus perseverante nobiscum Aristarcho Macedone Thessalonicense
ACTS|27|3|sequenti autem die devenimus Sidonem humane autem tractans Iulius Paulum permisit ad amicos ire et curam sui agere
ACTS|27|4|et inde cum sustulissemus subnavigavimus Cypro propterea quod essent venti contrarii
ACTS|27|5|et pelagus Ciliciae et Pamphiliae navigantes venimus Lystram quae est Lyciae
ACTS|27|6|et ibi inveniens centurio navem alexandrinam navigantem in Italiam transposuit nos in eam
ACTS|27|7|et cum multis diebus tarde navigaremus et vix devenissemus contra Cnidum prohibente nos vento adnavigavimus Cretae secundum Salmonem
ACTS|27|8|et vix iuxta navigantes venimus in locum quendam qui vocatur Boni portus cui iuxta erat civitas Thalassa
ACTS|27|9|multo autem tempore peracto et cum iam non esset tuta navigatio eo quod et ieiunium iam praeterisset consolabatur Paulus
ACTS|27|10|dicens eis viri video quoniam cum iniuria et multo damno non solum oneris et navis sed etiam animarum nostrarum incipit esse navigatio
ACTS|27|11|centurio autem gubernatori et nauclerio magis credebat quam his quae a Paulo dicebantur
ACTS|27|12|et cum aptus portus non esset ad hiemandum plurimi statuerunt consilium navigare inde si quo modo possent devenientes Phoenice hiemare portum Cretae respicientem ad africum et ad chorum
ACTS|27|13|adspirante autem austro aestimantes propositum se tenere cum sustulissent de Asson legebant Cretam
ACTS|27|14|non post multum autem misit se contra ipsam ventus typhonicus qui vocatur euroaquilo
ACTS|27|15|cumque arrepta esset navis et non posset conari in ventum data nave flatibus ferebamur
ACTS|27|16|insulam autem quandam decurrentes quae vocatur Caudam potuimus vix obtinere scapham
ACTS|27|17|qua sublata adiutoriis utebantur accingentes navem timentes ne in Syrtim inciderent submisso vase sic ferebantur
ACTS|27|18|valide autem nobis tempestate iactatis sequenti die iactum fecerunt
ACTS|27|19|et tertia die suis manibus armamenta navis proiecerunt
ACTS|27|20|neque sole autem neque sideribus apparentibus per plures dies et tempestate non exigua inminente iam ablata erat spes omnis salutis nostrae
ACTS|27|21|et cum multa ieiunatio fuisset tunc stans Paulus in medio eorum dixit oportebat quidem o viri audito me non tollere a Creta lucrique facere iniuriam hanc et iacturam
ACTS|27|22|et nunc suadeo vobis bono animo esse amissio enim nullius animae erit ex vobis praeterquam navis
ACTS|27|23|adstitit enim mihi hac nocte angelus Dei cuius sum ego et cui deservio
ACTS|27|24|dicens ne timeas Paule Caesari te oportet adsistere et ecce donavit tibi Deus omnes qui navigant tecum
ACTS|27|25|propter quod bono animo estote viri credo enim Deo quia sic erit quemadmodum dictum est mihi
ACTS|27|26|in insulam autem quandam oportet nos devenire
ACTS|27|27|sed posteaquam quartadecima nox supervenit navigantibus nobis in Hadria circa mediam noctem suspicabantur nautae apparere sibi aliquam regionem
ACTS|27|28|qui submittentes invenerunt passus viginti et pusillum inde separati invenerunt passus quindecim
ACTS|27|29|timentes autem ne in aspera loca incideremus de puppi mittentes anchoras quattuor optabant diem fieri
ACTS|27|30|nautis vero quaerentibus fugere de navi cum misissent scapham in mare sub obtentu quasi a prora inciperent anchoras extendere
ACTS|27|31|dixit Paulus centurioni et militibus nisi hii in navi manserint vos salvi fieri non potestis
ACTS|27|32|tunc absciderunt milites funes scaphae et passi sunt eam excidere
ACTS|27|33|et cum lux inciperet fieri rogabat Paulus omnes sumere cibum dicens quartadecima hodie die expectantes ieiuni permanetis nihil accipientes
ACTS|27|34|propter quod rogo vos accipere cibum pro salute vestra quia nullius vestrum capillus de capite peribit
ACTS|27|35|et cum haec dixisset sumens panem gratias egit Deo in conspectu omnium et cum fregisset coepit manducare
ACTS|27|36|animaequiores autem facti omnes et ipsi adsumpserunt cibum
ACTS|27|37|eramus vero universae animae in navi ducentae septuaginta sex
ACTS|27|38|et satiati cibo adleviabant navem iactantes triticum in mare
ACTS|27|39|cum autem dies factus esset terram non agnoscebant sinum vero quendam considerabant habentem litus in quem cogitabant si possent eicere navem
ACTS|27|40|et cum anchoras abstulissent committebant se mari simul laxantes iuncturas gubernaculorum et levato artemone secundum flatum aurae tendebant ad litus
ACTS|27|41|et cum incidissemus in locum bithalassum inpegerunt navem et prora quidem fixa manebat inmobilis puppis vero solvebatur a vi maris
ACTS|27|42|militum autem consilium fuit ut custodias occiderent ne quis cum enatasset effugeret
ACTS|27|43|centurio autem volens servare Paulum prohibuit fieri iussitque eos qui possent natare mittere se primos et evadere et ad terram exire
ACTS|27|44|et ceteros alios in tabulis ferebant quosdam super ea quae de navi essent et sic factum est ut omnes animae evaderent ad terram
ACTS|28|1|et cum evasissemus tunc cognovimus quia Militene insula vocatur barbari vero praestabant non modicam humanitatem nobis
ACTS|28|2|accensa enim pyra reficiebant nos omnes propter imbrem qui inminebat et frigus
ACTS|28|3|cum congregasset autem Paulus sarmentorum aliquantam multitudinem et inposuisset super ignem vipera a calore cum processisset invasit manum eius
ACTS|28|4|ut vero viderunt barbari pendentem bestiam de manu eius ad invicem dicebant utique homicida est homo hic qui cum evaserit de mari Ultio non sinit vivere
ACTS|28|5|et ille quidem excutiens bestiam in ignem nihil mali passus est
ACTS|28|6|at illi existimabant eum in tumorem convertendum et subito casurum et mori diu autem illis sperantibus et videntibus nihil mali in eo fieri convertentes se dicebant eum esse deum
ACTS|28|7|in locis autem illis erant praedia principis insulae nomine Publii qui nos suscipiens triduo benigne exhibuit
ACTS|28|8|contigit autem patrem Publii febribus et dysenteria vexatum iacere ad quem Paulus intravit et cum orasset et inposuisset ei manus salvavit eum
ACTS|28|9|quo facto et omnes qui in insula habebant infirmitates accedebant et curabantur
ACTS|28|10|qui etiam multis honoribus nos honoraverunt et navigantibus inposuerunt quae necessaria erant
ACTS|28|11|post menses autem tres navigavimus in nave alexandrina quae in insula hiemaverat cui erat insigne Castorum
ACTS|28|12|et cum venissemus Syracusam mansimus ibi triduo
ACTS|28|13|inde circumlegentes devenimus Regium et post unum diem flante austro secunda die venimus Puteolos
ACTS|28|14|ubi inventis fratribus rogati sumus manere apud eos dies septem et sic venimus Romam
ACTS|28|15|et inde cum audissent fratres occurrerunt nobis usque ad Appii Forum et Tribus Tabernis quos cum vidisset Paulus gratias agens Deo accepit fiduciam
ACTS|28|16|cum venissemus autem Romam permissum est Paulo manere sibimet cum custodiente se milite
ACTS|28|17|post tertium autem diem convocavit primos Iudaeorum cumque convenissent dicebat eis ego viri fratres nihil adversus plebem faciens aut morem paternum vinctus ab Hierosolymis traditus sum in manus Romanorum
ACTS|28|18|qui cum interrogationem de me habuissent voluerunt me dimittere eo quod nulla causa esset mortis in me
ACTS|28|19|contradicentibus autem Iudaeis coactus sum appellare Caesarem non quasi gentem meam habens aliquid accusare
ACTS|28|20|propter hanc igitur causam rogavi vos videre et adloqui propter spem enim Israhel catena hac circumdatus sum
ACTS|28|21|at illi dixerunt ad eum nos neque litteras accepimus de te a Iudaea neque adveniens aliquis fratrum nuntiavit aut locutus est quid de te malum
ACTS|28|22|rogamus autem a te audire quae sentis nam de secta hac notum est nobis quia ubique ei contradicitur
ACTS|28|23|cum constituissent autem illi diem venerunt ad eum in hospitium plures quibus exponebat testificans regnum Dei suadensque eos de Iesu ex lege Mosi et prophetis a mane usque ad vesperam
ACTS|28|24|et quidam credebant his quae dicebantur quidam vero non credebant
ACTS|28|25|cumque invicem non essent consentientes discedebant dicente Paulo unum verbum quia bene Spiritus Sanctus locutus est per Esaiam prophetam ad patres nostros
ACTS|28|26|dicens vade ad populum istum et dic aure audietis et non intellegetis et videntes videbitis et non perspicietis
ACTS|28|27|incrassatum est enim cor populi huius et auribus graviter audierunt et oculos suos conpresserunt ne forte videant oculis et auribus audiant et corde intellegant et convertantur et sanem illos
ACTS|28|28|notum ergo sit vobis quoniam gentibus missum est hoc salutare Dei ipsi et audient
ACTS|28|29|
ACTS|28|30|mansit autem biennio toto in suo conducto et suscipiebat omnes qui ingrediebantur ad eum
ACTS|28|31|praedicans regnum Dei et docens quae sunt de Domino Iesu Christo cum omni fiducia sine prohibitione
