HEB|1|1|Multifariam et multis modis olim Deus locutus patribus in prophetis,
HEB|1|2|in novissimis his diebus locutus est nobis in Filio, quem constituit heredem universorum, per quem fecit et saecula;
HEB|1|3|qui, cum sit splendor gloriae et figura substantiae eius et portet omnia verbo virtutis suae, purgatione peccatorum facta, consedit ad dexteram maiestatis in excelsis,
HEB|1|4|tanto melior angelis effectus, quanto differentius prae illis nomen hereditavit.
HEB|1|5|Cui enim dixit aliquando angelorum: Filius meus es tu;ego hodie genui te "et rursum: " Ego ero illi in patrem, et ipse erit mihi in filium "?
HEB|1|6|Cum autem iterum introducit primogenitum in orbem terrae, dicit: Et adorent eum omnes angeli Dei ".
HEB|1|7|Et ad angelos quidem dicit: Qui facit angelos suos spirituset ministros suos flammam ignis ";
HEB|1|8|ad Filium autem: Thronus tuus, Deus, in saeculum saeculi,et virga aequitatis virga regni tui.
HEB|1|9|Dilexisti iustitiam et odisti iniquitatem,propterea unxit te Deus, Deus tuus,oleo exsultationis prae participibus tuis "
HEB|1|10|et: Tu in principio, Domine, terram fundasti;et opera manuum tuarum sunt caeli.
HEB|1|11|Ipsi peribunt, tu autem permanes;et omnes ut vestimentum veterascent,
HEB|1|12|et velut amictum involves eos,sicut vestimentum et mutabuntur.Tu autem idem es, et anni tui non deficient ".
HEB|1|13|Ad quem autem angelorum dixit aliquando: Sede a dextris meis,donec ponam inimicos tuos scabellum pedum tuorum "?
HEB|1|14|Nonne omnes sunt administratorii spiritus, qui in ministerium mittuntur propter eos, qui hereditatem capient salutis?
HEB|2|1|Propterea abundantius oportet observare nos ea, quae audivi mus, ne forte praeterfluamus.
HEB|2|2|Si enim, qui per angelos dictus est, sermo factus est firmus, et omnis praevaricatio et inoboedientia accepit iustam mercedis retributionem,
HEB|2|3|quomodo nos effugiemus, si tantam neglexerimus salutem? Quae, cum initium accepisset enarrari per Dominum, ab eis, qui audierunt, in nos confirmata est,
HEB|2|4|contestante Deo signis et portentis et variis virtutibus et Spiritus Sancti distributionibus secundum suam voluntatem.
HEB|2|5|Non enim angelis subiecit orbem terrae futurum, de quo loquimur.
HEB|2|6|Testatus est autem in quodam loco quis dicens: Quid est homo, quod memor es eius,aut filius hominis, quoniam visitas eum?
HEB|2|7|Minuisti eum paulo minus ab angelis,gloria et honore coronasti eum,
HEB|2|8|omnia subiecisti sub pedibus eius ".In eo enim quod ei omnia subiecit, nihil dimisit non subiectibile ei. Nunc autem necdum videmus omnia subiecta ei;
HEB|2|9|eum autem, qui paulo minus ab angelis minoratus est, videmus Iesum propter passionem mortis gloria et honore coronatum, ut gratia Dei pro omnibus gustaverit mortem.
HEB|2|10|Decebat enim eum, propter quem omnia et per quem omnia, qui multos filios in gloriam adduxit, ducem salutis eorum per passiones consummare.
HEB|2|11|Qui enim sanctificat et qui sanctificantur, ex uno omnes; propter quam causam non erubescit fratres eos vocare
HEB|2|12|dicens: Nuntiabo nomen tuum fratribus meis,in medio ecclesiae laudabo te";
HEB|2|13|et iterum: " Ego ero fidens in eum ";et iterum: " Ecce ego et pueri, quos mihi dedit Deus ".
HEB|2|14|Quia ergo pueri communicaverunt sanguini et carni, et ipse similiter participavit iisdem, ut per mortem destrueret eum, qui habebat mortis imperium, id est Diabolum,
HEB|2|15|et liberaret eos, qui timore mortis per totam vitam obnoxii erant servituti.
HEB|2|16|Nusquam enim angelos apprehendit, sed semen Abrahae apprehendit.
HEB|2|17|Unde debuit per omnia fratribus similari, ut misericors fieret et fidelis pontifex in iis,quae sunt ad Deum, ut repropitiaret delicta populi;
HEB|2|18|in quo enim passus est ipse tentatus, po tens est eis, qui tentantur, auxiliari.
HEB|3|1|Unde, fratres sancti, vocationis caelestis participes, considerate apostolum et pontificem confessionis nostrae Iesum,
HEB|3|2|qui fidelis est ei, qui fecit illum, sicut et Moyses in tota domo illius.
HEB|3|3|Amplioris enim gloriae iste prae Moyse dignus est habitus, quanto ampliorem honorem habet quam domus, qui fabricavit illam.
HEB|3|4|Omnis namque domus fabricatur ab aliquo; qui autem omnia fabricavit, Deus est.
HEB|3|5|Et Moyses quidem fidelis erat in tota domo eius tamquam famulus in testimonium eorum, quae dicenda erant,
HEB|3|6|Christus vero tamquam Filius super domum illius; cuius domus sumus nos, si fiduciam et gloriationem spei retineamus.
HEB|3|7|Quapropter, sicut dicit Spiritus Sanctus: Hodie, si vocem eius audieritis,
HEB|3|8|nolite obdurare corda vestra sicut in exacerbatione,secundum diem tentationis in deserto,
HEB|3|9|ubi tentaverunt me patres vestri in probationeet viderunt opera mea
HEB|3|10|quadraginta annos. Propter quod infensus fui generationi huic et dixi: Semper errant corde.Ipsi autem non cognoverunt vias meas;
HEB|3|11|sicut icut iuravi in ira mea:Non introibunt in requiem meam ".
HEB|3|12|Videte, fratres, ne forte sit in aliquo vestrum cor malum incredulitatis discedendi a Deo vivo,
HEB|3|13|sed adhortamini vosmetipsos per singulos dies, donec illud " hodie " vocatur, ut non obduretur quis ex vobis fallacia peccati;
HEB|3|14|participes enim Christi effecti sumus, si tamen initium substantiae usque ad finem firmum retineamus,
HEB|3|15|dum dicitur: Hodie, si vocem eius audieritis,nolite obdurare corda vestra quemadmodum in illa exacerbatione ".
HEB|3|16|Qui sunt enim qui audientes exacerbaverunt? Nonne universi, qui profecti sunt ab Aegypto per Moysen?
HEB|3|17|Quibus autem infensus fuit quadraginta annos? Nonne illis, qui peccaverunt, quorum membra ceciderunt in deserto?
HEB|3|18|Quibus autem iuravit non introire in requiem ipsius, nisi illis, qui increduli fuerunt?
HEB|3|19|Et videmus quia non potuerunt introire propter incredulitatem.
HEB|4|1|Timeamus ergo, ne forte, relicta pollicitatione introeundi in re quiem eius, existimetur aliquis ex vobis deesse;
HEB|4|2|etenim et nobis evangelizatum est quemadmodum et illis, sed non profuit illis sermo auditus, non commixtis fide cum iis, qui audierant.
HEB|4|3|Ingredimur enim in requiem, qui credidimus, quemadmodum dixit: Sicut iuravi in ira mea:Non introibunt in requiem meam ",et quidem operibus ab institutione mundi factis.
HEB|4|4|Dixit enim quodam loco de die septima sic: "Et requievit Deus die septima ab omnibus operibus suis ";
HEB|4|5|et in isto rursum: " Non introibunt in requiem meam ".
HEB|4|6|Quoniam ergo superest quosdam introire in illam, et hi, quibus prioribus evangelizatum est, non introierunt propter inoboedientiam,
HEB|4|7|iterum terminat diem quendam, " Hodie ", in David dicendo post tantum temporis, sicut supra dictum est: Hodie, si vocem eius audieritis,nolite obdurare corda vestra ".
HEB|4|8|Nam, si eis Iesus requiem praestitisset, non de alio loqueretur posthac die.
HEB|4|9|Itaque relinquitur sabbatismus populo Dei;
HEB|4|10|qui enim ingressus est in requiem eius, etiam ipse requievit ab operibus suis, sicut a suis Deus.
HEB|4|11|Festinemus ergo ingredi in illam requiem, ut ne in idipsum quis incidat inoboedientiae exemplum.
HEB|4|12|Vivus est enim Dei sermo et efficax et penetrabilior omni gladio ancipiti et pertingens usque ad divisionem animae ac spiritus, compagum quoque et medullarum, et discretor cogitationum et intentionum cordis;
HEB|4|13|et non est creatura invisibilis in conspectu eius, omnia autem nuda et aperta sunt oculis eius, ad quem nobis sermo.
HEB|4|14|Habentes ergo pontificem magnum, qui penetravit caelos, Iesum Filium Dei, teneamus confessionem.
HEB|4|15|Non enim habemus pontificem, qui non possit compati infirmitatibus nostris, tentatum autem per omnia secundum similitudinem absque peccato;
HEB|4|16|adeamus ergo cum fiducia ad thronum gratiae, ut misericordiam consequamur et gratiam inveniamus in auxilium opportunum.
HEB|5|1|Omnis namque pontifex ex hominibus assumptus pro homi nibus constituitur in his, quae sunt ad Deum, ut offerat dona et sacrificia pro peccatis;
HEB|5|2|qui aeque condolere possit his, qui ignorant et errant, quoniam et ipse circumdatus est infirmitate
HEB|5|3|et propter eam debet, quemadmodum et pro populo, ita etiam pro semetipso offerre pro peccatis.
HEB|5|4|Nec quisquam sumit sibi illum honorem, sed qui vocatur a Deo tamquam et Aaron.
HEB|5|5|Sic et Christus non semetipsum glorificavit, ut pontifex fieret, sed qui locutus est ad eum: Filius meus es tu;ego hodie genui te ";
HEB|5|6|quemadmodum et in alio dicit: Tu es sacerdos in aeternum secundum ordinem Melchisedech ".
HEB|5|7|Qui in diebus carnis suae, preces supplicationesque ad eum, qui possit salvum illum a morte facere, cum clamore valido et lacrimis offerens et exauditus pro sua reverentia,
HEB|5|8|et quidem cum esset Filius, didicit ex his, quae passus est, oboedientiam;
HEB|5|9|et, consummatus, factus est omnibus oboedientibus sibi auctor salutis aeternae,
HEB|5|10|appellatus a Deo pontifex iuxta ordinem Melchisedech.
HEB|5|11|De quo grandis nobis sermo et ininterpretabilis ad dicendum, quoniam segnes facti estis ad audiendum.
HEB|5|12|Etenim cum deberetis magistri esse propter tempus, rursum indigetis, ut vos doceat aliquis elementa exordii sermonum Dei, et facti estis, quibus lacte opus sit, non solido cibo.
HEB|5|13|Omnis enim, qui lactis est particeps, expers est sermonis iustitiae, parvulus enim est;
HEB|5|14|perfectorum autem est solidus cibus, eorum, qui pro consuetudine exercitatos habent sensus ad discretionem boni ac mali.
HEB|6|1|Quapropter praetermittentes inchoationis Christi sermonem ad perfectionem feramur, non rursum iacientes fundamentum paenitentiae ab operibus mortuis et fidei ad Deum,
HEB|6|2|baptismatum doctrinae, impositionis quoque manuum, ac resurrectionis mortuorum et iudicii aeterni.
HEB|6|3|Et hoc faciemus, si quidem permiserit Deus.
HEB|6|4|Impossibile est enim eos, qui semel sunt illuminati, gustaverunt etiam donum caeleste et participes sunt facti Spiritus Sancti
HEB|6|5|et bonum gustaverunt Dei verbum virtutesque saeculi venturi
HEB|6|6|et prolapsi sunt, rursus renovari ad paenitentiam, rursum crucifigentes sibimetipsis Filium Dei et ostentui habentes.
HEB|6|7|Terra enim saepe venientem super se bibens imbrem et generans herbam opportunam illis, propter quos et colitur, accipit benedictionem a Deo;
HEB|6|8|proferens autem spinas ac tribulos reproba est et maledicto proxima, cuius finis in combustionem.
HEB|6|9|Confidimus autem de vobis, dilectissimi, meliora et viciniora saluti, tametsi ita loquimur;
HEB|6|10|non enim iniustus Deus, ut obliviscatur operis vestri et dilectionis, quam ostendistis nomini ipsius, qui ministrastis sanctis et ministratis.
HEB|6|11|Cupimus autem unumquemque vestrum eandem ostentare sollicitudinem ad expletionem spei usque in finem,
HEB|6|12|ut non segnes efficiamini, verum imitatores eorum, qui fide et patientia hereditant promissiones.
HEB|6|13|Abrahae namque promittens Deus, quoniam neminem habuit, per quem iuraret maiorem, iuravit per semetipsum
HEB|6|14|dicens: " Utique benedicens benedicam te et multiplicans multiplicabo te ";
HEB|6|15|et sic longanimiter ferens adeptus est repromissionem.
HEB|6|16|Homines enim per maiorem sui iurant, et omnis controversiae eorum finis ad confirmationem est iuramentum;
HEB|6|17|in quo abundantius volens Deus ostendere pollicitationis heredibus immobilitatem consilii sui, se interposuit iure iurando,
HEB|6|18|ut per duas res immobiles, in quibus impossibile est mentiri Deum, fortissimum solacium habeamus, qui confugimus ad tenendam propositam spem;
HEB|6|19|quam sicut ancoram habemus animae, tutam ac firmam et incedentem usque in interiora velaminis,
HEB|6|20|ubi praecursor pro nobis introivit Iesus, secundum ordinem Melchisedech pontifex factus in aeternum.
HEB|7|1|Hic enim Melchisedech, rex Salem, sacerdos Dei summi, qui ob viavit Abrahae regresso a caede regum et benedixit ei,
HEB|7|2|cui et decimam omnium divisit Abraham, primum quidem, qui interpretatur rex iustitiae, deinde autem et rex Salem, quod est rex Pacis,
HEB|7|3|sine patre, sine matre, sine genealogia, neque initium dierum neque finem vitae habens, assimilatus autem Filio Dei, manet sacerdos in perpetuum.
HEB|7|4|Intuemini autem quantus sit hic, cui et decimam dedit de praecipuis Abraham patriarcha.
HEB|7|5|Et illi quidem, qui de filiis Levi sacerdotium accipiunt, mandatum habent decimas sumere a populo secundum legem, id est a fratribus suis, quamquam et ipsi exierunt de lumbis Abrahae;
HEB|7|6|hic autem, cuius generatio non annumeratur in eis, decimam sumpsit ab Abraham et eum, qui habebat repromissiones, benedixit.
HEB|7|7|Sine ulla autem contradictione, quod minus est, a meliore benedicitur.
HEB|7|8|Et hic quidem decimas morientes homines sumunt; ibi autem testimonium accipiens quia vivit.
HEB|7|9|Et, ut ita dictum sit, per Abraham et Levi, qui decimas accipit, decimatus est;
HEB|7|10|adhuc enim in lumbis patris erat, quando obviavit ei Melchisedech.
HEB|7|11|Si ergo consummatio per sacerdotium leviticum erat, populus enim sub ipso legem accepit, quid adhuc necessarium secundum ordinem Melchisedech alium surgere sacerdotem et non secundum ordinem Aaron dici?
HEB|7|12|Translato enim sacerdotio, necesse est, ut et legis translatio fiat.
HEB|7|13|De quo enim haec dicuntur, ex alia tribu est, ex qua nullus altari praesto fuit;
HEB|7|14|manifestum enim quod ex Iuda ortus sit Dominus noster, in quam tribum nihil de sacerdotibus Moyses locutus est.
HEB|7|15|Et amplius adhuc manifestum est, si secundum similitudinem Melchisedech exsurgit alius sacerdos,
HEB|7|16|qui non secundum legem mandati carnalis factus est sed secundum virtutem vitae insolubilis,
HEB|7|17|testimonium enim accipit: Tu es sacerdos in aeternum secundum ordinem Melchisedech ".
HEB|7|18|Reprobatio quidem fit praecedentis mandati propter infirmitatem eius et inutilitatem,
HEB|7|19|nihil enim ad perfectum adduxit lex; introductio vero melioris spei, per quam proximamus ad Deum.
HEB|7|20|Et quantum non est sine iure iurando; illi quidem sine iure iurando sacerdotes facti sunt,
HEB|7|21|hic autem cum iure iurando per eum, qui dicit ad illum: Iuravit Dominus et non paenitebit eum: Tu es sacerdos in aeternum ",
HEB|7|22|in tantum et melioris testamenti sponsor factus est Iesus.
HEB|7|23|Et illi quidem plures facti sunt sacerdotes, idcirco quod morte prohibebantur permanere;
HEB|7|24|hic autem eo quod manet in aeternum, intransgressibile habet sacerdotium;
HEB|7|25|unde et salvare in perpetuum potest accedentes per semetipsum ad Deum, semper vivens ad interpellandum pro eis.
HEB|7|26|Talis enim et decebat ut nobis esset pontifex, sanctus, innocens, impollutus, segregatus a peccatoribus et excelsior caelis factus;
HEB|7|27|qui non habet necessitatem cotidie, quemadmodum pontifices, prius pro suis delictis hostias offerre, deinde pro populi; hoc enim fecit semel semetipsum offerendo.
HEB|7|28|Lex enim homines constituit pontifices infirmitatem habentes; sermo autem iuris iurandi, quod post legem est, Filium in aeternum consummatum.
HEB|8|1|Caput autem super ea, quae dicuntur: talem habemus ponti ficem, qui consedit in dextera throni Maiestatis in caelis,
HEB|8|2|sanctorum minister et tabernaculi veri, quod fixit Dominus, non homo.
HEB|8|3|Omnis enim pontifex ad offerenda munera et hostias constituitur; unde necesse erat et hunc habere aliquid, quod offerret.
HEB|8|4|Si ergo esset super terram, nec esset sacerdos, cum sint qui offerant secundum legem munera;
HEB|8|5|qui figurae et umbrae deserviunt caelestium, sicut responsum est Moysi, cum consummaturus esset tabernaculum: " Vide enim, inquit, omnia facies secundum exemplar, quod tibi ostensum est in monte ".
HEB|8|6|Nunc autem differentius sortitus est ministerium, quanto et melioris testamenti mediator est, quod in melioribus repromissionibus sancitum est.
HEB|8|7|Nam si illud prius culpa vacasset, non secundi locus inquireretur;
HEB|8|8|vituperans enim eos dicit: " Ecce dies veniunt, dicit Dominus, et consummabo super domum Israel et super domum Iudae testamentum novum;
HEB|8|9|non secundum testamentum, quod feci patribus eorum in die, qua apprehendi manum illorum, ut educerem illos de terra Aegypti; quoniam ipsi non permanserunt in testamento meo, et ego neglexi eos, dicit Dominus.
HEB|8|10|Quia hoc est testamentum, quod testabor domui Israel post dies illos, dicit Dominus, dando leges meas in mentem eorum, et in corde eorum superscribam eas; et ero eis in Deum, et ipsi erunt mihi in populum.
HEB|8|11|Et non docebit unusquisque civem suum, et unusquisque fratrem suum dicens: "Cognosce Dominum"; quoniam omnes scient me, a minore usque ad maiorem eorum,
HEB|8|12|quia propitius ero iniquitatibus eorum et peccatorum illorum iam non memorabor ".
HEB|8|13|Dicendo " novum " veteravit prius; quod autem antiquatur et senescit, prope interitum est.
HEB|9|1|Habuit ergo et prius praecepta cultus et Sanctum huius saeculi.
HEB|9|2|Tabernaculum enim praeparatum est primum, in quo inerat candelabrum et mensa et propositio panum, quod dicitur Sancta;
HEB|9|3|post secundum autem velamentum, tabernaculum, quod dicitur Sancta Sanctorum,
HEB|9|4|aureum habens turibulum et arcam testamenti circumtectam ex omni parte auro, in qua urna aurea habens manna et virga Aaron, quae fronduerat, et tabulae testamenti,
HEB|9|5|superque eam cherubim gloriae obumbrantia propitiatorium; de quibus non est modo dicendum per singula.
HEB|9|6|His vero ita praeparatis, in prius quidem tabernaculum semper intrant sacerdotes sacrorum officia consummantes;
HEB|9|7|in secundum autem semel in anno solus pontifex, non sine sanguine, quem offert pro suis et populi ignorantiis;
HEB|9|8|hoc significante Spiritu Sancto, nondum propalatam esse sanctorum viam, adhuc priore tabernaculo habente statum;
HEB|9|9|quae parabola est temporis instantis, iuxta quam munera et hostiae offeruntur, quae non possunt iuxta conscientiam perfectum facere servientem,
HEB|9|10|solummodo in cibis et in potibus et variis baptismis, quae sunt praecepta carnis usque ad tempus correctionis imposita.
HEB|9|11|Christus autem cum advenit pontifex futurorum bonorum, per amplius et perfectius tabernaculum, non manufactum, id est non huius creationis,
HEB|9|12|neque per sanguinem hircorum et vitulorum sed per proprium sanguinem introivit semel in Sancta, aeterna redemptione inventa.
HEB|9|13|Si enim sanguis hircorum et taurorum et cinis vitulae aspersus inquinatos sanctificat ad emundationem carnis,
HEB|9|14|quanto magis sanguis Christi, qui per Spiritum aeternum semetipsum obtulit immaculatum Deo, emundabit conscientiam nostram ab operibus mortuis ad serviendum Deo viventi.
HEB|9|15|Et ideo novi testamenti mediator est, ut, morte intercedente in redemptionem earum praevaricationum, quae erant sub priore testamento, repromissionem accipiant, qui vocati sunt aeternae hereditatis.
HEB|9|16|Ubi enim testamentum, mors necesse est afferatur testatoris;
HEB|9|17|testamentum autem in mortuis est confirmatum, nondum enim valet, dum vivit, qui testatus est.
HEB|9|18|Unde ne prius quidem sine sanguine dedicatum est;
HEB|9|19|enuntiato enim omni mandato secundum legem a Moyse universo populo, accipiens sanguinem vitulorum et hircorum cum aqua et lana coccinea et hyssopo, ipsum librum et omnem populum aspersit
HEB|9|20|dicens: " Hic sanguis testamenti, quod mandavit ad vos Deus ";
HEB|9|21|etiam tabernaculum et omnia vasa ministerii sanguine similiter aspersit.
HEB|9|22|Et omnia paene in sanguine mundantur secundum legem, et sine sanguinis effusione non fit remissio.
HEB|9|23|Necesse erat ergo figuras quidem caelestium his mundari, ipsa autem caelestia melioribus hostiis quam istis.
HEB|9|24|Non enim in manufacta Sancta Christus introivit, quae sunt similitudo verorum, sed in ipsum caelum, ut appareat nunc vultui Dei pro nobis;
HEB|9|25|neque ut saepe offerat semetipsum, quemadmodum pontifex intrat in Sancta per singulos annos in sanguine alieno.
HEB|9|26|Alioquin oportebat eum frequenter pati ab origine mundi; nunc autem semel in consummatione saeculorum ad destitutionem peccati per sacrificium sui manifestatus est.
HEB|9|27|Et quemadmodum statutum est hominibus semel mori, post hoc autem iudicium,
HEB|9|28|sic et Christus, semel oblatus ad multorum auferenda peccata, secundo sine peccato apparebit exspectantibus se in salutem.
HEB|10|1|Umbram enim habens lex bonorum futurorum, non ip sam imaginem rerum, per singulos annos iisdem ipsis hostiis, quas offerunt indesinenter, numquam potest accedentes perfectos facere.
HEB|10|2|Alioquin nonne cessassent offerri, ideo quod nullam haberent ultra conscientiam peccatorum cultores semel mundati?
HEB|10|3|Sed in ipsis commemoratio peccatorum per singulos annos fit.
HEB|10|4|Impossibile enim est sanguinem taurorum et hircorum auferre peccata.
HEB|10|5|Ideo ingrediens mundum dicit: Hostiam et oblationem noluisti,corpus autem aptasti mihi;
HEB|10|6|holocautomata et sacrificia pro peccatonon tibi placuerunt.
HEB|10|7|Tunc dixi: Ecce venio,in capitulo libri scriptum est de me,ut faciam, Deus, voluntatem tuam ".
HEB|10|8|Superius dicens: " Hostias et oblationes et holocautomata et sacrificia pro peccato noluisti, nec placuerunt tibi ", quae secundum legem offeruntur,
HEB|10|9|tunc dixit: " Ecce venio, ut faciam voluntatem tuam ". Aufert primum, ut secundum statuat;
HEB|10|10|in qua voluntate sanctificati sumus per oblationem corporis Christi Iesu in semel.
HEB|10|11|Et omnis quidem sacerdos stat cotidie ministrans et easdem saepe offerens hostias, quae numquam possunt auferre peccata.
HEB|10|12|Hic autem, una pro peccatis oblata hostia, in sempiternum consedit in dextera Dei,
HEB|10|13|de cetero exspectans, donec ponantur inimici eius scabellum pedum eius;
HEB|10|14|una enim oblatione consummavit in sempiternum eos, qui sanctificantur.
HEB|10|15|Testificatur autem nobis et Spiritus Sanctus; postquam enim dixit:
HEB|10|16|" Hoc est testamentum, quod testabor ad illos post dies illos, dicit Dominus, dando leges meas in cordibus eorum, et in mente eorum superscribam eas;
HEB|10|17|et peccatorum eorum et iniquitatum eorum iam non recordabor amplius ".
HEB|10|18|Ubi autem horum remissio, iam non oblatio pro peccato.
HEB|10|19|Habentes itaque, fratres, fiduciam in introitum Sanctorum in sanguine Iesu,
HEB|10|20|quam initiavit nobis viam novam et viventem per velamen, id est carnem suam,
HEB|10|21|et sacerdotem magnum super domum Dei,
HEB|10|22|accedamus cum vero corde in plenitudine fidei, aspersi corda a conscientia mala et abluti corpus aqua munda;
HEB|10|23|teneamus spei confessionem indeclinabilem, fidelis enim est, qui repromisit;
HEB|10|24|et consideremus invicem in provocationem caritatis et bonorum operum,
HEB|10|25|non deserentes congregationem nostram, sicut est consuetudinis quibusdam, sed exhortantes, et tanto magis quanto videtis appropinquantem diem.
HEB|10|26|Voluntarie enim peccantibus nobis, post acceptam notitiam veritatis, iam non relinquitur pro peccatis hostia,
HEB|10|27|terribilis autem quaedam exspectatio iudicii, et ignis aemulatio, quae consumptura est adversarios.
HEB|10|28|Irritam quis faciens legem Moysis, sine ulla miseratione duobus vel tribus testibus moritur;
HEB|10|29|quanto deteriora putatis merebitur supplicia, qui Filium Dei conculcaverit et sanguinem testamenti communem duxerit, in quo sanctificatus est, et Spiritui gratiae contumeliam fecerit?
HEB|10|30|Scimus enim eum, qui dixit: " Mihi vindicta, ego retribuam "; et iterum: " Iudicabit Dominus populum suum ".
HEB|10|31|Horrendum est incidere in manus Dei viventis.
HEB|10|32|Rememoramini autem pristinos dies, in quibus illuminati magnum certamen sustinuistis passionum,
HEB|10|33|in altero quidem opprobriis et tribulationibus spectaculum facti, in altero autem socii taliter conversantium effecti;
HEB|10|34|nam et vinctis compassi estis et rapinam bonorum vestrorum cum gaudio suscepistis, cognoscentes vos habere meliorem substantiam et manentem.
HEB|10|35|Nolite itaque abicere confidentiam vestram, quae magnam habet remunerationem;
HEB|10|36|patientia enim vobis necessaria est, ut voluntatem Dei facientes reportetis promissionem.
HEB|10|37|Adhuc enim modicum quantulum,qui venturus est, veniet et non tardabit.
HEB|10|38|Iustus autem meus ex fide vivet;quod si subtraxerit se,non sibi complacet in eo anima mea.
HEB|10|39|Nos autem non sumus subtractionis in perditionem, sed fidei in acquisitionem animae.
HEB|11|1|Est autem fides sperando rum substantia, rerum argu mentum non apparentium.
HEB|11|2|In hac enim testimonium consecuti sunt seniores.
HEB|11|3|Fide intellegimus aptata esse saecula verbo Dei, ut ex invisibilibus visibilia facta sint.
HEB|11|4|Fide ampliorem hostiam Abel quam Cain obtulit Deo, per quam testimonium consecutus est esse iustus, testimonium perhibente muneribus eius Deo; et per illam defunctus adhuc loquitur.
HEB|11|5|Fide Henoch translatus est, ne videret mortem, et non inveniebatur, quia transtulit illum Deus; ante translationem enim testimonium accepit placuisse Deo.
HEB|11|6|Sine fide autem impossibile placere; credere enim oportet accedentem ad Deum quia est et inquirentibus se remunerator fit.
HEB|11|7|Fide Noe, responso accepto de his, quae adhuc non videbantur, reveritus aptavit arcam in salutem domus suae; per quam damnavit mundum, et iustitiae, quae secundum fidem est, heres est institutus.
HEB|11|8|Fide vocatus Abraham oboedivit in locum exire, quem accepturus erat in hereditatem; et exivit nesciens quo iret.
HEB|11|9|Fide peregrinatus est in terra promissionis tamquam in aliena, in casulis habitando cum Isaac et Iacob, coheredibus promissionis eiusdem;
HEB|11|10|exspectabat enim fundamenta habentem civitatem, cuius artifex et conditor Deus.
HEB|11|11|Fide - et ipsa Sara sterilis - virtutem in conceptionem seminis accepit etiam praeter tempus aetatis, quoniam fidelem credidit esse, qui promiserat;
HEB|11|12|propter quod et ab uno orti sunt, et hoc emortuo, tamquam sidera caeli in multitudine, et sicut arena, quae est ad oram maris, innumerabilis.
HEB|11|13|Iuxta fidem defuncti sunt omnes isti, non acceptis promissionibus, sed a longe eas aspicientes et salutantes, et confitentes quia peregrini et hospites sunt supra terram;
HEB|11|14|qui enim haec dicunt, significant se patriam inquirere.
HEB|11|15|Et si quidem illius meminissent, de qua exierant, habebant utique tempus revertendi;
HEB|11|16|nunc autem meliorem appetunt, id est caelestem. Ideo non confunditur Deus vocari Deus eorum, paravit enim illis civitatem.
HEB|11|17|Fide obtulit Abraham Isaac, cum tentaretur; et unigenitum offerebat ille, qui susceperat promissiones,
HEB|11|18|ad quem dictum erat: " In Isaac vocabitur tibi semen ",
HEB|11|19|arbitratus quia et a mortuis suscitare potens est Deus; unde eum et in parabola reportavit.
HEB|11|20|Fide et de futuris benedixit Isaac Iacob et Esau.
HEB|11|21|Fide Iacob moriens singulis filiorum Ioseph benedixit et adoravit super fastigium virgae suae.
HEB|11|22|Fide Ioseph moriens de profectione filiorum Israel memoratus est et de ossibus suis mandavit.
HEB|11|23|Fide Moyses natus occultatus est mensibus tribus a parentibus suis, eo quod vidissent formosum infantem et non timuerunt regis edictum.
HEB|11|24|Fide Moyses grandis factus negavit se dici filium filiae pharaonis,
HEB|11|25|magis eligens affligi cum populo Dei quam temporalem peccati habere iucunditatem,
HEB|11|26|maiores divitias aestimans thesauris Aegypti improperium Christi; aspiciebat enim in remunerationem.
HEB|11|27|Fide reliquit Aegyptum non veritus animositatem regis, invisibilem enim tamquam videns sustinuit.
HEB|11|28|Fide celebravit Pascha et sanguinis effusionem, ne, qui vastabat primogenita, tangeret ea.
HEB|11|29|Fide transierunt mare Rubrum tamquam per aridam terram, quod experti Aegyptii devorati sunt.
HEB|11|30|Fide muri Iericho ruerunt circuiti diebus septem.
HEB|11|31|Fide Rahab meretrix non periit cum incredulis, quia exceperat exploratores cum pace.
HEB|11|32|Et quid adhuc dicam? Deficiet enim me tempus enarrantem de Gedeon, Barac, Samson, Iephte, David et Samuel atque prophetis,
HEB|11|33|qui per fidem devicerunt regna, operati sunt iustitiam, adepti sunt repromissiones, obturaverunt ora leonum,
HEB|11|34|exstinxerunt impetum ignis, effugerunt aciem gladii, convaluerunt de infirmitate, fortes facti sunt in bello, castra verterunt exterorum;
HEB|11|35|acceperunt mulieres de resurrectione mortuos suos; alii autem distenti sunt, non suscipientes redemptionem, ut meliorem invenirent resurrectionem;
HEB|11|36|alii vero ludibria et verbera experti sunt, insuper et vincula et carcerem;
HEB|11|37|lapidati sunt, secti sunt, in occisione gladii mortui sunt, circumierunt in melotis, in pellibus caprinis, egentes, angustiati, afflicti,
HEB|11|38|quibus dignus non erat mundus, in solitudinibus errantes et montibus et speluncis et in cavernis terrae.
HEB|11|39|Et hi omnes testimonium per fidem consecuti non reportaverunt promissionem,
HEB|11|40|Deo pro nobis melius aliquid providente, ut ne sine nobis consummarentur.
HEB|12|1|Ideoque et nos tantam ha bentes circumpositam nobis nubem testium, deponentes omne pondus et circumstans nos peccatum, per patientiam curramus propositum nobis certamen,
HEB|12|2|aspicientes in ducem fidei et consummatorem Iesum, qui pro gaudio sibi proposito sustinuit crucem, confusione contempta, atque in dextera throni Dei sedet.
HEB|12|3|Recogitate enim eum, qui talem sustinuit a peccatoribus adversum semetipsum contradictionem, ut ne fatigemini animis vestris deficientes.
HEB|12|4|Nondum usque ad sanguinem restitistis adversus peccatum repugnantes;
HEB|12|5|et obliti estis exhortationis, quae vobis tamquam filiis loquitur: Fili mi, noli neglegere disciplinam Dominineque deficias, dum ab eo argueris:
HEB|12|6|quem enim diligit, Dominus castigat,flagellat autem omnem filium, quem recipit ".
HEB|12|7|Ad disciplinam suffertis; tamquam filios vos tractat Deus. Quis enim filius, quem non corripit pater?
HEB|12|8|Quod si extra disciplinam estis, cuius participes facti sunt omnes, ergo adulterini et non filii estis!
HEB|12|9|Deinde patres quidem carnis nostrae habebamus eruditores et reverebamur; non multo magis obtemperabimus Patri spirituum et vivemus?
HEB|12|10|Et illi quidem ad tempus paucorum dierum, secundum quod videbatur illis, castigabant; hic autem ad id, quod utile est ad participandam sanctitatem eius.
HEB|12|11|Omnis autem disciplina in praesenti quidem videtur non esse gaudii sed maeroris; postea autem fructum pacificum exercitatis per eam reddit iustitiae.
HEB|12|12|Propter quod remissas manus et soluta genua erigite
HEB|12|13|et gressus rectos facite pedibus vestris, ut, quod claudum est, non extorqueatur, magis autem sanetur.
HEB|12|14|Pacem sectamini cum omnibus et sanctificationem, sine qua nemo videbit Dominum,
HEB|12|15|providentes, ne quis desit gratiae Dei, ne qua radix amaritudinis sursum germinans perturbet, et per illam inquinentur multi;
HEB|12|16|ne quis fornicator aut profanus ut Esau, qui propter unam escam vendidit primogenita sua.
HEB|12|17|Scitis enim quoniam et postea cupiens hereditare benedictionem reprobatus est; non enim invenit paenitentiae locum, quamquam cum lacrimis inquisisset eam.
HEB|12|18|Non enim accessistis ad tractabilem et ardentem ignem et turbinem et caliginem et procellam
HEB|12|19|et tubae sonum et vocem verborum, quam qui audierunt, recusaverunt, ne ultra eis fieret verbum;
HEB|12|20|non enim portabant mandatum: " Et si bestia tetigerit montem, lapidabitur";
HEB|12|21|et ita terribile erat, quod videbatur, Moyses dixit: " Exterritus sum et tremebundus ".
HEB|12|22|Sed accessistis ad Sion montem et civitatem Dei viventis, Ierusalem caelestem, et multa milia angelorum, frequentiam
HEB|12|23|et ecclesiam primogenitorum, qui conscripti sunt in caelis, et iudicem Deum omnium et spiritus iustorum, qui consummati sunt,
HEB|12|24|et testamenti novi mediatorem Iesum et sanguinem aspersionis, melius loquentem quam Abel.
HEB|12|25|Videte, ne recusetis loquentem; si enim illi non effugerunt recusantes eum, qui super terram loquebatur, multo magis nos, qui de caelis loquentem avertimus;
HEB|12|26|cuius vox movit terram tunc, modo autem pronuntiavit dicens: " Adhuc semel ego movebo non solum terram sed et caelum ".
HEB|12|27|Hoc autem " adhuc semel " declarat mobilium translationem tamquam factorum, ut maneant ea, quae sunt immobilia.
HEB|12|28|Itaque, regnum immobile suscipientes, habeamus gratiam, per quam serviamus placentes Deo cum reverentia et metu;
HEB|12|29|etenim Deus noster ignis consumens est.
HEB|13|1|Caritas fraternitatis maneat.
HEB|13|2|Hospitalitatem nolite obli visci; per hanc enim quidam nescientes hospitio receperunt angelos.
HEB|13|3|Mementote vinctorum tamquam simul vincti, laborantium tamquam et ipsi in corpore morantes.
HEB|13|4|Honorabile conubium in omnibus, et torus immaculatus; fornicatores enim et adulteros iudicabit Deus.
HEB|13|5|Sint mores sine avaritia; contenti praesentibus. Ipse enim dixit: " Non te deseram neque derelinquam ",
HEB|13|6|ita ut confidenter dicamus: Dominus mihi adiutor est, non timebo; quid faciet mihi homo? ".
HEB|13|7|Mementote praepositorum vestrorum, qui vobis locuti sunt verbum Dei; quorum intuentes exitum conversationis, imitamini fidem.
HEB|13|8|Iesus Christus heri et hodie idem, et in saecula!
HEB|13|9|Doctrinis variis et peregrinis nolite abduci; optimum enim est gratia stabiliri cor, non escis, quae non profuerunt ambulantibus in eis.
HEB|13|10|Habemus altare, de quo edere non habent potestatem, qui tabernaculo deserviunt.
HEB|13|11|Quorum enim animalium infertur sanguis pro peccato in Sancta per pontificem, horum corpora cremantur extra castra.
HEB|13|12|Propter quod et Iesus, ut sanctificaret per suum sanguinem populum, extra portam passus est.
HEB|13|13|Exeamus igitur ad eum extra castra, improperium eius portantes;
HEB|13|14|non enim habemus hic manentem civitatem, sed futuram inquirimus.
HEB|13|15|Per ipsum ergo offeramus hostiam laudis semper Deo, id est fructum labiorum confitentium nomini eius.
HEB|13|16|Beneficientiae autem et communionis nolite oblivisci; talibus enim hostiis oblectatur Deus.
HEB|13|17|Oboedite praepositis vestris et subiacete eis; ipsi enim pervigilant pro animabus vestris quasi rationem reddituri, ut cum gaudio hoc faciant et non gementes; hoc enim non expedit vobis.
HEB|13|18|Orate pro nobis; confidimus enim quia bonam conscientiam habemus, in omnibus bene volentes conversari.
HEB|13|19|Amplius autem deprecor vos hoc facere, ut quo celerius restituar vobis.
HEB|13|20|Deus autem pacis, qui eduxit de mortuis pastorem magnum ovium in sanguine testamenti aeterni, Dominum nostrum Iesum,
HEB|13|21|aptet vos in omni bono, ut faciatis voluntatem eius, faciens in nobis, quod placeat coram se per Iesum Christum, cui gloria in saecula saeculorum. Amen.
HEB|13|22|Rogo autem vos, fratres, sufferte sermonem exhortationis; etenim perpaucis scripsi vobis.
HEB|13|23|Cognoscite fratrem nostrum Timotheum dimissum esse; cum quo, si celerius venerit, videbo vos.
HEB|13|24|Salutate omnes praepositos vestros et omnes sanctos. Salutant vos, qui de Italia sunt.
HEB|13|25|Gratia cum omnibus vobis.
