1COR|1|1|Павло, волею Божою покликаний за апостола Ісуса Христа, і брат Состен,
1COR|1|2|Божій Церкві, що в Коринті, посвяченим у Христі Ісусі, покликаним святим, зо всіма, що на всякому місті прикликають Ім'я Господа нашого Ісуса Христа, їхнього і нашого,
1COR|1|3|благодать вам і мир від Бога Отця нашого й Господа Ісуса Христа!
1COR|1|4|Я завжди дякую моєму Богові за вас, через Божу благодать, що була вам дана в Христі Ісусі,
1COR|1|5|бо ви всім збагатилися в Ньому, словом усяким і всяким знанням,
1COR|1|6|бо свідоцтво Христове між вами утвердилось,
1COR|1|7|так що не маєте недостачі в жаднім дарі благодаті ви, що очікуєте з'явлення Господа нашого Ісуса Христа.
1COR|1|8|Він вас утвердить до кінця неповинними бути дня Господа нашого Ісуса Христа!
1COR|1|9|Вірний Бог, що ви через Нього покликані до спільноти Сина Його Ісуса Христа, Господа нашого.
1COR|1|10|Тож благаю вас, браття, Ім'ям Господа нашого Ісуса Христа, щоб ви всі говорили те саме, і щоб не було поміж вами поділення, але щоб були ви поєднані в однім розумінні та в думці одній!
1COR|1|11|Бо стало відомо мені про вас, мої браття, від Хлоїних, що між вами суперечки.
1COR|1|12|А кажу я про те, що з вас кожен говорить: я ж Павлів, а я Аполлосів, а я Кифин, а я Христів.
1COR|1|13|Чи ж Христос поділився? Чи ж Павло був розп'ятий за вас? Чи в Павлове ім'я ви христились?
1COR|1|14|Дякую Богові, що я ані одного з вас не христив, окрім Кріспа та Гая,
1COR|1|15|щоб ніхто не сказав, ніби я охристив був у ймення своє.
1COR|1|16|Охристив же був я й дім Степанів; більш не знаю, чи христив кого іншого я.
1COR|1|17|Бо Христос не послав мене, щоб христити, а звіщати Євангелію, і то не в мудрості слова, щоб безсилим не став хрест Христа.
1COR|1|18|Бож слово про хреста тим, що гинуть, то глупота, а для нас, що спасаємось, Сила Божа!
1COR|1|19|Бо написано: Я погублю мудрість премудрих, а розум розумних відкину!
1COR|1|20|Де мудрий? Де книжник? Де дослідувач віку цього? Хіба Бог мудрість світу цього не змінив на глупоту?
1COR|1|21|Через те ж, що світ мудрістю не зрозумів Бога в мудрості Божій, то Богові вгодно було спасти віруючих через дурість проповіді.
1COR|1|22|Бо й юдеї жадають ознак, і греки пошукують мудрости,
1COR|1|23|а ми проповідуємо Христа розп'ятого, для юдеїв згіршення, а для греків безумство,
1COR|1|24|а для самих покликаних юдеїв та греків Христа, Божу силу та Божую мудрість!
1COR|1|25|Бо Боже й немудре розумніше воно від людей, а Боже немічне сильніше воно від людей!
1COR|1|26|Дивіться бо, браття, на ваших покликаних, що небагато-хто мудрі за тілом, небагато-хто сильні, небагато-хто шляхетні.
1COR|1|27|Але Бог вибрав немудре світу, щоб засоромити мудрих, і немічне світу Бог вибрав, щоб засоромити сильне,
1COR|1|28|і простих світу, і погорджених, і незначних вибрав Бог, щоб значне знівечити,
1COR|1|29|так щоб не хвалилося перед Богом жадне тіло.
1COR|1|30|А з Нього ви в Христі Ісусі, що став нам мудрістю від Бога, праведністю ж, і освяченням, і відкупленням,
1COR|1|31|щоб було, як написано: Хто хвалиться, нехай хвалиться Господом!
1COR|2|1|А я, як прийшов до вас, браття, не прийшов вам звіщати про Боже свідоцтво з добірною мовою або мудрістю,
1COR|2|2|бо я надумавсь нічого між вами не знати, крім Ісуса Христа, і Того розп'ятого...
1COR|2|3|І я в вас був у немочі, і в страху, і в великім тремтінні.
1COR|2|4|І слово моє й моя проповідь не в словах переконливих людської мудрости, але в доказі духа та сили,
1COR|2|5|щоб була віра ваша не в мудрості людській, але в силі Божій!
1COR|2|6|А ми говоримо про мудрість між досконалими, але мудрість не віку цього, ані володарів цього віку, що гинуть,
1COR|2|7|але ми говоримо Божу мудрість у таємниці, приховану, яку Бог перед віками призначив нам на славу,
1COR|2|8|яку ніхто з володарів цього віку не пізнав; коли б бо пізнали були, то не розп'яли б вони Господа слави!
1COR|2|9|Але, як написано: Чого око не бачило й вухо не чуло, і що на серце людині не впало, те Бог приготував був тим, хто любить Його!
1COR|2|10|А нам Бог відкрив це Своїм Духом, усе бо досліджує Дух, навіть Божі глибини.
1COR|2|11|Хто бо з людей знає речі людські, окрім людського духа, що в нім проживає? Так само не знає ніхто й речей Божих, окрім Духа Божого.
1COR|2|12|А ми прийняли духа не світу, але Духа, що з Бога, щоб знати про речі, від Бога даровані нам,
1COR|2|13|що й говоримо не вивченими словами людської мудрости, але вивченими від Духа Святого, порівнюючи духовне до духовного.
1COR|2|14|А людина тілесна не приймає речей, що від Божого Духа, бо їй це глупота, і вона зрозуміти їх не може, бо вони розуміються тільки духовно.
1COR|2|15|Духовна ж людина судить усе, а її судити не може ніхто.
1COR|2|16|Бо хто розум Господній пізнав, який би його міг навчати? А ми маємо розум Христів!
1COR|3|1|І я, браття, не міг говорити до вас, як до духовних, але як до тілесних, як до немовлят у Христі.
1COR|3|2|Я вас годував молоком, а не твердою їжею, бо ви не могли її їсти, та й тепер ще не можете,
1COR|3|3|бо ви ще тілесні. Бо коли заздрість та суперечки між вами, то чи ж ви не тілесні, і хіба не полюдському робите?
1COR|3|4|Бо коли хто каже: Я ж Павлів, а інший: Я Аполлосів, то чи ж ви не тілесні?
1COR|3|5|Бо хто ж Аполлос? Або хто то Павло? Вони тільки служителі, що ви ввірували через них, і то скільки кому дав Господь.
1COR|3|6|Я посадив, Аполлос поливав, Бог же зростив,
1COR|3|7|тому ані той, хто садить, ані хто поливає, є щось, але Бог, що родить!
1COR|3|8|І хто садить, і хто поливає одне, і кожен одержить свою нагороду за працею своєю!
1COR|3|9|Бо ми співробітники Божі, а ви Боже поле, Божа будівля.
1COR|3|10|Я за благодаттю Божою, що дана мені, як мудрий будівничий, основу поклав, а інший будує на ній; але нехай кожен пильнує, як він будує на ній!
1COR|3|11|Ніхто бо не може покласти іншої основи, окрім покладеної, а вона Ісус Христос.
1COR|3|12|А коли хто на цій основі будує з золота, срібла, дорогоцінного каміння, із дерева, сіна, соломи,
1COR|3|13|то буде виявлене діло кожного, бо виявить день, тому що він огнем об'являється, і огонь діло кожного випробує, яке воно є.
1COR|3|14|І коли чиє діло, яке збудував хто, устоїть, то той нагороду одержить;
1COR|3|15|коли ж діло згорить, той матиме шкоду, та сам він спасеться, але так, як через огонь.
1COR|3|16|Чи не знаєте ви, що ви Божий храм, і Дух Божий у вас пробуває?
1COR|3|17|Як хто нівечить Божого храма, того знівечить Бог, бо храм Божий святий, а храм той то ви!
1COR|3|18|Хай не зводить ніхто сам себе. Як кому з вас здається, що він мудрий в цім віці, нехай стане нерозумним, щоб бути премудрим.
1COR|3|19|Цьогосвітня бо мудрість у Бога глупота, бо написано: Він ловить премудрих у хитрощах їхніх!
1COR|3|20|І знову: Знає Господь думки мудрих, що марнотні вони!
1COR|3|21|Тож нехай ніхто не хвалиться людьми, бо все ваше:
1COR|3|22|чи Павло, чи Аполлос, чи Кифа, чи світ, чи життя, чи смерть, чи теперішнє, чи майбутнє усе ваше,
1COR|3|23|ви ж Христові, а Христос Божий!
1COR|4|1|Нехай кожен нас так уважає, якби служителів Христових і доморядників Божих таємниць;
1COR|4|2|а що ще шукається в доморядниках, щоб кожен був знайдений вірним.
1COR|4|3|А для мене то найменше, щоб судили мене ви чи суд людський, бо я й сам не суджу себе.
1COR|4|4|Я бо проти себе нічого не знаю, але цим не виправдуюсь; Той же, Хто судить мене, то Господь.
1COR|4|5|Тому не судіть передчасно нічого, аж поки не прийде Господь, що й висвітлить таємниці темряви та виявить задуми сердець, і тоді кожному буде похвала від Бога.
1COR|4|6|Оце ж усе, браття, приклав я до себе й Аполлоса ради вас, щоб від нас ви навчилися думати не більш, як написано, щоб ви не чванились один за одним перед іншим.
1COR|4|7|Хто бо тебе вирізняє? Що ти маєш, чого б ти не взяв? А коли ж бо ти взяв, чого чванишся, ніби не взяв?
1COR|4|8|Ви вже нагодовані, ви вже збагатилися, без нас ви царюєте. І коли б то ви стали царювати, щоб і ми царювали з вами!
1COR|4|9|Бо я думаю, що Бог нас, апостолів, поставив за найостанніших, мов на смерть засуджених, бо ми стали дивовищем світові, і Анголам, і людям.
1COR|4|10|Ми нерозумні Христа ради, а ви мудрі в Христі; ми слабі, ви ж міцні; ви славні, а ми безчесні!
1COR|4|11|Ми до цього часу і голодуємо, і прагнемо, і нагі ми, і катовані, і тиняємось,
1COR|4|12|і трудимось, працюючи своїми руками. Коли нас лихословлять, ми благословляємо; як нас переслідують, ми терпимо;
1COR|4|13|як лають, ми молимось; ми стали, як сміття те для світу, аж досі ми всім, як ті викидки!
1COR|4|14|Не пишу це для того, щоб вас осоромити, але остерігаю, як своїх любих дітей.
1COR|4|15|Бо хоч би ви мали десять тисяч наставників у Христі, та отців не багато; а я вас породив у Христі Ісусі через Євангелію...
1COR|4|16|Тож благаю я вас: будьте наслідувачами мене!
1COR|4|17|Для цього послав я до вас Тимофія, що для мене улюблений і вірний син у Господі, він вам нагадає шляхи мої в Христі Ісусі, як навчаю я скрізь у кожній Церкві.
1COR|4|18|Деякі згорділи, так немов би не мав я прийти до вас.
1COR|4|19|Та небавом прийду до вас, як захоче Господь, і пізнаю не слово згорділих, але силу.
1COR|4|20|Бо Царство Боже не в слові, а в силі.
1COR|4|21|Чого хочете? Чи прийти до вас з києм, чи з любов'ю та з духом лагідности?
1COR|5|1|Всюди чути, що між вами перелюб, і то такий перелюб, який і між поганами незнаний, що хтось має за дружину собі дружину батькову...
1COR|5|2|І ви завеличалися, а не засмутились радніш, щоб був вилучений з-поміж вас, хто цей учинок зробив.
1COR|5|3|Отож я, відсутній тілом, та присутній духом, уже розсудив, як присутній між вами: того, хто так учинив це,
1COR|5|4|у Ім'я Господа Ісуса, як зберетеся ви та мій дух, із силою Господа нашого Ісуса,
1COR|5|5|віддати такого сатані на погибіль тіла, щоб дух спасся Господнього дня!
1COR|5|6|Величання ваше не добре. Хіба ви не знаєте, що мала розчина все тісто заквашує?
1COR|5|7|Отож, очистьте стару розчину, щоб стати вам новим тістом, бо ви прісні, бо наша Пасха, Христос, за нас у жертву принесений.
1COR|5|8|Тому святкуймо не в давній розчині, ані в розчині злоби й лукавства, але в опрісноках чистости та правди!
1COR|5|9|Я писав вам у листі не єднатися з перелюбниками,
1COR|5|10|але не взагалі з цьогосвітніми перелюбниками, чи з користолюбцями, чи з хижаками, чи з ідолянами, бо ви мусіли були б відійти від світу.
1COR|5|11|А тепер я писав вам не єднатися з тим, хто зветься братом, та є перелюбник, чи користолюбець, чи ідолянин, чи злоріка, чи п'яниця, чи хижак, із такими навіть не їсти!
1COR|5|12|Бо що ж мені судити й чужих? Чи ви не судите своїх?
1COR|5|13|А чужих судить Бог. Тож вилучіть лукавого з-поміж себе самих!
1COR|6|1|Чи посміє хто з вас, маючи справу до іншого, судитися в неправедних, а не в святих?
1COR|6|2|Хіба ви не знаєте, що святі світ судитимуть? Коли ж будете ви світ судити, то чи ж ви негідні судити незначні справи?
1COR|6|3|Хіба ви не знаєте, що ми будем судити Анголів, а не тільки життєве?
1COR|6|4|А ви, коли маєте суд за життєве, то ставите суддями тих, хто нічого не значить у Церкві.
1COR|6|5|Я на сором це вам говорю. Чи ж між вами немає ні одного мудрого, щоб він міг розсудити між братами своїми?
1COR|6|6|Та брат судиться з братом, і то перед невірними!
1COR|6|7|Тож уже для вас сором зовсім, що суди між собою ви маєте. Чому краще не терпите кривди? Чому краще не маєте шкоди?
1COR|6|8|Але ви самі кривду чините та обдираєте, та ще братів...
1COR|6|9|Хіба ви не знаєте, що неправедні не вспадкують Божого Царства? Не обманюйте себе: ні розпусники, ні ідоляни, ні перелюбники, ні блудодійники, ні мужоложники,
1COR|6|10|ні злодії, ні користолюбці, ні п'яниці, ні злоріки, ні хижаки Царства Божого не вспадкують вони!
1COR|6|11|І такими були дехто з вас, але ви обмились, але освятились, але виправдались Іменем Господа Ісуса Христа й Духом нашого Бога.
1COR|6|12|Усе мені можна, та не все на пожиток. Усе мені можна, але мною ніщо володіти не повинно.
1COR|6|13|Їжа для черева, і черево для їжі, але Бог одне й друге понищить. А тіло не для розпусти, але для Господа, і Господь для тіла.
1COR|6|14|Бог же й Господа воскресив, воскресить Він і нас Своєю силою!
1COR|6|15|Хіба ви не знаєте, що ваші тіла то члени Христові? Отож, узявши члени Христові, зроблю їх членами розпусниці? Зовсім ні!
1COR|6|16|Хіба ви не знаєте, що той, хто злучується з розпусницею, стає одним тілом із нею? Бо каже: Обидва ви будете тілом одним.
1COR|6|17|А хто з Господом злучується, стає одним духом із Ним.
1COR|6|18|Утікайте від розпусти. Усякий бо гріх, що його чинить людина, є поза тілом. А хто чинить розпусту, той грішить проти власного тіла.
1COR|6|19|Хіба ви не знаєте, що ваше тіло то храм Духа Святого, що живе Він у вас, якого від Бога ви маєте, і ви не свої?
1COR|6|20|Бо дорого куплені ви. Отож прославляйте Бога в тілі своєму та в дусі своєму, що Божі вони!
1COR|7|1|А про що ви писали мені, то добре було б чоловікові не дотикатися жінки.
1COR|7|2|Але щоб уникнути розпусти, нехай кожен муж має дружину свою, і кожна жінка хай має свого чоловіка.
1COR|7|3|Нехай віддає чоловік своїй дружині потрібну любов, так же само й чоловікові дружина.
1COR|7|4|Дружина не володіє над тілом своїм, але чоловік; так же само й чоловік не володіє над тілом своїм, але дружина.
1COR|7|5|Не вхиляйтесь одне від одного, хібащо дочасно за згодою, щоб бути в пості та молитві, та й сходьтеся знову докупи, щоб вас сатана не спокушував вашим нестриманням.
1COR|7|6|А це говорю вам як раду, а не як наказа.
1COR|7|7|Бо хочу, щоб усі чоловіки були, як і я; але кожен має від Бога свій дар, один так, інший так.
1COR|7|8|Говорю ж неодруженим і вдовам: добре їм, як вони позостануться так, як і я.
1COR|7|9|Коли ж не втримаються, нехай одружуються, бо краще женитися, ніж розпалятися.
1COR|7|10|А тим, що побрались, наказую не я, а Господь: Нехай не розлучається дружина з своїм чоловіком!
1COR|7|11|А коли ж і розлучиться, хай зостається незаміжня, або з чоловіком своїм хай помириться, і не відпускати чоловікові дружини!
1COR|7|12|Іншим же я говорю, не Господь: коли який брат має дружину невіруючу, і згідна вона жити з ним, нехай він не лишає її.
1COR|7|13|І жінка, як має чоловіка невіруючого, а той згоден жити з нею, нехай не лишає його.
1COR|7|14|Чоловік бо невіруючий освячується в дружині, а дружина невіруюча освячується в чоловікові. А інакше нечисті були б ваші діти, тепер же святі.
1COR|7|15|А як хоче невіруючий розлучитися, хай розлучиться, не неволиться брат чи сестра в такім разі, бо покликав нас Бог до миру.
1COR|7|16|Звідки знаєш ти, дружино, чи не спасеш чоловіка? Або звідки знаєш, чоловіче, чи не спасеш дружини?
1COR|7|17|Нехай тільки так ходить кожен, як кому Бог призначив, як Господь покликав його. І так усім Церквам я наказую.
1COR|7|18|Хто покликаний був в обрізанні, нехай він того не цурається; чи покликаний хто в необрізанні, нехай не обрізується.
1COR|7|19|Обрізання ніщо, і ніщо необрізання, а важливе дотримування Божих заповідей.
1COR|7|20|Нехай кожен лишається в стані такому, в якому покликаний був.
1COR|7|21|Чи покликаний був ти рабом? Не турбуйся про те. Але коли й можеш стати вільним, то використай краще це.
1COR|7|22|Бо покликаний в Господі раб визволенець Господній; так само покликаний і визволенець він раб Христа.
1COR|7|23|Ви дорого куплені, тож не ставайте рабами людей!
1COR|7|24|Браття, кожен із вас, в якім стані покликаний був, хай у тім перед Богом лишається!
1COR|7|25|Про дівчат же не маю наказу Господнього, але даю раду як той, хто одержав від Господа милість буть вірним.
1COR|7|26|Отож за сучасного утиску добрим уважаю я те, що чоловікові добре лишатися так.
1COR|7|27|Ти зв'язаний з дружиною? Не шукай розв'язання. Розв'язався від дружини? Не шукай дружини.
1COR|7|28|А коли ти й оженишся, то не згрішив; і як дівчина заміж піде, вона не згрішить. Та муку тілесну такі будуть мати, а мені шкода вас.
1COR|7|29|А це, браття, кажу я, бо час позосталий короткий, щоб і ті, що мають дружин, були, як ті, що не мають,
1COR|7|30|а хто плаче, як ті, хто не плаче, а хто тішиться, як ті, хто не тішиться; і хто купує, як би не набули,
1COR|7|31|а хто цьогосвітнім користується, як би не користувались, бо минає стан світу цього.
1COR|7|32|А я хочу, щоб ви безклопітні були. Неодружений про речі Господні клопочеться, як догодити Господеві,
1COR|7|33|а одружений про речі життєві клопочеться, як догодити своїй дружині,
1COR|7|34|і він поділений. Незаміжня ж жінка та дівчина про речі Господні клопочеться, щоб бути святою ті тілом, і духом. А заміжня про речі життєві клопочеться, як догодити чоловікові.
1COR|7|35|А це я кажу вам самим на пожиток, а не щоб сильце вам накинути, але щоб пристойно й горливо держались ви Господа.
1COR|7|36|А як думає хто про дівчину свою, що соромно, як вона переросте, і так мала б лишатись, нехай робить, що хоче, не згрішить: нехай заміж виходять.
1COR|7|37|А хто в серці своїм стоїть міцно, не має конечности, владу ж має над своєю волею, і це постановив він у серці своєму берегти свою дівчину, той робить добре.
1COR|7|38|Тому й той, хто віддає свою дівчину заміж, добре робить, а хто не віддає робить краще.
1COR|7|39|Дружина законом прив'язана, поки живе чоловік її; коли ж чоловік її вмре, вона вільна виходити заміж, за кого захоче, аби тільки в Господі.
1COR|7|40|Блаженніша вона, коли так позостанеться за моєю порадою, бо міркую, що й я маю Божого Духа.
1COR|8|1|А щодо ідольських жертов, то ми знаємо, що всі маємо знання. Знання ж надимає, любов же будує!
1COR|8|2|Коли хто думає, ніби щось знає, той нічого не знає ще так, як знати повинно.
1COR|8|3|Коли ж любить хто Бога, той пізнаний Ним.
1COR|8|4|Тож про споживання ідольських жертов ми знаємо, що ідол у світі ніщо, і що іншого Бога нема, окрім Бога Одного.
1COR|8|5|Бо хоч і існують так звані боги чи на небі, чи то на землі, як існує багато богів і багато панів,
1COR|8|6|та для нас один Бог Отець, що з Нього походить усе, ми ж для Нього, і один Господь Ісус Христос, що все сталося Ним, і ми Ним.
1COR|8|7|Та не всі таке мають знання, бо деякі мають призвичаєння до ідола й досі, і їдять, як ідольську жертву, і їхнє сумління, бувши недуже, споганюється.
1COR|8|8|Їжа ж нас до Бога не зближує: бо коли не їмо, то нічого не тратимо, а коли ми їмо, то не набуваєм нічого.
1COR|8|9|Але стережіться, щоб ця ваша воля не стала якось за спотикання слабим!
1COR|8|10|Коли бо хто бачить тебе, маючого знання, як ти в ідольській божниці сидиш за столом, чи ж сумління його, бувши слабе, не буде спонукане їсти ідольські жертви?
1COR|8|11|І через знання твоє згине недужий твій брат, що за нього Христос був умер!
1COR|8|12|Грішачи так проти братів та вражаючи їхнє слабе сумління, ви проти Христа грішите.
1COR|8|13|Ось тому, коли їжа спокушує брата мого, то повік я не їстиму м'яса, щоб не спокусити брата свого!
1COR|9|1|Хіба ж я не вільний? Чи ж я не апостол? Хіба я не бачив Ісуса Христа, Господа нашого? Хіба ви, то не справа моя перед Господом?
1COR|9|2|Коли я не апостол для інших, то для вас я апостол, ви бо печать мого апостольства в Господі.
1COR|9|3|Оце оборона моя перед тими, хто судить мене.
1COR|9|4|Чи ми права не маємо їсти та пити?
1COR|9|5|Чи ми права не маємо водити з собою сестру, дружину, як і інші апостоли, і Господні брати, і Кифа?
1COR|9|6|Хіба я один і Варнава не маємо права, щоб не працювати?
1COR|9|7|Хто коштом своїм коли служить у війську? Або хто виноградника садить, і не їсть з його плоду? Або хто отару пасе, і не їсть молока від отари?
1COR|9|8|Чи я тільки по-людському це говорю? Хіба ж і Закон не говорить цього?
1COR|9|9|Бо в Законі Мойсеєвім писано: Не в'яжи рота волові, що молотить. Хіба за волів Бог турбується?
1COR|9|10|Чи говорить Він зовсім для нас? Для нас, бо написано, що з надією мусить орати орач, а молотник молотити з надією мати частку в своїм сподіванні.
1COR|9|11|Коли ми сіяли вам духовне, чи ж велика то річ, як пожнемо ми ваше тілесне?
1COR|9|12|Як право на вас мають інші, то тим більше ми. Але ми не вжили цього права, та все терпимо, аби перешкоди якої Христовій Євангелії ми не вчинили.
1COR|9|13|Хіба ви не знаєте, що священнослужителі від святині годуються? Що ті, хто служить вівтареві, із вівтаря мають частку?
1COR|9|14|Так і Господь наказав проповідникам Євангелії жити з Євангелії.
1COR|9|15|Але з того нічого не вжив я. А цього не писав я для того, щоб для мене так було. Бо мені краще вмерти, аніж щоб хто знівечив хвалу мою!
1COR|9|16|Бо коли я звіщаю Євангелію, то нема чим хвалитись мені, це бо повинність моя. І горе мені, коли я не звіщаю Євангелії!
1COR|9|17|Тож коли це роблю добровільно, я маю нагороду; коли ж недобровільно, то виконую службу доручену.
1COR|9|18|Яка ж нагорода мені? Та, що, благовістячи, я безкорисливо проповідував Христову Євангелію, не використовуючи особистих прав щодо благовістя.
1COR|9|19|Від усіх бувши вільний, я зробився рабом для всіх, щоб найбільше придбати.
1COR|9|20|Для юдеїв я був, як юдей, щоб юдеїв придбати; для підзаконних був, як підзаконний, хоч сам підзаконним не бувши, щоб придбати підзаконних.
1COR|9|21|Для тих, хто без Закону, я був беззаконний, не бувши беззаконний Богові, а законний Христові, щоб придбати беззаконних.
1COR|9|22|Для слабих, як слабий, щоб придбати слабих. Для всіх я був усе, щоб спасти бодай деяких.
1COR|9|23|А це я роблю для Євангелії, щоб стати її спільником.
1COR|9|24|Хіба ви не знаєте, що ті, хто на перегонах біжить, усі біжать, але нагороду приймає один? Біжіть так, щоб одержали ви!
1COR|9|25|І кожен змагун від усього стримується; вони ж щоб тлінний прийняти вінок, але ми щоб нетлінний.
1COR|9|26|Тож біжу я не так, немов на непевне, борюся не так, немов би повітря б'ючи.
1COR|9|27|Але вмертвляю й неволю я тіло своє, щоб, звіщаючи іншим, не стати самому негідним.
1COR|10|1|Не хочу я, браття, щоб ви не знали, що під хмарою всі отці наші були, і всі перейшли через море,
1COR|10|2|і всі охристилися в хмарі та в морі в Мойсея,
1COR|10|3|і всі їли ту саму поживу духовну,
1COR|10|4|і пили всі той самий духовний напій, бо пили від духовної скелі, що йшла вслід за ними, а та скеля був Христос!
1COR|10|5|Але їх багатьох не вподобав був Бог, бо понищив Він їх у пустині.
1COR|10|6|А це були приклади нам, щоб ми пожадливі на зле не були, як були пожадливі й вони.
1COR|10|7|Не будьте також ідолянами, як деякі з них, як написано: Люди сіли, щоб їсти та пити, і встали, щоб грати.
1COR|10|8|Не станьмо чинити блуду, як деякі з них блудодіяли, і полягло їх одного дня двадцять три тисячі.
1COR|10|9|Ані не випробовуймо Христа, як деякі з них випробовували, та й від зміїв загинули.
1COR|10|10|Ані не нарікайте, як деякі з них нарікали, і загинули від погубителя.
1COR|10|11|Усе це трапилось з ними, як приклади, а написане нам на науку, бо за нашого часу кінець віку прийшов.
1COR|10|12|Тому то, хто думає, ніби стоїть він, нехай стережеться, щоб не впасти!
1COR|10|13|Досягла вас спроба не інша, тільки людська; але вірний Бог, Який не попустить, щоб ви випробовувалися більше, ніж можете, але при спробі й полегшення дасть, щоб знести могли ви її.
1COR|10|14|Тому, мої любі, утікайте від служіння ідолам.
1COR|10|15|Кажу, як розумним; судіть самі, що кажу я.
1COR|10|16|Чаша благословення, яку благословляємо, чи не спільнота то крови Христової? Хліб, який ломимо, чи не спільнота він тіла Христового?
1COR|10|17|Тому що один хліб, тіло одне нас багато, бо ми всі спільники хліба одного.
1COR|10|18|Погляньте на Ізраїля за тілом: чи ж ті, що жертви їдять, не спільники вівтаря?
1COR|10|19|Тож що я кажу? Що ідольська жертва є щось? Чи що ідол є щось?
1COR|10|20|Ні, але те, що в жертву приносять, демонам, а не Богові в жертву приносять. Я ж не хочу, щоб ви спільниками для демонів стали.
1COR|10|21|Бо не можете пити чаші Господньої та чаші демонської; не можете бути спільниками Господнього столу й столу демонського.
1COR|10|22|Чи ми дратуватимем Господа? Хіба ми потужніші за Нього?
1COR|10|23|Усе мені можна, та не все на пожиток. Усе мені можна, та будує не все!
1COR|10|24|Нехай не шукає ніхто свого власного, але кожен для ближнього!
1COR|10|25|Їжте все, що на ятках м'ясних продається, за сумління зовсім не турбуючись,
1COR|10|26|Бо Господня земля, і все, що на ній!
1COR|10|27|Як покличе вас хтось із невіруючих, і ви захочете піти, їжте все, що дадуть вам, за сумління зовсім не турбуючись.
1COR|10|28|Коли ж скаже вам хтось: Це ідольська жертва, не їжте тоді через того, хто сказав, та через сумління!
1COR|10|29|Говорю ж не про власне сумління, але іншого, чого б моя воля судилась сумлінням чужим?
1COR|10|30|Коли я стаю спільником їжі з подякою, чому мене зневажають за те, за що дякую я?
1COR|10|31|Тож, коли ви їсте, чи коли ви п'єте, або коли інше що робите, усе на Божу славу робіть!
1COR|10|32|Не робіть спокуси юдеям та гелленам, та Церкві Божій,
1COR|10|33|як догоджую й я всім у всьому, не шукаючи в тому пожитку свого, але пожитку для багатьох, щоб спаслися вони.
1COR|11|1|Будьте наслідувачами мене, як і я Христа!
1COR|11|2|Похваляю ж вас, браття, що ви все моє пам'ятаєте, і заховуєте так передання, як я вам передав.
1COR|11|3|Хочу ж я, щоб ви знали, що всякому чоловікові голова Христос, а жінці голова чоловік, голова ж Христові Бог.
1COR|11|4|Кожен чоловік, що молиться чи пророкує з головою покритою, осоромлює він свою голову.
1COR|11|5|І кожна жінка, що молиться чи пророкує з головою відкритою, осоромлює тим свою голову, бо це є те саме, як була б вона виголена.
1COR|11|6|Бо коли жінка не покривається, хай стрижеться вона; коли ж жінці сором стригтися чи голитися, нехай покривається!
1COR|11|7|Отож, чоловік покривати голови не повинен, бо він образ і слава Бога, а жінка чоловікові слава.
1COR|11|8|Бо чоловік не походить від жінки, але жінка від чоловіка,
1COR|11|9|не створений бо чоловік ради жінки, але жінка ради чоловіка.
1COR|11|10|Тому жінка повина мати на голові знака влади над нею, ради Анголів.
1COR|11|11|Одначе в Господі ані чоловік без жінки, ані жінка без чоловіка.
1COR|11|12|Бо як жінка від чоловіка, так і чоловік через жінку; а все від Бога.
1COR|11|13|Поміркуйте самі між собою, чи пристойне воно, щоб жінка молилася Богові непокрита?
1COR|11|14|Чи ж природа сама вас не вчить, що коли чоловік запускає волосся, то безчестя для нього?
1COR|11|15|Коли ж жінка косу запускає, це слава для неї, бо замість покривала дана коса їй.
1COR|11|16|Коли ж хто сперечатися хоче, ми такого звичаю не маємо, ані Церкви Божі.
1COR|11|17|Пропонуючи це вам, я не хвалю, що збираєтесь ви не на ліпше, а на гірше.
1COR|11|18|Бо найперше, я чую, що як сходитесь ви на збори, то між вами бувають поділення, у що почасти я й вірю.
1COR|11|19|Бо мусять між вами й поділи бути, щоб відкрились між вами й досвідчені.
1COR|11|20|А далі, коли ви збираєтесь разом, то не на те, щоб їсти Господню Вечерю.
1COR|11|21|Бо кожен спішить з'їсти власну вечерю, і один голодує, а другий впивається.
1COR|11|22|Хіба ж ви не маєте хат, щоб їсти та пити? Чи ви зневажаєте Божу Церкву, і осоромлюєте немаючих? Що маю сказати вам? Чи за це похвалю вас? Не похвалю!
1COR|11|23|Бо прийняв я від Господа, що й вам передав, що Господь Ісус ночі тієї, як виданий був, узяв хліб,
1COR|11|24|подяку віддав, і переломив, і сказав: Прийміть, споживайте, це тіло Моє, що за вас ломається. Це робіть на спомин про Мене!
1COR|11|25|Так само і чашу взяв Він по Вечері й сказав: Ця чаша Новий Заповіт у Моїй крові. Це робіть, коли тільки будете пити, на спомин про Мене!
1COR|11|26|Бо кожного разу, як будете їсти цей хліб та чашу цю пити, смерть Господню звіщаєте, аж доки Він прийде.
1COR|11|27|Тому то, хто їстиме хліб цей чи питиме чашу Господню негідно, буде винний супроти тіла та крови Господньої!
1COR|11|28|Нехай же людина випробовує себе, і так нехай хліб їсть і з чаші хай п'є.
1COR|11|29|Бо хто їсть і п'є негідно, не розважаючи про тіло, той суд собі їсть і п'є!
1COR|11|30|Через це поміж вами багато недужих та хворих, і багато-хто заснули.
1COR|11|31|Бо коли б ми самі судили себе, то засуджені ми не були б.
1COR|11|32|Та засуджені від Господа, караємося, щоб нас не засуджено з світом.
1COR|11|33|Ось тому, мої браття, сходячись на поживу, чекайте один одного.
1COR|11|34|А коли хто голодний, нехай вдома він їсть, щоб не сходилися ви на осуд. А про інше, як прийду, заряджу.
1COR|12|1|А щодо духовних дарів, то не хочу я, браття, щоб не відали ви.
1COR|12|2|Знаєте, що коли ви поганами були, то ходили до німих ідолів, ніби воджено вас.
1COR|12|3|Тому то кажу вам, що ніхто, хто говорить Духом Божим, не скаже: Нехай анатема буде на Ісуса, і не може сказати ніхто: Ісус то Господь, як тільки Духом Святим.
1COR|12|4|Є різниця між дарами милости, Дух же той Самий.
1COR|12|5|Є й різниця між служіннями, та Господь той же Самий.
1COR|12|6|Є різниця й між діями, але Бог той же Самий, що в усіх робить усе.
1COR|12|7|І кожному дається виявлення Духа на користь.
1COR|12|8|Одному бо Духом дається слово мудрости, а другому слово знання тим же Духом,
1COR|12|9|а іншому віра тим же Духом, а іншому дари вздоровлення тим же Духом,
1COR|12|10|а іншому роблення чуд, а іншому пророкування, а іншому розпізнавання духів, а тому різні мови, а іншому вияснення мов.
1COR|12|11|А все оце чинить один і той Самий Дух, уділяючи кожному осібно, як Він хоче.
1COR|12|12|Бо як тіло одне, але має членів багато, усі ж члени тіла, хоч їх багато, то тіло одне, так і Христос.
1COR|12|13|Бо ми всі одним Духом охрищені в тіло одне, чи то юдеї, чи геллени, чи раби, чи то вільні, і всі ми напоєні Духом одним.
1COR|12|14|Бо тіло не є один член, а багато.
1COR|12|15|Коли скаже нога, що я не від тіла, бо я не рука, то хіба через це не від тіла вона?
1COR|12|16|І коли скаже вухо, що я не від тіла, бо я не око, то хіба через це не від тіла воно?
1COR|12|17|Коли б оком було ціле тіло, то де був би слух? А коли б усе слух, то де був би нюх?
1COR|12|18|Та нині Бог розклав члени в тілі, кожного з них, як хотів.
1COR|12|19|Якби всі одним членом були, то де тіло було б?
1COR|12|20|Отож, тепер членів багато, та тіло одне.
1COR|12|21|Бо око не може сказати руці: Ти мені непотрібна; або голова знов ногам: Ви мені непотрібні.
1COR|12|22|Але члени тіла, що здаються слабіші, значно більше потрібні.
1COR|12|23|А тим, що вважаємо їх за зовсім нешановані в тілі, таким честь найбільшу приносимо, і бридкі наші члени отримують пристойність найбільшу,
1COR|12|24|а нашим пристойним того не потрібно. Та Бог змішав тіло, і честь більшу дав нижчому членові,
1COR|12|25|щоб поділення в тілі не було, а щоб члени однаково дбали один про одного.
1COR|12|26|І коли терпить один член, то всі члени з ним терплять; і коли один член пошанований, то всі члени з ним тішаться.
1COR|12|27|І ви тіло Христове, а зосібна ви члени!
1COR|12|28|А інших поставив Бог у Церкві поперше апостолами, подруге пророками, потретє учителями, потім дав сили, також дари вздоровлення, допомоги, управління, різні мови.
1COR|12|29|Чи ж усі апостоли? Чи ж усі пророки? Чи ж усі вчителі? Чи ж усі сили чудодійні?
1COR|12|30|Чи ж усі мають дари вздоровлення? Чи ж мовами всі розмовляють? Чи ж усі виясняють?
1COR|12|31|Тож дбайте ревно про ліпші дари, а я вам покажу путь іще кращу!
1COR|13|1|Коли я говорю мовами людськими й ангольськими, та любови не маю, то став я як мідь та дзвінка або бубон гудячий!
1COR|13|2|І коли маю дара пророкувати, і знаю всі таємниці й усе знання, і коли маю всю віру, щоб навіть гори переставляти, та любови не маю, то я ніщо!
1COR|13|3|І коли я роздам усі маєтки свої, і коли я віддам своє тіло на спалення, та любови не маю, то пожитку не матиму жадного!
1COR|13|4|Любов довготерпить, любов милосердствує, не заздрить, любов не величається, не надимається,
1COR|13|5|не поводиться нечемно, не шукає тільки свого, не рветься до гніву, не думає лихого,
1COR|13|6|не радіє з неправди, але тішиться правдою,
1COR|13|7|усе зносить, вірить у все, сподівається всього, усе терпить!
1COR|13|8|Ніколи любов не перестає! Хоч пророцтва й існують, та припиняться, хоч мови існують, замовкнуть, хоч існує знання, та скасується.
1COR|13|9|Бо ми знаємо частинно, і пророкуємо частинно;
1COR|13|10|коли ж досконале настане, тоді зупиниться те, що частинне.
1COR|13|11|Коли я дитиною був, то я говорив, як дитина, як дитина я думав, розумів, як дитина. Коли ж мужем я став, то відкинув дитяче.
1COR|13|12|Отож, тепер бачимо ми ніби у дзеркалі, у загадці, але потім обличчям в обличчя; тепер розумію частинно, а потім пізнаю, як і пізнаний я.
1COR|13|13|А тепер залишаються віра, надія, любов, оці три. А найбільша між ними любов!
1COR|14|1|Дбайте про любов, і про духовне пильнуйте, а найбільше щоб пророкувати.
1COR|14|2|Як говорить хто чужою мовою, той не людям говорить, а Богові, бо ніхто його не розуміє, і він духом говорить таємне.
1COR|14|3|А хто пророкує, той людям говорить на збудування, і на умовлення, і на розраду.
1COR|14|4|Як говорить хто чужою мовою, той будує тільки самого себе, а хто пророкує, той Церкву будує.
1COR|14|5|Я ж хочу, щоб мовами говорили всі, а ліпше щоб пророкували: більший бо той, хто пророкує, аніж той, хто говорить мовами, хібащо пояснює, щоб будувалася Церква.
1COR|14|6|А тепер, як прийду я до вас, браття, і до вас говорити буду чужою мовою, то який вам пожиток зроблю, коли не поясню вам чи то відкриттям, чи знанням, чи пророцтвом, чи наукою?
1COR|14|7|Бо навіть і речі бездушні, що звук видають, як сопілка чи лютня, коли б не видавали вони різних звуків, як пізнати б тоді, що бринить або грає?
1COR|14|8|Бо коли сурма звук невиразний дає, хто до бою готовитись буде?
1COR|14|9|Так і ви, коли мовою не подасте зрозумілого слова, як пізнати, що кажете? Ви говоритимете на вітер!
1COR|14|10|Як багато, наприклад, різних мов є на світі, і жадна з них не без значення!
1COR|14|11|І коли я не знатиму значення слів, то я буду чужинцем промовцеві, і промовець чужинцем мені.
1COR|14|12|Так і ви, що пильнуєте про духовні дари, дбайте, щоб збагачуватись через них на збудування Церкви!
1COR|14|13|Ось тому, хто говорить чужою мовою, нехай молиться, щоб умів виясняти.
1COR|14|14|Бо коли я молюся чужою мовою, то молиться дух мій, а мій розум без плоду!
1COR|14|15|Ну, то що ж? Буду молитися духом, і буду молитися й розумом, співатиму духом, і співатиму й розумом.
1COR|14|16|Бо коли благословлятимеш духом, то як той, що займає місце простої людини, промовить амінь на подяку твою? Не знає бо він, що ти кажеш.
1COR|14|17|Ти дякуєш добре, але не будується інший.
1COR|14|18|Дякую Богові моєму, розмовляю я мовами більше всіх вас.
1COR|14|19|Але в Церкві волію п'ять слів зрозумілих сказати, щоб і інших навчити, аніж десять тисяч слів чужою мовою!
1COR|14|20|Браття, не будьте дітьми своїм розумом, будьте в лихому дітьми, а в розумі досконалими будьте!
1COR|14|21|У Законі написано: Іншими мовами й іншими устами Я говоритиму людям оцим, та Мене вони й так не послухають, каже Господь.
1COR|14|22|Отож, мови існують на знак не для віруючих, але для невіруючих, а пророцтво для віруючих, а не для невіруючих.
1COR|14|23|А як зійдеться Церква вся разом, і всі говоритимуть чужими мовами, і ввійдуть туди й сторонні чи невіруючі, чи ж не скажуть вони, що біснуєтесь ви?
1COR|14|24|Коли ж усі пророкують, а ввійде якийсь невіруючий чи сторонній, то всі докоряють йому, усі судять його,
1COR|14|25|і так таємниці серця його виявляються, і так він падає ницьма і вклоняється Богові й каже: Бог справді між вами!
1COR|14|26|То що ж, браття? Коли сходитесь ви, то кожен із вас псалом має, має науку, має мову, об'явлення має, має вияснення, нехай буде все це на збудування!
1COR|14|27|Як говорить хто чужою мовою, говоріть по двох, чи найбільше по трьох, і то за чергою, а один нехай перекладає!
1COR|14|28|А коли б не було перекладача, то нехай він у Церкві мовчить, а говорить нехай собі й Богові!
1COR|14|29|А пророки нехай промовляють по двох чи по трьох, а інші нехай розпізнають.
1COR|14|30|Коли ж відкриття буде іншому з тих, хто сидить, нехай перший замовкне!
1COR|14|31|Бо можете пророкувати ви всі по одному, щоб училися всі й усі тішилися!
1COR|14|32|І коряться духи пророчі пророкам,
1COR|14|33|бо Бог не є Богом безладу, але миру. Як по всіх Церквах у святих,
1COR|14|34|нехай у Церкві мовчать жінки ваші! Бо їм говорити не позволено, тільки коритись, як каже й Закон.
1COR|14|35|Коли ж вони хочуть навчитись чогось, нехай вдома питають своїх чоловіків, непристойно бо жінці говорити в Церкві!
1COR|14|36|Хіба вийшло від вас Слово Боже? Чи прийшло воно тільки до вас?
1COR|14|37|Коли хто вважає себе за пророка або за духовного, нехай розуміє, що я пишу вам, бо Господня це заповідь!
1COR|14|38|Коли б же хто не розумів, нехай не розуміє!
1COR|14|39|Отож, браття мої, майте ревність пророкувати, та не бороніть говорити й мовами!
1COR|14|40|Але все нехай буде добропристойно і статечно!
1COR|15|1|Звіщаю ж вам, браття, Євангелію, яку я вам благовістив, і яку прийняли ви, в якій і стоїте,
1COR|15|2|Якою й спасаєтесь, коли пам'ятаєте, яким словом я благовістив вам, якщо тільки ви ввірували не наосліп.
1COR|15|3|Бо я передав вам найперш, що й прийняв, що Христос був умер ради наших гріхів за Писанням,
1COR|15|4|і що Він був похований, і що третього дня Він воскрес за Писанням,
1COR|15|5|і що з'явився Він Кифі, потім Дванадцятьом.
1COR|15|6|А потім з'явився нараз більше як п'ятистам браттям, що більшість із них живе й досі, а дехто й спочили.
1COR|15|7|Потому з'явився Він Якову, опісля усім апостолам.
1COR|15|8|А по всіх Він з'явився й мені, мов якому недородкові.
1COR|15|9|Я бо найменший з апостолів, що негідний зватись апостолом, бо я переслідував був Божу Церкву.
1COR|15|10|Та благодаттю Божою я те, що є, і благодать Його, що в мені, не даремна була, але я працював більше всіх їх, правда не я, але Божа благодать, що зо мною вона.
1COR|15|11|Тож чи я, чи вони, ми так проповідуємо, і так ви ввірували.
1COR|15|12|Коли ж про Христа проповідується, що воскрес Він із мертвих, як же дехто між вами говорять, що немає воскресення мертвих?
1COR|15|13|Як немає ж воскресення мертвих, то й Христос не воскрес!
1COR|15|14|оли ж бо Христос не воскрес, то проповідь наша даремна, даремна також віра ваша!
1COR|15|15|Ми знайшлися б тоді неправдивими свідками Божими, бо про Бога ми свідчили, що воскресив Він Христа, Якого Він не воскресив, якщо не воскресають померлі.
1COR|15|16|Бо як мертві не воскресають, то й Христос не воскрес!
1COR|15|17|Коли ж бо Христос не воскрес, тоді віра ваша даремна, ви в своїх ще гріхах,
1COR|15|18|тоді то загинули й ті, що в Христі упокоїлись!
1COR|15|19|Коли ми надіємося на Христа тільки в цьому житті, то ми найнещасніші від усіх людей!
1COR|15|20|Та нині Христос воскрес із мертвих, первісток серед покійних.
1COR|15|21|Смерть бо через людину, і через Людину воскресення мертвих.
1COR|15|22|Бо так, як в Адамі вмирають усі, так само в Христі всі оживуть,
1COR|15|23|кожен у своєму порядку: первісток Христос, потім ті, що Христові, під час Його приходу.
1COR|15|24|А потому кінець, коли Він передасть царство Богові й Отцеві, коли Він зруйнує всякий уряд, і владу всяку та силу.
1COR|15|25|Бо належить Йому царювати, аж доки Він не покладе всіх Своїх ворогів під ногами Своїми!
1COR|15|26|Як ворог останній смерть знищиться,
1COR|15|27|бо під ноги Його Він усе впокорив. Коли ж каже, що впокорено все, то ясно, що все, окрім Того, Хто впокорив Йому все.
1COR|15|28|А коли Йому все Він упокорить, тоді й Сам Син упокориться Тому, Хто все впокорив Йому, щоб Бог був у всьому все.
1COR|15|29|Бо що зроблять ті, хто христяться ради мертвих? Коли мертві не воскресають зовсім, то нащо вони ради мертвих і христяться?
1COR|15|30|Для чого й ми повсякчас наражаємось на небезпеки?
1COR|15|31|Я щодень умираю. Так свідчу, браття, вашою хвалою, що маю її в Христі Ісусі, Господі нашім.
1COR|15|32|Коли я зо звірами боровся в Ефесі, яка мені по-людському користь, коли мертві не воскресають? Будем їсти та пити, бо ми взавтра вмрем!...
1COR|15|33|Не дайте себе звести, товариство лихе псує добрі звичаї!
1COR|15|34|Протверезіться правдиво, та й не грішіть, бо деякі Бога не знають, говорю вам на сором!
1COR|15|35|Але дехто скаже: Як мертві воскреснуть? І в якім тілі прийдуть?
1COR|15|36|Нерозумний, що ти сієш, те не оживе, як не вмре.
1COR|15|37|І коли сієш, то сієш не тіло майбутнє, але голе зерно, яке трапиться, пшениці або чого іншого,
1COR|15|38|і Бог йому тіло дає, як захоче, і кожному зерняті тіло його.
1COR|15|39|Не кожне тіло однакове тіло, але ж інше в людей, та інше тіло в скотини, та інше тіло в пташок, та інше у риб.
1COR|15|40|Є небесні тіла й тіла земні, але ж інша слава небесним, а інша земним.
1COR|15|41|Інша слава для сонця, та інша слава для місяця, та інша слава для зір, бо зоря від зорі відрізняється славою!
1COR|15|42|Так само й воскресення мертвих: сіється в тління, в нетління встає,
1COR|15|43|сіється в неславу, у славі встає, сіється в немочі, у силі встає,
1COR|15|44|сіється тіло звичайне, встає тіло духовне. Є тіло звичайне, є й тіло духовне.
1COR|15|45|Так і написано: Перша людина Адам став душею живою, а останній Адам то дух оживляючий.
1COR|15|46|Та не перше духовне, але звичайне, а потім духовне.
1COR|15|47|Перша людина з землі, земна, друга Людина із неба Господь.
1COR|15|48|Який земний, такі й земні, і Який небесний, такі й небесні.
1COR|15|49|І, як носили ми образ земного, так і образ небесного будемо носити.
1COR|15|50|І це скажу, браття, що тіло й кров посісти Божого Царства не можуть, ані тління нетління не посяде.
1COR|15|51|Ось кажу я вам таємницю: не всі ми заснемо, та всі перемінимось,
1COR|15|52|раптом, як оком змигнути, при останній сурмі: бо засурмить вона і мертві воскреснуть, а ми перемінимось!...
1COR|15|53|Мусить бо тлінне оце зодягнутись в нетління, а смертне оце зодягтися в безсмертя.
1COR|15|54|А коли оце тлінне в нетління зодягнеться, і оце смертне в безсмертя зодягнеться, тоді збудеться слово написане: Поглинута смерть перемогою!
1COR|15|55|Де, смерте, твоя перемога? Де твоє, смерте, жало?
1COR|15|56|Жало ж смерти то гріх, а сила гріха то Закон.
1COR|15|57|А Богові дяка, що Він Господом нашим Ісусом Христом перемогу нам дав.
1COR|15|58|Отож, брати любі мої, будьте міцні, непохитні, збагачуйтесь завжди в Господньому ділі, знаючи, що ваша праця не марнотна у Господі!
1COR|16|1|А щодо складок на святих, то й ви робіть так, як я постановив для Церков галатійських.
1COR|16|2|А першого дня в тижні нехай кожен із вас відкладає собі та збирає, згідно з тим, як ведеться йому, щоб складок не робити тоді, аж коли я прийду.
1COR|16|3|А коли я прийду, тоді тих, кого виберете, тих пошлю я з листами, щоб вони ваш дар любови віднесли до Єрусалиму.
1COR|16|4|А коли ж і мені випадатиме йти, то зо мною підуть.
1COR|16|5|Я прибуду до вас, коли перейду Македонію, бо проходжу через Македонію.
1COR|16|6|А в вас, коли трапиться, я поживу або й перезимую, щоб мене провели ви, куди я піду.
1COR|16|7|Не хочу я бачитись з вами тепер мимохідь, але сподіваюся деякий час перебути у вас, як дозволить Господь.
1COR|16|8|А в Ефесі пробуду я до П'ятдесятниці,
1COR|16|9|бо двері великі й широкі мені відчинилися, та багато противників...
1COR|16|10|Коли ж прийде до вас Тимофій, то пильнуйте, щоб він був безпечний у вас, бо діло Господнє він робить, як і я.
1COR|16|11|Тому то нехай ним ніхто не погорджує, але відпровадьте його з миром, щоб прийшов він до мене, бо чекаю його з братами.
1COR|16|12|А щодо брата Аполлоса, то я дуже благав був його, щоб прийшов до вас з братами, та охоти не мав він прибути тепер, але прийде, як матиме час відповідний.
1COR|16|13|Пильнуйте, стійте у вірі, будьте мужні, будьте міцні,
1COR|16|14|хай з любов'ю все робиться в вас!
1COR|16|15|Благаю ж вас, браття, знаєте ви дім Степанів, що в Ахаї він первісток, і що службі святим присвятились вони,
1COR|16|16|і ви підкоряйтесь таким, також кожному, хто помагає та працює.
1COR|16|17|Я тішусь з приходу Степана, і Фортуната, і Ахаїка, бо вашу відсутність вони заступили,
1COR|16|18|бо вони заспокоїли духа мого й вашого. Тож шануйте таких!
1COR|16|19|Вітають вас азійські Церкви; Акила й Прискилла з домашньою Церквою їхньою гаряче вітають у Господі вас.
1COR|16|20|Вітають вас усі брати. Вітайте один одного святим поцілунком.
1COR|16|21|Привітання моєю рукою Павловою.
1COR|16|22|Коли хто не любить Господа, нехай буде проклятий! Марана та!
1COR|16|23|Благодать Господа нашого Ісуса нехай буде з вами!
1COR|16|24|Любов моя з вами всіма у Христі Ісусі, амінь!
