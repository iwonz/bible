EPH|1|1|奉上帝旨意作基督耶稣使徒的 保罗 ，写信给在 以弗所 的 众圣徒，就是在基督耶稣里忠心的人。
EPH|1|2|愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
EPH|1|3|愿颂赞归给我们主耶稣基督的父上帝。他在基督里曾把天上各样属灵的福气赐给我们。
EPH|1|4|因为他从创世以前，在基督里拣选了我们，使我们在他面前成为圣洁，没有瑕疵，满有爱心。
EPH|1|5|他按着自己旨意所喜悦的 ，预定我们藉着耶稣基督得儿子的名分，
EPH|1|6|使他荣耀的恩典得到称赞；这恩典是他在爱子里白白赐给我们的。
EPH|1|7|我们藉着这爱子的血得蒙救赎，过犯得以赦免，这是照他丰富的恩典，
EPH|1|8|充充足足地赏给我们的。他以诸般的智慧聪明，
EPH|1|9|照自己在基督里所立定的美意，使我们知道他旨意的奥秘，
EPH|1|10|要照着所安排的，在时机成熟的时候，使天上、地上、一切所有的，都在基督里面同归于一。
EPH|1|11|我们也在他里面得了基业；这原是那位随己意行万事的上帝照着自己的旨意所预定的，
EPH|1|12|为要使我们，这些首先把希望寄托在基督里的人，颂赞他的荣耀。
EPH|1|13|在基督里你们听见真理的道，就是那使你们得救的福音，你们也信了他，就受了所应许的圣灵为印记。
EPH|1|14|这圣灵是我们得基业的凭据，直等到上帝的子民得救赎，使他的荣耀得到称赞。
EPH|1|15|因此，我既然听见你们对主耶稣有信心，对众圣徒有爱心，
EPH|1|16|就不住地为你们感谢上帝，祷告的时候常常提到你们，
EPH|1|17|求我们主耶稣基督的上帝，荣耀的父，把那赐人智慧和启示的灵赐给你们，使你们真正认识他，
EPH|1|18|照亮你们心中的眼睛，使你们知道他呼召你们来得的指望是什么，他在圣徒中所得荣耀的基业是何等丰盛，
EPH|1|19|并知道他向我们这些信的人所显的能力是何等浩大，这是照他的大能大力运行的。
EPH|1|20|这大能曾运行在基督身上，使他从死人中复活，又使他在天上坐在自己的右边，
EPH|1|21|远超越一切执政的、掌权的、有权能的、统治的和一切有名号的；不但是今世的，连来世的也都超越了。
EPH|1|22|上帝使万有服在他的脚下，又使他为了教会作万有之首；
EPH|1|23|教会是他的身体，是那充满万有者所充满的。
EPH|2|1|从前，你们因着自己的过犯罪恶而死了。
EPH|2|2|那时，你们在过犯罪恶中生活，随从今世的风俗，顺服空中掌权者的领袖，就是现今在悖逆的人心中运行的邪灵。
EPH|2|3|我们从前也都生活在他们当中，放纵肉体的私欲，随着肉体和心中的意念去做，和别人一样，生来就是该受惩罚的人。
EPH|2|4|然而，上帝有丰富的怜悯，因着他爱我们的大爱，
EPH|2|5|竟在我们因过犯而死了的时候，使我们与基督一同活过来—可见你们得救是本乎恩—
EPH|2|6|他又使我们在基督耶稣里与他一同复活，一同坐在天上，
EPH|2|7|为要把他极丰富的恩典，就是他在基督耶稣里向我们所施的恩慈，显明给后来的世代。
EPH|2|8|你们得救是本乎恩，也因着信；这并不是出于自己，而是上帝所赐的；
EPH|2|9|也不是出于行为，免得有人自夸。
EPH|2|10|我们是他所造之物，在基督耶稣里创造的，为要使我们行善，就是上帝早已预备好要我们做的。
EPH|2|11|所以，你们要记得：从前你们按肉体是外邦人，是“没受割礼的”；这名字是那些凭人手在肉身上“受割礼的人”所取的。
EPH|2|12|要记得那时候，你们与基督无关，与 以色列 选民团体隔绝，在所应许的约上是局外人，而且在世上没有指望，没有上帝。
EPH|2|13|从前你们是远离上帝的人，如今却在基督耶稣里，靠着他的血，已经得以亲近了。
EPH|2|14|因为他自己是我们的和平 ，使双方合而为一，拆毁了中间隔绝的墙，而且以自己的身体终止了冤仇，
EPH|2|15|废掉那记在律法上的规条，为要使两方藉着自己造成一个新人，促成了和平；
EPH|2|16|既在十字架上消灭了冤仇，就藉这十字架使双方归为一体，与上帝和好，
EPH|2|17|并且来传和平的福音给你们远处的人，也传和平给那些近处的人，
EPH|2|18|因为我们双方藉着他，在同一位圣灵里得以进到父面前。
EPH|2|19|这样，你们不再是外人或客旅，是与圣徒同国，是上帝家里的人了，
EPH|2|20|被建造在使徒和先知的根基上，而基督耶稣自己为房角石，
EPH|2|21|靠着他整座房子连接得紧凑，渐渐成为在主里的圣殿。
EPH|2|22|你们也靠他同被建造，成为上帝藉着圣灵居住的所在。
EPH|3|1|因此，我— 保罗 为你们外邦人作了基督耶稣 囚徒的，替你们祈祷 。
EPH|3|2|想你们必曾听见上帝赐恩给我，把关切你们的职分托付我，
EPH|3|3|用启示让我知道福音的奥秘，正如我以前略略写过的。
EPH|3|4|你们读了，就会知道我深深了解基督的奥秘；
EPH|3|5|这奥秘在以前的世代没有让人知道，像如今藉着圣灵向他的圣使徒和先知启示一样，
EPH|3|6|就是外邦人在基督耶稣里，藉着福音，得以同为后嗣，同为一体，同为蒙应许的人。
EPH|3|7|我作了这福音的仆役，是照着上帝的恩赐，是照他运行的大能赐给我的。
EPH|3|8|虽然我比众圣徒中最小的还小，他还赐我这恩典，让我把基督那测不透的丰富传给外邦人，
EPH|3|9|又使众人都明白 什么是历代以来隐藏在创造万物之上帝里的奥秘，
EPH|3|10|为要在现今藉着教会使天上执政的、掌权的知道上帝百般的智慧。
EPH|3|11|这是照着上帝在我们主基督耶稣里所完成的永恒的计划。
EPH|3|12|我们因信耶稣 ，就在他里面放胆无惧，满有自信地进到上帝面前。
EPH|3|13|所以我求你们，不要因我为你们所受的患难丧胆；这原是你们的光荣。
EPH|3|14|因此，我在父面前屈膝—
EPH|3|15|天上地上的各家都是从他得名的－
EPH|3|16|为要他按着他丰盛的荣耀，藉着他的灵，使你们内心的力量刚强起来；
EPH|3|17|又要他使基督因着你们的信住在你们心里，使你们既在爱中生根立基，
EPH|3|18|能够和众圣徒一同明白基督的爱是何等的长、阔、高、深，并知道这爱是超过人的知识所能测度的，为要使你们充满上帝一切的丰盛。
EPH|3|19|
EPH|3|20|上帝能照着运行在我们心里的大能充充足足地成就一切，超过我们所求所想的。
EPH|3|21|愿他在教会中，并在基督耶稣里，得着荣耀，直到世世代代，永永远远。阿们！
EPH|4|1|我为主作囚徒的劝你们，既然蒙召，行事为人就要与你们所蒙的呼召相称。
EPH|4|2|凡事要谦虚、温柔、忍耐，用爱心互相宽容，
EPH|4|3|以和平彼此联系，竭力保持圣灵所赐的合一。
EPH|4|4|身体只有一个，圣灵只有一位，正如你们蒙召，是为同有一个指望而蒙召，
EPH|4|5|一主，一信，一洗，
EPH|4|6|一上帝－就是万人之父，超越万有之上，贯通万有，在万有之中。
EPH|4|7|我们每个人蒙恩都是照基督所量给每个人的恩赐。
EPH|4|8|所以有话说： “他升上高天的时候，掳掠了俘虏， 将各样的恩赐赏给人。”
EPH|4|9|既说“他升上”，岂不是指他曾降到地底下吗？
EPH|4|10|那降下的，就是高升远超越诸天之上的，为要充满万有。
EPH|4|11|他所赐的有使徒，有先知，有传福音的，有牧者和教师，
EPH|4|12|为要装备圣徒，做事奉的工作，建立基督的身体，
EPH|4|13|直等到我们众人在信仰上同归于一，认识上帝的儿子，得以长大成人，达到基督完全长成的身量。
EPH|4|14|这样，我们不再作小孩子，中了人的诡计和欺骗的法术，被一切邪说之风摇动，飘来飘去。
EPH|4|15|我们反而要用爱心说诚实话，各方面向着基督长进，连于元首基督，
EPH|4|16|靠着他全身都连接得紧凑，百节各按各职，照着各体的功用彼此相助，使身体渐渐增长，在爱中建立自己。
EPH|4|17|所以我这样说，且在主里郑重地说，你们行事为人，不要再像外邦人存虚妄的心而活。
EPH|4|18|他们心地昏昧，因自己无知，心里刚硬而与上帝所赐的生命隔绝了。
EPH|4|19|既然他们已经麻木，就放纵情欲，贪婪地行种种污秽的事。
EPH|4|20|但你们从基督学的不是这样。
EPH|4|21|如果你们听过他的道，领了他的教，因为真理就在耶稣里，
EPH|4|22|你们要脱去从前的行为，脱去旧我；这旧我是因私欲的迷惑而渐渐败坏的。
EPH|4|23|你们要把自己的心志更新，
EPH|4|24|并且穿上新我；这新我是照着上帝的形像造的，有从真理来的公义和圣洁。
EPH|4|25|所以，你们要弃绝谎言，每个人要与邻舍说诚实话，因为我们是互为肢体。
EPH|4|26|即使生气也不要犯罪；不可含怒到日落，
EPH|4|27|不可给魔鬼留地步。
EPH|4|28|偷窃的，不要再偷；总要勤劳，亲手 做正当的事，这样才可以把自己有的，分给有缺乏的人。
EPH|4|29|一句坏话也不可出口，只要随着需要说造就人的好话，让听见的人得益处。
EPH|4|30|不要使上帝的圣灵担忧，你们原是受了他的印记，等候得救赎的日子来到。
EPH|4|31|一切苦毒、愤怒、恼恨、嚷闹、毁谤，和一切的恶毒都要从你们中间除掉。
EPH|4|32|要仁慈相待，存怜悯的心，彼此饶恕，正如上帝在基督里饶恕了你们一样。
EPH|5|1|所以，作为蒙慈爱的儿女，你们该效法上帝。
EPH|5|2|要凭爱心行事，正如基督爱我们，为我们舍了自己，当作馨香的供物和祭物献给上帝。
EPH|5|3|至于淫乱和一切污秽，或是贪婪，在你们中间连提都不可，这才合乎圣徒的体统。
EPH|5|4|淫词、妄语和粗俗的俏皮话都不合宜；总要说感谢的话。
EPH|5|5|要确实知道，无论是淫乱的，是污秽的，是贪心的（贪心的就是拜偶像的），在基督和上帝的国里都得不到基业。
EPH|5|6|不要被人虚浮的话欺骗了，因这些事，上帝的愤怒必临到那些悖逆的人。
EPH|5|7|所以，不要与他们同伙。
EPH|5|8|从前你们是暗昧的，但如今在主里面是光明的，行事为人要像光明的子女—
EPH|5|9|光明所结的果子就是一切的良善、公义、诚实。
EPH|5|10|总要察验什么是主所喜悦的事。
EPH|5|11|那暗昧无益的事，不可参与，倒要把这种事揭发出来。
EPH|5|12|因为，他们暗中所做的，就是连提起来都是可耻的。
EPH|5|13|凡被光所照明的都显露出来，
EPH|5|14|因为使一切显露出来的就是光。所以有话说： “你这睡着的人醒过来吧！ 要从死人中复活， 基督要光照你了。”
EPH|5|15|你们要谨慎行事，不要像无知的人，要像智慧的人。
EPH|5|16|要把握时机 ，因为现今的世代邪恶。
EPH|5|17|不要作糊涂人，要明白主的旨意如何。
EPH|5|18|不要醉酒，酒能使人放荡；要被圣灵充满。
EPH|5|19|要用诗篇、赞美诗、灵歌彼此对说，口唱心和地赞美主。
EPH|5|20|凡事要奉我们主耶稣基督的名常常感谢父上帝。
EPH|5|21|要存敬畏基督的心彼此顺服。
EPH|5|22|作妻子的，你们要顺服自己的丈夫，如同顺服主。
EPH|5|23|因为丈夫是妻子的头，如同基督是教会的头；他又是这身体的救主。
EPH|5|24|教会怎样顺服基督，妻子也要怎样凡事顺服丈夫。
EPH|5|25|作丈夫的，你们要爱自己的妻子，正如基督爱教会，为教会舍己，
EPH|5|26|以水藉着道把教会洗净，使她成为圣洁，
EPH|5|27|好献给自己，作荣耀的教会，毫无玷污、皱纹等类的缺陷，而是圣洁没有瑕疵的。
EPH|5|28|丈夫也应当照样爱妻子，如同爱自己的身体；爱妻子就是爱自己了。
EPH|5|29|从来没有人恨恶自己的身体，总是保养爱惜，正像基督待教会一样，
EPH|5|30|因我们是他身体的肢体。
EPH|5|31|“为这个缘故，人要离开父母，与妻子结合，二人成为一体。”
EPH|5|32|这是极大的奥秘，而我是指基督和教会说的。
EPH|5|33|然而，你们每个人都要爱妻子，如同爱自己一样；妻子也要敬重她的丈夫。
EPH|6|1|作儿女的，你们要在主里 听从父母，这是理所当然的。
EPH|6|2|当孝敬父母，使你得福，在世长寿。这是第一条带应许的诫命。
EPH|6|3|
EPH|6|4|作父亲的，你们不要激怒儿女，但要照着主的教导和劝戒养育他们。
EPH|6|5|作仆人的，你们要惧怕战兢，用诚实的心听从你们肉身的主人，好像听从基督一般；
EPH|6|6|不要只在人的眼前这样做，像仅是讨人的喜欢，而是作基督的仆人，从心里遵行上帝的旨意，
EPH|6|7|甘心服侍，好像服侍主，不像服侍人，
EPH|6|8|因为知道每个人所做的善事，不论是为奴的或是自主的，都必按所做的从主得到赏赐。
EPH|6|9|作主人的，你们待仆人也是一样，不要威吓他们，因为知道他们和你们在天上同有一位主，他并不偏待人。
EPH|6|10|最后，你们要靠着主，依赖他的大能大力作刚强的人。
EPH|6|11|要穿戴上帝所赐的全副军装，好抵挡魔鬼的诡计。
EPH|6|12|因为我们的争战并不是对抗有血有肉的人，而是对抗那些执政的、掌权的、管辖这幽暗世界的，以及天空灵界的恶魔。
EPH|6|13|所以，要拿起上帝所赐的全副军装，好在邪恶的日子能抵挡仇敌，并且完成了一切后还能站立得住。
EPH|6|14|所以，要站稳了，用真理当作带子束腰，用公义当作护心镜遮胸，
EPH|6|15|又用和平的福音当作预备走路的鞋穿在脚上。
EPH|6|16|此外，要拿信德当作盾牌，用来扑灭那恶者一切烧着的箭。
EPH|6|17|要戴上救恩的头盔，拿着圣灵的宝剑—就是上帝的道。
EPH|6|18|要靠着圣灵，随时多方祷告祈求，并要为此警醒不倦，为众圣徒祈求。
EPH|6|19|也要为我祈求，让我有口才，能放胆开口讲明福音的奥秘，
EPH|6|20|我为这福音的奥秘作了带铁链的使者，让我能照着当尽的本分放胆宣讲。
EPH|6|21|今有亲爱、忠心服事主的弟兄 推基古 ，为了你们也明白我的事情和我的景况，他会让你们知道一切的事。
EPH|6|22|我特意打发他到你们那里去，好让你们知道我们的情况，又让他安慰你们的心。
EPH|6|23|愿平安 、慈爱、信心从父上帝和主耶稣基督归给弟兄们。
EPH|6|24|愿所有恒心爱我们主耶稣基督的人都蒙恩惠。
