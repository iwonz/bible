MARK|1|1|Початок Євангелії Ісуса Христа, Сина Божого.
MARK|1|2|Як у пророка Ісаї написано: Ось перед обличчя Твоє посилаю Свого посланця, який перед Тобою дорогу Твою приготує.
MARK|1|3|Голос того, хто кличе: У пустині готуйте дорогу для Господа, рівняйте стежки Йому!
MARK|1|4|виступив був так Іван, що в пустині христив та проповідував хрищення на покаяння для прощення гріхів.
MARK|1|5|І до нього приходила вся країна Юдейська та всі єрусалимляни, і в річці Йордані від нього христились вони, і визнавали гріхи свої.
MARK|1|6|А Іван зодягався в одежу з верблюжого волосу, і мав пояс ремінний на стегнах своїх, а їв сарану та мед польовий.
MARK|1|7|І він проповідував, кажучи: Услід за мною йде он Потужніший від мене, що Йому я негідний, нагнувшись, розв'язати ремінця від узуття Його.
MARK|1|8|Я христив вас водою, а Той вас христитиме Духом Святим.
MARK|1|9|І сталося тими днями, прийшов Ісус з Назарету Галілейського, і від Івана христився в Йордані.
MARK|1|10|І зараз, коли Він виходив із води, то побачив Іван небо розкрите, і Духа, як голуба, що сходив на Нього.
MARK|1|11|І голос із неба почувся: Ти Син Мій Улюблений, що Я вподобав Його!
MARK|1|12|І зараз повів Його Дух у пустиню.
MARK|1|13|І Він був сорок днів у пустині, випробовуваний від сатани, і перебував зо звіриною. І служили Йому Анголи.
MARK|1|14|А коли Іван виданий був, то прийшов Ісус до Галілеї, і проповідував Божу Євангелію,
MARK|1|15|і говорив: Збулися часи, і Боже Царство наблизилось. Покайтеся, і віруйте в Євангелію!
MARK|1|16|А коли Він проходив біля Галілейського моря, то побачив Симона та Андрія, брата Симонового, що невода в море закидали, бо рибалки були.
MARK|1|17|І сказав їм Ісус: Ідіть услід за Мною, і зроблю, що станете ви ловцями людей.
MARK|1|18|І зараз вони свого невода кинули, та й пішли вслід за Ним.
MARK|1|19|А коли недалеко прийшов, то побачив Він Якова Зеведеєвого та брата його Івана, що й вони в човні невода лагодили.
MARK|1|20|І зараз покликав Він їх. І вони залишили батька свого Зеведея в човні з робітниками, і пішли вслід за Ним.
MARK|1|21|І приходять вони в Капернаум. І негайно в суботу ввійшов Він у синагогу, і навчати зачав.
MARK|1|22|І дивувались науці Його, бо навчав Він їх, як можновладний, а не як ті книжники.
MARK|1|23|І зараз у їхній синагозі знайшовся один чоловік, що мав духа нечистого, і він закричав,
MARK|1|24|і сказав: Що Тобі до нас, Ісусе Назарянине? Ти прийшов погубити нас. Я знаю Тебе, хто Ти, Божий Святий.
MARK|1|25|Ісус же йому заказав: Замовчи, і вийди з нього!
MARK|1|26|І затряс дух нечистий того, і, скрикнувши голосом гучним, вийшов із нього.
MARK|1|27|І жахнулися всі, аж питали вони один одного, кажучи: Що це таке? Нова наука із потугою! Навіть духам нечистим наказує Він, і вони Його слухають.
MARK|1|28|І чутка про Нього пішла хвилі тієї по всій Галілейській країні.
MARK|1|29|І вийшли вони із синагоги небавом, і прийшли з Яковом та Іваном до дому Симонового й Андрієвого.
MARK|1|30|А теща Симонова лежала в гарячці; і зараз сказали про неї Йому.
MARK|1|31|І Він підійшов і підвів її, узявши за руку, і гарячка покинула ту, і вона зачала прислуговувати їм.
MARK|1|32|А як вечір настав, коли сонце зайшло, то стали приносити до Нього недужих усіх та біснуватих.
MARK|1|33|І все місто зібралося перед дверима.
MARK|1|34|І Він уздоровив багатьох, на різні хвороби недужих, і багатьох демонів повиганяв. А демонам не дозволяв Він казати, що знають Його.
MARK|1|35|А над ранком, як дуже ще темно було, уставши, Він вийшов і пішов у місце самітне, і там молився.
MARK|1|36|А Симон та ті, що були з ним, поспішили за Ним.
MARK|1|37|І, знайшовши Його, вони кажуть Йому: Усі шукають Тебе.
MARK|1|38|А Він промовляє до них: Ходім в інше місце, до сіл та околишніх міст, щоб і там проповідувати, бо на те Я прийшов.
MARK|1|39|І пішов, і проповідував в їхніх синагогах по всій Галілеї. І демонів Він виганяв.
MARK|1|40|І приходить до Нього прокажений, благає Його, і на коліна впадає та й каже Йому: Коли хочеш, Ти можеш очистити мене!
MARK|1|41|І змилосердився Він, простяг руку Свою, і доторкнувся до нього, та й каже йому: Хочу, будь чистий!
MARK|1|42|І проказа зійшла з нього хвилі тієї, і чистим він став.
MARK|1|43|А Він, погрозивши йому, зараз вислав його,
MARK|1|44|і йому наказав: Гляди, не оповідай нічого нікому. Але йди, покажися священикові, і принеси за своє очищення, що Мойсей заповів, їм на свідоцтво.
MARK|1|45|А він, вийшовши, став багато оповідати й говорити про подію, так що Він не міг явно ввійти вже до міста, але перебував віддалік по самітних місцях. І сходилися звідусюди до Нього.
MARK|2|1|Коли ж Він по кількох днях прийшов знов до Капернауму, то чутка пішла, що Він удома.
MARK|2|2|І зібралось багато, аж вони не вміщалися навіть при дверях. А Він їм виголошував слово.
MARK|2|3|І прийшли ось до Нього, несучи розслабленого, якого несли четверо.
MARK|2|4|А що через народ до Нього наблизитися не могли, то стелю розкрили, де Він був, і пробравши, звісили ложе, що на ньому лежав розслаблений.
MARK|2|5|А Ісус, віру їхню побачивши, каже розслабленому: Відпускаються, сину, гріхи тобі!
MARK|2|6|Там же сиділи дехто з книжників, і в серцях своїх думали:
MARK|2|7|Чого Він говорить отак? Зневажає Він Бога... Хто може прощати гріхи, окрім Бога Самого?
MARK|2|8|І зараз Ісус відчув Духом Своїм, що вони так міркують собі, і сказав їм: Що таке ви в серцях своїх думаєте?
MARK|2|9|Що легше: сказати розслабленому: Гріхи відпускаються тобі, чи сказати: Уставай, візьми ложе своє та й ходи?
MARK|2|10|Але щоб ви знали, що Син Людський має владу прощати гріхи на землі, каже розслабленому:
MARK|2|11|Тобі Я наказую: Уставай, візьми ложе своє, та й іди у свій дім!
MARK|2|12|І той устав, і негайно взяв ложе, і вийшов перед усіма, так що всі дивувались і славили Бога, й казали: Ніколи такого не бачили ми!
MARK|2|13|І вийшов над море Він знов. А ввесь натовп до Нього приходив, і Він їх навчав.
MARK|2|14|А коли Він проходив, то побачив Левія Алфієвого, що сидів на митниці, і каже йому: Іди за Мною! Той устав, і пішов услід за Ним.
MARK|2|15|Коли ж Він сидів при столі в його домі, то багато митників і грішників сиділи з Ісусом та з учнями Його; бо було їх багато, і вони ходили за Ним.
MARK|2|16|Як побачили ж книжники та фарисеї, що Він їсть із грішниками та з митниками, то сказали до учнів Його: Чому то Він їсть із митниками та з грішниками?
MARK|2|17|А Ісус, як почув, промовляє до них: Лікаря не потребують здорові, а слабі. Я не прийшов кликати праведних, але грішників на покаяння.
MARK|2|18|А учні Іванові та фарисейські постили. І приходять вони, та й говорять до Нього: Чому учні Іванові та фарисейські постять, а учні Твої не постять?
MARK|2|19|Ісус же промовив до них: Хіба постити можуть гості весільні, поки з ними ще є молодий? Доки мають вони молодого з собою, то постити не можуть.
MARK|2|20|Але прийдуть ті дні, коли заберуть молодого від них, то й постити будуть вони за тих днів.
MARK|2|21|І не пришиває ніхто до старої одежі латки з сукна сирового, а як ні, то край латки нової одірветься там від старого, і дірка стане ще гірша.
MARK|2|22|І ніхто не вливає вина молодого в старі бурдюки, а то попрориває вино бурдюки, і вино й бурдюки пропадуть, а вливають вино молоде до нових бурдюків.
MARK|2|23|І сталось, як Він переходив ланами в суботу, Його учні дорогою йшли, та й стали колосся зривати.
MARK|2|24|Фарисеї ж казали Йому: Подивись, чому роблять у суботу вони, чого не годиться?
MARK|2|25|А Він їм відказав: Чи ж ви не читали ніколи, що зробив був Давид, як потребу він мав та сам зголоднів був і ті, що були з ним?
MARK|2|26|Як він увійшов був до Божого дому за первосвященика Авіятара, і спожив хліби показні, яких їсти не можна було, тільки священикам, і дав він і тим, хто був із ним?
MARK|2|27|І сказав Він до них: Субота постала для чоловіка, а не чоловік для суботи,
MARK|2|28|а тому то Син Людський Господь і суботі.
MARK|3|1|І Він знову до синагоги ввійшов. І був там один чоловік, який мав суху руку.
MARK|3|2|І, щоб обвинуватити Його, наглядали за Ним, чи Він у суботу того не вздоровить.
MARK|3|3|І говорить Він до чоловіка з сухою рукою: Стань посередині!
MARK|3|4|А до них промовляє: У суботу годиться робити добре, чи робити лихе, життя зберегти, чи погубити? Вони ж мовчали.
MARK|3|5|І споглянув Він із гнівом на них, засмучений закам'янілістю їхніх сердець, і сказав чоловікові: Простягни свою руку! І той простяг, і рука йому стала здорова!
MARK|3|6|Фарисеї ж негайно пішли та з іродіянами раду зробили на Нього, як Його погубити.
MARK|3|7|А Ісус із Своїми учнями вийшов над море. І натовп великий ішов вслід за Ним із Галілеї й з Юдеї,
MARK|3|8|і з Єрусалиму, і з Ідумеї, і з-за Йордання, і з Тиру й Сидону. Натовп великий, прочувши, як багато чинив Він, зібрався до Нього.
MARK|3|9|І сказав Він до учнів Своїх наготовити човна Йому, через натовп, щоб до Нього не тиснулись.
MARK|3|10|Бо Він багатьох уздоровив, так що хто тільки немочі мав, то тислись до Нього, щоб Його доторкнутись.
MARK|3|11|І духи нечисті, як тільки вбачали Його, то падали ницьма перед Ним, і кричали й казали: Ти Син Божий!
MARK|3|12|А Він їм суворо наказував, щоб вони Його не виявляли.
MARK|3|13|І Він вийшов на гору, і покликав, кого Сам хотів; вони ж приступили до Нього.
MARK|3|14|І визначив Дванадцятьох, щоб із Ним перебували, і щоб послати на проповідь їх,
MARK|3|15|і щоб мали вони владу вздоровляти недуги й вигонити демонів.
MARK|3|16|І визначив Він оцих Дванадцятьох: Симона, і дав йому ймення Петро,
MARK|3|17|і Якова Зеведеєвого, і Івана, брата Якова, і дав їм імена Воанергес, цебто сини громові,
MARK|3|18|і Андрія, і Пилипа, і Варфоломія, і Матвія, і Хому, і Якова Алфієвого, і Тадея, і Симона Кананіта
MARK|3|19|та Юду Іскаріотського, що й видав Його.
MARK|3|20|І приходять до дому вони. І знову зібралось народу, що вони не могли навіть хліба з'їсти.
MARK|3|21|І коли Його ближчі почули, то вийшли, щоб узяти Його, бо говорено, ніби Він несамовитий.
MARK|3|22|А книжники, що поприходили з Єрусалиму, казали: Має Він Вельзевула, і виганяє демонів силою князя демонів.
MARK|3|23|І, закликавши їх, Він у притчах до них промовляв: Як може сатана сатану виганяти?
MARK|3|24|І коли царство поділиться супроти себе, не може встояти те царство.
MARK|3|25|І коли дім поділиться супроти себе, не може встояти той дім.
MARK|3|26|І коли б сатана сам на себе повстав і поділився, то не зможе встояти він, але згине.
MARK|3|27|Ніхто бо не може вдертись у дім дужого, та й пограбувати добро його, якщо перше не зв'яже дужого, і аж тоді пограбує господу його.
MARK|3|28|Поправді кажу вам, що простяться людським синам усі прогріхи та богозневаги, хоч би як вони богозневажали.
MARK|3|29|Але, хто богозневажить Духа Святого, повіки йому не відпуститься, але гріху вічному він підпадає.
MARK|3|30|Бож казали вони: Він духа нечистого має.
MARK|3|31|І поприходили мати Його та брати Його, і, осторонь ставши, послали до Нього і Його викликали.
MARK|3|32|А народ кругом Нього сидів. І сказали Йому: Ото мати Твоя, і брати Твої, і сестри Твої он про Тебе питаються осторонь.
MARK|3|33|А Він їм відповів і сказав: Хто Моя мати й брати?
MARK|3|34|І поглянув на тих, що круг Нього сиділи, і промовив: Ось мати Моя та браття Мої!
MARK|3|35|Бо хто Божу волю чинитиме, той Мені брат, і сестра, і мати.
MARK|4|1|І знову почав Він навчати над морем. І зібралось до Нього багато народу, так що Сам Він до човна на морі ввійшов і сидів, а народ увесь був на землі покрай моря.
MARK|4|2|І багато навчав Він їх притчами, і в науці Своїй їм казав:
MARK|4|3|Слухайте, вийшов сіяч ось, щоб сіяти.
MARK|4|4|І як сіяв, упало зерно одне край дороги, і налетіли пташки, і його повидзьобували.
MARK|4|5|Друге ж упало на ґрунт кам'янистий, де не мало багато землі, і негайно зійшло, бо земля неглибока була;
MARK|4|6|а як сонце зійшло то зів'яло, і, коріння не мавши, усохло.
MARK|4|7|А інше впало між терен, і вигнався терен, і його поглушив, і плоду воно не дало.
MARK|4|8|Інше ж упало на добрую землю, і дало плід, що посходив і ріс; і видало втридцятеро, у шістдесят і в сто раз.
MARK|4|9|І сказав: Хто має вуха, щоб слухати, нехай слухає!
MARK|4|10|І, як остався Він насамоті, Його запитали найближчі з Дванадцятьма про цю притчу.
MARK|4|11|І Він їм відповів: Вам дано пізнати таємниці Божого Царства, а тим, що за вами, усе відбувається в притчах,
MARK|4|12|щоб оком дивились вони і не бачили, вухом слухали і не зрозуміли, щоб коли вони не навернулися, і відпущені будуть гріхи їм!
MARK|4|13|І Він їх запитав: Ви не розумієте притчі цієї? І як вам зрозуміти всі притчі!
MARK|4|14|Сіяч сіє слово.
MARK|4|15|А котрі край дороги, де сіється слово, це ті, що як тільки почують, то зараз приходить до них сатана, і забирає слово, посіяне в них.
MARK|4|16|Так само й посіяні на кам'янистому ґрунті, вони, як почують те слово, то з радістю зараз приймають його,
MARK|4|17|та коріння не мають у собі й непостійні; а згодом, як утиск або переслідування наступає за слово, вони спокушаються зараз.
MARK|4|18|А між терен посіяне, це ті, що слухають слово,
MARK|4|19|але клопоти цьогосвітні й омана багатства та різні бажання ввіходять, та й заглушують слово, і плоду воно не дає.
MARK|4|20|А посіяне в добрую землю це ті, що слухають слово й приймають, і родять утридцятеро, у шістдесят і в сто раз.
MARK|4|21|І сказав Він до них: Чи світильника приносять на те, щоб поставити його під посудину, чи може під ліжко? А не щоб поставити на свічнику?
MARK|4|22|Бо немає нічого захованого, що не виявиться, і немає таємного, що не вийде наяв.
MARK|4|23|Хто має вуха, щоб слухати, нехай слухає!
MARK|4|24|І сказав Він до них: Уважайте, що чуєте: Якою мірою будете міряти, такою відміряють вам, і додадуть вам.
MARK|4|25|Бо хто має, то дасться йому, хто ж не має, забереться від нього й те, що він має.
MARK|4|26|І сказав Він: Так і Боже Царство, як той чоловік, що кидає в землю насіння,
MARK|4|27|і чи спить, чи встає він удень та вночі, а насіння пускає паростки та росте, хоч не знає він, як.
MARK|4|28|Бо родить земля сама з себе: перше вруна, потім колос, а тоді повне збіжжя на колосі.
MARK|4|29|А коли плід доспіє, зараз він посилає серпа, бо настали жнива.
MARK|4|30|І сказав Він: До чого прирівняємо Царство Боже? Або в якій притчі представим його?
MARK|4|31|Воно як те зерно гірчичне, яке, коли сіється в землю, найдрібніше за всі земні насіння.
MARK|4|32|Як посіяне ж буде, виростає, і стає над усі зілля більше, і віття пускає велике таке, що кублитись може в тіні його птаство небесне.
MARK|4|33|І такими притчами багатьома Він їм слово звіщав, поскільки вони могли слухати.
MARK|4|34|І без притчі нічого Він їм не казав, а учням Своїм самотою вияснював усе.
MARK|4|35|І сказав Він до них того дня, коли вечір настав: Переплиньмо на той бік.
MARK|4|36|І, лишивши народ, узяли із собою Його, як у човні Він був; і інші човни були з Ним.
MARK|4|37|І знялася ось буря велика, а хвилі вливалися в човен, аж човен водою вже був переповнився!
MARK|4|38|А Він спав на кормі на подушці... І вони розбудили Його та й сказали Йому: Учителю, чи Тобі байдуже, що ми гинемо?...
MARK|4|39|Тоді Він устав, і вітрові заборонив, і до моря сказав: Мовчи, перестань! І стих вітер, і тиша велика настала...
MARK|4|40|І сказав Він до них: Чого ви такі полохливі? Чому віри не маєте?
MARK|4|41|А вони налякалися страхом великим, і говорили один до одного: Хто ж це такий, що вітер і море слухняні Йому?
MARK|5|1|І на другий бік моря вони прибули, до землі Гадаринської.
MARK|5|2|І як вийшов Він із човна, то зараз Його перестрів чоловік із могильних печер, що мав духа нечистого.
MARK|5|3|Він мешкання мав у гробах, і ніхто й ланцюгами зв'язати не міг його,
MARK|5|4|бо часто кайданами та ланцюгами в'язали його, але він розривав ланцюги та кайдани торощив, і ніхто не міг угамувати його.
MARK|5|5|І він повсякчас перебував день і ніч у гробах та в горах, і кричав, і бився об каміння...
MARK|5|6|А коли він Ісуса побачив здалека, то прибіг, і вклонився Йому,
MARK|5|7|і закричав гучним голосом, кажучи: Що до мене Тобі, Ісусе, Сину Бога Всевишнього? Богом Тебе заклинаю, не муч Ти мене!
MARK|5|8|Бо сказав Він йому: Вийди, душе нечистий, із людини!
MARK|5|9|І запитав Він його: Як тобі на ім'я? А той відповів: Леґіон мені ймення багато бо нас.
MARK|5|10|І він Його дуже просив, щоб їх не висилав із тієї землі.
MARK|5|11|Пасся ж там на горі гурт великий свиней.
MARK|5|12|І просилися демони, кажучи: Пошли нас у свиней, щоб у них ми ввійшли.
MARK|5|13|І дозволив Він їм. І повиходили духи нечисті, і в свиней увійшли. І гурт кинувся з кручі до моря, а було зо дві тисячі їх і вони потопилися в морі...
MARK|5|14|А їхні пастухи повтікали та в місті й по селах звістили. І повиходили люди побачити, що сталось.
MARK|5|15|І прийшли до Ісуса й побачили, що той біснуватий, що мав леґіона, убраний сидів, і при умі, і полякались вони...
MARK|5|16|Самовидці ж їм розповіли, що сталося з тим біснуватим, також про свиней.
MARK|5|17|І вони стали благати Його, щоб пішов Собі з їхнього краю.
MARK|5|18|А як Він сів до човна, то біснуватий став просити Його, щоб залишитися з Ним.
MARK|5|19|Ісус же йому не дозволив, а промовив до нього: Іди до дому свого, до своїх, і їм розповіж, які речі великі Господь учинив тобі, і як змилувався над тобою!
MARK|5|20|І пішов він та в Десятимісті зачав проповідувати, які речі великі Ісус учинив йому. І всі дивувались!
MARK|5|21|І коли переплив Ісус човном на той бік ізнов, то до Нього зібралось багато народу. І був Він над морем.
MARK|5|22|І приходить один із старших синагоги, на ймення Яір, і, як побачив Його, припадає до ніг Йому,
MARK|5|23|і дуже благає Його та говорить: Моя дочка кінчається. Прийди ж, поклади Свої руки на неї, щоб видужала та жила!...
MARK|5|24|І пішов Він із ним. За Ним натовп великий ішов, і тиснувсь до Нього.
MARK|5|25|А жінка одна, що дванадцять років хворою на кровотечу була,
MARK|5|26|що чимало натерпілася від багатьох лікарів, і витратила все добро своє, та ніякої помочі з того не мала, а прийшла ще до гіршого,
MARK|5|27|як зачула вона про Ісуса, підійшла через натовп іззаду, і доторкнулась до одежі Його...
MARK|5|28|Бо вона говорила про себе: Коли хоч доторкнусь до одежі Його, то одужаю...
MARK|5|29|І висохло хвилі тієї джерело кровотечі її, і тілом відчула вона, що видужала від недуги!
MARK|5|30|І в ту мить Ісус вичув у Собі, що вийшла з Нього сила. І Він до народу звернувся й спитав: Хто доторкнувсь до Моєї одежі?
MARK|5|31|І відказали Йому Його учні: Ти бачиш, що тисне на Тебе народ, а питаєшся: Хто доторкнувся до Мене?
MARK|5|32|А Він навкруги поглядав, щоб побачити ту, що зробила оце.
MARK|5|33|І жінка злякалась та затрусилась, бо знала, що сталося їй. І вона підійшла, і впала ницьма перед Ним, і всю правду Йому розповіла...
MARK|5|34|А Він їй сказав: Твоя віра, о дочко, спасла тебе; іди з миром, і здоровою будь від своєї недуги!
MARK|5|35|Як Він ще говорив, приходять ось від старшини синагоги та й кажуть: Дочка твоя вмерла; чого ще турбуєш Учителя?...
MARK|5|36|А Ісус, як почув слово сказане, промовляє до старшини синагоги: Не лякайсь, тільки віруй!
MARK|5|37|І Він не дозволив іти за Собою нікому, тільки Петрові та Якову, та Іванові, братові Якова.
MARK|5|38|І приходять у дім старшини синагоги, і Він бачить метушню та людей, що плакали та голосили.
MARK|5|39|А ввійшовши, сказав Він до них: Чого ви метушитеся та плачете? Не вмерло дівча, але спить!
MARK|5|40|І вони насміхалися з Нього. А Він усіх випровадив, узяв батька дівчати та матір, та тих, хто був із Ним, і ввійшов, де лежало дівча.
MARK|5|41|І взяв Він за руку дівча та й промовив до нього: Таліта, кумі що значить: Дівчатко, кажу тобі встань!
MARK|5|42|І в ту мить підвелося й ходило дівча; а років мало з дванадцять. І всі зараз жахнулися з дива великого!...
MARK|5|43|А Він наказав їм суворо, щоб ніхто не довідавсь про це. І дати їй їсти звелів.
MARK|6|1|І, вийшовши звідти, Він прийшов до Своєї батьківщини, а за Ним ішли учні Його.
MARK|6|2|Як настала ж субота, Він навчати почав у синагозі. І багато-хто, чувши, дивуватися стали й питали: Звідки в Нього оце? І що за мудрість, що дана Йому? І що за чуда, що стаються руками Його?
MARK|6|3|Хіба ж Він не тесля, син Маріїн, брат же Якову, і Йосипу, і Юді та Симонові? А сестри Його хіба тут не між нами? І вони спокушалися Ним...
MARK|6|4|А Ісус їм сказав: Пророка нема без пошани, хіба тільки в вітчизні своїй, та в родині своїй, та в домі своїм.
MARK|6|5|І Він тут учинити не міг чуда жадного, тільки деяких хворих, руки поклавши на них, уздоровив.
MARK|6|6|І Він дивувавсь їх невірству. І ходив Він по селах навкруг та навчав.
MARK|6|7|І, закликавши Дванадцятьох, зачав їх по двох посилати, і владу їм дав над нечистими духами.
MARK|6|8|І звелів їм нічого в дорогу не брати, крім палиці тільки самої: ні торби, ні хліба, ані мідяків у свій черес,
MARK|6|9|а ходити в сандалях, і двох убрань не носити.
MARK|6|10|І промовив до них: Коли ви де ввійдете в дім, залишайтеся там, аж поки не вийдете звідти.
MARK|6|11|А як місто яке вас не прийме, і не послухають вас, то, виходячи звідти, обтрусіть порох, що в вас під ногами, на свідчення супроти них. Поправді кажу вам, легше буде Содому й Гоморрі дня судного, аніж місту тому!
MARK|6|12|І вийшли вони, і проповідували, щоб каялися.
MARK|6|13|І багато вигонили демонів, і оливою хворих багато намащували і вздоровляли.
MARK|6|14|І прочув про Ісуса цар Ірод, бо ім'я Його стало загально відоме, і сказав, що то Іван Христитель із мертвих воскрес, і тому творяться чуда від нього.
MARK|6|15|Інші впевняли, що Ілля Він, а знов інші казали, що пророк, або як один із пророків.
MARK|6|16|А Ірод, прочувши, сказав: Іван, якому я голову стяв був, оце він воскрес!
MARK|6|17|Той бо Ірод, пославши, схопив був Івана, і в в'язниці закув його, через Іродіяду, дружину брата свого Пилипа, бо він одружився був із нею.
MARK|6|18|Бо Іван казав Іродові: Не годиться тобі мати за дружину жінку брата свого!
MARK|6|19|А Іродіяда лютилась на нього, і хотіла йому смерть заподіяти, та не могла.
MARK|6|20|Бо Ірод боявся Івана, знавши, що він муж праведний і святий, і беріг його. І, його слухаючи, він дуже бентежився, але слухав його залюбки.
MARK|6|21|Та настав день догідний, коли дня народження Ірод справляв був бенкета вельможам своїм, і тисячникам, і галілейській старшині,
MARK|6|22|і коли прийшла дочка тієї Іродіяди, і танцювала, і сподобалася Іродові та присутнім із ним при столі, тоді цар промовив до дівчини: Проси в мене, чого хочеш, і дам я тобі!
MARK|6|23|І поклявся він їй: Чого тільки від мене попросиш, то дам я тобі, хоча б і півцарства мого!
MARK|6|24|Вона ж вийшла, і спиталася матері своєї: Чого маю просити? А та відказала: Голови Івана Христителя...
MARK|6|25|І зараз квапливо вернулась вона до царя, і просила, говорячи: Я хочу, щоб дав ти негайно мені на полумиску голову Івана Христителя!
MARK|6|26|І засмутився цар, але через клятву й з-за тих, що з ним були при столі, не схотів їй відмовити.
MARK|6|27|І цар зараз послав вояка, і звелів принести Іванову голову.
MARK|6|28|І пішов він, і стяв у в'язниці Івана, і приніс його голову на полумискові, і дівчаті віддав, а дівча віддало її своїй матері...
MARK|6|29|А коли його учні зачули, то прийшли, і взяли його тіло, і до гробу поклали його.
MARK|6|30|І посходилися до Ісуса апостоли, і розповіли Йому все, як багато зробили вони, і як багато навчили.
MARK|6|31|І сказав Він до них: Ідіть осібно самі до безлюдного місця, та трохи спочиньте. Бо багато народу приходило та відбувало, аж навіть не мали коли й поживитись.
MARK|6|32|І відпливли вони човном окремо до місця безлюдного.
MARK|6|33|І побачили їх, коли плинули, і багато-хто їх розпізнали. І пішки побігли туди з усіх міст, та й їх випередили.
MARK|6|34|І, як вийшов Ісус, Він побачив багато народу, і змилувався над ними, бо були, немов вівці, що не мають пастуха. І зачав їх багато навчати.
MARK|6|35|І, як минуло вже часу доволі, підійшли Його учні до Нього та й кажуть: Це місце безлюдне, а година вже пізня.
MARK|6|36|Відпусти їх, нехай підуть в осади та села близькі, і куплять собі чого їсти.
MARK|6|37|А Він відповів і сказав їм: Дайте їсти їм ви. Вони ж відказали Йому: Чи ми маємо піти та хліба купити на двісті динаріїв, і дати їм їсти?
MARK|6|38|А Він їх запитав: Скільки маєте хліба? Ідіть, побачте! І розізнавши, сказали: П'ять хлібів та дві рибі.
MARK|6|39|І звелів їм усіх на зеленій траві посадити один біля одного.
MARK|6|40|І розсілись рядами вони, по сто та по п'ятдесят.
MARK|6|41|І Він узяв п'ять хлібів та дві рибі, споглянув на небо, поблагословив, і поламав ті хліби, і дав учням, щоб клали перед ними, і дві рибі на всіх поділив.
MARK|6|42|І всі їли й наїлися!
MARK|6|43|А з кусків позосталих та з риб назбирали дванадцять повних кошів.
MARK|6|44|А тих, хто хліб споживав, було тисяч із п'ять чоловіка!
MARK|6|45|І зараз звелів Своїм учням до човна сідати, і на той бік поплинути до Віфсаїди, раніше Його, поки Сам Він відпустить народ.
MARK|6|46|І Він їх відпустив, та й пішов помолитись на гору.
MARK|6|47|А як вечір настав, човен був серед моря, а Він Сам один на землі.
MARK|6|48|Коли ж Він побачив, як вони веслуванням мордуються, бо вітер їм був супротивний, о четвертій сторожі вночі підійшов Він до них, по морю йдучи, і хотів їх минути.
MARK|6|49|А вони, як побачили, що йде Він по морю, подумали, що то мара, та й стали кричати,
MARK|6|50|бо Його всі побачили та налякались. А Він зараз до них обізвався й сказав їм: Будьте смілі, це Я, не лякайтесь!
MARK|6|51|І ввійшов Він у човен до них, і вітер затих. А вони здивувалися дуже в собі,
MARK|6|52|бо не зрозуміли чуда про хліби, бо серце їхнє було затверділе.
MARK|6|53|Перепливши ж вони, прибули в землю Генісаретську й причалили.
MARK|6|54|І, як вони повиходили з човна, люди зараз пізнали Його,
MARK|6|55|і порозбігались по всій тій околиці, і стали на ложах недужих приносити, де тільки прочули були, що Він є.
MARK|6|56|І куди тільки Він прибував до сіл, чи до міст, чи до осель, клали недужих на майданах, і благали Його, щоб могли доторкнутись хоч краю одежі Його. І хто тільки до Нього доторкувався, той був уздоровлений!
MARK|7|1|І зібрались до Нього фарисеї та деякі з книжників, які прибули із Єрусалиму,
MARK|7|2|і побачили, що деякі з учнів Його їли хліб руками нечистими, цебто невмитими.
MARK|7|3|Бо фарисеї й усі юдеї, зберігаючи передання старших, не їдять, як старанно не вимиють рук;
MARK|7|4|а вернувшися з ринку, вони ні їдять, поки не вмиються. Багато є й іншого, що вони прийняли, щоб додержувати: миття чаш, і глеків, і мідяного посуду.
MARK|7|5|І запитали Його фарисеї та книжники: Чому учні Твої не живуть за переданням старших, але хліб споживають руками нечистими?
MARK|7|6|А Він їм відказав: Добре пророкував про вас, лицемірів, Ісая, як написано: Оці люди устами шанують Мене, серце ж їхнє далеко від Мене...
MARK|7|7|Та однак надаремне шанують Мене, бо навчають наук людських заповідей.
MARK|7|8|Занехаявши заповідь Божу, передань людських ви тримаєтесь: обмиваєте глеки та чаші, і багато такого подібного й іншого робите ви.
MARK|7|9|І сказав Він до них: Спритно відкидаєте ви заповідь Божу, аби зберегти своє передання.
MARK|7|10|Бо Мойсей наказав: Шануй батька свого та матір свою, та: Хто злорічить на батька чи матір, нехай смертю помре.
MARK|7|11|А ви кажете: Коли скаже хто батьку чи матері: Корван, чи дар Богові те, чим би ти скористатись від мене хотів,
MARK|7|12|то вже вільно йому не робити нічого для батька чи матері,
MARK|7|13|порушуючи Боже Слово вашим переданням, що його ви самі встановили. І багато такого ви іншого робите.
MARK|7|14|І Він знову покликав народ і промовив до нього: Послухайте Мене всі, і зрозумійте!
MARK|7|15|Немає нічого назовні людини, що, увіходячи в неї, могло б опоганити її; що ж із неї виходить, те людину опоганює.
MARK|7|16|Коли має хто вуха, щоб слухати, нехай слухає!
MARK|7|17|А коли від народу ввійшов Він до дому, тоді учні Його запиталися в Нього про притчу.
MARK|7|18|І Він їм відказав: Чи ж і ви розуміння не маєте? Хіба ж не розумієте ви, що все те, що входить іззовні в людину, не може опоганити її?
MARK|7|19|Бо не входить до серця йому, але до живота, і виходить назовні, очищуючи всяку їжу.
MARK|7|20|А далі сказав Він: Що з людини виходить, те людину опоганює.
MARK|7|21|Бо зсередини, із людського серця виходять лихі думки, розпуста, крадіж, душогубства,
MARK|7|22|перелюби, здирства, лукавства, підступ, безстидства, завидющеє око, богозневага, гордощі, безум.
MARK|7|23|Усе зле це виходить зсередини, і людину опоганює!
MARK|7|24|І встав Він, і звідти пішов у землю тирську й сидонську. І, ввійшовши до дому, Він хотів, щоб ніхто не довідавсь, та не міг утаїтись.
MARK|7|25|Негайно бо жінка одна, якої дочка мала духа нечистого, прочула про Нього, і прийшла, та й припала до ніг Йому.
MARK|7|26|А ця жінка грекиня була, родом сирофінікіянка. Вона стала благати Його, щоб із дочки її демона вигнав.
MARK|7|27|А Він їй сказав: Дай, щоб перше наїлися діти, не годиться бо хліб забирати в дітей, і кинути щенятам!
MARK|7|28|А вона Йому в відповідь каже: Так, Господи! Але навіть щенята їдять під столом від дитячих кришок...
MARK|7|29|І Він їй сказав: За слово оце йди собі, демон вийшов із твоєї дочки!
MARK|7|30|А коли вона в дім свій вернулась, то знайшла, що дочка на постелі лежала, а демон вийшов із неї.
MARK|7|31|І вийшов Він знов із країв тирських і сидонських, і подався шляхом на Сидон над море Галілейське, через околиці Десятимістя.
MARK|7|32|І приводять до Нього глухого немову, і благають Його, щоб руку на нього поклав.
MARK|7|33|І взяв Він його від народу самого, і вклав пальці Свої йому в вуха, і, сплюнувши, доторкнувся його язика.
MARK|7|34|І, на небо споглянувши, Він зідхнув і промовив до нього: Еффата; цебто: Відкрийся!
MARK|7|35|І відкрилися вуха йому, і путо його язика розв'язалось негайно, і він став говорити виразно!
MARK|7|36|А Він їм звелів, щоб нікому цього не розповідали. Та що більше наказував їм, то ще більш розголошували.
MARK|7|37|І дуже всі дивувалися та говорили: Він добре все робить: глухим дає чути, а німим говорити!
MARK|8|1|Тими днями, коли було знову багато народу, а їсти не мали чого, покликав Він учнів Своїх та й промовив до них:
MARK|8|2|Жаль мені тих людей, що вже три дні зо Мною знаходяться, та їсти не мають чого.
MARK|8|3|А коли відпущу їх голодних до їхніх домівок, то ослабнуть у дорозі, бо деякі з них поприходили здалека.
MARK|8|4|І відказали Йому Його учні: Звідки зможе хто нагодувати їх хлібом отут у пустині?
MARK|8|5|А Він їх запитав: Скільки маєте хліба? Вони ж повідомили: Семеро.
MARK|8|6|Тоді Він народу звелів на землі посідати. І, взявши семеро хліба, віддавши подяку, Він поламав і дав учням Своїм, щоб роздати. А вони роздавали народові.
MARK|8|7|І мали вони трохи рибок; і Він їх поблагословив, і роздати звелів також їх.
MARK|8|8|І всі їли й наїлися, а з позосталих кусків сім кошів назбирали...
MARK|8|9|А їдців було тисяч з чотири!
MARK|8|10|І всів Він негайно до човна з Своїми учнями, та й прибув до землі Далманутської.
MARK|8|11|І вийшли фарисеї, і почали сперечатися з Ним, і, Його випробовуючи, хотіли від Нього ознаки із неба.
MARK|8|12|А Він тяжко зідхнув у Своїм дусі й промовив: Якої ознаки цей рід вимагає? Поправді кажу вам, що родові цьому ознака не буде дана!
MARK|8|13|І покинув Він їх, усів знову до човна, і на той бік відбув.
MARK|8|14|І забули вони взяти хліба, і крім одного буханця, у човні не мали з собою нічого.
MARK|8|15|А Він їм наказував та говорив: Стережіться уважливо фарисейської розчини й розчини Іродової!
MARK|8|16|Вони ж міркували й казали один до одного, що хліба не мають вони.
MARK|8|17|А Ісус, знавши те, промовляє до них: Чого ви міркуєте, що хліба не маєте? Чи ви ще не знаєте й не розумієте? Чи ще маєте серце своє затверділим?
MARK|8|18|Мавши очі не бачите, і мавши вуха не чуєте? І не пам'ятаєте,
MARK|8|19|коли п'ять хлібів Я ламав на п'ять тисяч, скільки повних кошів із кусків ви зібрали? Вони кажуть до Нього: Дванадцять.
MARK|8|20|А як сім на чотири тисячі, скільки кошиків повних з кусків ви зібрали? І відказують: Сім.
MARK|8|21|І сказав Він до них: Ви ще не розумієте?...
MARK|8|22|І приходять вони в Віфсаїду. І приводять до Нього сліпого, і благають Його, щоб доторкнувся до нього.
MARK|8|23|І взяв Він сліпого за руку, та й вивів його за село. І послинивши очі йому, поклав руки на нього, і питався його, чи що бачить.
MARK|8|24|І, зиркнувши, сказав той: Я бачу людей, які ходять, немов би дерева...
MARK|8|25|Потім знов Він поклав Свої руки на очі йому, і прозрів той, і одужав, і виразно став бачити все!
MARK|8|26|І послав Він додому його й наказав: До села й не заходь, і нікому в селі не розповідай!
MARK|8|27|Потому пішов Ісус й учні Його до сіл Кесарії Пилипової, а в дорозі питав Своїх учнів, говорячи їм: За кого Мене люди вважають?
MARK|8|28|Вони ж відповіли Йому, кажучи: За Івана Христителя, другі за Іллю, а інші за одного з пророків.
MARK|8|29|І Він запитав їх: А ви за кого Мене маєте? Петро Йому в відповідь каже: Ти Христос!
MARK|8|30|І Він заборонив їм, щоб нікому про Нього вони не казали!
MARK|8|31|І почав їх навчати, що Синові Людському треба багато страждати, і Його відцураються старші, і первосвященики, і книжники, і Він буде вбитий, але третього дня Він воскресне.
MARK|8|32|І те слово казав Він відкрито. А Петро узяв набік Його, і Йому став перечити.
MARK|8|33|А Він обернувся й поглянув на учнів Своїх, та й Петру докорив і сказав: Відступись, сатано, від Мене, бо думаєш ти не про Боже, а про людське!
MARK|8|34|І Він покликав народ із Своїми учнями, та й промовив до них: Коли хоче хто йти вслід за Мною, хай зречеться самого себе, і хай візьме свого хреста та й за Мною йде!
MARK|8|35|Бо хто хоче душу свою зберегти, той погубить її, а хто згубить душу свою ради Мене та Євангелії, той її збереже.
MARK|8|36|Яка ж користь людині, що здобуде ввесь світ, але душу свою занапастить?
MARK|8|37|Або що назамін дасть людина за душу свою?
MARK|8|38|Бо хто буде Мене та Моєї науки соромитися в роді цім перелюбнім та грішнім, того посоромиться також Син Людський, як прийде у славі Свого Отця з Анголами святими.
MARK|9|1|І сказав Він до них: Поправді кажу вам, що деякі з тут-о приявних не скуштують смерти, аж поки не бачитимуть Царства Божого, що прийшло воно в силі.
MARK|9|2|А через шість день забирає Ісус Петра, і Якова, і Івана, та й веде їх осібно на гору високу самих. І Він переобразивсь перед ними.
MARK|9|3|І стала одежа Його осяйна, дуже біла, як сніг, якої білильник не зміг би так вибілити на землі!
MARK|9|4|І з'явивсь їм Ілля та Мойсей, і розмовляли з Ісусом.
MARK|9|5|І озвався Петро та й сказав до Ісуса: Учителю, добре бути нам тут! Поставмо ж собі три шатрі: для Тебе одне, і одне для Мойсея, і одне для Іллі...
MARK|9|6|Бо не знав, що казати, бо були перелякані.
MARK|9|7|Та хмара ось їх заслонила, і голос почувся із хмари: Це Син Мій Улюблений, Його слухайтеся!
MARK|9|8|І зараз, звівши очі свої, вони вже нікого з собою не бачили, крім Самого Ісуса.
MARK|9|9|А коли з гори сходили, Він їм наказав, щоб нікому того не казали, що бачили, аж поки Син Людський із мертвих воскресне.
MARK|9|10|І вони заховали те слово в собі, сперечаючися, що то є: воскреснути з мертвих.
MARK|9|11|І вони запитали Його та сказали: Що це книжники кажуть, ніби треба Іллі перш прийти?
MARK|9|12|А Він відказав їм: Тож Ілля, коли прийде попереду, усе приготує. Та як же про Людського Сина написано, що мусить багато Він витерпіти, і буде зневажений?
MARK|9|13|Але вам кажу, що й Ілля був прийшов, та зробили йому, що тільки хотіли, як про нього написано...
MARK|9|14|А коли повернулись до учнів, коло них вони вгледіли безліч народу та книжників, що сперечалися з ними.
MARK|9|15|І негайно ввесь натовп, як побачив Його, сполохнувся із дива, і назустріч побіг, і став вітати Його.
MARK|9|16|І запитався Він їх: Про що сперечаєтесь з ними?
MARK|9|17|І Йому відповів один із натовпу: Учителю, привів я до Тебе ось сина свого, що духа німого він має.
MARK|9|18|А як він де схопить його, то об землю кидає ним, і він піну пускає й зубами скрегоче та сохне. Я казав Твоїм учням, щоб прогнали його, та вони не змогли.
MARK|9|19|А Він їм у відповідь каже: О, роде невірний, доки буду Я з вами? Доки вас Я терпітиму? Приведіть до Мене його!
MARK|9|20|І до Нього того привели. І як тільки побачив Його, то дух зараз затряс ним. А той, повалившись на землю, став качатися та заливатися піною...
MARK|9|21|І Він запитав його батька: Як давно йому сталося це? Той сказав: Із дитинства.
MARK|9|22|І почасту кидав він ним і в огонь, і до води, щоб його погубити. Але коли можеш що Ти, то змилуйсь над нами, і нам поможи!
MARK|9|23|Ісус же йому відказав: Щодо того твого коли можеш, то тому, хто вірує, все можливе!
MARK|9|24|Зараз батько хлоп'яти з слізьми закричав і сказав: Вірую, Господи, поможи недовірству моєму!
MARK|9|25|А Ісус, як побачив, що натовп збігається, то нечистому духові заказав, і сказав йому: Душе німий і глухий, тобі Я наказую: вийди з нього, і більше у нього не входь!
MARK|9|26|І, закричавши та міцно затрясши, той вийшов. І він став, немов мертвий, аж багато-хто стали казати, що помер він...
MARK|9|27|А Ісус узяв за руку його та й підвів його, і той устав.
MARK|9|28|Коли ж Він до дому прийшов, то учні питали Його самотою: Чому ми не могли його вигнати?
MARK|9|29|А Він їм сказав: Цей рід не виходить інакше, як тільки від молитви та посту.
MARK|9|30|І вони вийшли звідти, і проходили по Галілеї. А Він не хотів, щоб довідався хто.
MARK|9|31|Бо Він Своїх учнів навчав і казав їм: Людський Син буде виданий людям до рук, і вони Його вб'ють, але вбитий, воскресне Він третього дня!
MARK|9|32|Вони ж не зрозуміли цього слова, та боялись Його запитати.
MARK|9|33|І прибули вони в Капернаум. А як був Він у домі, то їх запитав: Про що міркували в дорозі?
MARK|9|34|І мовчали вони, сперечалися бо проміж себе в дорозі, хто найбільший.
MARK|9|35|А як сів, то покликав Він Дванадцятьох, і промовив до них: Коли хто бути першим бажає, нехай буде найменшим із усіх і слуга всім!
MARK|9|36|І взяв Він дитину, і поставив її серед них. І, обнявши її, Він промовив до них:
MARK|9|37|Коли хто в Ім'я Моє прийме одне з дітей таких, той приймає Мене. Хто ж приймає Мене, не Мене він приймає, а Того, Хто послав Мене!
MARK|9|38|Обізвався до нього Іван: Учителю, ми бачили одного чоловіка, який з нами не ходить, що виганяє Ім'ям Твоїм демонів; і ми заборонили йому, бо він із нами не ходить.
MARK|9|39|А Ісус відказав: Не забороняйте йому, бо немає такого, що Ім'ям Моїм чудо зробив би, і зміг би небаром лихословити Мене.
MARK|9|40|Хто бо не супроти нас, той за нас!
MARK|9|41|І коли хто напоїть вас кухлем води в Ім'я Моє ради того, що ви Христові, поправді кажу вам: той не згубить своєї нагороди!
MARK|9|42|Хто ж спокусить одного з малих цих, що вірять, то краще б такому було, коли б жорно млинове на шию йому почепити, та й кинути в море!
MARK|9|43|І коли рука твоя спокушає тебе, відітни її: краще тобі ввійти до життя одноруким, ніж з обома руками ввійти до геєнни, до огню невгасимого,
MARK|9|44|де їхній червяк не вмирає, і не гасне огонь.
MARK|9|45|І коли нога твоя спокушає тебе, відітни її: краще тобі ввійти до життя одноногим, ніж з обома ногами бути вкиненому до геєнни, до огню невгасимого,
MARK|9|46|де їхній червяк не вмирає, і не гасне огонь.
MARK|9|47|І коли твоє око тебе спокушає, вибери його: краще тобі однооким ввійти в Царство Боже, ніж з обома очима бути вкиненому до геєнни огненної,
MARK|9|48|де їхній червяк не вмирає, і не гасне огонь!
MARK|9|49|Бо посолиться кожен огнем, і кожна жертва посолиться сіллю.
MARK|9|50|Сіль добра річ. Коли ж сіль несолоною стане, чим поправити її? Майте сіль у собі, майте й мир між собою!
MARK|10|1|І, вийшовши звідти, Він приходить у землю Юдейську, на той бік Йордану. І знову зібралися юрби до Нього, і знов Він навчав їх, звичаєм Своїм.
MARK|10|2|І підійшли фарисеї й спитали, Його випробовуючи: Чи дозволено чоловікові дружину свою відпустити?
MARK|10|3|А Він відповів і сказав їм: Що Мойсей заповів вам?
MARK|10|4|Вони ж відказали: Мойсей заповів написати листа розводового, та й відпустити.
MARK|10|5|Ісус же промовив до них: То за ваше жорстокосердя він вам написав оцю заповідь.
MARK|10|6|Бог же з початку творіння створив чоловіком і жінкою їх.
MARK|10|7|Покине тому чоловік свого батька та матір,
MARK|10|8|і стануть обоє вони одним тілом, тим то немає вже двох, але одне тіло.
MARK|10|9|Тож, що Бог спарував, людина нехай не розлучує!
MARK|10|10|А вдома про це учні знов запитали Його.
MARK|10|11|І Він їм відказав: Хто дружину відпустить свою, та й одружиться з іншою, той чинить перелюб із нею.
MARK|10|12|І коли дружина покине свого чоловіка, і вийде заміж за іншого, то чинить перелюб вона.
MARK|10|13|Тоді поприносили діток до Нього, щоб Він доторкнувся до них, учні ж їм докоряли.
MARK|10|14|А коли спостеріг це Ісус, то обурився, та й промовив до них: Пустіть діток до Мене приходити, і не бороніть їм, бо таких Царство Боже!
MARK|10|15|Поправді кажу вам: Хто Божого Царства не прийме, немов те дитя, той у нього не ввійде.
MARK|10|16|І Він їх пригорнув, і поблагословив, на них руки поклавши.
MARK|10|17|І коли вирушав Він у путь, то швидко наблизивсь один, упав перед Ним на коліна, і спитався Його: Учителю Добрий, що робити мені, щоб вічне життя вспадкувати?
MARK|10|18|Ісус же йому відказав: Чого звеш Мене Добрим? Ніхто не є Добрий, крім Бога Самого.
MARK|10|19|Знаєш заповіді: Не вбивай, не чини перелюбу, не кради, не свідкуй неправдиво, не кривди, шануй свого батька та матір.
MARK|10|20|А він відказав Йому: Учителю, це все виконав я ще змалку.
MARK|10|21|Ісус же поглянув на нього з любов'ю, і промовив йому: Одного бракує тобі: іди, розпродай, що маєш, та вбогим роздай, і матимеш скарб ти на небі! Потому приходь та й іди вслід за Мною, узявши хреста.
MARK|10|22|А він засмутився тим словом, і пішов, зажурившись, бо великі маєтки він мав!
MARK|10|23|І поглянув довкола Ісус, та й сказав Своїм учням: Як тяжко отим, хто має багатство, увійти в Царство Боже!
MARK|10|24|І учні жахнулись від слів Його. А Ісус знов у відповідь каже до них: Мої діти, як тяжко отим, хто надію кладе на багатство, увійти в Царство Боже!
MARK|10|25|Верблюдові легше пройти через голчине вушко, ніж багатому в Божеє Царство ввійти!
MARK|10|26|А вони здивувалися дуже, і казали один до одного: Хто ж тоді може спастися?
MARK|10|27|Ісус же поглянув на них і промовив: Неможливе це людям, а не Богові. Бо для Бога можливе все!
MARK|10|28|А Петро став казати Йому: От усе ми покинули, та й пішли за Тобою слідом.
MARK|10|29|Ісус відказав: Поправді кажу вам: Немає такого, щоб дім полишив, чи братів, чи сестер, або матір, чи батька, або діти, чи поля ради Мене та ради Євангелії,
MARK|10|30|і не одержав би в сто раз більше тепер, цього часу, серед переслідувань, домів, і братів, і сестер, і матерів, і дітей, і піль, а в віці наступному вічне життя.
MARK|10|31|І багато-хто з перших стануть останніми, а останні першими.
MARK|10|32|Були ж у дорозі вони, простуючи в Єрусалим. А Ісус ішов попереду них, аж дуже вони дивувались, а ті, що йшли вслід за Ним, боялись. І, взявши знов Дванадцятьох, почав їм розповідати, що з Ним статися має:
MARK|10|33|Оце в Єрусалим ми йдемо, і первосвященикам і книжникам виданий буде Син Людський, і засудять на смерть Його, і поганам Його видадуть,
MARK|10|34|і насміхатися будуть із Нього, і будуть плювати на Нього, і будуть Його бичувати, і вб'ють, але третього дня Він воскресне!
MARK|10|35|І підходять до Нього Яків та Іван, сини Зеведеєві, та й кажуть Йому: Учителю, ми хочемо, щоб Ти зробив нам, про що будемо просити Тебе.
MARK|10|36|А Він їх поспитав: Чого ж хочете, щоб Я вам зробив?
MARK|10|37|Вони ж відказали Йому: Дай нам, щоб у славі Твоїй ми сиділи праворуч від Тебе один, і ліворуч один!
MARK|10|38|А Ісус відказав їм: Не знаєте, чого просите. Чи ж можете ви пити чашу, що Я її п'ю, і христитися хрищенням, що Я ним хрищуся?
MARK|10|39|Вони відказали Йому: Можемо. А Ісус їм сказав: Чашу, що Я її п'ю, ви питимете, і хрищенням, що Я ним хрищусь, ви охриститеся.
MARK|10|40|А сидіти праворуч Мене та ліворуч не Моє це давати, а кому уготовано.
MARK|10|41|Як почули ж це Десятеро, то обурились на Якова та на Івана.
MARK|10|42|А Ісус їх покликав, і промовив до них: Ви знаєте, що ті, що вважають себе за князів у народів, панують над ними, а їхні вельможі їх тиснуть.
MARK|10|43|Не так буде між вами, але хто з вас великим бути хоче, нехай буде він вам за слугу.
MARK|10|44|А хто з вас бути першим бажає, нехай буде всім за раба.
MARK|10|45|Бо Син Людський прийшов не на те, щоб служили Йому, але щоб послужити, і душу Свою дати на викуп за багатьох.
MARK|10|46|І приходять вони в Єрихон. А коли з Єрихону виходив Він разом із Своїми учнями й з безліччю люду, сидів і просив при дорозі сліпий Вартимей, син Тимеїв.
MARK|10|47|І, прочувши, що то Ісус Назарянин, почав кликати та говорити: Сину Давидів, Ісусе, змилуйся надо мною!
MARK|10|48|І сварились на нього багато-хто, щоб мовчав, а він іще більше кричав: Сину Давидів, змилуйся надо мною!
MARK|10|49|І спинився Ісус та й сказав: Покличте його! І кличуть сліпого та й кажуть йому: Будь бадьорий, устань, Він кличе тебе.
MARK|10|50|А той скинув плаща свого, і скочив із місця, і прибіг до Ісуса.
MARK|10|51|А Ісус відповів і сказав йому: Що ти хочеш, щоб зробив Я тобі? Сліпий же Йому відказав: Учителю, нехай я прозрю!
MARK|10|52|Ісус же до нього промовив: Іди, твоя віра спасла тебе! І той зараз прозрів, і пішов за Ісусом дорогою.
MARK|11|1|І коли вони наблизились до Єрусалиму, до Вітфагії й Віфанії, на Оливній горі, тоді Він посилає двох учнів Своїх,
MARK|11|2|і каже до них: Ідіть у село, яке перед вами, і, входячи в нього, ви знайдете зараз прив'язане осля, що на нього ніхто ще з людей не сідав. Відв'яжіть його, і приведіть.
MARK|11|3|Коли ж скаже хто вам: Що це ви робите? відкажіть: Господь потребує його, і відішле його сюди зараз.
MARK|11|4|І вони відійшли, і знайшли те осля, що прив'язане коло воріт ізнадвору було при дорозі, і відв'язали його.
MARK|11|5|А деякі з тих, що стояли там, сказали до них: Що ви робите? Пощо осля ви відв'язуєте?
MARK|11|6|Вони ж їм відказали, як звелів їм Ісус, і відпущено їх.
MARK|11|7|І вони привели до Ісуса осля, і поклали на нього плащі свої, а Він сів на нього.
MARK|11|8|Багато ж народу стелили одежу свою по дорозі, а інші стелили дорогою зелень, натяту в полях.
MARK|11|9|А ті, що йшли перед Ним і позаду, викрикували: Осанна! Благословенний, хто йде у Господнє Ім'я!
MARK|11|10|Благословенне Царство, що надходить, Отця нашого Давида! Осанна на висоті!
MARK|11|11|Потому ввійшов Він до Єрусалиму, і в храм. А оглянувши все, як година вже пізня була, Він пішов у Віфанію з Дванадцятьма.
MARK|11|12|А назавтра, коли вони вийшли з Віфанії, Він зголоднів був.
MARK|11|13|І, побачивши здалека фіґове дерево, вкрите листями, Він підійшов, чи не знайде на ньому чого. І, прийшовши до нього, не знайшов нічого, крім листя самого, не пора бо на фіґи була.
MARK|11|14|І озвався Ісус і промовив до нього: Щоб більше ніхто твого плоду не з'їв аж повіки! А учні Його все те чули.
MARK|11|15|І прийшли вони в Єрусалим. А як Він у храм увійшов, то став виганяти продавців і покупців у храмі, і поперевертав столи грошомінам та ослони продавцям голубів.
MARK|11|16|І Він не дозволяв, щоб хто річ яку носив через храм.
MARK|11|17|І Він їх навчав і казав їм: Хіба не написано: Дім Мій буде домом молитви в народів усіх, ви ж із нього зробили печеру розбійників!
MARK|11|18|І почули це первосвященики й книжники, і шукали, як Його погубити, бо боялись Його, увесь бо народ дивувався науці Його.
MARK|11|19|А як пізно ставало, вони поза місто виходили.
MARK|11|20|А проходячи вранці, побачили фіґове дерево, усохле від кореня.
MARK|11|21|І, згадавши Петро, говорить Йому: Учителю, глянь фіґове дерево, що прокляв Ти, усохло!
MARK|11|22|А Ісус їм у відповідь каже: Майте віру Божу!
MARK|11|23|Поправді кажу вам: Як хто скаже горі цій: Порушся та й кинься до моря, і не матиме сумніву в серці своїм, але матиме віру, що станеться так, як говорить, то буде йому!
MARK|11|24|Через це говорю вам: Усе, чого ви в молитві попросите, вірте, що одержите, і сповниться вам.
MARK|11|25|І коли стоїте на молитві, то прощайте, як маєте що проти кого, щоб і Отець ваш Небесний пробачив вам прогріхи ваші.
MARK|11|26|Коли ж не прощаєте ви, то й Отець ваш Небесний не простить вам прогріхів ваших.
MARK|11|27|І знову прийшли вони в Єрусалим. Коли ж Він у храмі ходив, поприходили первосвященики й книжники, і старшини до Нього,
MARK|11|28|і сказали Йому: Якою Ти владою все оце чиниш? І хто Тобі владу цю дав, щоб Ти це робив?
MARK|11|29|А Ісус відказав їм: Запитаю й Я вас одне слово, і відповідайте Мені, то й Я відкажу вам, якою Я владою це все чиню.
MARK|11|30|Іванове хрищення з неба було, чи від людей? Відповідайте Мені!
MARK|11|31|Вони ж міркували собі й говорили: Коли скажемо: Із неба, відкаже: Чого ж ви йому не повірили?
MARK|11|32|А як скажемо: Від людей, то боялись народу, бо всі вважали, що Іван був поправді пророк.
MARK|11|33|І сказали Ісусові в відповідь: Не знаємо... А Ісус їм відказує: То й Я не скажу вам, якою Я владою це все чиню.
MARK|12|1|І почав Він у притчах до них промовляти: Насадив був один чоловік виноградника, муром обгородив, видовбав у ньому чавило, башту поставив, і віддав його винарям, та й пішов.
MARK|12|2|А певного часу послав він раба до своїх винарів, щоб прийняти частину плоду з виноградника в тих винарів.
MARK|12|3|Та вони схопили його та й побили, і відіслали ні з чим.
MARK|12|4|І знову послав він до них раба іншого, та й того вони зранили в голову та зневажили.
MARK|12|5|Тоді вислав він іншого, і того вони вбили. І багатьох іще інших, набили одних, а одних повбивали.
MARK|12|6|І він мав ще одного, сина улюбленого. Наостанок послав і того він до них і сказав: Посоромляться сина мого!
MARK|12|7|А ті винарі міркували собі: Це спадкоємець; ходім, замордуймо його, і нашою спадщина буде!
MARK|12|8|І вони схопили його та й убили, і викинули його за виноградник...
MARK|12|9|Отож, що пан виноградника зробить? Він прибуде та й вигубить тих винарів, і віддасть виноградника іншим.
MARK|12|10|Чи ви не читали в Писанні: Камінь, що його будівничі відкинули, той наріжним став каменем!
MARK|12|11|Від Господа сталося це, і дивне воно в очах наших.
MARK|12|12|І шукали Його, щоб схопити, але побоялись народу. Бо вони зрозуміли, що про них Він цю притчу сказав. І, лишивши Його, відійшли.
MARK|12|13|І вони вислали деяких із фарисеїв та іродіянів до Нього, щоб зловити на слові Його.
MARK|12|14|Ті ж прийшли та й говорять Йому: Учителю, знаємо ми, що Ти справедливий, і не зважаєш зовсім ні на кого, бо на людське обличчя не дивишся, а наставляєш на Божу дорогу правдиво. Чи годиться давати податок для кесаря, чи ні? Давати нам, чи не давати?
MARK|12|15|А Ісус, знавши їх лицемірство, сказав їм: Чого ви Мене випробовуєте? Принесіть Мені гріш податковий, щоб бачити.
MARK|12|16|І принесли вони. А Він каже до них: Чий це образ і напис? Ті ж Йому відказали: Кесарів.
MARK|12|17|Ісус тоді каже в відповідь їм: Віддайте кесареве кесареві, а Богові Боже! І дивувалися з Нього вони...
MARK|12|18|І прийшли до Нього ті саддукеї, що твердять, ніби нема воскресення, і запитали Його та сказали:
MARK|12|19|Учителю, Мойсей написав нам: Як помре кому брат, і полишить дружину, а дитини не лишить, то нехай його брат візьме дружину його, та й відновить насіння для брата свого.
MARK|12|20|Було сім братів. І перший взяв дружину й умер, не лишивши дітей.
MARK|12|21|Другий теж її взяв та й помер, і він не лишив дітей. Так само і третій.
MARK|12|22|І всі семеро не полишили дітей. А по всіх вмерла й жінка.
MARK|12|23|А в воскресенні, як воскреснуть вони, то котрому із них вона дружиною буде? Бо семеро мали за дружину її.
MARK|12|24|Ісус їм відказав: Чи ви не тому помиляєтесь, що не знаєте ані Писання, ані Божої сили?
MARK|12|25|Бо як із мертвих воскреснуть, то не будуть женитись, ані заміж виходити, але будуть, немов Анголи ті на небі.
MARK|12|26|Щождо мертвих, що воскреснуть, чи ж ви не читали в Мойсеєвій книзі, як при кущі сказав йому Бог, промовляючи: Я Бог Авраамів, і Бог Ісаків, і Бог Яковів,
MARK|12|27|Бо Він є Бог не мертвих, а живих! Тим то ви помиляєтесь дуже.
MARK|12|28|А один із тих книжників, що чув, як вони сперечались, та бачив, як добре Він відповідав їм, приступив та й спитався Його: Котра заповідь перша з усіх?
MARK|12|29|Ісус відповів: Перша: Слухай, Ізраїлю: наш Господь Бог Бог єдиний.
MARK|12|30|І: Люби Господа, Бога свого, усім серцем своїм, і всією душею своєю, і всім своїм розумом, і з цілої сили своєї! Це заповідь перша!
MARK|12|31|А друга однакова з нею: Люби свого ближнього, як самого себе! Нема іншої більшої заповіді над оці!
MARK|12|32|І сказав Йому книжник: Добре, Учителю! Ти поправді сказав, що Один Він, і нема іншого, окрім Нього,
MARK|12|33|і що Любити Його всім серцем, і всім розумом, і всією душею, і з цілої сили, і що Любити свого ближнього, як самого себе, це важливіше за всі цілопалення й жертви!
MARK|12|34|Ісус же, побачивши, що розумно той відповідь дав, промовив до нього: Ти недалеко від Божого Царства! І ніхто не насмілювався вже питати Його.
MARK|12|35|Потому Ісус відповів і промовив, у храмі навчаючи: Як то книжники кажуть, що ніби Христос син Давидів?
MARK|12|36|Адже той Давид Святим Духом сказав: Промовив Господь Господеві моєму: сядь праворуч Мене, доки не покладу Я Твоїх ворогів підніжком ногам Твоїм!
MARK|12|37|Сам Давид Його Господом зве, як же Він йому син? І багато людей залюбки Його слухали.
MARK|12|38|Він же казав у науці Своїй: Стережіться тих книжників, що люблять у довгих одежах проходжуватись, і привіти на ринках,
MARK|12|39|і перші лавки в синагогах, і перші місця на прийняттях,
MARK|12|40|що вдовині хати поїдають, і моляться довго напоказ, вони тяжче осудження приймуть!
MARK|12|41|І сів Він навпроти скарбниці, і дививсь, як народ мідяки до скарбниці вкидає. І багато заможних укидали багато.
MARK|12|42|І підійшла одна вбога вдовиця, і поклала дві лепті, цебто гріш.
MARK|12|43|І покликав Він учнів Своїх та й промовив до них: Поправді кажу вам, що ця вбога вдовиця поклала найбільше за всіх, хто клав у скарбницю.
MARK|12|44|Бо всі клали від лишка свого, а вона поклала з убозтва свого все, що мала, свій прожиток увесь...
MARK|13|1|І коли Він виходив із храму, говорить Йому один із учнів Його: Подивися, Учителю яке то каміння та що за будівлі!
MARK|13|2|Ісус же до нього сказав: Чи ти бачиш великі будинки оці? Не залишиться тут навіть камінь на камені, який не зруйнується!
MARK|13|3|Коли ж Він сидів на Оливній горі, проти храму, питали Його насамоті Петро, і Яків, і Іван, і Андрій:
MARK|13|4|Скажи нам, коли станеться це? І яка буде ознака, коли все те виконатись має?
MARK|13|5|Ісус же почав промовляти до них: Стережіться, щоб вас хто не звів.
MARK|13|6|Бо багато-хто прийдуть в Ім'я Моє, кажучи: Це Я. І зведуть багатьох.
MARK|13|7|І як про війни почуєте ви, і про воєнні чутки, не лякайтесь, бо статись належить тому. Та це ще не кінець.
MARK|13|8|Бо повстане народ на народ, і царство на царство, будуть землетруси місцями, буде голод. Це початок терпінь породільних.
MARK|13|9|Пильнуйте ж самі, бо вас на суди видаватимуть, і бичуватимуть вас у синагогах, і поведуть до правителів та до царів ради Мене, на свідчення їм.
MARK|13|10|Але перше Євангелія мусить бути народам усім проповідувана.
MARK|13|11|Коли ж видадуть вас і поведуть, не турбуйтеся заздалегідь, що вам говорити, а що дане вам буде тієї години, то те говоріть: бо не ви промовлятимете, але Дух Святий.
MARK|13|12|І видасть на смерть брата брат, а батько дитину. І діти повстануть навпроти батьків, і їм смерть заподіють.
MARK|13|13|І за Ім'я Моє будуть усі вас ненавидіти. А хто витерпить аж до кінця, той буде спасений!
MARK|13|14|Коли ж ви побачите ту гидоту спустошення, що про неї звіщав пророк Даниїл, що вона залягла, де не слід, хто читає, нехай розуміє, тоді ті, хто в Юдеї, нехай в гори втікають.
MARK|13|15|І хто на покрівлі, нехай той не сходить, і нехай не входить узяти щось із дому свого.
MARK|13|16|І хто на полі, хай назад не вертається взяти одежу свою.
MARK|13|17|Горе ж вагітним і тим, хто годує грудьми, у ті дні!
MARK|13|18|Моліться ж, щоб не трапилося це зимою!
MARK|13|19|Будуть бо ті дні такою скорботою, що її не було з первопочину світу, що його Бог створив, аж досі, і не буде.
MARK|13|20|І коли б Господь не вкоротив був тих днів, не спаслася б ніяка людина; але ради вибраних, кого вибрав, укоротив Він ті дні.
MARK|13|21|Тоді ж, як хто скаже до вас: Ото, Христос тут, Ото там, не йміть віри.
MARK|13|22|Бо повстануть христи неправдиві, і неправдиві пророки, і будуть чинити ознаки та чуда, щоб спокусити, як можна, і вибраних.
MARK|13|23|Але ви стережіться! Я сказав вам усе наперед.
MARK|13|24|Але за тих днів, по скорботі отій, сонце затьмиться, і місяць не дасть свого світла.
MARK|13|25|і зорі спадатимуть з неба, і сили небесні порушаться...
MARK|13|26|І побачать тоді Сина Людського, що йтиме на хмарах із великою потугою й славою.
MARK|13|27|І тоді Він пошле Анголів і зберуть Його вибраних від вітрів чотирьох, від краю землі до край-неба.
MARK|13|28|Від дерева ж фіґового навчіться прикладу: коли віття його вже розпукується, і кинеться листя, то знаєте, що близько літо.
MARK|13|29|Так і ви: коли тільки побачите, що діється це, то знайте, що близько, під дверима.
MARK|13|30|Поправді кажу вам: не перейде цей рід, аж усе оце станеться!
MARK|13|31|Небо й земля проминуться, але не минуться слова Мої!
MARK|13|32|Про день же той чи про годину не знає ніхто: ні Анголи на небі, ні Син, тільки Отець.
MARK|13|33|Уважайте, чувайте й моліться: бо не знаєте, коли час той настане!
MARK|13|34|Як той чоловік, що від'їхав, і залишив свій дім, і дав рабам своїм владу й кожному працю свою, а воротареві звелів пильнувати.
MARK|13|35|Тож пильнуйте, не знаєте бо, коли прийде пан дому: увечорі, чи опівночі, чи як півні співатимуть, чи ранком.
MARK|13|36|Щоб вас не застав, що спите, коли вернеться він несподівано.
MARK|13|37|А що вам Я кажу, те всім Я кажу: Пильнуйте!
MARK|14|1|За два ж дні була Пасха й Опрісноки. А первосвященики й книжники стали шукати, як би підступом взяти Його та забити.
MARK|14|2|Вони говорили: Та не в свято, щоб бува колотнеча в народі не сталась.
MARK|14|3|Коли ж Ісус був у Віфанії, у домі Симона, на проказу слабого, і сидів при столі, підійшла одна жінка, алябастрову пляшечку маючи щирого нардового дуже цінного мира. І розбила вона алябастрову пляшечку, і вилила миро на голову Йому!
MARK|14|4|А дехто обурювались між собою й казали: Нащо таке марнотратство на миро?
MARK|14|5|Бо можна було б це миро продати більше, як за три сотні динаріїв, і вбогим роздати. І нарікали на неї.
MARK|14|6|Ісус же сказав: Залишіть її! Чого прикрість їй робите? Вона добрий учинок зробила Мені.
MARK|14|7|Бо вбогих ви маєте завжди з собою, і коли схочете, можете їм робити добро, Мене ж не постійно ви маєте.
MARK|14|8|Що могла, те зробила вона: заздалегідь намастила Моє тіло на похорон...
MARK|14|9|Поправді кажу вам: де тільки ця Євангелія проповідувана буде в цілому світі, на пам'ятку їй буде сказане й те, що зробила вона!
MARK|14|10|Юда ж Іскаріотський, один із Дванадцятьох, подався до первосвящеників, щоб їм Його видати.
MARK|14|11|А вони, як почули, зраділи, і обіцяли йому срібняків за те дати. І він став вишукувати, як би слушного часу їм видати Його.
MARK|14|12|А першого дня Опрісноків, коли пасху приношено в жертву, сказали Йому Його учні: Куди хочеш, щоб пішли й приготували ми Тобі пасху спожити?
MARK|14|13|І посилає Він двох із Своїх учнів, і каже до них: Підіть до міста, і стріне вас чоловік, що нестиме в глекові воду, то йдіть за ним.
MARK|14|14|І там, куди він увійде, скажіть до господаря дому: Учитель питає: Де кімната Моя, в якій Я споживу зо Своїми учнями пасху?
MARK|14|15|І він вам покаже великую горницю, вистелену та готову: там приготуйте для нас.
MARK|14|16|І учні пішли, і до міста прийшли, і знайшли, як Він їм сказав, і зачали вони пасху готувати.
MARK|14|17|А коли настав вечір, Він приходить із Дванадцятьма.
MARK|14|18|І як сиділи вони при столі й споживали, промовив Ісус: Поправді кажу вам, що один з-поміж вас, який споживає зо Мною, видасть Мене...
MARK|14|19|Вони зачали сумувати, і один по одному питати Його: Чи не я?
MARK|14|20|А Він їм сказав: Один із Дванадцятьох, що в миску мачає зо Мною...
MARK|14|21|Людський Син справді йде, як про Нього написано; та горе тому чоловікові, що видасть він Людського Сина! Було б краще тому чоловікові, коли б він не родився!...
MARK|14|22|Як вони ж споживали, Ісус узяв хліб, і поблагословив, поламав, і дав їм, і сказав: Прийміть, споживайте, це тіло Моє!
MARK|14|23|І взяв Він чашу, і, вчинивши подяку, подав їм, і пили з неї всі.
MARK|14|24|І промовив до них: Це кров Моя Нового Заповіту, що за багатьох проливається.
MARK|14|25|Поправді кажу вам, що віднині не питиму Я від плоду виноградного до того дня, як новим буду пити його в Царстві Божім!
MARK|14|26|А коли відспівали вони, на гору Оливну пішли.
MARK|14|27|Промовляє тоді їм Ісус: Усі ви спокуситесь ночі цієї, як написано: Уражу пастиря, і розпорошаться вівці!
MARK|14|28|По воскресенні ж Своїм Я вас випереджу в Галілеї.
MARK|14|29|І відізвався до Нього Петро: Хоч спокусяться й усі, та не я!
MARK|14|30|Ісус же йому відказав: Поправді кажу тобі, що сьогодні, цієї ось ночі, перше ніж заспіває півень двічі, відречешся ти тричі від Мене!
MARK|14|31|А він ще сильніш запевняв: Коли б мені й умерти з Тобою, я не відречуся Тебе! Так же само сказали й усі...
MARK|14|32|І приходять вони до місцевости, на ім'я Гефсиманія, і каже Він учням Своїм: Посидьте ви тут, поки Я помолюся.
MARK|14|33|І, взявши з Собою Петра, і Якова та Івана, Він зачав сумувати й тужити...
MARK|14|34|І сказав Він до них: Обгорнена сумом смертельним душа Моя! Залишіться тут і пильнуйте!
MARK|14|35|І Він відійшов трохи далі, припав до землі, та й благав, щоб, як можна, минула Його ця година.
MARK|14|36|І благав Він: Авва-Отче, Тобі все можливе: пронеси мимо Мене цю чашу!... А проте, не чого хочу Я, але чого Ти...
MARK|14|37|І вернувся, і знайшов їх, що спали, та й каже Петрові: Симоне, спиш ти? Однієї години не зміг попильнувати?
MARK|14|38|Пильнуйте й моліться, щоб не впасти в спокусу, бадьорий бо дух, але немічне тіло!
MARK|14|39|І знову пішов і молився, те саме промовивши слово.
MARK|14|40|А вернувшись, ізнову знайшов їх, що спали, бо зважніли їм очі були. І не знали вони, що Йому відказати...
MARK|14|41|І вернувсь Він утретє, та й каже до них: Ви ще далі спите й спочиваєте? Скінчено, надійшла та година: у руки грішникам ось видається Син Людський!...
MARK|14|42|Уставайте, ходім, ось наблизивсь Мій зрадник...
MARK|14|43|І зараз, як Він ще говорив, прийшов Юда, один із Дванадцятьох, а з ним люди з мечами та киями від первосвящеників, і книжників, і старших.
MARK|14|44|А зрадник Його дав був знака їм, кажучи: Кого я поцілую, то Він, беріть Його, і обережно ведіть.
MARK|14|45|І, прийшовши, підійшов він негайно та й каже: Учителю! І поцілував Його...
MARK|14|46|Вони ж руки свої наклали на Нього, і схопили Його.
MARK|14|47|А один із тих, що стояли навколо, меча вихопив та й рубонув раба первосвященика, і відтяв йому вухо.
MARK|14|48|А Ісус їм промовив у відповідь: Немов на розбійника вийшли з мечами та киями, щоб узяти Мене.
MARK|14|49|Я щодня був із вами у храмі, навчаючи, і Мене не взяли ви. Але, щоб збулися Писання.
MARK|14|50|Тоді всі полишили Його й повтікали...
MARK|14|51|Один же юнак, по нагому загорнений у покривало, ішов услід за Ним. І хапають його.
MARK|14|52|Але він, покривало покинувши, утік нагий.
MARK|14|53|А Ісуса вони повели до первосвященика. І зійшлися всі первосвященики й старші та книжники.
MARK|14|54|Петро ж здалека йшов услід за Ним до середини двору первосвященика; і сидів він із службою, і грівсь при огні.
MARK|14|55|А первосвященики та ввесь синедріон шукали посвідчення на Ісуса, щоб Йому заподіяти смерть, і не знаходили.
MARK|14|56|Бо багато-хто свідчив фальшиво на Нього, але не було згідних свідчень.
MARK|14|57|Тоді деякі встали, і кривосвідчили супроти Нього й казали:
MARK|14|58|Ми чули, як Він говорив: Я зруйную цей храм рукотворний, і за три дні збудую інший, нерукотворний.
MARK|14|59|Але й так не було їхнє свідчення згідне.
MARK|14|60|Тоді встав насередині первосвященик, та й Ісуса спитав і сказав: Ти нічого не відповідаєш, що свідчать вони проти Тебе?
MARK|14|61|Він же мовчав, і нічого не відповідав. Первосвященик ізнову спитав Його, до Нього говорячи: Чи Христос Ти, Син Благословенного?
MARK|14|62|А Ісус відказав: Я! І побачите ви Сина Людського, що сидітиме по правиці сили Божої, і на хмарах небесних приходитиме!
MARK|14|63|Роздер тоді первосвященик одежу свою та й сказав: На що нам ще свідки потрібні?
MARK|14|64|Ви чули цю богозневагу. Як вам здається? Вони ж усі присудили, що Він умерти повинен...
MARK|14|65|Тоді деякі стали плювати на Нього, і закривати обличчя Йому, і бити Його та казати Йому: Пророкуй! Служба теж Його била по щоках...
MARK|14|66|А коли Петро був на подвір'ї надолі, приходить одна із служниць первосвященика,
MARK|14|67|і як Петра вона вгледіла, що грівся, подивилась на нього та й каже: І ти був із Ісусом Назарянином!
MARK|14|68|Він же відрікся, говорячи: Не відаю, і не розумію, що кажеш... І вийшов назовні, на переддвір'я. І заспівав тоді півень.
MARK|14|69|Служниця ж, коли його вгледіла, стала знов говорити приявним: Цей із них!
MARK|14|70|І він знову відрікся. Незабаром же знов говорили приявні Петрові: Поправді, ти з них, бо ти галілеянин. Та й мова твоя така сама.
MARK|14|71|А він став клястись та божитись: Не знаю Цього Чоловіка, про Якого говорите ви!
MARK|14|72|І заспівав півень хвилі тієї подруге. І згадав Петро слово, що Ісус був промовив йому: Перше ніж заспіває півень двічі, відречешся ти тричі від Мене. І кинувся він, та й плакати став...
MARK|15|1|А первосвященики з старшими й книжниками, та ввесь синедріон, зараз уранці, нараду вчинивши, зв'язали Ісуса, повели та й Пилатові видали.
MARK|15|2|А Пилат запитався Його: Чи Ти Цар Юдейський? А Він йому в відповідь каже: Сам ти кажеш...
MARK|15|3|А первосвященики міцно Його винуватили.
MARK|15|4|Тоді Пилат знову Його запитав і сказав: Ти нічого не відповідаєш? Дивись, як багато проти Тебе свідкують!
MARK|15|5|А Ісус більш нічого не відповідав, так що Пилат дивувався.
MARK|15|6|На свято ж він їм відпускав був одного із в'язнів, котрого просили вони.
MARK|15|7|Був же один, що звався Варавва, ув'язнений разом із повстанцями, які за повстання вчинили були душогубство.
MARK|15|8|Коли ж натовп зібрався, він став просити Пилата зробити, як він завжди робив їм.
MARK|15|9|Пилат же сказав їм у відповідь: Хочете, відпущу вам Царя Юдейського?
MARK|15|10|Бо він знав, що Його через заздрощі видали первосвященики.
MARK|15|11|А первосвященики натовп підмовили, щоб краще пустив їм Варавву.
MARK|15|12|Пилат же промовив ізнов їм у відповідь: А що ж я чинитиму з Тим, що Його ви Юдейським Царем називаєте?
MARK|15|13|Вони ж стали кричати знов: Розіпни Його!
MARK|15|14|Пилат же сказав їм: Яке ж зло вчинив Він? А вони ще сильніше кричали: Розіпни Його!...
MARK|15|15|Пилат же хотів догодити народові, і відпустив їм Варавву. І видав Ісуса, збичувавши, щоб розп'ятий був.
MARK|15|16|Вояки ж повели Його до середини двору, цебто в преторій, і цілий відділ скликають.
MARK|15|17|І вони зодягли Його в багряницю і, сплівши з тернини вінка, поклали на Нього.
MARK|15|18|І вітати Його зачали: Радій, Царю Юдейський!
MARK|15|19|І тростиною по голові Його били, і плювали на Нього. І навколішки кидалися та вклонялись Йому...
MARK|15|20|І коли назнущалися з Нього, зняли з Нього багряницю, і наділи на Нього одежу Його. І Його повели, щоб розп'ясти Його.
MARK|15|21|І одного перехожого, що з поля вертався, Симона Кірінеянина, батька Олександра та Руфа, змусили, щоб хреста Йому ніс.
MARK|15|22|І Його привели на місце Голгофу, що значить Череповище.
MARK|15|23|І давали Йому пити вина, із миррою змішаного, але Він не прийняв.
MARK|15|24|І Його розп'яли, і поділили одежу Його, кинувши жереб про неї, хто що візьме.
MARK|15|25|Була ж третя година, як Його розп'яли.
MARK|15|26|І був написаний напис провини Його: Цар Юдейський.
MARK|15|27|Тоді розп'ято з Ним двох розбійників, одного праворуч, і одного ліворуч Його.
MARK|15|28|І збулося Писання, що каже: До злочинців Його зараховано!
MARK|15|29|А хто побіч проходив, то Його лихословили, головами своїми хитали й казали: Отак! Ти, що храма руйнуєш та за три дні будуєш,
MARK|15|30|зійди із хреста, та спаси Самого Себе!
MARK|15|31|Теж і первосвященики з книжниками глузували й один до одного казали: Він інших спасав, а Самого Себе не може спасти!
MARK|15|32|Христос, Цар Ізраїлів, нехай зійде тепер із хреста, щоб побачили ми та й увірували. Навіть ті, що разом із Ним були розп'яті, насміхалися з Нього...
MARK|15|33|А як шоста година настала, то аж до години дев'ятої темрява стала по цілій землі.
MARK|15|34|О годині ж дев'ятій Ісус скрикнув голосом гучним та й вимовив: Елої, Елої, лама савахтані, що в перекладі значить: Боже Мій, Боже Мій, нащо Мене Ти покинув?
MARK|15|35|Дехто ж із тих, що стояли навколо, це почули й казали: Ось Він кличе Іллю!
MARK|15|36|А один із них побіг, намочив губку оцтом, настромив на тростину, і давав Йому пити й казав: Чекайте, побачим, чи прийде Ілля Його зняти!
MARK|15|37|А Ісус скрикнув голосом гучним, і духа віддав!...
MARK|15|38|І в храмі завіса роздерлась надвоє, від верху аж додолу.
MARK|15|39|А сотник, що насупроти Нього стояв, як побачив, що Він отак духа віддав, то промовив: Чоловік Цей був справді Син Божий!
MARK|15|40|Були ж і жінки, що дивились здалека, між ними Марія Магдалина, і Марія, мати Якова Молодшого та Йосії, і Саломія,
MARK|15|41|що вони, як Він був у Галілеї, ходили за Ним та Йому прислуговували; і інших багато, що до Єрусалиму прийшли з Ним.
MARK|15|42|А коли настав вечір, через те, що було Приготовлення, цебто перед суботою,
MARK|15|43|прийшов Йосип із Ариматеї, радник поважний, що сам сподівавсь Царства Божого, і сміливо ввійшов до Пилата, і просив тіла Ісусового.
MARK|15|44|А Пилат здивувався, щоб Він міг уже вмерти. І, покликавши сотника, запитався його, чи давно вже Розп'ятий помер.
MARK|15|45|І, дізнавшись від сотника, він подарував тіло Йосипові.
MARK|15|46|А Йосип купив плащаницю, і, знявши Його, обгорнув плащаницею, та й поклав Його в гробі, що в скелі був висічений. І каменя привалив до могильних дверей.
MARK|15|47|Марія ж Магдалина й Марія, мати Йосієва, дивилися, де ховали Його.
MARK|16|1|Як минула ж субота, Марія Магдалина, і Марія Яковова, і Саломія накупили пахощів, щоб піти й намастити Його.
MARK|16|2|І на світанку дня першого в тижні, як сходило сонце, до гробу вони прибули,
MARK|16|3|і говорили одна одній: Хто відвалить нам каменя від могильних дверей?
MARK|16|4|А зиркнувши, побачили, що камінь відвалений; був же він дуже великий...
MARK|16|5|І, ввійшовши до гробу, побачили там юнака, що праворуч сидів, і був одягнений в білу одежу, і жахнулись вони...
MARK|16|6|А він промовляє до них: Не жахайтесь! Ви шукаєте Розп'ятого, Ісуса Назарянина. Він воскрес, нема Його тут! Ось місце, де Його поховали були.
MARK|16|7|Але йдіть, скажіть учням Його та Петрові: Він іде в Галілею попереду вас, там Його ви побачите, як Він вам говорив.
MARK|16|8|А як вийшли вони, то побігли від гробу, бо їх трепет та страх обгорнув. І не сказали нікому нічого, бо боялись...
MARK|16|9|Як воскрес Він уранці дня першого в тижні, то з'явився найперше Марії Магдалині, із якої був вигнав сім демонів.
MARK|16|10|Пішовши вона, повідомила тих, що були з Ним, які сумували та плакали.
MARK|16|11|А вони, як почули, що живий Він, і вона Його бачила, не йняли тому віри.
MARK|16|12|По цьому з'явився Він двом із них у постаті іншій в дорозі, як ішли вони на село.
MARK|16|13|А вони, як вернулися, інших про те сповістили, але не повірено й їм.
MARK|16|14|Нарешті, Він з'явився Одинадцятьом, як сиділи вони при столі, і докоряв їм за недовірство їхнє та твердосердя, що вони не йняли віри тим, хто воскреслого бачив Його.
MARK|16|15|І казав Він до них: Ідіть по цілому світові, та всьому створінню Євангелію проповідуйте!
MARK|16|16|Хто увірує й охриститься, буде спасений, а хто не ввірує засуджений буде.
MARK|16|17|А тих, хто ввірує, супроводити будуть ознаки такі: у Ім'я Моє демонів будуть вигонити, говоритимуть мовами новими,
MARK|16|18|братимуть змій; а коли смертодійне що вип'ють, не буде їм шкодити; кластимуть руки на хворих, і добре їм буде!
MARK|16|19|Господь же Ісус, по розмові із ними, вознісся на небо, і сів по Божій правиці.
MARK|16|20|І пішли вони, і скрізь проповідували. А Господь помагав їм, і стверджував слово ознаками, що його супроводили. Амінь.
