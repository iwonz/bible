ROM|1|1|基督耶稣的仆人 保罗 ，蒙召为使徒，奉派传上帝的福音。
ROM|1|2|这福音是上帝从前藉众先知，在圣经上所应许的。
ROM|1|3|论到他儿子－我主耶稣基督，按肉体说，是从 大卫 后裔生的；按神圣的灵说，因从死人中复活，用大能显明他是上帝的儿子。
ROM|1|4|
ROM|1|5|我们从他蒙恩受了使徒的职分，为他的名在万国中使人因信而顺服，
ROM|1|6|其中也有你们这蒙召属耶稣基督的人。
ROM|1|7|我写信给你们在 罗马 、为上帝所爱、蒙召作圣徒的众人。愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
ROM|1|8|首先，我靠着耶稣基督，为你们众人感谢我的上帝，因你们的信德传遍了天下。
ROM|1|9|我在他儿子的福音上，用心灵所事奉的上帝可以见证，我怎样不住地提到你们，
ROM|1|10|在我的祷告中常常恳求，或许照上帝的旨意，最终我能毫无阻碍地往你们那里去。
ROM|1|11|因为我迫切地想见你们，要把一些属灵的恩赐分给你们，使你们得以坚固，
ROM|1|12|也可以说，我在你们中间，因你我彼此的信心而同得安慰。
ROM|1|13|弟兄们，我不愿意你们不知道，我屡次计划往你们那里去，要在你们中间得些果子，如同在其余的外邦人中一样，只是到如今仍有拦阻。
ROM|1|14|无论是 希腊 人、未开化的人、聪明人、愚拙人，我都欠他们的债，
ROM|1|15|所以愿意尽我的力量把福音也传给你们在 罗马 的人。
ROM|1|16|我不以福音为耻；这福音本是上帝的大能，要救一切相信的，先是 犹太 人，后是 希腊 人。
ROM|1|17|因为上帝的义正在这福音上显明出来；这义是本于信，以至于信。如经上所记：“义人必因信得生。”
ROM|1|18|原来，上帝的愤怒从天上显明在一切不虔不义的人身上，就是那些行不义压制真理的人。
ROM|1|19|上帝的事情，人所能知道的，原显明在人心里，因为上帝已经向他们显明。
ROM|1|20|自从造天地以来，上帝的永能和神性是明明可知的，虽然眼不能见，但藉着所造之物就可以了解看见，叫人无可推诿。
ROM|1|21|因为，他们虽然知道上帝，却不把他当作上帝荣耀他，也不感谢他。他们的思想变为虚妄，无知的心昏暗了。
ROM|1|22|他们自以为聪明，反成了愚昧，
ROM|1|23|将不能朽坏之上帝的荣耀变为偶像，仿照必朽坏的人、飞禽、走兽、爬虫的形像。
ROM|1|24|所以，上帝任凭他们随着心里的情欲行污秽的事，以致彼此羞辱自己的身体。
ROM|1|25|他们将上帝的真实变为虚谎，去敬拜事奉受造之物，不敬奉那造物的主—主是可称颂的，直到永远。阿们！
ROM|1|26|因此，上帝任凭他们放纵可羞耻的情欲。他们的女人把自然的关系变成违反自然的；
ROM|1|27|男人也是如此，放弃了和女人自然的关系，欲火攻心，男的和男的彼此贪恋，行可耻的事，就在自己身上受这逆性行为当得的报应。
ROM|1|28|他们既然故意不认识上帝，上帝就任凭他们存扭曲的心，做那些不该做的事，
ROM|1|29|装满了各样不义 、邪恶、贪婪、恶毒，满心是嫉妒、凶杀、纷争、诡诈、毒恨，又是毁谤的、
ROM|1|30|说人坏话的、怨恨上帝的 、侮辱人的、狂傲的、自夸的、制造是非的、忤逆父母的、
ROM|1|31|顽梗不化的、言而无信的、无情无义的、不怜悯人的。
ROM|1|32|他们虽知道上帝判定做这样事的人是该死的，然而他们不但自己去做，还赞同别人去做。
ROM|2|1|所以，你这评断人的人哪，无论你是谁，都无可推诿。你在什么事上评断人，就在什么事上定自己的罪。因你这评断人的，自己所做的却和别人一样。
ROM|2|2|我们知道这样做的人，上帝必公平地审判他。
ROM|2|3|你这个人哪，你评断做这样事的人，自己所做的却和别人一样，你以为能逃脱上帝的审判吗？
ROM|2|4|还是你藐视他丰富的恩慈、宽容、忍耐，不知道他的恩慈是领你悔改吗？
ROM|2|5|你竟放任你刚硬不悔改的心，为自己累积愤怒！在愤怒的日子，上帝公义的审判要显示出来。
ROM|2|6|他要照各人的行为报应各人。
ROM|2|7|凡恒心行善，寻求荣耀、尊贵和不能朽坏的，就有永生报偿他们；
ROM|2|8|但是那些自私自利、不顺从真理、反顺从不义的人，就有恼恨、愤怒报应他们。
ROM|2|9|他要把患难、困苦加给一切作恶的人，先是 犹太 人，后是 希腊 人；
ROM|2|10|却把荣耀、尊贵、平安加给一切行善的人，先是 犹太 人，后是 希腊 人。
ROM|2|11|因为上帝不偏待人。
ROM|2|12|凡在律法之外犯了罪的，将在律法之外灭亡；凡在律法之内犯了罪的，将按律法受审判。
ROM|2|13|原来在上帝面前，不是听律法的为义，而是行律法的称义。
ROM|2|14|没有律法的外邦人若顺着本性行律法上的事，他们虽然没有律法，自己就是自己的律法。
ROM|2|15|他们显明律法的功用刻在他们心里，他们的良心一同作证—他们的内心挣扎，有时自责，有时为自己辩护。
ROM|2|16|在那日，上帝要藉着基督耶稣 ，按照我所传的福音，审判人隐藏的事。
ROM|2|17|但是你，你既自称为 犹太 人，倚靠律法，以上帝夸口，
ROM|2|18|知道上帝的旨意，从律法受了教导而能分辨是非；
ROM|2|19|你既深信自己是给盲人领路的，是在黑暗中人的光，
ROM|2|20|是无知的人的师傅，是小孩子的老师，体现了律法中的知识和真理；
ROM|2|21|那么，你这教导别人的，还不教导自己吗？你这宣讲不可偷窃的，自己还偷窃吗？
ROM|2|22|你这说不可奸淫的，自己还奸淫吗？你这厌恶偶像的，自己还抢劫庙中之物吗？
ROM|2|23|你这以律法夸口的，自己倒违犯律法，羞辱上帝！
ROM|2|24|上帝的名在外邦人中因你们受了亵渎，正如经上所记的。
ROM|2|25|你若遵行律法，割礼固然于你有益；若违犯律法，你的割礼就算不得割礼。
ROM|2|26|所以，那未受割礼的，若遵守律法的要求，他虽然未受割礼，岂不算是受了割礼吗？
ROM|2|27|而且那本来未受割礼的，若能全守律法，岂不是要审判你这有仪文和割礼，竟违犯律法的人吗？
ROM|2|28|因为外表是 犹太 人的不是真 犹太 人；外表肉身的割礼也不是真割礼。
ROM|2|29|惟有内心作 犹太 人的才是真 犹太 人，真割礼也是心里的，在乎圣灵 ，不在乎仪文。这样的人所受的称赞不是从人来的，而是从上帝来的。
ROM|3|1|这样说来， 犹太 人有什么比别人强呢？割礼有什么益处呢？
ROM|3|2|很多，各方面都有。首先，上帝的圣言交托他们。
ROM|3|3|即使有不信的，这又何妨呢？难道他们的不信就废掉上帝的信实吗？
ROM|3|4|绝对不会！不如说，上帝是真实的，而人都是虚谎的。如经上所记： “以致你责备的时候显为公义； 你被指控的时候一定胜诉。”
ROM|3|5|我姑且照着人的看法来说，我们的不义若显出上帝的义来，我们要怎么说呢？上帝降怒是他不义吗？
ROM|3|6|绝对不是！若是这样，上帝怎能审判世界呢？
ROM|3|7|若上帝的真实因我的虚谎越发显出他的荣耀，为什么我还像罪人一样受审判呢？
ROM|3|8|为什么不说，我们可以作恶以成善呢？有人毁谤我们，说我们讲过这话；这等人被定罪是应该的。
ROM|3|9|那又怎么样呢？我们比他们强吗？绝不是！因我们已经指证： 犹太 人和 希腊 人都在罪恶之下。
ROM|3|10|就如经上所记： “没有义人，连一个也没有。
ROM|3|11|没有明白的， 没有寻求上帝的。
ROM|3|12|人人偏离正路，一同走向败坏。 没有行善的，连一个也没有 。
ROM|3|13|他们的喉咙是敞开的坟墓； 他们的舌头玩弄诡诈。 他们的嘴唇里有毒蛇的毒液，
ROM|3|14|满口是咒骂苦毒。
ROM|3|15|他们的脚为杀人流血飞跑；
ROM|3|16|他们的路留下毁坏和灾难。
ROM|3|17|和平的路，他们不认识；
ROM|3|18|他们眼中不怕上帝。”
ROM|3|19|我们知道律法所说的话都是对律法之下的人说的，好塞住各人的口，使普世的人都伏在上帝的审判之下。
ROM|3|20|所以，凡血肉之躯没有一个能因律法的行为而在上帝面前称义，因为律法本是要人认识罪。
ROM|3|21|但如今，上帝的义在律法之外已经显明出来，有律法和先知为证：
ROM|3|22|就是上帝的义，因信耶稣基督 加给一切信的人。这并没有分别，
ROM|3|23|因为世人都犯了罪，亏缺了上帝的荣耀，
ROM|3|24|如今却蒙上帝的恩典，藉着在基督耶稣里的救赎，就白白地得称为义。
ROM|3|25|上帝设立耶稣作赎罪祭，是凭耶稣的血，藉着信，要显明上帝的义；因为他用忍耐的心宽容人先前所犯的罪，好使今时显明他的义，让人知道他自己为义，也称信耶稣的人为义 。
ROM|3|26|
ROM|3|27|既是这样，哪里可夸口呢？没有可夸的。是藉什么法呢？功德吗？不是！是藉信主之法。
ROM|3|28|所以我们认定，人称义是因着信，不在于律法的行为。
ROM|3|29|难道上帝只是 犹太 人的吗？不也是外邦人的吗？是的，他也是外邦人的上帝。
ROM|3|30|既然上帝是一位，他就要本于信称那受割礼的为义，也要藉着信称那未受割礼的为义。
ROM|3|31|这样，我们藉着信废了律法吗？绝对不是！更是巩固律法。
ROM|4|1|这样，那按肉体作我们祖宗的 亚伯拉罕 ，我们要怎么说呢？
ROM|4|2|倘若 亚伯拉罕 是因行为称义，他就有可夸的，但是在上帝面前他一无可夸。
ROM|4|3|经上说什么呢？“ 亚伯拉罕 信了上帝，这就算他为义。”
ROM|4|4|做工的得工资不算是恩典，而是应得的；
ROM|4|5|但那不做工的，只信那位称不敬虔之人为义的，他的信就算为义。
ROM|4|6|正如 大卫 称那在行为之外蒙上帝算为义的人是有福的：
ROM|4|7|“过犯得赦免，罪恶蒙遮盖的人有福了！
ROM|4|8|主不算为有罪的，这样的人有福了！”
ROM|4|9|如此看来，这福只加给那受割礼的人吗？不也加给那未受割礼的人吗？我们说，因着信，就算 亚伯拉罕 为义。
ROM|4|10|那么，这是怎么算的呢？是在他受割礼的时候呢？还是在他未受割礼的时候呢？不是在受割礼的时候，而是在未受割礼的时候。
ROM|4|11|并且，他受了割礼的记号，作他未受割礼的时候因信称义的印证，为使他作一切未受割礼而信之人的父，使他们也算为义，
ROM|4|12|也使他作受割礼之人的父，就是那些不但受割礼，而且跟随我们的祖宗 亚伯拉罕 未受割礼而信的足迹的人。
ROM|4|13|因为上帝给 亚伯拉罕 和他后裔承受世界的应许不是藉着律法，而是藉着信而得的义。
ROM|4|14|若是属于律法的人才是后嗣，信就落空了，应许也就失效了。
ROM|4|15|因为律法是惹动愤怒的，哪里没有律法，哪里就没有过犯。
ROM|4|16|所以，人作后嗣是出于信，因此就属乎恩，以致应许保证归给所有的后裔，不但归给那属于律法的，也归给那效法 亚伯拉罕 之信的人。 亚伯拉罕 所信的是那叫死人复活、使无变为有的上帝，在这位上帝面前 亚伯拉罕 成为我们众人的父，如经上所记：“我已经立你作多国之父。”
ROM|4|17|
ROM|4|18|他在没有盼望的时候，仍存着盼望来相信，就得以作多国之父，正如先前所说：“你的后裔将要如此。”
ROM|4|19|他将近百岁的时候，虽然想到 自己的身体如同已死， 撒拉 也不可能生育，他的信心还是不软弱，
ROM|4|20|仍仰望上帝的应许，总没有因不信而起疑惑，反倒因信而刚强，将荣耀归给上帝，
ROM|4|21|且满心相信上帝所应许的必能成就。
ROM|4|22|所以这也 就算他为义。
ROM|4|23|“算他为义”这句话不是单为他写的，
ROM|4|24|也是为我们将来得算为义的人写的，就是为我们这些信上帝使我们的主耶稣从死人中复活的人写的。
ROM|4|25|耶稣被出卖，是为我们的过犯；他复活，是为使我们称义。
ROM|5|1|所以，我们既因信称义，就藉着我们的主耶稣基督得以与上帝和好。
ROM|5|2|我们又藉着他，因信 得以进入现在所站立的这恩典中，并且欢欢喜喜盼望上帝的荣耀。
ROM|5|3|不但如此，就是在患难中也是欢欢喜喜的，因为知道患难生忍耐，
ROM|5|4|忍耐生老练，老练生盼望，
ROM|5|5|盼望不至于落空，因为上帝的爱，已藉着所赐给我们的圣灵，浇灌在我们心里。
ROM|5|6|我们还软弱的时候，基督就在特定的时刻为不敬虔之人死。
ROM|5|7|为义人死，是少有的；为仁人死，或者有敢做的。
ROM|5|8|惟有基督在我们还作罪人的时候为我们死，上帝的爱就在此向我们显明了。
ROM|5|9|现在我们既靠着他的血称义，就更要藉着他得救，免受上帝的愤怒。
ROM|5|10|因为我们作仇敌的时候，尚且藉着上帝儿子的死得以与上帝和好，既已和好，就更要因他的生得救了。
ROM|5|11|不但如此，我们既藉着我们的主耶稣基督得以与上帝和好，也就藉着他以上帝为乐。
ROM|5|12|为此，正如罪是从一人进入世界，死又从罪而来，于是死就临到所有的人，因为人人都犯了罪。
ROM|5|13|没有律法之前，罪已经在世上，但没有律法，罪也不算罪。
ROM|5|14|然而，从 亚当 到 摩西 ，死就掌了权，连那些不与 亚当 犯一样罪过的，也在死的权下。 亚当 是那以后要来之人的预像。
ROM|5|15|但是过犯不如恩赐，若因一人的过犯，众人都死了，那么，上帝的恩典，与那因耶稣基督一人而来的恩典中的赏赐，岂不加倍地临到众人吗？
ROM|5|16|因一人犯罪而来的后果，也不如赏赐，原来审判是由一人而定罪，恩赐乃是由许多过犯而称义。
ROM|5|17|若因一人的过犯，死就因这一人掌权，那些受洪恩又蒙所赐之义的，岂不更要因耶稣基督一人在他们生命中掌权吗？
ROM|5|18|这样看来，因一次的过犯，所有的人都被定罪；照样，因一次的义行，所有的人也就被称义而得生命了。
ROM|5|19|因一人的悖逆，众人成为罪人；照样，因一人的顺从，众人也成为义了。
ROM|5|20|而且加添了律法，使得过犯增加，只是罪在哪里增加，恩典就在哪里越发丰盛了。
ROM|5|21|所以，正如罪藉着死掌权；照样，恩典也藉着义掌权，使人因我们的主耶稣基督得永生。
ROM|6|1|这样，我们要怎么说呢？我们可以仍在罪中使恩典增多吗？
ROM|6|2|绝对不可！我们向罪死了的人，岂可仍在罪中活着呢？
ROM|6|3|难道你们不知道，我们这受洗归入基督耶稣的人，就是受洗归入他的死吗？
ROM|6|4|所以，我们藉着洗礼归入死，和他一同埋葬，是要我们行事为人都有新生的样子，像基督藉着父的荣耀从死人中复活一样。
ROM|6|5|我们若与他合一，经历与他一样的死，也将经历与他一样的复活。
ROM|6|6|我们知道，我们的旧人和他同钉十字架，使罪身灭绝，叫我们不再作罪的奴隶，
ROM|6|7|因为已死的人是脱离了罪。
ROM|6|8|我们若与基督同死，我们信也必与他同活，
ROM|6|9|因为知道基督既从死人中复活，就不再死，死也不再作他的主了。
ROM|6|10|他死了，是对罪死，只这一次；他活，是对上帝活着。
ROM|6|11|这样，你们也要看自己对罪是死的，在基督耶稣里对上帝却是活的。
ROM|6|12|所以，不要让罪在你们必死的身上掌权，使你们顺从身体的私欲。
ROM|6|13|也不要把你们的肢体献给罪作不义的工具，倒要像从死人中活着的人，把自己献给上帝，并把你们的肢体献给上帝作义的工具。
ROM|6|14|罪必不能作你们的主，因你们不在律法之下，而是在恩典之下。
ROM|6|15|那又怎么样呢？我们在恩典之下，不在律法之下，就可以犯罪吗？绝对不可！
ROM|6|16|难道你们不知道，你们献自己作奴仆，顺从谁就作谁的奴仆吗？或作罪的奴隶，以至于死；或作顺服的奴仆，以至于成义。
ROM|6|17|感谢上帝！因为你们从前虽然作罪的奴隶，现在却从心里顺服了所传给你们教导的典范。
ROM|6|18|你们既从罪里得了释放，就作了义的奴仆。
ROM|6|19|我因你们肉体的软弱，就以人的观点来说。你们从前怎样把肢体献给不洁不法作奴隶，以至于不法；现在也要照样将肢体献给义作奴仆，以至于成圣。
ROM|6|20|因为你们作罪的奴隶时，不被义所约束。
ROM|6|21|那么，你们现在所看为羞耻的事，当时有什么果子呢？那些事的结局就是死。
ROM|6|22|但如今，你们既从罪里得了释放，作了上帝的奴仆，就结出果子，以至于成圣，那结局就是永生。
ROM|6|23|因为罪的工价乃是死；惟有上帝的恩赐，在我们的主基督耶稣里，乃是永生。
ROM|7|1|弟兄们，我对你们这些明白律法的人说，你们岂不知道律法约束人是在他活着的时候吗？
ROM|7|2|就如女人有了丈夫，丈夫还活着，她就被律法约束；丈夫若死了，她就从丈夫的律法中解脱了。
ROM|7|3|所以丈夫还活着，她若跟了别的男人，就叫淫妇；丈夫若死了，她就脱离了律法，虽然跟了别的男人，也不是淫妇。
ROM|7|4|我的弟兄们，这样说来，你们藉着基督的身体对律法也是死了，使你们归于另一位，就是归于那从死人中复活的，为要使我们结果子给上帝。
ROM|7|5|因为我们属肉体的时候，那因律法而生犯罪的欲望在我们肢体中发动，以致结出死亡的果子。
ROM|7|6|但如今，我们既然在捆绑我们的律法上死了，就从律法中解脱，使我们服侍主，要按着圣灵 的新样，不按着仪文的旧样。
ROM|7|7|这样，我们要怎么说呢？律法是罪吗？绝对不是！但是，若不是藉着律法，我就不知何为罪；若不是律法说“不可贪心”，我就不知何为贪心。
ROM|7|8|然而，罪趁着机会，藉着诫命，使各样的贪心在我里头发动，因为没有律法，罪是死的。
ROM|7|9|以前没有律法的时候，我是活的；但是诫命来到，罪活起来，
ROM|7|10|我就死了。那本该叫人活的诫命反而叫我死。
ROM|7|11|因为罪趁着机会，藉着诫命诱惑我，并且藉着诫命杀了我。
ROM|7|12|这样看来，律法是圣的，诫命也是圣的、义的、善的。
ROM|7|13|那么，那善的是叫我死吗？绝对不是！叫我死的是罪。罪藉着那善的叫我死，为要显出这真是罪，以致罪藉着诫命更显出是恶极了。
ROM|7|14|我们原知道律法是属灵的，我却是属肉体的，是已经卖给罪了。
ROM|7|15|因为我所做的，我自己不明白。我所愿意的，我并不做；我所恨恶的，我反而去做。
ROM|7|16|如果我所做的是我所不愿意的，我得承认律法是善的。
ROM|7|17|事实上，这不是我做的，而是住在我里面的罪做的。
ROM|7|18|我也知道，住在我里面的，就是我肉体之中，没有善。因为立志为善由得我，只是行出来由不得我。
ROM|7|19|我所愿意的善，我不去做；我所不愿意的恶，我反而去做。
ROM|7|20|如果我去做我不愿意做的，就不是我做的，而是住在我里面的罪做的。
ROM|7|21|我觉得有个律，就是我愿意行善的时候，就有恶缠着我。
ROM|7|22|因为，按着我里面的人，我喜欢上帝的律，
ROM|7|23|但我看出肢体中另有个律和我内心的律交战，把我掳去，使我附从那肢体中罪的律。
ROM|7|24|我真苦啊！谁能救我脱离这必死的身体呢？
ROM|7|25|感谢上帝，靠着我们的主耶稣基督就能！这样看来，一方面，我内心顺服上帝的律，另一方面，肉体却顺服罪的律了。
ROM|8|1|如今，那些在基督耶稣里的人就不被定罪了。
ROM|8|2|因为赐生命的圣灵的律，在基督耶稣里从罪和死的律中把你释放出来。
ROM|8|3|律法既因肉体软弱而无能为力，上帝就差遣自己的儿子成为罪身的样子，为了对付罪 ，在肉体中定了罪，
ROM|8|4|为要使律法要求的义，实现在我们这不随从肉体、只随从圣灵去行的人身上。
ROM|8|5|因为，随从肉体的人体贴肉体的事；随从圣灵的人体贴圣灵的事。
ROM|8|6|体贴肉体就是死；体贴圣灵就是生命和平安 。
ROM|8|7|因为体贴肉体就是与上帝为敌，对上帝的律法不顺服，事实上也无法顺服。
ROM|8|8|属肉体的人无法使上帝喜悦。
ROM|8|9|如果上帝的灵住在你们里面，你们就不属肉体，而是属圣灵了。人若没有基督的灵，就不是属基督的。
ROM|8|10|基督若在你们里面，身体就因罪而死，灵却因义而活。
ROM|8|11|然而，使耶稣从死人中复活的上帝的灵若住在你们里面，那使基督从死人中复活的，也必藉着住在你们里面的圣灵使你们必死的身体又活过来。
ROM|8|12|弟兄们，这样看来，我们不是欠肉体的债去顺从肉体而活。
ROM|8|13|你们若顺从肉体活着，必定会死；若靠着圣灵把身体的恶行处死，就必存活。
ROM|8|14|因为凡被上帝的灵引导的都是上帝的儿子。
ROM|8|15|你们所领受的不是奴仆的灵，仍旧害怕；所领受的是儿子名分的灵，因此我们呼叫：“阿爸，父！”
ROM|8|16|圣灵自己与我们的灵一同见证我们是上帝的儿女。
ROM|8|17|若是儿女，就是后嗣，是上帝的后嗣，和基督同作后嗣。如果我们和他一同受苦，是要我们和他一同得荣耀。
ROM|8|18|我认为，现在的苦楚，若比起将来要显示给我们的荣耀，是不足介意的。
ROM|8|19|受造之物切望等候上帝的众子显出来。
ROM|8|20|因为受造之物屈服在虚空之下，不是自己愿意，而是因那使它屈服的叫他如此。但受造之物仍然指望从败坏的辖制下得释放，得享上帝儿女荣耀的自由。
ROM|8|21|
ROM|8|22|我们知道，一切受造之物一同呻吟，一同忍受阵痛，直到如今。
ROM|8|23|不但如此，就是我们这有圣灵作初熟果子的，也是自己内心呻吟，等候得着儿子的名分，就是我们的身体得救赎。
ROM|8|24|我们得救是在于盼望；可是看得见的盼望就不是盼望。谁还去盼望他所看得见的呢？
ROM|8|25|但我们若盼望那看不见的，我们就耐心等候。
ROM|8|26|同样，我们的软弱有圣灵帮助。我们本不知道当怎样祷告，但是圣灵亲自用无可言喻的叹息替我们祈求。
ROM|8|27|那鉴察人心的知道圣灵所体贴的，因为圣灵照着上帝的旨意替圣徒祈求。
ROM|8|28|我们知道，万事 都互相效力，叫爱上帝的人得益处，就是按他旨意被召的人。
ROM|8|29|因为他所预知的人，他也预定他们效法他儿子的榜样，使他儿子在许多弟兄中作长子 。
ROM|8|30|他所预定的人，他又召他们来；所召来的人，他又称他们为义；所称为义的人，他又叫他们得荣耀。
ROM|8|31|既是这样，我们对这些事还要怎么说呢？上帝若帮助我们，谁能抵挡我们呢？
ROM|8|32|上帝既不顾惜自己的儿子，为我们众人舍了他，岂不也把万物和他一同白白地赐给我们吗？
ROM|8|33|谁能控告上帝所拣选的人呢？有上帝称他们为义了。
ROM|8|34|谁能定他们的罪呢？有基督耶稣 已经死了，而且复活了，现今在上帝的右边，也替我们祈求。
ROM|8|35|谁能使我们与基督的爱隔绝呢？难道是患难吗？是困苦吗？是迫害吗？是饥饿吗？是赤身露体吗？是危险吗？是刀剑吗？
ROM|8|36|如经上所记： “我们为你的缘故终日被杀； 人看我们如将宰的羊。”
ROM|8|37|然而，靠着爱我们的主，在这一切的事上，我们已经得胜有余了。
ROM|8|38|因为我深信，无论是死，是活，是天使，是掌权的，是有权能的 ，是现在的事，是将来的事，
ROM|8|39|是高处的，是深处的，是别的受造之物，都不能使我们与上帝的爱隔绝，这爱是在我们的主基督耶稣里的。
ROM|9|1|我在基督里说真话，不说谎话；我的良心被圣灵感动为我作证。
ROM|9|2|我非常忧愁，心里时常伤痛。
ROM|9|3|为我弟兄，我骨肉之亲，就是自己被诅咒，与基督分离，我也愿意。
ROM|9|4|他们是 以色列 人，那儿子的名分、荣耀、诸约、律法的颁布、敬拜的礼仪、应许都是给他们的。
ROM|9|5|列祖是他们的，基督按肉体说也是从他们出来的。愿在万有之上的上帝被称颂，直到永远 。阿们！
ROM|9|6|这不是说上帝的话落了空。因为从 以色列 生的不都是 以色列 人，
ROM|9|7|也不因为是 亚伯拉罕 的后裔就都是他的儿女；惟独“从 以撒 生的才要称为你的后裔。”
ROM|9|8|这就是说，肉身所生的儿女不是上帝的儿女，惟独那应许的儿女才算是后裔。
ROM|9|9|因为所应许的话是这样：“到明年这时候我要来， 撒拉 必会生一个儿子。”
ROM|9|10|不但如此， 利百加 也是这样。她从一个人，就是从我们的祖宗 以撒 怀了孕。
ROM|9|11|双胞胎还没有生下来，善恶还没有行出来，为要贯彻上帝拣选人的旨意，
ROM|9|12|不是凭着人的行为，而是凭着那呼召人的，上帝就对 利百加 说：“将来，大的要服侍小的。”
ROM|9|13|正如经上所记：“ 雅各 是我所爱的； 以扫 是我所恶的。”
ROM|9|14|这样，我们要怎么说呢？难道上帝有什么不义吗？绝对没有！
ROM|9|15|因他对 摩西 说： “我要怜悯谁就怜悯谁， 要恩待谁就恩待谁。”
ROM|9|16|由此看来，这不靠人的意愿，也不靠人的努力，只靠上帝的怜悯。
ROM|9|17|因为经上有话对法老说：“我将你兴起来，特要在你身上彰显我的权能，为要使我的名传遍全地。”
ROM|9|18|由此看来，上帝要怜悯谁就怜悯谁，要使谁刚硬就使谁刚硬。
ROM|9|19|这样，你会对我说：“那么，他为什么还指责人呢？有谁能抗拒他的旨意呢？”
ROM|9|20|你这个人哪，你是谁，竟敢向上帝顶嘴呢？受造之物岂会对造他的说：“你为什么把我造成这样呢？”
ROM|9|21|难道陶匠没有权从一团泥里拿一块做成贵重的器皿，又拿一块做成卑贱的器皿吗？
ROM|9|22|倘若上帝要显明他的愤怒，彰显他的权能，难道不可多多忍耐宽容那应受愤怒、预备遭毁灭的器皿吗？
ROM|9|23|这是为了要把他丰盛的荣耀彰显在那蒙怜悯、早预备得荣耀的器皿上。
ROM|9|24|这器皿也就是我们这些蒙上帝所召的，不但是从 犹太 人中，也是从外邦人中召来的。
ROM|9|25|正如上帝在《何西阿书》上说： “那本来不是我子民的， 我要称为‘我的子民’； 本来不是蒙爱的， 我要称为‘蒙爱的’。
ROM|9|26|从前在什么地方对他们说： 你们不是我的子民， 将来就在那里称他们为‘永生上帝的儿子’。”
ROM|9|27|关于 以色列 人， 以赛亚 喊着：“虽然 以色列 人多如海沙，得救的将是剩下的余数，
ROM|9|28|因为主要在地上施行他的话，彻底而又迅速。”
ROM|9|29|又如 以赛亚 先前说过： “若不是万军之主给我们存留余种， 我们早已变成 所多玛 ，像 蛾摩拉 一样了。”
ROM|9|30|这样，我们要怎么说呢？那不追求义的外邦人却获得了义，就是因信而获得的义。
ROM|9|31|但 以色列 人追求律法的义，反而达不到律法的义。
ROM|9|32|这是什么缘故呢？是因为他们不凭着信心，而是凭着行为，他们正跌在那绊脚石上。
ROM|9|33|就如经上所记： “我在 锡安 放一块绊脚的石头，使人跌倒的磐石； 信靠他的人必不蒙羞。”
ROM|10|1|弟兄们，我心里所渴望的和向上帝所求的，是要 以色列 人得救。
ROM|10|2|我为他们作证，他们对上帝有热心，但不是按着真知识。
ROM|10|3|因为不明白上帝的义，想要立自己的义，他们就不服上帝的义了。
ROM|10|4|律法的总结就是基督，使所有信他的人都得着义。
ROM|10|5|论到出于律法的义， 摩西 写着：“行这些事的人，就必因此得生。”
ROM|10|6|但出于信的义却如此说：“你不要心里说：谁要升到天上去呢？（就是说，把基督领下来。）
ROM|10|7|或说：谁要下到阴间去呢？（就是说，把基督从死人中领上来。）”
ROM|10|8|他到底怎么说呢？ “这话语就离你近， 就在你口中，在你心里，” （就是说，我们传扬所信的话语。）
ROM|10|9|你若口里宣认耶稣为主，心里信上帝叫他从死人中复活，就必得救。
ROM|10|10|因为，人心里信就可以称义，口里宣认就可以得救。
ROM|10|11|经上说：“凡信靠他的人必不蒙羞。”
ROM|10|12|犹太 人和 希腊 人并没有分别，因为人人都有同一位主，他也厚待求告他的每一个人。
ROM|10|13|因为“凡求告主名的就必得救”。
ROM|10|14|然而，人未曾信他，怎能求告他呢？未曾听见他，怎能信他呢？没有传道的，怎能听见呢？
ROM|10|15|若没有奉差遣，怎能传道呢？如经上所记：“报福音、传喜信的人，他们的脚踪何等佳美！”
ROM|10|16|但不是每一个人都听从福音，因为 以赛亚 说：“主啊，我们所传的有谁信呢？”
ROM|10|17|可见，信道是从听道来的，听道是从基督的话来的。
ROM|10|18|但我要问，人没有听见吗？当然听见了。 “他们的声音传遍全地； 他们的言语传到地极。”
ROM|10|19|我再问， 以色列 人不知道吗？先有 摩西 说： “我要以不成国的激起你们嫉妒； 我要以愚顽的国惹起你们发怒。”
ROM|10|20|又有 以赛亚 放胆说： “没有寻找我的，我要让他们寻见； 没有求问我的，我要向他们显现。”
ROM|10|21|关于 以色列 人，他说：“我整天向那悖逆顶嘴的百姓招手。”
ROM|11|1|那么，我要问，上帝弃绝了他的百姓吗？绝对没有！因为我也是 以色列 人， 亚伯拉罕 的后裔，属 便雅悯 支派的。
ROM|11|2|上帝并没有弃绝他预先所知道的百姓。你们岂不知道经上论到 以利亚 是怎么说的呢？他在上帝面前怎样控告 以色列 人说：
ROM|11|3|“主啊，他们杀了你的先知，拆了你的祭坛，只剩下我一个人，他们还要我的命。”
ROM|11|4|但上帝的指示是怎么对他说的呢？他说：“我为自己留下七千人，是未曾向 巴力 屈膝的。”
ROM|11|5|现在这时刻也是这样，照着出于恩典的拣选，还有所留的余数。
ROM|11|6|既是靠恩典，就不凭行为，不然，恩典就不再是恩典了。
ROM|11|7|那又怎么说呢？ 以色列 人所寻求的，他们没有得着。但是蒙拣选的人得着了，其余的人却成了顽梗不化的。
ROM|11|8|如经上所记： “上帝给他们昏沉的灵， 眼睛看不见， 耳朵听不到， 直到今日。”
ROM|11|9|大卫 也说： “愿他们的宴席变为罗网，变为陷阱， 变为绊脚石，作他们的报应。
ROM|11|10|愿他们的眼睛昏花，看不见； 愿你时常弯下他们的腰。”
ROM|11|11|那么，我再问，他们失足是要他们跌倒吗？绝对不是！因他们的过犯，救恩反而临到外邦人，要激起他们嫉妒的心。
ROM|11|12|如果他们的过犯成为世界的富足，他们的缺乏成为外邦人的富足，更何况他们全数得救呢？
ROM|11|13|我对你们外邦人说，正因为我是外邦人的使徒，我敬重我的职分，
ROM|11|14|希望可以激起我骨肉之亲的嫉妒，好救他们一些人。
ROM|11|15|如果他们被丢弃，世界因而得以与上帝和好；他们被收纳，岂不就是从死人中复生吗？
ROM|11|16|所献的新面若圣洁，整个面团都圣洁了；树根若圣洁，树枝也圣洁了。
ROM|11|17|若有几根枝子被折下来，你这野橄榄枝接上去，同享橄榄根的肥汁，
ROM|11|18|你就不可向旧枝子夸口；若是夸口，该知道不是你托着根，而是根托着你。
ROM|11|19|你会说，那些枝子被折下来是为了使我接上去。
ROM|11|20|不错。他们因为不信，所以被折下来；你因为信，所以立得住。你不可自高，反要战战兢兢。
ROM|11|21|上帝既然不顾惜原来的枝子，岂会顾惜你？
ROM|11|22|可见，上帝又恩慈又严厉：对那跌倒的人是严厉的；对你是恩慈的，只要你长久在他的恩慈里，不然，你也要被砍下来。
ROM|11|23|而且，他们若不是长久不信，仍要被接上，因为上帝能够重新把他们接上去。
ROM|11|24|你是从那天生的野橄榄上砍下来的，尚且违反自然地接在好橄榄上，何况这些原来的枝子岂不更要接在原树上吗？
ROM|11|25|弟兄们，我不愿意你们不知道这奥秘，恐怕你们自以为聪明。这奥秘就是有一部分 以色列 人是硬心的，等到外邦人的数目添满了，
ROM|11|26|以色列 全家都要得救。如经上所记： “必有一位救主从 锡安 出来， 要消除 雅各 家一切不虔不敬。”
ROM|11|27|“这就是我与他们所立的约， 那时我要除去他们的罪。”
ROM|11|28|就福音来说，他们为你们的缘故是仇敌；就拣选来说，他们因列祖的缘故是蒙爱的。
ROM|11|29|因为上帝的恩赐和选召是不会撤回的。
ROM|11|30|你们从前不顺服上帝，如今因他们的不顺服，你们倒蒙了怜悯。
ROM|11|31|同样，他们现在也是不顺服，叫他们因着施给你们的怜悯，现在 也就蒙怜悯。
ROM|11|32|因为上帝把众人都圈在不顺服中，为的是要怜悯众人。
ROM|11|33|深哉，上帝的丰富、智慧和知识！ 他的判断何其难测！ 他的踪迹何其难寻！
ROM|11|34|谁知道主的心？ 谁作过他的谋士？
ROM|11|35|谁先给了他， 使他后来偿还呢？
ROM|11|36|因为万有都是本于他， 倚靠他，归于他。 愿荣耀归给他，直到永远。阿们！
ROM|12|1|所以，弟兄们，我以上帝的慈悲劝你们，将身体献上当作活祭，是圣洁的，是上帝所喜悦的，你们如此事奉乃是理所当然的 。
ROM|12|2|不要效法这个世界，只要心意更新而变化，叫你们察验何为上帝的善良、纯全、可喜悦的旨意。
ROM|12|3|我凭着所赐我的恩对你们每一位说：不要把自己看得太高，要照着上帝所分给各人的信心来衡量，看得合乎中道。
ROM|12|4|正如我们一个身子上有好些肢体，肢体也不都有一样的用处。
ROM|12|5|这样，我们许多人在基督里是一个身体，互相联络作肢体。
ROM|12|6|按着所得的恩典，我们各有不同的恩赐：或说预言，要按着信心的程度说预言；
ROM|12|7|或服事的，要专一服事；或教导的，要专一教导；
ROM|12|8|或劝勉的，要专一劝勉；施舍的，要诚实；治理的，要殷勤；怜悯人的，要乐意。
ROM|12|9|爱，不可虚假；恶，要厌恶；善，要亲近。
ROM|12|10|爱弟兄，要相亲相爱；恭敬人，要彼此推让；
ROM|12|11|殷勤，不可懒惰。要灵里火热；常常服侍主。
ROM|12|12|在盼望中要喜乐；在患难中要忍耐；祷告要恒切。
ROM|12|13|圣徒有缺乏，要供给；异乡客，要殷勤款待。
ROM|12|14|要祝福迫害你们 的，要祝福，不可诅咒。
ROM|12|15|要与喜乐的人同乐；要与哀哭的人同哭。
ROM|12|16|要彼此同心，不要心高气傲，倒要俯就卑微的人。不要自以为聪明。
ROM|12|17|不要以恶报恶，众人以为美的事要留心去做。
ROM|12|18|若是可行，总要尽力与众人和睦。
ROM|12|19|各位亲爱的，不要自己伸冤，宁可给主的愤怒留地步，因为经上记着：“主说：‘伸冤在我，我必报应。’”
ROM|12|20|不但如此，“你的仇敌若饿了，就给他吃；若渴了，就给他喝。因为你这样做，就是把炭火堆在他的头上。”
ROM|12|21|不要被恶所胜，反要以善胜恶。
ROM|13|1|在上有权柄的，人人要顺服，因为没有权柄不是来自上帝的。掌权的都是上帝所立的。
ROM|13|2|所以，抗拒掌权的就是抗拒上帝所立的；抗拒的人必自招审判。
ROM|13|3|作官的原不是要使行善的惧怕，而是要使作恶的惧怕。你愿意不惧怕掌权的吗？只要行善，你就可得他的称赞；
ROM|13|4|因为他是上帝的用人，是与你有益的。你若作恶，就该惧怕，因为他不是徒然佩剑；他是上帝的用人，为上帝的愤怒，报应作恶的。
ROM|13|5|所以，你们必须顺服，不但是因上帝的愤怒，也是因着良心。
ROM|13|6|你们纳粮也为这个缘故，因他们是上帝的仆役，专管这事。
ROM|13|7|凡人所当得的，就给他。当得粮的，给他纳粮；当得税的，给他上税；当惧怕的，惧怕他；当恭敬的，恭敬他。
ROM|13|8|你们除了彼此相爱，对任何人都不可亏欠什么，因为那爱人的就成全了律法。
ROM|13|9|那不可奸淫，不可杀人，不可偷盗，不可贪婪，或别的诫命，都包括在“爱邻 如己”这一句话之内了。
ROM|13|10|爱是不对邻人作恶，所以爱就成全了律法。
ROM|13|11|还有，你们要知道，现在正是该从睡梦中醒来的时候了；因为我们得救，现在比初信的时候更近了。
ROM|13|12|黑夜已深，白昼将近。所以我们该除去暗昧的行为，带上光明的兵器。
ROM|13|13|行事为人要端正，好像在白昼行走。不可荒宴醉酒；不可好色淫荡；不可纷争嫉妒。
ROM|13|14|总要披戴主耶稣基督，不要只顾满足肉体，去放纵私欲。
ROM|14|1|信心软弱的，你们要接纳，不同的意见，不要争论。
ROM|14|2|有人信什么都可吃；但那软弱的，只吃蔬菜。
ROM|14|3|吃的人不可轻看不吃的人；不吃的人也不可评断吃的人，因为上帝已经接纳他了。
ROM|14|4|你是谁，竟评断别人的仆人呢？他或站立或跌倒，自有他的主人在，而且他也必会站立，因为主能使他站稳。
ROM|14|5|有人看这日比那日强；有人看日日都是一样。只是各人要在自己的心意上坚定。
ROM|14|6|守日子的人是为主守的。吃的人是为主吃的，因他感谢上帝；不吃的人是为主不吃的，他也感谢上帝。
ROM|14|7|我们没有一个人为自己而活，也没有一个人为自己而死。
ROM|14|8|我们若活，是为主而活；我们若死，是为主而死。所以，我们或死或活总是主的人。
ROM|14|9|为此，基督死了，又活了，为要作死人和活人的主。
ROM|14|10|可是你，你为什么评断弟兄呢？你又为什么轻看弟兄呢？因我们都要站在上帝的审判台前。
ROM|14|11|经上写着： “主说，我指着我的永生起誓： 万膝必向我跪拜； 万口必称颂上帝。”
ROM|14|12|这样看来，我们各人一定要把自己的事在上帝面前 交代。
ROM|14|13|所以，我们不可再彼此评断，宁可决意不给弟兄放置障碍或绊脚石。
ROM|14|14|我凭着主耶稣确知深信，凡物本来没有不洁净的，除非人以为不洁净的，在他就不洁净了。
ROM|14|15|你若因食物使弟兄忧愁，就不是按着爱心行事。基督已经为他死，你不可因你的食物使他败坏。
ROM|14|16|所以，不可让你们的善被人毁谤。
ROM|14|17|因为上帝的国不在乎饮食，而在乎公义、和平及圣灵中的喜乐 。
ROM|14|18|凡这样服侍基督的，就为上帝所喜悦，又为人所赞许。
ROM|14|19|所以，我们务要追求 和平与彼此造就的事。
ROM|14|20|不可因食物毁坏上帝的工作。一切都是洁净的，但有人因食物使人跌倒，这在他就是恶了。
ROM|14|21|无论是吃肉是喝酒，是什么别的事，使弟兄跌倒，一概不做，才是善的。
ROM|14|22|你有信心，就要在上帝面前持守。人能在自己以为可行的事上不自责就有福了。
ROM|14|23|若有人疑惑而吃的，就被定罪，因为他吃不是出于信心。凡不出于信心的都是罪。
ROM|15|1|我们坚强的人应该分担不坚强的人的软弱，不求自己的喜悦。
ROM|15|2|我们各人务必要让邻人喜悦，使他得益处，得造就。
ROM|15|3|因为基督也不求自己的喜悦，如经上所记：“辱骂你的人的辱骂都落在我身上。”
ROM|15|4|从前所写的圣经都是为教导我们写的，要使我们藉着忍耐和因圣经所生的安慰，得着盼望。
ROM|15|5|但愿赐忍耐和安慰的上帝使你们彼此同心，效法基督耶稣，
ROM|15|6|为使你们同心同声荣耀我们主耶稣基督的父上帝！
ROM|15|7|所以，你们要彼此接纳，如同基督接纳你们一样，归荣耀给上帝。
ROM|15|8|我说，基督是为上帝真理作了受割礼的人的执事，要证实所应许列祖的话，
ROM|15|9|并使外邦人，因他的怜悯，荣耀上帝。如经上所记： “因此，我要在外邦中称颂你， 歌颂你的名。”
ROM|15|10|又说： “外邦人哪，你们要与主的子民一同欢乐。”
ROM|15|11|又说： “列邦啊，你们要赞美主！ 万民哪，你们都要颂赞他！”
ROM|15|12|又有 以赛亚 说： “将来有 耶西 的根， 就是那兴起来要治理列邦的； 外邦人要仰望他。”
ROM|15|13|愿赐盼望的上帝，因你们的信把各样的喜乐、平安 充满你们的心，使你们藉着圣灵的能力大有盼望！
ROM|15|14|我的弟兄们，我本人也深信你们自己充满良善，有各种丰富的知识，也能彼此劝戒。
ROM|15|15|但我更大胆写信给你们，是要在一些事上提醒你们，我因上帝所赐我的恩，
ROM|15|16|使我为外邦人作基督耶稣的仆役，作上帝福音的祭司，使所献上的外邦人因着圣灵成为圣洁，可蒙悦纳。
ROM|15|17|所以，有关上帝面前的事奉，我在基督耶稣里是有可夸的。
ROM|15|18|除了基督藉我做的那些事，我什么都不敢提，只提他藉我的言语作为，用神迹奇事的能力，并上帝的灵 的能力，使外邦人顺服；甚至我从 耶路撒冷 ，直转到 以利哩古 ，到处传了基督的福音。
ROM|15|19|
ROM|15|20|这样，我立了志向，不在基督的名已经传扬过的地方传福音，免得建造在别人的根基上；
ROM|15|21|却如经上所记： “未曾传给他们的，他们必看见； 未曾听见过的事，他们要明白。”
ROM|15|22|因此我多次被拦阻，不能到你们那里去。
ROM|15|23|但如今，在这一带再没有可传的地方，而且这许多年来，我迫切想去你们那里，
ROM|15|24|盼望到 西班牙 去的时候经过，得见你们，先与你们彼此交往，心里稍得满足，然后蒙你们为我送行。
ROM|15|25|但如今我要到 耶路撒冷 去，供应圣徒的需要。
ROM|15|26|因为 马其顿 和 亚该亚 人乐意凑出一些捐款给 耶路撒冷 圣徒中的穷人。
ROM|15|27|这固然是他们乐意的，其实也算是所欠的债；因为外邦人既然分享了他们灵性上的好处，就当把肉体上的需用供给他们。
ROM|15|28|等我办完了这事，把这笔捐款 交付给他们，我就要路过你们那里，到 西班牙 去。
ROM|15|29|我也知道去你们那里的时候，我将带着基督丰盛的恩典去。
ROM|15|30|弟兄们，我藉着我们的主耶稣基督，又藉着圣灵的爱，劝你们与我一同竭力为我祈求上帝，
ROM|15|31|使我脱离在 犹太 不顺从的人，也让我在 耶路撒冷 的事奉可蒙圣徒悦纳，
ROM|15|32|并使我照着上帝的旨意欢欢喜喜地到你们那里，与你们同得安息。
ROM|15|33|愿赐平安的上帝与你们众人同在。阿们！
ROM|16|1|我对你们推荐我们的姊妹 非比 ，她是 坚革哩 教会中的执事。
ROM|16|2|请你们在主里用合乎圣徒的方式来接待她。她在任何事上需要你们帮助，你们就帮助她；因她素来帮助许多人，也帮助了我。
ROM|16|3|请向 百基拉 和 亚居拉 问安。他们在基督耶稣里作我的同工，
ROM|16|4|也为我的性命把自己的生死置之度外；不但我感谢他们，就是外邦的众教会也感谢他们。
ROM|16|5|又向在他们家中的教会问安。向我所亲爱的 以拜尼土 问安，他是 亚细亚 归于基督的初结果子。
ROM|16|6|又向 马利亚 问安，她为你们非常辛劳。
ROM|16|7|又向与我一同坐监的亲戚 安多尼古 和 犹尼亚 问安，他们在使徒中是有名望的，也是比我先在基督里的。
ROM|16|8|又向我在主里面所亲爱的 暗伯利 问安。
ROM|16|9|又向我们在基督里的同工 耳巴奴 和我所亲爱的 士大古 问安。
ROM|16|10|又向在基督里经过考验的 亚比利 问安。向 亚利多布 家里的人问安。
ROM|16|11|又向我亲戚 希罗天 问安。向 拿其数 家在主里的人问安。
ROM|16|12|又向为主辛劳的 土非拿 和 土富撒 问安。向所亲爱、为主非常辛劳的 彼息 问安。
ROM|16|13|又向在主里蒙拣选的 鲁孚 和他母亲问安，他的母亲就是我的母亲。
ROM|16|14|又向 亚逊其土 、 弗勒干 、 黑米 、 八罗巴 、 黑马 ，和跟他们在一起的弟兄们问安。
ROM|16|15|又向 非罗罗古 和 犹利亚 ， 尼利亚 和他姊妹， 阿林巴 和跟他们在一起的众圣徒问安。
ROM|16|16|你们要以圣洁的吻彼此问安。基督的众教会都向你们问安！
ROM|16|17|弟兄们，那些离间你们、使你们跌倒、违背所学之道的人，我劝你们要留意躲避他们。
ROM|16|18|因为这样的人不服侍我们的主基督，只服侍自己的肚腹，用花言巧语诱惑老实人的心。
ROM|16|19|你们的顺服已经传于众人，所以我为你们欢喜；但我愿你们在善上聪明，在恶上愚拙。
ROM|16|20|那赐平安 的上帝快要把撒但践踏在你们脚下。愿我们主耶稣基督的恩与你们同在！
ROM|16|21|我的同工 提摩太 ，和我的亲戚 路求 、 耶孙 、 所西巴德 ，向你们问安。
ROM|16|22|我这代笔写信的 德提 ，在主里向你们问安。
ROM|16|23|那接待我，也接待全教会的 该犹 ，向你们问安。城里的财务官 以拉都 和弟兄 括土 向你们问安。
ROM|16|24|
ROM|16|25|惟有上帝能照我所传的福音和所讲的耶稣基督，并照历代以来隐藏的奥秘的启示，坚固你们。
ROM|16|26|这奥秘如今显示出来，而且按着永生上帝的命令，藉众先知的书指示万民，使他们因信而顺服。
ROM|16|27|愿荣耀，藉着耶稣基督，归给独一全智的上帝，直到永远。阿们！
