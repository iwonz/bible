PHIL|1|1|Paulus et Timotheus servi Christi Iesu omnibus sanctis in Christo Iesu, qui sunt Philippis, cum episcopis et diaconis:
PHIL|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
PHIL|1|3|Gratias ago Deo meo in omni memoria vestri,
PHIL|1|4|semper in omni oratione mea pro omnibus vobis cum gaudio deprecationem faciens
PHIL|1|5|super communione vestra in evangelio a prima die usque nunc;
PHIL|1|6|confidens hoc ipsum, quia, qui coepit in vobis opus bonum, perficiet usque in diem Christi Iesu;
PHIL|1|7|sicut est mihi iustum hoc sentire pro omnibus vobis, eo quod habeam in corde vos et in vinculis meis et in defensione et confirmatione evangelii socios gratiae meae omnes vos esse.
PHIL|1|8|Testis enim mihi Deus, quomodo cupiam omnes vos in visceribus Christi Iesu.
PHIL|1|9|Et hoc oro, ut caritas vestra magis ac magis abundet in scientia et omni sensu,
PHIL|1|10|ut probetis potiora, ut sitis sinceri et sine offensa in diem Christi,
PHIL|1|11|repleti fructu iustitiae, qui est per Iesum Christum, in gloriam et laudem Dei.
PHIL|1|12|Scire autem vos volo, fratres, quia, quae circa me sunt, magis ad profectum venerunt evangelii,
PHIL|1|13|ita ut vincula mea manifesta fierent in Christo in omni praetorio et in ceteris omnibus;
PHIL|1|14|et plures e fratribus in Domino confidentes vinculis meis, abundantius audere sine timore verbum loqui.
PHIL|1|15|Quidam quidem et propter invidiam et contentionem, quidam autem et propter bonam voluntatem Christum praedicant;
PHIL|1|16|hi quidem ex caritate scientes quoniam in defensionem evangelii positus sum,
PHIL|1|17|illi autem ex contentione Christum annuntiant, non sincere, existimantes pressuram se suscitare vinculis meis.
PHIL|1|18|Quid enim? Dum omni modo, sive sub obtentu sive in veritate, Christus annuntietur, et in hoc gaudeo; sed et gaudebo,
PHIL|1|19|scio enim quia hoc mihi proveniet in salutem per vestram orationem et subministrationem Spiritus Iesu Christi,
PHIL|1|20|secundum exspectationem et spem meam quia in nullo confundar, sed in omni fiducia, sicut semper et nunc, magnificabitur Christus in corpore meo, sive per vitam sive per mortem.
PHIL|1|21|Mihi enim vivere Christus est et mori lucrum.
PHIL|1|22|Quod si vivere in carne, hic mihi fructus operis est, et quid eligam ignoro.
PHIL|1|23|Coartor autem ex his duobus: desiderium habens dissolvi et cum Christo esse, multo magis melius;
PHIL|1|24|permanere autem in carne, magis necessarium est propter vos.
PHIL|1|25|Et hoc confidens, scio quia manebo et permanebo omnibus vobis ad profectum vestrum et gaudium fidei,
PHIL|1|26|ut gloriatio vestra abundet in Christo Iesu in me, per meum adventum iterum ad vos.
PHIL|1|27|Tantum digne evangelio Christi conversamini, ut sive cum venero et videro vos, sive absens audiam de vobis quia statis in uno Spiritu unanimes, concertantes fide evangelii;
PHIL|1|28|et in nullo perterriti ab adversariis, quod est illis indicium perditionis, vobis autem salutis, et hoc a Deo;
PHIL|1|29|quia vobis hoc donatum est pro Christo, non solum ut in eum credatis, sed ut etiam pro illo patiamini
PHIL|1|30|idem certamen habentes, quale vidistis in me et nunc auditis in me.
PHIL|2|1|Si qua ergo consolatio in Christo, si quod solacium cari tatis, si qua communio spiritus, si quae viscera et miserationes,
PHIL|2|2|implete gaudium meum, ut idem sapiatis, eandem caritatem habentes, unanimes, id ipsum sapientes;
PHIL|2|3|nihil per contentionem neque per inanem gloriam, sed in humilitate superiores sibi invicem arbitrantes;
PHIL|2|4|non, quae sua sunt, singuli considerantes, sed et ea, quae aliorum.
PHIL|2|5|Hoc sentite in vobis, quod et in Christo Iesu:
PHIL|2|6|qui cum in forma Dei esset,non rapinam arbitratus est esse se aequalem Deo,
PHIL|2|7|sed semetipsum exinanivit formam servi accipiens,in similitudinem hominum factus;et habitu inventus ut homo,
PHIL|2|8|humiliavit semetipsum factus oboediens usque ad mortem,mortem autem crucis.
PHIL|2|9|Propter quod et Deus illum exaltavitet donavit illi nomen,quod est super omne nomen,
PHIL|2|10|ut in nomine Iesu omne genu flectaturcaelestium et terrestrium et infernorum,
PHIL|2|11|et omnis lingua confiteatur Dominus Iesus Christus! ",in gloriam Dei Patris.
PHIL|2|12|Itaque, carissimi mei, sicut semper oboedistis, non ut in praesentia mei tantum sed multo magis nunc in absentia mea, cum metu et tremore vestram salutem operamini;
PHIL|2|13|Deus est enim, qui operatur in vobis et velle et perficere pro suo beneplacito.
PHIL|2|14|Omnia facite sine murmurationibus et haesitationibus,
PHIL|2|15|ut efficiamini sine querela et simplices, filii Dei sine reprehensione in medio generationis pravae et perversae, inter quos lucetis sicut luminaria in mundo,
PHIL|2|16|verbum vitae firmiter tenentes ad gloriam meam in die Christi, quia non in vacuum cucurri neque in vacuum laboravi.
PHIL|2|17|Sed et si delibor supra sacrificium et obsequium fidei vestrae, gaudeo et congaudeo omnibus vobis;
PHIL|2|18|idipsum autem et vos gaudete et congaudete mihi.
PHIL|2|19|Spero autem in Domino Iesu Timotheum cito me mittere ad vos, ut et ego bono animo sim, cognitis, quae circa vos sunt.
PHIL|2|20|Neminem enim habeo tam unanimem, qui sincere pro vobis sollicitus sit;
PHIL|2|21|omnes enim sua quaerunt, non quae sunt Iesu Christi.
PHIL|2|22|Probationem autem eius cognoscitis, quoniam sicut patri filius mecum servivit in evangelium.
PHIL|2|23|Hunc igitur spero me mittere, mox ut videro, quae circa me sunt;
PHIL|2|24|confido autem in Domino, quoniam et ipse cito veniam.
PHIL|2|25|Necessarium autem existimavi Epaphroditum fratrem et cooperatorem et commilitonem meum, vestrum autem apostolum et ministrum necessitatis meae, mittere ad vos,
PHIL|2|26|quoniam omnes vos desiderabat et maestus erat, propterea quod audieratis illum infirmatum.
PHIL|2|27|Nam et infirmatus est usque ad mortem, sed Deus misertus est eius; non solum autem eius, verum et mei, ne tristitiam super tristitiam haberem.
PHIL|2|28|Festinantius ergo misi illum, ut, viso eo, iterum gaudeatis, et ego sine tristitia sim.
PHIL|2|29|Excipite itaque illum in Domino cum omni gaudio et eiusmodi cum honore habetote,
PHIL|2|30|quoniam propter opus Christi usque ad mortem accessit in interitum tradens animam suam, ut suppleret id, quod vobis deerat ministerii erga me.
PHIL|3|1|De cetero, fratres mei, gaudete in Domino. Eadem vobis scribe re mihi quidem non pigrum, vobis autem securum.
PHIL|3|2|Videte canes, videte malos operarios, videte concisionem!
PHIL|3|3|Nos enim sumus circumcisio, qui Spiritu Dei servimus et gloriamur in Christo Iesu et non in carne fiduciam habentes,
PHIL|3|4|quamquam ego habeam confidentiam et in carne. Si quis alius videtur confidere in carne, ego magis:
PHIL|3|5|circumcisus octava die, ex genere Israel, de tribu Beniamin, Hebraeus ex Hebraeis, secundum legem pharisaeus,
PHIL|3|6|secundum aemulationem persequens ecclesiam, secundum iustitiam, quae in lege est, conversatus sine querela.
PHIL|3|7|Sed, quae mihi erant lucra, haec arbitratus sum propter Christum detrimentum.
PHIL|3|8|Verumtamen existimo omnia detrimentum esse propter eminentiam scientiae Christi Iesu Domini mei, propter quem omnia detrimentum feci et arbitror ut stercora, ut Christum lucrifaciam
PHIL|3|9|et inveniar in illo non habens meam iustitiam, quae ex lege est, sed illam, quae per fidem est Christi, quae ex Deo est iustitia in fide;
PHIL|3|10|ad cognoscendum illum et virtutem resurrectionis eius et communionem passionum illius, conformans me morti eius,
PHIL|3|11|si quo modo occurram ad resurrectionem, quae est ex mortuis.
PHIL|3|12|Non quod iam acceperim aut iam perfectus sim; persequor autem si umquam comprehendam, sicut et comprehensus sum a Christo Iesu.
PHIL|3|13|Fratres, ego me non arbitror comprehendisse; unum autem: quae quidem retro sunt, obliviscens, ad ea vero, quae ante sunt, extendens me
PHIL|3|14|ad destinatum persequor, ad bravium supernae vocationis Dei in Christo Iesu.
PHIL|3|15|Quicumque ergo perfecti, hoc sentiamus; et si quid aliter sapitis, et hoc vobis Deus revelabit;
PHIL|3|16|verumtamen, ad quod pervenimus, in eodem ambulemus.
PHIL|3|17|Coimitatores mei estote, fratres, et observate eos, qui ita ambulant, sicut habetis formam nos.
PHIL|3|18|Multi enim ambulant, quos saepe dicebam vobis, nunc autem et flens dico, inimicos crucis Christi,
PHIL|3|19|quorum finis interitus, quorum deus venter et gloria in confusione ipsorum, qui terrena sapiunt.
PHIL|3|20|Noster enim municipatus in caelis est, unde etiam salvatorem exspectamus Dominum Iesum Christum,
PHIL|3|21|qui transfigurabit corpus humilitatis nostrae, ut illud conforme faciat corpori gloriae suae secundum operationem, qua possit etiam subicere sibi omnia.
PHIL|4|1|Itaque, fratres mei carissimi et desideratissimi, gaudium et co rona mea, sic state in Domino, carissimi!
PHIL|4|2|Evodiam rogo et Syntychen deprecor idipsum sapere in Domino.
PHIL|4|3|Etiam rogo et te, germane compar, adiuva illas, quae mecum concertaverunt in evangelio cum Clemente et ceteris adiutoribus meis, quorum nomina sunt in libro vitae.
PHIL|4|4|Gaudete in Domino semper. Iterum dico: Gaudete!
PHIL|4|5|Modestia vestra nota sit omnibus hominibus. Dominus prope.
PHIL|4|6|Nihil solliciti sitis, sed in omnibus oratione et obsecratione cum gratiarum actione petitiones vestrae innotescant apud Deum.
PHIL|4|7|Et pax Dei, quae exsuperat omnem sensum, custodiet corda vestra et intellegentias vestras in Christo Iesu.
PHIL|4|8|De cetero, fratres, quaecumque sunt vera, quaecumque pudica, quaecumque iusta, quaecumque casta, quaecumque amabilia, quaecumque bonae famae, si qua virtus et si qua laus, haec cogitate;
PHIL|4|9|quae et didicistis et accepistis et audistis et vidistis in me, haec agite; et Deus pacis erit vobiscum.
PHIL|4|10|Gavisus sum autem in Domino vehementer, quoniam tandem aliquando refloruistis pro me sentire, sicut et sentiebatis, opportunitate autem carebatis.
PHIL|4|11|Non quasi propter penuriam dico, ego enim didici, in quibus sum, sufficiens esse.
PHIL|4|12|Scio et humiliari, scio et abundare; ubique et in omnibus institutus sum et satiari et esurire et abundare et penuriam pati.
PHIL|4|13|Omnia possum in eo, qui me confortat.
PHIL|4|14|Verumtamen bene fecistis communicantes tribulationi meae.
PHIL|4|15|Scitis autem et vos, Philippenses, quod in principio evangelii, quando profectus sum a Macedonia, nulla mihi ecclesia communicavit in ratione dati et accepti, nisi vos soli;
PHIL|4|16|quia et Thessalonicam et semel et bis in usum mihi misistis.
PHIL|4|17|Non quia quaero datum, sed requiro fructum, qui abundet in rationem vestram.
PHIL|4|18|Accepi autem omnia et abundo; repletus sum acceptis ab Epaphrodito, quae misistis odorem suavitatis, hostiam acceptam, placentem Deo.
PHIL|4|19|Deus autem meus implebit omne desiderium vestrum secundum divitias suas in gloria in Christo Iesu.
PHIL|4|20|Deo autem et Patri nostro gloria in saecula saeculorum. Amen.
PHIL|4|21|Salutate omnem sanctum in Christo Iesu. Salutant vos, qui mecum sunt, fratres.
PHIL|4|22|Salutant vos omnes sancti, maxime autem, qui de Caesaris domo sunt.
PHIL|4|23|Gratia Domini Iesu Christi cum spiritu vestro. Amen.
