2JOHN|1|1|Presbyter electae dominae et filiis eius, quos ego diligo in veritate, et non ego solus, sed et omnes, qui noverunt veritatem,
2JOHN|1|2|propter veritatem, quae permanet in nobis et nobiscum erit in sempiternum.
2JOHN|1|3|Erit nobiscum gratia, misericordia, pax a Deo Patre et a Iesu Christo, Filio Patris, in veritate et caritate.
2JOHN|1|4|Gavisus sum valde, quoniam inveni de filiis tuis ambulantes in veritate, sicut mandatum accepimus a Patre.
2JOHN|1|5|Et nunc rogo te, domina, non tamquam mandatum novum scribens tibi, sed quod habuimus ab initio, ut diligamus alterutrum.
2JOHN|1|6|Et haec est caritas, ut ambulemus secundum mandata eius; hoc mandatum est, quemadmodum audistis ab initio, ut in eo ambuletis.
2JOHN|1|7|Quoniam multi seductores prodierunt in mundum, qui non confitentur Iesum Christum venientem in carne; hic est seductor et antichristus.
2JOHN|1|8|Videte vosmetipsos, ne perdatis, quae operati estis, sed ut mercedem plenam accipiatis.
2JOHN|1|9|Omnis, qui ultra procedit et non manet in doctrina Christi, Deum non habet; qui permanet in doctri na, hic et Patrem et Filium habet.
2JOHN|1|10|Si quis venit ad vos et hanc doctrinam non affert, nolite accipere eum in domum nec " Ave " ei dixeritis;
2JOHN|1|11|qui enim dicit illi: " Ave ", communicat operibus illius malignis.
2JOHN|1|12|Plura habens vobis scribere, nolui per chartam et atramentum; spero enim me futurum apud vos, et os ad os loqui, ut gaudium nostrum plenum sit.
2JOHN|1|13|Salutant te filii sororis tuae electae.
