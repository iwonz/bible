EZEK|1|1|在三十年四月初五，我在 迦巴鲁河 边被掳的人当中，那时天开了，我看见上帝的异象。
EZEK|1|2|正是 约雅斤 王被掳的第五年四月初五，
EZEK|1|3|在 迦勒底 人之地的 迦巴鲁河 边，耶和华的话特地临到 布西 的儿子 以西结 祭司，耶和华的手按在他身上。
EZEK|1|4|我观看，看哪，狂风从北方刮来，有一朵大云闪烁着火，周围有光辉，其中的火好像闪耀的金属；
EZEK|1|5|又从其中显出四个活物的形像。他们的形状是这样：有人的形像，
EZEK|1|6|各有四张脸，四个翅膀。
EZEK|1|7|他们的腿是直的，脚掌好像牛犊的蹄，灿烂如磨亮的铜。
EZEK|1|8|在四面的翅膀以下有人的手。这四个活物的脸和翅膀是这样：
EZEK|1|9|翅膀彼此相接，行走时并不转弯，各自往前直行。
EZEK|1|10|至于脸的形像：四个活物各有人的脸，右面有狮子的脸，左面有牛的脸，也有鹰的脸；
EZEK|1|11|这就是他们的脸 。他们的翅膀向上张开，各有两个翅膀彼此相接，用另外两个翅膀遮体。
EZEK|1|12|他们各自往前直行。灵往哪里去，他们就往哪里去，行走时并不转弯。
EZEK|1|13|至于四活物的形像，就如烧着火炭的形状，又如火把的形状。有火在四活物中间来回移动，这火有光辉，从火中发出闪电。
EZEK|1|14|这些活物往来奔走，好像电光一闪。
EZEK|1|15|我观看活物，看哪，有四张脸的活物旁边各有一个轮子在地上。
EZEK|1|16|轮子的形状结构 好像耀眼的水苍玉。四轮都是一个样式，形状 结构好像轮中套轮。
EZEK|1|17|轮子行走的时候，向四方直行，行走时并不转弯。
EZEK|1|18|至于轮圈，高而可畏；四个轮圈周围布满眼睛。
EZEK|1|19|活物行走，轮子也在旁边行走；活物离地上升，轮子也上升。
EZEK|1|20|灵往哪里去，活物就往哪里去；轮子在活物旁边上升，因为活物的灵在轮中。
EZEK|1|21|活物行走，轮子也行走；活物站住，轮子也站住；活物离地上升，轮子也在旁边上升，因为活物的灵在轮中。
EZEK|1|22|活物的头上面有穹苍的形像，像耀眼惊人的水晶，铺张在活物的头顶上。
EZEK|1|23|穹苍之下，活物的翅膀伸直，彼此相对，每个活物用两个翅膀遮住自己；每个活物用两个翅膀遮住自己 ，就是自己的身体。
EZEK|1|24|活物行走的时候，我听见翅膀的响声，像大水的声音，像全能者的声音，又像军队闹哄的声音。活物站住的时候，翅膀垂下。
EZEK|1|25|在他们头上的穹苍之上有声音。他们站住的时候，翅膀垂下。
EZEK|1|26|在他们头上的穹苍之上有宝座的形像，仿佛蓝宝石的样子；宝座的形像上方有仿佛人的样子的形像。
EZEK|1|27|我见他的腰以上有仿佛闪耀的金属，周围有仿佛火的形状，又见他的腰以下有仿佛火的形状，周围也有光辉。
EZEK|1|28|下雨的日子，云中彩虹的形状怎样，周围光辉的形状也是怎样。 这就是耶和华荣耀形像的样式，我一看见就脸伏于地。我又听见一位说话者的声音。
EZEK|2|1|他对我说：“人子啊，你站起来，我要和你说话。”
EZEK|2|2|他对我说话的时候，灵进入我里面，使我站起来，我就听见他对我说话。
EZEK|2|3|他对我说：“人子啊，我差你往悖逆我的国家， 以色列 人那里去，他们是悖逆我的。他们和他们的祖先违背我，直到今日。
EZEK|2|4|这些人厚着脸皮，心里刚硬。我差你到他们那里去，你要对他们说：‘主耶和华如此说。’
EZEK|2|5|他们是悖逆之家，他们或听，或不听，必知道在他们中间有了先知。
EZEK|2|6|你，人子啊，虽有荆棘和蒺藜在你那里，你又住在蝎子中间，总不要怕他们，也不要怕他们的话；他们虽是悖逆之家，但你不要怕他们的话，也不要因他们的脸色惊惶。
EZEK|2|7|他们或听，或不听，你只管将我的话告诉他们；他们是极其悖逆的。
EZEK|2|8|“但是你，人子啊，要听我对你说的话，不要像那悖逆之家一样悖逆，要开口吃我所赐给你的。”
EZEK|2|9|我观看，看哪，有一只手向我伸来；看哪，手中有一书卷。
EZEK|2|10|他在我面前展开书卷，它内外都写着字，上面所写的有哀号、叹息、悲痛的话。
EZEK|3|1|他对我说：“人子啊，要吃你所得到的，吃下这书卷；然后要去，对 以色列 家宣讲。”
EZEK|3|2|于是我张开了口，他就使我吃这书卷。
EZEK|3|3|他对我说：“人子啊，要吃我所赐给你的这书卷，塞满你的肚腹。”我就吃了，口中觉得其甜如蜜。
EZEK|3|4|他对我说：“人子啊，你要到 以色列 家那里去，对他们传讲我的话。
EZEK|3|5|你奉差遣不是往那说话艰涩、言语难懂的民那里，而是往 以色列 家去；
EZEK|3|6|你不是往那说话艰涩、言语难懂的许多民族那里去，他们的话你不懂。然而，我若差你往他们那里去，他们会听从你。
EZEK|3|7|以色列 家却不肯听从你，因为他们不肯听从我；原来 以色列 全家是额头坚硬、心里刚愎的人。
EZEK|3|8|看哪，我使你的脸坚硬，对抗他们的脸；使你的额头坚硬，对抗他们的额头。
EZEK|3|9|我使你的额头像金刚石，比火石更坚硬。他们虽是悖逆之家，但你不要怕他们，也不要因他们的脸色而惊惶。”
EZEK|3|10|他又对我说：“人子啊，我对你说的一切话，你心里要领会，耳朵要听。
EZEK|3|11|要到被掳的人，到你本国百姓那里去，他们或听，或不听，你要对他们宣讲，告诉他们这是主耶和华说的。”
EZEK|3|12|那时，灵将我举起，我就听见在我身后有极大震动的声音：“耶和华的荣耀，从他所在之处，是应当称颂的！”
EZEK|3|13|有活物的翅膀相碰的声音，也有活物旁边轮子的声音，是极大震动的声音。
EZEK|3|14|于是灵将我举起，带着我走。我就去了，十分苦恼，我的灵火热；耶和华的手重重地按在我身上。
EZEK|3|15|我就来到 提勒．亚毕 那些住在 迦巴鲁河 边被掳的人那里，到他们住的地方 ，在他们中间惊愕地坐了七日。
EZEK|3|16|过了七日，耶和华的话临到我，说：
EZEK|3|17|“人子啊，我立你作 以色列 家的守望者，所以你要听我口中的话，替我警戒他们。
EZEK|3|18|我何时指着恶人说：‘他必要死’；你若不警戒他，也不劝告他，使他离开恶行，拯救他的性命，这恶人必死在罪孽之中；我却要从你手里讨他的血债。
EZEK|3|19|倘若你警戒恶人，他仍不转离罪恶，也不离开恶行，他必死在罪孽之中，你却救了自己的命。
EZEK|3|20|但是义人若转离他的义而作恶，我要把绊脚石放在他面前，他必死亡；因你没有警戒他，他必死在罪中，他素来所行的义不被记念；我却要从你手里讨他的血债。
EZEK|3|21|倘若你警戒义人，使他不犯罪，他就不犯罪；他因领受警戒就必存活，你也救了自己的命。”
EZEK|3|22|在那里耶和华的手按在我身上。他对我说：“起来，到平原去，我要在那里和你说话。”
EZEK|3|23|于是我起来，到平原去，看哪，耶和华的荣耀停在那里，正如我在 迦巴鲁河 边所见到的一样，我就脸伏于地。
EZEK|3|24|灵进入我里面，使我站起来。耶和华对我说：“你进屋里去，把门关上。
EZEK|3|25|你，人子，看哪，人要用绳索捆绑你，使你不能出去到他们中间。
EZEK|3|26|我必使你的舌头贴住上膛，以致你哑口，不能作责备他们的人；他们原是悖逆之家。
EZEK|3|27|但我对你说话的时候，必使你开口，你就要对他们说：‘主耶和华如此说。’听的，让他听；不听的，任他不听，因为他们是悖逆之家。”
EZEK|4|1|“你，人子啊，拿一块砖，摆在你面前，将一座城 耶路撒冷 画在上面。
EZEK|4|2|你要围攻这城，筑堡垒，建土堆，安营攻击，周围设撞城槌攻城，
EZEK|4|3|又要拿一个铁盘放在你和城的中间，作为铁墙。你要把你的脸对着这城，使城被困。你要围攻这城，这要成为 以色列 家的预兆。
EZEK|4|4|“你要向左侧卧，承担 以色列 家的罪孽；按你向左侧卧的日数，担当他们的罪孽。
EZEK|4|5|我已将他们作恶的年数定了日期，就是三百九十天，你要如此担当 以色列 家的罪孽。
EZEK|4|6|这些日子结束之后，你还要向右侧卧，担当 犹大 家的罪孽。我为你定了四十天，一天顶一年。
EZEK|4|7|你要把你的脸对着被困的 耶路撒冷 ，露出膀臂，说预言攻击这城。
EZEK|4|8|看哪，我用绳索捆绑你，使你不能从这边翻到那边，直等到你围困的日子结束。
EZEK|4|9|“你要取小麦、大麦、豆子、红豆、小米、粗麦，装在一个器皿里，为自己做饼；在你侧卧的三百九十天吃这饼。
EZEK|4|10|你所吃食物的量是每天二十舍客勒，要按时吃。
EZEK|4|11|你喝水的量是每天六分之一欣，要按时喝。
EZEK|4|12|你要吃这饼像大麦饼一样，在众人眼前用人的粪烤它。”
EZEK|4|13|耶和华说：“ 以色列 人在我赶他们到的列国中，也必这样吃不洁净的食物。”
EZEK|4|14|我说：“唉！主耶和华，看哪，我从来未曾被玷污，从幼年到如今没有吃过自然死的，或被野兽撕裂的，那不洁净的肉也未曾入我的口。”
EZEK|4|15|于是他对我说：“看，我给你牛粪代替人粪，你要在上面烤你的饼。”
EZEK|4|16|他又对我说：“人子，看哪，我必断绝 耶路撒冷 粮食的供应 。他们要带着忧虑限量吃饼；带着惊惶限量喝水。
EZEK|4|17|他们因缺粮缺水，彼此惊惶，在自己的罪孽中消灭。”
EZEK|5|1|“你，人子啊，拿一把快刀当作剃刀，用这刀剃你的头发和胡须，然后用天平将须发分成几份。
EZEK|5|2|围困的日子满了，你要把三分之一放在城中用火焚烧；三分之一放在城的四围用刀砍碎；三分之一任风吹散，我要拔刀追赶它们。
EZEK|5|3|你要从其中取几根须发，用衣服的边包起来，
EZEK|5|4|再从其中取一些扔在火里，在火中焚烧；必有火从其中出来烧尽 以色列 全家。
EZEK|5|5|主耶和华如此说：这就是 耶路撒冷 。我曾将它安置在列国中，列邦都在它的四围。
EZEK|5|6|耶路撒冷 行恶，违背我的典章，过于列国；干犯我的律例，过于四围的列邦。它弃绝我的典章，也没有遵行我的律例。
EZEK|5|7|所以主耶和华如此说：因为你们混乱，过于四围的列国，不遵行我的律例，不顺从我的典章，甚至也不顺从四围列国的规条 ，
EZEK|5|8|所以主耶和华如此说：看哪，我，我必与你为敌，必在列国眼前，在你中间施行审判；
EZEK|5|9|并且因你一切可憎的事，我要在你中间行未曾行过，将来也不会行的事。
EZEK|5|10|在你中间，父亲要吃儿子，儿子要吃父亲。我必向你施行审判，将你剩下的人分散四方 。
EZEK|5|11|主耶和华说：我指着我的永生起誓，因你用一切可憎之物、可厌的事玷污我的圣所，所以，我要把你剃光 ，我的眼必不顾惜你，也不可怜你。
EZEK|5|12|你的百姓三分之一必遭瘟疫而死，因饥荒在你们中间而消灭；三分之一必在你四围倒在刀下；我必将三分之一分散四方，要拔刀追赶他们。
EZEK|5|13|“我要这样发尽我的怒气；我向他们发的愤怒停止以后，自己就得到平息。当我向他们发尽我的愤怒时，他们就知道我─耶和华所说的是出于妒忌。
EZEK|5|14|在四围的列国中，我要使你成为荒凉，在所有过路人的眼前看为羞辱。
EZEK|5|15|这样，我必以怒气、愤怒和烈怒的责备，向你施行审判。那时，它 就在四围的列国中成为羞辱、讥刺、警戒、惊骇；这是我─耶和华说的。
EZEK|5|16|我向灭亡的人射出饥荒的恶箭，将它们射出，毁灭你们；那时，我要加重你们的饥荒，断绝你们粮食的供应。
EZEK|5|17|我要令饥荒和恶兽临到你，使你丧失儿女。瘟疫和流血的事必在你那里盛行，我也要使刀剑临到你。这是我─耶和华说的。”
EZEK|6|1|耶和华的话临到我，说：
EZEK|6|2|“人子啊，你要面向 以色列 的众山说预言。
EZEK|6|3|你要说： 以色列 的众山哪，要听主耶和华的话。主耶和华对大山、小冈、水沟、山谷如此说：看哪，我要使刀剑临到你们，也必毁坏你们的丘坛。
EZEK|6|4|你们的祭坛要荒废，香坛必打碎。我要使你们当中被杀的人仆倒在你们的偶像面前，
EZEK|6|5|将 以色列 人的尸首放在他们的偶像面前，把你们的骸骨抛散在祭坛的四周围。
EZEK|6|6|无论你们住在何处，城镇要变为废墟，丘坛也必毁坏，以至于你们的祭坛荒废，被定罪 ，偶像打碎消除，香坛砍倒；你们所做的被涂去。
EZEK|6|7|被杀的人必仆倒在你们中间，你们就知道我是耶和华。
EZEK|6|8|“我必留下一些人，你们中有人得以在列国中脱离刀剑，分散在列邦。
EZEK|6|9|那些逃脱的人，必在被掳所到的各国中记得我，我心里何等伤痛，因他们起淫心，离弃我，淫荡的眼追随偶像。他们因所做一切可憎的恶事，必厌恶自己。
EZEK|6|10|他们必知道我是耶和华；我说过要使这灾祸临到他们身上，并非空话。
EZEK|6|11|“主耶和华如此说：你当击掌顿足，说：哀哉！ 以色列 家做了这一切可憎的恶事，必仆倒在刀剑、饥荒、瘟疫之下。
EZEK|6|12|在远方的，必遭瘟疫而死；在近处的，必倒在刀剑之下；那存留被围困的，必因饥荒而死；我要在他们身上发尽我的愤怒。
EZEK|6|13|被杀的要仆倒在祭坛四围的偶像中，在各高冈、各山顶、各青翠的树下，和各茂密的橡树下，就是他们献馨香的祭给一切偶像的地方。那时，他们就知道我是耶和华。
EZEK|6|14|我必伸手攻击他们，使他们的地荒废，从 第伯拉他 的旷野起 ，一切的住处都荒凉。他们就知道我是耶和华。”
EZEK|7|1|耶和华的话又临到我，说：
EZEK|7|2|“你，人子啊，主耶和华对 以色列 地如此说：结局，结局临到了地的四境！
EZEK|7|3|现在你的结局已经来临；我要使我的怒气临到你，也要按你的行为审判你，照你所做一切可憎的事惩罚你。
EZEK|7|4|我的眼必不顾惜你，也不可怜你，却要按你所做的报应你，照你们中间可憎的事惩罚你；你就知道我是耶和华。
EZEK|7|5|“主耶和华如此说：灾难，惟一的灾难 ，看哪，临近了！
EZEK|7|6|结局到了，结局到了，它要醒起来攻击你。看哪，它已来到！
EZEK|7|7|境内的居民哪，厄运临到你；时候到了，日子近了，有闹哄，但不是山上欢呼的声音。
EZEK|7|8|我快要将我的愤怒倾倒在你身上，向你发尽我的怒气，按你的行为审判你，照你所做一切可憎的事惩罚你。
EZEK|7|9|我的眼必不顾惜你，也不可怜你，必按你所做的报应你，照你中间可憎的事惩罚你；你就知道击打你的是我─耶和华。
EZEK|7|10|“看哪，那日子！看哪，已来到！厄运已经发生！杖已开花，骄傲已发芽。
EZEK|7|11|残暴兴起，成了罚恶的杖。他们将一无所有，他们的富足 、他们的财宝 都不复存在；他们中间也不再有尊荣。
EZEK|7|12|时候到了，日子近了，买主不可欢喜，卖主也不用愁烦，因为烈怒已经临到他们众人身上。
EZEK|7|13|卖主即使存活，也不能讨回所卖的，因为这异象关乎他们众人；谁都不能讨回，也没有人能在罪孽中使自己的生命刚强。”
EZEK|7|14|“他们吹了角，预备齐全，却无一人出战，因为我的烈怒临到他们众人身上。
EZEK|7|15|外有刀剑，内有瘟疫、饥荒。在田野的，必因刀剑而死；在城中的，必遭饥荒、瘟疫吞灭。
EZEK|7|16|其中幸存的要逃脱，各人因自己的罪孽在山上发出悲声，如谷中的鸽子哀鸣；
EZEK|7|17|双手发软，膝盖软弱如水，
EZEK|7|18|腰束麻布，战栗笼罩他们；各人脸上羞愧，头上光秃。
EZEK|7|19|他们要把银子抛弃在街上，看金子如污秽之物。正当耶和华发怒的日子，金银不能拯救他们，不能满足食欲，也不能使肚腹饱满，反倒成了自己罪孽的绊脚石。
EZEK|7|20|他们用所夸耀华美的妆饰制造可憎可厌的偶像，所以我使他们看它如污秽之物。
EZEK|7|21|我必将它交给外邦人为掠物，交给地上的恶人为掳物；他们要亵渎它。
EZEK|7|22|他们亵渎我宝贵之所 ，强盗也进去亵渎它。我必转脸不顾 以色列 人 。
EZEK|7|23|“要制造锁链；因为遍地都有流血的罪，满城都是残暴的事。
EZEK|7|24|所以，我要使列国中最凶恶的人前来占据他们的房屋；我要止息残暴人的骄傲，他们的圣所也要被亵渎。
EZEK|7|25|毁灭来到；他们求平安，却没有平安。
EZEK|7|26|灾害加上灾害，风声接连风声；他们要向先知寻求异象，但祭司的教诲、长老的谋略都必断绝。
EZEK|7|27|君王要悲哀，官长要披绝望为衣，这地百姓的手都发颤。我必照他们所做的待他们，按他们所应得的审判他们，他们就知道我是耶和华。”
EZEK|8|1|第六年六月初五，我坐在家中； 犹大 的众长老坐在我面前。在那里主耶和华的手降在我身上。
EZEK|8|2|我观看，看哪，有形像仿佛火 的形状，从他腰部以下形状是火，从他腰部以上有光辉的形状，好像闪耀的金属。
EZEK|8|3|他伸出一只手的样式，抓住我的一绺头发，灵就将我举到天地中间；在上帝的异象中，他带我到 耶路撒冷 朝北的内院门口，在那里有惹动妒忌的偶像的座位，它惹动了妒忌。
EZEK|8|4|看哪，在那里有 以色列 上帝的荣耀，形状与我在平原所见的一样。
EZEK|8|5|上帝对我说：“人子啊，你举目向北观看。”我就举目向北观看，看哪，祭坛门北边的门口有那惹动妒忌的偶像。
EZEK|8|6|他又对我说：“人子啊，你看见 以色列 家所做的吗？他们在这里做了极其可憎的事，使我远离我的圣所。你还要看见另有极其可憎的事。”
EZEK|8|7|他领我到院子门口。我观看，看哪，墙上有一个洞。
EZEK|8|8|他对我说：“人子啊，你要挖墙。”我就挖墙。看哪，有一扇门。
EZEK|8|9|他说：“你进去，看他们在这里所做可憎的恶事。”
EZEK|8|10|于是我进去看。看哪，四面墙上刻着各样爬行的动物、可憎的走兽和 以色列 家各样的偶像。
EZEK|8|11|以色列 家的七十个长老站在这些像前， 沙番 的儿子 雅撒尼亚 也站在其中，各人手拿他的香炉，烟云的香气上腾。
EZEK|8|12|他对我说：“人子啊，你看见 以色列 家的长老，暗中在自己偶像的房间里所做的吗？因为他们说：‘耶和华看不见我们；耶和华已经离弃这地。’”
EZEK|8|13|他又说：“你还要看见他们所做另外极其可憎的事。”
EZEK|8|14|他领我到耶和华殿朝北的门口。看哪，在那里有妇女们坐着，为 搭模斯 哭泣。
EZEK|8|15|他对我说：“人子啊，你看见了吗？你还要看见比这更可憎的事。”
EZEK|8|16|然后他领我到耶和华殿的内院。看哪，在耶和华殿门口、走廊和祭坛中间，约有二十五个人背向耶和华的殿，面向东方，向东拜太阳。
EZEK|8|17|他对我说：“人子啊，你看见了吗？ 犹大 家在这里行可憎的事还算为小吗？他们遍地行残暴，再三惹我发怒。看哪，他们手拿枝条举向鼻前 ！
EZEK|8|18|因此，我也要以愤怒行事。我的眼必不顾惜，也不可怜他们；他们虽在我耳边大声呼求，我还是不听。”
EZEK|9|1|他在我耳边大声喊叫，说：“上前来啊，惩罚这城的人，手中要各拿毁灭的兵器。”
EZEK|9|2|看哪，有六个人从朝北的 上门 而来，各人手里拿着致命的兵器；他们当中有一人身穿细麻衣，腰间系着文士用的墨盒。他们进来，站在铜的祭坛旁。
EZEK|9|3|在基路伯之上， 以色列 上帝的荣耀从那里上升，到殿的入口处。上帝召那身穿细麻衣、腰间系着墨盒的人前来。
EZEK|9|4|耶和华对他说：“你去走遍 耶路撒冷 全城，那些为城中所做可憎之事叹息哀哭的人，你要在他们额上做记号。”
EZEK|9|5|我耳中听见耶和华对其余的人说：“要跟随他走遍全城去击杀。你们的眼不要顾惜，也不要可怜他们。
EZEK|9|6|要将年老的、年轻的、少女、孩童和妇女，从我的圣所开始全都杀尽，只是不可挨近凡有记号的人。”于是他们从殿前的长老杀起。
EZEK|9|7|他对他们说：“要使这殿污秽，使院中遍满被杀的人。你们出去吧！”他们就出去，在城中击杀。
EZEK|9|8|他们击杀的时候，只剩我一人，我就脸伏在地上，呼喊说：“唉！主耶和华啊，你将愤怒倾倒在 耶路撒冷 ，岂要把 以色列 所剩余的人都灭绝吗？”
EZEK|9|9|他对我说：“ 以色列 家和 犹大 家的罪孽极其重大。遍地都有流血的事，满城有冤屈，因为他们说：‘耶和华已经离弃这地，他看不见我们。’
EZEK|9|10|因此，我的眼必不顾惜，也不可怜他们，要照他们所做的报应在他们头上。”
EZEK|9|11|看哪，那身穿细麻衣、腰间系着墨盒的人回覆这事说：“我已经照你所吩咐的做了。”
EZEK|10|1|我观看，看哪，在穹苍之中，也就是基路伯的头上，有蓝宝石的形状，仿佛宝座的形像显在他们上面。
EZEK|10|2|耶和华对那身穿细麻衣的人说：“你进到基路伯下面旋转的轮子中，从基路伯之间取出火炭装满两手掌，撒在城上。” 我亲眼看见他进去。
EZEK|10|3|那人进去的时候，基路伯站在殿的南边，云彩充满了内院。
EZEK|10|4|耶和华的荣耀从基路伯那里上升，到殿的入口处；殿内满布云彩，院子也充满了耶和华荣耀的光辉。
EZEK|10|5|基路伯翅膀的响声传到外院，好像全能上帝说话的声音。
EZEK|10|6|耶和华吩咐那身穿细麻衣的人说：“要从基路伯之间旋转的轮子中取火。”那人就进去站在一个轮子旁边。
EZEK|10|7|基路伯中的一个基路伯伸手到基路伯中间的火那里，取一些放在那身穿细麻衣人的手掌中，那人拿了就出去。
EZEK|10|8|在基路伯翅膀以下，显出有人手的样式。
EZEK|10|9|我又观看，看哪，这些基路伯的旁边有四个轮子。一个基路伯旁有一个轮子，另一个基路伯旁也有一个轮子；轮子的形状好像水苍玉石。
EZEK|10|10|至于四轮的形状，都是一个样式，好像轮中套轮。
EZEK|10|11|轮子行走的时候，向四方都能直行，行走时并不转弯。头转向何方，它们也随着向何方行走，行走时并不转弯。
EZEK|10|12|基路伯的全身，连背带手和翅膀，并轮子周围都布满眼睛。他们四个的轮子都是如此。
EZEK|10|13|我耳中听见这些轮子称为“旋转的轮”。
EZEK|10|14|基路伯各有四张脸：第一是基路伯的脸，第二是人的脸，第三是狮子的脸，第四是鹰的脸。
EZEK|10|15|基路伯升上去了；这就是我在 迦巴鲁河 边所看见的活物。
EZEK|10|16|基路伯行走，轮子也在旁边行走。基路伯展开翅膀，离地上升，轮子也不转离他们的旁边。
EZEK|10|17|基路伯站住，轮子也站住；基路伯上升，轮子也跟着上升，因为活物的灵在轮中。
EZEK|10|18|耶和华的荣耀离开殿的入口处，停在基路伯之上。
EZEK|10|19|基路伯展开翅膀，在我眼前离地上升；他们离去的时候，轮子在旁边，都停在耶和华殿的东门口。在他们上面有 以色列 上帝的荣耀。
EZEK|10|20|这是我在 迦巴鲁河 边所见的活物，他们在 以色列 上帝之下；因此我知道他们是基路伯。
EZEK|10|21|他们各有四张脸、四个翅膀，翅膀以下有人手的样式。
EZEK|10|22|至于他们脸的模样，以及身体的形像 ，正是我从前在 迦巴鲁河 边所看见的。他们各自往前直行。
EZEK|11|1|灵将我举起，带我到耶和华圣殿面向东方的东门。看哪，门口有二十五个人。我见其中有百姓的领袖 押朔 的儿子 雅撒尼亚 和 比拿雅 的儿子 毗拉提 。
EZEK|11|2|耶和华对我说：“人子啊，他们就是图谋罪孽，在这城中设计恶谋的人。
EZEK|11|3|他们说：‘盖房屋的时候尚未临近；这城是锅，我们是肉。’
EZEK|11|4|人子啊，因此你当说预言，说预言攻击他们。”
EZEK|11|5|耶和华的灵降在我身上，对我说：“你当说，耶和华如此说： 以色列 家啊，你们所说的，你们心里所想的，我都知道。
EZEK|11|6|你们在这城里大行屠杀，被杀的人遍满街道。
EZEK|11|7|所以主耶和华如此说：你们在城中杀的人是肉，这城是锅；你们却要从其中被带出去。
EZEK|11|8|你们怕刀剑，我却要使刀剑临到你们。这是主耶和华说的。
EZEK|11|9|我要把你们从这城中带出去，交在外邦人的手里，且要在你们中间施行审判。
EZEK|11|10|你们要仆倒在刀下；我必在 以色列 的边界审判你们，你们就知道我是耶和华。
EZEK|11|11|这城必不作你们的锅，你们也不作锅中的肉。我要在 以色列 的边界审判你们，
EZEK|11|12|你们就知道我是耶和华；因为你们不遵行我的律例，也不顺从我的典章，却随从你们四围列国的规条。”
EZEK|11|13|我正说预言的时候， 比拿雅 的儿子 毗拉提 死了。于是我脸伏在地，大声呼叫说：“唉！主耶和华啊，你要把 以色列 剩余的人都灭绝净尽吗？”
EZEK|11|14|耶和华的话临到我，说：
EZEK|11|15|“人子啊， 耶路撒冷 的居民对你的兄弟、你的本家、你的亲属、 以色列 全家所有的人说：‘你们远离耶和华吧！这地是赐给我们为业的。’
EZEK|11|16|所以你当说：‘主耶和华如此说：我虽将 以色列 全家远远流放到列国，使他们分散在列邦，我却要在他们所到的列邦，暂时作他们的圣所。’
EZEK|11|17|你当说：‘主耶和华如此说：我必从万民中召集你们，从分散的列邦中聚集你们，又将 以色列 地赐给你们。’
EZEK|11|18|他们到了那里，必从其中除掉一切可憎之物、可厌的事。
EZEK|11|19|我要使他们有合一的心，也要将新灵放在你们 里面，又从他们的肉体中除掉石心，赐给他们肉心，
EZEK|11|20|使他们顺从我的律例，谨守遵行我的典章。他们要作我的子民，我要作他们的上帝。
EZEK|11|21|至于那些心中随从可憎之物、可厌的事的人，我必照他们所做的报应在他们头上。这是主耶和华说的。”
EZEK|11|22|于是，基路伯展开翅膀，轮子都在他们旁边；在他们上面有 以色列 上帝的荣耀。
EZEK|11|23|耶和华的荣耀从城中上升，停在城东的那座山上。
EZEK|11|24|灵将我举起，在异象中上帝的灵将我带回 迦勒底 地，到被掳的人那里；之后我所见的异象就离我上升去了。
EZEK|11|25|我就把耶和华指示我的一切事都说给被掳的人听。
EZEK|12|1|耶和华的话临到我，说：
EZEK|12|2|“人子啊，你住在悖逆之家中；他们有眼可看却看不见，有耳可听却听不到，因为他们是悖逆之家。
EZEK|12|3|所以人子啊，你要收拾被掳时需用的物件，白天在他们眼前离去，在他们眼前离开你所住的地方，移到别处去；他们虽是悖逆之家，或者可以领悟。
EZEK|12|4|你要白天在他们眼前拿出你被掳时需用的物件。到了晚上，要在他们眼前离去，像被掳的人离去一样。
EZEK|12|5|你要在他们眼前挖通墙壁，从其中将物件带出去 。
EZEK|12|6|到天黑时，在他们眼前背在肩上带走 ，并要蒙住脸看不见地，因为我要使你成为 以色列 家的预兆。”
EZEK|12|7|我就照着所吩咐的去做，白天拿出被掳时需用的物件。到了晚上，用手挖通墙壁；天黑的时候，在他们眼前背在肩上带走。
EZEK|12|8|次日早晨，耶和华的话临到我，说：
EZEK|12|9|“人子啊， 以色列 家，就是那悖逆之家，岂不是问你说：‘你在做什么呢？’
EZEK|12|10|你要对他们说：‘主耶和华如此说：这是关乎 耶路撒冷 君王和其中 以色列 全家的默示。’
EZEK|12|11|你要说：‘我是你们的预兆：我怎样做，他们所遭遇的也必这样，他们必被掳去，作俘虏。’
EZEK|12|12|他们中间的君王也必在天黑时把物件背在肩上带走。他们要挖通墙壁，从其中带出去 。他必蒙住脸，眼看不见地。
EZEK|12|13|我要把我的网撒在他身上，他就被我的罗网缠住。我要带他到 迦勒底 人之地的 巴比伦 ；他没有看见那地，就死在那里。
EZEK|12|14|我要把四围帮助他的和他所有的军队分散到四方 ，也要拔刀追赶他们。
EZEK|12|15|我把他们驱逐到列国，分散在列邦的时候，他们就知道我是耶和华。
EZEK|12|16|我却要留下他们当中几个人得免刀剑、饥荒、瘟疫，使他们在所到的列国述说自己所做一切可憎的事；他们就知道我是耶和华。”
EZEK|12|17|耶和华的话临到我，说：
EZEK|12|18|“人子啊，你吃饭时必战抖，喝水时必惊惶忧虑。
EZEK|12|19|你要对这地的百姓说：主耶和华论 以色列 地的 耶路撒冷 居民如此说，他们吃饭时必忧虑，喝水时必惊惶，因其中居民所行残暴的事，这地必然荒废，一无所存。
EZEK|12|20|有人居住的城镇必变为废墟，地必荒凉；你们就知道我是耶和华。”
EZEK|12|21|耶和华的话临到我，说：
EZEK|12|22|“人子啊，在 以色列 地你们怎么有这俗语说：‘日子延长，一切异象却落了空’呢？
EZEK|12|23|你要告诉他们说：‘主耶和华如此说：我必令这俗语止息， 以色列 中不再有人引用这俗语。’你却要对他们说：‘日子临近，一切的异象都必应验。’
EZEK|12|24|从此以后， 以色列 家不再有虚假的异象和奉承的占卜。
EZEK|12|25|我─耶和华说话，所说的必定实现，不再耽延。你们这悖逆之家啊，你们在世的日子，我所说的话必定实现。这是主耶和华说的。”
EZEK|12|26|耶和华的话临到我，说：
EZEK|12|27|“人子，看哪， 以色列 家的人说：‘他所见的异象是许多日子以后的事，所说的预言是指着遥远的时候。’
EZEK|12|28|所以你要对他们说：‘主耶和华如此说：我的话不再有一句耽延，我所说的话必定实现。’这是主耶和华说的。”
EZEK|13|1|耶和华的话临到我，说：
EZEK|13|2|“人子啊，你要说预言，攻击 以色列 中说预言的先知，对那些随心说预言的人说：‘你们当听耶和华的话。’”
EZEK|13|3|主耶和华如此说：“祸哉！那些愚顽的先知，随从自己的心意，却一无所见
EZEK|13|4|以色列 啊，你的先知好像废墟中的狐狸，
EZEK|13|5|没有上去堵住缺口，也没有为 以色列 家重修城墙，使它在耶和华的日子来临时，可以在战争中站得住。
EZEK|13|6|他们看见的是虚假，是谎诈的占卜，说是耶和华说的；其实耶和华并没有差遣他们，他们却指望那话必站立得住。
EZEK|13|7|你们岂不是见了虚假的异象吗？岂不是说了谎诈的占卜吗？你们说，这是耶和华说的，其实我没有说过。”
EZEK|13|8|所以主耶和华如此说：“因你们说的是虚假，见的是谎诈，所以，看哪，我要敌对你们。这是主耶和华说的。
EZEK|13|9|我的手必攻击那见虚假异象、用谎诈占卜的先知，他们必不列在我百姓的会中，不录在 以色列 家的名册上，也不能进入 以色列 地；你们就知道我是主耶和华。
EZEK|13|10|他们诱惑我的百姓，说：‘平安！’其实没有平安，就像有人筑墙壁，看哪，他们倒去粉刷它。
EZEK|13|11|所以你要对那些粉刷的人说：‘墙要倒塌，暴雨漫过。你们大冰雹啊，要降下 ，狂风要吹裂这墙。’
EZEK|13|12|看哪，这墙倒塌，人岂不是要问你们说：‘你们所粉刷的在哪里呢？’”
EZEK|13|13|所以主耶和华如此说：“我要发怒，使狂风吹裂它，在怒中令暴雨漫过，又发怒降下大冰雹，毁坏它。
EZEK|13|14|我要这样拆毁你们那粉饰的墙，把它夷为平地，以致根基露出；墙一倒塌，你们也要在其中灭亡。你们就知道我是耶和华。
EZEK|13|15|我要对墙和粉刷它的人发尽我的愤怒，我 要对你们说：‘墙没有了！粉刷它的人也没有了！’
EZEK|13|16|这就是 以色列 的先知，他们指着 耶路撒冷 说预言，见到这城平安的异象，其实没有平安。这是主耶和华说的。”
EZEK|13|17|“你，人子啊，要面向你百姓中随心说预言的妇女们，说预言攻击她们，
EZEK|13|18|说，主耶和华如此说：‘这些妇女有祸了！她们为众人的手腕缝驱邪带，替身材高矮不同的人做头巾，为要猎取人的性命。难道你们要猎取我百姓的性命，使自己存活吗？
EZEK|13|19|你们为几把大麦、几块饼，在我的百姓中亵渎我，对那肯听谎言的百姓说谎言，让不该死的人死，让不该活的人活。’”
EZEK|13|20|所以主耶和华如此说：“看哪，我要对付你们那用以猎取人，如猎飞鸟般的驱邪带。我要把驱邪带从你们的手腕扯去，释放那些如飞鸟被你们猎取的人。
EZEK|13|21|我也必撕裂你们的头巾，救我百姓脱离你们的手，使他们不再被猎取，落在你们手中；你们就知道我是耶和华。
EZEK|13|22|我未曾使义人伤心，你们却以谎话使他伤心，且又坚固恶人的手，不使他回转离开恶道得以存活。
EZEK|13|23|所以，你们必不再看见虚假的异象，也不再行占卜的事；我要救我的百姓脱离你们的手；你们就知道我是耶和华。”
EZEK|14|1|有几个 以色列 的长老到我这里来，坐在我面前。
EZEK|14|2|耶和华的话临到我，说：
EZEK|14|3|“人子啊，这些人在心中设立偶像，把陷自己于罪的绊脚石放在面前，我真的能让他们求问吗？
EZEK|14|4|所以你要告诉他们，对他们说：‘主耶和华如此说： 以色列 家的人，凡在心中设立偶像，把陷自己于罪的绊脚石放在面前，却来到先知那里的，我─耶和华在他所求的事上，必因他拜许多偶像向他施行报应 ，
EZEK|14|5|为要夺回 以色列 家的心，他们全都拜偶像，与我疏远了。’
EZEK|14|6|“所以你要对 以色列 家说：‘主耶和华如此说：回转吧！回转离开你们的偶像，转脸离开一切可憎的事。’
EZEK|14|7|因为 以色列 家的人，或在 以色列 中寄居的外人，凡与我隔绝，在心中设立偶像，把陷自己于罪的绊脚石放在面前，却来到先知那里，要为自己的事求问我的，我─耶和华必亲自报应他。
EZEK|14|8|我要向那人变脸，使他成为警戒和笑柄，并且我要把他从我民中剪除；你们就知道我是耶和华。
EZEK|14|9|先知若被骗说了一句预言，是我─耶和华骗了那先知，我要伸手攻击他，把他从我百姓 以色列 中除灭。
EZEK|14|10|他们必担当自己的罪孽。先知的罪孽和求问之人的罪孽都一样，
EZEK|14|11|使 以色列 家不再走迷离开我，也不再因各样的罪过玷污自己，却要作我的子民，我也作他们的上帝。这是主耶和华说的。”
EZEK|14|12|耶和华的话临到我，说：
EZEK|14|13|“人子啊，若有一国犯罪干犯我，我也伸手攻击它，断绝他们粮食的供应，使饥荒临到那地，将人与牲畜从其中剪除；
EZEK|14|14|虽有 挪亚 、 但以理 、 约伯 这三人在那里，他们只能因自己的义救自己的命。这是主耶和华说的。
EZEK|14|15|我若使恶兽经过那地，大肆蹂躏，使地荒凉，以致因这些兽，人都不得经过；
EZEK|14|16|虽有这三人在其中，主耶和华说：我指着我的永生起誓，他们不能救儿子女儿，只有他们自己可以得救，那地仍然荒凉。
EZEK|14|17|或者我使刀剑临到那地，说：‘让刀剑穿越那地’，以致我把人与牲畜从其中剪除；
EZEK|14|18|虽有这三人在其中，主耶和华说：我指着我的永生起誓，他们不能救儿子女儿，只有他们自己可以得救。
EZEK|14|19|或者我叫瘟疫流行那地，把我的愤怒带着血倾在其中，好使人与牲畜从其中剪除；
EZEK|14|20|虽有 挪亚 、 但以理 、 约伯 在那里，主耶和华说：我指着我的永生起誓，他们不能救儿子女儿，只能因自己的义救自己的命。
EZEK|14|21|“主耶和华如此说：我若将这四样大灾，就是刀剑、饥荒、恶兽、瘟疫降在 耶路撒冷 ，将人与牲畜从其中剪除，岂不是更严重吗？
EZEK|14|22|看哪，在那里必有幸免于难的人带着儿子女儿；看哪，他们来到你们这里；你们看见他们的所作所为，就会因我降给 耶路撒冷 的灾祸，因我降给它的一切，得到安慰。
EZEK|14|23|你们因看见他们的所作所为，得到安慰，就会知道我在 耶路撒冷 所做的并非毫无缘故。这是主耶和华说的。”
EZEK|15|1|耶和华的话临到我，说：
EZEK|15|2|“人子啊，葡萄树比一切其他的树，就是树林里众树木的树枝，有什么长处呢？
EZEK|15|3|可以从其中取木料来做工吗？人可以拿来做钉子，挂东西在上面吗？
EZEK|15|4|看哪，它已经抛在火中当柴烧，火既烧了两头，中间也烧焦了，它还有什么用处呢？
EZEK|15|5|看哪，它完整的时候尚且不能拿来做工，何况被火烧焦了，还能拿来做工吗？
EZEK|15|6|所以，主耶和华如此说：我怎样使林中树里的葡萄树在火中当柴烧，我也必照样对待 耶路撒冷 的居民。
EZEK|15|7|我必向他们变脸；他们虽从火中逃出来，火仍要烧灭他们。我向他们变脸的时候，你们就知道我是耶和华。
EZEK|15|8|我必使这地荒凉，因为他们做了背叛的事。这是主耶和华说的。”
EZEK|16|1|耶和华的话临到我，说：
EZEK|16|2|“人子啊，你要使 耶路撒冷 知道它那些可憎的事。
EZEK|16|3|你要说，主耶和华对 耶路撒冷 如此说：你的根源，你的出身，是在 迦南 地；你的父亲是 亚摩利 人，母亲是 赫 人。
EZEK|16|4|论到你出世的景况，在你出生的日子没有人为你断脐带，也没有用水清洗，使你洁净；没有人撒盐在你身上，也没有人用布包你。
EZEK|16|5|没有人顾惜你，为你做一件这样的事来可怜你。你却被扔在田野上面，因你出生的日子就被厌恶。
EZEK|16|6|“我从你旁边经过，见你在血中打滚，就对你说：‘你虽在血中，却要活下去！’我又说：‘你虽在血中，却要活下去！’
EZEK|16|7|我使你成长如田间所生长的；你就渐长，美而又美 ，两乳成形，头发秀长，但你仍然赤身露体。
EZEK|16|8|“我从你旁边经过看见你，看哪，正是你渴慕爱情的时候，我就用我衣服的边搭在你身上，遮盖你的赤体；又向你起誓，与你立约，你就归我。这是主耶和华说的。
EZEK|16|9|那时我用水洗你，洗净你身上的血，又用油抹你。
EZEK|16|10|我使你身穿锦绣衣裳，脚穿海狗皮鞋，用细麻布裹着你，精致衣料披在你身上。
EZEK|16|11|我用首饰打扮你：我把手镯戴在你手上，项链在你颈上，
EZEK|16|12|我也把环子戴在你鼻上，耳环在你耳上，华冠在你头上。
EZEK|16|13|这样，你就有金银的首饰，穿的是细麻衣和精致衣料，以及锦绣衣裳；吃的是细面、蜂蜜和油。你也极其美貌，配登王后之位。
EZEK|16|14|你美貌的名声传到列国，因我加给你荣华，使你完美。这是主耶和华说的。
EZEK|16|15|“只是你仗着自己美貌，又凭着你的名声行淫。你向路人纵情淫乱，你的美貌就属于他的了 。
EZEK|16|16|你拿你的衣服为自己做成彩色丘坛，在其上行淫。这样的事本不该有，以后也不该发生。
EZEK|16|17|你拿我所赐给你的那些美丽的金银宝物，为自己制造男性的偶像，与它们行淫；
EZEK|16|18|你拿你的锦绣衣裳为它们披上，把我的膏油和香料摆在它们面前；
EZEK|16|19|你把我赐给你的食物，就是我赐给你享用的细面、油和蜂蜜，都摆在它们面前作为馨香的供物。事情就是这样。这是主耶和华说的。
EZEK|16|20|你拿你为我所生的儿女献给它们吞噬。你的淫乱岂是小事？
EZEK|16|21|你竟把我的儿女杀了，使他们经火献给它们！
EZEK|16|22|你做这一切可憎和淫乱的事，并未追念你幼年的日子，那时你赤身露体，在血中打滚。”
EZEK|16|23|“你有祸了！你有祸了！这是主耶和华说的。你做这一切恶事之后，
EZEK|16|24|又为自己建造土墩，在各广场上筑起高台。
EZEK|16|25|你在各个街头建造高台，使你的美貌变为可憎；又向所有过路的人招手 ，多行淫乱。
EZEK|16|26|你也和你那放纵情欲的邻邦 埃及 人行淫，增添你的淫乱，惹我发怒。
EZEK|16|27|看哪，我伸手攻击你，减少你的福分，却将你交给恨恶你的 非利士 人 ，让他们任意待你。他们为你的淫行也感到羞耻。
EZEK|16|28|你尚且不满意，又与 亚述 人行淫，但与他们行淫之后，仍不满足；
EZEK|16|29|于是你与那称为贸易之地的 迦勒底 多行淫乱，即使这样，你仍不满足。
EZEK|16|30|“你的心何等脆弱！这是主耶和华说的。你做这一切事，都是不知羞耻的妓女所做的，
EZEK|16|31|在各个街头建造土墩，在各广场上筑高台；但你藐视行淫的赏金，又不像妓女。
EZEK|16|32|你这行淫的妻子啊，竟然接外人，替代丈夫。
EZEK|16|33|凡妓女都是得人赠礼，你反倒馈赠你所爱的人，倒贴他们，使他们从四围来与你行淫。
EZEK|16|34|你的淫行与其他妇女相反，不是人要求与你行淫；是你给人赏金，不是人给你赏金；你是相反的。”
EZEK|16|35|“你这妓女啊，要听耶和华的话。
EZEK|16|36|主耶和华如此说：因你放纵情欲，露出下体，与你所爱的行淫，因你敬拜一切可憎的偶像，就像 自己儿女的血献给它们，
EZEK|16|37|所以，看哪，我要聚集所有与你交欢的情人，不论是你所爱的或你所恨的，聚集他们从四围到你那里来；我要在他们面前暴露你的下体，使他们看尽你的下体。
EZEK|16|38|我也要审判你，如审判淫妇和流人血的妇女一样。我要在愤怒和妒忌中使流血的罪归到你身上。
EZEK|16|39|我要把你交在他们手中；他们必拆毁你的土墩，毁坏你的高台，剥去你的衣服，夺取你美丽的宝物，留下你赤身露体。
EZEK|16|40|他们必聚集众人攻击你，用石头打死你，用刀剑刺透你，
EZEK|16|41|用火焚烧你的房屋，在许多妇女眼前审判你。我必使你不再行淫，你也不再给赏金。
EZEK|16|42|我止息了向你所发的愤怒，我的妒忌也离开了你；这样，我就平静，不再恼怒。
EZEK|16|43|因你不追念幼年的日子，反而在这一切的事上惹我发烈怒，所以，看哪，我必照你所做的报应在你头上。在你一切可憎的事上，你不是还行了淫乱吗？这是主耶和华说的。”
EZEK|16|44|“看哪，凡说俗语的必用这俗语攻击你，说：‘有其母必有其女。’
EZEK|16|45|你实在是你母亲的女儿，厌弃丈夫和儿女；你也是你姊妹的姊妹，厌弃丈夫和儿女。你的母亲是 赫 人，父亲是 亚摩利 人。
EZEK|16|46|你的姊姊是 撒玛利亚 ，她和她的女儿们住在你北边；你的妹妹是 所多玛 ，她和她的女儿们住在你南边。
EZEK|16|47|你不只效法她们的行为，照她们可憎的事去做，不消多时 ，你所做的一切就比她们更恶。
EZEK|16|48|主耶和华说：我指着我的永生起誓，你的妹妹 所多玛 与她的女儿们并未做你和你女儿们所做的事。
EZEK|16|49|看哪，你的妹妹 所多玛 的罪孽是这样：她和她的女儿们都骄傲，粮源充足，大享安逸，却不扶持困苦和贫穷人的手。
EZEK|16|50|她们狂傲，在我面前做可憎的事，我看见了就把她们除掉。
EZEK|16|51|撒玛利亚 所犯的罪不及你的一半，你所做可憎的事比她更多；比起你所做这一切可憎的事，你的姊妹倒显为义。
EZEK|16|52|你既为你的姊妹辩护，就要担当自己的羞辱。因你所犯的罪比她们更可憎，她们比你倒显为义；你既使你的姊妹显为义，就要抱愧，担当自己的羞辱。”
EZEK|16|53|“我必使她们被掳的归回，使 所多玛 和她的女儿们、 撒玛利亚 和她的女儿们，并与你一起被掳的都归回；
EZEK|16|54|好使你担当自己的羞辱，为所做的一切抱愧，让她们得到安慰。
EZEK|16|55|你的妹妹 所多玛 和她的女儿们必回复原状； 撒玛利亚 和她的女儿们必回复原状；你和你的女儿们也必回复原状。
EZEK|16|56|在你骄傲的日子，你的妹妹 所多玛 岂不是你口中的笑柄吗？
EZEK|16|57|在你的恶行显露以前，那受了凌辱的 亚兰 女儿们和 亚兰 四围 非利士 的女儿们，都在四围藐视你。
EZEK|16|58|耶和华说：你的淫荡和可憎之事，你自己要担当。”
EZEK|16|59|“主耶和华如此说：你这轻看誓言而背约的，我必照你所做的报应你。
EZEK|16|60|然而我要追念在你幼年时我与你所立的约，也要与你立定永约。
EZEK|16|61|当你接纳你的姊姊和妹妹时，你要追念你所行的，自觉惭愧；并且我要将她们赏给你做女儿，却不是按着我与你所立的约。
EZEK|16|62|我要坚定与你所立的约，你就知道我是耶和华，
EZEK|16|63|使你在我赦免你一切恶行时，心中追念，自觉惭愧，又因羞辱就不再开口。这是主耶和华说的。”
EZEK|17|1|耶和华的话临到我，说：
EZEK|17|2|“人子啊，你要向 以色列 家出谜语，设比喻，
EZEK|17|3|说，主耶和华如此说：有一只大鹰，翅膀大，翎毛长，羽毛丰满，色彩缤纷；它飞到 黎巴嫩 ，啄去香柏树梢，
EZEK|17|4|啄断它顶端的嫩枝，叼到贸易之地，放在商业城中。
EZEK|17|5|它又从这地取了一些种子，种在肥沃的田里，栽于丰沛的水源旁，如种植柳树。
EZEK|17|6|它渐渐生长，成为低矮蔓生的葡萄树；树枝伸向那鹰，根部在它下面。这样，它就长成了一棵葡萄树，生出枝子，长出枝干。
EZEK|17|7|“有一只 大鹰，翅膀大，羽毛多。看哪，葡萄树从栽种它的苗圃向这鹰伸出根来，长出枝子，期盼从它得到浇灌。
EZEK|17|8|这棵树栽于肥田丰沛的水源旁，原是为了生枝、结果，成为佳美的葡萄树。
EZEK|17|9|你要说，主耶和华如此说：这棵葡萄树岂能发旺呢？鹰岂不拔出它的根来，摘光它的果子，使它枯干，连长出的嫩叶都枯萎了吗？要把它连根拔除，并不需要费大力或动用许多人。
EZEK|17|10|看哪，葡萄树虽然栽种了，岂能发旺呢？一经东风击打，岂不全然枯干了吗？它必在生长的苗圃中枯干了。”
EZEK|17|11|耶和华的话临到我，说：
EZEK|17|12|“你要对那悖逆之家说：你们不知道这些事是什么意思吗？你要这样说，看哪， 巴比伦 王曾到 耶路撒冷 ，把其中的君王和官长带到 巴比伦 去，
EZEK|17|13|又从 以色列 王室后裔中选取一人，与他立约，令他发誓，又掳走国中有势力的人，
EZEK|17|14|使王国衰弱，不再强盛，只能靠守盟约方得生存。
EZEK|17|15|他却背叛 巴比伦 王，差派使者前往 埃及 ，要求 埃及 人给他马匹和许多人。他岂能亨通呢？这样做的人岂能逃脱呢？他背了约岂能逃脱呢？
EZEK|17|16|主耶和华说：我指着我的永生起誓，他定要死在 巴比伦 ，就是 巴比伦 王所在之处；因为 巴比伦 王立他为王，他竟轻看向王所起的誓，背弃王与他所立的约。
EZEK|17|17|当敌人建土堆，筑堡垒，要歼灭许多人时，法老虽有强大军队和大批人马，在战场上还是不能帮助他。
EZEK|17|18|他轻看誓言，背弃盟约，看哪，虽已投降 ，却又做这一切的事，他必不能逃脱。
EZEK|17|19|所以主耶和华如此说：我指着我的永生起誓，他既轻看我的誓言，背弃我的约，我必使这罪归到他头上。
EZEK|17|20|我要把我的网撒在他身上，他就被我的罗网缠住。我要带他到 巴比伦 ，在那里因他背叛我的罪惩罚他。
EZEK|17|21|所有逃跑的 军队必倒在刀下；剩余的也必分散四方 。你们就知道说这话的是我─耶和华。”
EZEK|17|22|主耶和华如此说：“我要从香柏树高高的树梢摘取并栽上，从顶端的嫩枝中折下一嫩枝，栽于极高的山上，
EZEK|17|23|栽在 以色列 高处的山上。它就生枝、结果，成为高大的香柏树，各类飞禽中的鸟都来宿在其下，宿在枝子的荫下 。
EZEK|17|24|田野的树木因此就知道是我─耶和华使高树矮小，使矮树高大，使绿树枯干，使枯树发旺。我─耶和华说了这话，就必成就。”
EZEK|18|1|耶和华的话又临到我，说：
EZEK|18|2|“你们在 以色列 地何以有这俗语，‘父亲吃了酸葡萄，儿子牙齿就酸倒’呢？
EZEK|18|3|主耶和华说：我指着我的永生起誓，你们在 以色列 必不再引用这俗语。
EZEK|18|4|看哪，所有的生命都是属我的；父亲的生命怎样属我，儿子的生命也照样属我；然而犯罪的，他必定死。
EZEK|18|5|“人若是公义，行公平公义的事：
EZEK|18|6|未曾在山上吃祭物，未曾向 以色列 家的偶像举目；未曾污辱邻舍的妻，也未曾在妇人的经期间亲近她；
EZEK|18|7|未曾亏负人，而是将欠债之人的抵押品还给他；未曾抢夺人的物件，却把食物给饥饿的人吃，把衣服给赤身的人穿；
EZEK|18|8|未曾向人取利息，也未曾索取高利，反倒缩手不作恶，在人与人之间施行诚实的判断；
EZEK|18|9|遵行我的律例，谨守我的典章，按诚实行事 ；这人是公义的，必要存活。这是主耶和华说的。
EZEK|18|10|“他若生了儿子，儿子作强盗，流人的血，作父亲的 虽然未犯此过，儿子却对弟兄 行了以上所说的恶，在山上吃祭物，污辱邻舍的妻；
EZEK|18|11|
EZEK|18|12|亏负困苦和贫穷的人，抢夺别人的物件，不归还抵押品，却向偶像举目，做可憎的事；
EZEK|18|13|向人取利息，索取高利，这人岂能存活呢？他不能存活。他因做这一切可憎的事，必要死亡，他的血要归到自己身上。
EZEK|18|14|“看哪，他若生了儿子，儿子见父亲所犯的一切罪，他见了，却不照样去做；
EZEK|18|15|他未曾在山上吃祭物，未曾向 以色列 家的偶像举目，未曾污辱邻舍的妻；
EZEK|18|16|也未曾亏负人，未曾取人的抵押品，未曾抢夺人的物件，却把食物给饥饿的人吃，把衣服给赤身的人穿，
EZEK|18|17|缩手不害困苦人，未曾向人索取利息或高利；反倒顺从我的典章，遵行我的律例；如此，他必不因父亲的罪孽死亡，定要存活。
EZEK|18|18|至于他父亲，因为施行欺压，抢夺弟兄，在百姓中行不善，看哪，他必因自己的罪孽死亡。
EZEK|18|19|“你们还说：‘儿子为什么不担当父亲的罪孽呢？’儿子若行公平公义的事，谨守遵行我一切的律例，他必要存活。
EZEK|18|20|惟有犯罪的，却必死亡。儿子不担当父亲的罪孽，父亲也不担当儿子的罪孽。义人的善果要归自己，恶人的恶报也要归自己。
EZEK|18|21|“恶人若回转离开所做的一切罪恶，谨守我的一切律例，行公平公义的事，他必要存活，不致死亡。
EZEK|18|22|他所犯的一切罪过都不被记念；他因所行的义，必要存活。
EZEK|18|23|恶人死亡，岂是我所喜悦的呢？我岂不是喜悦他回转离开所行的道而存活吗？这是主耶和华说的。
EZEK|18|24|至于义人，他若转离义行而作恶，照着恶人所做一切可憎的事去做，岂能存活呢？他所行的一切义都不被记念；反而因所行的恶、所犯的罪死亡。
EZEK|18|25|“你们却说：‘主的道不公平！’ 以色列 家啊，你们要听，我的道不公平吗？你们的道不是不公平吗？
EZEK|18|26|义人若转离义行而作恶，他就因这些恶而死亡。他要死在他所作的恶中。
EZEK|18|27|恶人若回转离开所行的恶，行公平公义的事，他必救自己的命；
EZEK|18|28|因为他省察，回转离开所犯的一切罪过，他必要存活，不致死亡。
EZEK|18|29|以色列 家还说：‘主的道不公平！’ 以色列 家啊，我的道不公平吗？你们的道不是不公平吗？
EZEK|18|30|所以， 以色列 家啊，我必按你们各人所做的审判你们。当回转，回转离开你们一切的罪过，免得罪孽成为你们的绊脚石。这是主耶和华说的。
EZEK|18|31|你们要把所犯的一切罪过尽行抛弃，为自己造一个新的心和新的灵。 以色列 家啊，你们为什么要死呢？
EZEK|18|32|我不喜欢有任何人死亡，所以你们当回转，要存活！这是主耶和华说的。”
EZEK|19|1|你当为 以色列 的领袖们唱哀歌，
EZEK|19|2|说： 你的母亲在狮子中 是怎样的母狮呢？ 它蹲伏在少壮狮子中， 养育小狮子。
EZEK|19|3|它养大了其中一只小狮子， 成了少壮狮子， 学会抓食， 它就吃人。
EZEK|19|4|列国听见了就把它逮住在他们的坑里， 用钩子拉它到 埃及 地去。
EZEK|19|5|母狮见自己等候， 期望落空， 就从小狮子中取一只 ， 养为少壮狮子；
EZEK|19|6|它在众狮子中徜徉， 长大成为少壮狮子， 学会抓食， 它就吃人。
EZEK|19|7|它拆毁他们的宫殿 ， 使他们的城镇变为废墟； 因它咆哮的声音， 遍地和其中所充满的都荒废了。
EZEK|19|8|于是四围列国 从各省前来攻击它， 把网撒在它身上， 把它逮住在他们的坑里。
EZEK|19|9|他们又用钩子钩住它，把它放入笼中， 带到 巴比伦 王那里， 把它押进城堡， 以色列 山上就不再听见它的声音。
EZEK|19|10|你的母亲如葡萄树， 在葡萄园中 ， 栽于水边，因为水多， 就多结果子，多生枝子；
EZEK|19|11|它长出坚固的枝干， 可作统治者的权杖。 这枝干高举在茂密的树枝中， 可见树身高大，枝子繁多。
EZEK|19|12|但在烈怒中它被拔出，摔在地上； 东风吹干其果子， 那坚固的枝干因折断而枯干， 被火烧毁；
EZEK|19|13|如今这葡萄树移植于旷野， 在干旱无水之地，
EZEK|19|14|火从枝干中发出， 烧灭它的枝条和它的果子 ， 以致不再有坚固的枝干， 可作统治者的权杖。 这是哀伤之歌，成为一首哀歌。
EZEK|20|1|第七年五月初十，有 以色列 的几个长老前来求问耶和华，坐在我面前。
EZEK|20|2|耶和华的话临到我，说：
EZEK|20|3|“人子啊，你要告诉 以色列 的长老，对他们说，主耶和华如此说：你们来是为求问我吗？主耶和华说：我指着我的永生起誓，我必不让你们求问。
EZEK|20|4|人子啊，你要审问他们吗？你要审问吗？你当使他们知道他们祖先那些可憎的事；
EZEK|20|5|你要对他们说，主耶和华如此说：当日我拣选 以色列 ，对 雅各 家的后裔起誓，在 埃及 地向他们显现，起誓说：我是耶和华─你们的上帝；
EZEK|20|6|那日我向他们起誓，要领他们出 埃及 地，到我为他们所找到的流奶与蜜之地，就是全地中最美好之地。
EZEK|20|7|我对他们说，你们各人要抛弃眼中所喜爱的可憎之物，不可用 埃及 的偶像玷污自己。我是耶和华─你们的上帝。
EZEK|20|8|他们却悖逆我，不肯听从我，不抛弃他们眼中所喜爱的可憎之物，离弃 埃及 的偶像。 “我就说，在 埃及 地，我要把我的愤怒倾倒在他们身上，向他们发尽我的怒气。
EZEK|20|9|我这么做是为了我名的缘故，免得我的名在他们所居住之列国眼中被亵渎；我曾在这些列国眼前向他们显现，领他们出了 埃及 地。
EZEK|20|10|我领他们出 埃及 地，带他们到旷野。
EZEK|20|11|我将我的律例赐给他们，将我的典章指示他们；人若遵行就必因此存活。
EZEK|20|12|我将我的安息日赐给他们，在我与他们中间作记号，让他们知道我─耶和华是使他们分别为圣的。
EZEK|20|13|以色列 家却在旷野中悖逆我，不顺从我的律例，厌弃我的典章；人若遵行就必因此存活。他们却大大干犯我的安息日。 “因此我说，我要在旷野把我的愤怒倾倒在他们身上，灭绝他们。
EZEK|20|14|我这么做是为了我名的缘故，免得我的名在列国眼中被亵渎，因为在这些列国眼前我领了他们出来。
EZEK|20|15|并且我在旷野向他们起誓，必不领他们进入我所赐的流奶与蜜之地，就是全地中最美好之地；
EZEK|20|16|因为他们厌弃我的典章，不顺从我的律例，干犯我的安息日，他们的心随从自己的偶像。
EZEK|20|17|虽然如此，我的眼仍顾惜他们，不毁灭他们，不在旷野把他们灭绝净尽。
EZEK|20|18|“我在旷野对他们的儿女说：‘不要遵行你们祖先的律例，不要谨守他们的规条，也不要用他们的偶像玷污自己。
EZEK|20|19|我是耶和华─你们的上帝，你们要顺从我的律例，谨守遵行我的典章，
EZEK|20|20|且以我的安息日为圣。这日必在我与你们中间作记号，使你们知道我是耶和华─你们的上帝。’
EZEK|20|21|只是他们的儿女悖逆我，不顺从我的律例，也不谨守遵行我的典章；人若遵行就必因此存活。他们却干犯我的安息日。 “因此我说，我要在旷野把我的愤怒倾倒在他们身上，向他们发尽我的怒气。
EZEK|20|22|但我却缩手而未如此行；我这么做是为了我名的缘故，免得我的名在列国眼中被亵渎，因为在这些列国眼前我领了他们出来。
EZEK|20|23|并且我在旷野向他们起誓，要把他们驱散到列国，分散在列邦；
EZEK|20|24|因为他们不遵行我的典章，厌弃我的律例，干犯我的安息日，眼目向着他们祖先的偶像。
EZEK|20|25|我也任他们遵行那无益的律例，随从那不能使人存活的规条。
EZEK|20|26|他们使所有头生的经火，我就任凭他们在这供物上玷污自己；我令他们惊恐，他们就知道我是耶和华。
EZEK|20|27|“人子啊，你要告诉 以色列 家，对他们说，主耶和华如此说：你们的祖先在背叛我的事上再次亵渎了我；
EZEK|20|28|我领他们到我起誓应许赐给他们的地，他们看见各高冈、各茂密的树，就在那里献祭，献上惹我发怒的供物，也在那里焚烧馨香的祭，献浇酒祭。
EZEK|20|29|我就对他们说：你们去的那丘坛叫什么呢？它名叫 巴麻 ，直到今日。
EZEK|20|30|所以你要对 以色列 家说，主耶和华如此说：你们仍要照你们祖先所做的玷污自己吗？还要照他们可憎的事行淫吗？
EZEK|20|31|当你们献上供物，使你们儿子经火的时候，你们仍用各样的偶像玷污自己，直到今日。 以色列 家啊，我岂能让你们求问呢？主耶和华说：我指着我的永生起誓，我必不让你们求问。
EZEK|20|32|“你们说：‘我们要像列国和列邦的宗族一样，去事奉木头与石头。’你们所起的心意万不能成就。”
EZEK|20|33|“主耶和华说：我指着我的永生起誓，我要作王，用大能的手和伸出的膀臂，并倾倒出来的愤怒治理你们。
EZEK|20|34|我必用大能的手和伸出的膀臂，并倾倒出来的愤怒，把你们从万民中领出来，从被赶散到的列邦聚集你们。
EZEK|20|35|我必带你们到万民的旷野，在那里当面审判你们。
EZEK|20|36|我怎样在 埃及 地的旷野审判你们的祖先，也必照样审判你们。这是主耶和华说的。
EZEK|20|37|我要使你们从杖下经过，按着约的拘束 带领你们。
EZEK|20|38|我必从你们中间除尽叛逆和得罪我的人；我将他们从所寄居的地方领出来，他们却不得进入 以色列 地，你们就知道我是耶和华。
EZEK|20|39|“你们， 以色列 家啊，主耶和华如此说：你们若不听从我，从今以后就让各人去事奉他的偶像吧，只是不可再以你们的供物和偶像亵渎我的圣名。
EZEK|20|40|“在我的圣山，就是 以色列 高处的山， 以色列 全家，那地所有的人，都要在那里事奉我。在那里我悦纳他们，并要你们献供物和初熟的土产，以及一切的圣物。这是主耶和华说的。
EZEK|20|41|我把你们从万民中领出来，从被赶散到的列邦聚集你们，那时我必悦纳你们如同悦纳馨香之祭，我要在列国眼前，在你们中间显为圣。
EZEK|20|42|我领你们进入 以色列 地，就是我起誓应许赐给你们列祖之地，那时你们就知道我是耶和华。
EZEK|20|43|你们在那里要追念那玷污自己的所作所为，又要因所行的一切恶事厌恶自己。
EZEK|20|44|以色列 家啊，我为我名的缘故，没有照着你们的恶行和你们的败坏对待你们；你们就知道我是耶和华。这是主耶和华说的。”
EZEK|20|45|耶和华的话临到我，说：
EZEK|20|46|“人子啊，你要面向南方，向南方传讲 ，向 尼革夫 田野的树林说预言。
EZEK|20|47|你要对 尼革夫 的树林说，要听耶和华的话。主耶和华如此说：看哪，我要在你那里点火，烧灭你们中间所有的绿树和枯树，猛烈的火焰必不熄灭；从南到北，人的脸都被烧焦。
EZEK|20|48|凡血肉之躯都知道是我─耶和华点了火，这火必不熄灭。”
EZEK|20|49|于是我说：“唉！主耶和华啊，人都指着我说：他不是说比喻的人吗？”
EZEK|21|1|耶和华的话临到我，说：
EZEK|21|2|“人子啊，把你的脸正对着 耶路撒冷 ，对着圣所 传讲 ，向 以色列 地说预言。
EZEK|21|3|你要向 以色列 地说，耶和华如此说：看哪，我与你为敌，拔刀出鞘，把义人和恶人从你中间剪除。
EZEK|21|4|因为我要剪除你当中的义人和恶人，所以我的刀要出鞘，从南到北攻击所有的血肉之躯；
EZEK|21|5|凡血肉之躯都知道我─耶和华已拔刀出鞘，刀必不再入鞘。
EZEK|21|6|你，人子啊，要叹息，在他们眼前断了腰，愁苦地叹息。
EZEK|21|7|若有人对你说：‘你为什么叹息呢？’你就说：‘因为有风声传来，人心惶惶，双手发软，精神衰败，膝弱如水。看哪，它临近了，一定会发生。’这是主耶和华说的。”
EZEK|21|8|耶和华的话临到我，说：
EZEK|21|9|“人子啊，你要预言说，耶和华如此吩咐，你要说： 有刀，刀已磨快， 又擦亮了；
EZEK|21|10|磨快为要大大杀戮， 擦亮为要像闪电。 我们岂能快乐呢？ 它藐视我儿的权杖和一切的木头 。
EZEK|21|11|它已经交给人擦亮，可以掌握使用；这刀已经磨快擦亮，好交在行杀戮的人手中。
EZEK|21|12|人子啊，你要呼喊哀号，因为这刀将临到我的百姓，临到 以色列 所有的领袖身上。他们和我的百姓都要交在刀下，所以你要捶胸 。
EZEK|21|13|因为这是一个考验，若它藐视权杖，也不算一回事，又怎么样呢？这是主耶和华说的。”
EZEK|21|14|“人子啊，你要拍掌预言，使这刀三番两次临到；这是致人死伤的刀，就是包围人，使人大受死伤的刀。
EZEK|21|15|我设立这恐吓 的刀，攻击他们一切的城门，为要使他们的心惊慌害怕，许多人因而跌倒。唉！它 造得像闪电，磨得尖利 ，要行杀戮。
EZEK|21|16|刀啊，要行动一致 ，向右边，或指向左边；面向哪方，就向哪方。
EZEK|21|17|我也要拍掌，使我的愤怒平息。这是我─耶和华说的。”
EZEK|21|18|耶和华的话临到我，说：
EZEK|21|19|“人子啊，你要画定两条路线，使 巴比伦 王的刀过来，这两条路必从同一地分出来；要在通往城里的路口画手作指标。
EZEK|21|20|你要划定一条路，使刀来到 亚扪 人的 拉巴 ，来到 犹大 ，在坚固城 耶路撒冷 。
EZEK|21|21|因为 巴比伦 王站在岔路上，在两条路口占卜。他摇签 求问神像，察看肝脏；
EZEK|21|22|右手是 耶路撒冷 的占卜，以便安设撞城槌，张口喊杀 ，扬声呼叫，建土堆，筑堡垒，以撞城槌攻打城门。
EZEK|21|23|在那些曾郑重起誓的 犹大 人眼中，这是虚假的占卜；但 巴比伦 王要使他们想起自己的罪孽，以便俘掳他们。”
EZEK|21|24|于是，主耶和华如此说：“因你们的过犯显露，你们的罪孽被记得，以致你们的罪恶在你们一切的行为上都彰显出来；你们既被记得，就被掳在掌中。
EZEK|21|25|你这亵渎行恶的 以色列 王啊，你的日子，最后惩罚的时刻已来临。
EZEK|21|26|主耶和华如此说：当除掉荣冕，摘下华冠，景况已不复从前；要使卑者升为高，使高者降为卑。
EZEK|21|27|我要将这国倾覆，倾覆，再倾覆；这国必不存在，直等到那应得的人来到，我就将国赐给他。”
EZEK|21|28|“人子啊，你要说预言；你要说，论到 亚扪 人和他们的凌辱，主耶和华吩咐我如此说：有刀，拔出来的刀，已经擦亮，为了行杀戮；它亮如闪电以行吞灭。
EZEK|21|29|他们为你见虚假的异象，行谎诈的占卜，使你倒在亵渎之恶人的颈项上；他们的日子，最后惩罚的时刻已来临。
EZEK|21|30|你收刀入鞘吧！我要在你受造之处、生长之地惩罚你。
EZEK|21|31|我要把我的愤怒倾倒在你身上，把我烈怒的火喷在你身上；又将你交在善于杀灭、畜牲一般的人手中。
EZEK|21|32|你要成为火中之柴，你的血必在地里；你必不再被记得，因为这是我─耶和华说的。”
EZEK|22|1|耶和华的话临到我，说：
EZEK|22|2|“你，人子啊，你要审问，审问这流人血的城吗？要使它知道它一切可憎的事。
EZEK|22|3|你要说，主耶和华如此说：那在其中流人血的城啊，它的时刻已到，它制造偶像玷污了自己。
EZEK|22|4|你因流了人的血，算为有罪；因所制造的偶像，玷污自己；你使你的日子临近，你的年数已来到 。所以我使你承受列国的凌辱和列邦的讥诮。
EZEK|22|5|你这恶名昭彰、混乱的城啊，离你或远或近的国家都必讥诮你。
EZEK|22|6|“看哪， 以色列 的领袖在你那里，为了流人的血各逞其能。
EZEK|22|7|你那里有轻慢父母的，在你当中有欺压寄居者的，你那里也有亏负孤儿寡妇的。
EZEK|22|8|你藐视我的圣物，干犯我的安息日。
EZEK|22|9|你那里有为流人血而毁谤人的，你那里有在山上吃祭物的，在你当中也有行淫乱的，
EZEK|22|10|有露父亲下体的 ，有玷辱经期中不洁净之妇人的。
EZEK|22|11|这人与邻舍的妻子行可憎的事，那人行淫污辱媳妇，在你那里还有人污辱他的姊妹，父亲的女儿。
EZEK|22|12|你那里有收取报酬而流人血的。你取利息，又索取高利；欺压邻舍，夺取财物；你竟然忘了我。这是主耶和华说的。
EZEK|22|13|“看哪，我因你所得不义之财和你们中间所流的血，就击打手掌。
EZEK|22|14|到了我对付你的日子，你的心岂能忍受呢？你的手还能有力吗？我─耶和华说了这话，就必成就。
EZEK|22|15|我要把你驱散到列国，分散在列邦。我也必除掉你们中间的污秽。
EZEK|22|16|你在列国眼前因自己所做的被侮辱 ，你就知道我是耶和华。”
EZEK|22|17|耶和华的话临到我，说：
EZEK|22|18|“人子啊，我看 以色列 家为渣滓。他们是炉中的铜、锡、铁、铅，是炼银的渣滓 。
EZEK|22|19|所以主耶和华如此说：因你们全都成为渣滓，所以，看哪，我必将你们聚集在 耶路撒冷 中。
EZEK|22|20|人怎样把银、铜、铁、铅、锡聚在炉中，吹火使它镕化；照样，我也要在我的怒气和愤怒中聚集你们，把你们安置在城中，使你们镕化。
EZEK|22|21|我必聚集你们，把我烈怒的火吹在你们身上，你们就在其中镕化。
EZEK|22|22|银子怎样在炉中镕化，你们也必照样在城中镕化，因此就知道是我─耶和华把愤怒倾倒在你们身上。”
EZEK|22|23|耶和华的话临到我，说：
EZEK|22|24|“人子啊，你要向这地说：你是未被洁净 之地，在我盛怒的日子，没有雨水在其上。
EZEK|22|25|其中的先知同谋背叛 ，如咆哮的狮子抓撕掠物。他们吞灭人命，抢夺财宝，使这地寡妇增多。
EZEK|22|26|其中的祭司曲解我的律法，亵渎我的圣物，不分别圣与俗，也不使人分辨洁净和不洁净，又遮眼不顾我的安息日；在他们中间连我也被亵慢了。
EZEK|22|27|其中的领袖仿佛野狼抓撕掠物，流人的血，伤害人命，为得不义之财。
EZEK|22|28|其中的先知为他们粉刷，见虚假的异象，行谎诈的占卜，说：‘主耶和华如此说’，其实耶和华并没有说。
EZEK|22|29|这地的百姓惯行欺压抢夺之事，亏负困苦和贫穷的人，欺压寄居者，没有公平。
EZEK|22|30|我在他们中间寻找一人重修城墙，在我面前为这地站在缺口上，使我不致灭绝它，却连一个也找不着。
EZEK|22|31|所以我把愤怒倾倒在他们身上，用烈怒之火消灭他们，照他们所做的报应在他们头上。这是主耶和华说的。”
EZEK|23|1|耶和华的话临到我，说：
EZEK|23|2|“人子啊，有两个女子，是一母所生，
EZEK|23|3|她们在 埃及 行淫，年少时就开始行淫；在那里任人拥抱胸怀，抚弄她们少女的乳房。
EZEK|23|4|她们的名字，大的叫 阿荷拉 ，妹妹叫 阿荷利巴 。她们都归于我，生了儿女。论到她们的名字， 阿荷拉 是 撒玛利亚 ， 阿荷利巴 是 耶路撒冷 。
EZEK|23|5|“ 阿荷拉 归我之后却仍行淫，恋慕所爱的人，就是 亚述 人，都是战士 ，
EZEK|23|6|穿着蓝衣，作省长、副省长，全都是俊美的年轻人，骑着马的骑士。
EZEK|23|7|阿荷拉 与 亚述 人中所有的美男子放纵淫行，她因拜所恋慕之人的一切偶像，玷污了自己。
EZEK|23|8|她从 埃及 的时候，就没有离开过淫乱；因为她年轻时，有人与她同寝，抚弄她少女的乳房，和她纵欲行淫。
EZEK|23|9|因此，我把她交在她所爱的人手中，就是她所恋慕的 亚述 人手中。
EZEK|23|10|他们暴露她的下体，掳掠她的儿女，用刀杀了她；他们向她施行审判，使她在妇女中留下臭名。
EZEK|23|11|“她妹妹 阿荷利巴 虽然看见了，却还是纵欲，比姊姊更加腐败，行淫乱比姊姊更甚。
EZEK|23|12|她恋慕 亚述 人，就是省长和副省长，披挂整齐的战士，骑着马的骑士，全都是俊美的年轻人。
EZEK|23|13|我看见她被污辱，姊妹二人同行一路。
EZEK|23|14|阿荷利巴 又加增淫行，她看见墙上刻有人像，就是鲜红色的 迦勒底 人雕刻的像。
EZEK|23|15|它们腰间系着带子，头上有飘扬的裹头巾，都是将军的样子， 巴比伦 人的形像； 迦勒底 是他们的出生地。
EZEK|23|16|阿荷利巴 一看见就恋慕他们，派遣使者往 迦勒底 他们那里去。
EZEK|23|17|巴比伦 人来到她那里，上了她爱情的床，与她行淫污辱她。她被污辱，随后她的心却与他们生疏。
EZEK|23|18|这样，她既暴露淫行，暴露下体；我的心就与她生疏，像先前与她的姊姊生疏一样。
EZEK|23|19|她仍继续增添淫行，追念她年轻时在 埃及 地行淫的日子，
EZEK|23|20|恋慕情人的身壮精足，如驴似马。
EZEK|23|21|这样，你就渴望年轻时的淫荡；那时， 埃及 人因你年轻时的胸怀，抚弄你的乳房 。”
EZEK|23|22|阿荷利巴 啊，主耶和华如此说：“看哪，我要激起先前你喜爱，而后生疏的人前来攻击你。我必使他们前来，在你四围攻击你；
EZEK|23|23|有 巴比伦 人、 迦勒底 众人、 比割 人、 书亚 人、 哥亚 人，还有 亚述 众人与他们一起，都是俊美的年轻人。他们是省长、副省长、将军、有名声的，全都骑着马。
EZEK|23|24|他们用兵器、 战车、辎重车，率领大军前来攻击你。他们要拿大小盾牌，戴着头盔，在你四围摆阵攻击你。我要把审判交给他们，他们必按着自己的规条审判你。
EZEK|23|25|我要向你倾泄我的妒忌，使他们以愤怒对待你。他们必割去你的鼻子和耳朵，你剩余的人必倒在刀下。他们必掳去你的儿女，你所剩余的必被火焚烧。
EZEK|23|26|他们必剥去你的衣服，夺取你美丽的宝物。
EZEK|23|27|这样，我必止息你的淫行和你从 埃及 地就开始犯的淫乱，使你不再仰望 亚述 ，也不再追念 埃及 。
EZEK|23|28|主耶和华如此说：看哪，我必把你交在你所恨恶的人手中，就是你心与他生疏的人手中。
EZEK|23|29|他们要以恨恶对待你，夺取你劳碌得来的一切，留下你赤身露体。你淫乱的下体，连你的淫行和淫荡，都必显露。
EZEK|23|30|人必向你行这些事；因为你随从外邦人行淫，用他们的偶像玷污自己。
EZEK|23|31|你走了你姊姊的路，所以我必把她的杯交在你的手中。”
EZEK|23|32|主耶和华如此说： “你必喝你姊姊的杯， 那杯又深又广， 盛得很多， 使你遭受嗤笑讥刺。
EZEK|23|33|你必酩酊大醉， 满有愁苦。 你姊姊 撒玛利亚 的杯， 惊骇和凄凉的杯，
EZEK|23|34|你必喝它，并且喝干。 甚至咀嚼杯片， 撕裂自己的胸脯； 因为我曾说过。 这是主耶和华说的。”
EZEK|23|35|主耶和华如此说：“因你忘记我，将我丢在背后，所以你要担当你的淫行和淫荡。”
EZEK|23|36|耶和华对我说：“人子啊，你要审问 阿荷拉 与 阿荷利巴 吗？要指出她们所做可憎的事。
EZEK|23|37|她们行奸淫，手中有血。她们与偶像行奸淫，使她们为我所生的儿女经火，给它们当食物。
EZEK|23|38|此外，她们还向我这样做：同一天又玷污我的圣所，干犯我的安息日。
EZEK|23|39|她们杀了儿女献给偶像，当天又进入我的圣所，亵渎了它。看哪，这就是她们在我殿中所做的。
EZEK|23|40|“况且你们两姊妹派人从远方召人来。使者到了他们那里，看哪，他们就来了。为了他们，你们沐浴，画眼影，佩戴首饰，
EZEK|23|41|坐在华美的床上，前面摆设桌子，把我的香料和膏油放在其上。
EZEK|23|42|在那里有一群人欢乐的声音；有许多的平民，从旷野来的醉汉 ，把镯子戴在她们手上，把华冠戴在她们头上。
EZEK|23|43|“我论到这久行奸淫而色衰的妇人说：现在人们还要与她行淫，她也要与人行淫。
EZEK|23|44|人去到 阿荷拉 和 阿荷利巴 二淫妇那里 ，好像与妓女行淫。
EZEK|23|45|义人必按照审判淫妇和流人血之妇人的规条，审判她们；因为她们是淫妇，她们的手中有血。”
EZEK|23|46|主耶和华如此说：“我要让军队上来攻击她们，使她们惊骇，成为掳物。
EZEK|23|47|这军队必用石头打死她们，用刀剑杀害她们，又杀戮她们的儿女，用火焚烧她们的房屋。
EZEK|23|48|我必使这地不再有淫行，所有的妇女都受警戒，不再效法你们的淫行 。
EZEK|23|49|人必因你们的淫行报应你们；你们要担当拜偶像的罪，因此你们就知道我是主耶和华。”
EZEK|24|1|第九年十月初十，耶和华的话临到我，说：
EZEK|24|2|“人子啊，你要记录这一天的名称，这特别的一天， 巴比伦 王围困 耶路撒冷 ，就在这特别的一天。
EZEK|24|3|你要向这悖逆之家设比喻，对他们说，主耶和华如此说： 把锅放在火上， 放好了，倒水在其中；
EZEK|24|4|要将肉块，一切肥美的肉块， 腿和肩都放在锅里， 要装满上等的骨头；
EZEK|24|5|要取羊群中最好的， 把柴 堆在下面， 把它煮开， 骨头煮在其中。
EZEK|24|6|“主耶和华如此说：祸哉！这流人血的城，就是长锈的锅。它的锈未曾除掉，要将肉块从其中一一取出，不必抽签。
EZEK|24|7|这城所流的血还在城中，血倒在光滑的磐石上，没有倒在地上，用土掩盖；
EZEK|24|8|是我使这城所流的血倒在光滑的磐石上，不得掩盖，为要惹动愤怒，施行报应。
EZEK|24|9|所以主耶和华如此说：祸哉！这流人血的城，我必亲自加大柴堆。
EZEK|24|10|你要添上木柴，使火着旺，将肉煮烂，加上香料 ，烤焦骨头；
EZEK|24|11|你要把空锅放在炭火上，将锅烧热，把铜烧红，镕化其中的污秽，除净其上的锈。
EZEK|24|12|然而这一切劳碌无效 ，它厚厚的锈，即使用火也除不掉。
EZEK|24|13|虽然我想洁净你污秽的淫行，你却不洁净，你的污秽再也不能洁净，直等我止息了向你发的愤怒。
EZEK|24|14|我─耶和华说了这话，时候到了，就必成就；必不退缩，不顾惜，也不怜悯。人必照你的所作所为审判你。这是主耶和华说的。”
EZEK|24|15|耶和华的话临到我，说：
EZEK|24|16|“人子，看哪，我要以灾病夺取你眼中所喜爱的，你却不可悲哀哭泣，也不可流泪，
EZEK|24|17|只可叹息，不可出声，不可办理丧事；裹上头巾，脚上穿鞋，不可捂着胡须，也不可吃一般人的食物 。”
EZEK|24|18|到了早晨我把这事告诉百姓，晚上我的妻子就死了。次日早晨我就遵命而行。
EZEK|24|19|百姓对我说：“你这样做跟我们有什么关系，你不告诉我们吗？”
EZEK|24|20|我对他们说：“耶和华的话临到我，说：
EZEK|24|21|‘你告诉 以色列 家，主耶和华如此说：我要使我的圣所被亵渎，就是你们凭势力所夸耀、眼里所喜爱、心中所爱惜的；并且你们所遗留的儿女必倒在刀下。
EZEK|24|22|那时，你们要照我所做的去做。你们不可捂着胡须，也不可吃一般人的食物。
EZEK|24|23|你们头要裹上头巾，脚要穿上鞋；不可悲哀哭泣。你们必因自己的罪孽衰残，相对叹息。
EZEK|24|24|以西结 必这样成为你们的预兆；凡他所做的，你们也必照样做。那事来到，你们就知道我是主耶和华。’”
EZEK|24|25|“你，人子啊，那日当我除掉他们所倚靠的保障、所欢喜的荣耀，并眼中所喜爱的，心里所重看的儿女时，
EZEK|24|26|逃脱的人岂不来到你这里，使你耳闻这事吗？
EZEK|24|27|那日你要向逃脱的人开口说话，不再哑口无言。你必这样成为他们的预兆，他们就知道我是耶和华。”
EZEK|25|1|耶和华的话临到我，说：
EZEK|25|2|“人子啊，你要面向 亚扪 人说预言，攻击他们。
EZEK|25|3|你要对 亚扪 人说，当听主耶和华的话。主耶和华如此说：我的圣所遭亵渎， 以色列 地变荒凉， 犹大 家被掳掠；那时，你因这些事说‘啊哈’，
EZEK|25|4|所以，看哪，我要把你交给东方人为业；他们必在你中间安营居住，设立居所，吃你的果子，喝你的奶。
EZEK|25|5|我必使 拉巴 成为牧放骆驼之地，使 亚扪 成为羊群躺卧之处，你们就知道我是耶和华。
EZEK|25|6|主耶和华如此说：因你们拍手顿足，幸灾乐祸，藐视 以色列 地，
EZEK|25|7|所以，看哪，我要伸手攻击你，把你交给列国作为掳物。我必从万民中剪除你，从列邦中消灭你。我必除灭你，你就知道我是耶和华。”
EZEK|25|8|“主耶和华如此说：因 摩押 和 西珥 人说‘看哪， 犹大 家与列国无异’，
EZEK|25|9|所以，看哪，我要破开 摩押 边界的城镇，就是 摩押 人所夸耀的城镇， 伯．耶施末 、 巴力．免 、 基列亭 ，
EZEK|25|10|令东方人前来攻击 亚扪 人。我必将 亚扪 交给他们为业，使 亚扪 人在列国中不再被记念。
EZEK|25|11|我也必向 摩押 施行审判，他们就知道我是耶和华。”
EZEK|25|12|“主耶和华如此说：因为 以东 向 犹大 家报仇，因向他们报仇而大大显为有罪，
EZEK|25|13|所以主耶和华如此说：我要伸手攻击 以东 ，将人与牲畜剪除，使 以东 从 提幔 起，直到 底但 ，地变荒凉，人也都倒在刀下。
EZEK|25|14|我要藉我子民 以色列 的手报复 以东 ；他们必照我的怒气，按我的愤怒对待 以东 ， 以东 人就知道施报的是我。这是主耶和华说的。”
EZEK|25|15|“主耶和华如此说：因 非利士 人报仇，就是心存轻蔑报仇；他们永怀仇恨，意图毁灭，
EZEK|25|16|所以主耶和华如此说：看哪，我要伸手攻击 非利士 人，剪除 基利提 人，灭绝沿海剩余的居民。
EZEK|25|17|我要大大报复他们，发怒斥责他们。我报复他们的时候，他们就知道我是耶和华。”
EZEK|26|1|第十一年某月初一，耶和华的话临到我，说：
EZEK|26|2|“人子啊，因 推罗 向 耶路撒冷 说：‘啊哈！那众民之门已经破坏，向我敞开；它既变为废墟，我必丰盛。’
EZEK|26|3|所以，主耶和华如此说： 推罗 ，看哪，我与你为敌，使许多国家涌上攻击你，如同海洋使波浪涌上一样。
EZEK|26|4|他们要破坏 推罗 的城墙，拆毁它的城楼。我也要刮净它的尘土，使它成为光滑的磐石。
EZEK|26|5|推罗 必成为海中的晒网场，因为我曾说过， 这是主耶和华说的。它必成为列国的掳物，
EZEK|26|6|推罗 乡间邻近的城镇 必遭刀剑灭绝，他们就知道我是耶和华。”
EZEK|26|7|主耶和华如此说：“看哪，我必使诸王之王，就是 巴比伦 王 尼布甲尼撒 ，率领马匹、战车、骑兵、军队和许多人从北方来攻击 推罗 。
EZEK|26|8|他必用刀剑杀灭你乡间邻近的城镇，也必筑堡垒，建土堆，举盾牌攻击你。
EZEK|26|9|他要安设撞城槌攻破你的城墙，以刀剑拆毁你的城楼。
EZEK|26|10|因他马匹众多，尘土必扬起遮蔽你。他进入你的城门，如同进入已有缺口之城。那时，你的城墙必因骑兵、车轮和战车的响声震动。
EZEK|26|11|他的马蹄必践踏你所有的街道；他必用刀剑杀戮你的居民。你坚固的柱子 必倒在地上。
EZEK|26|12|人必掳获你的财宝，掠夺你的货财；他们要破坏你的城墙，拆毁你华美的房屋，将你的石头、木头、尘土都抛在水中。
EZEK|26|13|我要使你唱歌的声音止息；人不再听见你弹琴的声音。
EZEK|26|14|我必使你成为光滑的磐石，作晒网的场所。你不得再被建造，因为我─耶和华已这样说了。这是主耶和华说的。”
EZEK|26|15|主耶和华对 推罗 如此说：“在你中间行杀戮，受伤的人唉哼时，海岛岂不都因你倾倒的响声震动吗？
EZEK|26|16|那时沿海的君王都要从宝座下来，除去朝服，脱下锦衣，披上战兢，坐在地上，不停发抖，为你而惊骇。
EZEK|26|17|他们必为你作哀歌，向你说： ‘你这闻名之城， 航海之人居住， 海上最为坚固的， 你和居民使所有住在沿海的人 无不惊恐， 现在竟然毁灭了！
EZEK|26|18|如今在你倾覆的日子， 海岛都要战兢； 海中的群岛见你归于无有 就都惊惶。’”
EZEK|26|19|主耶和华如此说：“ 推罗 啊 ，我要使你变为荒凉，如无人居住的城镇；又使深水漫过你，大水淹没你。
EZEK|26|20|那时，我要使你和下到地府的人同去，到古时候的人那里；我要使你和下到地府的人一同住在地的深处，在久已荒废的地方，使你那里不再有人居住；我要在活人之地显荣耀 。
EZEK|26|21|我必叫你令人惊恐，使你不再存留于世；人虽寻找你，却永不寻见。这是主耶和华说的。”
EZEK|27|1|耶和华的话临到我，说：
EZEK|27|2|“人子啊，要为 推罗 作哀歌。
EZEK|27|3|你要对位于海口，跟许多海岛的百姓做生意的 推罗 说，主耶和华如此说： 推罗 啊，你曾说： ‘我全然美丽。’
EZEK|27|4|你的疆界在海的中心， 造你的使你全然美丽。
EZEK|27|5|他们用 示尼珥 的松树作你的甲板， 用 黎巴嫩 的香柏树作桅杆，
EZEK|27|6|用 巴珊 的橡树作你的桨， 用镶嵌象牙的 基提 海岛黄杨木 为舱板。
EZEK|27|7|你的帆是用 埃及 绣花细麻布做的， 可作你的大旗； 你的篷是用 以利沙岛 的蓝色和紫色布做的。
EZEK|27|8|西顿 和 亚发 的居民为你划桨； 推罗 啊，你们中间的智慧人为你掌舵。
EZEK|27|9|迦巴勒 的长者和智者 在你中间修补裂缝； 海上一切的船只和水手 都在你那里进行货物交易。
EZEK|27|10|“ 波斯 人、 路德 人、 弗 人在你的军营中作战士；他们在你们中间悬挂盾牌和头盔，彰显你的尊荣。
EZEK|27|11|亚发 人和你的军队都驻守在四围的城墙上，你的城楼上也有勇士；他们悬挂盾牌，成全你的美丽。
EZEK|27|12|“ 他施 因你多有财物，就作你的客商，他们带着银、铁、锡、铅前来换你的商品。
EZEK|27|13|雅完 、 土巴 、 米设 都与你交易，以人口和铜器换你的货物。
EZEK|27|14|陀迦玛 族用马匹、战马和骡子换你的商品。
EZEK|27|15|底但 人与你交易，许多海岛成为你的码头；他们拿象牙、黑檀木与你交换。
EZEK|27|16|亚兰 因你货品充裕，就作你的客商；他们用绿宝石、紫色布、刺绣、细麻布、珊瑚、红宝石换你的商品。
EZEK|27|17|犹大 和 以色列 地都与你交易；他们用 米匿 的小麦、饼、蜜、油、乳香换你的货物。
EZEK|27|18|大马士革 也因你货品充裕，多有各类财物，就带来 黑本 酒和白羊毛与你交易。
EZEK|27|19|威但 和从 乌萨 来的 雅完 人 为了你的货物，以加工的铁、桂皮、香菖蒲换你的商品。
EZEK|27|20|底但 以骑马用的座垫毯子与你交换。
EZEK|27|21|阿拉伯 和 基达 所有的领袖都作你的客商，用羔羊、公绵羊、公山羊与你交换。
EZEK|27|22|示巴 和 拉玛 的商人也来与你交易，他们用各类上好的香料、各类的宝石和黄金换你的商品。
EZEK|27|23|哈兰 、 干尼 、 伊甸 、 示巴 商人、 亚述 和 基抹 都与你交易。
EZEK|27|24|这些商人将美好的货物包在蓝色的绣花包袱内，又将华丽的衣服装在香柏木的箱子里，用绳索捆着，以此与你交易 。
EZEK|27|25|他施 的船只为你运货， 你在海中满载货物，极其沉重。
EZEK|27|26|划桨的把你划到水深之处， 东风在海中将你击破。
EZEK|27|27|你的财宝、商品、货物、 水手、掌舵的、 修补船缝的、进行货物交易的， 并你那里所有的战士 和你中间所有的军队， 在你倾覆的日子都必沉在海底。
EZEK|27|28|因掌舵者的呼声， 郊野就必震动。
EZEK|27|29|所有划桨的 都从他们的船下来； 水手和所有在海上掌舵的， 都要登岸。
EZEK|27|30|他们必为你放声痛哭， 撒尘土于头上， 在灰中打滚；
EZEK|27|31|又为你使头光秃， 用麻布束腰， 号啕痛哭， 痛苦至极。
EZEK|27|32|他们哀号的时候， 为你作哀歌， 为你痛哭： 有何城如 推罗 ， 在海中沉寂呢？
EZEK|27|33|你由海上运出商品， 使许多民族充裕； 你以许多财宝货物 令地上的君王丰富。
EZEK|27|34|在深水中被海浪打破的时候， 你的货物和你中间所有的军队都下沉。
EZEK|27|35|海岛所有的居民为你惊奇， 他们的君王都甚恐慌，面带愁容。
EZEK|27|36|万民中的商人向你发嘘声； 你令人惊恐， 不再存留于世，直到永远。”
EZEK|28|1|耶和华的话临到我，说：
EZEK|28|2|“人子啊，你要对 推罗 的君王说，主耶和华如此说： 你心里高傲，说：‘我是神明； 我在海中坐诸神之位。’ 虽然你把你的心比作神明的心， 你却不过是人，并不是神明！
EZEK|28|3|看哪，你比 但以理 更有智慧， 任何秘密都不能向你隐藏。
EZEK|28|4|你靠自己的智慧聪明得了财宝， 把金银收入库房；
EZEK|28|5|你靠自己的大智慧以贸易增添财宝， 又因你的财宝心里高傲；
EZEK|28|6|所以主耶和华如此说： 因你把你的心比作神明的心，
EZEK|28|7|所以，看哪，我必使外国人， 就是列国中凶暴的人临到你这里； 他们要拔刀摧毁你用智慧得来的美物， 污损你的荣光。
EZEK|28|8|他们必使你坠入地府； 你要像被刺杀之人的死，死在海中。
EZEK|28|9|在杀你的人面前， 你还能说‘我是神明’吗？ 在杀害你的人手中， 你不过是人，并不是神明。
EZEK|28|10|你要死在陌生人手中， 像未受割礼之人的死， 因为我曾说过， 这是主耶和华说的。”
EZEK|28|11|耶和华的话临到我，说：
EZEK|28|12|“人子啊，要为 推罗 王作哀歌，对他说，主耶和华如此说： 你曾是完美的典范， 智慧充足，全然美丽。
EZEK|28|13|你在 伊甸 ─上帝的园中， 佩戴各样宝石， 就是红宝石、红璧玺、金刚石、 水苍玉、红玛瑙、碧玉、 蓝宝石、绿宝石、红玉； 你的宝石有黄金的底座，手工精巧 ， 都是在你受造之日预备的。
EZEK|28|14|我指定你为受膏的基路伯， 看守保护； 你在上帝的圣山上； 往来在如火的宝石中。
EZEK|28|15|你从受造之日起行为正直， 直到后来查出你的不义。
EZEK|28|16|你因贸易发达， 暴力充斥其中，以致犯罪， 所以我污辱你，使你离开上帝的山。 守护者基路伯啊， 我已将你从如火的宝石中歼灭。
EZEK|28|17|你因美丽心中高傲， 因荣光而败坏智慧， 我已将你抛弃在地， 把你摆在君王面前， 好叫他们目睹眼见。
EZEK|28|18|你因罪孽众多，贸易不公， 亵渎了你的圣所； 因此我使火从你中间发出， 烧灭了你， 使你在所有观看的人眼前 变为地上的灰烬。
EZEK|28|19|万民中凡认识你的 都必为你惊奇。 你令人惊恐， 不再存留于世，直到永远。”
EZEK|28|20|耶和华的话临到我，说：
EZEK|28|21|“人子啊，你要面向 西顿 ，向它说预言。
EZEK|28|22|你要说，主耶和华如此说： ‘ 西顿 ，看哪，我与你为敌， 我要在你中间得荣耀。’ 我在它中间施行审判、显为圣的时候， 人就知道我是耶和华。
EZEK|28|23|我必令瘟疫进入 西顿 ， 使血流在街上。 刀剑从四围临到它， 被杀的要仆倒在其中； 人就知道我是耶和华。”
EZEK|28|24|“四围恨恶 以色列 家的人，对他们必不再如刺人的荆棘、伤人的蒺藜；他们就知道我是主耶和华。”
EZEK|28|25|主耶和华如此说：“我将分散在万民中的 以色列 家召集回来，在列国眼前向他们显为圣的时候，他们仍可在我所赐给我仆人 雅各 之地居住。
EZEK|28|26|他们要在这地上安然居住。我向四围恨恶他们的众人施行审判之后，他们要建造房屋，栽葡萄园，安然居住，他们就知道我是耶和华─他们的上帝。”
EZEK|29|1|第十年十月十二日，耶和华的话临到我，说：
EZEK|29|2|“人子啊，你要面向 埃及 王法老，向他和 埃及 全地说预言。
EZEK|29|3|你要说，主耶和华如此说： 埃及 王法老， 你这卧在自己江河中的海怪， 看哪，我与你为敌。 你曾说：‘我的 尼罗河 是我的， 是我为自己造的。’
EZEK|29|4|我必用钩子钩住你的腮颊， 令江河中的鱼贴住你的鳞甲； 我要把你和所有贴着鳞甲的鱼 从你的江河中拉上来。
EZEK|29|5|我要把你和江河中的鱼全都抛弃在旷野； 你必仆倒在田间， 无人收殓，无人掩埋。 我已将你给了地上的走兽、空中的飞鸟作食物。
EZEK|29|6|“ 埃及 所有的居民必定知道我是耶和华。因为你已成为 以色列 家芦苇的杖；
EZEK|29|7|他们用手掌一握，你就断裂，伤了他们的肩；他们靠着你，你却折断，闪了他们的腰 。
EZEK|29|8|所以主耶和华如此说：我必使刀剑临到你，把人与牲畜从你中间剪除。
EZEK|29|9|埃及 地必荒芜废弃，他们就知道我是耶和华。 “因为法老说‘ 尼罗河 是我的，是我所造的’，
EZEK|29|10|所以，看哪，我必与你和你的江河为敌，使 埃及 地，从 密夺 到 色弗尼 ，直到 古实 边界，全然废弃荒芜。
EZEK|29|11|人的脚不经过，兽的蹄也不经过，四十年之久无人居住。
EZEK|29|12|我要使 埃及 地成为荒芜中最荒芜的地，使它的城镇变为荒废中最荒废的城镇，共四十年之久。我必将 埃及 人分散到列国，四散在列邦。
EZEK|29|13|“主耶和华如此说：满了四十年后，我必招聚分散在万民中的 埃及 人。
EZEK|29|14|我要令 埃及 被掳的人归回，使他们回到本地 巴特罗 。在那里，他们必成为弱小的国家，
EZEK|29|15|成为列国中最低微的，不再自高于列邦之上。我必使他们变为小国，不再辖制列邦。
EZEK|29|16|埃及 必不再作 以色列 家的倚靠，却使 以色列 家想起他们仰赖 埃及 的罪。他们就知道我是主耶和华。”
EZEK|29|17|第二十七年正月初一，耶和华的话临到我，说：
EZEK|29|18|“人子啊， 巴比伦 王 尼布甲尼撒 令他的军兵大力攻打 推罗 ，以致头都光秃，肩都磨破；然而他和军兵虽然为攻打 推罗 花这么多力气，却没有从那里得到什么犒赏。
EZEK|29|19|所以主耶和华如此说：我要将 埃及 地赐给 巴比伦 王 尼布甲尼撒 ；他必掳掠 埃及 的财富，抢夺它的掳物，掳掠它的掠物，用以犒赏他的军兵。
EZEK|29|20|我将 埃及 地赐给他，犒赏他，因他们为我效劳。这是主耶和华说的。
EZEK|29|21|“当那日，我必使 以色列 家壮大 ，又必使你─ 以西结 在他们中间开口；他们就知道我是耶和华。”
EZEK|30|1|耶和华的话临到我，说：
EZEK|30|2|“人子啊，你要说预言；你要说，主耶和华如此说： 哀哉这日！你们应当哭号，
EZEK|30|3|因为日子近了， 耶和华的日子临近了； 那是密云之日， 是列国受罚 之期。
EZEK|30|4|必有刀剑临到 埃及 ； 被杀的人仆倒在 埃及 时， 古实 人颤惊不已。 埃及 的财富遭掳掠， 根基被拆毁。
EZEK|30|5|古实 人、 弗 人、 路德 人、混居的各族和 古伯 人，以及盟国的人都要与 埃及 人一同倒在刀下。”
EZEK|30|6|耶和华如此说： 扶助 埃及 的必倾倒， 埃及 骄傲的权势必降为卑， 从 密夺 到 色弗尼 ，人必倒在刀下。 这是主耶和华说的。
EZEK|30|7|埃及 成为荒凉中最荒凉的国， 它的城镇变为荒废中最荒废的城镇。
EZEK|30|8|我在 埃及 放火， 帮助 埃及 的，都遭灭绝； 那时，他们就知道我是耶和华。
EZEK|30|9|“到那日，必有使者从我面前乘船出去，使安逸无虑的 古实 人惊惧；当 埃及 遭难的日子，痛苦也必临到他们。看哪，这事临近了！
EZEK|30|10|主耶和华如此说： 我要藉 巴比伦 王 尼布甲尼撒 的手 除灭 埃及 的军队。
EZEK|30|11|他和随从他的人， 就是列国中凶暴的人， 要前来毁灭这地， 拔刀攻击 埃及 ， 使遍地布满被杀的人。
EZEK|30|12|我要使江河干涸， 将这地卖在恶人手中； 我要藉外国人的手， 使这地和其中所充满的变为荒芜； 这是我─耶和华说的。
EZEK|30|13|“主耶和华如此说： 我要毁灭偶像， 从 挪弗 除掉神像； 不再有君王出自 埃及 地， 我要使 埃及 地的人惧怕。
EZEK|30|14|我必令 巴特罗 荒凉， 在 琐安 放火， 向 挪 施行审判。
EZEK|30|15|我要将我的愤怒倾倒在 训 ， 埃及 的堡垒上， 要剪除 挪 的众民。
EZEK|30|16|我必在 埃及 放火， 训 必大大痛苦， 挪 被攻破， 挪弗 终日遭敌侵袭。
EZEK|30|17|亚文 和 比．伯实 的年轻人必倒在刀下， 这些城镇将被掳掠。
EZEK|30|18|我在 答比匿 折断 埃及 的轭 ， 使它骄傲的权势止息。 那时，日光必退去； 至于这城，必有密云遮蔽， 邻近的城镇 也遭掳掠。
EZEK|30|19|我要如此向 埃及 施行审判， 他们就知道我是耶和华。”
EZEK|30|20|第十一年正月初七，耶和华的话临到我，说：
EZEK|30|21|“人子啊，我已折断 埃及 王法老的一只膀臂；看哪，无人为他敷药，也无人为他包扎绷带，使他有力持刀。
EZEK|30|22|因此，主耶和华如此说：看哪，我与 埃及 王法老为敌，要折断他的膀臂，折断强壮的和已受伤的，使刀从他手中掉落。
EZEK|30|23|我必将 埃及 人分散到列国，四散在列邦。
EZEK|30|24|我要使 巴比伦 王的膀臂有力，把我的刀交在他手中；却要折断法老的膀臂，使他在 巴比伦 王面前呻吟，如同被杀的人一样。
EZEK|30|25|我要使 巴比伦 王的膀臂强壮，法老的膀臂却要下垂；当我把我的刀交在 巴比伦 王手中时，他要举刀攻击 埃及 地，他们就知道我是耶和华。
EZEK|30|26|我必将 埃及 人分散到列国，四散在列邦；他们就知道我是耶和华。”
EZEK|31|1|第十一年三月初一，耶和华的话临到我，说：
EZEK|31|2|“人子啊，你要对 埃及 王法老和他的军队说： 论到你的强盛，谁能与你相比呢？
EZEK|31|3|看哪， 亚述 是 黎巴嫩 的香柏树， 枝条荣美，荫密如林， 极其高大，树顶高耸入云。
EZEK|31|4|众水使它生长， 深水使它长高； 所栽之地有江河环绕， 汊出的水道流至田野的树木。
EZEK|31|5|所以它高大超过田野的树木； 生长时因水源丰沛， 枝子繁多，枝条增长。
EZEK|31|6|空中所有的飞鸟在枝子上搭窝， 野地所有的走兽在枝条下生子， 所有的大国也在它的荫下居住。
EZEK|31|7|它树大枝长，极为荣美， 因它的根在众水之旁。
EZEK|31|8|上帝园中的香柏树不能遮蔽它； 松树不及它的枝子， 枫树不及它的枝条， 上帝园中的树都没有它荣美。
EZEK|31|9|我使它枝条繁多， 极为荣美； 在上帝的园中， 伊甸 所有的树都嫉妒它。”
EZEK|31|10|所以主耶和华如此说：“因它 高大，树顶高耸入云，心高气傲，
EZEK|31|11|我要把它交给 列国中强人的手里，他们必定按它的罪恶惩治它。我已经驱逐它。
EZEK|31|12|外国人，就是列国中凶暴的人，已把它砍断抛弃。它的枝条掉落山间和一切谷中，枝子折断，落在地上一切河道。地上的万民都离开它的遮荫，抛弃了它。
EZEK|31|13|空中的飞鸟都栖身在掉落的树干上，野地的走兽也都躺卧在它的枝条中。
EZEK|31|14|为了要使水边的树木枝干不再长高，树顶也不再高耸入云；那些得水滋润的，不再屹立于其中。因为它们和下到地府的人一起，都被交与死亡，到了地底下。”
EZEK|31|15|主耶和华如此说：“它坠落阴间的那日，我为它遮盖深渊，拦住江河，使众水停流，以表哀悼。我使 黎巴嫩 为它悲哀，田野的树木都因它枯萎。
EZEK|31|16|我把它扔到阴间，与下到地府的人一同坠落。那时，列国听见坠落的响声就震惊； 伊甸 一切的树木，就是 黎巴嫩 中得水滋润、最佳最美的树，在地底下都得了安慰。
EZEK|31|17|这些树也要与它同下阴间，到被刀所杀的人那里；它们曾作它的膀臂 ，在列国中曾居住在它的荫下。
EZEK|31|18|在这样的荣耀与威势中， 伊甸 树木有谁能与你相比呢？然而你要与 伊甸 的树木一同到地底下；在未受割礼的人中，与被刀所杀的人一同躺下。 “法老和他的军队正是如此。这是主耶和华说的。”
EZEK|32|1|第十二年十二月初一，耶和华的话临到我，说：
EZEK|32|2|“人子啊，你要为 埃及 王法老作哀歌，说： 你在列国中，如同少壮狮子， 却像海里的海怪， 冲出江河， 以爪搅动诸水， 使江河浑浊。
EZEK|32|3|主耶和华如此说： 许多民族聚集时， 我要将我的网撒在你身上， 他们要把你拉上来。
EZEK|32|4|我要把你丢在地上， 抛在田野， 使空中的飞鸟落在你身上， 遍地的野兽因你得以饱足。
EZEK|32|5|我要将你的肉丢在山间， 用你巨大的尸首 填满山谷。
EZEK|32|6|我要以你所流的血 浸透大地， 漫过山顶， 溢满河道。
EZEK|32|7|我毁灭你时， 要遮蔽诸天， 使众星昏暗； 我必以密云遮掩太阳， 月亮也不放光。
EZEK|32|8|我要使天上发亮的光体 在你上面变为昏暗， 使你的地也变为黑暗。 这是主耶和华说的。
EZEK|32|9|“我使你在列国，在你所不认识的列邦中灭亡 。那时，我必使许多民族的心因你愁烦。
EZEK|32|10|当我在他们面前举起我的刀，我要使许多民族因你惊恐，他们的君王也必因你极其恐慌。在你仆倒的日子，他们各人为自己的性命时时战兢。
EZEK|32|11|主耶和华如此说： 巴比伦 王的刀必临到你。
EZEK|32|12|我必藉勇士的刀使你的军队仆倒；这些勇士都是列国中凶暴的人。 他们必使 埃及 的骄傲归于无有， 埃及 的军队必被灭绝。
EZEK|32|13|我要除灭众水旁一切的走兽， 人的脚必不再搅浑这水， 兽的蹄也不搅浑这水。
EZEK|32|14|那时，我必使他们的水澄清， 使他们的江河像油缓流。 这是主耶和华说的。
EZEK|32|15|我使 埃及 地荒废， 使这地空无一物， 又击杀其中所有的居民； 那时，他们就知道我是耶和华。
EZEK|32|16|“这是一首为人所吟唱的哀歌；列国的女子要唱这哀歌，她们要为 埃及 和它的军队唱这哀歌。这是主耶和华说的。”
EZEK|32|17|第十二年某月 十五日，耶和华的话临到我，说：
EZEK|32|18|“人子啊，你要为 埃及 的军队哀号，把他们和强盛之国 一同扔到地底下，与那些下到地府的人在一起。
EZEK|32|19|‘你的美丽胜过谁呢？ 坠落吧，与未受割礼的人躺在一起！’
EZEK|32|20|他们要仆倒在被刀所杀的人当中。 埃及 被交给刀剑，人要把它和它的军队拉走。
EZEK|32|21|强壮的勇士要在阴间对 埃及 王和他的盟友说话；他们未受割礼，被刀剑所杀，已经坠落躺下。
EZEK|32|22|“ 亚述 和它的全军在那里，四围都是坟墓；他们全都是被杀倒在刀下的人。
EZEK|32|23|他们的坟墓在地府极深之处，它的众军环绕它的坟墓，他们全都是被杀倒在刀下的人，曾在活人之地使人惊恐。
EZEK|32|24|“ 以拦 在那里，它的全军环绕它的坟墓；他们全都是被杀倒在刀下、未受割礼而到地底下的，曾在活人之地使人惊恐；他们与下到地府的人一同担当羞辱。
EZEK|32|25|人为它和它的军队在被杀的人中设立床榻，四围都是坟墓；他们都是未受割礼被刀所杀的，曾在活人之地使人惊恐；他们与下到地府的人一同担当羞辱。 以拦 已列在被杀的人中。
EZEK|32|26|“ 米设 、 土巴 和他们的全军都在那里，四围都是坟墓；他们都是未受割礼被刀所杀的，曾在活人之地使人惊恐。
EZEK|32|27|他们不得与那未受割礼 仆倒的勇士躺在一起；这些勇士带着兵器下到阴间，头枕着刀剑，骨头带着本身的罪孽，曾在活人之地使人惊恐。
EZEK|32|28|法老啊，你必与未受割礼的人一起毁灭，与被刀所杀的人躺在一起。
EZEK|32|29|“ 以东 在那里，它的君王和所有官长虽然英勇，还是与被刀所杀的人同列；他们必与未受割礼的和下到地府的人躺在一起。
EZEK|32|30|“在那里有北方的众王子和所有的 西顿 人，全都与被杀的人一同下去。他们虽然英勇，使人惊恐，还是蒙羞。他们未受割礼，和被刀所杀的人躺在一起，与下到地府的人一同担当羞辱。
EZEK|32|31|“法老看见他们，就为他的军兵，就是被刀所杀属法老的人和他的全军感到安慰。这是主耶和华说的。
EZEK|32|32|我任凭法老在活人之地使人惊恐，法老和他的军兵必躺在未受割礼和被刀所杀的人中。这是主耶和华说的。”
EZEK|33|1|耶和华的话临到我，说：
EZEK|33|2|“人子啊，你要吩咐本国的百姓，对他们说：我使刀剑临到哪一国，哪一国的百姓从他们中间选立一人，作为守望者。
EZEK|33|3|守望者见刀剑临到那地，若吹角警戒百姓，
EZEK|33|4|有人听见角声却不受警戒，刀剑来除灭了他，这人的血必归到自己头上。
EZEK|33|5|他听见角声，不受警戒，他的血必归到自己身上；他若受警戒，就救了自己的命。
EZEK|33|6|倘若守望者见刀剑临到，却不吹角，以致百姓未受警戒，刀剑来杀了他们中间的一个人，这人虽然因自己的罪孽而死，我却要从守望者的手里讨他的血债。
EZEK|33|7|“人子啊，我照样立你作 以色列 家的守望者；你要听我口中的话，替我警戒他们。
EZEK|33|8|我对恶人说：‘恶人哪，你必要死！’你若不开口警戒恶人，使他离开所行的道，这恶人必因自己的罪孽而死，我却要从你手里讨他的血债。
EZEK|33|9|但是你，你若警戒恶人，叫他离弃所行的道，他仍不转离，他必因自己的罪孽而死，你却救了自己的命。”
EZEK|33|10|“人子啊，你要对 以色列 家说：你们曾这样说：‘我们的过犯罪恶在自己身上，我们必因此消灭，怎能存活呢？’
EZEK|33|11|你要对他们说，主耶和华说：我指着我的永生起誓，我断不喜悦恶人死亡，惟喜悦恶人转离他所行的道而存活。 以色列 家啊，你们回转，回转离开恶道吧！何必死亡呢？
EZEK|33|12|人子啊，你要对本国的百姓说：义人的义，在他犯罪之日不能救他；至于恶人的恶，在他转离恶行之日不会使他倾倒；义人在他犯罪之日不能因自己的义存活。
EZEK|33|13|我对义人说：‘你必存活！’他若倚靠自己的义作恶，所行的义就不被记念；他必因所作的恶死亡。
EZEK|33|14|我对恶人说：‘你必死亡！’他若转离他的罪恶，行公平公义的事；
EZEK|33|15|恶人若归还抵押品，归回所抢夺的东西，遵行生命的律例，不再作恶；他必存活，不致死亡。
EZEK|33|16|他所犯的一切罪必不被记念；他行了公平公义的事，必要存活。
EZEK|33|17|“你本国的百姓说：‘主的道不公平。’其实他们，他们的道才是不公平。
EZEK|33|18|义人转离自己的义作恶，他必因此而死亡。
EZEK|33|19|恶人转离他的恶，行公平公义的事，他必因此而存活。
EZEK|33|20|你们还说：‘主的道不公平。’ 以色列 家啊，我必按你们各人所行的审判你们。”
EZEK|33|21|我们被掳后第十二年的十月初五，有人从 耶路撒冷 逃到我这里，说：“城已被攻破。”
EZEK|33|22|逃来的人到的前一天晚上，耶和华的手按在我身上，开我的口。第二天早晨，等那人来到我这里，我的口就开了，不再说不出话来。
EZEK|33|23|耶和华的话临到我，说：
EZEK|33|24|“人子啊，住在 以色列 荒废之地的人说：‘ 亚伯拉罕 一人能得这地为业，我们人数众多，这地更是给我们为业的。’
EZEK|33|25|所以你要对他们说，主耶和华如此说：你们吃带血的食物，向偶像举目，并且流人的血，你们还能得这地为业吗？
EZEK|33|26|你们倚靠自己的刀剑行可憎的事，人人污辱邻舍的妻，你们还能得这地为业吗？
EZEK|33|27|你要对他们这样说，主耶和华如此说：我指着我的永生起誓，在废墟的，必倒在刀下；在田野的，必交给野兽吞吃；在堡垒和洞中的，必遭瘟疫而死。
EZEK|33|28|我必使这地荒废荒凉，它骄傲的权势也必止息； 以色列 的山都必荒废，无人经过。
EZEK|33|29|我因他们所做一切可憎的事，使地荒废荒凉；那时，他们就知道我是耶和华。”
EZEK|33|30|“你，人子啊，你本国的百姓在城墙旁边、在房屋门口谈论你。弟兄对弟兄彼此说：‘来吧！听听有什么话从耶和华而出。’
EZEK|33|31|他们如同百姓前来，来到你这里，坐在你面前仿佛是我的子民。他们听了你的话，却不实行；因为他们口里说爱，心却追随财利。
EZEK|33|32|看哪，他们看你如同一个唱情歌的人 ，声音优雅、善于奏乐；他们听了你的话，却不实行。
EZEK|33|33|看哪，这话就要应验；应验时，他们就知道在他们中间有了先知。”
EZEK|34|1|耶和华的话临到我，说：
EZEK|34|2|“人子啊，你要向 以色列 的牧人说预言，对他们说，主耶和华如此说：祸哉！ 以色列 的牧人只知牧养自己。牧人岂不当牧养群羊吗？
EZEK|34|3|你们吃肥油 、穿羊毛、宰杀肥羊，却不牧养群羊。
EZEK|34|4|瘦弱的，你们不调养；有病的，你们不医治；受伤的，你们未包扎；被逐的，你们不去领回；失丧的，你们不寻找；却用暴力严严地辖制它们 。
EZEK|34|5|它们因无牧人就分散；既分散，就成为一切野兽的食物。
EZEK|34|6|我的羊流落众山之间和各高冈上，分散在全地，无人去寻，无人去找。
EZEK|34|7|“所以，你们这些牧人要听耶和华的话。
EZEK|34|8|主耶和华说：我指着我的永生起誓，我的羊因无牧人就成为掠物，也作了一切野兽的食物。我的牧人不寻找我的羊；这些牧人只知喂养自己，并不喂养我的羊。
EZEK|34|9|所以你们这些牧人要听耶和华的话。
EZEK|34|10|主耶和华如此说：看哪，我必与牧人为敌，从他们手里讨回我的羊，使他们不再牧放群羊；牧人也不再喂养自己。我必救我的羊脱离他们的口，不再作他们的食物。”
EZEK|34|11|“主耶和华如此说：‘看哪，我必亲自寻找我的羊，将它们寻见。
EZEK|34|12|牧人在羊群四散的日子怎样寻找他的羊，我必照样寻找我的羊。这些羊在密云黑暗的日子散在各处，我要从那里救回它们。
EZEK|34|13|我要从万民中领出它们，从各国聚集它们，引领它们归回故土。我要在 以色列 山上，在一切溪水旁边，在境内所有可居住的地牧养它们。
EZEK|34|14|我要在肥美的草场牧养它们。它们的圈必在 以色列 高处的山上，它们必躺卧在佳美的圈内，在 以色列 山肥美的草场上吃草。
EZEK|34|15|我要亲自牧养我的群羊，使它们得以躺卧。这是主耶和华说的。
EZEK|34|16|失丧的，我必寻找；被逐的，我必领回；受伤的，我必包扎；有病的，我必医治；只是肥的壮的，我要除灭 ；我必秉公牧养它们。’
EZEK|34|17|“我的羊群哪，论到你们，主耶和华如此说：看哪，我要在羊与羊中间、公绵羊与公山羊中间施行审判。
EZEK|34|18|你们在肥美的草场上吃草还以为是小事吗？竟用你们的脚践踏剩下的草；你们喝了清水，竟用你们的脚搅浑剩下的水。
EZEK|34|19|至于我的羊，只能吃你们所践踏的，喝你们所搅浑的。
EZEK|34|20|“所以，主耶和华对它们如此说：看哪，我要亲自在肥羊和瘦羊中间施行审判。
EZEK|34|21|因为你们用侧边用肩推挤一切瘦弱的羊，又用角抵撞，使它们四散在外；
EZEK|34|22|所以，我要拯救我的群羊，它们必不再作掠物；我也要在羊和羊中间施行审判。
EZEK|34|23|我必在他们之上立一牧人 ，就是我的仆人 大卫 ，牧养它们；他必牧养他们，作他们的牧人。
EZEK|34|24|我─耶和华必作他们的上帝，我的仆人 大卫 要在他们中间作王。这是我─耶和华说的。
EZEK|34|25|“我要与他们立平安的约，使恶兽从境内断绝；他们在旷野也能安然居住，在树林也能躺卧。
EZEK|34|26|我要使他们和我山冈的四围蒙福；我也必叫时雨落下，使福如甘霖降下。
EZEK|34|27|田野的树木必结果子，地也必有出产；他们要在自己的土地安然居住。我折断他们所负的轭，救他们脱离奴役他们之人的手；那时，他们就知道我是耶和华。
EZEK|34|28|他们必不再作外邦人的掠物，地上的野兽也不再吞吃他们；他们却要安然居住，无人使他们惊吓。
EZEK|34|29|我必为他们建立闻名的 栽种之地；他们在境内就不再为饥荒所灭，也不再受列国的羞辱。
EZEK|34|30|他们必知道我─耶和华他们的上帝与他们同在，并知道他们， 以色列 家，是我的子民。这是主耶和华说的。
EZEK|34|31|你们这些人，你们是我的羊，我草场上的羊；我是你们的上帝。这是主耶和华说的。”
EZEK|35|1|耶和华的话临到我，说：
EZEK|35|2|“人子啊，你要面向 西珥山 ，向它说预言，
EZEK|35|3|对它说，主耶和华如此说： 西珥山 ，看哪，我与你为敌，必伸手攻击你，使你荒凉荒废。
EZEK|35|4|我必使你的城镇变为废墟，使你成为荒凉；你就知道我是耶和华。
EZEK|35|5|因为你永怀仇恨，在 以色列 人遭遇灾难、罪孽到了尽头时，把他们交给刀剑，
EZEK|35|6|所以主耶和华说：我指着我的永生起誓，我必使你遭遇血的报应，血必追赶你；你既不恨恶血，血必追赶你。
EZEK|35|7|我要使 西珥山 荒凉荒废，把来往经过的人从它那里剪除。
EZEK|35|8|我要使 西珥山 布满被杀的人。被刀杀的要倒在小山和山谷，并一切的溪水中。
EZEK|35|9|我必使你永远荒凉，使你的城镇无人居住，你们就知道我是耶和华。
EZEK|35|10|“因为你曾说‘这二国、这二邦必归我，我们必得为业’，其实耶和华仍在那里；
EZEK|35|11|所以主耶和华说：我指着我的永生起誓，我必照你因仇恨向他们发的怒气和嫉妒对待你；我审判你的时候，要在他们中间显明自己。
EZEK|35|12|你必知道我─耶和华已听见你一切凌辱的话，是针对 以色列 群山说的：‘这些山荒凉了，它们是给我们作食物的。’
EZEK|35|13|你们用口向我说夸大的话，增多与我敌对的话，我都听见了。
EZEK|35|14|主耶和华如此说：全地欢乐的时候，我必使你荒凉。
EZEK|35|15|你怎样因 以色列 家的地业荒凉而喜乐，我也要照你所做的对待你。 西珥山 哪，你和 以东 全地都必荒凉；人就知道 我是耶和华。”
EZEK|36|1|“人子啊，你要对 以色列 群山说预言： 以色列 群山哪，要听耶和华的话。
EZEK|36|2|主耶和华如此说，因仇敌说：‘啊哈！这古老的丘坛都归我们为业了！’
EZEK|36|3|所以你要预言，说：主耶和华如此说：因为敌人使你荒凉，四围践踏你，要叫你归其余的列国为业，使你们成为各族的话柄与百姓的笑谈；
EZEK|36|4|因此， 以色列 群山哪，要听主耶和华的话。对那遭四围其余列国占据、讥刺的大山小冈、水沟山谷、荒废之地、被弃之城，主耶和华如此说；
EZEK|36|5|所以，主耶和华如此说：我因妒火中烧，就责备其余的列国和 以东 的众人。他们快乐满怀，心存恨恶，将我的地占为己有，视为被抛弃的掠物。
EZEK|36|6|所以，你要指着 以色列 地说预言，对大山小冈、水沟山谷说，主耶和华如此说：看哪，我在妒忌和愤怒中宣布：因你们曾受列国的羞辱，
EZEK|36|7|所以我起誓说，你们四围的列国要担当自己的羞辱。这是主耶和华说的。
EZEK|36|8|“ 以色列 群山哪，要长出枝条，为我子民 以色列 结出果子，因为他们即将来到。
EZEK|36|9|看哪，我是帮助你们的，我要转向你们，使你们得以耕作栽种。
EZEK|36|10|我要使 以色列 全家在你们那里人数增多，城镇有人居住，废墟重新建造。
EZEK|36|11|我要使人丁和牲畜在你们那里加增，他们必生养众多。我要使你们那里像以前一样有人居住，并要赐福，比先前更多；你们就知道我是耶和华。
EZEK|36|12|我要使我的子民 以色列 在你们那里行走，他们必得你为业；你就成为他们的产业，不再使他们丧失儿女。
EZEK|36|13|主耶和华如此说，因为人对你们说‘你是吞吃人的，又使国民丧失儿女’，
EZEK|36|14|所以你必不再吞吃人，也不再使国民丧失儿女。这是主耶和华说的。
EZEK|36|15|我使你不再听见列国的羞辱；你必不再受万民的辱骂，也不再使国民绊跌。这是主耶和华说的。”
EZEK|36|16|耶和华的话临到我，说：
EZEK|36|17|“人子啊， 以色列 家住本地的时候，所作所为使那地玷污。他们的行为在我面前，好像妇人在经期中那样污秽。
EZEK|36|18|所以我因他们在那地流人的血，且以偶像使那地玷污，就把我的愤怒倾倒在他们身上。
EZEK|36|19|我将他们分散到列国，四散在列邦，按他们的所作所为惩罚他们。
EZEK|36|20|他们到了 所去的列国，使我的圣名被亵渎；因为人谈论他们说，这是耶和华的子民，却从耶和华的地出来。
EZEK|36|21|但我顾惜我的圣名，就是 以色列 家在所到的列国中亵渎的。
EZEK|36|22|“所以，你要对 以色列 家说，主耶和华如此说： 以色列 家啊，我做这事不是为你们，而是为了我的圣名，就是你们在所到的列国中亵渎的。
EZEK|36|23|我要使我至大的名显为圣；这名在列国中已遭亵渎，是你们在他们中间亵渎的。我在他们眼前，在你们身上显为圣的时候，他们就知道我是耶和华。这是主耶和华说的。
EZEK|36|24|我必从列国带领你们，从列邦聚集你们，领你们回到本地。
EZEK|36|25|我必洒清水在你们身上，你们就洁净了。我要洁净你们，使你们脱离一切的污秽，弃绝一切的偶像。
EZEK|36|26|我也要赐给你们一颗新心，将新灵放在你们里面，又从你们的肉体中除掉石心，赐给你们肉心。
EZEK|36|27|我必将我的灵放在你们里面，使你们顺从我的律例，谨守遵行我的典章。
EZEK|36|28|你们必住在我所赐给你们祖先之地；你们要作我的子民，我要作你们的上帝。
EZEK|36|29|我要救你们脱离一切的污秽，也要令五谷丰登，使你们不再遭遇饥荒。
EZEK|36|30|我要使树木多结果子，田地多出土产，好叫你们不再因饥荒被列国凌辱。
EZEK|36|31|那时，你们必追念自己的恶行和不好的作为，就因你们的罪孽和可憎的事厌恶自己。
EZEK|36|32|你们要知道，我这样做不是为你们。 以色列 家啊，你们当为自己的行为抱愧蒙羞。这是主耶和华说的。
EZEK|36|33|“主耶和华如此说：我洁净你们，使你们脱离一切罪孽的日子，必使城镇有人居住，废墟重新建造。
EZEK|36|34|这荒芜的土地，曾被过路的人看为荒芜，现今却得以耕种。
EZEK|36|35|他们必说：‘这荒芜之地，现在成了像 伊甸园 一样；这荒凉、荒废、毁坏的城镇，现今坚固，有人居住。’
EZEK|36|36|那时，在你们四围其余的列国必知道，我─耶和华修造那毁坏之处，开垦那荒芜之地。我─耶和华说了这话，就必成就。
EZEK|36|37|“主耶和华如此说：我要回应 以色列 家的求问，成全他们，增添他们的人数，使他们多如羊群。
EZEK|36|38|在 耶路撒冷 守节时，作为祭物所献的羊群有多少，照样，荒凉的城镇必为人群所充满；他们就知道我是耶和华。”
EZEK|37|1|耶和华的手按在我身上。耶和华藉着他的灵带我出去，把我放在平原中，平原遍满骸骨。
EZEK|37|2|他使我从骸骨的四围经过，看哪，平原上面的骸骨甚多，看哪，极其枯干。
EZEK|37|3|他对我说：“人子啊，这些骸骨能活过来吗？”我说：“主耶和华啊，你是知道的。”
EZEK|37|4|他又对我说：“你要向这些骸骨说预言，对它们说：枯干的骸骨啊，要听耶和华的话。
EZEK|37|5|主耶和华对这些骸骨如此说：‘看哪，我必使气息 进入你们里面，你们就要活过来。
EZEK|37|6|我要给你们加上筋，长出肉，又给你们包上皮，使气息进入你们里面，你们就要活过来；你们就知道我是耶和华。’”
EZEK|37|7|于是，我遵命说预言。正说预言的时候，有响声，看哪，有地震；骨与骨彼此接连。
EZEK|37|8|我观看，看哪，骸骨上面有筋，长了肉，又包上皮，只是里面还没有气息。
EZEK|37|9|耶和华对我说：“人子啊，你要说预言，向风 说预言。你要说，耶和华如此说：气息啊，要从四方 而来，吹在这些被杀的人身上，使他们活过来。”
EZEK|37|10|于是我遵命说预言，气息就进入骸骨，骸骨就活过来，并且用脚站起来，成为极大的军队。
EZEK|37|11|他对我说：“人子啊，这些骸骨就是 以色列 全家。他们说：‘看哪，我们的骨头枯干了，我们的指望失去了，我们灭绝净尽了！’
EZEK|37|12|所以你要说预言，对他们说，主耶和华如此说：我的子民，看哪，我要打开你们的坟墓，把你们带出坟墓，领你们进入 以色列 地。
EZEK|37|13|我的子民哪，我打开你们的坟墓，把你们带出坟墓时，你们就知道我是耶和华。
EZEK|37|14|我必将我的灵放在你们里面，你们就要活过来。我把你们安置在本地，你们就知道我─耶和华说了这话，就必成就。这是耶和华说的。”
EZEK|37|15|耶和华的话临到我，说：
EZEK|37|16|“人子啊，你要取一根木杖，在其上写‘为 犹大 和他的盟友 以色列 人’；又取一根 木杖，在其上写‘为 约瑟 ，就是 以法莲 的杖，和他的盟友 以色列 全家’。
EZEK|37|17|你要将这两根木杖彼此相接，连成一根，使它们在你手中合而为一。
EZEK|37|18|当你本国的子民对你说：‘你这是什么意思，你不指示我们吗？’
EZEK|37|19|你就对他们说，主耶和华如此说：看哪，我要将 约瑟 和他的盟友 以色列 支派的杖，就是在 以法莲 手中的那根，与 犹大 的杖接连成为一根，在我手中合而为一。
EZEK|37|20|你要在他们眼前，把写了字的那两根杖拿在手中，
EZEK|37|21|对他们说，主耶和华如此说：看哪，我要从 以色列 人所到的列国带领他们，从四围聚集他们，领他们回到本地。
EZEK|37|22|我要使他们在这地，在 以色列 群山上成为一国，必有一王作他们全体的王。他们不再成为二国，绝不再分为二国。
EZEK|37|23|他们不再因偶像和可憎的物，并一切的罪过玷污自己。我却要救他们离开一切犯罪所住的地方 ；我要洁净他们，如此，他们要作我的子民，我要作他们的上帝。’
EZEK|37|24|“我的仆人 大卫 要作他们的王；他们全体必归一个牧人。他们必顺从我的典章，谨守遵行我的律例。
EZEK|37|25|他们要住在我赐给我仆人 雅各 的地上，就是你们列祖所住之地。他们和他们的子孙，并子孙的子孙，都永远住在那里。我的仆人 大卫 要作他们的王，直到永远；
EZEK|37|26|并且我要与他们立平安的约，作为永约。我要安顿他们，使他们人数增多，又在他们中间设立我的圣所，直到永远。
EZEK|37|27|我的居所必在他们中间；我要作他们的上帝，他们要作我的子民。
EZEK|37|28|我的圣所在 以色列 人中间直到永远，列国就知道是我─耶和华使 以色列 分别为圣。”
EZEK|38|1|耶和华的话临到我，说：
EZEK|38|2|“人子啊，你要面向 玛各 地的 歌革 ，就是 米设 和 土巴 的大王，向他说预言。
EZEK|38|3|你要说，主耶和华如此说： 米设 和 土巴 的大王 歌革 ，看哪，我与你为敌。
EZEK|38|4|我要把你掉转过来，用钩子钩住你的腮颊，把你和你的军兵、马匹、骑兵都带走。他们全都披挂整齐，成为大军，佩带大小盾牌，各人拿着刀剑；
EZEK|38|5|他们当中有 波斯 人、 古实 人和 弗 人，都带着盾牌和头盔；
EZEK|38|6|还有 歌篾 人和他的军队，北方极远的 陀迦玛 族和他的军队，这许多民族都跟着你。
EZEK|38|7|“你和聚集到你那里的军队都要预备，预备妥当，你要作他们的守卫。
EZEK|38|8|过了多日，你必被差派；到末后之年，你要来到那脱离刀剑、从列国召集回来的人所住之地，来到 以色列 常久荒凉的山上；他们都从列国中被领出，在那里安然居住。
EZEK|38|9|你和你的全军，并跟随你的许多民族都要上来，如暴风刮来，如密云遮盖地面。
EZEK|38|10|“主耶和华如此说：那时，你的心必起意念，图谋恶计，
EZEK|38|11|说：‘我要上那无墙的乡村之地，到那安静的居民那里，他们无墙，无门、无闩，安然居住。
EZEK|38|12|我去那里要抢财为掳物，夺货为掠物，反手攻击那从前荒凉、现在有人居住之地，又攻击那从列国招聚出来、得了牲畜财货、住在地的高处的百姓。’
EZEK|38|13|示巴 人、 底但 人、 他施 的商人和他们的少壮狮子都对你说：‘你来是要抢财为掳物吗？你聚集军队是要夺货为掠物，夺取金银，掳去牲畜、财货，抢夺许多财宝为掳物吗？’
EZEK|38|14|“人子啊，你要因此说预言，对 歌革 说，主耶和华如此说：我的子民 以色列 安然居住时，你是知道的。
EZEK|38|15|你从你的地方，从北方极远处率领许多民族前来，他们都骑着马，是一队强而多的军兵。
EZEK|38|16|歌革 啊，你必上来攻击我的子民 以色列 ，如密云遮盖地面。末后的日子，我必领你来攻击我的地，我藉你在列国眼前显为圣的时候，他们就要认识我。
EZEK|38|17|主耶和华如此说：我在古时藉我仆人 以色列 众先知所说的，不就是你吗？ 他们在那些日子，多年说预言，我必领你来攻击 以色列 人。”
EZEK|38|18|“主耶和华说： 歌革 上来攻击 以色列 地的时候，我的怒气要从鼻孔里发出。
EZEK|38|19|我在妒忌和如火的烈怒中说：那日在 以色列 地必有大震动，
EZEK|38|20|甚至海中的鱼、天空的鸟、野地的兽，和地上爬的各种爬行动物，并地面上的众人，因见我的面就都震动；山岭崩裂，陡岩塌陷，一切的墙都必坍塌。
EZEK|38|21|我必令刀剑在我的众山攻击 歌革 ；人要用刀剑杀害弟兄。这是主耶和华说的。
EZEK|38|22|我要用瘟疫和血惩罚他。我也必降暴雨、大冰雹、火及硫磺在他和他的军队，并跟随他的许多民族身上。
EZEK|38|23|我必显为大，显为圣，在许多国家眼前显明自己；他们就知道我是耶和华。”
EZEK|39|1|“你，人子啊，要向 歌革 说预言。你要说，主耶和华如此说： 米设 和 土巴 的大王 歌革 ，看哪，我与你为敌。
EZEK|39|2|我要把你调转过来，带领你，从北方极远的地方上来，带你到 以色列 的群山上。
EZEK|39|3|我要打落你左手的弓，打掉你右手的箭。
EZEK|39|4|你和你的全军，并跟随你的列国的人，都必倒在 以色列 的群山上。我要将你给各类攫食的飞鸟和野地的走兽作食物。
EZEK|39|5|你必倒在田野，因为我曾说过，这是主耶和华说的。
EZEK|39|6|我要降火在 玛各 和海岛安然居住的人身上，他们就知道我是耶和华。
EZEK|39|7|“我要在我的子民 以色列 中彰显我的圣名，不容我的圣名再被亵渎，列国就知道我─耶和华是 以色列 中的圣者。
EZEK|39|8|看哪，时候到了，必然成就，这就是我曾说过的日子。这是主耶和华说的。
EZEK|39|9|“住 以色列 城镇的人要出去生火，用军器燃烧，就是大小盾牌、弓箭、棍棒、枪矛；用它们来烧火，直烧了七年。
EZEK|39|10|他们不必从田野捡柴，也不必从森林伐木，因为他们要用这些军器烧火。他们要抢夺那抢夺他们的人，掳掠那掳掠他们的人。这是主耶和华说的。”
EZEK|39|11|“当那日，我要把 以色列 境内、海东边的 旅人谷 给 歌革 在那里作坟地 ，阻挡了旅行的人 。在那里，人要埋葬 歌革 和他的军兵，称那地为 哈们．歌革谷 。
EZEK|39|12|以色列 家的人要用七个月埋葬他们，好使那地洁净。
EZEK|39|13|那地所有的百姓都来埋葬他们。当我得荣耀的日子，这事必叫百姓得名声。这是主耶和华说的。
EZEK|39|14|他们要分派人专职巡查遍地，埋葬那遗留在地面上入侵者的尸首，好洁净全地。过了七个月，他们还要再巡查。
EZEK|39|15|巡查的人要遍行全地，见有人的骸骨，就在旁边立一标记，等埋葬的人来将骸骨葬在 哈们．歌革谷 ，
EZEK|39|16|且有一城要取名为 哈摩那 。他们必这样洁净那地。
EZEK|39|17|“你，人子啊，主耶和华如此说：你要向各类的飞鸟和野地的走兽说：你们要聚集，来吧，从四方聚集来吃我为你们准备的祭物，就是在 以色列 的群山上丰盛的祭物，叫你们吃肉、喝血。
EZEK|39|18|你们要吃勇士的肉，喝地上领袖的血，如吃公绵羊、羔羊、公山羊、公牛；他们全都是 巴珊 的肥畜。
EZEK|39|19|你们吃我为你们准备的祭物，必吃油脂直到饱了，喝血直到醉了。
EZEK|39|20|你们要因我席上的马匹、骑兵、勇士和所有的战士而饱足。这是主耶和华说的。”
EZEK|39|21|“我要在列国中彰显我的荣耀，万国就必看见我怎样把手加在他们身上，施行审判。
EZEK|39|22|从那日以后， 以色列 家就知道我是耶和华─他们的上帝，
EZEK|39|23|列国也必知道， 以色列 家被掳掠是因他们的罪孽。他们得罪我，我就转脸不顾他们，将他们交在敌人手中，使他们全都倒在刀下。
EZEK|39|24|我照他们的污秽和罪过待他们，转脸不顾他们。
EZEK|39|25|“所以主耶和华如此说：现在，我要使 雅各 被掳的人归回，要怜悯 以色列 全家，又为我的圣名发热心。
EZEK|39|26|我将他们从万民中领回，从仇敌之地召来，在许多国家的眼前，在他们身上显为圣，他们在本地安然居住，无人使他们惊吓，那时，他们要担当 自己的羞辱和干犯我的一切罪。
EZEK|39|27|
EZEK|39|28|我使他们被掳到列国，后又聚集他们回到本地，不再留一人在那里，那时他们就知道我是耶和华─他们的上帝。
EZEK|39|29|我不再转脸不顾他们，因我已将我的灵浇灌 以色列 家。这是主耶和华说的。”
EZEK|40|1|我们被掳的第二十五年， 耶路撒冷城 攻破后十四年，正在年初，某月初十，就在那一天，耶和华的手按在我身上，把我带到那里。
EZEK|40|2|在上帝的异象中，他带我到 以色列 地，把我安置在一座极高的山上；在山的南边有仿佛一座城的建筑物。
EZEK|40|3|他带我到那里，看哪，有一人面貌 如铜，手拿麻绳和丈量的芦苇竿，站在门口。
EZEK|40|4|那人对我说：“人子啊，凡我所指示你的，你都要用眼看，用耳听，并要放在心上。我带你到这里来，为要指示你；凡你所见的，都要告诉 以色列 家。”
EZEK|40|5|看哪，殿外四围有墙。那人手拿丈量的芦苇竿，长六肘，每肘再加一掌。他量围墙，宽一竿，高一竿。
EZEK|40|6|他到了朝东的门，就上台阶，量这门的门槛，宽一竿；这门槛宽一竿。
EZEK|40|7|又有守卫房，每间长一竿，宽一竿，守卫房之间相隔五肘。挨着通往殿之门走廊的门槛，一竿。
EZEK|40|8|他量通往殿之门的走廊，一竿。
EZEK|40|9|他量门的走廊，八肘；墙柱，二肘；门的走廊通往殿那里。
EZEK|40|10|往东的门有守卫房：这旁三间，那旁三间，大小都一样；这边和那边的墙柱，大小也一样。
EZEK|40|11|他量门的入口，宽十肘，门长十三肘。
EZEK|40|12|守卫房前有矮墙，一肘，那边的矮墙也是一肘；守卫房这边六肘，那边也是六肘。
EZEK|40|13|他量门，从守卫房这边的房顶到那边的房顶，宽二十五肘；入口与入口相对。
EZEK|40|14|他量墙柱，六十肘，院子的四周围有挨着墙柱的门。
EZEK|40|15|从大门入口到里面门的走廊，五十肘。
EZEK|40|16|守卫房和四围挨着墙柱的门，都有嵌壁式的窗户，廊子也有；里面到处都有窗户，墙柱上雕刻着棕树。
EZEK|40|17|他带我到外院，看哪，院子的四围有房间，有石板地；石板地上有三十个房间。
EZEK|40|18|沿着门侧边的石板地，就是下面的石板地，与门的长度相同。
EZEK|40|19|他量宽度，从下门的前面到内院外的前面，东向北向一百肘。
EZEK|40|20|他量外院朝北的门的长和宽。
EZEK|40|21|门的守卫房，这旁三间，那旁三间；墙柱和廊子，与第一个门的大小一样。长五十肘，宽二十五肘。
EZEK|40|22|其窗户和廊子，并雕刻的棕树，与朝东的门大小一样。要登七个台阶才能上到这门，前面 有廊子。
EZEK|40|23|内院有门与这门相对，北面东面都是如此。他从这门量到那门，共一百肘。
EZEK|40|24|他带我往南去，看哪，朝南有门，他量门的墙柱 和廊子，大小与先前一样。
EZEK|40|25|门两旁与廊子的周围都有窗户，和先前量的窗户一样。门长五十肘，宽二十五肘。
EZEK|40|26|要登七个台阶才能上到这门，前面 有廊子；墙柱上雕刻着棕树，这边一棵，那边一棵。
EZEK|40|27|内院朝南也有门，从这门量到朝南的那门，共一百肘。
EZEK|40|28|他带我从南门到内院，他量南门，大小与先前一样。
EZEK|40|29|守卫房和墙柱、廊子，大小与先前一样。门两旁与廊子的周围都有窗户。门长五十肘，宽二十五肘。
EZEK|40|30|周围有廊子，长二十五肘，宽五肘。
EZEK|40|31|廊子朝着外院，墙柱上雕刻着棕树。要登八个台阶才能上到这门。
EZEK|40|32|他带我到内院的东边，他量那门，大小与先前一样。
EZEK|40|33|守卫房和墙柱、廊子，大小与先前一样。门两旁与廊子的周围都有窗户。长五十肘，宽二十五肘。
EZEK|40|34|廊子朝着外院。墙柱两边都雕刻着棕树。要登八个台阶才能上到这门。
EZEK|40|35|他带我到北门，他量了，大小与先前一样，
EZEK|40|36|就是量守卫房和墙柱、廊子。门的周围都有窗户；门长五十肘，宽二十五肘。
EZEK|40|37|墙柱 朝着外院。墙柱两边都雕刻着棕树。要登八个台阶才能上到这门。
EZEK|40|38|有房间和它的入口在门的墙柱 旁，那里是洗燔祭牲的地方。
EZEK|40|39|在门的走廊内，这边有两张桌子，那边也有两张桌子，其上可宰杀燔祭牲、赎罪祭牲和赎愆祭牲。
EZEK|40|40|上到北门的入口，朝向外面的这边有两张桌子，门的走廊那边也有两张桌子。
EZEK|40|41|门这边有四张桌子，那边也有四张桌子，共八张，在其上宰杀祭牲。
EZEK|40|42|为燔祭牲的四张桌子是用石头凿成的，长一肘半，宽一肘半，高一肘。宰杀燔祭牲和其他祭牲所用的器皿可放在其上。
EZEK|40|43|有钩子，宽一掌，挂在廊内的四周围。桌子上可放祭牲的肉。
EZEK|40|44|从外面进到内门，内院里有房间，为歌唱的人而设 ；一间在北门旁，朝南，又有一间在南 门旁，朝北。
EZEK|40|45|他对我说：“这朝南的房间是为了圣殿供职的祭司，
EZEK|40|46|那朝北的房间是为了祭坛前供职的祭司；这些祭司是 利未 人中 撒督 的子孙，近前来事奉耶和华的。”
EZEK|40|47|他又量内院，长一百肘，宽一百肘，是正方的。祭坛就在殿前。
EZEK|40|48|于是他带我到殿前的走廊，量走廊的墙柱。这面宽五肘，那面宽五肘。 门的两旁，这边三肘，那边三肘。
EZEK|40|49|走廊长二十肘，宽十一肘 。要登台阶 才能上到走廊。靠近墙柱又有柱子，这边一根，那边一根。
EZEK|41|1|他带我到殿那里，他量墙柱：这面宽六肘，那面宽六肘，宽窄与会幕相同 。
EZEK|41|2|门口宽十肘。门的两旁，这边五肘，那边五肘。他又量了殿，长四十肘，宽二十肘。
EZEK|41|3|他到内殿量门的墙柱，二肘，门口六肘，门的两旁各宽七肘。
EZEK|41|4|他量内殿，长二十肘，宽二十肘。他对我说：“这是至圣所。”
EZEK|41|5|他又量殿的墙，六肘；围着殿有厢房，各宽四肘。
EZEK|41|6|厢房有三层，层叠而上，每层排列三十间。殿的墙四周有凸出的墙支撑厢房，厢房就不必以殿的墙为支柱。
EZEK|41|7|这围绕着殿的厢房越高越宽；厢房围着殿悬叠而上，所以越上面越宽，从下一层，到中一层，到上一层。
EZEK|41|8|我又见有高台围绕着殿，作为厢房的根基，高足足有一竿，就是六大肘。
EZEK|41|9|厢房的外墙宽五肘。殿的厢房和那边的房间中间还有空地，宽二十肘，围绕着殿。
EZEK|41|10|
EZEK|41|11|厢房的门口向着空地：一门向北，一门向南。周围的空地宽五肘。
EZEK|41|12|在西边空地之后有房子，宽七十肘，长九十肘，墙四围厚五肘。
EZEK|41|13|这样，他量了殿，长一百肘，又量空地和那房子并墙，共长一百肘。
EZEK|41|14|殿的前面和东边的空地，宽一百肘。
EZEK|41|15|他量了空地后面的那房子，并两旁的楼廊，共长一百肘。 内殿、院的走廊、
EZEK|41|16|门槛 、嵌壁式的窗户，并对着门槛的三层楼廊，周围都镶上木板；地板到窗户，窗户都关着，
EZEK|41|17|直到门以上，就是到内殿和外殿内外四围墙壁，都这样测量。
EZEK|41|18|墙上雕刻基路伯和棕树，基路伯和基路伯之间有一棵棕树，每基路伯有两张脸；
EZEK|41|19|人的脸向着这边的棕树，狮子的脸向着那边的棕树，殿内四周围都是如此。
EZEK|41|20|从地板到门的上面，都有基路伯和棕树。殿的墙就是这样。
EZEK|41|21|殿的门柱是方的。至圣所的前面有个东西形状像
EZEK|41|22|木头做的坛，高三肘，长二肘 。坛角和底座 ，并四面，都是木头做的。他对我说：“这是耶和华面前的供桌。”
EZEK|41|23|殿和圣所各有一个双层门。
EZEK|41|24|每个门有两扇，每扇又有两个摺叠页；这一扇有两页，另一扇也有两页。
EZEK|41|25|殿的门扇上雕刻着基路伯和棕树，与刻在墙上的一样。在外面门的走廊前有木头做的飞檐。
EZEK|41|26|门的走廊这边和那边都有嵌壁式的窗户和棕树；殿的厢房和飞檐也是这样。
EZEK|42|1|他带我出来往北，到外院，又带我进入一个房间，一面对着空地，一面对着北边的房子。
EZEK|42|2|前面长一百肘，宽五十肘，有门向北；
EZEK|42|3|对着内院那二十肘 ，又对着外院的石板地，在第三层楼有楼廊对着楼廊。
EZEK|42|4|那些房间前有一条走道，宽十肘，往里面有宽一肘的通道 。房门都向北。
EZEK|42|5|房间因为楼廊占掉一些地方，所以房子的上层比中下两层窄。
EZEK|42|6|房间分三层，却不像外院的屋子用柱子支撑，而是从地面往上，所以一层比一层更窄。
EZEK|42|7|外面有一道墙，长五十肘，在房间前面，与朝外院的房间平行。
EZEK|42|8|靠着外院的房间长五十肘，看哪，朝圣殿的长一百肘。
EZEK|42|9|这些房间下面的东边有一个入口，从外院可由此进入；
EZEK|42|10|其宽如院墙。朝东 也有房间，一面对着空地，一面对着房子。
EZEK|42|11|这些房间前的通道与北边房间的通道一样；长、宽、出口、样式和入口都相同。
EZEK|42|12|在东边通道的开端，正对着那道墙有门可以进入，与向南边房间的门一样。
EZEK|42|13|他对我说：“面对空地南边的房间和北边的房间，都是圣的房间；亲近耶和华的祭司当在那里吃至圣的东西，也当在那里存放至圣的东西，就是素祭、赎罪祭和赎愆祭，因此处为圣。
EZEK|42|14|祭司进圣所，出来的时候，不可直接到外院，要在那里放下他们供职的衣服，因为这是圣衣；要穿上别的衣服才可以到百姓所在之处。”
EZEK|42|15|他量完了内殿的大小，就带我出朝东的门，去量院的四周围。
EZEK|42|16|他用丈量的芦苇竿量东面，五百竿 ；又转去
EZEK|42|17|用丈量的芦苇竿量北面，五百竿；又转去
EZEK|42|18|用丈量的芦苇竿量南面，五百竿。
EZEK|42|19|他又转到西面，用丈量的芦苇竿去量，五百竿。
EZEK|42|20|他量四面，长五百，宽五百，四周围有墙，为要分别圣与俗。
EZEK|43|1|以后，他带我到一座门，就是朝东的门。
EZEK|43|2|看哪， 以色列 上帝的荣光从东而来，他的声音如同众水的响声，地因他的荣耀发光。
EZEK|43|3|我所见的异象如同从前我 来灭城的时候所见的异象，又如我在 迦巴鲁河 边所见的异象，我就脸伏于地。
EZEK|43|4|耶和华的荣光从朝东的门照入殿中。
EZEK|43|5|灵将我举起，带入内院，看哪，耶和华的荣光充满了殿。
EZEK|43|6|我听见有一位从殿中向我说话，有一人站在我旁边。
EZEK|43|7|他对我说：“人子啊，这是我宝座之地，是我脚掌所踏之地。我要住在这里，住在 以色列 人中间直到永远。 以色列 家和他们的君王不可再以淫行，或在高处以君王的尸首 玷污我的圣名。
EZEK|43|8|因他们使自己的门槛挨近我的门槛，使自己的门框挨近我的门框，又使他们与我之间仅隔一墙，并且行可憎的事，玷污我的圣名，所以我发怒灭绝他们。
EZEK|43|9|现在，他们当从我面前远离淫行和君王的尸首，我就要住在他们中间，直到永远。
EZEK|43|10|“你，人子啊，要将这殿指示 以色列 家，让他们量殿的大小 ，使他们因自己的罪孽羞愧。
EZEK|43|11|他们若因自己所做的一切感到羞愧，你就要将殿的规模、样式、出口、入口，以及有关整体规模的条例、礼仪、律法指示他们 ，在他们眼前写下，使他们遵照殿整体的规模和条例去做。
EZEK|43|12|这是殿的律法：山顶上四周围的全地界都称为至圣；看哪，这就是殿的律法 。”
EZEK|43|13|这些是祭坛的大小，以肘来量，这肘是一肘一掌。底座高一肘，边宽一肘，四周围有边，高一虎口；这是祭坛的座 。
EZEK|43|14|从底座到下层的台座，二肘，边宽一肘。从小台座到大台座，四肘，边宽一肘。
EZEK|43|15|坛上的炉台，高四肘，从炉台向上突起四个角。
EZEK|43|16|这炉台长十二肘，宽十二肘，四面见方。
EZEK|43|17|台座长十四肘，宽十四肘，四面见方。四周围有边，高半肘，底座四围的边宽一肘。有台阶朝东。
EZEK|43|18|他对我说：“人子啊，主耶和华如此说：这些是建造祭坛，为要在其上献燔祭，把血洒在上面的条例：
EZEK|43|19|你要将一头公牛犊作为赎罪祭，交给那近前来事奉我的 利未 家的祭司 撒督 的后裔；这是主耶和华说的。
EZEK|43|20|你要取那公牛犊的一些血，抹在坛的四角和台座的四角，并周围的边上。你要这样洁净坛，为坛赎罪。
EZEK|43|21|你又要将那作赎罪祭的公牛烧在圣所外面，殿的预定之处。
EZEK|43|22|次日，要将无残疾的公山羊献为赎罪祭；要洁净坛，像用公牛洁净一样。
EZEK|43|23|你洁净了坛，就要将一头无残疾的公牛犊和羊群中一只无残疾的公绵羊
EZEK|43|24|奉到耶和华面前。祭司要撒盐在其上，献给耶和华为燔祭。
EZEK|43|25|七日内，你要每日献一只公山羊为赎罪祭，也要献一头公牛犊和羊群中的一只公绵羊，都要没有残疾的。
EZEK|43|26|七日内祭司要为坛赎罪，使它洁净，把它分别为圣。
EZEK|43|27|满了七日，自八日以后，祭司要在坛上献你们的燔祭和平安祭；我必悦纳你们。这是主耶和华说的。”
EZEK|44|1|他又带我回到圣所朝东的外门，那门关闭了。
EZEK|44|2|耶和华对我说：“这门必须关闭，不可敞开，谁也不可由其中进入；因为耶和华─ 以色列 的上帝已经由其中进入，所以必须关闭。
EZEK|44|3|至于君王，他必按君王的位分坐在其内，在耶和华面前吃饼。他必由这门的走廊而入，也必由此而出。”
EZEK|44|4|他又带我由北门来到殿前。我观看，看哪，耶和华的荣光充满耶和华的殿，我就脸伏于地。
EZEK|44|5|耶和华对我说：“人子啊，我对你所说耶和华殿中一切的条例和律法，你要留心，用眼看，用耳听，要留心殿的入口和圣所一切的出口。
EZEK|44|6|你要对那悖逆的 以色列 家说，主耶和华如此说： 以色列 家啊，你们行这一切可憎的事，够了吧！
EZEK|44|7|你们把我的食物，就是脂肪和血献上的时候，竟把心和肉体未受割礼的外邦人领进我的圣所，玷污我的殿；你们行这一切可憎的事，违背了我的约。
EZEK|44|8|你们未尽看守我圣物的职责，竟派别人在我的圣所替你们尽看守之责。
EZEK|44|9|“主耶和华如此说：所有心和肉体未受割礼的外邦人，就是住在 以色列 中间的任何外邦人，都不可进入我的圣所。”
EZEK|44|10|“ 以色列 人走迷的时候， 利未 人远离我，随从他们的偶像走迷离开我，他们必担当自己的罪孽。
EZEK|44|11|他们必在我的圣所当仆役，照管殿门，在殿里伺候；他们要为百姓宰杀燔祭牲和其他祭牲，站在百姓面前伺候他们。
EZEK|44|12|因为这些 利未 人曾在偶像前伺候他们，成了 以色列 家罪孽的绊脚石，所以我向他们起誓：他们必担当自己的罪孽。这是主耶和华说的。
EZEK|44|13|他们不可亲近我，作事奉我的祭司，也不可挨近我任何一件圣物，就是至圣的物；他们却要担当自己的羞辱和所行可憎之事的报应。
EZEK|44|14|我要指派他们在殿里看守，办理殿中一切事务，做一切当做的工。”
EZEK|44|15|“ 以色列 人走迷离开我的时候， 利未 家的祭司 撒督 的子孙仍然尽看守我圣所的职责；因此他们必亲近我，事奉我，并且侍立在我面前，把脂肪与血献给我。这是主耶和华说的。
EZEK|44|16|只有他们可以进我的圣所，来到我的桌前事奉我，守我吩咐的职责。
EZEK|44|17|他们进内院的门要穿细麻衣，在内院门和殿内供职时不可穿羊毛衣服。
EZEK|44|18|他们要头戴细麻布的头巾，腰穿细麻布的裤子；不可穿容易出汗的衣服。
EZEK|44|19|他们出到外院，到外院 百姓那里，要脱下供职所穿的衣服，放在圣的房间内，换上别的衣服，免得因他们的衣服使百姓成为圣。
EZEK|44|20|他们不可剃头，也不可留长发，头发一定要修剪。
EZEK|44|21|祭司进内院时不可喝酒。
EZEK|44|22|他们不可娶寡妇或被休的妇人为妻，只可娶 以色列 后裔中的处女，或祭司的寡妇。
EZEK|44|23|他们要教导我的子民分辨圣与俗，使他们知道洁净和不洁净的分别。
EZEK|44|24|有争讼的事，他们应当审判，按我的典章审判。他们要在我的节期守我的律法和条例，也当以我的安息日为圣日。
EZEK|44|25|祭司不可挨近死尸使自己不洁净，只可为父亲、母亲、儿子、女儿、兄弟和未出嫁的姊妹使自己不洁净。
EZEK|44|26|他洁净之后，他们必须再为他计算七天。
EZEK|44|27|当他进内院，入圣所，在圣所中事奉的日子，要为自己献上赎罪祭。这是主耶和华说的。
EZEK|44|28|“祭司必有产业，我就是他们的产业。不可在 以色列 中给他们基业，我就是他们的基业。
EZEK|44|29|素祭、赎罪祭和赎愆祭他们都可以吃， 以色列 中一切永献的祭物都归他们。
EZEK|44|30|各样上好的初熟之物和所献的供物，都要归祭司。你们也要将最先的面团给祭司；这样，福气就必临到你们的家。
EZEK|44|31|无论是鸟是兽，凡自然死去的，或是被撕裂的，祭司都不可吃。”
EZEK|45|1|你们抽签分地为业，要献上一份作为献给耶和华的圣地，长二万五千肘 ，宽二万 肘。整个地区都作为圣地。
EZEK|45|2|再从其中划出一块作为圣所，长五百肘，宽五百肘，四面见方；四围再加五十肘的空地。
EZEK|45|3|从这整个范围要划出长二万五千肘，宽一万肘的地，其中要有圣所，是至圣的。
EZEK|45|4|这是地上的一块圣地，要归给在圣所供职、亲近事奉耶和华的祭司，作为他们房屋用地与圣所的圣地。
EZEK|45|5|其余长二万五千肘，宽一万肘，要归给在殿中供职的 利未 人，作为他们二十间房屋 的地业。
EZEK|45|6|在那块献上的圣地旁边，你们要划分造城的地业，宽五千肘，长二万五千肘，归 以色列 全家。
EZEK|45|7|划归君王的地要在献上的圣地和城用地的两旁，面对着圣地，又面对城的用地，西至西边的疆界，东至东边的疆界，从西到东，长度与每支派所分得的一样。
EZEK|45|8|这地要在 以色列 中归君王为业。我所立的君王必不再欺压我的子民，却要按支派把地分给 以色列 家。
EZEK|45|9|主耶和华如此说：“ 以色列 的王啊，你们够了吧！要除掉残暴和抢夺的事，行公平和公义，不可再勒索我的百姓。这是主耶和华说的。
EZEK|45|10|“你们要用公道的天平、公道的伊法、公道的罢特。
EZEK|45|11|伊法要与罢特等量；一罢特为贺梅珥的十分之一，一伊法也是贺梅珥的十分之一，都以贺梅珥为计算单位。
EZEK|45|12|一舍客勒是二十季拉；二十舍客勒，二十五舍客勒，十五舍客勒，合起来为你们的一弥那。
EZEK|45|13|“你们当献的供物是这样：一贺梅珥麦子要献六分之一伊法，一贺梅珥大麦也要献六分之一伊法。
EZEK|45|14|献油的条例是这样，按油的罢特：每一歌珥油，即十罢特或一贺梅珥，要献十分之一罢特，原来十罢特等于一贺梅珥。
EZEK|45|15|从 以色列 水源丰沛的草场上，每二百只羊中要献一只羔羊。这都可作素祭、燔祭、平安祭，来为民赎罪。这是主耶和华说的。
EZEK|45|16|这地所有的百姓都要带这些供物到 以色列 王那里。
EZEK|45|17|王的本分是在节期、初一、安息日，就是 以色列 家一切的盛会，奉上燔祭、素祭、浇酒祭。他要献上赎罪祭、素祭、燔祭和平安祭，为 以色列 家赎罪。”
EZEK|45|18|主耶和华如此说：“正月初一，你要取无残疾的公牛犊，洁净圣所。
EZEK|45|19|祭司要取一些赎罪祭牲的血，抹在殿的门柱上和祭坛台座的四角上，并内院的门框上。
EZEK|45|20|本月初七，你也要为误犯罪的和因无知而犯罪的这样做；你们要为圣殿赎罪。
EZEK|45|21|“正月十四日，你们要守逾越节，七天的节期都要吃无酵饼。
EZEK|45|22|当日，王要为自己和全国百姓预备一头公牛作赎罪祭。
EZEK|45|23|节期的七天内，每天他要预备无残疾的七头公牛、七只公绵羊，给耶和华为燔祭；每天又要预备一只公山羊为赎罪祭。
EZEK|45|24|他也要预备素祭，为一头公牛同献一伊法细面，为一只公绵羊同献一伊法细面，每一伊法加一欣油。
EZEK|45|25|七月十五日守节的时候，七天他都要像这样预备赎罪祭、燔祭、素祭和油。”
EZEK|46|1|主耶和华如此说：“内院朝东的门，在六个工作的日子必须关闭；惟有安息日和初一要敞开。
EZEK|46|2|王从外面要由门的走廊进入，站在门框旁边；祭司要为他预备燔祭和平安祭，王要在门的门槛那里敬拜，然后退出。这门直到晚上不可关闭。
EZEK|46|3|安息日和初一，这地的百姓要在这门口，在耶和华面前敬拜。
EZEK|46|4|安息日，王要用六只无残疾的羔羊、一只无残疾的公绵羊，献给耶和华为燔祭；
EZEK|46|5|同献的素祭，要为公绵羊献一伊法细面，为羔羊则按照他的力量献，一伊法要加一欣油。
EZEK|46|6|初一，他要献一头无残疾的公牛犊、六只羔羊、一只公绵羊，全都要用无残疾的。
EZEK|46|7|他也要预备素祭，为公牛献一伊法细面，为公绵羊献一伊法细面，为羔羊则按照他的力量献，一伊法要加一欣油。
EZEK|46|8|王进入的时候要由这门的走廊而入，也要从原路出去。
EZEK|46|9|“在各节期，这地的百姓朝见耶和华的时候，从北门进入敬拜的，要由南门而出；从南门进入的，要由北门而出。不可从进入的门出去，要往前直行，从对面的门出去。
EZEK|46|10|他们进入时，王也跟他们一同进入；他们出去，他也要出去。
EZEK|46|11|“在节期和盛会的日子同献的素祭，要为一头公牛献一伊法细面，为一只公绵羊献一伊法细面，为羔羊则按照各人的力量献，一伊法要加一欣油。
EZEK|46|12|王奉献甘心祭，就是向耶和华甘心献的燔祭或平安祭时，当有人为他开朝东的门。他就献上燔祭和平安祭，与安息日所献的一样，然后退出。他出去之后，当有人将门关闭。”
EZEK|46|13|“每日，你要取一只无残疾一岁的羔羊献给耶和华为燔祭；要每天早晨献上。
EZEK|46|14|每天早晨你也要预备同献的素祭，六分之一伊法细面，并三分之一欣油，调和细面。这素祭要经常献给耶和华，作为永远的定例。
EZEK|46|15|每天早晨要这样献上羔羊、素祭和油，为经常献的燔祭。”
EZEK|46|16|主耶和华如此说：“王若将礼物赐给他的任何一个儿子，这就成为儿子的产业，可留给子孙，是他们所承受的地业。
EZEK|46|17|倘若王将他产业的一份赐给他的一个臣仆，这就成为他臣仆的产业，直到自由之年，然后地要归还王；王的产业终究要归自己的儿子。
EZEK|46|18|王不可夺取百姓的产业，以致赶逐他们离开自己的地业；他应该从自己的地业中将产业赐给子孙，免得我的子民离开自己的地业，四散各处。”
EZEK|46|19|他带领我从大门旁边的入口，进到朝北为祭司所预备圣的房间，看哪，西边尽头有一块土地。
EZEK|46|20|他对我说：“这是祭司煮赎愆祭牲、赎罪祭牲，烤素祭的地方，免得带出外院，使百姓成为圣。”
EZEK|46|21|他又带我出到外院，使我经过院子的四个角落，看哪，院子的每个角落都有一个小院子。
EZEK|46|22|院子四个角落有小院子，周围有墙，每个小院子长四十肘 ，宽三十肘；四个角落的小院子大小都一样，
EZEK|46|23|小院子周围各有一排石墙，每排石墙下面有炉灶。
EZEK|46|24|他对我说：“这些是煮肉用的屋子，殿内的仆役要在这里煮百姓的祭物。”
EZEK|47|1|他带我回到殿门，看哪，有水从殿的门槛下面往东流出，因为这殿是朝东的。水从殿的侧面，就是右边，从祭坛的南边往下流。
EZEK|47|2|他带我出北门，又领我从外边转到朝东的外门，看哪，水从右边流出。
EZEK|47|3|他手拿绳子往东出去，量了一千肘，使我涉水而过，水到脚踝。
EZEK|47|4|他又量了一千，使我涉水而过，水就到膝；再量了一千，使我过去，水就到腰；
EZEK|47|5|又量了一千，水已成河，无法过去；因为水势高涨成河，只能游泳，无法走过。
EZEK|47|6|他对我说：“人子啊，你看见了吗？” 他带我回到河边。
EZEK|47|7|我回到河边时，看哪，河这边与那边的岸上有极多的树木。
EZEK|47|8|他对我说：“这水往东方流，下到 亚拉巴 ，直到海。所流出来的水，一入海 就使水变淡 。
EZEK|47|9|这两条河 所到之处，凡滋生的动物都必存活；这水流到那里，使那里的水变淡，因此里面有极多的鱼。这河水所到之处，百物都必存活。
EZEK|47|10|必有渔夫站在河边，从 隐．基底 直到 隐．以革莲 ，全都成了晒 网的场所。那里的鱼各从其类，好像大海的鱼甚多。
EZEK|47|11|但是沼泽与池塘的水无法变淡，只能作产盐之用。
EZEK|47|12|河这边与那边的岸上必生长各类树木，可作食物；叶子不枯干，果子不断绝。每月必结新果子，因为这水是从圣所流出来的。树上的果子必作食物，叶子可以治病。”
EZEK|47|13|主耶和华如此说：“这是你们按 以色列 十二支派分地为业的地界， 约瑟 要得两份。
EZEK|47|14|你们承受这地为业，要彼此均分；我曾起誓应许将这地赐给你们的列祖，这地必归你们为业。
EZEK|47|15|“这地的疆界如下：北界从 大海 往 希特伦 ，直到 西达达 口；
EZEK|47|16|又往 哈马 、 比罗他 、 西伯莲 ( 西伯莲 在 大马士革 的边界与 哈马 的边界中间)，到 浩兰 边界的 哈撒．哈提干 。
EZEK|47|17|这样，疆界是从 大海 往 大马士革 地界上的 哈萨．以难 ，北边以 哈马 为界。这是北界。
EZEK|47|18|“东界在 浩兰 和 大马士革 中间， 基列 和 以色列 地的中间，以 约旦河 为界。你们要量疆界直到东海 。这是东界。
EZEK|47|19|“南界是从 他玛 到 加低斯 的 米利巴 水，经 埃及 溪谷 ，直到 大海 。这是南界。
EZEK|47|20|“西界就是 大海 ，从南界直到 哈马口 对面。这是西界。
EZEK|47|21|“你们要为自己按 以色列 的支派分这地。
EZEK|47|22|要抽签分这地为业，归自己和那在你们中间寄居，生儿育女的外人。你们要看他们如本地出生的 以色列 人，他们要在 以色列 支派中与你们同得地业。
EZEK|47|23|外人寄居在哪个支派，你们就在哪里将地业分给他们。这是主耶和华说的。”
EZEK|48|1|众支派的名字如下：从北边尽头，由 希特伦 往 哈马 口，到 大马士革 地界上的 哈萨．以难 。北边靠着 哈马 地，从东到西是 但 的一份。
EZEK|48|2|靠着 但 的地界，从东到西，是 亚设 的一份。
EZEK|48|3|靠着 亚设 的地界，从东到西，是 拿弗他利 的一份。
EZEK|48|4|靠着 拿弗他利 的地界，从东到西，是 玛拿西 的一份。
EZEK|48|5|靠着 玛拿西 的地界，从东到西，是 以法莲 的一份。
EZEK|48|6|靠着 以法莲 的地界，从东到西，是 吕便 的一份。
EZEK|48|7|靠着 吕便 的地界，从东到西，是 犹大 的一份。
EZEK|48|8|靠着 犹大 的地界，从东到西，必有你们所当献的圣地，宽二万五千肘 ；长短与各族从东到西所分的地相同，圣所当在其中。
EZEK|48|9|你们献给耶和华的圣地要长二万五千肘，宽一万肘。
EZEK|48|10|这圣地要归祭司，北长二万五千肘，西宽一万肘，东宽一万肘，南长二万五千肘。耶和华的圣所当在其中。
EZEK|48|11|这地要归 撒督 的子孙中成为圣的祭司，他们谨守我所吩咐的；当 以色列 人走迷的时候，他们不像那些 利未 人走迷了。
EZEK|48|12|在圣地中要特别保留一份归他们，为至圣，紧邻着 利未 人的地界。
EZEK|48|13|利未 人所得的地长二万五千肘，宽一万肘，与祭司的地界相等，都长二万五千肘，宽一万肘。
EZEK|48|14|这地不可卖，不可换；这上好的部分不可转让给别人，因为它归耶和华为圣。
EZEK|48|15|剩下的地长二万五千肘、宽五千肘，要作公用，为造城、盖房、空地之用；城要在中间。
EZEK|48|16|以下是城的大小：北面四千五百肘，南面四千五百肘，东面四千五百肘，西面四千五百肘。
EZEK|48|17|城要有空地，向北二百五十肘，向南二百五十肘，向东二百五十肘，向西二百五十肘。
EZEK|48|18|靠着圣地并排剩余的，东长一万肘，西长一万肘；它与圣地并排，其中所出产的要作城内工人的食物。
EZEK|48|19|以色列 支派中所有在城内做工的，都要耕种这地。
EZEK|48|20|你们要将整块四方的圣地，长二万五千肘，宽二万五千肘，连同城的用地都献作圣地。
EZEK|48|21|圣地和城的用地两边剩余的要归给王。地的东边，南北二万五千肘，东至东界；西边，南北二万五千肘，西至西界；靠着各支派所分的地，都要归给王。圣地和殿的圣所要在其中。
EZEK|48|22|利未 人的地与城的用地都在王的地中间， 犹大 边界和 便雅悯 边界之间，要归给王。
EZEK|48|23|论到其余的支派，从东到西，是 便雅悯 的一份。
EZEK|48|24|靠着 便雅悯 的地界，从东到西，是 西缅 的一份。
EZEK|48|25|靠着 西缅 的地界，从东到西，是 以萨迦 的一份。
EZEK|48|26|靠着 以萨迦 的地界，从东到西，是 西布伦 的一份。
EZEK|48|27|靠着 西布伦 的地界，从东到西，是 迦得 的一份。
EZEK|48|28|靠着 迦得 南边的地界，界限从 他玛 到 加低斯 的 米利巴 水，经 埃及 溪谷 ，直到 大海 。
EZEK|48|29|这就是你们要抽签分给 以色列 支派为业之地，是他们各支派所得的份。这是主耶和华说的。
EZEK|48|30|以下是城的出口：北面四千五百肘，
EZEK|48|31|城的各门要按 以色列 的支派命名。北面有三个门，一为 吕便 门，一为 犹大 门，一为 利未 门。
EZEK|48|32|东面四千五百肘，有三个门，一为 约瑟 门，一为 便雅悯 门，一为 但 门。
EZEK|48|33|南面四千五百肘，有三个门，一为 西缅 门，一为 以萨迦 门，一为 西布伦 门。
EZEK|48|34|西面四千五百肘，有三个门，一为 迦得 门，一为 亚设 门，一为 拿弗他利 门。
EZEK|48|35|城的周围共一万八千肘。从此以后，这城的名字必称为“耶和华的所在”。
