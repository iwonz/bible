PHLM|1|1|Paul, a prisoner for Christ Jesus, and Timothy our brother, To Philemon our beloved fellow worker
PHLM|1|2|and Apphia our sister and Archippus our fellow soldier, and the church in your house:
PHLM|1|3|Grace to you and peace from God our Father and the Lord Jesus Christ.
PHLM|1|4|I thank my God always when I remember you in my prayers,
PHLM|1|5|because I hear of your love and of the faith that you have toward the Lord Jesus and all the saints,
PHLM|1|6|and I pray that the sharing of your faith may become effective for the full knowledge of every good thing that is in us for the sake of Christ.
PHLM|1|7|For I have derived much joy and comfort from your love, my brother, because the hearts of the saints have been refreshed through you.
PHLM|1|8|Accordingly, though I am bold enough in Christ to command you to do what is required,
PHLM|1|9|yet for love's sake I prefer to appeal to you- I, Paul, an old man and now a prisoner also for Christ Jesus-
PHLM|1|10|I appeal to you for my child, Onesimus, whose father I became in my imprisonment.
PHLM|1|11|(Formerly he was useless to you, but now he is indeed useful to you and to me.)
PHLM|1|12|I am sending him back to you, sending my very heart.
PHLM|1|13|I would have been glad to keep him with me, in order that he might serve me on your behalf during my imprisonment for the gospel,
PHLM|1|14|but I preferred to do nothing without your consent in order that your goodness might not be by compulsion but of your own free will.
PHLM|1|15|For this perhaps is why he was parted from you for a while, that you might have him back forever,
PHLM|1|16|no longer as a slave but more than a slave, as a beloved brother- especially to me, but how much more to you, both in the flesh and in the Lord.
PHLM|1|17|So if you consider me your partner, receive him as you would receive me.
PHLM|1|18|If he has wronged you at all, or owes you anything, charge that to my account.
PHLM|1|19|I, Paul, write this with my own hand: I will repay it- to say nothing of your owing me even your own self.
PHLM|1|20|Yes, brother, I want some benefit from you in the Lord. Refresh my heart in Christ.
PHLM|1|21|Confident of your obedience, I write to you, knowing that you will do even more than I say.
PHLM|1|22|At the same time, prepare a guest room for me, for I am hoping that through your prayers I will be graciously given to you.
PHLM|1|23|Epaphras, my fellow prisoner in Christ Jesus, sends greetings to you,
PHLM|1|24|and so do Mark, Aristarchus, Demas, and Luke, my fellow workers.
PHLM|1|25|The grace of the Lord Jesus Christ be with your spirit.
