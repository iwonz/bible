2TIM|1|1|Павло, з волі Божої апостол Христа Ісуса, за обітницею життя, що в Христі Ісусі,
2TIM|1|2|до Тимофія, сина улюбленого: благодать, милість, мир від Бога Отця й Христа Ісуса, Господа нашого!
2TIM|1|3|Дякую Богові, Якому служу від предків чистим сумлінням, що тебе пам'ятаю я завжди в молитвах своїх день і ніч.
2TIM|1|4|Я бажаю побачити тебе, пам'ятаючи сльози твої, щоб наповнитись радістю.
2TIM|1|5|Я приводжу на пам'ять собі твою нелицемірну віру, що перше була оселилася в бабі твоїй Лоіді та в твоїй матері Евнікії; певен же я, що й у тобі вона оселилась.
2TIM|1|6|З цієї причини я нагадую тобі, що ти розгрівав Божого дара, який у тобі через покладання рук моїх.
2TIM|1|7|Бо не дав нам Бог духа страху, але сили, і любови, і здорового розуму.
2TIM|1|8|Тож, не соромся засвідчення Господа нашого, ні мене, Його в'язня, але страждай з Євангелією за силою Бога,
2TIM|1|9|що нас спас і покликав святим покликом, не за наші діла, але з волі Своєї та з благодаті, що нам дана в Христі Ісусі попереду вічних часів.
2TIM|1|10|А тепер об'явилась через з'явлення Спасителя нашого Христа Ісуса, що й смерть зруйнував, і вивів на світло життя та нетління Євангелією,
2TIM|1|11|що для неї я був настановлений за проповідника, апостола й учителя.
2TIM|1|12|З цієї причини й терплю я оце, але не соромлюсь, бо знаю, в Кого я ввірував та впевнився, що має Він силу заховати на той день заставу мою.
2TIM|1|13|Май же за взір здорових слів ті, які від мене почув ти у вірі й любові, що в Христі Ісусі вона.
2TIM|1|14|Добро припоручене стережи Святим Духом, що в нас пробуває.
2TIM|1|15|Ти знаєш оце, що відвернулись від мене всі, хто в Азії, а між ними Фігел та Гермоген.
2TIM|1|16|Хай Господь подасть милосердя Онисифоровому дому, бо він часто мене підкріпляв і кайданів моїх не соромився.
2TIM|1|17|А коли він до Риму прибув, шукав мене пильно й знайшов,
2TIM|1|18|хай Господь йому дасть знайти милість від Господа в день той, скільки ж він послужив був в Ефесі мені, ти відаєш краще!
2TIM|2|1|Отож, сину мій, зміцняйся в благодаті, що в Христі Ісусі вона!
2TIM|2|2|А що чув ти від мене при багатьох свідках, те передай вірним людям, що будуть спроможні й інших навчити.
2TIM|2|3|А ти терпи лихо, як добрий вояк Христа Ісуса!
2TIM|2|4|Бо жаден вояк не в'яжеться в справи життя, аби догодити тому, хто військо збирає.
2TIM|2|5|А як хто йде на змаги, то вінка не одержує, якщо незаконно змагається.
2TIM|2|6|Трудящому хліборобові належиться першому покуштувати з плоду.
2TIM|2|7|Розумій, що я говорю. А Господь нехай дасть тобі розум у всьому.
2TIM|2|8|Пам'ятай про Ісуса Христа з насіння Давидового, що воскрес із мертвих, за моєю Євангелією,
2TIM|2|9|за яку я терплю муки аж до ув'язнення, як той злочинець. Але Слова Божого не ув'язнити!
2TIM|2|10|Через це переношу я все ради вибраних, щоб і вони доступили спасіння, що в Христі Ісусі, зо славою вічною.
2TIM|2|11|Вірне слово: коли разом із Ним ми померли, то й житимемо разом із Ним!
2TIM|2|12|А коли терпимо, то будемо разом також царювати. А коли відцураємось, то й Він відцурається нас!
2TIM|2|13|А коли ми невірні, зостається Він вірним, бо не може зректися Самого Себе!
2TIM|2|14|Нагадуй про це й заклинай перед Богом, щоб не сперечались словами, бо нінащо воно, хіба слухачам на руїну.
2TIM|2|15|Силкуйся поставити себе перед Богом гідним, працівником бездоганним, що вірно навчає науки правди.
2TIM|2|16|Стережися ж базікань марних, бо вони ще більше провадять до безбожности,
2TIM|2|17|а їхнє слово, як рак, буде ширитися. Від таких Гіменей і Філіт,
2TIM|2|18|що вони погрішилися в правді, казавши, що воскресіння було вже, і віру деяких руйнують.
2TIM|2|19|Та однако стоїть міцна Божа основа та має печатку оцю: Господь знає тих, хто Його, та: Нехай від неправди відступиться всякий, хто Господнє Ім'я називає!
2TIM|2|20|А в великому домі знаходиться посуд не тільки золотий та срібний, але й дерев'яний та глиняний, і одні посудини на честь, а другі на нечесть.
2TIM|2|21|Отож, хто від цього очистить себе, буде посуд на честь, освячений, потрібний Володареві, приготований на всяке добре діло.
2TIM|2|22|Стережися молодечих пожадливостей, тримайся правди, віри, любови, миру з тими, хто Господа кличе від чистого серця.
2TIM|2|23|А від нерозумних та від невчених змагань ухиляйся, знавши, що вони родять сварки.
2TIM|2|24|А раб Господній не повинен сваритись, але бути привітним до всіх, навчальним, до лиха терплячим,
2TIM|2|25|що навчав би противників із лагідністю, чи Бог їм не дасть покаяння, щоб правду пізнати,
2TIM|2|26|щоб визволитися від сітки диявола, що він уловив їх для роблення волі своєї.
2TIM|3|1|Знай же ти це, що останніми днями настануть тяжкі часи.
2TIM|3|2|Будуть бо люди тоді самолюбні, грошолюбні, зарозумілі, горді, богозневажники, батькам неслухняні, невдячні, непобожні,
2TIM|3|3|нелюбовні, запеклі, осудливі, нестримливі, жорстокі, ненависники добра,
2TIM|3|4|зрадники, нахабні, бундючні, що більше люблять розкоші, аніж люблять Бога,
2TIM|3|5|вони мають вигляд благочестя, але сили його відреклися. Відвертайсь від таких!
2TIM|3|6|До них бо належать і ті, хто пролазить до хат та зводить жінок, гріхами обтяжених, ведених усякими пожадливостями,
2TIM|3|7|що вони завжди вчаться, та ніколи не можуть прийти до пізнання правди.
2TIM|3|8|Як Янній та Ямврій протиставилися були Мойсеєві, так і ці протиставляться правді, люди зіпсутого розуму, неуки щодо віри.
2TIM|3|9|Та більше не матимуть успіху, бо всім виявиться їхній безум, як і з тими було.
2TIM|3|10|Ти ж пішов услід за мною наукою, поступованням, заміром, вірою, витривалістю, любов'ю, терпеливістю,
2TIM|3|11|переслідуваннями та стражданнями, що спіткали були мене в Антіохії, в Іконії, у Лістрах, такі переслідування переніс я, та Господь від усіх мене визволив.
2TIM|3|12|Та й усі, хто хоче жити побожно у Христі Ісусі, будуть переслідувані.
2TIM|3|13|А люди лихі та дурисвіти матимуть успіх у злому, зводячи й зведені бувши.
2TIM|3|14|А ти в тім пробувай, чого тебе навчено, і що тобі звірено, відаючи тих, від кого навчився був ти.
2TIM|3|15|І ти знаєш з дитинства Писання святе, що може зробити тебе мудрим на спасіння вірою в Христа Ісуса.
2TIM|3|16|Усе Писання Богом надхнене, і корисне до навчання, до докору, до направи, до виховання в праведності,
2TIM|3|17|щоб Божа людина була досконала, до всякого доброго діла готова.
2TIM|4|1|Отже, я свідкую тобі перед Богом і Христом Ісусом, що Він має судити живих і мертвих за Свого приходу та за Свого Царства.
2TIM|4|2|Проповідуй Слово, допоминайся вчасно-невчасно, докоряй, забороняй, переконуй з терпеливістю та з наукою.
2TIM|4|3|Настане бо час, коли здорової науки не будуть триматись, але за своїми пожадливостями виберуть собі вчителів, щоб вони їхні вуха влещували.
2TIM|4|4|Вони слух свій від правди відвернуть та до байок нахиляться.
2TIM|4|5|Але ти будь пильний у всьому, терпи лихо, виконуй працю благовісника, сповняй свою службу.
2TIM|4|6|Бо я вже за жертву стаю, і час відходу мого вже настав.
2TIM|4|7|Я змагався добрим змагом, свій біг закінчив, віру зберіг.
2TIM|4|8|Наостанку мені призначається вінок праведности, якого мені того дня дасть Господь, Суддя праведний; і не тільки мені, але й усім, хто прихід Його полюбив.
2TIM|4|9|Подбай незабаром прибути до мене.
2TIM|4|10|Бо Димас мене кинув, цей вік полюбивши, і пішов до Солуня, Крискент до Галатії, Тит до Далматії.
2TIM|4|11|Зо мною сам тільки Лука. Візьми Марка, і приведи з собою, бо мені він потрібний для служби.
2TIM|4|12|А Тихика послав я в Ефес.
2TIM|4|13|Як будеш іти, то плаща принеси, що його я в Троаді зоставив у Карпа, і книжки, особливо пергаменові.
2TIM|4|14|Котляр Олександер накоїв був лиха чимало мені... Нехай Господь йому віддасть за його вчинками!
2TIM|4|15|Стережись його й ти, бо він міцно противився нашим словам!
2TIM|4|16|При першій моїй обороні жаден не був при мені, але всі покинули мене... Хай Господь їм того не полічить!
2TIM|4|17|Але Господь став при мені та й мене підкріпив, щоб проповідь виконалась через мене, та щоб усі погани почули її. І я визволився з пащі лев'ячої...
2TIM|4|18|А від усякого вчинку лихого Господь мене визволить та збереже для Свого Небесного Царства. Йому слава на віки вічні, амінь!
2TIM|4|19|Поздоров Прискиллу й Акилу та дім Онисифора.
2TIM|4|20|Ераст позостався в Коринті, а Трохима лишив я слабого в Мілеті.
2TIM|4|21|Попильнуй прийти до зими. Вітає тебе Еввул, і Пуд, і Лин, і Клавдія, і вся браття.
2TIM|4|22|Господь з твоїм духом! Благодать з вами! Амінь.
