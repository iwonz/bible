MAL|1|1|The oracle of the word of the LORD to Israel by Malachi.
MAL|1|2|"I have loved you," says the LORD. But you say, "How have you loved us?" "Is not Esau Jacob's brother?" declares the LORD. "Yet I have loved Jacob
MAL|1|3|but Esau I have hated. I have laid waste his hill country and left his heritage to jackals of the desert."
MAL|1|4|If Edom says, "We are shattered but we will rebuild the ruins," the LORD of hosts says, "They may build, but I will tear down, and they will be called 'the wicked country,' and 'the people with whom the LORD is angry forever.'"
MAL|1|5|Your own eyes shall see this, and you shall say, "Great is the LORD beyond the border of Israel!"
MAL|1|6|"A son honors his father, and a servant his master. If then I am a father, where is my honor? And if I am a master, where is my fear? says the LORD of hosts to you, O priests, who despise my name. But you say, 'How have we despised your name?'
MAL|1|7|By offering polluted food upon my altar. But you say, 'How have we polluted you?' By saying that the LORD's table may be despised.
MAL|1|8|When you offer blind animals in sacrifice, is that not evil? And when you offer those that are lame or sick, is that not evil? Present that to your governor; will he accept you or show you favor? says the LORD of hosts.
MAL|1|9|And now entreat the favor of God, that he may be gracious to us. With such a gift from your hand, will he show favor to any of you? says the LORD of hosts.
MAL|1|10|Oh that there were one among you who would shut the doors, that you might not kindle fire on my altar in vain! I have no pleasure in you, says the LORD of hosts, and I will not accept an offering from your hand.
MAL|1|11|For from the rising of the sun to its setting my name will be great among the nations, and in every place incense will be offered to my name, and a pure offering. For my name will be great among the nations, says the LORD of hosts.
MAL|1|12|But you profane it when you say that the Lord's table is polluted, and its fruit, that is, its food may be despised.
MAL|1|13|But you say, 'What a weariness this is,' and you snort at it, says the LORD of hosts. You bring what has been taken by violence or is lame or sick, and this you bring as your offering! Shall I accept that from your hand? says the LORD.
MAL|1|14|Cursed be the cheat who has a male in his flock, and vows it, and yet sacrifices to the Lord what is blemished. For I am a great King, says the LORD of hosts, and my name will be feared among the nations.
MAL|2|1|"And now, O priests, this command is for you.
MAL|2|2|If you will not listen, if you will not take it to heart to give honor to my name, says the LORD of hosts, then I will send the curse upon you and I will curse your blessings. Indeed, I have already cursed them, because you do not lay it to heart.
MAL|2|3|Behold, I will rebuke your offspring, and spread dung on your faces, the dung of your offerings, and you shall be taken away with it.
MAL|2|4|So shall you know that I have sent this command to you, that my covenant with Levi may stand, says the LORD of hosts.
MAL|2|5|My covenant with him was one of life and peace, and I gave them to him. It was a covenant of fear, and he feared me. He stood in awe of my name.
MAL|2|6|True instruction was in his mouth, and no wrong was found on his lips. He walked with me in peace and uprightness, and he turned many from iniquity.
MAL|2|7|For the lips of a priest should guard knowledge, and people should seek instruction from his mouth, for he is the messenger of the LORD of hosts.
MAL|2|8|But you have turned aside from the way. You have caused many to stumble by your instruction. You have corrupted the covenant of Levi, says the LORD of hosts,
MAL|2|9|and so I make you despised and abased before all the people, inasmuch as you do not keep my ways but show partiality in your instruction."
MAL|2|10|Have we not all one Father? Has not one God created us? Why then are we faithless to one another, profaning the covenant of our fathers?
MAL|2|11|Judah has been faithless, and abomination has been committed in Israel and in Jerusalem. For Judah has profaned the sanctuary of the LORD, which he loves, and has married the daughter of a foreign god.
MAL|2|12|May the LORD cut off from the tents of Jacob, any descendant of the man who does this, who brings an offering to the LORD of hosts!
MAL|2|13|And this second thing you do. You cover the LORD's altar with tears, with weeping and groaning because he no longer regards the offering or accepts it with favor from your hand.
MAL|2|14|But you say, "Why does he not?" Because the LORD was witness between you and the wife of your youth, to whom you have been faithless, though she is your companion and your wife by covenant.
MAL|2|15|Did he not make them one, with a portion of the Spirit in their union? And what was the one God seeking? Godly offspring. So guard yourselves in your spirit, and let none of you be faithless to the wife of your youth.
MAL|2|16|"For the man who hates and divorces, says the LORD, the God of Israel, covers his garment with violence, says the LORD of hosts. So guard yourselves in your spirit, and do not be faithless."
MAL|2|17|You have wearied the LORD with your words. But you say, "How have we wearied him?" By saying, "Everyone who does evil is good in the sight of the LORD, and he delights in them." Or by asking, "Where is the God of justice?"
MAL|3|1|"Behold, I send my messenger and he will prepare the way before me. And the Lord whom you seek will suddenly come to his temple; and the messenger of the covenant in whom you delight, behold, he is coming, says the LORD of hosts.
MAL|3|2|But who can endure the day of his coming, and who can stand when he appears? For he is like a refiner's fire and like fullers' soap.
MAL|3|3|He will sit as a refiner and purifier of silver, and he will purify the sons of Levi and refine them like gold and silver, and they will bring offerings in righteousness to the LORD.
MAL|3|4|Then the offering of Judah and Jerusalem will be pleasing to the LORD as in the days of old and as in former years.
MAL|3|5|"Then I will draw near to you for judgment. I will be a swift witness against the sorcerers, against the adulterers, against those who swear falsely, against those who oppress the hired worker in his wages, the widow and the fatherless, against those who thrust aside the sojourner, and do not fear me, says the LORD of hosts.
MAL|3|6|"For I the LORD do not change; therefore you, O children of Jacob, are not consumed.
MAL|3|7|From the days of your fathers you have turned aside from my statutes and have not kept them. Return to me, and I will return to you, says the LORD of hosts. But you say, 'How shall we return?'
MAL|3|8|Will man rob God? Yet you are robbing me. But you say, 'How have we robbed you?' In your tithes and contributions.
MAL|3|9|You are cursed with a curse, for you are robbing me, the whole nation of you.
MAL|3|10|Bring the full tithes into the storehouse, that there may be food in my house. And thereby put me to the test, says the LORD of hosts, if I will not open the windows of heaven for you and pour down for you a blessing until there is no more need.
MAL|3|11|I will rebuke the devourer for you, so that it will not destroy the fruits of your soil, and your vine in the field shall not fail to bear, says the LORD of hosts.
MAL|3|12|Then all nations will call you blessed, for you will be a land of delight, says the LORD of hosts.
MAL|3|13|"Your words have been hard against me, says the LORD. But you say, 'How have we spoken against you?'
MAL|3|14|You have said, 'It is vain to serve God. What is the profit of our keeping his charge or of walking as in mourning before the LORD of hosts?
MAL|3|15|And now we call the arrogant blessed. Evildoers not only prosper but they put God to the test and they escape.'"
MAL|3|16|Then those who feared the LORD spoke with one another. The LORD paid attention and heard them, and a book of remembrance was written before him of those who feared the LORD and esteemed his name.
MAL|3|17|"They shall be mine, says the LORD of hosts, in the day when I make up my treasured possession, and I will spare them as a man spares his son who serves him.
MAL|3|18|Then once more you shall see the distinction between the righteous and the wicked, between one who serves God and one who does not serve him.
MAL|4|1|"For behold, the day is coming, burning like an oven, when all the arrogant and all evildoers will be stubble. The day that is coming shall set them ablaze, says the LORD of hosts, so that it will leave them neither root nor branch.
MAL|4|2|But for you who fear my name, the sun of righteousness shall rise with healing in its wings. You shall go out leaping like calves from the stall.
MAL|4|3|And you shall tread down the wicked, for they will be ashes under the soles of your feet, on the day when I act, says the LORD of hosts.
MAL|4|4|"Remember the law of my servant Moses, the statutes and rules that I commanded him at Horeb for all Israel.
MAL|4|5|"Behold, I will send you Elijah the prophet before the great and awesome day of the LORD comes.
MAL|4|6|And he will turn the hearts of fathers to their children and the hearts of children to their fathers, lest I come and strike the land with a decree of utter destruction."
