DEUT|1|1|These are the words Moses spoke to all Israel in the desert east of the Jordan-that is, in the Arabah-opposite Suph, between Paran and Tophel, Laban, Hazeroth and Dizahab.
DEUT|1|2|(It takes eleven days to go from Horeb to Kadesh Barnea by the Mount Seir road.)
DEUT|1|3|In the fortieth year, on the first day of the eleventh month, Moses proclaimed to the Israelites all that the LORD had commanded him concerning them.
DEUT|1|4|This was after he had defeated Sihon king of the Amorites, who reigned in Heshbon, and at Edrei had defeated Og king of Bashan, who reigned in Ashtaroth.
DEUT|1|5|East of the Jordan in the territory of Moab, Moses began to expound this law, saying:
DEUT|1|6|The LORD our God said to us at Horeb, "You have stayed long enough at this mountain.
DEUT|1|7|Break camp and advance into the hill country of the Amorites; go to all the neighboring peoples in the Arabah, in the mountains, in the western foothills, in the Negev and along the coast, to the land of the Canaanites and to Lebanon, as far as the great river, the Euphrates.
DEUT|1|8|See, I have given you this land. Go in and take possession of the land that the LORD swore he would give to your fathers-to Abraham, Isaac and Jacob-and to their descendants after them."
DEUT|1|9|At that time I said to you, "You are too heavy a burden for me to carry alone.
DEUT|1|10|The LORD your God has increased your numbers so that today you are as many as the stars in the sky.
DEUT|1|11|May the LORD, the God of your fathers, increase you a thousand times and bless you as he has promised!
DEUT|1|12|But how can I bear your problems and your burdens and your disputes all by myself?
DEUT|1|13|Choose some wise, understanding and respected men from each of your tribes, and I will set them over you."
DEUT|1|14|You answered me, "What you propose to do is good."
DEUT|1|15|So I took the leading men of your tribes, wise and respected men, and appointed them to have authority over you-as commanders of thousands, of hundreds, of fifties and of tens and as tribal officials.
DEUT|1|16|And I charged your judges at that time: Hear the disputes between your brothers and judge fairly, whether the case is between brother Israelites or between one of them and an alien.
DEUT|1|17|Do not show partiality in judging; hear both small and great alike. Do not be afraid of any man, for judgment belongs to God. Bring me any case too hard for you, and I will hear it.
DEUT|1|18|And at that time I told you everything you were to do.
DEUT|1|19|Then, as the LORD our God commanded us, we set out from Horeb and went toward the hill country of the Amorites through all that vast and dreadful desert that you have seen, and so we reached Kadesh Barnea.
DEUT|1|20|Then I said to you, "You have reached the hill country of the Amorites, which the LORD our God is giving us.
DEUT|1|21|See, the LORD your God has given you the land. Go up and take possession of it as the LORD, the God of your fathers, told you. Do not be afraid; do not be discouraged."
DEUT|1|22|Then all of you came to me and said, "Let us send men ahead to spy out the land for us and bring back a report about the route we are to take and the towns we will come to."
DEUT|1|23|The idea seemed good to me; so I selected twelve of you, one man from each tribe.
DEUT|1|24|They left and went up into the hill country, and came to the Valley of Eshcol and explored it.
DEUT|1|25|Taking with them some of the fruit of the land, they brought it down to us and reported, "It is a good land that the LORD our God is giving us."
DEUT|1|26|But you were unwilling to go up; you rebelled against the command of the LORD your God.
DEUT|1|27|You grumbled in your tents and said, "The LORD hates us; so he brought us out of Egypt to deliver us into the hands of the Amorites to destroy us.
DEUT|1|28|Where can we go? Our brothers have made us lose heart. They say, 'The people are stronger and taller than we are; the cities are large, with walls up to the sky. We even saw the Anakites there.'"
DEUT|1|29|Then I said to you, "Do not be terrified; do not be afraid of them.
DEUT|1|30|The LORD your God, who is going before you, will fight for you, as he did for you in Egypt, before your very eyes,
DEUT|1|31|and in the desert. There you saw how the LORD your God carried you, as a father carries his son, all the way you went until you reached this place."
DEUT|1|32|In spite of this, you did not trust in the LORD your God,
DEUT|1|33|who went ahead of you on your journey, in fire by night and in a cloud by day, to search out places for you to camp and to show you the way you should go.
DEUT|1|34|When the LORD heard what you said, he was angry and solemnly swore:
DEUT|1|35|"Not a man of this evil generation shall see the good land I swore to give your forefathers,
DEUT|1|36|except Caleb son of Jephunneh. He will see it, and I will give him and his descendants the land he set his feet on, because he followed the LORD wholeheartedly."
DEUT|1|37|Because of you the LORD became angry with me also and said, "You shall not enter it, either.
DEUT|1|38|But your assistant, Joshua son of Nun, will enter it. Encourage him, because he will lead Israel to inherit it.
DEUT|1|39|And the little ones that you said would be taken captive, your children who do not yet know good from bad-they will enter the land. I will give it to them and they will take possession of it.
DEUT|1|40|But as for you, turn around and set out toward the desert along the route to the Red Sea. "
DEUT|1|41|Then you replied, "We have sinned against the LORD. We will go up and fight, as the LORD our God commanded us." So every one of you put on his weapons, thinking it easy to go up into the hill country.
DEUT|1|42|But the LORD said to me, "Tell them, 'Do not go up and fight, because I will not be with you. You will be defeated by your enemies.'"
DEUT|1|43|So I told you, but you would not listen. You rebelled against the LORD's command and in your arrogance you marched up into the hill country.
DEUT|1|44|The Amorites who lived in those hills came out against you; they chased you like a swarm of bees and beat you down from Seir all the way to Hormah.
DEUT|1|45|You came back and wept before the LORD, but he paid no attention to your weeping and turned a deaf ear to you.
DEUT|1|46|And so you stayed in Kadesh many days-all the time you spent there.
DEUT|2|1|Then we turned back and set out toward the desert along the route to the Red Sea, as the LORD had directed me. For a long time we made our way around the hill country of Seir.
DEUT|2|2|Then the LORD said to me,
DEUT|2|3|"You have made your way around this hill country long enough; now turn north.
DEUT|2|4|Give the people these orders: 'You are about to pass through the territory of your brothers the descendants of Esau, who live in Seir. They will be afraid of you, but be very careful.
DEUT|2|5|Do not provoke them to war, for I will not give you any of their land, not even enough to put your foot on. I have given Esau the hill country of Seir as his own.
DEUT|2|6|You are to pay them in silver for the food you eat and the water you drink.'"
DEUT|2|7|The LORD your God has blessed you in all the work of your hands. He has watched over your journey through this vast desert. These forty years the LORD your God has been with you, and you have not lacked anything.
DEUT|2|8|So we went on past our brothers the descendants of Esau, who live in Seir. We turned from the Arabah road, which comes up from Elath and Ezion Geber, and traveled along the desert road of Moab.
DEUT|2|9|Then the LORD said to me, "Do not harass the Moabites or provoke them to war, for I will not give you any part of their land. I have given Ar to the descendants of Lot as a possession."
DEUT|2|10|(The Emites used to live there-a people strong and numerous, and as tall as the Anakites.
DEUT|2|11|Like the Anakites, they too were considered Rephaites, but the Moabites called them Emites.
DEUT|2|12|Horites used to live in Seir, but the descendants of Esau drove them out. They destroyed the Horites from before them and settled in their place, just as Israel did in the land the LORD gave them as their possession.)
DEUT|2|13|And the LORD said, "Now get up and cross the Zered Valley." So we crossed the valley.
DEUT|2|14|Thirty-eight years passed from the time we left Kadesh Barnea until we crossed the Zered Valley. By then, that entire generation of fighting men had perished from the camp, as the LORD had sworn to them.
DEUT|2|15|The LORD's hand was against them until he had completely eliminated them from the camp.
DEUT|2|16|Now when the last of these fighting men among the people had died,
DEUT|2|17|the LORD said to me,
DEUT|2|18|"Today you are to pass by the region of Moab at Ar.
DEUT|2|19|When you come to the Ammonites, do not harass them or provoke them to war, for I will not give you possession of any land belonging to the Ammonites. I have given it as a possession to the descendants of Lot."
DEUT|2|20|(That too was considered a land of the Rephaites, who used to live there; but the Ammonites called them Zamzummites.
DEUT|2|21|They were a people strong and numerous, and as tall as the Anakites. The LORD destroyed them from before the Ammonites, who drove them out and settled in their place.
DEUT|2|22|The LORD had done the same for the descendants of Esau, who lived in Seir, when he destroyed the Horites from before them. They drove them out and have lived in their place to this day.
DEUT|2|23|And as for the Avvites who lived in villages as far as Gaza, the Caphtorites coming out from Caphtor destroyed them and settled in their place.)
DEUT|2|24|"Set out now and cross the Arnon Gorge. See, I have given into your hand Sihon the Amorite, king of Heshbon, and his country. Begin to take possession of it and engage him in battle.
DEUT|2|25|This very day I will begin to put the terror and fear of you on all the nations under heaven. They will hear reports of you and will tremble and be in anguish because of you."
DEUT|2|26|From the desert of Kedemoth I sent messengers to Sihon king of Heshbon offering peace and saying,
DEUT|2|27|"Let us pass through your country. We will stay on the main road; we will not turn aside to the right or to the left.
DEUT|2|28|Sell us food to eat and water to drink for their price in silver. Only let us pass through on foot-
DEUT|2|29|as the descendants of Esau, who live in Seir, and the Moabites, who live in Ar, did for us-until we cross the Jordan into the land the LORD our God is giving us."
DEUT|2|30|But Sihon king of Heshbon refused to let us pass through. For the LORD your God had made his spirit stubborn and his heart obstinate in order to give him into your hands, as he has now done.
DEUT|2|31|The LORD said to me, "See, I have begun to deliver Sihon and his country over to you. Now begin to conquer and possess his land."
DEUT|2|32|When Sihon and all his army came out to meet us in battle at Jahaz,
DEUT|2|33|the LORD our God delivered him over to us and we struck him down, together with his sons and his whole army.
DEUT|2|34|At that time we took all his towns and completely destroyed them-men, women and children. We left no survivors.
DEUT|2|35|But the livestock and the plunder from the towns we had captured we carried off for ourselves.
DEUT|2|36|From Aroer on the rim of the Arnon Gorge, and from the town in the gorge, even as far as Gilead, not one town was too strong for us. The LORD our God gave us all of them.
DEUT|2|37|But in accordance with the command of the LORD our God, you did not encroach on any of the land of the Ammonites, neither the land along the course of the Jabbok nor that around the towns in the hills.
DEUT|3|1|Next we turned and went up along the road toward Bashan, and Og king of Bashan with his whole army marched out to meet us in battle at Edrei.
DEUT|3|2|The LORD said to me, "Do not be afraid of him, for I have handed him over to you with his whole army and his land. Do to him what you did to Sihon king of the Amorites, who reigned in Heshbon."
DEUT|3|3|So the LORD our God also gave into our hands Og king of Bashan and all his army. We struck them down, leaving no survivors.
DEUT|3|4|At that time we took all his cities. There was not one of the sixty cities that we did not take from them-the whole region of Argob, Og's kingdom in Bashan.
DEUT|3|5|All these cities were fortified with high walls and with gates and bars, and there were also a great many unwalled villages.
DEUT|3|6|We completely destroyed them, as we had done with Sihon king of Heshbon, destroying every city-men, women and children.
DEUT|3|7|But all the livestock and the plunder from their cities we carried off for ourselves.
DEUT|3|8|So at that time we took from these two kings of the Amorites the territory east of the Jordan, from the Arnon Gorge as far as Mount Hermon.
DEUT|3|9|(Hermon is called Sirion by the Sidonians; the Amorites call it Senir.)
DEUT|3|10|We took all the towns on the plateau, and all Gilead, and all Bashan as far as Salecah and Edrei, towns of Og's kingdom in Bashan.
DEUT|3|11|(Only Og king of Bashan was left of the remnant of the Rephaites. His bed was made of iron and was more than thirteen feet long and six feet wide. It is still in Rabbah of the Ammonites.)
DEUT|3|12|Of the land that we took over at that time, I gave the Reubenites and the Gadites the territory north of Aroer by the Arnon Gorge, including half the hill country of Gilead, together with its towns.
DEUT|3|13|The rest of Gilead and also all of Bashan, the kingdom of Og, I gave to the half tribe of Manasseh. (The whole region of Argob in Bashan used to be known as a land of the Rephaites.
DEUT|3|14|Jair, a descendant of Manasseh, took the whole region of Argob as far as the border of the Geshurites and the Maacathites; it was named after him, so that to this day Bashan is called Havvoth Jair. )
DEUT|3|15|And I gave Gilead to Makir.
DEUT|3|16|But to the Reubenites and the Gadites I gave the territory extending from Gilead down to the Arnon Gorge (the middle of the gorge being the border) and out to the Jabbok River, which is the border of the Ammonites.
DEUT|3|17|Its western border was the Jordan in the Arabah, from Kinnereth to the Sea of the Arabah (the Salt Sea ), below the slopes of Pisgah.
DEUT|3|18|I commanded you at that time: "The LORD your God has given you this land to take possession of it. But all your able-bodied men, armed for battle, must cross over ahead of your brother Israelites.
DEUT|3|19|However, your wives, your children and your livestock (I know you have much livestock) may stay in the towns I have given you,
DEUT|3|20|until the LORD gives rest to your brothers as he has to you, and they too have taken over the land that the LORD your God is giving them, across the Jordan. After that, each of you may go back to the possession I have given you."
DEUT|3|21|At that time I commanded Joshua: "You have seen with your own eyes all that the LORD your God has done to these two kings. The LORD will do the same to all the kingdoms over there where you are going.
DEUT|3|22|Do not be afraid of them; the LORD your God himself will fight for you."
DEUT|3|23|At that time I pleaded with the LORD:
DEUT|3|24|"O Sovereign LORD, you have begun to show to your servant your greatness and your strong hand. For what god is there in heaven or on earth who can do the deeds and mighty works you do?
DEUT|3|25|Let me go over and see the good land beyond the Jordan-that fine hill country and Lebanon."
DEUT|3|26|But because of you the LORD was angry with me and would not listen to me. "That is enough," the LORD said. "Do not speak to me anymore about this matter.
DEUT|3|27|Go up to the top of Pisgah and look west and north and south and east. Look at the land with your own eyes, since you are not going to cross this Jordan.
DEUT|3|28|But commission Joshua, and encourage and strengthen him, for he will lead this people across and will cause them to inherit the land that you will see."
DEUT|3|29|So we stayed in the valley near Beth Peor.
DEUT|4|1|Hear now, O Israel, the decrees and laws I am about to teach you. Follow them so that you may live and may go in and take possession of the land that the LORD, the God of your fathers, is giving you.
DEUT|4|2|Do not add to what I command you and do not subtract from it, but keep the commands of the LORD your God that I give you.
DEUT|4|3|You saw with your own eyes what the LORD did at Baal Peor. The LORD your God destroyed from among you everyone who followed the Baal of Peor,
DEUT|4|4|but all of you who held fast to the LORD your God are still alive today.
DEUT|4|5|See, I have taught you decrees and laws as the LORD my God commanded me, so that you may follow them in the land you are entering to take possession of it.
DEUT|4|6|Observe them carefully, for this will show your wisdom and understanding to the nations, who will hear about all these decrees and say, "Surely this great nation is a wise and understanding people."
DEUT|4|7|What other nation is so great as to have their gods near them the way the LORD our God is near us whenever we pray to him?
DEUT|4|8|And what other nation is so great as to have such righteous decrees and laws as this body of laws I am setting before you today?
DEUT|4|9|Only be careful, and watch yourselves closely so that you do not forget the things your eyes have seen or let them slip from your heart as long as you live. Teach them to your children and to their children after them.
DEUT|4|10|Remember the day you stood before the LORD your God at Horeb, when he said to me, "Assemble the people before me to hear my words so that they may learn to revere me as long as they live in the land and may teach them to their children."
DEUT|4|11|You came near and stood at the foot of the mountain while it blazed with fire to the very heavens, with black clouds and deep darkness.
DEUT|4|12|Then the LORD spoke to you out of the fire. You heard the sound of words but saw no form; there was only a voice.
DEUT|4|13|He declared to you his covenant, the Ten Commandments, which he commanded you to follow and then wrote them on two stone tablets.
DEUT|4|14|And the LORD directed me at that time to teach you the decrees and laws you are to follow in the land that you are crossing the Jordan to possess.
DEUT|4|15|You saw no form of any kind the day the LORD spoke to you at Horeb out of the fire. Therefore watch yourselves very carefully,
DEUT|4|16|so that you do not become corrupt and make for yourselves an idol, an image of any shape, whether formed like a man or a woman,
DEUT|4|17|or like any animal on earth or any bird that flies in the air,
DEUT|4|18|or like any creature that moves along the ground or any fish in the waters below.
DEUT|4|19|And when you look up to the sky and see the sun, the moon and the stars-all the heavenly array-do not be enticed into bowing down to them and worshiping things the LORD your God has apportioned to all the nations under heaven.
DEUT|4|20|But as for you, the LORD took you and brought you out of the iron-smelting furnace, out of Egypt, to be the people of his inheritance, as you now are.
DEUT|4|21|The LORD was angry with me because of you, and he solemnly swore that I would not cross the Jordan and enter the good land the LORD your God is giving you as your inheritance.
DEUT|4|22|I will die in this land; I will not cross the Jordan; but you are about to cross over and take possession of that good land.
DEUT|4|23|Be careful not to forget the covenant of the LORD your God that he made with you; do not make for yourselves an idol in the form of anything the LORD your God has forbidden.
DEUT|4|24|For the LORD your God is a consuming fire, a jealous God.
DEUT|4|25|After you have had children and grandchildren and have lived in the land a long time-if you then become corrupt and make any kind of idol, doing evil in the eyes of the LORD your God and provoking him to anger,
DEUT|4|26|I call heaven and earth as witnesses against you this day that you will quickly perish from the land that you are crossing the Jordan to possess. You will not live there long but will certainly be destroyed.
DEUT|4|27|The LORD will scatter you among the peoples, and only a few of you will survive among the nations to which the LORD will drive you.
DEUT|4|28|There you will worship man-made gods of wood and stone, which cannot see or hear or eat or smell.
DEUT|4|29|But if from there you seek the LORD your God, you will find him if you look for him with all your heart and with all your soul.
DEUT|4|30|When you are in distress and all these things have happened to you, then in later days you will return to the LORD your God and obey him.
DEUT|4|31|For the LORD your God is a merciful God; he will not abandon or destroy you or forget the covenant with your forefathers, which he confirmed to them by oath.
DEUT|4|32|Ask now about the former days, long before your time, from the day God created man on the earth; ask from one end of the heavens to the other. Has anything so great as this ever happened, or has anything like it ever been heard of?
DEUT|4|33|Has any other people heard the voice of God speaking out of fire, as you have, and lived?
DEUT|4|34|Has any god ever tried to take for himself one nation out of another nation, by testings, by miraculous signs and wonders, by war, by a mighty hand and an outstretched arm, or by great and awesome deeds, like all the things the LORD your God did for you in Egypt before your very eyes?
DEUT|4|35|You were shown these things so that you might know that the LORD is God; besides him there is no other.
DEUT|4|36|From heaven he made you hear his voice to discipline you. On earth he showed you his great fire, and you heard his words from out of the fire.
DEUT|4|37|Because he loved your forefathers and chose their descendants after them, he brought you out of Egypt by his Presence and his great strength,
DEUT|4|38|to drive out before you nations greater and stronger than you and to bring you into their land to give it to you for your inheritance, as it is today.
DEUT|4|39|Acknowledge and take to heart this day that the LORD is God in heaven above and on the earth below. There is no other.
DEUT|4|40|Keep his decrees and commands, which I am giving you today, so that it may go well with you and your children after you and that you may live long in the land the LORD your God gives you for all time.
DEUT|4|41|Then Moses set aside three cities east of the Jordan,
DEUT|4|42|to which anyone who had killed a person could flee if he had unintentionally killed his neighbor without malice aforethought. He could flee into one of these cities and save his life.
DEUT|4|43|The cities were these: Bezer in the desert plateau, for the Reubenites; Ramoth in Gilead, for the Gadites; and Golan in Bashan, for the Manassites.
DEUT|4|44|This is the law Moses set before the Israelites.
DEUT|4|45|These are the stipulations, decrees and laws Moses gave them when they came out of Egypt
DEUT|4|46|and were in the valley near Beth Peor east of the Jordan, in the land of Sihon king of the Amorites, who reigned in Heshbon and was defeated by Moses and the Israelites as they came out of Egypt.
DEUT|4|47|They took possession of his land and the land of Og king of Bashan, the two Amorite kings east of the Jordan.
DEUT|4|48|This land extended from Aroer on the rim of the Arnon Gorge to Mount Siyon (that is, Hermon),
DEUT|4|49|and included all the Arabah east of the Jordan, as far as the Sea of the Arabah, below the slopes of Pisgah.
DEUT|5|1|Moses summoned all Israel and said: Hear, O Israel, the decrees and laws I declare in your hearing today. Learn them and be sure to follow them.
DEUT|5|2|The LORD our God made a covenant with us at Horeb.
DEUT|5|3|It was not with our fathers that the LORD made this covenant, but with us, with all of us who are alive here today.
DEUT|5|4|The LORD spoke to you face to face out of the fire on the mountain.
DEUT|5|5|(At that time I stood between the LORD and you to declare to you the word of the LORD, because you were afraid of the fire and did not go up the mountain.) And he said:
DEUT|5|6|"I am the LORD your God, who brought you out of Egypt, out of the land of slavery.
DEUT|5|7|"You shall have no other gods before me.
DEUT|5|8|"You shall not make for yourself an idol in the form of anything in heaven above or on the earth beneath or in the waters below.
DEUT|5|9|You shall not bow down to them or worship them; for I, the LORD your God, am a jealous God, punishing the children for the sin of the fathers to the third and fourth generation of those who hate me,
DEUT|5|10|but showing love to a thousand generations of those who love me and keep my commandments.
DEUT|5|11|"You shall not misuse the name of the LORD your God, for the LORD will not hold anyone guiltless who misuses his name.
DEUT|5|12|"Observe the Sabbath day by keeping it holy, as the LORD your God has commanded you.
DEUT|5|13|Six days you shall labor and do all your work,
DEUT|5|14|but the seventh day is a Sabbath to the LORD your God. On it you shall not do any work, neither you, nor your son or daughter, nor your manservant or maidservant, nor your ox, your donkey or any of your animals, nor the alien within your gates, so that your manservant and maidservant may rest, as you do.
DEUT|5|15|Remember that you were slaves in Egypt and that the LORD your God brought you out of there with a mighty hand and an outstretched arm. Therefore the LORD your God has commanded you to observe the Sabbath day.
DEUT|5|16|"Honor your father and your mother, as the LORD your God has commanded you, so that you may live long and that it may go well with you in the land the LORD your God is giving you.
DEUT|5|17|"You shall not murder.
DEUT|5|18|"You shall not commit adultery.
DEUT|5|19|"You shall not steal.
DEUT|5|20|"You shall not give false testimony against your neighbor.
DEUT|5|21|"You shall not covet your neighbor's wife. You shall not set your desire on your neighbor's house or land, his manservant or maidservant, his ox or donkey, or anything that belongs to your neighbor."
DEUT|5|22|These are the commandments the LORD proclaimed in a loud voice to your whole assembly there on the mountain from out of the fire, the cloud and the deep darkness; and he added nothing more. Then he wrote them on two stone tablets and gave them to me.
DEUT|5|23|When you heard the voice out of the darkness, while the mountain was ablaze with fire, all the leading men of your tribes and your elders came to me.
DEUT|5|24|And you said, "The LORD our God has shown us his glory and his majesty, and we have heard his voice from the fire. Today we have seen that a man can live even if God speaks with him.
DEUT|5|25|But now, why should we die? This great fire will consume us, and we will die if we hear the voice of the LORD our God any longer.
DEUT|5|26|For what mortal man has ever heard the voice of the living God speaking out of fire, as we have, and survived?
DEUT|5|27|Go near and listen to all that the LORD our God says. Then tell us whatever the LORD our God tells you. We will listen and obey."
DEUT|5|28|The LORD heard you when you spoke to me and the LORD said to me, "I have heard what this people said to you. Everything they said was good.
DEUT|5|29|Oh, that their hearts would be inclined to fear me and keep all my commands always, so that it might go well with them and their children forever!
DEUT|5|30|"Go, tell them to return to their tents.
DEUT|5|31|But you stay here with me so that I may give you all the commands, decrees and laws you are to teach them to follow in the land I am giving them to possess."
DEUT|5|32|So be careful to do what the LORD your God has commanded you; do not turn aside to the right or to the left.
DEUT|5|33|Walk in all the way that the LORD your God has commanded you, so that you may live and prosper and prolong your days in the land that you will possess.
DEUT|6|1|These are the commands, decrees and laws the LORD your God directed me to teach you to observe in the land that you are crossing the Jordan to possess,
DEUT|6|2|so that you, your children and their children after them may fear the LORD your God as long as you live by keeping all his decrees and commands that I give you, and so that you may enjoy long life.
DEUT|6|3|Hear, O Israel, and be careful to obey so that it may go well with you and that you may increase greatly in a land flowing with milk and honey, just as the LORD, the God of your fathers, promised you.
DEUT|6|4|Hear, O Israel: The LORD our God, the LORD is one.
DEUT|6|5|Love the LORD your God with all your heart and with all your soul and with all your strength.
DEUT|6|6|These commandments that I give you today are to be upon your hearts.
DEUT|6|7|Impress them on your children. Talk about them when you sit at home and when you walk along the road, when you lie down and when you get up.
DEUT|6|8|Tie them as symbols on your hands and bind them on your foreheads.
DEUT|6|9|Write them on the doorframes of your houses and on your gates.
DEUT|6|10|When the LORD your God brings you into the land he swore to your fathers, to Abraham, Isaac and Jacob, to give you-a land with large, flourishing cities you did not build,
DEUT|6|11|houses filled with all kinds of good things you did not provide, wells you did not dig, and vineyards and olive groves you did not plant-then when you eat and are satisfied,
DEUT|6|12|be careful that you do not forget the LORD, who brought you out of Egypt, out of the land of slavery.
DEUT|6|13|Fear the LORD your God, serve him only and take your oaths in his name.
DEUT|6|14|Do not follow other gods, the gods of the peoples around you;
DEUT|6|15|for the LORD your God, who is among you, is a jealous God and his anger will burn against you, and he will destroy you from the face of the land.
DEUT|6|16|Do not test the LORD your God as you did at Massah.
DEUT|6|17|Be sure to keep the commands of the LORD your God and the stipulations and decrees he has given you.
DEUT|6|18|Do what is right and good in the LORD's sight, so that it may go well with you and you may go in and take over the good land that the LORD promised on oath to your forefathers,
DEUT|6|19|thrusting out all your enemies before you, as the LORD said.
DEUT|6|20|In the future, when your son asks you, "What is the meaning of the stipulations, decrees and laws the LORD our God has commanded you?"
DEUT|6|21|tell him: "We were slaves of Pharaoh in Egypt, but the LORD brought us out of Egypt with a mighty hand.
DEUT|6|22|Before our eyes the LORD sent miraculous signs and wonders-great and terrible-upon Egypt and Pharaoh and his whole household.
DEUT|6|23|But he brought us out from there to bring us in and give us the land that he promised on oath to our forefathers.
DEUT|6|24|The LORD commanded us to obey all these decrees and to fear the LORD our God, so that we might always prosper and be kept alive, as is the case today.
DEUT|6|25|And if we are careful to obey all this law before the LORD our God, as he has commanded us, that will be our righteousness."
DEUT|7|1|When the LORD your God brings you into the land you are entering to possess and drives out before you many nations-the Hittites, Girgashites, Amorites, Canaanites, Perizzites, Hivites and Jebusites, seven nations larger and stronger than you-
DEUT|7|2|and when the LORD your God has delivered them over to you and you have defeated them, then you must destroy them totally. Make no treaty with them, and show them no mercy.
DEUT|7|3|Do not intermarry with them. Do not give your daughters to their sons or take their daughters for your sons,
DEUT|7|4|for they will turn your sons away from following me to serve other gods, and the LORD's anger will burn against you and will quickly destroy you.
DEUT|7|5|This is what you are to do to them: Break down their altars, smash their sacred stones, cut down their Asherah poles and burn their idols in the fire.
DEUT|7|6|For you are a people holy to the LORD your God. The LORD your God has chosen you out of all the peoples on the face of the earth to be his people, his treasured possession.
DEUT|7|7|The LORD did not set his affection on you and choose you because you were more numerous than other peoples, for you were the fewest of all peoples.
DEUT|7|8|But it was because the LORD loved you and kept the oath he swore to your forefathers that he brought you out with a mighty hand and redeemed you from the land of slavery, from the power of Pharaoh king of Egypt.
DEUT|7|9|Know therefore that the LORD your God is God; he is the faithful God, keeping his covenant of love to a thousand generations of those who love him and keep his commands.
DEUT|7|10|But those who hate him he will repay to their face by destruction; he will not be slow to repay to their face those who hate him.
DEUT|7|11|Therefore, take care to follow the commands, decrees and laws I give you today.
DEUT|7|12|If you pay attention to these laws and are careful to follow them, then the LORD your God will keep his covenant of love with you, as he swore to your forefathers.
DEUT|7|13|He will love you and bless you and increase your numbers. He will bless the fruit of your womb, the crops of your land-your grain, new wine and oil-the calves of your herds and the lambs of your flocks in the land that he swore to your forefathers to give you.
DEUT|7|14|You will be blessed more than any other people; none of your men or women will be childless, nor any of your livestock without young.
DEUT|7|15|The LORD will keep you free from every disease. He will not inflict on you the horrible diseases you knew in Egypt, but he will inflict them on all who hate you.
DEUT|7|16|You must destroy all the peoples the LORD your God gives over to you. Do not look on them with pity and do not serve their gods, for that will be a snare to you.
DEUT|7|17|You may say to yourselves, "These nations are stronger than we are. How can we drive them out?"
DEUT|7|18|But do not be afraid of them; remember well what the LORD your God did to Pharaoh and to all Egypt.
DEUT|7|19|You saw with your own eyes the great trials, the miraculous signs and wonders, the mighty hand and outstretched arm, with which the LORD your God brought you out. The LORD your God will do the same to all the peoples you now fear.
DEUT|7|20|Moreover, the LORD your God will send the hornet among them until even the survivors who hide from you have perished.
DEUT|7|21|Do not be terrified by them, for the LORD your God, who is among you, is a great and awesome God.
DEUT|7|22|The LORD your God will drive out those nations before you, little by little. You will not be allowed to eliminate them all at once, or the wild animals will multiply around you.
DEUT|7|23|But the LORD your God will deliver them over to you, throwing them into great confusion until they are destroyed.
DEUT|7|24|He will give their kings into your hand, and you will wipe out their names from under heaven. No one will be able to stand up against you; you will destroy them.
DEUT|7|25|The images of their gods you are to burn in the fire. Do not covet the silver and gold on them, and do not take it for yourselves, or you will be ensnared by it, for it is detestable to the LORD your God.
DEUT|7|26|Do not bring a detestable thing into your house or you, like it, will be set apart for destruction. Utterly abhor and detest it, for it is set apart for destruction.
DEUT|8|1|Be careful to follow every command I am giving you today, so that you may live and increase and may enter and possess the land that the LORD promised on oath to your forefathers.
DEUT|8|2|Remember how the LORD your God led you all the way in the desert these forty years, to humble you and to test you in order to know what was in your heart, whether or not you would keep his commands.
DEUT|8|3|He humbled you, causing you to hunger and then feeding you with manna, which neither you nor your fathers had known, to teach you that man does not live on bread alone but on every word that comes from the mouth of the LORD.
DEUT|8|4|Your clothes did not wear out and your feet did not swell during these forty years.
DEUT|8|5|Know then in your heart that as a man disciplines his son, so the LORD your God disciplines you.
DEUT|8|6|Observe the commands of the LORD your God, walking in his ways and revering him.
DEUT|8|7|For the LORD your God is bringing you into a good land-a land with streams and pools of water, with springs flowing in the valleys and hills;
DEUT|8|8|a land with wheat and barley, vines and fig trees, pomegranates, olive oil and honey;
DEUT|8|9|a land where bread will not be scarce and you will lack nothing; a land where the rocks are iron and you can dig copper out of the hills.
DEUT|8|10|When you have eaten and are satisfied, praise the LORD your God for the good land he has given you.
DEUT|8|11|Be careful that you do not forget the LORD your God, failing to observe his commands, his laws and his decrees that I am giving you this day.
DEUT|8|12|Otherwise, when you eat and are satisfied, when you build fine houses and settle down,
DEUT|8|13|and when your herds and flocks grow large and your silver and gold increase and all you have is multiplied,
DEUT|8|14|then your heart will become proud and you will forget the LORD your God, who brought you out of Egypt, out of the land of slavery.
DEUT|8|15|He led you through the vast and dreadful desert, that thirsty and waterless land, with its venomous snakes and scorpions. He brought you water out of hard rock.
DEUT|8|16|He gave you manna to eat in the desert, something your fathers had never known, to humble and to test you so that in the end it might go well with you.
DEUT|8|17|You may say to yourself, "My power and the strength of my hands have produced this wealth for me."
DEUT|8|18|But remember the LORD your God, for it is he who gives you the ability to produce wealth, and so confirms his covenant, which he swore to your forefathers, as it is today.
DEUT|8|19|If you ever forget the LORD your God and follow other gods and worship and bow down to them, I testify against you today that you will surely be destroyed.
DEUT|8|20|Like the nations the LORD destroyed before you, so you will be destroyed for not obeying the LORD your God.
DEUT|9|1|Hear, O Israel. You are now about to cross the Jordan to go in and dispossess nations greater and stronger than you, with large cities that have walls up to the sky.
DEUT|9|2|The people are strong and tall-Anakites! You know about them and have heard it said: "Who can stand up against the Anakites?"
DEUT|9|3|But be assured today that the LORD your God is the one who goes across ahead of you like a devouring fire. He will destroy them; he will subdue them before you. And you will drive them out and annihilate them quickly, as the LORD has promised you.
DEUT|9|4|After the LORD your God has driven them out before you, do not say to yourself, "The LORD has brought me here to take possession of this land because of my righteousness." No, it is on account of the wickedness of these nations that the LORD is going to drive them out before you.
DEUT|9|5|It is not because of your righteousness or your integrity that you are going in to take possession of their land; but on account of the wickedness of these nations, the LORD your God will drive them out before you, to accomplish what he swore to your fathers, to Abraham, Isaac and Jacob.
DEUT|9|6|Understand, then, that it is not because of your righteousness that the LORD your God is giving you this good land to possess, for you are a stiff-necked people.
DEUT|9|7|Remember this and never forget how you provoked the LORD your God to anger in the desert. From the day you left Egypt until you arrived here, you have been rebellious against the LORD.
DEUT|9|8|At Horeb you aroused the LORD's wrath so that he was angry enough to destroy you.
DEUT|9|9|When I went up on the mountain to receive the tablets of stone, the tablets of the covenant that the LORD had made with you, I stayed on the mountain forty days and forty nights; I ate no bread and drank no water.
DEUT|9|10|The LORD gave me two stone tablets inscribed by the finger of God. On them were all the commandments the LORD proclaimed to you on the mountain out of the fire, on the day of the assembly.
DEUT|9|11|At the end of the forty days and forty nights, the LORD gave me the two stone tablets, the tablets of the covenant.
DEUT|9|12|Then the LORD told me, "Go down from here at once, because your people whom you brought out of Egypt have become corrupt. They have turned away quickly from what I commanded them and have made a cast idol for themselves."
DEUT|9|13|And the LORD said to me, "I have seen this people, and they are a stiff-necked people indeed!
DEUT|9|14|Let me alone, so that I may destroy them and blot out their name from under heaven. And I will make you into a nation stronger and more numerous than they."
DEUT|9|15|So I turned and went down from the mountain while it was ablaze with fire. And the two tablets of the covenant were in my hands.
DEUT|9|16|When I looked, I saw that you had sinned against the LORD your God; you had made for yourselves an idol cast in the shape of a calf. You had turned aside quickly from the way that the LORD had commanded you.
DEUT|9|17|So I took the two tablets and threw them out of my hands, breaking them to pieces before your eyes.
DEUT|9|18|Then once again I fell prostrate before the LORD for forty days and forty nights; I ate no bread and drank no water, because of all the sin you had committed, doing what was evil in the LORD's sight and so provoking him to anger.
DEUT|9|19|I feared the anger and wrath of the LORD, for he was angry enough with you to destroy you. But again the LORD listened to me.
DEUT|9|20|And the LORD was angry enough with Aaron to destroy him, but at that time I prayed for Aaron too.
DEUT|9|21|Also I took that sinful thing of yours, the calf you had made, and burned it in the fire. Then I crushed it and ground it to powder as fine as dust and threw the dust into a stream that flowed down the mountain.
DEUT|9|22|You also made the LORD angry at Taberah, at Massah and at Kibroth Hattaavah.
DEUT|9|23|And when the LORD sent you out from Kadesh Barnea, he said, "Go up and take possession of the land I have given you." But you rebelled against the command of the LORD your God. You did not trust him or obey him.
DEUT|9|24|You have been rebellious against the LORD ever since I have known you.
DEUT|9|25|I lay prostrate before the LORD those forty days and forty nights because the LORD had said he would destroy you.
DEUT|9|26|I prayed to the LORD and said, "O Sovereign LORD, do not destroy your people, your own inheritance that you redeemed by your great power and brought out of Egypt with a mighty hand.
DEUT|9|27|Remember your servants Abraham, Isaac and Jacob. Overlook the stubbornness of this people, their wickedness and their sin.
DEUT|9|28|Otherwise, the country from which you brought us will say, 'Because the LORD was not able to take them into the land he had promised them, and because he hated them, he brought them out to put them to death in the desert.'
DEUT|9|29|But they are your people, your inheritance that you brought out by your great power and your outstretched arm."
DEUT|10|1|At that time the LORD said to me, "Chisel out two stone tablets like the first ones and come up to me on the mountain. Also make a wooden chest.
DEUT|10|2|I will write on the tablets the words that were on the first tablets, which you broke. Then you are to put them in the chest."
DEUT|10|3|So I made the ark out of acacia wood and chiseled out two stone tablets like the first ones, and I went up on the mountain with the two tablets in my hands.
DEUT|10|4|The LORD wrote on these tablets what he had written before, the Ten Commandments he had proclaimed to you on the mountain, out of the fire, on the day of the assembly. And the LORD gave them to me.
DEUT|10|5|Then I came back down the mountain and put the tablets in the ark I had made, as the LORD commanded me, and they are there now.
DEUT|10|6|(The Israelites traveled from the wells of the Jaakanites to Moserah. There Aaron died and was buried, and Eleazar his son succeeded him as priest.
DEUT|10|7|From there they traveled to Gudgodah and on to Jotbathah, a land with streams of water.
DEUT|10|8|At that time the LORD set apart the tribe of Levi to carry the ark of the covenant of the LORD, to stand before the LORD to minister and to pronounce blessings in his name, as they still do today.
DEUT|10|9|That is why the Levites have no share or inheritance among their brothers; the LORD is their inheritance, as the LORD your God told them.)
DEUT|10|10|Now I had stayed on the mountain forty days and nights, as I did the first time, and the LORD listened to me at this time also. It was not his will to destroy you.
DEUT|10|11|"Go," the LORD said to me, "and lead the people on their way, so that they may enter and possess the land that I swore to their fathers to give them."
DEUT|10|12|And now, O Israel, what does the LORD your God ask of you but to fear the LORD your God, to walk in all his ways, to love him, to serve the LORD your God with all your heart and with all your soul,
DEUT|10|13|and to observe the LORD's commands and decrees that I am giving you today for your own good?
DEUT|10|14|To the LORD your God belong the heavens, even the highest heavens, the earth and everything in it.
DEUT|10|15|Yet the LORD set his affection on your forefathers and loved them, and he chose you, their descendants, above all the nations, as it is today.
DEUT|10|16|Circumcise your hearts, therefore, and do not be stiff-necked any longer.
DEUT|10|17|For the LORD your God is God of gods and Lord of lords, the great God, mighty and awesome, who shows no partiality and accepts no bribes.
DEUT|10|18|He defends the cause of the fatherless and the widow, and loves the alien, giving him food and clothing.
DEUT|10|19|And you are to love those who are aliens, for you yourselves were aliens in Egypt.
DEUT|10|20|Fear the LORD your God and serve him. Hold fast to him and take your oaths in his name.
DEUT|10|21|He is your praise; he is your God, who performed for you those great and awesome wonders you saw with your own eyes.
DEUT|10|22|Your forefathers who went down into Egypt were seventy in all, and now the LORD your God has made you as numerous as the stars in the sky.
DEUT|11|1|Love the LORD your God and keep his requirements, his decrees, his laws and his commands always.
DEUT|11|2|Remember today that your children were not the ones who saw and experienced the discipline of the LORD your God: his majesty, his mighty hand, his outstretched arm;
DEUT|11|3|the signs he performed and the things he did in the heart of Egypt, both to Pharaoh king of Egypt and to his whole country;
DEUT|11|4|what he did to the Egyptian army, to its horses and chariots, how he overwhelmed them with the waters of the Red Sea as they were pursuing you, and how the LORD brought lasting ruin on them.
DEUT|11|5|It was not your children who saw what he did for you in the desert until you arrived at this place,
DEUT|11|6|and what he did to Dathan and Abiram, sons of Eliab the Reubenite, when the earth opened its mouth right in the middle of all Israel and swallowed them up with their households, their tents and every living thing that belonged to them.
DEUT|11|7|But it was your own eyes that saw all these great things the LORD has done.
DEUT|11|8|Observe therefore all the commands I am giving you today, so that you may have the strength to go in and take over the land that you are crossing the Jordan to possess,
DEUT|11|9|and so that you may live long in the land that the LORD swore to your forefathers to give to them and their descendants, a land flowing with milk and honey.
DEUT|11|10|The land you are entering to take over is not like the land of Egypt, from which you have come, where you planted your seed and irrigated it by foot as in a vegetable garden.
DEUT|11|11|But the land you are crossing the Jordan to take possession of is a land of mountains and valleys that drinks rain from heaven.
DEUT|11|12|It is a land the LORD your God cares for; the eyes of the LORD your God are continually on it from the beginning of the year to its end.
DEUT|11|13|So if you faithfully obey the commands I am giving you today-to love the LORD your God and to serve him with all your heart and with all your soul-
DEUT|11|14|then I will send rain on your land in its season, both autumn and spring rains, so that you may gather in your grain, new wine and oil.
DEUT|11|15|I will provide grass in the fields for your cattle, and you will eat and be satisfied.
DEUT|11|16|Be careful, or you will be enticed to turn away and worship other gods and bow down to them.
DEUT|11|17|Then the LORD's anger will burn against you, and he will shut the heavens so that it will not rain and the ground will yield no produce, and you will soon perish from the good land the LORD is giving you.
DEUT|11|18|Fix these words of mine in your hearts and minds; tie them as symbols on your hands and bind them on your foreheads.
DEUT|11|19|Teach them to your children, talking about them when you sit at home and when you walk along the road, when you lie down and when you get up.
DEUT|11|20|Write them on the doorframes of your houses and on your gates,
DEUT|11|21|so that your days and the days of your children may be many in the land that the LORD swore to give your forefathers, as many as the days that the heavens are above the earth.
DEUT|11|22|If you carefully observe all these commands I am giving you to follow-to love the LORD your God, to walk in all his ways and to hold fast to him-
DEUT|11|23|then the LORD will drive out all these nations before you, and you will dispossess nations larger and stronger than you.
DEUT|11|24|Every place where you set your foot will be yours: Your territory will extend from the desert to Lebanon, and from the Euphrates River to the western sea.
DEUT|11|25|No man will be able to stand against you. The LORD your God, as he promised you, will put the terror and fear of you on the whole land, wherever you go.
DEUT|11|26|See, I am setting before you today a blessing and a curse-
DEUT|11|27|the blessing if you obey the commands of the LORD your God that I am giving you today;
DEUT|11|28|the curse if you disobey the commands of the LORD your God and turn from the way that I command you today by following other gods, which you have not known.
DEUT|11|29|When the LORD your God has brought you into the land you are entering to possess, you are to proclaim on Mount Gerizim the blessings, and on Mount Ebal the curses.
DEUT|11|30|As you know, these mountains are across the Jordan, west of the road, toward the setting sun, near the great trees of Moreh, in the territory of those Canaanites living in the Arabah in the vicinity of Gilgal.
DEUT|11|31|You are about to cross the Jordan to enter and take possession of the land the LORD your God is giving you. When you have taken it over and are living there,
DEUT|11|32|be sure that you obey all the decrees and laws I am setting before you today.
DEUT|12|1|These are the decrees and laws you must be careful to follow in the land that the LORD, the God of your fathers, has given you to possess-as long as you live in the land.
DEUT|12|2|Destroy completely all the places on the high mountains and on the hills and under every spreading tree where the nations you are dispossessing worship their gods.
DEUT|12|3|Break down their altars, smash their sacred stones and burn their Asherah poles in the fire; cut down the idols of their gods and wipe out their names from those places.
DEUT|12|4|You must not worship the LORD your God in their way.
DEUT|12|5|But you are to seek the place the LORD your God will choose from among all your tribes to put his Name there for his dwelling. To that place you must go;
DEUT|12|6|there bring your burnt offerings and sacrifices, your tithes and special gifts, what you have vowed to give and your freewill offerings, and the firstborn of your herds and flocks.
DEUT|12|7|There, in the presence of the LORD your God, you and your families shall eat and shall rejoice in everything you have put your hand to, because the LORD your God has blessed you.
DEUT|12|8|You are not to do as we do here today, everyone as he sees fit,
DEUT|12|9|since you have not yet reached the resting place and the inheritance the LORD your God is giving you.
DEUT|12|10|But you will cross the Jordan and settle in the land the LORD your God is giving you as an inheritance, and he will give you rest from all your enemies around you so that you will live in safety.
DEUT|12|11|Then to the place the LORD your God will choose as a dwelling for his Name-there you are to bring everything I command you: your burnt offerings and sacrifices, your tithes and special gifts, and all the choice possessions you have vowed to the LORD.
DEUT|12|12|And there rejoice before the LORD your God, you, your sons and daughters, your menservants and maidservants, and the Levites from your towns, who have no allotment or inheritance of their own.
DEUT|12|13|Be careful not to sacrifice your burnt offerings anywhere you please.
DEUT|12|14|Offer them only at the place the LORD will choose in one of your tribes, and there observe everything I command you.
DEUT|12|15|Nevertheless, you may slaughter your animals in any of your towns and eat as much of the meat as you want, as if it were gazelle or deer, according to the blessing the LORD your God gives you. Both the ceremonially unclean and the clean may eat it.
DEUT|12|16|But you must not eat the blood; pour it out on the ground like water.
DEUT|12|17|You must not eat in your own towns the tithe of your grain and new wine and oil, or the firstborn of your herds and flocks, or whatever you have vowed to give, or your freewill offerings or special gifts.
DEUT|12|18|Instead, you are to eat them in the presence of the LORD your God at the place the LORD your God will choose-you, your sons and daughters, your menservants and maidservants, and the Levites from your towns-and you are to rejoice before the LORD your God in everything you put your hand to.
DEUT|12|19|Be careful not to neglect the Levites as long as you live in your land.
DEUT|12|20|When the LORD your God has enlarged your territory as he promised you, and you crave meat and say, "I would like some meat," then you may eat as much of it as you want.
DEUT|12|21|If the place where the LORD your God chooses to put his Name is too far away from you, you may slaughter animals from the herds and flocks the LORD has given you, as I have commanded you, and in your own towns you may eat as much of them as you want.
DEUT|12|22|Eat them as you would gazelle or deer. Both the ceremonially unclean and the clean may eat.
DEUT|12|23|But be sure you do not eat the blood, because the blood is the life, and you must not eat the life with the meat.
DEUT|12|24|You must not eat the blood; pour it out on the ground like water.
DEUT|12|25|Do not eat it, so that it may go well with you and your children after you, because you will be doing what is right in the eyes of the LORD.
DEUT|12|26|But take your consecrated things and whatever you have vowed to give, and go to the place the LORD will choose.
DEUT|12|27|Present your burnt offerings on the altar of the LORD your God, both the meat and the blood. The blood of your sacrifices must be poured beside the altar of the LORD your God, but you may eat the meat.
DEUT|12|28|Be careful to obey all these regulations I am giving you, so that it may always go well with you and your children after you, because you will be doing what is good and right in the eyes of the LORD your God.
DEUT|12|29|The LORD your God will cut off before you the nations you are about to invade and dispossess. But when you have driven them out and settled in their land,
DEUT|12|30|and after they have been destroyed before you, be careful not to be ensnared by inquiring about their gods, saying, "How do these nations serve their gods? We will do the same."
DEUT|12|31|You must not worship the LORD your God in their way, because in worshiping their gods, they do all kinds of detestable things the LORD hates. They even burn their sons and daughters in the fire as sacrifices to their gods.
DEUT|12|32|See that you do all I command you; do not add to it or take away from it.
DEUT|13|1|If a prophet, or one who foretells by dreams, appears among you and announces to you a miraculous sign or wonder,
DEUT|13|2|and if the sign or wonder of which he has spoken takes place, and he says, "Let us follow other gods" (gods you have not known) "and let us worship them,"
DEUT|13|3|you must not listen to the words of that prophet or dreamer. The LORD your God is testing you to find out whether you love him with all your heart and with all your soul.
DEUT|13|4|It is the LORD your God you must follow, and him you must revere. Keep his commands and obey him; serve him and hold fast to him.
DEUT|13|5|That prophet or dreamer must be put to death, because he preached rebellion against the LORD your God, who brought you out of Egypt and redeemed you from the land of slavery; he has tried to turn you from the way the LORD your God commanded you to follow. You must purge the evil from among you.
DEUT|13|6|If your very own brother, or your son or daughter, or the wife you love, or your closest friend secretly entices you, saying, "Let us go and worship other gods" (gods that neither you nor your fathers have known,
DEUT|13|7|gods of the peoples around you, whether near or far, from one end of the land to the other),
DEUT|13|8|do not yield to him or listen to him. Show him no pity. Do not spare him or shield him.
DEUT|13|9|You must certainly put him to death. Your hand must be the first in putting him to death, and then the hands of all the people.
DEUT|13|10|Stone him to death, because he tried to turn you away from the LORD your God, who brought you out of Egypt, out of the land of slavery.
DEUT|13|11|Then all Israel will hear and be afraid, and no one among you will do such an evil thing again.
DEUT|13|12|If you hear it said about one of the towns the LORD your God is giving you to live in
DEUT|13|13|that wicked men have arisen among you and have led the people of their town astray, saying, "Let us go and worship other gods" (gods you have not known),
DEUT|13|14|then you must inquire, probe and investigate it thoroughly. And if it is true and it has been proved that this detestable thing has been done among you,
DEUT|13|15|you must certainly put to the sword all who live in that town. Destroy it completely, both its people and its livestock.
DEUT|13|16|Gather all the plunder of the town into the middle of the public square and completely burn the town and all its plunder as a whole burnt offering to the LORD your God. It is to remain a ruin forever, never to be rebuilt.
DEUT|13|17|None of those condemned things shall be found in your hands, so that the LORD will turn from his fierce anger; he will show you mercy, have compassion on you, and increase your numbers, as he promised on oath to your forefathers,
DEUT|13|18|because you obey the LORD your God, keeping all his commands that I am giving you today and doing what is right in his eyes.
DEUT|14|1|You are the children of the LORD your God. Do not cut yourselves or shave the front of your heads for the dead,
DEUT|14|2|for you are a people holy to the LORD your God. Out of all the peoples on the face of the earth, the LORD has chosen you to be his treasured possession.
DEUT|14|3|Do not eat any detestable thing.
DEUT|14|4|These are the animals you may eat: the ox, the sheep, the goat,
DEUT|14|5|the deer, the gazelle, the roe deer, the wild goat, the ibex, the antelope and the mountain sheep.
DEUT|14|6|You may eat any animal that has a split hoof divided in two and that chews the cud.
DEUT|14|7|However, of those that chew the cud or that have a split hoof completely divided you may not eat the camel, the rabbit or the coney. Although they chew the cud, they do not have a split hoof; they are ceremonially unclean for you.
DEUT|14|8|The pig is also unclean; although it has a split hoof, it does not chew the cud. You are not to eat their meat or touch their carcasses.
DEUT|14|9|Of all the creatures living in the water, you may eat any that has fins and scales.
DEUT|14|10|But anything that does not have fins and scales you may not eat; for you it is unclean.
DEUT|14|11|You may eat any clean bird.
DEUT|14|12|But these you may not eat: the eagle, the vulture, the black vulture,
DEUT|14|13|the red kite, the black kite, any kind of falcon,
DEUT|14|14|any kind of raven,
DEUT|14|15|the horned owl, the screech owl, the gull, any kind of hawk,
DEUT|14|16|the little owl, the great owl, the white owl,
DEUT|14|17|the desert owl, the osprey, the cormorant,
DEUT|14|18|the stork, any kind of heron, the hoopoe and the bat.
DEUT|14|19|All flying insects that swarm are unclean to you; do not eat them.
DEUT|14|20|But any winged creature that is clean you may eat.
DEUT|14|21|Do not eat anything you find already dead. You may give it to an alien living in any of your towns, and he may eat it, or you may sell it to a foreigner. But you are a people holy to the LORD your God. Do not cook a young goat in its mother's milk.
DEUT|14|22|Be sure to set aside a tenth of all that your fields produce each year.
DEUT|14|23|Eat the tithe of your grain, new wine and oil, and the firstborn of your herds and flocks in the presence of the LORD your God at the place he will choose as a dwelling for his Name, so that you may learn to revere the LORD your God always.
DEUT|14|24|But if that place is too distant and you have been blessed by the LORD your God and cannot carry your tithe (because the place where the LORD will choose to put his Name is so far away),
DEUT|14|25|then exchange your tithe for silver, and take the silver with you and go to the place the LORD your God will choose.
DEUT|14|26|Use the silver to buy whatever you like: cattle, sheep, wine or other fermented drink, or anything you wish. Then you and your household shall eat there in the presence of the LORD your God and rejoice.
DEUT|14|27|And do not neglect the Levites living in your towns, for they have no allotment or inheritance of their own.
DEUT|14|28|At the end of every three years, bring all the tithes of that year's produce and store it in your towns,
DEUT|14|29|so that the Levites (who have no allotment or inheritance of their own) and the aliens, the fatherless and the widows who live in your towns may come and eat and be satisfied, and so that the LORD your God may bless you in all the work of your hands.
DEUT|15|1|At the end of every seven years you must cancel debts.
DEUT|15|2|This is how it is to be done: Every creditor shall cancel the loan he has made to his fellow Israelite. He shall not require payment from his fellow Israelite or brother, because the LORD's time for canceling debts has been proclaimed.
DEUT|15|3|You may require payment from a foreigner, but you must cancel any debt your brother owes you.
DEUT|15|4|However, there should be no poor among you, for in the land the LORD your God is giving you to possess as your inheritance, he will richly bless you,
DEUT|15|5|if only you fully obey the LORD your God and are careful to follow all these commands I am giving you today.
DEUT|15|6|For the LORD your God will bless you as he has promised, and you will lend to many nations but will borrow from none. You will rule over many nations but none will rule over you.
DEUT|15|7|If there is a poor man among your brothers in any of the towns of the land that the LORD your God is giving you, do not be hardhearted or tightfisted toward your poor brother.
DEUT|15|8|Rather be openhanded and freely lend him whatever he needs.
DEUT|15|9|Be careful not to harbor this wicked thought: "The seventh year, the year for canceling debts, is near," so that you do not show ill will toward your needy brother and give him nothing. He may then appeal to the LORD against you, and you will be found guilty of sin.
DEUT|15|10|Give generously to him and do so without a grudging heart; then because of this the LORD your God will bless you in all your work and in everything you put your hand to.
DEUT|15|11|There will always be poor people in the land. Therefore I command you to be openhanded toward your brothers and toward the poor and needy in your land.
DEUT|15|12|If a fellow Hebrew, a man or a woman, sells himself to you and serves you six years, in the seventh year you must let him go free.
DEUT|15|13|And when you release him, do not send him away empty-handed.
DEUT|15|14|Supply him liberally from your flock, your threshing floor and your winepress. Give to him as the LORD your God has blessed you.
DEUT|15|15|Remember that you were slaves in Egypt and the LORD your God redeemed you. That is why I give you this command today.
DEUT|15|16|But if your servant says to you, "I do not want to leave you," because he loves you and your family and is well off with you,
DEUT|15|17|then take an awl and push it through his ear lobe into the door, and he will become your servant for life. Do the same for your maidservant.
DEUT|15|18|Do not consider it a hardship to set your servant free, because his service to you these six years has been worth twice as much as that of a hired hand. And the LORD your God will bless you in everything you do.
DEUT|15|19|Set apart for the LORD your God every firstborn male of your herds and flocks. Do not put the firstborn of your oxen to work, and do not shear the firstborn of your sheep.
DEUT|15|20|Each year you and your family are to eat them in the presence of the LORD your God at the place he will choose.
DEUT|15|21|If an animal has a defect, is lame or blind, or has any serious flaw, you must not sacrifice it to the LORD your God.
DEUT|15|22|You are to eat it in your own towns. Both the ceremonially unclean and the clean may eat it, as if it were gazelle or deer.
DEUT|15|23|But you must not eat the blood; pour it out on the ground like water.
DEUT|16|1|Observe the month of Abib and celebrate the Passover of the LORD your God, because in the month of Abib he brought you out of Egypt by night.
DEUT|16|2|Sacrifice as the Passover to the LORD your God an animal from your flock or herd at the place the LORD will choose as a dwelling for his Name.
DEUT|16|3|Do not eat it with bread made with yeast, but for seven days eat unleavened bread, the bread of affliction, because you left Egypt in haste-so that all the days of your life you may remember the time of your departure from Egypt.
DEUT|16|4|Let no yeast be found in your possession in all your land for seven days. Do not let any of the meat you sacrifice on the evening of the first day remain until morning.
DEUT|16|5|You must not sacrifice the Passover in any town the LORD your God gives you
DEUT|16|6|except in the place he will choose as a dwelling for his Name. There you must sacrifice the Passover in the evening, when the sun goes down, on the anniversary of your departure from Egypt.
DEUT|16|7|Roast it and eat it at the place the LORD your God will choose. Then in the morning return to your tents.
DEUT|16|8|For six days eat unleavened bread and on the seventh day hold an assembly to the LORD your God and do no work.
DEUT|16|9|Count off seven weeks from the time you begin to put the sickle to the standing grain.
DEUT|16|10|Then celebrate the Feast of Weeks to the LORD your God by giving a freewill offering in proportion to the blessings the LORD your God has given you.
DEUT|16|11|And rejoice before the LORD your God at the place he will choose as a dwelling for his Name-you, your sons and daughters, your menservants and maidservants, the Levites in your towns, and the aliens, the fatherless and the widows living among you.
DEUT|16|12|Remember that you were slaves in Egypt, and follow carefully these decrees.
DEUT|16|13|Celebrate the Feast of Tabernacles for seven days after you have gathered the produce of your threshing floor and your winepress.
DEUT|16|14|Be joyful at your Feast-you, your sons and daughters, your menservants and maidservants, and the Levites, the aliens, the fatherless and the widows who live in your towns.
DEUT|16|15|For seven days celebrate the Feast to the LORD your God at the place the LORD will choose. For the LORD your God will bless you in all your harvest and in all the work of your hands, and your joy will be complete.
DEUT|16|16|Three times a year all your men must appear before the LORD your God at the place he will choose: at the Feast of Unleavened Bread, the Feast of Weeks and the Feast of Tabernacles. No man should appear before the LORD empty-handed:
DEUT|16|17|Each of you must bring a gift in proportion to the way the LORD your God has blessed you.
DEUT|16|18|Appoint judges and officials for each of your tribes in every town the LORD your God is giving you, and they shall judge the people fairly.
DEUT|16|19|Do not pervert justice or show partiality. Do not accept a bribe, for a bribe blinds the eyes of the wise and twists the words of the righteous.
DEUT|16|20|Follow justice and justice alone, so that you may live and possess the land the LORD your God is giving you.
DEUT|16|21|Do not set up any wooden Asherah pole beside the altar you build to the LORD your God,
DEUT|16|22|and do not erect a sacred stone, for these the LORD your God hates.
DEUT|17|1|Do not sacrifice to the LORD your God an ox or a sheep that has any defect or flaw in it, for that would be detestable to him.
DEUT|17|2|If a man or woman living among you in one of the towns the LORD gives you is found doing evil in the eyes of the LORD your God in violation of his covenant,
DEUT|17|3|and contrary to my command has worshiped other gods, bowing down to them or to the sun or the moon or the stars of the sky,
DEUT|17|4|and this has been brought to your attention, then you must investigate it thoroughly. If it is true and it has been proved that this detestable thing has been done in Israel,
DEUT|17|5|take the man or woman who has done this evil deed to your city gate and stone that person to death.
DEUT|17|6|On the testimony of two or three witnesses a man shall be put to death, but no one shall be put to death on the testimony of only one witness.
DEUT|17|7|The hands of the witnesses must be the first in putting him to death, and then the hands of all the people. You must purge the evil from among you.
DEUT|17|8|If cases come before your courts that are too difficult for you to judge-whether bloodshed, lawsuits or assaults-take them to the place the LORD your God will choose.
DEUT|17|9|Go to the priests, who are Levites, and to the judge who is in office at that time. Inquire of them and they will give you the verdict.
DEUT|17|10|You must act according to the decisions they give you at the place the LORD will choose. Be careful to do everything they direct you to do.
DEUT|17|11|Act according to the law they teach you and the decisions they give you. Do not turn aside from what they tell you, to the right or to the left.
DEUT|17|12|The man who shows contempt for the judge or for the priest who stands ministering there to the LORD your God must be put to death. You must purge the evil from Israel.
DEUT|17|13|All the people will hear and be afraid, and will not be contemptuous again.
DEUT|17|14|When you enter the land the LORD your God is giving you and have taken possession of it and settled in it, and you say, "Let us set a king over us like all the nations around us,"
DEUT|17|15|be sure to appoint over you the king the LORD your God chooses. He must be from among your own brothers. Do not place a foreigner over you, one who is not a brother Israelite.
DEUT|17|16|The king, moreover, must not acquire great numbers of horses for himself or make the people return to Egypt to get more of them, for the LORD has told you, "You are not to go back that way again."
DEUT|17|17|He must not take many wives, or his heart will be led astray. He must not accumulate large amounts of silver and gold.
DEUT|17|18|When he takes the throne of his kingdom, he is to write for himself on a scroll a copy of this law, taken from that of the priests, who are Levites.
DEUT|17|19|It is to be with him, and he is to read it all the days of his life so that he may learn to revere the LORD his God and follow carefully all the words of this law and these decrees
DEUT|17|20|and not consider himself better than his brothers and turn from the law to the right or to the left. Then he and his descendants will reign a long time over his kingdom in Israel.
DEUT|18|1|The priests, who are Levites-indeed the whole tribe of Levi-are to have no allotment or inheritance with Israel. They shall live on the offerings made to the LORD by fire, for that is their inheritance.
DEUT|18|2|They shall have no inheritance among their brothers; the LORD is their inheritance, as he promised them.
DEUT|18|3|This is the share due the priests from the people who sacrifice a bull or a sheep: the shoulder, the jowls and the inner parts.
DEUT|18|4|You are to give them the firstfruits of your grain, new wine and oil, and the first wool from the shearing of your sheep,
DEUT|18|5|for the LORD your God has chosen them and their descendants out of all your tribes to stand and minister in the LORD's name always.
DEUT|18|6|If a Levite moves from one of your towns anywhere in Israel where he is living, and comes in all earnestness to the place the LORD will choose,
DEUT|18|7|he may minister in the name of the LORD his God like all his fellow Levites who serve there in the presence of the LORD.
DEUT|18|8|He is to share equally in their benefits, even though he has received money from the sale of family possessions.
DEUT|18|9|When you enter the land the LORD your God is giving you, do not learn to imitate the detestable ways of the nations there.
DEUT|18|10|Let no one be found among you who sacrifices his son or daughter in the fire, who practices divination or sorcery, interprets omens, engages in witchcraft,
DEUT|18|11|or casts spells, or who is a medium or spiritist or who consults the dead.
DEUT|18|12|Anyone who does these things is detestable to the LORD, and because of these detestable practices the LORD your God will drive out those nations before you.
DEUT|18|13|You must be blameless before the LORD your God.
DEUT|18|14|The nations you will dispossess listen to those who practice sorcery or divination. But as for you, the LORD your God has not permitted you to do so.
DEUT|18|15|The LORD your God will raise up for you a prophet like me from among your own brothers. You must listen to him.
DEUT|18|16|For this is what you asked of the LORD your God at Horeb on the day of the assembly when you said, "Let us not hear the voice of the LORD our God nor see this great fire anymore, or we will die."
DEUT|18|17|The LORD said to me: "What they say is good.
DEUT|18|18|I will raise up for them a prophet like you from among their brothers; I will put my words in his mouth, and he will tell them everything I command him.
DEUT|18|19|If anyone does not listen to my words that the prophet speaks in my name, I myself will call him to account.
DEUT|18|20|But a prophet who presumes to speak in my name anything I have not commanded him to say, or a prophet who speaks in the name of other gods, must be put to death."
DEUT|18|21|You may say to yourselves, "How can we know when a message has not been spoken by the LORD?"
DEUT|18|22|If what a prophet proclaims in the name of the LORD does not take place or come true, that is a message the LORD has not spoken. That prophet has spoken presumptuously. Do not be afraid of him.
DEUT|19|1|When the LORD your God has destroyed the nations whose land he is giving you, and when you have driven them out and settled in their towns and houses,
DEUT|19|2|then set aside for yourselves three cities centrally located in the land the LORD your God is giving you to possess.
DEUT|19|3|Build roads to them and divide into three parts the land the LORD your God is giving you as an inheritance, so that anyone who kills a man may flee there.
DEUT|19|4|This is the rule concerning the man who kills another and flees there to save his life-one who kills his neighbor unintentionally, without malice aforethought.
DEUT|19|5|For instance, a man may go into the forest with his neighbor to cut wood, and as he swings his ax to fell a tree, the head may fly off and hit his neighbor and kill him. That man may flee to one of these cities and save his life.
DEUT|19|6|Otherwise, the avenger of blood might pursue him in a rage, overtake him if the distance is too great, and kill him even though he is not deserving of death, since he did it to his neighbor without malice aforethought.
DEUT|19|7|This is why I command you to set aside for yourselves three cities.
DEUT|19|8|If the LORD your God enlarges your territory, as he promised on oath to your forefathers, and gives you the whole land he promised them,
DEUT|19|9|because you carefully follow all these laws I command you today-to love the LORD your God and to walk always in his ways-then you are to set aside three more cities.
DEUT|19|10|Do this so that innocent blood will not be shed in your land, which the LORD your God is giving you as your inheritance, and so that you will not be guilty of bloodshed.
DEUT|19|11|But if a man hates his neighbor and lies in wait for him, assaults and kills him, and then flees to one of these cities,
DEUT|19|12|the elders of his town shall send for him, bring him back from the city, and hand him over to the avenger of blood to die.
DEUT|19|13|Show him no pity. You must purge from Israel the guilt of shedding innocent blood, so that it may go well with you.
DEUT|19|14|Do not move your neighbor's boundary stone set up by your predecessors in the inheritance you receive in the land the LORD your God is giving you to possess.
DEUT|19|15|One witness is not enough to convict a man accused of any crime or offense he may have committed. A matter must be established by the testimony of two or three witnesses.
DEUT|19|16|If a malicious witness takes the stand to accuse a man of a crime,
DEUT|19|17|the two men involved in the dispute must stand in the presence of the LORD before the priests and the judges who are in office at the time.
DEUT|19|18|The judges must make a thorough investigation, and if the witness proves to be a liar, giving false testimony against his brother,
DEUT|19|19|then do to him as he intended to do to his brother. You must purge the evil from among you.
DEUT|19|20|The rest of the people will hear of this and be afraid, and never again will such an evil thing be done among you.
DEUT|19|21|Show no pity: life for life, eye for eye, tooth for tooth, hand for hand, foot for foot.
DEUT|20|1|When you go to war against your enemies and see horses and chariots and an army greater than yours, do not be afraid of them, because the LORD your God, who brought you up out of Egypt, will be with you.
DEUT|20|2|When you are about to go into battle, the priest shall come forward and address the army.
DEUT|20|3|He shall say: "Hear, O Israel, today you are going into battle against your enemies. Do not be fainthearted or afraid; do not be terrified or give way to panic before them.
DEUT|20|4|For the LORD your God is the one who goes with you to fight for you against your enemies to give you victory."
DEUT|20|5|The officers shall say to the army: "Has anyone built a new house and not dedicated it? Let him go home, or he may die in battle and someone else may dedicate it.
DEUT|20|6|Has anyone planted a vineyard and not begun to enjoy it? Let him go home, or he may die in battle and someone else enjoy it.
DEUT|20|7|Has anyone become pledged to a woman and not married her? Let him go home, or he may die in battle and someone else marry her."
DEUT|20|8|Then the officers shall add, "Is any man afraid or fainthearted? Let him go home so that his brothers will not become disheartened too."
DEUT|20|9|When the officers have finished speaking to the army, they shall appoint commanders over it.
DEUT|20|10|When you march up to attack a city, make its people an offer of peace.
DEUT|20|11|If they accept and open their gates, all the people in it shall be subject to forced labor and shall work for you.
DEUT|20|12|If they refuse to make peace and they engage you in battle, lay siege to that city.
DEUT|20|13|When the LORD your God delivers it into your hand, put to the sword all the men in it.
DEUT|20|14|As for the women, the children, the livestock and everything else in the city, you may take these as plunder for yourselves. And you may use the plunder the LORD your God gives you from your enemies.
DEUT|20|15|This is how you are to treat all the cities that are at a distance from you and do not belong to the nations nearby.
DEUT|20|16|However, in the cities of the nations the LORD your God is giving you as an inheritance, do not leave alive anything that breathes.
DEUT|20|17|Completely destroy them-the Hittites, Amorites, Canaanites, Perizzites, Hivites and Jebusites-as the LORD your God has commanded you.
DEUT|20|18|Otherwise, they will teach you to follow all the detestable things they do in worshiping their gods, and you will sin against the LORD your God.
DEUT|20|19|When you lay siege to a city for a long time, fighting against it to capture it, do not destroy its trees by putting an ax to them, because you can eat their fruit. Do not cut them down. Are the trees of the field people, that you should besiege them?
DEUT|20|20|However, you may cut down trees that you know are not fruit trees and use them to build siege works until the city at war with you falls.
DEUT|21|1|If a man is found slain, lying in a field in the land the LORD your God is giving you to possess, and it is not known who killed him,
DEUT|21|2|your elders and judges shall go out and measure the distance from the body to the neighboring towns.
DEUT|21|3|Then the elders of the town nearest the body shall take a heifer that has never been worked and has never worn a yoke
DEUT|21|4|and lead her down to a valley that has not been plowed or planted and where there is a flowing stream. There in the valley they are to break the heifer's neck.
DEUT|21|5|The priests, the sons of Levi, shall step forward, for the LORD your God has chosen them to minister and to pronounce blessings in the name of the LORD and to decide all cases of dispute and assault.
DEUT|21|6|Then all the elders of the town nearest the body shall wash their hands over the heifer whose neck was broken in the valley,
DEUT|21|7|and they shall declare: "Our hands did not shed this blood, nor did our eyes see it done.
DEUT|21|8|Accept this atonement for your people Israel, whom you have redeemed, O LORD, and do not hold your people guilty of the blood of an innocent man." And the bloodshed will be atoned for.
DEUT|21|9|So you will purge from yourselves the guilt of shedding innocent blood, since you have done what is right in the eyes of the LORD.
DEUT|21|10|When you go to war against your enemies and the LORD your God delivers them into your hands and you take captives,
DEUT|21|11|if you notice among the captives a beautiful woman and are attracted to her, you may take her as your wife.
DEUT|21|12|Bring her into your home and have her shave her head, trim her nails
DEUT|21|13|and put aside the clothes she was wearing when captured. After she has lived in your house and mourned her father and mother for a full month, then you may go to her and be her husband and she shall be your wife.
DEUT|21|14|If you are not pleased with her, let her go wherever she wishes. You must not sell her or treat her as a slave, since you have dishonored her.
DEUT|21|15|If a man has two wives, and he loves one but not the other, and both bear him sons but the firstborn is the son of the wife he does not love,
DEUT|21|16|when he wills his property to his sons, he must not give the rights of the firstborn to the son of the wife he loves in preference to his actual firstborn, the son of the wife he does not love.
DEUT|21|17|He must acknowledge the son of his unloved wife as the firstborn by giving him a double share of all he has. That son is the first sign of his father's strength. The right of the firstborn belongs to him.
DEUT|21|18|If a man has a stubborn and rebellious son who does not obey his father and mother and will not listen to them when they discipline him,
DEUT|21|19|his father and mother shall take hold of him and bring him to the elders at the gate of his town.
DEUT|21|20|They shall say to the elders, "This son of ours is stubborn and rebellious. He will not obey us. He is a profligate and a drunkard."
DEUT|21|21|Then all the men of his town shall stone him to death. You must purge the evil from among you. All Israel will hear of it and be afraid.
DEUT|21|22|If a man guilty of a capital offense is put to death and his body is hung on a tree,
DEUT|21|23|you must not leave his body on the tree overnight. Be sure to bury him that same day, because anyone who is hung on a tree is under God's curse. You must not desecrate the land the LORD your God is giving you as an inheritance.
DEUT|22|1|If you see your brother's ox or sheep straying, do not ignore it but be sure to take it back to him.
DEUT|22|2|If the brother does not live near you or if you do not know who he is, take it home with you and keep it until he comes looking for it. Then give it back to him.
DEUT|22|3|Do the same if you find your brother's donkey or his cloak or anything he loses. Do not ignore it.
DEUT|22|4|If you see your brother's donkey or his ox fallen on the road, do not ignore it. Help him get it to its feet.
DEUT|22|5|A woman must not wear men's clothing, nor a man wear women's clothing, for the LORD your God detests anyone who does this.
DEUT|22|6|If you come across a bird's nest beside the road, either in a tree or on the ground, and the mother is sitting on the young or on the eggs, do not take the mother with the young.
DEUT|22|7|You may take the young, but be sure to let the mother go, so that it may go well with you and you may have a long life.
DEUT|22|8|When you build a new house, make a parapet around your roof so that you may not bring the guilt of bloodshed on your house if someone falls from the roof.
DEUT|22|9|Do not plant two kinds of seed in your vineyard; if you do, not only the crops you plant but also the fruit of the vineyard will be defiled.
DEUT|22|10|Do not plow with an ox and a donkey yoked together.
DEUT|22|11|Do not wear clothes of wool and linen woven together.
DEUT|22|12|Make tassels on the four corners of the cloak you wear.
DEUT|22|13|If a man takes a wife and, after lying with her, dislikes her
DEUT|22|14|and slanders her and gives her a bad name, saying, "I married this woman, but when I approached her, I did not find proof of her virginity,"
DEUT|22|15|then the girl's father and mother shall bring proof that she was a virgin to the town elders at the gate.
DEUT|22|16|The girl's father will say to the elders, "I gave my daughter in marriage to this man, but he dislikes her.
DEUT|22|17|Now he has slandered her and said, 'I did not find your daughter to be a virgin.' But here is the proof of my daughter's virginity." Then her parents shall display the cloth before the elders of the town,
DEUT|22|18|and the elders shall take the man and punish him.
DEUT|22|19|They shall fine him a hundred shekels of silver and give them to the girl's father, because this man has given an Israelite virgin a bad name. She shall continue to be his wife; he must not divorce her as long as he lives.
DEUT|22|20|If, however, the charge is true and no proof of the girl's virginity can be found,
DEUT|22|21|she shall be brought to the door of her father's house and there the men of her town shall stone her to death. She has done a disgraceful thing in Israel by being promiscuous while still in her father's house. You must purge the evil from among you.
DEUT|22|22|If a man is found sleeping with another man's wife, both the man who slept with her and the woman must die. You must purge the evil from Israel.
DEUT|22|23|If a man happens to meet in a town a virgin pledged to be married and he sleeps with her,
DEUT|22|24|you shall take both of them to the gate of that town and stone them to death-the girl because she was in a town and did not scream for help, and the man because he violated another man's wife. You must purge the evil from among you.
DEUT|22|25|But if out in the country a man happens to meet a girl pledged to be married and rapes her, only the man who has done this shall die.
DEUT|22|26|Do nothing to the girl; she has committed no sin deserving death. This case is like that of someone who attacks and murders his neighbor,
DEUT|22|27|for the man found the girl out in the country, and though the betrothed girl screamed, there was no one to rescue her.
DEUT|22|28|If a man happens to meet a virgin who is not pledged to be married and rapes her and they are discovered,
DEUT|22|29|he shall pay the girl's father fifty shekels of silver. He must marry the girl, for he has violated her. He can never divorce her as long as he lives.
DEUT|22|30|A man is not to marry his father's wife; he must not dishonor his father's bed.
DEUT|23|1|No one who has been emasculated by crushing or cutting may enter the assembly of the LORD.
DEUT|23|2|No one born of a forbidden marriage nor any of his descendants may enter the assembly of the LORD, even down to the tenth generation.
DEUT|23|3|No Ammonite or Moabite or any of his descendants may enter the assembly of the LORD, even down to the tenth generation.
DEUT|23|4|For they did not come to meet you with bread and water on your way when you came out of Egypt, and they hired Balaam son of Beor from Pethor in Aram Naharaim to pronounce a curse on you.
DEUT|23|5|However, the LORD your God would not listen to Balaam but turned the curse into a blessing for you, because the LORD your God loves you.
DEUT|23|6|Do not seek a treaty of friendship with them as long as you live.
DEUT|23|7|Do not abhor an Edomite, for he is your brother. Do not abhor an Egyptian, because you lived as an alien in his country.
DEUT|23|8|The third generation of children born to them may enter the assembly of the LORD.
DEUT|23|9|When you are encamped against your enemies, keep away from everything impure.
DEUT|23|10|If one of your men is unclean because of a nocturnal emission, he is to go outside the camp and stay there.
DEUT|23|11|But as evening approaches he is to wash himself, and at sunset he may return to the camp.
DEUT|23|12|Designate a place outside the camp where you can go to relieve yourself.
DEUT|23|13|As part of your equipment have something to dig with, and when you relieve yourself, dig a hole and cover up your excrement.
DEUT|23|14|For the LORD your God moves about in your camp to protect you and to deliver your enemies to you. Your camp must be holy, so that he will not see among you anything indecent and turn away from you.
DEUT|23|15|If a slave has taken refuge with you, do not hand him over to his master.
DEUT|23|16|Let him live among you wherever he likes and in whatever town he chooses. Do not oppress him.
DEUT|23|17|No Israelite man or woman is to become a shrine prostitute.
DEUT|23|18|You must not bring the earnings of a female prostitute or of a male prostitute into the house of the LORD your God to pay any vow, because the LORD your God detests them both.
DEUT|23|19|Do not charge your brother interest, whether on money or food or anything else that may earn interest.
DEUT|23|20|You may charge a foreigner interest, but not a brother Israelite, so that the LORD your God may bless you in everything you put your hand to in the land you are entering to possess.
DEUT|23|21|If you make a vow to the LORD your God, do not be slow to pay it, for the LORD your God will certainly demand it of you and you will be guilty of sin.
DEUT|23|22|But if you refrain from making a vow, you will not be guilty.
DEUT|23|23|Whatever your lips utter you must be sure to do, because you made your vow freely to the LORD your God with your own mouth.
DEUT|23|24|If you enter your neighbor's vineyard, you may eat all the grapes you want, but do not put any in your basket.
DEUT|23|25|If you enter your neighbor's grainfield, you may pick kernels with your hands, but you must not put a sickle to his standing grain.
DEUT|24|1|If a man marries a woman who becomes displeasing to him because he finds something indecent about her, and he writes her a certificate of divorce, gives it to her and sends her from his house,
DEUT|24|2|and if after she leaves his house she becomes the wife of another man,
DEUT|24|3|and her second husband dislikes her and writes her a certificate of divorce, gives it to her and sends her from his house, or if he dies,
DEUT|24|4|then her first husband, who divorced her, is not allowed to marry her again after she has been defiled. That would be detestable in the eyes of the LORD. Do not bring sin upon the land the LORD your God is giving you as an inheritance.
DEUT|24|5|If a man has recently married, he must not be sent to war or have any other duty laid on him. For one year he is to be free to stay at home and bring happiness to the wife he has married.
DEUT|24|6|Do not take a pair of millstones-not even the upper one-as security for a debt, because that would be taking a man's livelihood as security.
DEUT|24|7|If a man is caught kidnapping one of his brother Israelites and treats him as a slave or sells him, the kidnapper must die. You must purge the evil from among you.
DEUT|24|8|In cases of leprous diseases be very careful to do exactly as the priests, who are Levites, instruct you. You must follow carefully what I have commanded them.
DEUT|24|9|Remember what the LORD your God did to Miriam along the way after you came out of Egypt.
DEUT|24|10|When you make a loan of any kind to your neighbor, do not go into his house to get what he is offering as a pledge.
DEUT|24|11|Stay outside and let the man to whom you are making the loan bring the pledge out to you.
DEUT|24|12|If the man is poor, do not go to sleep with his pledge in your possession.
DEUT|24|13|Return his cloak to him by sunset so that he may sleep in it. Then he will thank you, and it will be regarded as a righteous act in the sight of the LORD your God.
DEUT|24|14|Do not take advantage of a hired man who is poor and needy, whether he is a brother Israelite or an alien living in one of your towns.
DEUT|24|15|Pay him his wages each day before sunset, because he is poor and is counting on it. Otherwise he may cry to the LORD against you, and you will be guilty of sin.
DEUT|24|16|Fathers shall not be put to death for their children, nor children put to death for their fathers; each is to die for his own sin.
DEUT|24|17|Do not deprive the alien or the fatherless of justice, or take the cloak of the widow as a pledge.
DEUT|24|18|Remember that you were slaves in Egypt and the LORD your God redeemed you from there. That is why I command you to do this.
DEUT|24|19|When you are harvesting in your field and you overlook a sheaf, do not go back to get it. Leave it for the alien, the fatherless and the widow, so that the LORD your God may bless you in all the work of your hands.
DEUT|24|20|When you beat the olives from your trees, do not go over the branches a second time. Leave what remains for the alien, the fatherless and the widow.
DEUT|24|21|When you harvest the grapes in your vineyard, do not go over the vines again. Leave what remains for the alien, the fatherless and the widow.
DEUT|24|22|Remember that you were slaves in Egypt. That is why I command you to do this.
DEUT|25|1|When men have a dispute, they are to take it to court and the judges will decide the case, acquitting the innocent and condemning the guilty.
DEUT|25|2|If the guilty man deserves to be beaten, the judge shall make him lie down and have him flogged in his presence with the number of lashes his crime deserves,
DEUT|25|3|but he must not give him more than forty lashes. If he is flogged more than that, your brother will be degraded in your eyes.
DEUT|25|4|Do not muzzle an ox while it is treading out the grain.
DEUT|25|5|If brothers are living together and one of them dies without a son, his widow must not marry outside the family. Her husband's brother shall take her and marry her and fulfill the duty of a brother-in-law to her.
DEUT|25|6|The first son she bears shall carry on the name of the dead brother so that his name will not be blotted out from Israel.
DEUT|25|7|However, if a man does not want to marry his brother's wife, she shall go to the elders at the town gate and say, "My husband's brother refuses to carry on his brother's name in Israel. He will not fulfill the duty of a brother-in-law to me."
DEUT|25|8|Then the elders of his town shall summon him and talk to him. If he persists in saying, "I do not want to marry her,"
DEUT|25|9|his brother's widow shall go up to him in the presence of the elders, take off one of his sandals, spit in his face and say, "This is what is done to the man who will not build up his brother's family line."
DEUT|25|10|That man's line shall be known in Israel as The Family of the Unsandaled.
DEUT|25|11|If two men are fighting and the wife of one of them comes to rescue her husband from his assailant, and she reaches out and seizes him by his private parts,
DEUT|25|12|you shall cut off her hand. Show her no pity.
DEUT|25|13|Do not have two differing weights in your bag-one heavy, one light.
DEUT|25|14|Do not have two differing measures in your house-one large, one small.
DEUT|25|15|You must have accurate and honest weights and measures, so that you may live long in the land the LORD your God is giving you.
DEUT|25|16|For the LORD your God detests anyone who does these things, anyone who deals dishonestly.
DEUT|25|17|Remember what the Amalekites did to you along the way when you came out of Egypt.
DEUT|25|18|When you were weary and worn out, they met you on your journey and cut off all who were lagging behind; they had no fear of God.
DEUT|25|19|When the LORD your God gives you rest from all the enemies around you in the land he is giving you to possess as an inheritance, you shall blot out the memory of Amalek from under heaven. Do not forget!
DEUT|26|1|When you have entered the land the LORD your God is giving you as an inheritance and have taken possession of it and settled in it,
DEUT|26|2|take some of the firstfruits of all that you produce from the soil of the land the LORD your God is giving you and put them in a basket. Then go to the place the LORD your God will choose as a dwelling for his Name
DEUT|26|3|and say to the priest in office at the time, "I declare today to the LORD your God that I have come to the land the LORD swore to our forefathers to give us."
DEUT|26|4|The priest shall take the basket from your hands and set it down in front of the altar of the LORD your God.
DEUT|26|5|Then you shall declare before the LORD your God: "My father was a wandering Aramean, and he went down into Egypt with a few people and lived there and became a great nation, powerful and numerous.
DEUT|26|6|But the Egyptians mistreated us and made us suffer, putting us to hard labor.
DEUT|26|7|Then we cried out to the LORD, the God of our fathers, and the LORD heard our voice and saw our misery, toil and oppression.
DEUT|26|8|So the LORD brought us out of Egypt with a mighty hand and an outstretched arm, with great terror and with miraculous signs and wonders.
DEUT|26|9|He brought us to this place and gave us this land, a land flowing with milk and honey;
DEUT|26|10|and now I bring the firstfruits of the soil that you, O LORD, have given me." Place the basket before the LORD your God and bow down before him.
DEUT|26|11|And you and the Levites and the aliens among you shall rejoice in all the good things the LORD your God has given to you and your household.
DEUT|26|12|When you have finished setting aside a tenth of all your produce in the third year, the year of the tithe, you shall give it to the Levite, the alien, the fatherless and the widow, so that they may eat in your towns and be satisfied.
DEUT|26|13|Then say to the LORD your God: "I have removed from my house the sacred portion and have given it to the Levite, the alien, the fatherless and the widow, according to all you commanded. I have not turned aside from your commands nor have I forgotten any of them.
DEUT|26|14|I have not eaten any of the sacred portion while I was in mourning, nor have I removed any of it while I was unclean, nor have I offered any of it to the dead. I have obeyed the LORD my God; I have done everything you commanded me.
DEUT|26|15|Look down from heaven, your holy dwelling place, and bless your people Israel and the land you have given us as you promised on oath to our forefathers, a land flowing with milk and honey."
DEUT|26|16|The LORD your God commands you this day to follow these decrees and laws; carefully observe them with all your heart and with all your soul.
DEUT|26|17|You have declared this day that the LORD is your God and that you will walk in his ways, that you will keep his decrees, commands and laws, and that you will obey him.
DEUT|26|18|And the LORD has declared this day that you are his people, his treasured possession as he promised, and that you are to keep all his commands.
DEUT|26|19|He has declared that he will set you in praise, fame and honor high above all the nations he has made and that you will be a people holy to the LORD your God, as he promised.
DEUT|27|1|Moses and the elders of Israel commanded the people: "Keep all these commands that I give you today.
DEUT|27|2|When you have crossed the Jordan into the land the LORD your God is giving you, set up some large stones and coat them with plaster.
DEUT|27|3|Write on them all the words of this law when you have crossed over to enter the land the LORD your God is giving you, a land flowing with milk and honey, just as the LORD, the God of your fathers, promised you.
DEUT|27|4|And when you have crossed the Jordan, set up these stones on Mount Ebal, as I command you today, and coat them with plaster.
DEUT|27|5|Build there an altar to the LORD your God, an altar of stones. Do not use any iron tool upon them.
DEUT|27|6|Build the altar of the LORD your God with fieldstones and offer burnt offerings on it to the LORD your God.
DEUT|27|7|Sacrifice fellowship offerings there, eating them and rejoicing in the presence of the LORD your God.
DEUT|27|8|And you shall write very clearly all the words of this law on these stones you have set up."
DEUT|27|9|Then Moses and the priests, who are Levites, said to all Israel, "Be silent, O Israel, and listen! You have now become the people of the LORD your God.
DEUT|27|10|Obey the LORD your God and follow his commands and decrees that I give you today."
DEUT|27|11|On the same day Moses commanded the people:
DEUT|27|12|When you have crossed the Jordan, these tribes shall stand on Mount Gerizim to bless the people: Simeon, Levi, Judah, Issachar, Joseph and Benjamin.
DEUT|27|13|And these tribes shall stand on Mount Ebal to pronounce curses: Reuben, Gad, Asher, Zebulun, Dan and Naphtali.
DEUT|27|14|The Levites shall recite to all the people of Israel in a loud voice:
DEUT|27|15|"Cursed is the man who carves an image or casts an idol-a thing detestable to the LORD, the work of the craftsman's hands-and sets it up in secret." Then all the people shall say, "Amen!"
DEUT|27|16|"Cursed is the man who dishonors his father or his mother." Then all the people shall say, "Amen!"
DEUT|27|17|"Cursed is the man who moves his neighbor's boundary stone." Then all the people shall say, "Amen!"
DEUT|27|18|"Cursed is the man who leads the blind astray on the road." Then all the people shall say, "Amen!"
DEUT|27|19|"Cursed is the man who withholds justice from the alien, the fatherless or the widow." Then all the people shall say, "Amen!"
DEUT|27|20|"Cursed is the man who sleeps with his father's wife, for he dishonors his father's bed." Then all the people shall say, "Amen!"
DEUT|27|21|"Cursed is the man who has sexual relations with any animal." Then all the people shall say, "Amen!"
DEUT|27|22|"Cursed is the man who sleeps with his sister, the daughter of his father or the daughter of his mother." Then all the people shall say, "Amen!"
DEUT|27|23|"Cursed is the man who sleeps with his mother-in-law." Then all the people shall say, "Amen!"
DEUT|27|24|"Cursed is the man who kills his neighbor secretly." Then all the people shall say, "Amen!"
DEUT|27|25|"Cursed is the man who accepts a bribe to kill an innocent person." Then all the people shall say, "Amen!"
DEUT|27|26|"Cursed is the man who does not uphold the words of this law by carrying them out." Then all the people shall say, "Amen!"
DEUT|28|1|If you fully obey the LORD your God and carefully follow all his commands I give you today, the LORD your God will set you high above all the nations on earth.
DEUT|28|2|All these blessings will come upon you and accompany you if you obey the LORD your God:
DEUT|28|3|You will be blessed in the city and blessed in the country.
DEUT|28|4|The fruit of your womb will be blessed, and the crops of your land and the young of your livestock-the calves of your herds and the lambs of your flocks.
DEUT|28|5|Your basket and your kneading trough will be blessed.
DEUT|28|6|You will be blessed when you come in and blessed when you go out.
DEUT|28|7|The LORD will grant that the enemies who rise up against you will be defeated before you. They will come at you from one direction but flee from you in seven.
DEUT|28|8|The LORD will send a blessing on your barns and on everything you put your hand to. The LORD your God will bless you in the land he is giving you.
DEUT|28|9|The LORD will establish you as his holy people, as he promised you on oath, if you keep the commands of the LORD your God and walk in his ways.
DEUT|28|10|Then all the peoples on earth will see that you are called by the name of the LORD, and they will fear you.
DEUT|28|11|The LORD will grant you abundant prosperity-in the fruit of your womb, the young of your livestock and the crops of your ground-in the land he swore to your forefathers to give you.
DEUT|28|12|The LORD will open the heavens, the storehouse of his bounty, to send rain on your land in season and to bless all the work of your hands. You will lend to many nations but will borrow from none.
DEUT|28|13|The LORD will make you the head, not the tail. If you pay attention to the commands of the LORD your God that I give you this day and carefully follow them, you will always be at the top, never at the bottom.
DEUT|28|14|Do not turn aside from any of the commands I give you today, to the right or to the left, following other gods and serving them.
DEUT|28|15|However, if you do not obey the LORD your God and do not carefully follow all his commands and decrees I am giving you today, all these curses will come upon you and overtake you:
DEUT|28|16|You will be cursed in the city and cursed in the country.
DEUT|28|17|Your basket and your kneading trough will be cursed.
DEUT|28|18|The fruit of your womb will be cursed, and the crops of your land, and the calves of your herds and the lambs of your flocks.
DEUT|28|19|You will be cursed when you come in and cursed when you go out.
DEUT|28|20|The LORD will send on you curses, confusion and rebuke in everything you put your hand to, until you are destroyed and come to sudden ruin because of the evil you have done in forsaking him.
DEUT|28|21|The LORD will plague you with diseases until he has destroyed you from the land you are entering to possess.
DEUT|28|22|The LORD will strike you with wasting disease, with fever and inflammation, with scorching heat and drought, with blight and mildew, which will plague you until you perish.
DEUT|28|23|The sky over your head will be bronze, the ground beneath you iron.
DEUT|28|24|The LORD will turn the rain of your country into dust and powder; it will come down from the skies until you are destroyed.
DEUT|28|25|The LORD will cause you to be defeated before your enemies. You will come at them from one direction but flee from them in seven, and you will become a thing of horror to all the kingdoms on earth.
DEUT|28|26|Your carcasses will be food for all the birds of the air and the beasts of the earth, and there will be no one to frighten them away.
DEUT|28|27|The LORD will afflict you with the boils of Egypt and with tumors, festering sores and the itch, from which you cannot be cured.
DEUT|28|28|The LORD will afflict you with madness, blindness and confusion of mind.
DEUT|28|29|At midday you will grope about like a blind man in the dark. You will be unsuccessful in everything you do; day after day you will be oppressed and robbed, with no one to rescue you.
DEUT|28|30|You will be pledged to be married to a woman, but another will take her and ravish her. You will build a house, but you will not live in it. You will plant a vineyard, but you will not even begin to enjoy its fruit.
DEUT|28|31|Your ox will be slaughtered before your eyes, but you will eat none of it. Your donkey will be forcibly taken from you and will not be returned. Your sheep will be given to your enemies, and no one will rescue them.
DEUT|28|32|Your sons and daughters will be given to another nation, and you will wear out your eyes watching for them day after day, powerless to lift a hand.
DEUT|28|33|A people that you do not know will eat what your land and labor produce, and you will have nothing but cruel oppression all your days.
DEUT|28|34|The sights you see will drive you mad.
DEUT|28|35|The LORD will afflict your knees and legs with painful boils that cannot be cured, spreading from the soles of your feet to the top of your head.
DEUT|28|36|The LORD will drive you and the king you set over you to a nation unknown to you or your fathers. There you will worship other gods, gods of wood and stone.
DEUT|28|37|You will become a thing of horror and an object of scorn and ridicule to all the nations where the LORD will drive you.
DEUT|28|38|You will sow much seed in the field but you will harvest little, because locusts will devour it.
DEUT|28|39|You will plant vineyards and cultivate them but you will not drink the wine or gather the grapes, because worms will eat them.
DEUT|28|40|You will have olive trees throughout your country but you will not use the oil, because the olives will drop off.
DEUT|28|41|You will have sons and daughters but you will not keep them, because they will go into captivity.
DEUT|28|42|Swarms of locusts will take over all your trees and the crops of your land.
DEUT|28|43|The alien who lives among you will rise above you higher and higher, but you will sink lower and lower.
DEUT|28|44|He will lend to you, but you will not lend to him. He will be the head, but you will be the tail.
DEUT|28|45|All these curses will come upon you. They will pursue you and overtake you until you are destroyed, because you did not obey the LORD your God and observe the commands and decrees he gave you.
DEUT|28|46|They will be a sign and a wonder to you and your descendants forever.
DEUT|28|47|Because you did not serve the LORD your God joyfully and gladly in the time of prosperity,
DEUT|28|48|therefore in hunger and thirst, in nakedness and dire poverty, you will serve the enemies the LORD sends against you. He will put an iron yoke on your neck until he has destroyed you.
DEUT|28|49|The LORD will bring a nation against you from far away, from the ends of the earth, like an eagle swooping down, a nation whose language you will not understand,
DEUT|28|50|a fierce-looking nation without respect for the old or pity for the young.
DEUT|28|51|They will devour the young of your livestock and the crops of your land until you are destroyed. They will leave you no grain, new wine or oil, nor any calves of your herds or lambs of your flocks until you are ruined.
DEUT|28|52|They will lay siege to all the cities throughout your land until the high fortified walls in which you trust fall down. They will besiege all the cities throughout the land the LORD your God is giving you.
DEUT|28|53|Because of the suffering that your enemy will inflict on you during the siege, you will eat the fruit of the womb, the flesh of the sons and daughters the LORD your God has given you.
DEUT|28|54|Even the most gentle and sensitive man among you will have no compassion on his own brother or the wife he loves or his surviving children,
DEUT|28|55|and he will not give to one of them any of the flesh of his children that he is eating. It will be all he has left because of the suffering your enemy will inflict on you during the siege of all your cities.
DEUT|28|56|The most gentle and sensitive woman among you-so sensitive and gentle that she would not venture to touch the ground with the sole of her foot-will begrudge the husband she loves and her own son or daughter
DEUT|28|57|the afterbirth from her womb and the children she bears. For she intends to eat them secretly during the siege and in the distress that your enemy will inflict on you in your cities.
DEUT|28|58|If you do not carefully follow all the words of this law, which are written in this book, and do not revere this glorious and awesome name-the LORD your God-
DEUT|28|59|the LORD will send fearful plagues on you and your descendants, harsh and prolonged disasters, and severe and lingering illnesses.
DEUT|28|60|He will bring upon you all the diseases of Egypt that you dreaded, and they will cling to you.
DEUT|28|61|The LORD will also bring on you every kind of sickness and disaster not recorded in this Book of the Law, until you are destroyed.
DEUT|28|62|You who were as numerous as the stars in the sky will be left but few in number, because you did not obey the LORD your God.
DEUT|28|63|Just as it pleased the LORD to make you prosper and increase in number, so it will please him to ruin and destroy you. You will be uprooted from the land you are entering to possess.
DEUT|28|64|Then the LORD will scatter you among all nations, from one end of the earth to the other. There you will worship other gods-gods of wood and stone, which neither you nor your fathers have known.
DEUT|28|65|Among those nations you will find no repose, no resting place for the sole of your foot. There the LORD will give you an anxious mind, eyes weary with longing, and a despairing heart.
DEUT|28|66|You will live in constant suspense, filled with dread both night and day, never sure of your life.
DEUT|28|67|In the morning you will say, "If only it were evening!" and in the evening, "If only it were morning!"-because of the terror that will fill your hearts and the sights that your eyes will see.
DEUT|28|68|The LORD will send you back in ships to Egypt on a journey I said you should never make again. There you will offer yourselves for sale to your enemies as male and female slaves, but no one will buy you.
DEUT|29|1|These are the terms of the covenant the LORD commanded Moses to make with the Israelites in Moab, in addition to the covenant he had made with them at Horeb.
DEUT|29|2|Moses summoned all the Israelites and said to them: Your eyes have seen all that the LORD did in Egypt to Pharaoh, to all his officials and to all his land.
DEUT|29|3|With your own eyes you saw those great trials, those miraculous signs and great wonders.
DEUT|29|4|But to this day the LORD has not given you a mind that understands or eyes that see or ears that hear.
DEUT|29|5|During the forty years that I led you through the desert, your clothes did not wear out, nor did the sandals on your feet.
DEUT|29|6|You ate no bread and drank no wine or other fermented drink. I did this so that you might know that I am the LORD your God.
DEUT|29|7|When you reached this place, Sihon king of Heshbon and Og king of Bashan came out to fight against us, but we defeated them.
DEUT|29|8|We took their land and gave it as an inheritance to the Reubenites, the Gadites and the half-tribe of Manasseh.
DEUT|29|9|Carefully follow the terms of this covenant, so that you may prosper in everything you do.
DEUT|29|10|All of you are standing today in the presence of the LORD your God-your leaders and chief men, your elders and officials, and all the other men of Israel,
DEUT|29|11|together with your children and your wives, and the aliens living in your camps who chop your wood and carry your water.
DEUT|29|12|You are standing here in order to enter into a covenant with the LORD your God, a covenant the LORD is making with you this day and sealing with an oath,
DEUT|29|13|to confirm you this day as his people, that he may be your God as he promised you and as he swore to your fathers, Abraham, Isaac and Jacob.
DEUT|29|14|I am making this covenant, with its oath, not only with you
DEUT|29|15|who are standing here with us today in the presence of the LORD our God but also with those who are not here today.
DEUT|29|16|You yourselves know how we lived in Egypt and how we passed through the countries on the way here.
DEUT|29|17|You saw among them their detestable images and idols of wood and stone, of silver and gold.
DEUT|29|18|Make sure there is no man or woman, clan or tribe among you today whose heart turns away from the LORD our God to go and worship the gods of those nations; make sure there is no root among you that produces such bitter poison.
DEUT|29|19|When such a person hears the words of this oath, he invokes a blessing on himself and therefore thinks, "I will be safe, even though I persist in going my own way." This will bring disaster on the watered land as well as the dry.
DEUT|29|20|The LORD will never be willing to forgive him; his wrath and zeal will burn against that man. All the curses written in this book will fall upon him, and the LORD will blot out his name from under heaven.
DEUT|29|21|The LORD will single him out from all the tribes of Israel for disaster, according to all the curses of the covenant written in this Book of the Law.
DEUT|29|22|Your children who follow you in later generations and foreigners who come from distant lands will see the calamities that have fallen on the land and the diseases with which the LORD has afflicted it.
DEUT|29|23|The whole land will be a burning waste of salt and sulfur-nothing planted, nothing sprouting, no vegetation growing on it. It will be like the destruction of Sodom and Gomorrah, Admah and Zeboiim, which the LORD overthrew in fierce anger.
DEUT|29|24|All the nations will ask: "Why has the LORD done this to this land? Why this fierce, burning anger?"
DEUT|29|25|And the answer will be: "It is because this people abandoned the covenant of the LORD, the God of their fathers, the covenant he made with them when he brought them out of Egypt.
DEUT|29|26|They went off and worshiped other gods and bowed down to them, gods they did not know, gods he had not given them.
DEUT|29|27|Therefore the LORD's anger burned against this land, so that he brought on it all the curses written in this book.
DEUT|29|28|In furious anger and in great wrath the LORD uprooted them from their land and thrust them into another land, as it is now."
DEUT|29|29|The secret things belong to the LORD our God, but the things revealed belong to us and to our children forever, that we may follow all the words of this law.
DEUT|30|1|When all these blessings and curses I have set before you come upon you and you take them to heart wherever the LORD your God disperses you among the nations,
DEUT|30|2|and when you and your children return to the LORD your God and obey him with all your heart and with all your soul according to everything I command you today,
DEUT|30|3|then the LORD your God will restore your fortunes and have compassion on you and gather you again from all the nations where he scattered you.
DEUT|30|4|Even if you have been banished to the most distant land under the heavens, from there the LORD your God will gather you and bring you back.
DEUT|30|5|He will bring you to the land that belonged to your fathers, and you will take possession of it. He will make you more prosperous and numerous than your fathers.
DEUT|30|6|The LORD your God will circumcise your hearts and the hearts of your descendants, so that you may love him with all your heart and with all your soul, and live.
DEUT|30|7|The LORD your God will put all these curses on your enemies who hate and persecute you.
DEUT|30|8|You will again obey the LORD and follow all his commands I am giving you today.
DEUT|30|9|Then the LORD your God will make you most prosperous in all the work of your hands and in the fruit of your womb, the young of your livestock and the crops of your land. The LORD will again delight in you and make you prosperous, just as he delighted in your fathers,
DEUT|30|10|if you obey the LORD your God and keep his commands and decrees that are written in this Book of the Law and turn to the LORD your God with all your heart and with all your soul. The Offer of Life or Death
DEUT|30|11|Now what I am commanding you today is not too difficult for you or beyond your reach.
DEUT|30|12|It is not up in heaven, so that you have to ask, "Who will ascend into heaven to get it and proclaim it to us so we may obey it?"
DEUT|30|13|Nor is it beyond the sea, so that you have to ask, "Who will cross the sea to get it and proclaim it to us so we may obey it?"
DEUT|30|14|No, the word is very near you; it is in your mouth and in your heart so you may obey it.
DEUT|30|15|See, I set before you today life and prosperity, death and destruction.
DEUT|30|16|For I command you today to love the LORD your God, to walk in his ways, and to keep his commands, decrees and laws; then you will live and increase, and the LORD your God will bless you in the land you are entering to possess.
DEUT|30|17|But if your heart turns away and you are not obedient, and if you are drawn away to bow down to other gods and worship them,
DEUT|30|18|I declare to you this day that you will certainly be destroyed. You will not live long in the land you are crossing the Jordan to enter and possess.
DEUT|30|19|This day I call heaven and earth as witnesses against you that I have set before you life and death, blessings and curses. Now choose life, so that you and your children may live
DEUT|30|20|and that you may love the LORD your God, listen to his voice, and hold fast to him. For the LORD is your life, and he will give you many years in the land he swore to give to your fathers, Abraham, Isaac and Jacob.
DEUT|31|1|Then Moses went out and spoke these words to all Israel:
DEUT|31|2|"I am now a hundred and twenty years old and I am no longer able to lead you. The LORD has said to me, 'You shall not cross the Jordan.'
DEUT|31|3|The LORD your God himself will cross over ahead of you. He will destroy these nations before you, and you will take possession of their land. Joshua also will cross over ahead of you, as the LORD said.
DEUT|31|4|And the LORD will do to them what he did to Sihon and Og, the kings of the Amorites, whom he destroyed along with their land.
DEUT|31|5|The LORD will deliver them to you, and you must do to them all that I have commanded you.
DEUT|31|6|Be strong and courageous. Do not be afraid or terrified because of them, for the LORD your God goes with you; he will never leave you nor forsake you."
DEUT|31|7|Then Moses summoned Joshua and said to him in the presence of all Israel, "Be strong and courageous, for you must go with this people into the land that the LORD swore to their forefathers to give them, and you must divide it among them as their inheritance.
DEUT|31|8|The LORD himself goes before you and will be with you; he will never leave you nor forsake you. Do not be afraid; do not be discouraged."
DEUT|31|9|So Moses wrote down this law and gave it to the priests, the sons of Levi, who carried the ark of the covenant of the LORD, and to all the elders of Israel.
DEUT|31|10|Then Moses commanded them: "At the end of every seven years, in the year for canceling debts, during the Feast of Tabernacles,
DEUT|31|11|when all Israel comes to appear before the LORD your God at the place he will choose, you shall read this law before them in their hearing.
DEUT|31|12|Assemble the people-men, women and children, and the aliens living in your towns-so they can listen and learn to fear the LORD your God and follow carefully all the words of this law.
DEUT|31|13|Their children, who do not know this law, must hear it and learn to fear the LORD your God as long as you live in the land you are crossing the Jordan to possess."
DEUT|31|14|The LORD said to Moses, "Now the day of your death is near. Call Joshua and present yourselves at the Tent of Meeting, where I will commission him." So Moses and Joshua came and presented themselves at the Tent of Meeting.
DEUT|31|15|Then the LORD appeared at the Tent in a pillar of cloud, and the cloud stood over the entrance to the Tent.
DEUT|31|16|And the LORD said to Moses: "You are going to rest with your fathers, and these people will soon prostitute themselves to the foreign gods of the land they are entering. They will forsake me and break the covenant I made with them.
DEUT|31|17|On that day I will become angry with them and forsake them; I will hide my face from them, and they will be destroyed. Many disasters and difficulties will come upon them, and on that day they will ask, 'Have not these disasters come upon us because our God is not with us?'
DEUT|31|18|And I will certainly hide my face on that day because of all their wickedness in turning to other gods.
DEUT|31|19|"Now write down for yourselves this song and teach it to the Israelites and have them sing it, so that it may be a witness for me against them.
DEUT|31|20|When I have brought them into the land flowing with milk and honey, the land I promised on oath to their forefathers, and when they eat their fill and thrive, they will turn to other gods and worship them, rejecting me and breaking my covenant.
DEUT|31|21|And when many disasters and difficulties come upon them, this song will testify against them, because it will not be forgotten by their descendants. I know what they are disposed to do, even before I bring them into the land I promised them on oath."
DEUT|31|22|So Moses wrote down this song that day and taught it to the Israelites.
DEUT|31|23|The LORD gave this command to Joshua son of Nun: "Be strong and courageous, for you will bring the Israelites into the land I promised them on oath, and I myself will be with you."
DEUT|31|24|After Moses finished writing in a book the words of this law from beginning to end,
DEUT|31|25|he gave this command to the Levites who carried the ark of the covenant of the LORD:
DEUT|31|26|"Take this Book of the Law and place it beside the ark of the covenant of the LORD your God. There it will remain as a witness against you.
DEUT|31|27|For I know how rebellious and stiff-necked you are. If you have been rebellious against the LORD while I am still alive and with you, how much more will you rebel after I die!
DEUT|31|28|Assemble before me all the elders of your tribes and all your officials, so that I can speak these words in their hearing and call heaven and earth to testify against them.
DEUT|31|29|For I know that after my death you are sure to become utterly corrupt and to turn from the way I have commanded you. In days to come, disaster will fall upon you because you will do evil in the sight of the LORD and provoke him to anger by what your hands have made."
DEUT|31|30|And Moses recited the words of this song from beginning to end in the hearing of the whole assembly of Israel:
DEUT|32|1|Listen, O heavens, and I will speak; hear, O earth, the words of my mouth.
DEUT|32|2|Let my teaching fall like rain and my words descend like dew, like showers on new grass, like abundant rain on tender plants.
DEUT|32|3|I will proclaim the name of the LORD. Oh, praise the greatness of our God!
DEUT|32|4|He is the Rock, his works are perfect, and all his ways are just. A faithful God who does no wrong, upright and just is he.
DEUT|32|5|They have acted corruptly toward him; to their shame they are no longer his children, but a warped and crooked generation.
DEUT|32|6|Is this the way you repay the LORD, O foolish and unwise people? Is he not your Father, your Creator, who made you and formed you?
DEUT|32|7|Remember the days of old; consider the generations long past. Ask your father and he will tell you, your elders, and they will explain to you.
DEUT|32|8|When the Most High gave the nations their inheritance, when he divided all mankind, he set up boundaries for the peoples according to the number of the sons of Israel.
DEUT|32|9|For the LORD's portion is his people, Jacob his allotted inheritance.
DEUT|32|10|In a desert land he found him, in a barren and howling waste. He shielded him and cared for him; he guarded him as the apple of his eye,
DEUT|32|11|like an eagle that stirs up its nest and hovers over its young, that spreads its wings to catch them and carries them on its pinions.
DEUT|32|12|The LORD alone led him; no foreign god was with him.
DEUT|32|13|He made him ride on the heights of the land and fed him with the fruit of the fields. He nourished him with honey from the rock, and with oil from the flinty crag,
DEUT|32|14|with curds and milk from herd and flock and with fattened lambs and goats, with choice rams of Bashan and the finest kernels of wheat. You drank the foaming blood of the grape.
DEUT|32|15|Jeshurun grew fat and kicked; filled with food, he became heavy and sleek. He abandoned the God who made him and rejected the Rock his Savior.
DEUT|32|16|They made him jealous with their foreign gods and angered him with their detestable idols.
DEUT|32|17|They sacrificed to demons, which are not God- gods they had not known, gods that recently appeared, gods your fathers did not fear.
DEUT|32|18|You deserted the Rock, who fathered you; you forgot the God who gave you birth.
DEUT|32|19|The LORD saw this and rejected them because he was angered by his sons and daughters.
DEUT|32|20|"I will hide my face from them," he said, "and see what their end will be; for they are a perverse generation, children who are unfaithful.
DEUT|32|21|They made me jealous by what is no god and angered me with their worthless idols. I will make them envious by those who are not a people; I will make them angry by a nation that has no understanding.
DEUT|32|22|For a fire has been kindled by my wrath, one that burns to the realm of death below. It will devour the earth and its harvests and set afire the foundations of the mountains.
DEUT|32|23|"I will heap calamities upon them and spend my arrows against them.
DEUT|32|24|I will send wasting famine against them, consuming pestilence and deadly plague; I will send against them the fangs of wild beasts, the venom of vipers that glide in the dust.
DEUT|32|25|In the street the sword will make them childless; in their homes terror will reign. Young men and young women will perish, infants and gray-haired men.
DEUT|32|26|I said I would scatter them and blot out their memory from mankind,
DEUT|32|27|but I dreaded the taunt of the enemy, lest the adversary misunderstand and say, 'Our hand has triumphed; the LORD has not done all this.'"
DEUT|32|28|They are a nation without sense, there is no discernment in them.
DEUT|32|29|If only they were wise and would understand this and discern what their end will be!
DEUT|32|30|How could one man chase a thousand, or two put ten thousand to flight, unless their Rock had sold them, unless the LORD had given them up?
DEUT|32|31|For their rock is not like our Rock, as even our enemies concede.
DEUT|32|32|Their vine comes from the vine of Sodom and from the fields of Gomorrah. Their grapes are filled with poison, and their clusters with bitterness.
DEUT|32|33|Their wine is the venom of serpents, the deadly poison of cobras.
DEUT|32|34|"Have I not kept this in reserve and sealed it in my vaults?
DEUT|32|35|It is mine to avenge; I will repay. In due time their foot will slip; their day of disaster is near and their doom rushes upon them."
DEUT|32|36|The LORD will judge his people and have compassion on his servants when he sees their strength is gone and no one is left, slave or free.
DEUT|32|37|He will say: "Now where are their gods, the rock they took refuge in,
DEUT|32|38|the gods who ate the fat of their sacrifices and drank the wine of their drink offerings? Let them rise up to help you! Let them give you shelter!
DEUT|32|39|"See now that I myself am He! There is no god besides me. I put to death and I bring to life, I have wounded and I will heal, and no one can deliver out of my hand.
DEUT|32|40|I lift my hand to heaven and declare: As surely as I live forever,
DEUT|32|41|when I sharpen my flashing sword and my hand grasps it in judgment, I will take vengeance on my adversaries and repay those who hate me.
DEUT|32|42|I will make my arrows drunk with blood, while my sword devours flesh: the blood of the slain and the captives, the heads of the enemy leaders."
DEUT|32|43|Rejoice, O nations, with his people,, for he will avenge the blood of his servants; he will take vengeance on his enemies and make atonement for his land and people.
DEUT|32|44|Moses came with Joshua son of Nun and spoke all the words of this song in the hearing of the people.
DEUT|32|45|When Moses finished reciting all these words to all Israel,
DEUT|32|46|he said to them, "Take to heart all the words I have solemnly declared to you this day, so that you may command your children to obey carefully all the words of this law.
DEUT|32|47|They are not just idle words for you-they are your life. By them you will live long in the land you are crossing the Jordan to possess."
DEUT|32|48|On that same day the LORD told Moses,
DEUT|32|49|"Go up into the Abarim Range to Mount Nebo in Moab, across from Jericho, and view Canaan, the land I am giving the Israelites as their own possession.
DEUT|32|50|There on the mountain that you have climbed you will die and be gathered to your people, just as your brother Aaron died on Mount Hor and was gathered to his people.
DEUT|32|51|This is because both of you broke faith with me in the presence of the Israelites at the waters of Meribah Kadesh in the Desert of Zin and because you did not uphold my holiness among the Israelites.
DEUT|32|52|Therefore, you will see the land only from a distance; you will not enter the land I am giving to the people of Israel."
DEUT|33|1|This is the blessing that Moses the man of God pronounced on the Israelites before his death.
DEUT|33|2|He said: "The LORD came from Sinai and dawned over them from Seir; he shone forth from Mount Paran. He came with myriads of holy ones from the south, from his mountain slopes.
DEUT|33|3|Surely it is you who love the people; all the holy ones are in your hand. At your feet they all bow down, and from you receive instruction,
DEUT|33|4|the law that Moses gave us, the possession of the assembly of Jacob.
DEUT|33|5|He was king over Jeshurun when the leaders of the people assembled, along with the tribes of Israel.
DEUT|33|6|"Let Reuben live and not die, nor his men be few."
DEUT|33|7|And this he said about Judah: "Hear, O LORD, the cry of Judah; bring him to his people. With his own hands he defends his cause. Oh, be his help against his foes!"
DEUT|33|8|About Levi he said: "Your Thummim and Urim belong to the man you favored. You tested him at Massah; you contended with him at the waters of Meribah.
DEUT|33|9|He said of his father and mother, 'I have no regard for them.' He did not recognize his brothers or acknowledge his own children, but he watched over your word and guarded your covenant.
DEUT|33|10|He teaches your precepts to Jacob and your law to Israel. He offers incense before you and whole burnt offerings on your altar.
DEUT|33|11|Bless all his skills, O LORD, and be pleased with the work of his hands. Smite the loins of those who rise up against him; strike his foes till they rise no more."
DEUT|33|12|About Benjamin he said: "Let the beloved of the LORD rest secure in him, for he shields him all day long, and the one the LORD loves rests between his shoulders."
DEUT|33|13|About Joseph he said: "May the LORD bless his land with the precious dew from heaven above and with the deep waters that lie below;
DEUT|33|14|with the best the sun brings forth and the finest the moon can yield;
DEUT|33|15|with the choicest gifts of the ancient mountains and the fruitfulness of the everlasting hills;
DEUT|33|16|with the best gifts of the earth and its fullness and the favor of him who dwelt in the burning bush. Let all these rest on the head of Joseph, on the brow of the prince among his brothers.
DEUT|33|17|In majesty he is like a firstborn bull; his horns are the horns of a wild ox. With them he will gore the nations, even those at the ends of the earth. Such are the ten thousands of Ephraim; such are the thousands of Manasseh."
DEUT|33|18|About Zebulun he said: "Rejoice, Zebulun, in your going out, and you, Issachar, in your tents.
DEUT|33|19|They will summon peoples to the mountain and there offer sacrifices of righteousness; they will feast on the abundance of the seas, on the treasures hidden in the sand."
DEUT|33|20|About Gad he said: "Blessed is he who enlarges Gad's domain! Gad lives there like a lion, tearing at arm or head.
DEUT|33|21|He chose the best land for himself; the leader's portion was kept for him. When the heads of the people assembled, he carried out the LORD's righteous will, and his judgments concerning Israel."
DEUT|33|22|About Dan he said: "Dan is a lion's cub, springing out of Bashan."
DEUT|33|23|About Naphtali he said: "Naphtali is abounding with the favor of the LORD and is full of his blessing; he will inherit southward to the lake."
DEUT|33|24|About Asher he said: "Most blessed of sons is Asher; let him be favored by his brothers, and let him bathe his feet in oil.
DEUT|33|25|The bolts of your gates will be iron and bronze, and your strength will equal your days.
DEUT|33|26|"There is no one like the God of Jeshurun, who rides on the heavens to help you and on the clouds in his majesty.
DEUT|33|27|The eternal God is your refuge, and underneath are the everlasting arms. He will drive out your enemy before you, saying, 'Destroy him!'
DEUT|33|28|So Israel will live in safety alone; Jacob's spring is secure in a land of grain and new wine, where the heavens drop dew.
DEUT|33|29|Blessed are you, O Israel! Who is like you, a people saved by the LORD? He is your shield and helper and your glorious sword. Your enemies will cower before you, and you will trample down their high places. "
DEUT|34|1|Then Moses climbed Mount Nebo from the plains of Moab to the top of Pisgah, across from Jericho. There the LORD showed him the whole land-from Gilead to Dan,
DEUT|34|2|all of Naphtali, the territory of Ephraim and Manasseh, all the land of Judah as far as the western sea,
DEUT|34|3|the Negev and the whole region from the Valley of Jericho, the City of Palms, as far as Zoar.
DEUT|34|4|Then the LORD said to him, "This is the land I promised on oath to Abraham, Isaac and Jacob when I said, 'I will give it to your descendants.' I have let you see it with your eyes, but you will not cross over into it."
DEUT|34|5|And Moses the servant of the LORD died there in Moab, as the LORD had said.
DEUT|34|6|He buried him in Moab, in the valley opposite Beth Peor, but to this day no one knows where his grave is.
DEUT|34|7|Moses was a hundred and twenty years old when he died, yet his eyes were not weak nor his strength gone.
DEUT|34|8|The Israelites grieved for Moses in the plains of Moab thirty days, until the time of weeping and mourning was over.
DEUT|34|9|Now Joshua son of Nun was filled with the spirit of wisdom because Moses had laid his hands on him. So the Israelites listened to him and did what the LORD had commanded Moses.
DEUT|34|10|Since then, no prophet has risen in Israel like Moses, whom the LORD knew face to face,
DEUT|34|11|who did all those miraculous signs and wonders the LORD sent him to do in Egypt-to Pharaoh and to all his officials and to his whole land.
DEUT|34|12|For no one has ever shown the mighty power or performed the awesome deeds that Moses did in the sight of all Israel.
