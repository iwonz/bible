GEN|1|1|В начале сотворил Бог небо и землю.
GEN|1|2|Земля же была безвидна и пуста, и тьма над бездною, и Дух Божий носился над водою.
GEN|1|3|И сказал Бог: да будет свет. И стал свет.
GEN|1|4|И увидел Бог свет, что он хорош, и отделил Бог свет от тьмы.
GEN|1|5|И назвал Бог свет днем, а тьму ночью. И был вечер, и было утро: день один.
GEN|1|6|И сказал Бог: да будет твердь посреди воды, и да отделяет она воду от воды.
GEN|1|7|И создал Бог твердь, и отделил воду, которая под твердью, от воды, которая над твердью. И стало так.
GEN|1|8|И назвал Бог твердь небом. И был вечер, и было утро: день второй.
GEN|1|9|И сказал Бог: да соберется вода, которая под небом, в одно место, и да явится суша. И стало так.
GEN|1|10|И назвал Бог сушу землею, а собрание вод назвал морями. И увидел Бог, что [это] хорошо.
GEN|1|11|И сказал Бог: да произрастит земля зелень, траву, сеющую семя дерево плодовитое, приносящее по роду своему плод, в котором семя его на земле. И стало так.
GEN|1|12|И произвела земля зелень, траву, сеющую семя по роду ее, и дерево, приносящее плод, в котором семя его по роду его. И увидел Бог, что [это] хорошо.
GEN|1|13|И был вечер, и было утро: день третий.
GEN|1|14|И сказал Бог: да будут светила на тверди небесной для отделения дня от ночи, и для знамений, и времен, и дней, и годов;
GEN|1|15|и да будут они светильниками на тверди небесной, чтобы светить на землю. И стало так.
GEN|1|16|И создал Бог два светила великие: светило большее, для управления днем, и светило меньшее, для управления ночью, и звезды;
GEN|1|17|и поставил их Бог на тверди небесной, чтобы светить на землю,
GEN|1|18|и управлять днем и ночью, и отделять свет от тьмы. И увидел Бог, что [это] хорошо.
GEN|1|19|И был вечер, и было утро: день четвертый.
GEN|1|20|И сказал Бог: да произведет вода пресмыкающихся, душу живую; и птицы да полетят над землею, по тверди небесной.
GEN|1|21|И сотворил Бог рыб больших и всякую душу животных пресмыкающихся, которых произвела вода, по роду их, и всякую птицу пернатую по роду ее. И увидел Бог, что [это] хорошо.
GEN|1|22|И благословил их Бог, говоря: плодитесь и размножайтесь, и наполняйте воды в морях, и птицы да размножаются на земле.
GEN|1|23|И был вечер, и было утро: день пятый.
GEN|1|24|И сказал Бог: да произведет земля душу живую по роду ее, скотов, и гадов, и зверей земных по роду их. И стало так.
GEN|1|25|И создал Бог зверей земных по роду их, и скот по роду его, и всех гадов земных по роду их. И увидел Бог, что [это] хорошо.
GEN|1|26|И сказал Бог: сотворим человека по образу Нашему по подобию Нашему, и да владычествуют они над рыбами морскими, и над птицами небесными, и над скотом, и над всею землею, и над всеми гадами, пресмыкающимися по земле.
GEN|1|27|И сотворил Бог человека по образу Своему, по образу Божию сотворил его; мужчину и женщину сотворил их.
GEN|1|28|И благословил их Бог, и сказал им Бог: плодитесь и размножайтесь, и наполняйте землю, и обладайте ею, и владычествуйте над рыбами морскими и над птицами небесными, и над всяким животным, пресмыкающимся по земле.
GEN|1|29|И сказал Бог: вот, Я дал вам всякую траву, сеющую семя, какая есть на всей земле, и всякое дерево, у которого плод древесный, сеющий семя; – вам [сие] будет в пищу;
GEN|1|30|а всем зверям земным, и всем птицам небесным, и всякому пресмыкающемуся по земле, в котором душа живая, [дал] Я всю зелень травную в пищу. И стало так.
GEN|1|31|И увидел Бог все, что Он создал, и вот, хорошо весьма. И был вечер, и было утро: день шестой.
GEN|2|1|Так совершены небо и земля и все воинство их.
GEN|2|2|И совершил Бог к седьмому дню дела Свои, которые Он делал, и почил в день седьмый от всех дел Своих, которые делал.
GEN|2|3|И благословил Бог седьмой день, и освятил его, ибо в оный почил от всех дел Своих, которые Бог творил и созидал.
GEN|2|4|Вот происхождение неба и земли, при сотворении их, в то время, когда Господь Бог создал землю и небо,
GEN|2|5|и всякий полевой кустарник, которого еще не было на земле, и всякую полевую траву, которая еще не росла, ибо Господь Бог не посылал дождя на землю, и не было человека для возделывания земли,
GEN|2|6|но пар поднимался с земли и орошал все лице земли.
GEN|2|7|И создал Господь Бог человека из праха земного, и вдунул в лице его дыхание жизни, и стал человек душею живою.
GEN|2|8|И насадил Господь Бог рай в Едеме на востоке, и поместил там человека, которого создал.
GEN|2|9|И произрастил Господь Бог из земли всякое дерево, приятное на вид и хорошее для пищи, и дерево жизни посреди рая, и дерево познания добра и зла.
GEN|2|10|Из Едема выходила река для орошения рая; и потом разделялась на четыре реки.
GEN|2|11|Имя одной Фисон: она обтекает всю землю Хавила, ту, где золото;
GEN|2|12|и золото той земли хорошее; там бдолах и камень оникс.
GEN|2|13|Имя второй реки Гихон: она обтекает всю землю Куш.
GEN|2|14|Имя третьей реки Хиддекель: она протекает пред Ассириею. Четвертая река Евфрат.
GEN|2|15|И взял Господь Бог человека, и поселил его в саду Едемском, чтобы возделывать его и хранить его.
GEN|2|16|И заповедал Господь Бог человеку, говоря: от всякого дерева в саду ты будешь есть,
GEN|2|17|а от дерева познания добра и зла не ешь от него, ибо в день, в который ты вкусишь от него, смертью умрешь.
GEN|2|18|И сказал Господь Бог: не хорошо быть человеку одному; сотворим ему помощника, соответственного ему.
GEN|2|19|Господь Бог образовал из земли всех животных полевых и всех птиц небесных, и привел к человеку, чтобы видеть, как он назовет их, и чтобы, как наречет человек всякую душу живую, так и было имя ей.
GEN|2|20|И нарек человек имена всем скотам и птицам небесным и всем зверям полевым; но для человека не нашлось помощника, подобного ему.
GEN|2|21|И навел Господь Бог на человека крепкий сон; и, когда он уснул, взял одно из ребр его, и закрыл то место плотию.
GEN|2|22|И создал Господь Бог из ребра, взятого у человека, жену, и привел ее к человеку.
GEN|2|23|И сказал человек: вот, это кость от костей моих и плоть от плоти моей; она будет называться женою, ибо взята от мужа.
GEN|2|24|Потому оставит человек отца своего и мать свою и прилепится к жене своей; и будут одна плоть.
GEN|2|25|И были оба наги, Адам и жена его, и не стыдились.
GEN|3|1|Змей был хитрее всех зверей полевых, которых создал Господь Бог. И сказал змей жене: подлинно ли сказал Бог: не ешьте ни от какого дерева в раю?
GEN|3|2|И сказала жена змею: плоды с дерев мы можем есть,
GEN|3|3|только плодов дерева, которое среди рая, сказал Бог, не ешьте их и не прикасайтесь к ним, чтобы вам не умереть.
GEN|3|4|И сказал змей жене: нет, не умрете,
GEN|3|5|но знает Бог, что в день, в который вы вкусите их, откроются глаза ваши, и вы будете, как боги, знающие добро и зло.
GEN|3|6|И увидела жена, что дерево хорошо для пищи, и что оно приятно для глаз и вожделенно, потому что дает знание; и взяла плодов его и ела; и дала также мужу своему, и он ел.
GEN|3|7|И открылись глаза у них обоих, и узнали они, что наги, и сшили смоковные листья, и сделали себе опоясания.
GEN|3|8|И услышали голос Господа Бога, ходящего в раю во время прохлады дня; и скрылся Адам и жена его от лица Господа Бога между деревьями рая.
GEN|3|9|И воззвал Господь Бог к Адаму и сказал ему: где ты?
GEN|3|10|Он сказал: голос Твой я услышал в раю, и убоялся, потому что я наг, и скрылся.
GEN|3|11|И сказал: кто сказал тебе, что ты наг? не ел ли ты от дерева, с которого Я запретил тебе есть?
GEN|3|12|Адам сказал: жена, которую Ты мне дал, она дала мне от дерева, и я ел.
GEN|3|13|И сказал Господь Бог жене: что ты это сделала? Жена сказала: змей обольстил меня, и я ела.
GEN|3|14|И сказал Господь Бог змею: за то, что ты сделал это, проклят ты пред всеми скотами и пред всеми зверями полевыми; ты будешь ходить на чреве твоем, и будешь есть прах во все дни жизни твоей;
GEN|3|15|и вражду положу между тобою и между женою, и между семенем твоим и между семенем ее; оно будет поражать тебя в голову, а ты будешь жалить его в пяту.
GEN|3|16|Жене сказал: умножая умножу скорбь твою в беременности твоей; в болезни будешь рождать детей; и к мужу твоему влечение твое, и он будет господствовать над тобою.
GEN|3|17|Адаму же сказал: за то, что ты послушал голоса жены твоей и ел от дерева, о котором Я заповедал тебе, сказав: не ешь от него, проклята земля за тебя; со скорбью будешь питаться от нее во все дни жизни твоей;
GEN|3|18|терния и волчцы произрастит она тебе; и будешь питаться полевою травою;
GEN|3|19|в поте лица твоего будешь есть хлеб, доколе не возвратишься в землю, из которой ты взят, ибо прах ты и в прах возвратишься.
GEN|3|20|И нарек Адам имя жене своей: Ева, ибо она стала матерью всех живущих.
GEN|3|21|И сделал Господь Бог Адаму и жене его одежды кожаные и одел их.
GEN|3|22|И сказал Господь Бог: вот, Адам стал как один из Нас, зная добро и зло; и теперь как бы не простер он руки своей, и не взял также от дерева жизни, и не вкусил, и не стал жить вечно.
GEN|3|23|И выслал его Господь Бог из сада Едемского, чтобы возделывать землю, из которой он взят.
GEN|3|24|И изгнал Адама, и поставил на востоке у сада Едемского Херувима и пламенный меч обращающийся, чтобы охранять путь к дереву жизни.
GEN|4|1|Адам познал Еву, жену свою; и она зачала, и родила Каина, и сказала: приобрела я человека от Господа.
GEN|4|2|И еще родила брата его, Авеля. И был Авель пастырь овец, а Каин был земледелец.
GEN|4|3|Спустя несколько времени, Каин принес от плодов земли дар Господу,
GEN|4|4|и Авель также принес от первородных стада своего и от тука их. И призрел Господь на Авеля и на дар его,
GEN|4|5|а на Каина и на дар его не призрел. Каин сильно огорчился, и поникло лице его.
GEN|4|6|И сказал Господь Каину: почему ты огорчился? и отчего поникло лице твое?
GEN|4|7|если делаешь доброе, то не поднимаешь ли лица? а если не делаешь доброго, то у дверей грех лежит; он влечет тебя к себе, но ты господствуй над ним.
GEN|4|8|И сказал Каин Авелю, брату своему. И когда они были в поле, восстал Каин на Авеля, брата своего, и убил его.
GEN|4|9|И сказал Господь Каину: где Авель, брат твой? Он сказал: не знаю; разве я сторож брату моему?
GEN|4|10|И сказал: что ты сделал? голос крови брата твоего вопиет ко Мне от земли;
GEN|4|11|и ныне проклят ты от земли, которая отверзла уста свои принять кровь брата твоего от руки твоей;
GEN|4|12|когда ты будешь возделывать землю, она не станет более давать силы своей для тебя; ты будешь изгнанником и скитальцем на земле.
GEN|4|13|И сказал Каин Господу: наказание мое больше, нежели снести можно;
GEN|4|14|вот, Ты теперь сгоняешь меня с лица земли, и от лица Твоего я скроюсь, и буду изгнанником и скитальцем на земле; и всякий, кто встретится со мною, убьет меня.
GEN|4|15|И сказал ему Господь: за то всякому, кто убьет Каина, отмстится всемеро. И сделал Господь Каину знамение, чтобы никто, встретившись с ним, не убил его.
GEN|4|16|И пошел Каин от лица Господня и поселился в земле Нод, на восток от Едема.
GEN|4|17|И познал Каин жену свою; и она зачала и родила Еноха. И построил он город; и назвал город по имени сына своего: Енох.
GEN|4|18|У Еноха родился Ирад; Ирад родил Мехиаеля; Мехиаель родил Мафусала; Мафусал родил Ламеха.
GEN|4|19|И взял себе Ламех две жены: имя одной: Ада, и имя второй: Цилла.
GEN|4|20|Ада родила Иавала: он был отец живущих в шатрах со стадами.
GEN|4|21|Имя брату его Иувал: он был отец всех играющих на гуслях и свирели.
GEN|4|22|Цилла также родила Тувалкаина, который был ковачом всех орудий из меди и железа. И сестра Тувалкаина Ноема.
GEN|4|23|И сказал Ламех женам своим: Ада и Цилла! послушайте голоса моего; жены Ламеховы! внимайте словам моим: я убил мужа в язву мне и отрока в рану мне;
GEN|4|24|если за Каина отмстится всемеро, то за Ламеха в семьдесят раз всемеро.
GEN|4|25|И познал Адам еще жену свою, и она родила сына, и нарекла ему имя: Сиф, потому что, [говорила она], Бог положил мне другое семя, вместо Авеля, которого убил Каин.
GEN|4|26|У Сифа также родился сын, и он нарек ему имя: Енос; тогда начали призывать имя Господа.
GEN|5|1|Вот родословие Адама: когда Бог сотворил человека, по подобию Божию создал его,
GEN|5|2|мужчину и женщину сотворил их, и благословил их, и нарек им имя: человек, в день сотворения их.
GEN|5|3|Адам жил сто тридцать лет и родил [сына] по подобию своему по образу своему, и нарек ему имя: Сиф.
GEN|5|4|Дней Адама по рождении им Сифа было восемьсот лет, и родил он сынов и дочерей.
GEN|5|5|Всех же дней жизни Адамовой было девятьсот тридцать лет; и он умер.
GEN|5|6|Сиф жил сто пять лет и родил Еноса.
GEN|5|7|По рождении Еноса Сиф жил восемьсот семь лет и родил сынов и дочерей.
GEN|5|8|Всех же дней Сифовых было девятьсот двенадцать лет; и он умер.
GEN|5|9|Енос жил девяносто лет и родил Каинана.
GEN|5|10|По рождении Каинана Енос жил восемьсот пятнадцать лет и родил сынов и дочерей.
GEN|5|11|Всех же дней Еноса было девятьсот пять лет; и он умер.
GEN|5|12|Каинан жил семьдесят лет и родил Малелеила.
GEN|5|13|По рождении Малелеила Каинан жил восемьсот сорок лет и родил сынов и дочерей.
GEN|5|14|Всех же дней Каинана было девятьсот десять лет; и он умер.
GEN|5|15|Малелеил жил шестьдесят пять лет и родил Иареда.
GEN|5|16|По рождении Иареда Малелеил жил восемьсот тридцать лет и родил сынов и дочерей.
GEN|5|17|Всех же дней Малелеила было восемьсот девяносто пять лет; и он умер.
GEN|5|18|Иаред жил сто шестьдесят два года и родил Еноха.
GEN|5|19|По рождении Еноха Иаред жил восемьсот лет и родил сынов и дочерей.
GEN|5|20|Всех же дней Иареда было девятьсот шестьдесят два года; и он умер.
GEN|5|21|Енох жил шестьдесят пять лет и родил Мафусала.
GEN|5|22|И ходил Енох пред Богом, по рождении Мафусала, триста лет и родил сынов и дочерей.
GEN|5|23|Всех же дней Еноха было триста шестьдесят пять лет.
GEN|5|24|И ходил Енох пред Богом; и не стало его, потому что Бог взял его.
GEN|5|25|Мафусал жил сто восемьдесят семь лет и родил Ламеха.
GEN|5|26|По рождении Ламеха Мафусал жил семьсот восемьдесят два года и родил сынов и дочерей.
GEN|5|27|Всех же дней Мафусала было девятьсот шестьдесят девять лет; и он умер.
GEN|5|28|Ламех жил сто восемьдесят два года и родил сына,
GEN|5|29|и нарек ему имя: Ной, сказав: он утешит нас в работе нашей и в трудах рук наших при [возделывании] земли, которую проклял Господь.
GEN|5|30|И жил Ламех по рождении Ноя пятьсот девяносто пять лет и родил сынов и дочерей.
GEN|5|31|Всех же дней Ламеха было семьсот семьдесят семь лет; и он умер.
GEN|5|32|Ною было пятьсот лет и родил Ной Сима, Хама и Иафета.
GEN|6|1|Когда люди начали умножаться на земле и родились у них дочери,
GEN|6|2|тогда сыны Божии увидели дочерей человеческих, что они красивы, и брали [их] себе в жены, какую кто избрал.
GEN|6|3|И сказал Господь: не вечно Духу Моему быть пренебрегаемым человеками; потому что они плоть; пусть будут дни их сто двадцать лет.
GEN|6|4|В то время были на земле исполины, особенно же с того времени, как сыны Божии стали входить к дочерям человеческим, и они стали рождать им: это сильные, издревле славные люди.
GEN|6|5|И увидел Господь, что велико развращение человеков на земле, и что все мысли и помышления сердца их были зло во всякое время;
GEN|6|6|и раскаялся Господь, что создал человека на земле, и восскорбел в сердце Своем.
GEN|6|7|И сказал Господь: истреблю с лица земли человеков, которых Я сотворил, от человека до скотов, и гадов и птиц небесных истреблю, ибо Я раскаялся, что создал их.
GEN|6|8|Ной же обрел благодать пред очами Господа.
GEN|6|9|Вот житие Ноя: Ной был человек праведный и непорочный в роде своем; Ной ходил пред Богом.
GEN|6|10|Ной родил трех сынов: Сима, Хама и Иафета.
GEN|6|11|Но земля растлилась пред лицем Божиим, и наполнилась земля злодеяниями.
GEN|6|12|И воззрел Бог на землю, и вот, она растленна, ибо всякая плоть извратила путь свой на земле.
GEN|6|13|И сказал Бог Ною: конец всякой плоти пришел пред лице Мое, ибо земля наполнилась от них злодеяниями; и вот, Я истреблю их с земли.
GEN|6|14|Сделай себе ковчег из дерева гофер; отделения сделай в ковчеге и осмоли его смолою внутри и снаружи.
GEN|6|15|И сделай его так: длина ковчега триста локтей; ширина его пятьдесят локтей, а высота его тридцать локтей.
GEN|6|16|И сделай отверстие в ковчеге, и в локоть сведи его вверху, и дверь в ковчег сделай с боку его; устрой в нем нижнее, второе и третье [жилье].
GEN|6|17|И вот, Я наведу на землю потоп водный, чтоб истребить всякую плоть, в которой есть дух жизни, под небесами; все, что есть на земле, лишится жизни.
GEN|6|18|Но с тобою Я поставлю завет Мой, и войдешь в ковчег ты, и сыновья твои, и жена твоя, и жены сынов твоих с тобою.
GEN|6|19|Введи также в ковчег из всех животных, и от всякой плоти по паре, чтоб они остались с тобою в живых; мужеского пола и женского пусть они будут.
GEN|6|20|Из птиц по роду их, и из скотов по роду их, и из всех пресмыкающихся по земле по роду их, из всех по паре войдут к тебе, чтобы остались в живых.
GEN|6|21|Ты же возьми себе всякой пищи, какою питаются, и собери к себе; и будет она для тебя и для них пищею.
GEN|6|22|И сделал Ной все: как повелел ему Бог, так он и сделал.
GEN|7|1|И сказал Господь Ною: войди ты и все семейство твое в ковчег, ибо тебя увидел Я праведным предо Мною в роде сем;
GEN|7|2|и всякого скота чистого возьми по семи, мужеского пола и женского, а из скота нечистого по два, мужеского пола и женского;
GEN|7|3|также и из птиц небесных по семи, мужеского пола и женского, чтобы сохранить племя для всей земли,
GEN|7|4|ибо чрез семь дней Я буду изливать дождь на землю сорок дней и сорок ночей; и истреблю все существующее, что Я создал, с лица земли.
GEN|7|5|Ной сделал все, что Господь повелел ему.
GEN|7|6|Ной же был шестисот лет, как потоп водный пришел на землю.
GEN|7|7|И вошел Ной и сыновья его, и жена его, и жены сынов его с ним в ковчег от вод потопа.
GEN|7|8|И из скотов чистых и из скотов нечистых, и из всех пресмыкающихся по земле
GEN|7|9|по паре, мужеского пола и женского, вошли к Ною в ковчег, как Бог повелел Ною.
GEN|7|10|Чрез семь дней воды потопа пришли на землю.
GEN|7|11|В шестисотый год жизни Ноевой, во второй месяц, в семнадцатый день месяца, в сей день разверзлись все источники великой бездны, и окна небесные отворились;
GEN|7|12|и лился на землю дождь сорок дней и сорок ночей.
GEN|7|13|В сей самый день вошел в ковчег Ной, и Сим, Хам и Иафет, сыновья Ноевы, и жена Ноева, и три жены сынов его с ними.
GEN|7|14|Они, и все звери по роду их, и всякий скот по роду его, и все гады, пресмыкающиеся по земле, по роду их, и все летающие по роду их, все птицы, все крылатые,
GEN|7|15|и вошли к Ною в ковчег по паре от всякой плоти, в которой есть дух жизни;
GEN|7|16|и вошедшие мужеский и женский пол всякой плоти вошли, как повелел ему Бог. И затворил Господь за ним.
GEN|7|17|И продолжалось на земле наводнение сорок дней, и умножилась вода, и подняла ковчег, и он возвысился над землею;
GEN|7|18|вода же усиливалась и весьма умножалась на земле, и ковчег плавал по поверхности вод.
GEN|7|19|И усилилась вода на земле чрезвычайно, так что покрылись все высокие горы, какие есть под всем небом;
GEN|7|20|на пятнадцать локтей поднялась над ними вода, и покрылись горы.
GEN|7|21|И лишилась жизни всякая плоть, движущаяся по земле, и птицы, и скоты, и звери, и все гады, ползающие по земле, и все люди;
GEN|7|22|все, что имело дыхание духа жизни в ноздрях своих на суше, умерло.
GEN|7|23|Истребилось всякое существо, которое было на поверхности земли; от человека до скота, и гадов, и птиц небесных, – все истребилось с земли, остался только Ной и что [было] с ним в ковчеге.
GEN|7|24|Вода же усиливалась на земле сто пятьдесят дней.
GEN|8|1|И вспомнил Бог о Ное, и о всех зверях, и о всех скотах, (и о всех птицах, и о всех гадах пресмыкающихся,) бывших с ним в ковчеге; и навел Бог ветер на землю, и воды остановились.
GEN|8|2|И закрылись источники бездны и окна небесные, и перестал дождь с неба.
GEN|8|3|Вода же постепенно возвращалась с земли, и стала убывать вода по окончании ста пятидесяти дней.
GEN|8|4|И остановился ковчег в седьмом месяце, в семнадцатый день месяца, на горах Араратских.
GEN|8|5|Вода постоянно убывала до десятого месяца; в первый день десятого месяца показались верхи гор.
GEN|8|6|По прошествии сорока дней Ной открыл сделанное им окно ковчега
GEN|8|7|и выпустил ворона, который, вылетев, отлетал и прилетал, пока осушилась земля от воды.
GEN|8|8|Потом выпустил от себя голубя, чтобы видеть, сошла ли вода с лица земли,
GEN|8|9|но голубь не нашел места покоя для ног своих и возвратился к нему в ковчег, ибо вода была еще на поверхности всей земли; и он простер руку свою, и взял его, и принял к себе в ковчег.
GEN|8|10|И помедлил еще семь дней других и опять выпустил голубя из ковчега.
GEN|8|11|Голубь возвратился к нему в вечернее время, и вот, свежий масличный лист во рту у него, и Ной узнал, что вода сошла с земли.
GEN|8|12|Он помедлил еще семь дней других и выпустил голубя; и он уже не возвратился к нему.
GEN|8|13|Шестьсот первого года к первому [дню] первого месяца иссякла вода на земле; и открыл Ной кровлю ковчега и посмотрел, и вот, обсохла поверхность земли.
GEN|8|14|И во втором месяце, к двадцать седьмому дню месяца, земля высохла.
GEN|8|15|И сказал Бог Ною:
GEN|8|16|выйди из ковчега ты и жена твоя, и сыновья твои, и жены сынов твоих с тобою;
GEN|8|17|выведи с собою всех животных, которые с тобою, от всякой плоти, из птиц, и скотов, и всех гадов, пресмыкающихся по земле: пусть разойдутся они по земле, и пусть плодятся и размножаются на земле.
GEN|8|18|И вышел Ной и сыновья его, и жена его, и жены сынов его с ним;
GEN|8|19|все звери, и все гады, и все птицы, все движущееся по земле, по родам своим, вышли из ковчега.
GEN|8|20|И устроил Ной жертвенник Господу; и взял из всякого скота чистого и из всех птиц чистых и принес во всесожжение на жертвеннике.
GEN|8|21|И обонял Господь приятное благоухание, и сказал Господь в сердце Своем: не буду больше проклинать землю за человека, потому что помышление сердца человеческого – зло от юности его; и не буду больше поражать всего живущего, как Я сделал:
GEN|8|22|впредь во все дни земли сеяние и жатва, холод и зной, лето и зима, день и ночь не прекратятся.
GEN|9|1|И благословил Бог Ноя и сынов его и сказал им: плодитесь и размножайтесь, и наполняйте землю.
GEN|9|2|да страшатся и да трепещут вас все звери земные, и все птицы небесные, все, что движется на земле, и все рыбы морские: в ваши руки отданы они;
GEN|9|3|все движущееся, что живет, будет вам в пищу; как зелень травную даю вам все;
GEN|9|4|только плоти с душею ее, с кровью ее, не ешьте;
GEN|9|5|Я взыщу и вашу кровь, [в которой] жизнь ваша, взыщу ее от всякого зверя, взыщу также душу человека от руки человека, от руки брата его;
GEN|9|6|кто прольет кровь человеческую, того кровь прольется рукою человека: ибо человек создан по образу Божию;
GEN|9|7|вы же плодитесь и размножайтесь, и распространяйтесь по земле, и умножайтесь на ней.
GEN|9|8|И сказал Бог Ною и сынам его с ним:
GEN|9|9|вот, Я поставляю завет Мой с вами и с потомством вашим после вас,
GEN|9|10|и со всякою душею живою, которая с вами, с птицами и со скотами, и со всеми зверями земными, которые у вас, со всеми вышедшими из ковчега, со всеми животными земными;
GEN|9|11|поставляю завет Мой с вами, что не будет более истреблена всякая плоть водами потопа, и не будет уже потопа на опустошение земли.
GEN|9|12|И сказал Бог: вот знамение завета, который Я поставляю между Мною и между вами и между всякою душею живою, которая с вами, в роды навсегда:
GEN|9|13|Я полагаю радугу Мою в облаке, чтоб она была знамением завета между Мною и между землею.
GEN|9|14|И будет, когда Я наведу облако на землю, то явится радуга в облаке;
GEN|9|15|и Я вспомню завет Мой, который между Мною и между вами и между всякою душею живою во всякой плоти; и не будет более вода потопом на истребление всякой плоти.
GEN|9|16|И будет радуга в облаке, и Я увижу ее, и вспомню завет вечный между Богом и между всякою душею живою во всякой плоти, которая на земле.
GEN|9|17|И сказал Бог Ною: вот знамение завета, который Я поставил между Мною и между всякою плотью, которая на земле.
GEN|9|18|Сыновья Ноя, вышедшие из ковчега, были: Сим, Хам и Иафет. Хам же был отец Ханаана.
GEN|9|19|Сии трое были сыновья Ноевы, и от них населилась вся земля.
GEN|9|20|Ной начал возделывать землю и насадил виноградник;
GEN|9|21|и выпил он вина, и опьянел, и [лежал] обнаженным в шатре своем.
GEN|9|22|И увидел Хам, отец Ханаана, наготу отца своего, и выйдя рассказал двум братьям своим.
GEN|9|23|Сим же и Иафет взяли одежду и, положив ее на плечи свои, пошли задом и покрыли наготу отца своего; лица их были обращены назад, и они не видали наготы отца своего.
GEN|9|24|Ной проспался от вина своего и узнал, что сделал над ним меньший сын его,
GEN|9|25|и сказал: проклят Ханаан; раб рабов будет он у братьев своих.
GEN|9|26|Потом сказал: благословен Господь Бог Симов; Ханаан же будет рабом ему;
GEN|9|27|да распространит Бог Иафета, и да вселится он в шатрах Симовых; Ханаан же будет рабом ему.
GEN|9|28|И жил Ной после потопа триста пятьдесят лет.
GEN|9|29|Всех же дней Ноевых было девятьсот пятьдесят лет, и он умер.
GEN|10|1|Вот родословие сынов Ноевых: Сима, Хама и Иафета. После потопа родились у них дети.
GEN|10|2|Сыны Иафета: Гомер, Магог, Мадай, Иаван, Фувал, Мешех и Фирас.
GEN|10|3|Сыны Гомера: Аскеназ, Рифат и Фогарма.
GEN|10|4|Сыны Иавана: Елиса, Фарсис, Киттим и Доданим.
GEN|10|5|От сих населились острова народов в землях их, каждый по языку своему, по племенам своим, в народах своих.
GEN|10|6|Сыны Хама: Хуш, Мицраим, Фут и Ханаан.
GEN|10|7|Сыны Хуша: Сева, Хавила, Савта, Раама и Савтеха. Сыны Раамы: Шева и Дедан.
GEN|10|8|Хуш родил также Нимрода: сей начал быть силен на земле.
GEN|10|9|Он был сильный зверолов пред Господом; потому и говориться: сильный зверолов, как Нимрод, пред Господом.
GEN|10|10|Царство его вначале составляли: Вавилон, Эрех, Аккад и Халне, в земле Сеннаар.
GEN|10|11|Из сей земли вышел Ассур, и построил Ниневию, Реховофир, Калах.
GEN|10|12|И Ресен между Ниневию и между Калахом; это город великий.
GEN|10|13|От Мицраима произошли Лудим, Анамим, Легавим, Нафтухим,
GEN|10|14|Патрусим, Каслухим, откуда вышли Филистимляне, и Кафторим.
GEN|10|15|От Ханаана родились: Сидон, первенец его, Хет,
GEN|10|16|Иевусей, Аморей, Гергесей,
GEN|10|17|Евей, Аркей, Синей,
GEN|10|18|Арвадей, Цемарей и Химарей. В последствии племена Ханаанские рассеялись.
GEN|10|19|И были пределы Хананеев от Сидона к Герару до Газы, отсюда к Садому, Гаморре, Адме и Цевоиму до Лаши.
GEN|10|20|Это сыны Хамовы, по племенам их, по языкам их, в землях их, в народах их.
GEN|10|21|Были дети и у Сима, отца всех сынов Еверовых, старшего брата Иафетова.
GEN|10|22|Сыны Сима: Елам, Асур, Арфаксад, Луд, Арам.
GEN|10|23|Сыны Арама: Уц, Хул, Гефер и Маш.
GEN|10|24|Арфаксад родил Салу, Сала родил Евера.
GEN|10|25|У Евера родились два сына; имя одному: Фалек, потому что во дни его земля разделена; имя брата его: Иоктан.
GEN|10|26|Иоктан родил Алмодада, Шалефа, Хацармавефа, Иераха,
GEN|10|27|Гадорама, Узала, Диклу,
GEN|10|28|Овала, Авимаила, Шеву,
GEN|10|29|Офира, Хавилу и Иовава. Все эти сыновья Иоктана.
GEN|10|30|Поселения их были от Меши до Сефара, горы восточной.
GEN|10|31|Это сыновья Симовы по племенам их, по языкам их, в землях их, по народам их.
GEN|10|32|Вот племена сынов Ноевых, по родословию их, в народах их. От них распространились народы по земле после потопа.
GEN|11|1|На всей земле был один язык и одно наречие.
GEN|11|2|Двинувшись с востока, они нашли в земле Сеннаар равнину и поселились там.
GEN|11|3|И сказали друг другу: наделаем кирпичей и обожжем огнем. И стали у них кирпичи вместо камней, а земляная смола вместо извести.
GEN|11|4|И сказали они: построим себе город и башню, высотою до небес, и сделаем себе имя, прежде нежели рассеемся по лицу всей земли.
GEN|11|5|И сошел Господь посмотреть город и башню, которые строили сыны человеческие.
GEN|11|6|И сказал Господь: вот, один народ, и один у всех язык; и вот что начали они делать, и не отстанут они от того, что задумали делать;
GEN|11|7|сойдем же и смешаем там язык их, так чтобы один не понимал речи другого.
GEN|11|8|И рассеял их Господь оттуда по всей земле; и они перестали строить город.
GEN|11|9|Посему дано ему имя: Вавилон, ибо там смешал Господь язык всей земли, и оттуда рассеял их Господь по всей земле.
GEN|11|10|Вот родословие Сима: Сим был ста лет и родил Арфаксада, чрез два года после потопа;
GEN|11|11|по рождении Арфаксада Сим жил пятьсот лет и родил сынов и дочерей.
GEN|11|12|Арфаксад жил тридцать пять лет и родил Салу.
GEN|11|13|По рождении Салы Арфаксад жил четыреста три года и родил сынов и дочерей.
GEN|11|14|Сала жил тридцать лет и родил Евера.
GEN|11|15|По рождении Евера Сала жил четыреста три года и родил сынов и дочерей.
GEN|11|16|Евер жил тридцать четыре года и родил Фалека.
GEN|11|17|По рождении Фалека Евер жил четыреста тридцать лет и родил сынов и дочерей.
GEN|11|18|Фалек жил тридцать лет и родил Рагава.
GEN|11|19|По рождении Рагава Фалек жил двести девять лет и родил сынов и дочерей.
GEN|11|20|Рагав жил тридцать два года и родил Серуха.
GEN|11|21|По рождении Серуха Рагав жил двести семь лет и родил сынов и дочерей.
GEN|11|22|Серух жил тридцать лет и родил Нахора.
GEN|11|23|По рождении Нахора Серух жил двести лет и родил сынов и дочерей.
GEN|11|24|Нахор жил двадцать девять лет и родил Фарру.
GEN|11|25|По рождении Фарры Нахор жил сто девятнадцать лет и родил сынов и дочерей.
GEN|11|26|Фарра жил семьдесят лет и родил Аврама, Нахора и Арана.
GEN|11|27|Вот родословие Фарры: Фарра родил Аврама, Нахора и Арана. Аран родил Лота.
GEN|11|28|И умер Аран при Фарре, отце своем, в земле рождения своего, в Уре Халдейском.
GEN|11|29|Аврам и Нахор взяли себе жен; имя жены Аврамовой: Сара; имя жены Нахоровой: Милка, дочь Арана, отца Милки и отца Иски.
GEN|11|30|И Сара была неплодна и бездетна.
GEN|11|31|И взял Фарра Аврама, сына своего, и Лота, сына Аранова, внука своего, и Сару, невестку свою, жену Аврама, сына своего, и вышел с ними из Ура Халдейского, чтобы идти в землю Ханаанскую; но, дойдя до Харрана, они остановились там.
GEN|11|32|И было дней [жизни] Фарры двести пять лет, и умер Фарра в Харране.
GEN|12|1|И сказал Господь Авраму: пойди из земли твоей, от родства твоего и из дома отца твоего, в землю, которую Я укажу тебе;
GEN|12|2|и Я произведу от тебя великий народ, и благословлю тебя, и возвеличу имя твое, и будешь ты в благословение;
GEN|12|3|Я благословлю благословляющих тебя, и злословящих тебя прокляну; и благословятся в тебе все племена земные.
GEN|12|4|И пошел Аврам, как сказал ему Господь; и с ним пошел Лот. Аврам был семидесяти пяти лет, когда вышел из Харрана.
GEN|12|5|И взял Аврам с собою Сару, жену свою, Лота, сына брата своего, и все имение, которое они приобрели, и всех людей, которых они имели в Харране; и вышли, чтобы идти в землю Ханаанскую; и пришли в землю Ханаанскую.
GEN|12|6|И прошел Аврам по земле сей до места Сихема, до дубравы Море. В этой земле тогда [жили] Хананеи.
GEN|12|7|И явился Господь Авраму и сказал: потомству твоему отдам Я землю сию. И создал [он] там жертвенник Господу, Который явился ему.
GEN|12|8|Оттуда двинулся он к горе, на восток от Вефиля; и поставил шатер свой [так, что от него] Вефиль [был] на запад, а Гай на восток; и создал там жертвенник Господу и призвал имя Господа.
GEN|12|9|И поднялся Аврам и продолжал идти к югу.
GEN|12|10|И был голод в той земле. И сошел Аврам в Египет, пожить там, потому что усилился голод в земле той.
GEN|12|11|Когда же он приближался к Египту, то сказал Саре, жене своей: вот, я знаю, что ты женщина, прекрасная видом;
GEN|12|12|и когда Египтяне увидят тебя, то скажут: это жена его; и убьют меня, а тебя оставят в живых;
GEN|12|13|скажи же, что ты мне сестра, дабы мне хорошо было ради тебя, и дабы жива была душа моя чрез тебя.
GEN|12|14|И было, когда пришел Аврам в Египет, Египтяне увидели, что она женщина весьма красивая;
GEN|12|15|увидели ее и вельможи фараоновы и похвалили ее фараону; и взята была она в дом фараонов.
GEN|12|16|И Авраму хорошо было ради ее; и был у него мелкий и крупный скот и ослы, и рабы и рабыни, и лошаки и верблюды.
GEN|12|17|Но Господь поразил тяжкими ударами фараона и дом его за Сару, жену Аврамову.
GEN|12|18|И призвал фараон Аврама и сказал: что ты это сделал со мною? для чего не сказал мне, что она жена твоя?
GEN|12|19|для чего ты сказал: она сестра моя? и я взял было ее себе в жену. И теперь вот жена твоя; возьми и пойди.
GEN|12|20|И дал о нем фараон повеление людям, и проводили его, и жену его, и все, что у него было.
GEN|13|1|И поднялся Аврам из Египта, сам и жена его, и все, что у него было, и Лот с ним, на юг.
GEN|13|2|И был Аврам очень богат скотом, и серебром, и золотом.
GEN|13|3|И продолжал он переходы свои от юга до Вефиля, до места, где прежде был шатер его между Вефилем и между Гаем,
GEN|13|4|до места жертвенника, который он сделал там вначале; и там призвал Аврам имя Господа.
GEN|13|5|И у Лота, который ходил с Аврамом, также был мелкий и крупный скот и шатры.
GEN|13|6|И непоместительна была земля для них, чтобы жить вместе, ибо имущество их было так велико, что они не могли жить вместе.
GEN|13|7|И был спор между пастухами скота Аврамова и между пастухами скота Лотова; и Хананеи и Ферезеи жили тогда в той земле.
GEN|13|8|И сказал Аврам Лоту: да не будет раздора между мною и тобою, и между пастухами моими и пастухами твоими, ибо мы родственники;
GEN|13|9|не вся ли земля пред тобою? отделись же от меня: если ты налево, то я направо; а если ты направо, то я налево.
GEN|13|10|Лот возвел очи свои и увидел всю окрестность Иорданскую, что она, прежде нежели истребил Господь Содом и Гоморру, вся до Сигора орошалась водою, как сад Господень, как земля Египетская;
GEN|13|11|и избрал себе Лот всю окрестность Иорданскую; и двинулся Лот к востоку. И отделились они друг от друга.
GEN|13|12|Аврам стал жить на земле Ханаанской; а Лот стал жить в городах окрестности и раскинул шатры до Содома.
GEN|13|13|Жители же Содомские были злы и весьма грешны пред Господом.
GEN|13|14|И сказал Господь Авраму, после того как Лот отделился от него: возведи очи твои и с места, на котором ты теперь, посмотри к северу и к югу, и к востоку и к западу;
GEN|13|15|ибо всю землю, которую ты видишь, тебе дам Я и потомству твоему навеки,
GEN|13|16|и сделаю потомство твое, как песок земной; если кто может сосчитать песок земной, то и потомство твое сочтено будет;
GEN|13|17|встань, пройди по земле сей в долготу и в широту ее, ибо Я тебе дам ее.
GEN|13|18|И двинул Аврам шатер, и пошел, и поселился у дубравы Мамре, что в Хевроне; и создал там жертвенник Господу.
GEN|14|1|И было во дни Амрафела, царя Сеннаарского, Ариоха, царя Елласарского, Кедорлаомера, царя Еламского, и Фидала, царя Гоимского,
GEN|14|2|пошли они войною против Беры, царя Содомского, против Бирши, царя Гоморрского, Шинава, царя Адмы, Шемевера, царя Севоимского, и против царя Белы, которая есть Сигор.
GEN|14|3|Все сии соединились в долине Сиддим, где [ныне] море Соленое.
GEN|14|4|Двенадцать лет были они в порабощении у Кедорлаомера, а в тринадцатом году возмутились.
GEN|14|5|В четырнадцатом году пришел Кедорлаомер и цари, которые с ним, и поразили Рефаимов в Аштероф–Карнаиме, Зузимов в Гаме, Эмимов в Шаве–Кириафаиме,
GEN|14|6|и Хорреев в горе их Сеире, до Эл–Фарана, что при пустыне.
GEN|14|7|И возвратившись оттуда, они пришли к источнику Мишпат, который есть Кадес, и поразили всю страну Амаликитян, и также Аморреев, живущих в Хацацон–Фамаре.
GEN|14|8|И вышли царь Содомский, царь Гоморрский, царь Адмы, царь Севоимский и царь Белы, которая есть Сигор; и вступили в сражение с ними в долине Сиддим,
GEN|14|9|с Кедорлаомером, царем Еламским, Фидалом, царем Гоимским, Амрафелом, царем Сеннаарским, Ариохом, царем Елласарским, – четыре царя против пяти.
GEN|14|10|В долине же Сиддим было много смоляных ям. И цари Содомский и Гоморрский, обратившись в бегство, упали в них, а остальные убежали в горы.
GEN|14|11|[Победители] взяли все имущество Содома и Гоморры и весь запас их и ушли.
GEN|14|12|И взяли Лота, племянника Аврамова, жившего в Содоме, и имущество его и ушли.
GEN|14|13|И пришел один из уцелевших и известил Аврама Еврея, жившего тогда у дубравы Мамре, Аморреянина, брата Эшколу и брата Анеру, которые были союзники Аврамовы.
GEN|14|14|Аврам, услышав, что сродник его взят в плен, вооружил рабов своих, рожденных в доме его, триста восемнадцать, и преследовал [неприятелей] до Дана;
GEN|14|15|и, разделившись, [напал] на них ночью, сам и рабы его, и поразил их, и преследовал их до Ховы, что по левую сторону Дамаска;
GEN|14|16|и возвратил все имущество и Лота, сродника своего, и имущество его возвратил, также и женщин и народ.
GEN|14|17|Когда он возвращался после поражения Кедорлаомера и царей, бывших с ним, царь Содомский вышел ему навстречу в долину Шаве, что [ныне] долина царская;
GEN|14|18|и Мелхиседек, царь Салимский, вынес хлеб и вино, – он был священник Бога Всевышнего, –
GEN|14|19|и благословил его, и сказал: благословен Аврам от Бога Всевышнего, Владыки неба и земли;
GEN|14|20|и благословен Бог Всевышний, Который предал врагов твоих в руки твои. [Аврам] дал ему десятую часть из всего.
GEN|14|21|И сказал царь Содомский Авраму: отдай мне людей, а имение возьми себе.
GEN|14|22|Но Аврам сказал царю Содомскому: поднимаю руку мою к Господу Богу Всевышнему, Владыке неба и земли,
GEN|14|23|что даже нитки и ремня от обуви не возьму из всего твоего, чтобы ты не сказал: я обогатил Аврама;
GEN|14|24|кроме того, что съели отроки, и кроме доли, принадлежащей людям, которые ходили со мною; Анер, Эшкол и Мамрий пусть возьмут свою долю.
GEN|15|1|После сих происшествий было слово Господа к Авраму в видении, и сказано: не бойся, Аврам; Я твой щит; награда твоя весьма велика.
GEN|15|2|Аврам сказал: Владыка Господи! что Ты дашь мне? я остаюсь бездетным; распорядитель в доме моем этот Елиезер из Дамаска.
GEN|15|3|И сказал Аврам: вот, Ты не дал мне потомства, и вот, домочадец мой наследник мой.
GEN|15|4|И было слово Господа к нему, и сказано: не будет он твоим наследником, но тот, кто произойдет из чресл твоих, будет твоим наследником.
GEN|15|5|И вывел его вон и сказал: посмотри на небо и сосчитай звезды, если ты можешь счесть их. И сказал ему: столько будет у тебя потомков.
GEN|15|6|Аврам поверил Господу, и Он вменил ему это в праведность.
GEN|15|7|И сказал ему: Я Господь, Который вывел тебя из Ура Халдейского, чтобы дать тебе землю сию во владение.
GEN|15|8|Он сказал: Владыка Господи! по чему мне узнать, что я буду владеть ею?
GEN|15|9|[Господь] сказал ему: возьми Мне трехлетнюю телицу, трехлетнюю козу, трехлетнего овна, горлицу и молодого голубя.
GEN|15|10|Он взял всех их, рассек их пополам и положил одну часть против другой; только птиц не рассек.
GEN|15|11|И налетели на трупы хищные птицы; но Аврам отгонял их.
GEN|15|12|При захождении солнца крепкий сон напал на Аврама, и вот, напал на него ужас и мрак великий.
GEN|15|13|И сказал [Господь] Авраму: знай, что потомки твои будут пришельцами в земле не своей, и поработят их, и будут угнетать их четыреста лет,
GEN|15|14|но Я произведу суд над народом, у которого они будут в порабощении; после сего они выйдут с большим имуществом,
GEN|15|15|а ты отойдешь к отцам твоим в мире [и] будешь погребен в старости доброй;
GEN|15|16|в четвертом роде возвратятся они сюда: ибо [мера] беззаконий Аморреев доселе еще не наполнилась.
GEN|15|17|Когда зашло солнце и наступила тьма, вот, дым [как бы из] печи и пламя огня прошли между рассеченными [животными].
GEN|15|18|В этот день заключил Господь завет с Аврамом, сказав: потомству твоему даю Я землю сию, от реки Египетской до великой реки, реки Евфрата:
GEN|15|19|Кенеев, Кенезеев, Кедмонеев,
GEN|15|20|Хеттеев, Ферезеев, Рефаимов,
GEN|15|21|Аморреев, Хананеев, Гергесеев и Иевусеев.
GEN|16|1|Но Сара, жена Аврамова, не рождала ему. У ней была служанка Египтянка, именем Агарь.
GEN|16|2|И сказала Сара Авраму: вот, Господь заключил чрево мое, чтобы мне не рождать; войди же к служанке моей: может быть, я буду иметь детей от нее. Аврам послушался слов Сары.
GEN|16|3|И взяла Сара, жена Аврамова, служанку свою, Египтянку Агарь, по истечении десяти лет пребывания Аврамова в земле Ханаанской, и дала ее Авраму, мужу своему, в жену.
GEN|16|4|Он вошел к Агари, и она зачала. Увидев же, что зачала, она стала презирать госпожу свою.
GEN|16|5|И сказала Сара Авраму: в обиде моей ты виновен; я отдала служанку мою в недро твое; а она, увидев, что зачала, стала презирать меня; Господь пусть будет судьею между мною и между тобою.
GEN|16|6|Аврам сказал Саре: вот, служанка твоя в твоих руках; делай с нею, что тебе угодно. И Сара стала притеснять ее, и она убежала от нее.
GEN|16|7|И нашел ее Ангел Господень у источника воды в пустыне, у источника на дороге к Суру.
GEN|16|8|И сказал ей: Агарь, служанка Сарина! откуда ты пришла и куда идешь? Она сказала: я бегу от лица Сары, госпожи моей.
GEN|16|9|Ангел Господень сказал ей: возвратись к госпоже своей и покорись ей.
GEN|16|10|И сказал ей Ангел Господень: умножая умножу потомство твое, так что нельзя будет и счесть его от множества.
GEN|16|11|И еще сказал ей Ангел Господень: вот, ты беременна, и родишь сына, и наречешь ему имя Измаил, ибо услышал Господь страдание твое;
GEN|16|12|он будет [между] людьми, [как] дикий осел; руки его на всех, и руки всех на него; жить будет он пред лицем всех братьев своих.
GEN|16|13|И нарекла [Агарь] Господа, Который говорил к ней, [сим] именем: Ты Бог видящий меня. Ибо сказала она: точно я видела здесь в след видящего меня.
GEN|16|14|Посему источник [тот] называется: Беэр–лахай–рои. Он находится между Кадесом и между Баредом.
GEN|16|15|Агарь родила Авраму сына; и нарек [Аврам] имя сыну своему, рожденному от Агари: Измаил.
GEN|16|16|Аврам был восьмидесяти шести лет, когда Агарь родила Авраму Измаила.
GEN|17|1|Аврам был девяноста девяти лет, и Господь явился Авраму и сказал ему: Я Бог Всемогущий; ходи предо Мною и будь непорочен;
GEN|17|2|и поставлю завет Мой между Мною и тобою, и весьма, весьма размножу тебя.
GEN|17|3|И пал Аврам на лице свое. Бог продолжал говорить с ним и сказал:
GEN|17|4|Я – вот завет Мой с тобою: ты будешь отцом множества народов,
GEN|17|5|и не будешь ты больше называться Аврамом, но будет тебе имя: Авраам, ибо Я сделаю тебя отцом множества народов;
GEN|17|6|и весьма, весьма распложу тебя, и произведу от тебя народы, и цари произойдут от тебя;
GEN|17|7|и поставлю завет Мой между Мною и тобою и между потомками твоими после тебя в роды их, завет вечный в том, что Я буду Богом твоим и потомков твоих после тебя;
GEN|17|8|и дам тебе и потомкам твоим после тебя землю, по которой ты странствуешь, всю землю Ханаанскую, во владение вечное; и буду им Богом.
GEN|17|9|И сказал Бог Аврааму: ты же соблюди завет Мой, ты и потомки твои после тебя в роды их.
GEN|17|10|Сей есть завет Мой, который вы [должны] соблюдать между Мною и между вами и между потомками твоими после тебя: да будет у вас обрезан весь мужеский пол;
GEN|17|11|обрезывайте крайнюю плоть вашу: и сие будет знамением завета между Мною и вами.
GEN|17|12|Восьми дней от рождения да будет обрезан у вас в роды ваши всякий [младенец] мужеского пола, рожденный в доме и купленный за серебро у какого–нибудь иноплеменника, который не от твоего семени.
GEN|17|13|Непременно да будет обрезан рожденный в доме твоем и купленный за серебро твое, и будет завет Мой на теле вашем заветом вечным.
GEN|17|14|Необрезанный же мужеского пола, который не обрежет крайней плоти своей, истребится душа та из народа своего, [ибо] он нарушил завет Мой.
GEN|17|15|И сказал Бог Аврааму: Сару, жену твою, не называй Сарою, но да будет имя ей: Сарра;
GEN|17|16|Я благословлю ее и дам тебе от нее сына; благословлю ее, и произойдут от нее народы, и цари народов произойдут от нее.
GEN|17|17|И пал Авраам на лице свое, и рассмеялся, и сказал сам в себе: неужели от столетнего будет сын? и Сарра, девяностолетняя, неужели родит?
GEN|17|18|И сказал Авраам Богу: о, хотя бы Измаил был жив пред лицем Твоим!
GEN|17|19|Бог же сказал: именно Сарра, жена твоя, родит тебе сына, и ты наречешь ему имя: Исаак; и поставлю завет Мой с ним заветом вечным [и] потомству его после него.
GEN|17|20|И о Измаиле Я услышал тебя: вот, Я благословлю его, и возращу его, и весьма, весьма размножу; двенадцать князей родятся от него; и Я произведу от него великий народ.
GEN|17|21|Но завет Мой поставлю с Исааком, которого родит тебе Сарра в сие самое время на другой год.
GEN|17|22|И Бог перестал говорить с Авраамом и восшел от него.
GEN|17|23|И взял Авраам Измаила, сына своего, и всех рожденных в доме своем и всех купленных за серебро свое, весь мужеский пол людей дома Авраамова; и обрезал крайнюю плоть их в тот самый день, как сказал ему Бог.
GEN|17|24|Авраам был девяноста девяти лет, когда была обрезана крайняя плоть его.
GEN|17|25|А Измаил, сын его, был тринадцати лет, когда была обрезана крайняя плоть его.
GEN|17|26|В тот же самый день обрезаны были Авраам и Измаил, сын его,
GEN|17|27|и с ним обрезан был весь мужеский пол дома его, рожденные в доме и купленные за серебро у иноплеменников.
GEN|18|1|И явился ему Господь у дубравы Мамре, когда он сидел при входе в шатер, во время зноя дневного.
GEN|18|2|Он возвел очи свои и взглянул, и вот, три мужа стоят против него. Увидев, он побежал навстречу им от входа в шатер и поклонился до земли,
GEN|18|3|и сказал: Владыка! если я обрел благоволение пред очами Твоими, не пройди мимо раба Твоего;
GEN|18|4|и принесут немного воды, и омоют ноги ваши; и отдохните под сим деревом,
GEN|18|5|а я принесу хлеба, и вы подкрепите сердца ваши; потом пойдите; так как вы идете мимо раба вашего. Они сказали: сделай так, как говоришь.
GEN|18|6|И поспешил Авраам в шатер к Сарре и сказал: поскорее замеси три саты лучшей муки и сделай пресные хлебы.
GEN|18|7|И побежал Авраам к стаду, и взял теленка нежного и хорошего, и дал отроку, и тот поспешил приготовить его.
GEN|18|8|И взял масла и молока и теленка приготовленного, и поставил перед ними, а сам стоял подле них под деревом. И они ели.
GEN|18|9|И сказали ему: где Сарра, жена твоя? Он отвечал: здесь, в шатре.
GEN|18|10|И сказал [один из них]: Я опять буду у тебя в это же время, и будет сын у Сарры, жены твоей. А Сарра слушала у входа в шатер, сзади его.
GEN|18|11|Авраам же и Сарра были стары и в летах преклонных, и обыкновенное у женщин у Сарры прекратилось.
GEN|18|12|Сарра внутренно рассмеялась, сказав: мне ли, когда я состарилась, иметь сие утешение? и господин мой стар.
GEN|18|13|И сказал Господь Аврааму: отчего это рассмеялась Сарра, сказав: "неужели я действительно могу родить, когда я состарилась"?
GEN|18|14|Есть ли что трудное для Господа? В назначенный срок буду Я у тебя в следующем году, и у Сарры [будет] сын.
GEN|18|15|Сарра же не призналась, а сказала: я не смеялась. Ибо она испугалась. Но Он сказал: нет, ты рассмеялась.
GEN|18|16|И встали те мужи и оттуда отправились к Содому; Авраам же пошел с ними, проводить их.
GEN|18|17|И сказал Господь: утаю ли Я от Авраама, что хочу делать!
GEN|18|18|От Авраама точно произойдет народ великий и сильный, и благословятся в нем все народы земли,
GEN|18|19|ибо Я избрал его для того, чтобы он заповедал сынам своим и дому своему после себя, ходить путем Господним, творя правду и суд; и исполнит Господь над Авраамом, что сказал о нем.
GEN|18|20|И сказал Господь: вопль Содомский и Гоморрский, велик он, и грех их, тяжел он весьма;
GEN|18|21|сойду и посмотрю, точно ли они поступают так, каков вопль на них, восходящий ко Мне, или нет; узнаю.
GEN|18|22|И обратились мужи оттуда и пошли в Содом; Авраам же еще стоял пред лицем Господа.
GEN|18|23|И подошел Авраам и сказал: неужели Ты погубишь праведного с нечестивым?
GEN|18|24|может быть, есть в этом городе пятьдесят праведников? неужели Ты погубишь, и не пощадишь места сего ради пятидесяти праведников, в нем?
GEN|18|25|не может быть, чтобы Ты поступил так, чтобы Ты погубил праведного с нечестивым, чтобы то же было с праведником, что с нечестивым; не может быть от Тебя! Судия всей земли поступит ли неправосудно?
GEN|18|26|Господь сказал: если Я найду в городе Содоме пятьдесят праведников, то Я ради них пощажу все место сие.
GEN|18|27|Авраам сказал в ответ: вот, я решился говорить Владыке, я, прах и пепел:
GEN|18|28|может быть, до пятидесяти праведников недостанет пяти, неужели за [недостатком] пяти Ты истребишь весь город? Он сказал: не истреблю, если найду там сорок пять.
GEN|18|29|[Авраам] продолжал говорить с Ним и сказал: может быть, найдется там сорок? Он сказал: не сделаю [того] и ради сорока.
GEN|18|30|И сказал [Авраам]: да не прогневается Владыка, что я буду говорить: может быть, найдется там тридцать? Он сказал: не сделаю, если найдется там тридцать.
GEN|18|31|[Авраам] сказал: вот, я решился говорить Владыке: может быть, найдется там двадцать? Он сказал: не истреблю ради двадцати.
GEN|18|32|[Авраам] сказал: да не прогневается Владыка, что я скажу еще однажды: может быть, найдется там десять? Он сказал: не истреблю ради десяти.
GEN|18|33|И пошел Господь, перестав говорить с Авраамом; Авраам же возвратился в свое место.
GEN|19|1|И пришли те два Ангела в Содом вечером, когда Лот сидел у ворот Содома. Лот увидел, и встал, чтобы встретить их, и поклонился лицем до земли
GEN|19|2|и сказал: государи мои! зайдите в дом раба вашего и ночуйте, и умойте ноги ваши, и встаньте поутру и пойдете в путь свой. Но они сказали: нет, мы ночуем на улице.
GEN|19|3|Он же сильно упрашивал их; и они пошли к нему и пришли в дом его. Он сделал им угощение и испек пресные хлебы, и они ели.
GEN|19|4|Еще не легли они спать, как городские жители, Содомляне, от молодого до старого, весь народ со [всех] концов [города], окружили дом
GEN|19|5|и вызвали Лота и говорили ему: где люди, пришедшие к тебе на ночь? выведи их к нам; мы познаем их.
GEN|19|6|Лот вышел к ним ко входу, и запер за собою дверь,
GEN|19|7|и сказал: братья мои, не делайте зла;
GEN|19|8|вот у меня две дочери, которые не познали мужа; лучше я выведу их к вам, делайте с ними, что вам угодно, только людям сим не делайте ничего, так как они пришли под кров дома моего.
GEN|19|9|Но они сказали: пойди сюда. И сказали: вот пришлец, и хочет судить? теперь мы хуже поступим с тобою, нежели с ними. И очень приступали к человеку сему, к Лоту, и подошли, чтобы выломать дверь.
GEN|19|10|Тогда мужи те простерли руки свои и ввели Лота к себе в дом, и дверь заперли;
GEN|19|11|а людей, бывших при входе в дом, поразили слепотою, от малого до большого, так что они измучились, искав входа.
GEN|19|12|Сказали мужи те Лоту: кто у тебя есть еще здесь? зять ли, сыновья ли твои, дочери ли твои, и кто бы ни был у тебя в городе, всех выведи из сего места,
GEN|19|13|ибо мы истребим сие место, потому что велик вопль на жителей его к Господу, и Господь послал нас истребить его.
GEN|19|14|И вышел Лот, и говорил с зятьями своими, которые брали за себя дочерей его, и сказал: встаньте, выйдите из сего места, ибо Господь истребит сей город. Но зятьям его показалось, что он шутит.
GEN|19|15|Когда взошла заря, Ангелы начали торопить Лота, говоря: встань, возьми жену твою и двух дочерей твоих, которые у тебя, чтобы не погибнуть тебе за беззакония города.
GEN|19|16|И как он медлил, то мужи те, по милости к нему Господней, взяли за руку его и жену его, и двух дочерей его, и вывели его и поставили его вне города.
GEN|19|17|Когда же вывели их вон, [то один из них] сказал: спасай душу свою; не оглядывайся назад и нигде не останавливайся в окрестности сей; спасайся на гору, чтобы тебе не погибнуть.
GEN|19|18|Но Лот сказал им: нет, Владыка!
GEN|19|19|вот, раб Твой обрел благоволение пред очами Твоими, и велика милость Твоя, которую Ты сделал со мною, что спас жизнь мою; но я не могу спасаться на гору, чтоб не застигла меня беда и мне не умереть;
GEN|19|20|вот, ближе бежать в сей город, он же мал; побегу я туда, – он же мал; и сохранится жизнь моя.
GEN|19|21|И сказал ему: вот, в угодность тебе Я сделаю и это: не ниспровергну города, о котором ты говоришь;
GEN|19|22|поспешай, спасайся туда, ибо Я не могу сделать дела, доколе ты не придешь туда. Потому и назван город сей: Сигор.
GEN|19|23|Солнце взошло над землею, и Лот пришел в Сигор.
GEN|19|24|И пролил Господь на Содом и Гоморру дождем серу и огонь от Господа с неба,
GEN|19|25|и ниспроверг города сии, и всю окрестность сию, и всех жителей городов сих, и произрастания земли.
GEN|19|26|Жена же [Лотова] оглянулась позади его, и стала соляным столпом.
GEN|19|27|И встал Авраам рано утром и [пошел] на место, где стоял пред лицем Господа,
GEN|19|28|и посмотрел к Содому и Гоморре и на все пространство окрестности и увидел: вот, дым поднимается с земли, как дым из печи.
GEN|19|29|И было, когда Бог истреблял города окрестности сей, вспомнил Бог об Аврааме и выслал Лота из среды истребления, когда ниспровергал города, в которых жил Лот.
GEN|19|30|И вышел Лот из Сигора и стал жить в горе, и с ним две дочери его, ибо он боялся жить в Сигоре. И жил в пещере, и с ним две дочери его.
GEN|19|31|И сказала старшая младшей: отец наш стар, и нет человека на земле, который вошел бы к нам по обычаю всей земли;
GEN|19|32|итак напоим отца нашего вином, и переспим с ним, и восставим от отца нашего племя.
GEN|19|33|И напоили отца своего вином в ту ночь; и вошла старшая и спала с отцом своим: а он не знал, когда она легла и когда встала.
GEN|19|34|На другой день старшая сказала младшей: вот, я спала вчера с отцом моим; напоим его вином и в эту ночь; и ты войди, спи с ним, и восставим от отца нашего племя.
GEN|19|35|И напоили отца своего вином и в эту ночь; и вошла младшая и спала с ним; и он не знал, когда она легла и когда встала.
GEN|19|36|И сделались обе дочери Лотовы беременными от отца своего,
GEN|19|37|и родила старшая сына, и нарекла ему имя: Моав. Он отец Моавитян доныне.
GEN|19|38|И младшая также родила сына, и нарекла ему имя: Бен–Амми. Он отец Аммонитян доныне.
GEN|20|1|Авраам поднялся оттуда к югу и поселился между Кадесом и между Суром; и был на время в Гераре.
GEN|20|2|И сказал Авраам о Сарре, жене своей: она сестра моя. И послал Авимелех, царь Герарский, и взял Сарру.
GEN|20|3|И пришел Бог к Авимелеху ночью во сне и сказал ему: вот, ты умрешь за женщину, которую ты взял, ибо она имеет мужа.
GEN|20|4|Авимелех же не прикасался к ней и сказал: Владыка! неужели ты погубишь и невинный народ?
GEN|20|5|Не сам ли он сказал мне: она сестра моя? И она сама сказала: он брат мой. Я сделал это в простоте сердца моего и в чистоте рук моих.
GEN|20|6|И сказал ему Бог во сне: и Я знаю, что ты сделал сие в простоте сердца твоего, и удержал тебя от греха предо Мною, потому и не допустил тебя прикоснуться к ней;
GEN|20|7|теперь же возврати жену мужу, ибо он пророк и помолится о тебе, и ты будешь жив; а если не возвратишь, то знай, что непременно умрешь ты и все твои.
GEN|20|8|И встал Авимелех утром рано, и призвал всех рабов своих, и пересказал все слова сии в уши их; и люди сии весьма испугались.
GEN|20|9|И призвал Авимелех Авраама и сказал ему: что ты с нами сделал? чем согрешил я против тебя, что ты навел было на меня и на царство мое великий грех? Ты сделал со мною дела, каких не делают.
GEN|20|10|И сказал Авимелех Аврааму: что ты имел в виду, когда делал это дело?
GEN|20|11|Авраам сказал: я подумал, что нет на месте сем страха Божия, и убьют меня за жену мою;
GEN|20|12|да она и подлинно сестра мне: она дочь отца моего, только не дочь матери моей; и сделалась моею женою;
GEN|20|13|когда Бог повел меня странствовать из дома отца моего, то я сказал ей: сделай со мною сию милость, в какое ни придем мы место, везде говори обо мне: это брат мой.
GEN|20|14|И взял Авимелех мелкого и крупного скота, и рабов и рабынь, и дал Аврааму; и возвратил ему Сарру, жену его.
GEN|20|15|И сказал Авимелех: вот, земля моя пред тобою; живи, где тебе угодно.
GEN|20|16|И Сарре сказал: вот, я дал брату твоему тысячу [сиклей] серебра; вот, это тебе покрывало для очей пред всеми, которые с тобою, и пред всеми ты оправдана.
GEN|20|17|И помолился Авраам Богу, и исцелил Бог Авимелеха, и жену его, и рабынь его, и они стали рождать;
GEN|20|18|ибо заключил Господь всякое чрево в доме Авимелеха за Сарру, жену Авраамову.
GEN|21|1|И призрел Господь на Сарру, как сказал; и сделал Господь Сарре, как говорил.
GEN|21|2|Сарра зачала и родила Аврааму сына в старости его во время, о котором говорил ему Бог;
GEN|21|3|и нарек Авраам имя сыну своему, родившемуся у него, которого родила ему Сарра, Исаак;
GEN|21|4|и обрезал Авраам Исаака, сына своего, в восьмой день, как заповедал ему Бог.
GEN|21|5|Авраам был ста лет, когда родился у него Исаак, сын его.
GEN|21|6|И сказала Сарра: смех сделал мне Бог; кто ни услышит обо мне, рассмеется.
GEN|21|7|И сказала: кто сказал бы Аврааму: Сарра будет кормить детей грудью? ибо в старости его я родила сына.
GEN|21|8|Дитя выросло и отнято от груди; и Авраам сделал большой пир в тот день, когда Исаак отнят был от груди.
GEN|21|9|И увидела Сарра, что сын Агари Египтянки, которого она родила Аврааму, насмехается,
GEN|21|10|и сказала Аврааму: выгони эту рабыню и сына ее, ибо не наследует сын рабыни сей с сыном моим Исааком.
GEN|21|11|И показалось это Аврааму весьма неприятным ради сына его.
GEN|21|12|Но Бог сказал Аврааму: не огорчайся ради отрока и рабыни твоей; во всем, что скажет тебе Сарра, слушайся голоса ее, ибо в Исааке наречется тебе семя;
GEN|21|13|и от сына рабыни Я произведу народ, потому что он семя твое.
GEN|21|14|Авраам встал рано утром, и взял хлеба и мех воды, и дал Агари, положив ей на плечи, и отрока, и отпустил ее. Она пошла, и заблудилась в пустыне Вирсавии;
GEN|21|15|и не стало воды в мехе, и она оставила отрока под одним кустом
GEN|21|16|и пошла, села вдали, в расстоянии на [один] выстрел из лука. Ибо она сказала: не [хочу] видеть смерти отрока. И она села против, и подняла вопль, и плакала;
GEN|21|17|и услышал Бог голос отрока; и Ангел Божий с неба воззвал к Агари и сказал ей: что с тобою, Агарь? не бойся; Бог услышал голос отрока оттуда, где он находится;
GEN|21|18|встань, подними отрока и возьми его за руку, ибо Я произведу от него великий народ.
GEN|21|19|И Бог открыл глаза ее, и она увидела колодезь с водою, и пошла, наполнила мех водою и напоила отрока.
GEN|21|20|И Бог был с отроком; и он вырос, и стал жить в пустыне, и сделался стрелком из лука.
GEN|21|21|Он жил в пустыне Фаран; и мать его взяла ему жену из земли Египетской.
GEN|21|22|И было в то время, Авимелех с Фихолом, военачальником своим, сказал Аврааму: с тобою Бог во всем, что ты ни делаешь;
GEN|21|23|и теперь поклянись мне здесь Богом, что ты не обидишь ни меня, ни сына моего, ни внука моего; и как я хорошо поступал с тобою, так и ты будешь поступать со мною и землею, в которой ты гостишь.
GEN|21|24|И сказал Авраам: я клянусь.
GEN|21|25|И Авраам упрекал Авимелеха за колодезь с водою, который отняли рабы Авимелеховы.
GEN|21|26|Авимелех же сказал: не знаю, кто это сделал, и ты не сказал мне; я даже и не слыхал [о том] доныне.
GEN|21|27|И взял Авраам мелкого и крупного скота и дал Авимелеху, и они оба заключили союз.
GEN|21|28|И поставил Авраам семь агниц из [стада] мелкого скота особо.
GEN|21|29|Авимелех же сказал Аврааму: на что здесь сии семь агниц, которых ты поставил особо?
GEN|21|30|[он] сказал: семь агниц сих возьми от руки моей, чтобы они были мне свидетельством, что я выкопал этот колодезь.
GEN|21|31|Потому и назвал он сие место: Вирсавия, ибо тут оба они клялись
GEN|21|32|и заключили союз в Вирсавии. И встал Авимелех, и Фихол, военачальник его, и возвратились в землю Филистимскую.
GEN|21|33|И насадил [Авраам] при Вирсавии рощу и призвал там имя Господа, Бога вечного.
GEN|21|34|И жил Авраам в земле Филистимской, как странник, дни многие.
GEN|22|1|И было, после сих происшествий Бог искушал Авраама и сказал ему: Авраам! Он сказал: вот я.
GEN|22|2|[Бог] сказал: возьми сына твоего, единственного твоего, которого ты любишь, Исаака; и пойди в землю Мориа и там принеси его во всесожжение на одной из гор, о которой Я скажу тебе.
GEN|22|3|Авраам встал рано утром, оседлал осла своего, взял с собою двоих из отроков своих и Исаака, сына своего; наколол дров для всесожжения, и встав пошел на место, о котором сказал ему Бог.
GEN|22|4|На третий день Авраам возвел очи свои, и увидел то место издалека.
GEN|22|5|И сказал Авраам отрокам своим: останьтесь вы здесь с ослом, а я и сын пойдем туда и поклонимся, и возвратимся к вам.
GEN|22|6|И взял Авраам дрова для всесожжения, и возложил на Исаака, сына своего; взял в руки огонь и нож, и пошли оба вместе.
GEN|22|7|И начал Исаак говорить Аврааму, отцу своему, и сказал: отец мой! Он отвечал: вот я, сын мой. Он сказал: вот огонь и дрова, где же агнец для всесожжения?
GEN|22|8|Авраам сказал: Бог усмотрит Себе агнца для всесожжения, сын мой. И шли [далее] оба вместе.
GEN|22|9|И пришли на место, о котором сказал ему Бог; и устроил там Авраам жертвенник, разложил дрова и, связав сына своего Исаака, положил его на жертвенник поверх дров.
GEN|22|10|И простер Авраам руку свою и взял нож, чтобы заколоть сына своего.
GEN|22|11|Но Ангел Господень воззвал к нему с неба и сказал: Авраам! Авраам! Он сказал: вот я.
GEN|22|12|[Ангел] сказал: не поднимай руки твоей на отрока и не делай над ним ничего, ибо теперь Я знаю, что боишься ты Бога и не пожалел сына твоего, единственного твоего, для Меня.
GEN|22|13|И возвел Авраам очи свои и увидел: и вот, позади овен, запутавшийся в чаще рогами своими. Авраам пошел, взял овна и принес его во всесожжение вместо сына своего.
GEN|22|14|И нарек Авраам имя месту тому: Иегова–ире. Посему [и] ныне говорится: на горе Иеговы усмотрится.
GEN|22|15|И вторично воззвал к Аврааму Ангел Господень с неба
GEN|22|16|и сказал: Мною клянусь, говорит Господь, что, так как ты сделал сие дело, и не пожалел сына твоего, единственного твоего,
GEN|22|17|то Я благословляя благословлю тебя и умножая умножу семя твое, как звезды небесные и как песок на берегу моря; и овладеет семя твое городами врагов своих;
GEN|22|18|и благословятся в семени твоем все народы земли за то, что ты послушался гласа Моего.
GEN|22|19|И возвратился Авраам к отрокам своим, и встали и пошли вместе в Вирсавию; и жил Авраам в Вирсавии.
GEN|22|20|После сих происшествий Аврааму возвестили, сказав: вот, и Милка родила Нахору, брату твоему, сынов:
GEN|22|21|Уца, первенца его, Вуза, брата сему, Кемуила, отца Арамова,
GEN|22|22|Кеседа, Хазо, Пилдаша, Идлафа и Вафуила;
GEN|22|23|от Вафуила родилась Ревекка. Восьмерых сих родила Милка Нахору, брату Авраамову;
GEN|22|24|и наложница его, именем Реума, также родила Теваха, Гахама, Тахаша и Мааху.
GEN|23|1|Жизни Сарриной было сто двадцать семь лет: [вот] лета жизни Сарриной;
GEN|23|2|и умерла Сарра в Кириаф–Арбе, что [ныне] Хеврон, в земле Ханаанской. И пришел Авраам рыдать по Сарре и оплакивать ее.
GEN|23|3|И отошел Авраам от умершей своей, и говорил сынам Хетовым, и сказал:
GEN|23|4|я у вас пришлец и поселенец; дайте мне в собственность [место] [для] гроба между вами, чтобы мне умершую мою схоронить от глаз моих.
GEN|23|5|Сыны Хета отвечали Аврааму и сказали ему:
GEN|23|6|послушай нас, господин наш; ты князь Божий посреди нас; в лучшем из наших погребальных мест похорони умершую твою; никто из нас не откажет тебе в погребальном месте, для погребения умершей твоей.
GEN|23|7|Авраам встал и поклонился народу земли той, сынам Хетовым;
GEN|23|8|и говорил им и сказал: если вы согласны, чтобы я похоронил умершую мою, то послушайте меня, попросите за меня Ефрона, сына Цохарова,
GEN|23|9|чтобы он отдал мне пещеру Махпелу, которая у него на конце поля его, чтобы за довольную цену отдал ее мне посреди вас, в собственность для погребения.
GEN|23|10|Ефрон же сидел посреди сынов Хетовых; и отвечал Ефрон Хеттеянин Аврааму вслух сынов Хета, всех входящих во врата города его, и сказал:
GEN|23|11|нет, господин мой, послушай меня: я даю тебе поле и пещеру, которая на нем, даю тебе, пред очами сынов народа моего дарю тебе ее, похорони умершую твою.
GEN|23|12|Авраам поклонился пред народом земли той
GEN|23|13|и говорил Ефрону вслух народа земли той и сказал: если послушаешь, я даю тебе за поле серебро; возьми у меня, и я похороню там умершую мою.
GEN|23|14|Ефрон отвечал Аврааму и сказал ему:
GEN|23|15|господин мой! послушай меня: земля [стоит] четыреста сиклей серебра; для меня и для тебя что это? похорони умершую твою.
GEN|23|16|Авраам выслушал Ефрона; и отвесил Авраам Ефрону серебра, сколько он объявил вслух сынов Хетовых, четыреста сиклей серебра, какое ходит у купцов.
GEN|23|17|И стало поле Ефроново, которое при Махпеле, против Мамре, поле и пещера, которая на нем, и все деревья, которые на поле, во всех пределах его вокруг,
GEN|23|18|владением Авраамовым пред очами сынов Хета, всех входящих во врата города его.
GEN|23|19|После сего Авраам похоронил Сарру, жену свою, в пещере поля в Махпеле, против Мамре, что [ныне] Хеврон, в земле Ханаанской.
GEN|23|20|Так достались Аврааму от сынов Хетовых поле и пещера, которая на нем, в собственность для погребения.
GEN|24|1|Авраам был уже стар и в летах преклонных. Господь благословил Авраама всем.
GEN|24|2|И сказал Авраам рабу своему, старшему в доме его, управлявшему всем, что у него было: положи руку твою под стегно мое
GEN|24|3|и клянись мне Господом, Богом неба и Богом земли, что ты не возьмешь сыну моему жены из дочерей Хананеев, среди которых я живу,
GEN|24|4|но пойдешь в землю мою, на родину мою, и возьмешь жену сыну моему Исааку.
GEN|24|5|Раб сказал ему: может быть, не захочет женщина идти со мною в эту землю, должен ли я возвратить сына твоего в землю, из которой ты вышел?
GEN|24|6|Авраам сказал ему: берегись, не возвращай сына моего туда;
GEN|24|7|Господь, Бог неба, Который взял меня из дома отца моего и из земли рождения моего, Который говорил мне и Который клялся мне, говоря: "потомству твоему дам сию землю", – Он пошлет Ангела Своего пред тобою, и ты возьмешь жену сыну моему оттуда;
GEN|24|8|если же не захочет женщина идти с тобою, ты будешь свободен от сей клятвы моей; только сына моего не возвращай туда.
GEN|24|9|И положил раб руку свою под стегно Авраама, господина своего, и клялся ему в сем.
GEN|24|10|И взял раб из верблюдов господина своего десять верблюдов и пошел. В руках у него были также всякие сокровища господина его. Он встал и пошел в Месопотамию, в город Нахора,
GEN|24|11|и остановил верблюдов вне города, у колодезя воды, под вечер, в то время, когда выходят женщины черпать,
GEN|24|12|и сказал: Господи, Боже господина моего Авраама! пошли [ее] сегодня навстречу мне и сотвори милость с господином моим Авраамом;
GEN|24|13|вот, я стою у источника воды, и дочери жителей города выходят черпать воду;
GEN|24|14|и девица, которой я скажу: "наклони кувшин твой, я напьюсь", и которая скажет: "пей, я и верблюдам твоим дам пить", – вот та, которую Ты назначил рабу Твоему Исааку; и по сему узнаю я, что Ты творишь милость с господином моим.
GEN|24|15|Еще не перестал он говорить, и вот, вышла Ревекка, которая родилась от Вафуила, сына Милки, жены Нахора, брата Авраамова, и кувшин ее на плече ее;
GEN|24|16|девица [была] прекрасна видом, дева, которой не познал муж. Она сошла к источнику, наполнила кувшин свой и пошла вверх.
GEN|24|17|И побежал раб навстречу ей и сказал: дай мне испить немного воды из кувшина твоего.
GEN|24|18|Она сказала: пей, господин мой. И тотчас спустила кувшин свой на руку свою и напоила его.
GEN|24|19|И, когда напоила его, сказала: я стану черпать и для верблюдов твоих, пока не напьются.
GEN|24|20|И тотчас вылила воду из кувшина своего в поило и побежала опять к колодезю почерпнуть, и начерпала для всех верблюдов его.
GEN|24|21|Человек тот смотрел на нее с изумлением в молчании, желая уразуметь, благословил ли Господь путь его, или нет.
GEN|24|22|Когда верблюды перестали пить, тогда человек тот взял золотую серьгу, весом полсикля, и два запястья на руки ей, весом в десять [сиклей] золота;
GEN|24|23|И сказал: чья ты дочь? скажи мне, есть ли в доме отца твоего место нам ночевать?
GEN|24|24|Она сказала ему: я дочь Вафуила, сына Милки, которого она родила Нахору.
GEN|24|25|И еще сказала ему: у нас много соломы и корму, и [есть] место для ночлега.
GEN|24|26|И преклонился человек тот и поклонился Господу,
GEN|24|27|и сказал: благословен Господь Бог господина моего Авраама, Который не оставил господина моего милостью Своею и истиною Своею! Господь прямым путем привел меня к дому брата господина моего.
GEN|24|28|Девица побежала и рассказала об этом в доме матери своей.
GEN|24|29|У Ревекки был брат, именем Лаван. Лаван выбежал к тому человеку, к источнику.
GEN|24|30|И когда он увидел серьгу и запястья на руках у сестры своей и услышал слова Ревекки, сестры своей, которая говорила: так говорил со мною этот человек, – то пришел к человеку, и вот, он стоит при верблюдах у источника;
GEN|24|31|и сказал: войди, благословенный Господом; зачем ты стоишь вне? я приготовил дом и место для верблюдов.
GEN|24|32|И вошел человек. [Лаван] расседлал верблюдов и дал соломы и корму верблюдам, и воды умыть ноги ему и людям, которые были с ним;
GEN|24|33|и предложена была ему пища; но он сказал: не стану есть, доколе не скажу дела своего. И сказали: говори.
GEN|24|34|Он сказал: я раб Авраамов;
GEN|24|35|Господь весьма благословил господина моего, и он сделался великим: Он дал ему овец и волов, серебро и золото, рабов и рабынь, верблюдов и ослов;
GEN|24|36|Сарра, жена господина моего, уже состарившись, родила господину моему сына, которому он отдал все, что у него;
GEN|24|37|и взял с меня клятву господин мой, сказав: не бери жены сыну моему из дочерей Хананеев, в земле которых я живу,
GEN|24|38|а пойди в дом отца моего и к родственникам моим, и возьмешь жену сыну моему.
GEN|24|39|Я сказал господину моему: может быть, не пойдет женщина со мною.
GEN|24|40|Он сказал мне: Господь, пред лицем Которого я хожу, пошлет с тобою Ангела Своего и благоустроит путь твой, и возьмешь жену сыну моему из родных моих и из дома отца моего;
GEN|24|41|тогда будешь ты свободен от клятвы моей, когда сходишь к родственникам моим; и если они не дадут тебе, то будешь свободен от клятвы моей.
GEN|24|42|И пришел я ныне к источнику, и сказал: Господи, Боже господина моего Авраама! Если Ты благоустроишь путь, который я совершаю,
GEN|24|43|то вот, я стою у источника воды, и девица, которая выйдет почерпать, и которой я скажу: дай мне испить немного из кувшина твоего,
GEN|24|44|и которая скажет мне: "и ты пей, и верблюдам твоим я начерпаю" – вот жена, которую Господь назначил сыну господина моего.
GEN|24|45|Еще не перестал я говорить в уме моем, и вот вышла Ревекка, и кувшин ее на плече ее, и сошла к источнику и почерпнула; и я сказал ей: напой меня.
GEN|24|46|Она тотчас спустила с себя кувшин свой и сказала: пей, и верблюдов твоих я напою. И я пил, и верблюдов она напоила.
GEN|24|47|Я спросил ее и сказал: чья ты дочь? Она сказала: дочь Вафуила, сына Нахорова, которого родила ему Милка. И дал я серьги ей и запястья на руки ее.
GEN|24|48|И преклонился я и поклонился Господу, и благословил Господа, Бога господина моего Авраама, Который прямым путем привел меня, чтобы взять дочь брата господина моего за сына его.
GEN|24|49|И ныне скажите мне: намерены ли вы оказать милость и правду господину моему или нет? скажите мне, и я обращусь направо, или налево.
GEN|24|50|И отвечали Лаван и Вафуил и сказали: от Господа пришло это дело; мы не можем сказать тебе вопреки ни худого, ни доброго;
GEN|24|51|вот Ревекка пред тобою; возьми и пойди; пусть будет она женою сыну господина твоего, как сказал Господь.
GEN|24|52|Когда раб Авраамов услышал слова их, то поклонился Господу до земли.
GEN|24|53|И вынул раб серебряные вещи и золотые вещи и одежды и дал Ревекке; также и брату ее и матери ее дал богатые подарки.
GEN|24|54|И ели и пили он и люди, бывшие с ним, и переночевали. Когда же встали поутру, то он сказал: отпустите меня к господину моему.
GEN|24|55|Но брат ее и мать ее сказали: пусть побудет с нами девица дней хотя десять, потом пойдешь.
GEN|24|56|Он сказал им: не удерживайте меня, ибо Господь благоустроил путь мой; отпустите меня, и я пойду к господину моему.
GEN|24|57|Они сказали: призовем девицу и спросим, что она скажет.
GEN|24|58|И призвали Ревекку и сказали ей: пойдешь ли с этим человеком? Она сказала: пойду.
GEN|24|59|И отпустили Ревекку, сестру свою, и кормилицу ее, и раба Авраамова, и людей его.
GEN|24|60|И благословили Ревекку и сказали ей: сестра наша! да родятся от тебя тысячи тысяч, и да владеет потомство твое жилищами врагов твоих!
GEN|24|61|И встала Ревекка и служанки ее, и сели на верблюдов, и поехали за тем человеком. И раб взял Ревекку и пошел.
GEN|24|62|А Исаак пришел из Беэр–лахай–рои, ибо жил он в земле полуденной.
GEN|24|63|При наступлении вечера Исаак вышел в поле поразмыслить, и возвел очи свои, и увидел: вот, идут верблюды.
GEN|24|64|Ревекка взглянула, и увидела Исаака, и спустилась с верблюда.
GEN|24|65|И сказала рабу: кто этот человек, который идет по полю навстречу нам? Раб сказал: это господин мой. И она взяла покрывало и покрылась.
GEN|24|66|Раб же сказал Исааку все, что сделал.
GEN|24|67|И ввел ее Исаак в шатер Сарры, матери своей, и взял Ревекку, и она сделалась ему женою, и он возлюбил ее; и утешился Исаак в [печали] по матери своей.
GEN|25|1|И взял Авраам еще жену, именем Хеттуру.
GEN|25|2|Она родила ему Зимрана, Иокшана, Медана, Мадиана, Ишбака и Шуаха.
GEN|25|3|Иокшан родил Шеву и Дедана. Сыны Дедана были: Ашурим, Летушим и Леюмим.
GEN|25|4|Сыны Мадиана: Ефа, Ефер, Ханох, Авида и Елдага. Все сии сыны Хеттуры.
GEN|25|5|И отдал Авраам все, что было у него, Исааку,
GEN|25|6|а сынам наложниц, которые были у Авраама, дал Авраам подарки и отослал их от Исаака, сына своего, еще при жизни своей, на восток, в землю восточную.
GEN|25|7|Дней жизни Авраамовой, которые он прожил, было сто семьдесят пять лет;
GEN|25|8|и скончался Авраам, и умер в старости доброй, престарелый и насыщенный [жизнью], и приложился к народу своему.
GEN|25|9|И погребли его Исаак и Измаил, сыновья его, в пещере Махпеле, на поле Ефрона, сына Цохара, Хеттеянина, которое против Мамре,
GEN|25|10|на поле, которые Авраам приобрел от сынов Хетовых. Там погребены Авраам и Сарра, жена его.
GEN|25|11|По смерти Авраама Бог благословил Исаака, сына его. Исаак жил при Беэр–лахай–рои.
GEN|25|12|Вот родословие Измаила, сына Авраамова, которого родила Аврааму Агарь Египтянка, служанка Саррина;
GEN|25|13|и вот имена сынов Измаиловых, имена их по родословию их: первенец Измаилов Наваиоф, [за ним] Кедар, Адбеел, Мивсам,
GEN|25|14|Мишма, Дума, Масса,
GEN|25|15|Хадад, Фема, Иетур, Нафиш и Кедма.
GEN|25|16|Сии суть сыны Измаиловы, и сии имена их, в селениях их, в кочевьях их. [Это] двенадцать князей племен их.
GEN|25|17|Лет же жизни Измаиловой было сто тридцать семь лет; и скончался он, и умер, и приложился к народу своему.
GEN|25|18|Они жили от Хавилы до Сура, что пред Египтом, как идешь к Ассирии. Они поселились пред лицем всех братьев своих.
GEN|25|19|Вот родословие Исаака, сына Авраамова. Авраам родил Исаака.
GEN|25|20|Исаак был сорока лет, когда он взял себе в жену Ревекку, дочь Вафуила Арамеянина из Месопотамии, сестру Лавана Арамеянина.
GEN|25|21|И молился Исаак Господу о жене своей, потому что она была неплодна; и Господь услышал его, и зачала Ревекка, жена его.
GEN|25|22|Сыновья в утробе ее стали биться, и она сказала: если так будет, то для чего мне это? И пошла вопросить Господа.
GEN|25|23|Господь сказал ей: два племени во чреве твоем, и два различных народа произойдут из утробы твоей; один народ сделается сильнее другого, и больший будет служить меньшему.
GEN|25|24|И настало время родить ей: и вот близнецы в утробе ее.
GEN|25|25|Первый вышел красный, весь, как кожа, косматый; и нарекли ему имя Исав.
GEN|25|26|Потом вышел брат его, держась рукою своею за пяту Исава; и наречено ему имя Иаков. Исаак же был шестидесяти лет, когда они родились.
GEN|25|27|Дети выросли, и стал Исав человеком искусным в звероловстве, человеком полей; а Иаков человеком кротким, живущим в шатрах.
GEN|25|28|Исаак любил Исава, потому что дичь его была по вкусу его, а Ревекка любила Иакова.
GEN|25|29|И сварил Иаков кушанье; а Исав пришел с поля усталый.
GEN|25|30|И сказал Исав Иакову: дай мне поесть красного, красного этого, ибо я устал. От сего дано ему прозвание: Едом.
GEN|25|31|Но Иаков сказал: продай мне теперь же свое первородство.
GEN|25|32|Исав сказал: вот, я умираю, что мне в этом первородстве?
GEN|25|33|Иаков сказал: поклянись мне теперь же. Он поклялся ему, и продал первородство свое Иакову.
GEN|25|34|И дал Иаков Исаву хлеба и кушанья из чечевицы; и он ел и пил, и встал и пошел; и пренебрег Исав первородство.
GEN|26|1|Был голод в земле, сверх прежнего голода, который был во дни Авраама; и пошел Исаак к Авимелеху, царю Филистимскому, в Герар.
GEN|26|2|Господь явился ему и сказал: не ходи в Египет; живи в земле, о которой Я скажу тебе,
GEN|26|3|странствуй по сей земле, и Я буду с тобою и благословлю тебя, ибо тебе и потомству твоему дам все земли сии и исполню клятву, которою Я клялся Аврааму, отцу твоему;
GEN|26|4|умножу потомство твое, как звезды небесные, и дам потомству твоему все земли сии; благословятся в семени твоем все народы земные,
GEN|26|5|за то, что Авраам послушался гласа Моего и соблюдал, что Мною [заповедано] было соблюдать: повеления Мои, уставы Мои и законы Мои.
GEN|26|6|Исаак поселился в Гераре.
GEN|26|7|Жители места того спросили о жене его, и он сказал: это сестра моя; потому что боялся сказать: жена моя, чтобы не убили меня, [думал он], жители места сего за Ревекку, потому что она прекрасна видом.
GEN|26|8|Но когда уже много времени он там прожил, Авимелех, царь Филистимский, посмотрев в окно, увидел, что Исаак играет с Ревеккою, женою своею.
GEN|26|9|И призвал Авимелех Исаака и сказал: вот, это жена твоя; как же ты сказал: она сестра моя? Исаак сказал ему: потому что я думал, не умереть бы мне ради ее.
GEN|26|10|Но Авимелех сказал: что это ты сделал с нами? едва один из народа не совокупился с женою твоею, и ты ввел бы нас в грех.
GEN|26|11|И дал Авимелех повеление всему народу, сказав: кто прикоснется к сему человеку и к жене его, тот предан будет смерти.
GEN|26|12|И сеял Исаак в земле той и получил в тот год ячменя во сто крат: так благословил его Господь.
GEN|26|13|И стал великим человек сей и возвеличивался больше и больше до того, что стал весьма великим.
GEN|26|14|У него были стада мелкого и стада крупного скота и множество пахотных полей, и Филистимляне стали завидовать ему.
GEN|26|15|И все колодези, которые выкопали рабы отца его при жизни отца его Авраама, Филистимляне завалили и засыпали землею.
GEN|26|16|И Авимелех сказал Исааку: удались от нас, ибо ты сделался гораздо сильнее нас.
GEN|26|17|И Исаак удалился оттуда, и расположился шатрами в долине Герарской, и поселился там.
GEN|26|18|И вновь выкопал Исаак колодези воды, которые выкопаны были во дни Авраама, отца его, и которые завалили Филистимляне по смерти Авраама; и назвал их теми же именами, которыми назвал их отец его.
GEN|26|19|И копали рабы Исааковы в долине и нашли там колодезь воды живой.
GEN|26|20|И спорили пастухи Герарские с пастухами Исаака, говоря: наша вода. И он нарек колодезю имя: Есек, потому что спорили с ним.
GEN|26|21|выкопали другой колодезь; спорили также и о нем; и он нарек ему имя: Ситна.
GEN|26|22|И он двинулся отсюда и выкопал иной колодезь, о котором уже не спорили, и нарек ему имя: Реховоф, ибо, сказал он, теперь Господь дал нам пространное место, и мы размножимся на земле.
GEN|26|23|Оттуда перешел он в Вирсавию.
GEN|26|24|И в ту ночь явился ему Господь и сказал: Я Бог Авраама, отца твоего; не бойся, ибо Я с тобою; и благословлю тебя и умножу потомство твое, ради Авраама, раба Моего.
GEN|26|25|И он устроил там жертвенник и призвал имя Господа. И раскинул там шатер свой, и выкопали там рабы Исааковы колодезь.
GEN|26|26|Пришел к нему из Герара Авимелех и Ахузаф, друг его, и Фихол, военачальник его.
GEN|26|27|Исаак сказал им: для чего вы пришли ко мне, когда вы возненавидели меня и выслали меня от себя?
GEN|26|28|Они сказали: мы ясно увидели, что Господь с тобою, и потому мы сказали: поставим между нами и тобою клятву и заключим с тобою союз,
GEN|26|29|чтобы ты не делал нам зла, как и мы не коснулись до тебя, а делали тебе одно доброе и отпустили тебя с миром; теперь ты благословен Господом.
GEN|26|30|Он сделал им пиршество, и они ели и пили.
GEN|26|31|И встав рано утром, поклялись друг другу; и отпустил их Исаак, и они пошли от него с миром.
GEN|26|32|В тот же день пришли рабы Исааковы и известили его о колодезе, который копали они, и сказали ему: мы нашли воду.
GEN|26|33|И он назвал его: Шива. Посему имя городу тому Беэршива до сего дня.
GEN|26|34|И был Исав сорока лет, и взял себе в жены Иегудифу, дочь Беэра Хеттеянина, и Васемафу, дочь Елона Хеттеянина;
GEN|26|35|и они были в тягость Исааку и Ревекке.
GEN|27|1|Когда Исаак состарился и притупилось зрение глаз его, он призвал старшего сына своего Исава и сказал ему: сын мой! Тот сказал ему: вот я.
GEN|27|2|Он сказал: вот, я состарился; не знаю дня смерти моей;
GEN|27|3|возьми теперь орудия твои, колчан твой и лук твой, пойди в поле, и налови мне дичи,
GEN|27|4|и приготовь мне кушанье, какое я люблю, и принеси мне есть, чтобы благословила тебя душа моя, прежде нежели я умру.
GEN|27|5|Ревекка слышала, когда Исаак говорил сыну своему Исаву. И пошел Исав в поле достать и принести дичи;
GEN|27|6|а Ревекка сказала сыну своему Иакову: вот, я слышала, как отец твой говорил брату твоему Исаву:
GEN|27|7|принеси мне дичи и приготовь мне кушанье; я поем и благословлю тебя пред лицем Господним, пред смертью моею.
GEN|27|8|Теперь, сын мой, послушайся слов моих в том, что я прикажу тебе:
GEN|27|9|пойди в [стадо] и возьми мне оттуда два козленка хороших, и я приготовлю из них отцу твоему кушанье, какое он любит,
GEN|27|10|а ты принесешь отцу твоему, и он поест, чтобы благословить тебя пред смертью своею.
GEN|27|11|Иаков сказал Ревекке, матери своей: Исав, брат мой, человек косматый, а я человек гладкий;
GEN|27|12|может статься, ощупает меня отец мой, и я буду в глазах его обманщиком и наведу на себя проклятие, а не благословение.
GEN|27|13|Мать его сказала ему: на мне пусть будет проклятие твое, сын мой, только послушайся слов моих и пойди, принеси мне.
GEN|27|14|Он пошел, и взял, и принес матери своей; и мать его сделала кушанье, какое любил отец его.
GEN|27|15|И взяла Ревекка богатую одежду старшего сына своего Исава, бывшую у ней в доме, и одела [в нее] младшего сына своего Иакова;
GEN|27|16|а руки его и гладкую шею его обложила кожею козлят;
GEN|27|17|и дала кушанье и хлеб, которые она приготовила, в руки Иакову, сыну своему.
GEN|27|18|Он вошел к отцу своему и сказал: отец мой! Тот сказал: вот я; кто ты, сын мой?
GEN|27|19|Иаков сказал отцу своему: я Исав, первенец твой; я сделал, как ты сказал мне; встань, сядь и поешь дичи моей, чтобы благословила меня душа твоя.
GEN|27|20|И сказал Исаак сыну своему: что так скоро нашел ты, сын мой? Он сказал: потому что Господь Бог твой послал мне навстречу.
GEN|27|21|И сказал Исаак Иакову: подойди, я ощупаю тебя, сын мой, ты ли сын мой Исав, или нет?
GEN|27|22|Иаков подошел к Исааку, отцу своему, и он ощупал его и сказал: голос, голос Иакова; а руки, руки Исавовы.
GEN|27|23|И не узнал его, потому что руки его были, как руки Исава, брата его, косматые; и благословил его
GEN|27|24|и сказал: ты ли сын мой Исав? Он отвечал: я.
GEN|27|25|[Исаак] сказал: подай мне, я поем дичи сына моего, чтобы благословила тебя душа моя. [Иаков] подал ему, и он ел; принес ему и вина, и он пил.
GEN|27|26|Исаак, отец его, сказал ему: подойди, поцелуй меня, сын мой.
GEN|27|27|Он подошел и поцеловал его. И ощутил [Исаак] запах от одежды его и благословил его и сказал: вот, запах от сына моего, как запах от поля, которое благословил Господь;
GEN|27|28|да даст тебе Бог от росы небесной и от тука земли, и множество хлеба и вина;
GEN|27|29|да послужат тебе народы, и да поклонятся тебе племена; будь господином над братьями твоими, и да поклонятся тебе сыны матери твоей; проклинающие тебя – прокляты; благословляющие тебя – благословенны!
GEN|27|30|Как скоро совершил Исаак благословение над Иаковом, и как только вышел Иаков от лица Исаака, отца своего, Исав, брат его, пришел с ловли своей.
GEN|27|31|Приготовил и он кушанье, и принес отцу своему, и сказал отцу своему: встань, отец мой, и поешь дичи сына твоего, чтобы благословила меня душа твоя.
GEN|27|32|Исаак же, отец его, сказал ему: кто ты? Он сказал: я сын твой, первенец твой, Исав.
GEN|27|33|И вострепетал Исаак весьма великим трепетом, и сказал: кто ж это, который достал дичи и принес мне, и я ел от всего, прежде нежели ты пришел, и я благословил его? он и будет благословен.
GEN|27|34|Исав, выслушав слова отца своего, поднял громкий и весьма горький вопль и сказал отцу своему: отец мой! благослови и меня.
GEN|27|35|Но он сказал: брат твой пришел с хитростью и взял благословение твое.
GEN|27|36|И сказал он: не потому ли дано ему имя: Иаков, что он запнул меня уже два раза? Он взял первородство мое, и вот, теперь взял благословение мое. И [еще] сказал: неужели ты не оставил мне благословения?
GEN|27|37|Исаак отвечал Исаву: вот, я поставил его господином над тобою и всех братьев его отдал ему в рабы; одарил его хлебом и вином; что же я сделаю для тебя, сын мой?
GEN|27|38|Но Исав сказал отцу своему: неужели, отец мой, одно у тебя благословение? благослови и меня, отец мой! И возвысил Исав голос свой и заплакал.
GEN|27|39|И отвечал Исаак, отец его, и сказал ему: вот, от тука земли будет обитание твое и от росы небесной свыше;
GEN|27|40|и ты будешь жить мечом твоим и будешь служить брату твоему; будет же [время], когда воспротивишься и свергнешь иго его с выи твоей.
GEN|27|41|И возненавидел Исав Иакова за благословение, которым благословил его отец его; и сказал Исав в сердце своем: приближаются дни плача по отце моем, и я убью Иакова, брата моего.
GEN|27|42|И пересказаны были Ревекке слова Исава, старшего сына ее; и она послала, и призвала младшего сына своего Иакова, и сказала ему: вот, Исав, брат твой, грозит убить тебя;
GEN|27|43|и теперь, сын мой, послушайся слов моих, встань, беги к Лавану, брату моему, в Харран,
GEN|27|44|и поживи у него несколько времени, пока утолится ярость брата твоего,
GEN|27|45|пока утолится гнев брата твоего на тебя, и он позабудет, что ты сделал ему: тогда я пошлю и возьму тебя оттуда; для чего мне в один день лишиться обоих вас?
GEN|27|46|И сказала Ревекка Исааку: я жизни не рада от дочерей Хеттейских; если Иаков возьмет жену из дочерей Хеттейских, каковы эти, из дочерей этой земли, то к чему мне и жизнь?
GEN|28|1|И призвал Исаак Иакова и благословил его, и заповедал ему и сказал: не бери себе жены из дочерей Ханаанских;
GEN|28|2|встань, пойди в Месопотамию, в дом Вафуила, отца матери твоей, и возьми себе жену оттуда, из дочерей Лавана, брата матери твоей;
GEN|28|3|Бог же Всемогущий да благословит тебя, да расплодит тебя и да размножит тебя, и да будет от тебя множество народов,
GEN|28|4|и да даст тебе благословение Авраама, тебе и потомству твоему с тобою, чтобы тебе наследовать землю странствования твоего, которую Бог дал Аврааму!
GEN|28|5|И отпустил Исаак Иакова, и он пошел в Месопотамию к Лавану, сыну Вафуила Арамеянина, к брату Ревекки, матери Иакова и Исава.
GEN|28|6|Исав увидел, что Исаак благословил Иакова и благословляя послал его в Месопотамию, взять себе жену оттуда, и заповедал ему, сказав: не бери жены из дочерей Ханаанских;
GEN|28|7|и что Иаков послушался отца своего и матери своей и пошел в Месопотамию.
GEN|28|8|И увидел Исав, что дочери Ханаанские не угодны Исааку, отцу его;
GEN|28|9|и пошел Исав к Измаилу и взял себе жену Махалафу, дочь Измаила, сына Авраамова, сестру Наваиофову, сверх [других] жен своих.
GEN|28|10|Иаков же вышел из Вирсавии и пошел в Харран,
GEN|28|11|и пришел на [одно] место, и [остался] там ночевать, потому что зашло солнце. И взял [один] из камней того места, и положил себе изголовьем, и лег на том месте.
GEN|28|12|И увидел во сне: вот, лестница стоит на земле, а верх ее касается неба; и вот, Ангелы Божии восходят и нисходят по ней.
GEN|28|13|И вот, Господь стоит на ней и говорит: Я Господь, Бог Авраама, отца твоего, и Бог Исаака. Землю, на которой ты лежишь, Я дам тебе и потомству твоему;
GEN|28|14|и будет потомство твое, как песок земной; и распространишься к морю и к востоку, и к северу и к полудню; и благословятся в тебе и в семени твоем все племена земные;
GEN|28|15|и вот Я с тобою, и сохраню тебя везде, куда ты ни пойдешь; и возвращу тебя в сию землю, ибо Я не оставлю тебя, доколе не исполню того, что Я сказал тебе.
GEN|28|16|Иаков пробудился от сна своего и сказал: истинно Господь присутствует на месте сем; а я не знал!
GEN|28|17|И убоялся и сказал: как страшно сие место! это не иное что, как дом Божий, это врата небесные.
GEN|28|18|И встал Иаков рано утром, и взял камень, который он положил себе изголовьем, и поставил его памятником, и возлил елей на верх его.
GEN|28|19|И нарек имя месту тому: Вефиль, а прежнее имя того города было: Луз.
GEN|28|20|И положил Иаков обет, сказав: если Бог будет со мною и сохранит меня в пути сем, в который я иду, и даст мне хлеб есть и одежду одеться,
GEN|28|21|и я в мире возвращусь в дом отца моего, и будет Господь моим Богом, –
GEN|28|22|то этот камень, который я поставил памятником, будет домом Божиим; и из всего, что Ты, [Боже], даруешь мне, я дам Тебе десятую часть.
GEN|29|1|И встал Иаков и пошел в землю сынов востока.
GEN|29|2|И увидел: вот, на поле колодезь, и там три стада мелкого скота, лежавшие около него, потому что из того колодезя поили стада. Над устьем колодезя был большой камень.
GEN|29|3|Когда собирались туда все стада, отваливали камень от устья колодезя и поили овец; потом опять клали камень на свое место, на устье колодезя.
GEN|29|4|Иаков сказал им: братья мои! откуда вы? Они сказали: мы из Харрана.
GEN|29|5|Он сказал им: знаете ли вы Лавана, сына Нахорова? Они сказали: знаем.
GEN|29|6|Он еще сказал им: здравствует ли он? Они сказали: здравствует; и вот, Рахиль, дочь его, идет с овцами.
GEN|29|7|И сказал: вот, дня еще много; не время собирать скот; напойте овец и пойдите, пасите.
GEN|29|8|Они сказали: не можем, пока не соберутся все стада, и не отвалят камня от устья колодезя; тогда будем мы поить овец.
GEN|29|9|Еще он говорил с ними, как пришла Рахиль с мелким скотом отца своего, потому что она пасла.
GEN|29|10|Когда Иаков увидел Рахиль, дочь Лавана, брата матери своей, и овец Лавана, брата матери своей, то подошел Иаков, отвалил камень от устья колодезя и напоил овец Лавана, брата матери своей.
GEN|29|11|И поцеловал Иаков Рахиль и возвысил голос свой и заплакал.
GEN|29|12|И сказал Иаков Рахили, что он родственник отцу ее и что он сын Ревеккин. А она побежала и сказала отцу своему.
GEN|29|13|Лаван, услышав о Иакове, сыне сестры своей, выбежал ему навстречу, обнял его и поцеловал его, и ввел его в дом свой; и он рассказал Лавану все сие.
GEN|29|14|Лаван же сказал ему: подлинно ты кость моя и плоть моя. И жил у него [Иаков] целый месяц.
GEN|29|15|И Лаван сказал Иакову: неужели ты даром будешь служить мне, потому что ты родственник? скажи мне, что заплатить тебе?
GEN|29|16|У Лавана же было две дочери; имя старшей: Лия; имя младшей: Рахиль.
GEN|29|17|Лия была слаба глазами, а Рахиль была красива станом и красива лицем.
GEN|29|18|Иаков полюбил Рахиль и сказал: я буду служить тебе семь лет за Рахиль, младшую дочь твою.
GEN|29|19|Лаван сказал: лучше отдать мне ее за тебя, нежели отдать ее за другого кого; живи у меня.
GEN|29|20|И служил Иаков за Рахиль семь лет; и они показались ему за несколько дней, потому что он любил ее.
GEN|29|21|И сказал Иаков Лавану: дай жену мою, потому что мне уже исполнилось время, чтобы войти к ней.
GEN|29|22|Лаван созвал всех людей того места и сделал пир.
GEN|29|23|Вечером же взял дочь свою Лию и ввел ее к нему; и вошел к ней [Иаков].
GEN|29|24|И дал Лаван служанку свою Зелфу в служанки дочери своей Лии.
GEN|29|25|Утром же оказалось, что это Лия. И сказал Лавану: что это сделал ты со мною? не за Рахиль ли я служил у тебя? зачем ты обманул меня?
GEN|29|26|Лаван сказал: в нашем месте так не делают, чтобы младшую выдать прежде старшей;
GEN|29|27|окончи неделю этой, потом дадим тебе и ту за службу, которую ты будешь служить у меня еще семь лет других.
GEN|29|28|Иаков так и сделал и окончил неделю этой. И [Лаван] дал Рахиль, дочь свою, ему в жену.
GEN|29|29|И дал Лаван служанку свою Валлу в служанки дочери своей Рахили.
GEN|29|30|[Иаков] вошел и к Рахили, и любил Рахиль больше, нежели Лию; и служил у него еще семь лет других.
GEN|29|31|Господь узрел, что Лия была нелюбима, и отверз утробу ее, а Рахиль была неплодна.
GEN|29|32|Лия зачала и родила сына, и нарекла ему имя: Рувим, потому что сказала она: Господь призрел на мое бедствие; ибо теперь будет любить меня муж мой.
GEN|29|33|И зачала опять и родила сына, и сказала: Господь услышал, что я нелюбима, и дал мне и сего. И нарекла ему имя: Симеон.
GEN|29|34|И зачала еще и родила сына, и сказала: теперь–то прилепится ко мне муж мой, ибо я родила ему трех сынов. От сего наречено ему имя: Левий.
GEN|29|35|И еще зачала и родила сына, и сказала: теперь–то я восхвалю Господа. Посему нарекла ему имя Иуда. И перестала рождать.
GEN|30|1|И увидела Рахиль, что она не рождает детей Иакову, и позавидовала Рахиль сестре своей, и сказала Иакову: дай мне детей, а если не так, я умираю.
GEN|30|2|Иаков разгневался на Рахиль и сказал: разве я Бог, Который не дал тебе плода чрева?
GEN|30|3|Она сказала: вот служанка моя Валла; войди к ней; пусть она родит на колени мои, чтобы и я имела детей от нее.
GEN|30|4|И дала она Валлу, служанку свою, в жену ему; и вошел к ней Иаков.
GEN|30|5|Валла зачала и родила Иакову сына.
GEN|30|6|И сказала Рахиль: судил мне Бог, и услышал голос мой, и дал мне сына. Посему нарекла ему имя: Дан.
GEN|30|7|И еще зачала и родила Валла, служанка Рахилина, другого сына Иакову.
GEN|30|8|И сказала Рахиль: борьбою сильною боролась я с сестрою моею и превозмогла. И нарекла ему имя: Неффалим.
GEN|30|9|Лия увидела, что перестала рождать, и взяла служанку свою Зелфу, и дала ее Иакову в жену.
GEN|30|10|И Зелфа, служанка Лиина, родила Иакову сына.
GEN|30|11|И сказала Лия: прибавилось. И нарекла ему имя: Гад.
GEN|30|12|И родила Зелфа, служанка Лии, другого сына Иакову.
GEN|30|13|И сказала Лия: к благу моему, ибо блаженною будут называть меня женщины. И нарекла ему имя: Асир.
GEN|30|14|Рувим пошел во время жатвы пшеницы, и нашел мандрагоровые яблоки в поле, и принес их Лии, матери своей. И Рахиль сказала Лии: дай мне мандрагоров сына твоего.
GEN|30|15|Но она сказала ей: неужели мало тебе завладеть мужем моим, что ты домогаешься и мандрагоров сына моего? Рахиль сказала: так пусть он ляжет с тобою эту ночь, за мандрагоры сына твоего.
GEN|30|16|Иаков пришел с поля вечером, и Лия вышла ему навстречу и сказала: войди ко мне; ибо я купила тебя за мандрагоры сына моего. И лег он с нею в ту ночь.
GEN|30|17|И услышал Бог Лию, и она зачала и родила Иакову пятого сына.
GEN|30|18|И сказала Лия: Бог дал возмездие мне за то, что я отдала служанку мою мужу моему. И нарекла ему имя: Иссахар.
GEN|30|19|И еще зачала Лия и родила Иакову шестого сына.
GEN|30|20|И сказала Лия: Бог дал мне прекрасный дар; теперь будет жить у меня муж мой, ибо я родила ему шесть сынов. И нарекла ему имя: Завулон.
GEN|30|21|Потом родила дочь и нарекла ей имя: Дина.
GEN|30|22|И вспомнил Бог о Рахили, и услышал ее Бог, и отверз утробу ее.
GEN|30|23|Она зачала и родила сына, и сказала: снял Бог позор мой.
GEN|30|24|И нарекла ему имя: Иосиф, сказав: Господь даст мне и другого сына.
GEN|30|25|После того, как Рахиль родила Иосифа, Иаков сказал Лавану: отпусти меня, и пойду я в свое место, и в свою землю;
GEN|30|26|отдай жен моих и детей моих, за которых я служил тебе, и я пойду, ибо ты знаешь службу мою, какую я служил тебе.
GEN|30|27|И сказал ему Лаван: о, если бы я нашел благоволение пред очами твоими! я примечаю, что за тебя Господь благословил меня.
GEN|30|28|И сказал: назначь себе награду от меня, и я дам.
GEN|30|29|И сказал ему [Иаков]: ты знаешь, как я служил тебе, и каков стал скот твой при мне;
GEN|30|30|ибо мало было у тебя до меня, а стало много; Господь благословил тебя с приходом моим; когда же я буду работать для своего дома?
GEN|30|31|И сказал [Лаван]: что дать тебе? Иаков сказал: не давай мне ничего. Если только сделаешь мне, что я скажу, то я опять буду пасти и стеречь овец твоих.
GEN|30|32|Я пройду сегодня по всему [стаду] овец твоих; отдели из него всякий скот с крапинами и с пятнами, всякую скотину черную из овец, также с пятнами и с крапинами из коз. [Такой скот] будет наградою мне.
GEN|30|33|И будет говорить за меня пред тобою справедливость моя в следующее время, когда придешь посмотреть награду мою. Всякая из коз не с крапинами и не с пятнами, и из овец не черная, краденое это у меня.
GEN|30|34|Лаван сказал: хорошо, пусть будет по твоему слову.
GEN|30|35|И отделил в тот день козлов пестрых и с пятнами, и всех коз с крапинами и с пятнами, всех, на которых было [несколько] белого, и всех черных овец, и отдал на руки сыновьям своим;
GEN|30|36|и назначил расстояние между собою и между Иаковом на три дня пути. Иаков же пас остальной мелкий скот Лаванов.
GEN|30|37|И взял Иаков свежих прутьев тополевых, миндальных и яворовых, и вырезал на них белые полосы, сняв кору до белизны, которая на прутьях,
GEN|30|38|и положил прутья с нарезкою перед скотом в водопойных корытах, куда скот приходил пить, и где, приходя пить, зачинал пред прутьями.
GEN|30|39|И зачинал скот пред прутьями, и рождался скот пестрый, и с крапинами, и с пятнами.
GEN|30|40|И отделял Иаков ягнят и ставил скот лицем к пестрому и всему черному скоту Лаванову; и держал свои стада особо и не ставил их вместе со скотом Лавана.
GEN|30|41|Каждый раз, когда зачинал скот крепкий, Иаков клал прутья в корытах пред глазами скота, чтобы он зачинал пред прутьями.
GEN|30|42|А когда зачинал скот слабый, тогда он не клал. И доставался слабый [скот] Лавану, а крепкий Иакову.
GEN|30|43|И сделался этот человек весьма, весьма богатым, и было у него множество мелкого скота, и рабынь, и рабов, и верблюдов, и ослов.
GEN|31|1|И услышал [Иаков] слова сынов Лавановых, которые говорили: Иаков завладел всем, что было у отца нашего, и из имения отца нашего составил все богатство сие.
GEN|31|2|И увидел Иаков лице Лавана, и вот, оно не таково к нему, как было вчера и третьего дня.
GEN|31|3|И сказал Господь Иакову: возвратись в землю отцов твоих и на родину твою; и Я буду с тобою.
GEN|31|4|И послал Иаков, и призвал Рахиль и Лию в поле, к [стаду] мелкого скота своего,
GEN|31|5|и сказал им: я вижу лице отца вашего, что оно ко мне не таково, как было вчера и третьего дня; но Бог отца моего был со мною;
GEN|31|6|вы сами знаете, что я всеми силами служил отцу вашему,
GEN|31|7|а отец ваш обманывал меня и раз десять переменял награду мою; но Бог не попустил ему сделать мне зло.
GEN|31|8|Когда сказал он, что [скот] с крапинами будет тебе в награду, то скот весь родил с крапинами. А когда он сказал: пестрые будут тебе в награду, то скот весь и родил пестрых.
GEN|31|9|И отнял Бог скот у отца вашего и дал мне.
GEN|31|10|Однажды в такое время, когда скот зачинает, я взглянул и увидел во сне, и вот козлы, поднявшиеся на скот, пестрые с крапинами и пятнами.
GEN|31|11|Ангел Божий сказал мне во сне: Иаков! Я сказал: вот я.
GEN|31|12|Он сказал: возведи очи твои и посмотри: все козлы, поднявшиеся на скот, пестрые, с крапинами и с пятнами, ибо Я вижу все, что Лаван делает с тобою;
GEN|31|13|Я Бог [явившийся тебе] в Вефиле, где ты возлил елей на памятник и где ты дал Мне обет; теперь встань, выйди из земли сей и возвратись в землю родины твоей.
GEN|31|14|Рахиль и Лия сказали ему в ответ: есть ли еще нам доля и наследство в доме отца нашего?
GEN|31|15|не за чужих ли он нас почитает? ибо он продал нас и съел даже серебро наше;
GEN|31|16|посему все богатство, которое Бог отнял у отца нашего, есть наше и детей наших; итак делай все, что Бог сказал тебе.
GEN|31|17|И встал Иаков, и посадил детей своих и жен своих на верблюдов,
GEN|31|18|и взял с собою весь скот свой и все богатство свое, которое приобрел, скот собственный его, который он приобрел в Месопотамии, чтобы идти к Исааку, отцу своему, в землю Ханаанскую.
GEN|31|19|И как Лаван пошел стричь скот свой, то Рахиль похитила идолов, которые были у отца ее.
GEN|31|20|Иаков же похитил сердце у Лавана Арамеянина, потому что не известил его, что удаляется.
GEN|31|21|И ушел со всем, что у него было; и, встав, перешел реку и направился к горе Галаад.
GEN|31|22|На третий день сказали Лавану, что Иаков ушел.
GEN|31|23|Тогда он взял с собою родственников своих, и гнался за ним семь дней, и догнал его на горе Галаад.
GEN|31|24|И пришел Бог к Лавану Арамеянину ночью во сне и сказал ему: берегись, не говори Иакову ни доброго, ни худого.
GEN|31|25|И догнал Лаван Иакова; Иаков же поставил шатер свой на горе, и Лаван со сродниками своими поставил на горе Галаад.
GEN|31|26|И сказал Лаван Иакову: что ты сделал? для чего ты обманул меня, и увел дочерей моих, как плененных оружием?
GEN|31|27|зачем ты убежал тайно, и укрылся от меня, и не сказал мне? я отпустил бы тебя с веселием и с песнями, с тимпаном и с гуслями;
GEN|31|28|ты не позволил мне даже поцеловать внуков моих и дочерей моих; безрассудно ты сделал.
GEN|31|29|Есть в руке моей сила сделать вам зло; но Бог отца вашего вчера говорил ко мне и сказал: берегись, не говори Иакову ни хорошего, ни худого.
GEN|31|30|Но пусть бы ты ушел, потому что ты нетерпеливо захотел быть в доме отца твоего, – зачем ты украл богов моих?
GEN|31|31|Иаков отвечал Лавану и сказал: [я] боялся, ибо я думал, не отнял бы ты у меня дочерей своих.
GEN|31|32|у кого найдешь богов твоих, тот не будет жив; при родственниках наших узнавай, что у меня, и возьми себе. Иаков не знал, что Рахиль украла их.
GEN|31|33|И ходил Лаван в шатер Иакова, и в шатер Лии, и в шатер двух рабынь, но не нашел. И, выйдя из шатра Лии, вошел в шатер Рахили.
GEN|31|34|Рахиль же взяла идолов, и положила их под верблюжье седло и села на них. И обыскал Лаван весь шатер; но не нашел.
GEN|31|35|Она же сказала отцу своему: да не прогневается господин мой, что я не могу встать пред тобою, ибо у меня обыкновенное женское. И он искал, но не нашел идолов.
GEN|31|36|Иаков рассердился и вступил в спор с Лаваном. И начал Иаков говорить и сказал Лавану: какая вина моя, какой грех мой, что ты преследуешь меня?
GEN|31|37|ты осмотрел у меня все вещи, что нашел ты из всех вещей твоего дома? покажи здесь пред родственниками моими и пред родственниками твоими; пусть они рассудят между нами обоими.
GEN|31|38|Вот, двадцать лет я [был] у тебя; овцы твои и козы твои не выкидывали; овнов стада твоего я не ел;
GEN|31|39|растерзанного зверем я не приносил к тебе, это был мой убыток; ты с меня взыскивал, днем ли что пропадало, ночью ли пропадало;
GEN|31|40|я томился днем от жара, а ночью от стужи, и сон мой убегал от глаз моих.
GEN|31|41|Таковы мои двадцать лет в доме твоем. Я служил тебе четырнадцать лет за двух дочерей твоих и шесть лет за скот твой, а ты десять раз переменял награду мою.
GEN|31|42|Если бы не был со мною Бог отца моего, Бог Авраама и страх Исаака, ты бы теперь отпустил меня ни с чем. Бог увидел бедствие мое и труд рук моих и вступился [за меня] вчера.
GEN|31|43|И отвечал Лаван и сказал Иакову: дочери – мои дочери; дети – мои дети; скот – мой скот, и все, что ты видишь, это мое: могу ли я что сделать теперь с дочерями моими и с детьми их, которые рождены ими?
GEN|31|44|Теперь заключим союз я и ты, и это будет свидетельством между мною и тобою.
GEN|31|45|И взял Иаков камень и поставил его памятником.
GEN|31|46|И сказал Иаков родственникам своим: наберите камней. Они взяли камни, и сделали холм, и ели там на холме.
GEN|31|47|И назвал его Лаван: Иегар–Сагадуфа; а Иаков назвал его Галаадом.
GEN|31|48|И сказал Лаван: сегодня этот холм между мною и тобою свидетель. Посему и наречено ему имя: Галаад,
GEN|31|49|[также]: Мицпа, от того, что Лаван сказал: да надзирает Господь надо мною и над тобою, когда мы скроемся друг от друга;
GEN|31|50|если ты будешь худо поступать с дочерями моими, или если возьмешь жен сверх дочерей моих, то, хотя нет человека между нами, но смотри, Бог свидетель между мною и между тобою.
GEN|31|51|И сказал Лаван Иакову: вот холм сей и вот памятник, который я поставил между мною и тобою;
GEN|31|52|этот холм свидетель, и этот памятник свидетель, что ни я не перейду к тебе за этот холм, ни ты не перейдешь ко мне за этот холм и за этот памятник, для зла;
GEN|31|53|Бог Авраамов и Бог Нахоров да судит между нами, Бог отца их. Иаков поклялся страхом отца своего Исаака.
GEN|31|54|И заколол Иаков жертву на горе и позвал родственников своих есть хлеб; и они ели хлеб и ночевали на горе.
GEN|32|1|И встал Лаван рано утром и поцеловал внуков своих и дочерей своих, и благословил их. И пошел и возвратился Лаван в свое место.
GEN|32|2|А Иаков пошел путем своим. И встретили его Ангелы Божии.
GEN|32|3|Иаков, увидев их, сказал: это ополчение Божие. И нарек имя месту тому: Маханаим.
GEN|32|4|И послал Иаков пред собою вестников к брату своему Исаву в землю Сеир, в область Едом,
GEN|32|5|и приказал им, сказав: так скажите господину моему Исаву: вот что говорит раб твой Иаков: я жил у Лавана и прожил доныне;
GEN|32|6|и есть у меня волы и ослы и мелкий скот, и рабы и рабыни; и я послал известить [о себе] господина моего, дабы приобрести благоволение пред очами твоими.
GEN|32|7|И возвратились вестники к Иакову и сказали: мы ходили к брату твоему Исаву; он идет навстречу тебе, и с ним четыреста человек.
GEN|32|8|Иаков очень испугался и смутился; и разделил людей, бывших с ним, и скот мелкий и крупный и верблюдов на два стана.
GEN|32|9|И сказал: если Исав нападет на один стан и побьет его, то остальной стан может спастись.
GEN|32|10|И сказал Иаков: Боже отца моего Авраама и Боже отца моего Исаака, Господи, сказавший мне: возвратись в землю твою, на родину твою, и Я буду благотворить тебе!
GEN|32|11|Недостоин я всех милостей и всех благодеяний, которые Ты сотворил рабу Твоему, ибо я с посохом моим перешел этот Иордан, а теперь у меня два стана.
GEN|32|12|Избавь меня от руки брата моего, от руки Исава, ибо я боюсь его, чтобы он, придя, не убил меня [и] матери с детьми.
GEN|32|13|Ты сказал: Я буду благотворить тебе и сделаю потомство твое, как песок морской, которого не исчислить от множества.
GEN|32|14|И ночевал там [Иаков] в ту ночь. И взял из того, что у него было, в подарок Исаву, брату своему:
GEN|32|15|двести коз, двадцать козлов, двести овец, двадцать овнов,
GEN|32|16|тридцать верблюдиц дойных с жеребятами их, сорок коров, десять волов, двадцать ослиц, десять ослов.
GEN|32|17|И дал в руки рабам своим каждое стадо особо и сказал рабам своим: пойдите предо мною и оставляйте расстояние от стада до стада.
GEN|32|18|И приказал первому, сказав: когда брат мой Исав встретится тебе и спросит тебя, говоря: чей ты? и куда идешь? и чье это [стадо] пред тобою?
GEN|32|19|то скажи: раба твоего Иакова; это подарок, посланный господину моему Исаву; вот, и сам он за нами.
GEN|32|20|То же приказал он и второму, и третьему, и всем, которые шли за стадами, говоря: так скажите Исаву, когда встретите его;
GEN|32|21|и скажите: вот, и раб твой Иаков за нами. Ибо он сказал [сам в себе]: умилостивлю его дарами, которые идут предо мною, и потом увижу лице его; может быть, и примет меня.
GEN|32|22|И пошли дары пред ним, а он ту ночь ночевал в стане.
GEN|32|23|И встал в ту ночь, и, взяв двух жен своих и двух рабынь своих, и одиннадцать сынов своих, перешел через Иавок вброд;
GEN|32|24|и, взяв их, перевел через поток, и перевел все, что у него [было].
GEN|32|25|И остался Иаков один. И боролся Некто с ним до появления зари;
GEN|32|26|и, увидев, что не одолевает его, коснулся состава бедра его и повредил состав бедра у Иакова, когда он боролся с Ним.
GEN|32|27|И сказал: отпусти Меня, ибо взошла заря. Иаков сказал: не отпущу Тебя, пока не благословишь меня.
GEN|32|28|И сказал: как имя твое? Он сказал: Иаков.
GEN|32|29|И сказал: отныне имя тебе будет не Иаков, а Израиль, ибо ты боролся с Богом, и человеков одолевать будешь.
GEN|32|30|Спросил и Иаков, говоря: скажи имя Твое. И Он сказал: на что ты спрашиваешь о имени Моем? И благословил его там.
GEN|32|31|И нарек Иаков имя месту тому: Пенуэл; ибо, [говорил он], я видел Бога лицем к лицу, и сохранилась душа моя.
GEN|32|32|И взошло солнце, когда он проходил Пенуэл; и хромал он на бедро свое.
GEN|32|33|Поэтому и доныне сыны Израилевы не едят жилы, которая на составе бедра, потому что [Боровшийся] коснулся жилы на составе бедра Иакова.
GEN|33|1|Взглянул Иаков и увидел, и вот, идет Исав, и с ним четыреста человек. И разделил детей Лии, Рахили и двух служанок.
GEN|33|2|И поставил служанок и детей их впереди, Лию и детей ее за ними, а Рахиль и Иосифа позади.
GEN|33|3|А сам пошел пред ними и поклонился до земли семь раз, подходя к брату своему.
GEN|33|4|И побежал Исав к нему навстречу и обнял его, и пал на шею его и целовал его, и плакали.
GEN|33|5|И взглянул и увидел жен и детей и сказал: кто это у тебя? [Иаков] сказал: дети, которых Бог даровал рабу твоему.
GEN|33|6|И подошли служанки и дети их и поклонились;
GEN|33|7|подошла и Лия и дети ее и поклонились; наконец подошли Иосиф и Рахиль и поклонились.
GEN|33|8|И сказал Исав: для чего у тебя это множество, которое я встретил? И сказал Иаков: дабы приобрести благоволение в очах господина моего.
GEN|33|9|Исав сказал: у меня много, брат мой; пусть будет твое у тебя.
GEN|33|10|Иаков сказал: нет, если я приобрел благоволение в очах твоих, прими дар мой от руки моей, ибо я увидел лице твое, как бы кто увидел лице Божие, и ты был благосклонен ко мне;
GEN|33|11|прими благословение мое, которое я принес тебе, потому что Бог даровал мне, и есть у меня все. И упросил его, и тот взял
GEN|33|12|и сказал: поднимемся и пойдем; и я пойду пред тобою.
GEN|33|13|Иаков сказал ему: господин мой знает, что дети нежны, а мелкий и крупный скот у меня дойный: если погнать его один день, то помрет весь скот;
GEN|33|14|пусть господин мой пойдет впереди раба своего, а я пойду медленно, как пойдет скот, который предо мною, и как пойдут дети, и приду к господину моему в Сеир.
GEN|33|15|Исав сказал: оставлю я с тобою [несколько] из людей, которые при мне. Иаков сказал: к чему это? только бы мне приобрести благоволение в очах господина моего!
GEN|33|16|И возвратился Исав в тот же день путем своим в Сеир.
GEN|33|17|А Иаков двинулся в Сокхоф, и построил себе дом, и для скота своего сделал шалаши. От сего он нарек имя месту: Сокхоф.
GEN|33|18|Иаков, возвратившись из Месопотамии, благополучно пришел в город Сихем, который в земле Ханаанской, и расположился пред городом.
GEN|33|19|И купил часть поля, на котором раскинул шатер свой, у сынов Еммора, отца Сихемова, за сто монет.
GEN|33|20|И поставил там жертвенник, и призвал имя Господа Бога Израилева.
GEN|34|1|Дина, дочь Лии, которую она родила Иакову, вышла посмотреть на дочерей земли той.
GEN|34|2|И увидел ее Сихем, сын Еммора Евеянина, князя земли той, и взял ее, и спал с нею, и сделал ей насилие.
GEN|34|3|И прилепилась душа его в Дине, дочери Иакова, и он полюбил девицу и говорил по сердцу девицы.
GEN|34|4|И сказал Сихем Еммору, отцу своему, говоря: возьми мне эту девицу в жену.
GEN|34|5|Иаков слышал, что [сын Емморов] обесчестил Дину, дочь его, но как сыновья его были со скотом его в поле, то Иаков молчал, пока не пришли они.
GEN|34|6|И вышел Еммор, отец Сихемов, к Иакову, поговорить с ним.
GEN|34|7|Сыновья же Иакова пришли с поля, и когда услышали, то огорчились мужи те и воспылали гневом, потому что бесчестие сделал он Израилю, переспав с дочерью Иакова, а так не надлежало делать.
GEN|34|8|Еммор стал говорить им, и сказал: Сихем, сын мой, прилепился душею к дочери вашей; дайте же ее в жену ему;
GEN|34|9|породнитесь с нами; отдавайте за нас дочерей ваших, а наших дочерей берите себе.
GEN|34|10|и живите с нами; земля сия пред вами, живите и промышляйте на ней и приобретайте ее во владение.
GEN|34|11|Сихем же сказал отцу ее и братьям ее: только бы мне найти благоволение в очах ваших, я дам, что ни скажете мне;
GEN|34|12|назначьте самое большое вено и дары; я дам, что ни скажете мне, только отдайте мне девицу в жену.
GEN|34|13|И отвечали сыновья Иакова Сихему и Еммору, отцу его, с лукавством; а говорили так потому, что он обесчестил Дину, сестру их;
GEN|34|14|и сказали им: не можем этого сделать, выдать сестру нашу за человека, который необрезан, ибо это бесчестно для нас;
GEN|34|15|только на том условии мы согласимся с вами, если вы будете как мы, чтобы и у вас весь мужеский пол был обрезан;
GEN|34|16|и будем отдавать за вас дочерей наших и брать за себя ваших дочерей, и будем жить с вами, и составим один народ;
GEN|34|17|а если не послушаетесь нас в том, чтобы обрезаться, то мы возьмем дочь нашу и удалимся.
GEN|34|18|И понравились слова сии Еммору и Сихему, сыну Емморову.
GEN|34|19|Юноша не умедлил исполнить это, потому что любил дочь Иакова. А он более всех уважаем был из дома отца своего.
GEN|34|20|И пришел Еммор и Сихем, сын его, к воротам города своего, и стали говорить жителям города своего и сказали:
GEN|34|21|сии люди мирны с нами; пусть они селятся на земле и промышляют на ней; земля же вот пространна пред ними. Станем брать дочерей их себе в жены и наших дочерей выдавать за них.
GEN|34|22|Только на том условии сии люди соглашаются жить с нами и быть одним народом, чтобы и у нас обрезан был весь мужеский пол, как они обрезаны.
GEN|34|23|Не для нас ли стада их, и имение их, и весь скот их? Только согласимся с ними, и будут жить с нами.
GEN|34|24|И послушались Еммора и Сихема, сына его, все выходящие из ворот города его: и обрезан был весь мужеский пол, – все выходящие из ворот города его.
GEN|34|25|На третий день, когда они были в болезни, два сына Иакова, Симеон и Левий, братья Динины, взяли каждый свой меч, и смело напали на город, и умертвили весь мужеский пол;
GEN|34|26|и самого Еммора и Сихема, сына его, убили мечом; и взяли Дину из дома Сихемова и вышли.
GEN|34|27|Сыновья Иакова пришли к убитым и разграбили город за то, что обесчестили сестру их.
GEN|34|28|Они взяли мелкий и крупный скот их, и ослов их, и что ни было в городе, и что ни было в поле;
GEN|34|29|и все богатство их, и всех детей их, и жен их взяли в плен, и разграбили все, что было в домах.
GEN|34|30|И сказал Иаков Симеону и Левию: вы возмутили меня, сделав меня ненавистным для жителей сей земли, для Хананеев и Ферезеев. У меня людей мало; соберутся против меня, поразят меня, и истреблен буду я и дом мой.
GEN|34|31|Они же сказали: а разве можно поступать с сестрою нашею, как с блудницею!
GEN|35|1|Бог сказал Иакову: встань, пойди в Вефиль и живи там, и устрой там жертвенник Богу, явившемуся тебе, когда ты бежал от лица Исава, брата твоего.
GEN|35|2|И сказал Иаков дому своему и всем бывшим с ним: бросьте богов чужих, находящихся у вас, и очиститесь, и перемените одежды ваши;
GEN|35|3|встанем и пойдем в Вефиль; там устрою я жертвенник Богу, Который услышал меня в день бедствия моего и был со мною в пути, которым я ходил.
GEN|35|4|И отдали Иакову всех богов чужих, бывших в руках их, и серьги, бывшие в ушах у них, и закопал их Иаков под дубом, который близ Сихема.
GEN|35|5|И отправились они. И был ужас Божий на окрестных городах, и не преследовали сынов Иаковлевых.
GEN|35|6|И пришел Иаков в Луз, что в земле Ханаанской, то есть в Вефиль, сам и все люди, бывшие с ним,
GEN|35|7|и устроил там жертвенник, и назвал сие место: Эл–Вефиль, ибо тут явился ему Бог, когда он бежал от лица брата своего.
GEN|35|8|И умерла Девора, кормилица Ревеккина, и погребена ниже Вефиля под дубом, который и назвал [Иаков] дубом плача.
GEN|35|9|И явился Бог Иакову по возвращении его из Месопотамии, и благословил его,
GEN|35|10|и сказал ему Бог: имя твое Иаков; отныне ты не будешь называться Иаковом, но будет имя тебе: Израиль. И нарек ему имя: Израиль.
GEN|35|11|И сказал ему Бог: Я Бог Всемогущий; плодись и умножайся; народ и множество народов будет от тебя, и цари произойдут из чресл твоих;
GEN|35|12|землю, которую Я дал Аврааму и Исааку, Я дам тебе, и потомству твоему по тебе дам землю сию.
GEN|35|13|И восшел от него Бог с места, на котором говорил ему.
GEN|35|14|И поставил Иаков памятник на месте, на котором говорил ему [Бог], памятник каменный, и возлил на него возлияние, и возлил на него елей;
GEN|35|15|и нарек Иаков имя месту, на котором Бог говорил ему: Вефиль.
GEN|35|16|И отправились из Вефиля. И когда еще оставалось некоторое расстояние земли до Ефрафы, Рахиль родила, и роды ее были трудны.
GEN|35|17|Когда же она страдала в родах, повивальная бабка сказала ей: не бойся, ибо и это тебе сын.
GEN|35|18|И когда выходила из нее душа, ибо она умирала, то нарекла ему имя: Бенони. Но отец его назвал его Вениамином.
GEN|35|19|И умерла Рахиль, и погребена на дороге в Ефрафу, то есть Вифлеем.
GEN|35|20|Иаков поставил над гробом ее памятник. Это надгробный памятник Рахили до сего дня.
GEN|35|21|И отправился Израиль и раскинул шатер свой за башнею Гадер.
GEN|35|22|Во время пребывания Израиля в той стране, Рувим пошел и переспал с Валлою, наложницею отца своего. И услышал Израиль. Сынов же у Иакова было двенадцать.
GEN|35|23|Сыновья Лии: первенец Иакова Рувим, [по нем] Симеон, Левий, Иуда, Иссахар и Завулон.
GEN|35|24|Сыновья Рахили: Иосиф и Вениамин.
GEN|35|25|Сыновья Валлы, служанки Рахилиной: Дан и Неффалим.
GEN|35|26|Сыновья Зелфы, служанки Лииной: Гад и Асир. Сии сыновья Иакова, родившиеся ему в Месопотамии.
GEN|35|27|И пришел Иаков к Исааку, отцу своему, в Мамре, в Кириаф–Арбу, то есть Хеврон где странствовал Авраам и Исаак.
GEN|35|28|И было дней [жизни] Исааковой сто восемьдесят лет.
GEN|35|29|И испустил Исаак дух и умер, и приложился к народу своему, будучи стар и насыщен жизнью; и погребли его Исав и Иаков, сыновья его.
GEN|36|1|Вот родословие Исава, он же Едом.
GEN|36|2|Исав взял себе жен из дочерей Ханаанских: Аду, дочь Елона Хеттеянина, и Оливему, дочь Аны, сына Цивеона Евеянина,
GEN|36|3|и Васемафу, дочь Измаила, сестру Наваиофа.
GEN|36|4|Ада родила Исаву Елифаза, Васемафа родила Рагуила,
GEN|36|5|Оливема родила Иеуса, Иеглома и Корея. Это сыновья Исава, родившиеся ему в земле Ханаанской.
GEN|36|6|И взял Исав жен своих и сыновей своих, и дочерей своих, и всех людей дома своего, и стада свои, и весь скот свой, и все имение свое, которое он приобрел в земле Ханаанской, и пошел в [другую] землю от лица Иакова, брата своего,
GEN|36|7|ибо имение их было так велико, что они не могли жить вместе, и земля странствования их не вмещала их, по множеству стад их.
GEN|36|8|И поселился Исав на горе Сеир, Исав, он же Едом.
GEN|36|9|И вот родословие Исава, отца Идумеев, на горе Сеир.
GEN|36|10|Вот имена сынов Исава: Елифаз, сын Ады, жены Исавовой, и Рагуил, сын Васемафы, жены Исавовой.
GEN|36|11|У Елифаза были сыновья: Феман, Омар, Цефо, Гафам и Кеназ.
GEN|36|12|Фамна же была наложница Елифаза, сына Исавова, и родила Елифазу Амалика. Вот сыновья Ады, жены Исавовой.
GEN|36|13|И вот сыновья Рагуила: Нахаф и Зерах, Шамма и Миза. Это сыновья Васемафы, жены Исавовой.
GEN|36|14|И сии были сыновья Оливемы, дочери Аны, сына Цивеонова, жены Исавовой: она родила Исаву Иеуса, Иеглома и Корея.
GEN|36|15|Вот старейшины сынов Исавовых. Сыновья Елифаза, первенца Исавова: старейшина Феман, старейшина Омар, старейшина Цефо, старейшина Кеназ,
GEN|36|16|старейшина Корей, старейшина Гафам, старейшина Амалик. Сии старейшины Елифазовы в земле Едома; сии сыновья Ады.
GEN|36|17|Сии сыновья Рагуила, сына Исавова: старейшина Нахаф, старейшина Зерах, старейшина Шамма, старейшина Миза. Сии старейшины Рагуиловы в земле Едома; сии сыновья Васемафы, жены Исавовой.
GEN|36|18|Сии сыновья Оливемы, жены Исавовой: старейшина Иеус, старейшина Иеглом, старейшина Корей. Сии старейшины Оливемы, дочери Аны, жены Исавовой.
GEN|36|19|Вот сыновья Исава, и вот старейшины их. Это Едом.
GEN|36|20|Сии сыновья Сеира Хорреянина, жившие в земле той: Лотан, Шовал, Цивеон, Ана,
GEN|36|21|Дишон, Эцер и Дишан. Сии старейшины Хорреев, сынов Сеира, в земле Едома.
GEN|36|22|Сыновья Лотана были: Хори и Геман; а сестра у Лотана: Фамна.
GEN|36|23|Сии сыновья Шовала: Алван, Манахаф, Эвал, Шефо и Онам.
GEN|36|24|Сии сыновья Цивеона: Аиа и Ана. Это тот Ана, который нашел теплые воды в пустыне, когда пас ослов Цивеона, отца своего.
GEN|36|25|Сии дети Аны: Дишон и Оливема, дочь Аны.
GEN|36|26|Сии сыновья Дишона: Хемдан, Эшбан, Ифран и Херан.
GEN|36|27|Сии сыновья Эцера: Билган, Зааван, и Акан.
GEN|36|28|Сии сыновья Дишана: Уц и Аран.
GEN|36|29|Сии старейшины Хорреев: старейшина Лотан, старейшина Шовал, старейшина Цивеон, старейшина Ана,
GEN|36|30|старейшина Дишон, старейшина Эцер, старейшина Дишан. Вот старейшины Хорреев, по старшинствам их в земле Сеир.
GEN|36|31|Вот цари, царствовавшие в земле Едома, прежде царствования царей у сынов Израилевых:
GEN|36|32|царствовал в Едоме Бела, сын Веоров, а имя городу его Дингава.
GEN|36|33|И умер Бела, и воцарился по нем Иовав, сын Зераха, из Восоры.
GEN|36|34|Умер Иовав, и воцарился по нем Хушам, из земли Феманитян.
GEN|36|35|И умер Хушам, и воцарился по нем Гадад, сын Бедадов, который поразил Мадианитян на поле Моава; имя городу его Авиф.
GEN|36|36|И умер Гадад, и воцарился по нем Самла из Масреки.
GEN|36|37|И умер Самла, и воцарился по нем Саул из Реховофа, что при реке.
GEN|36|38|И умер Саул, и воцарился по нем Баал–Ханан, сын Ахбора.
GEN|36|39|И умер Баал–Ханан, сын Ахбора, и воцарился по нем Гадар: имя городу его Пау; имя жене его Мегетавеель, дочь Матреды, сына Мезагава.
GEN|36|40|Сии имена старейшин Исавовых, по племенам их, по местам их, по именам их: старейшина Фимна, старейшина Алва, старейшина Иетеф,
GEN|36|41|старейшина Оливема, старейшина Эла, старейшина Пинон,
GEN|36|42|старейшина Кеназ, старейшина Феман, старейшина Мивцар,
GEN|36|43|старейшина Магдиил, старейшина Ирам. Вот старейшины Идумейские, по их селениям, в земле обладания их. Вот Исав, отец Идумеев.
GEN|37|1|Иаков жил в земле странствования отца своего, в земле Ханаанской.
GEN|37|2|Вот житие Иакова. Иосиф, семнадцати лет, пас скот вместе с братьями своими, будучи отроком, с сыновьями Валлы и с сыновьями Зелфы, жен отца своего. И доводил Иосиф худые о них слухи до отца их.
GEN|37|3|Израиль любил Иосифа более всех сыновей своих, потому что он был сын старости его, – и сделал ему разноцветную одежду.
GEN|37|4|И увидели братья его, что отец их любит его более всех братьев его; и возненавидели его и не могли говорить с ним дружелюбно.
GEN|37|5|И видел Иосиф сон, и рассказал братьям своим: и они возненавидели его еще более.
GEN|37|6|Он сказал им: выслушайте сон, который я видел:
GEN|37|7|вот, мы вяжем снопы посреди поля; и вот, мой сноп встал и стал прямо; и вот, ваши снопы стали кругом и поклонились моему снопу.
GEN|37|8|И сказали ему братья его: неужели ты будешь царствовать над нами? неужели будешь владеть нами? И возненавидели его еще более за сны его и за слова его.
GEN|37|9|И видел он еще другой сон и рассказал его братьям своим, говоря: вот, я видел еще сон: вот, солнце и луна и одиннадцать звезд поклоняются мне.
GEN|37|10|И он рассказал отцу своему и братьям своим; и побранил его отец его и сказал ему: что это за сон, который ты видел? неужели я и твоя мать, и твои братья придем поклониться тебе до земли?
GEN|37|11|Братья его досадовали на него, а отец его заметил это слово.
GEN|37|12|Братья его пошли пасти скот отца своего в Сихем.
GEN|37|13|И сказал Израиль Иосифу: братья твои не пасут ли в Сихеме? пойди, я пошлю тебя к ним. Он отвечал ему: вот я.
GEN|37|14|И сказал ему: пойди, посмотри, здоровы ли братья твои и цел ли скот, и принеси мне ответ. И послал его из долины Хевронской; и он пришел в Сихем.
GEN|37|15|И нашел его некто блуждающим в поле, и спросил его тот человек, говоря: чего ты ищешь?
GEN|37|16|Он сказал: я ищу братьев моих; скажи мне, где они пасут?
GEN|37|17|И сказал тот человек: они ушли отсюда, ибо я слышал, как они говорили: пойдем в Дофан. И пошел Иосиф за братьями своими и нашел их в Дофане.
GEN|37|18|И увидели они его издали, и прежде нежели он приблизился к ним, стали умышлять против него, чтобы убить его.
GEN|37|19|И сказали друг другу: вот, идет сновидец;
GEN|37|20|пойдем теперь, и убьем его, и бросим его в какой–нибудь ров, и скажем, что хищный зверь съел его; и увидим, что будет из его снов.
GEN|37|21|И услышал [сие] Рувим и избавил его от рук их, сказав: не убьем его.
GEN|37|22|И сказал им Рувим: не проливайте крови; бросьте его в ров, который в пустыне, а руки не налагайте на него. [Сие говорил он], чтобы избавить его от рук их и возвратить его к отцу его.
GEN|37|23|Когда Иосиф пришел к братьям своим, они сняли с Иосифа одежду его, одежду разноцветную, которая была на нем,
GEN|37|24|и взяли его и бросили его в ров; ров же тот был пуст; воды в нем не было.
GEN|37|25|И сели они есть хлеб, и, взглянув, увидели, вот, идет из Галаада караван Измаильтян, и верблюды их несут стираксу, бальзам и ладан: идут они отвезти это в Египет.
GEN|37|26|И сказал Иуда братьям своим: что пользы, если мы убьем брата нашего и скроем кровь его?
GEN|37|27|Пойдем, продадим его Измаильтянам, а руки наши да не будут на нем, ибо он брат наш, плоть наша. Братья его послушались
GEN|37|28|и, когда проходили купцы Мадиамские, вытащили Иосифа изо рва и продали Иосифа Измаильтянам за двадцать сребренников; а они отвели Иосифа в Египет.
GEN|37|29|Рувим же пришел опять ко рву; и вот, нет Иосифа во рве. И разодрал он одежды свои,
GEN|37|30|и возвратился к братьям своим, и сказал: отрока нет, а я, куда я денусь?
GEN|37|31|И взяли одежду Иосифа, и закололи козла, и вымарали одежду кровью;
GEN|37|32|и послали разноцветную одежду, и доставили к отцу своему, и сказали: мы это нашли; посмотри, сына ли твоего эта одежда, или нет.
GEN|37|33|Он узнал ее и сказал: [это] одежда сына моего; хищный зверь съел его; верно, растерзан Иосиф.
GEN|37|34|И разодрал Иаков одежды свои, и возложил вретище на чресла свои, и оплакивал сына своего многие дни.
GEN|37|35|И собрались все сыновья его и все дочери его, чтобы утешить его; но он не хотел утешиться и сказал: с печалью сойду к сыну моему в преисподнюю. Так оплакивал его отец его.
GEN|37|36|Мадианитяне же продали его в Египте Потифару, царедворцу фараонову, начальнику телохранителей.
GEN|38|1|В то время Иуда отошел от братьев своих и поселился близ одного Одолламитянина, которому имя: Хира.
GEN|38|2|И увидел там Иуда дочь одного Хананеянина, которому имя: Шуа; и взял ее и вошел к ней.
GEN|38|3|Она зачала и родила сына; и он нарек ему имя: Ир.
GEN|38|4|И зачала опять, и родила сына, и нарекла ему имя: Онан.
GEN|38|5|И еще родила сына и нарекла ему имя: Шела. Иуда был в Хезиве, когда она родила его.
GEN|38|6|И взял Иуда жену Иру, первенцу своему; имя ей Фамарь.
GEN|38|7|Ир, первенец Иудин, был неугоден пред очами Господа, и умертвил его Господь.
GEN|38|8|И сказал Иуда Онану: войди к жене брата твоего, женись на ней, как деверь, и восстанови семя брату твоему.
GEN|38|9|Онан знал, что семя будет не ему, и потому, когда входил к жене брата своего, изливал на землю, чтобы не дать семени брату своему.
GEN|38|10|Зло было пред очами Господа то, что он делал; и Он умертвил и его.
GEN|38|11|И сказал Иуда Фамари, невестке своей: живи вдовою в доме отца твоего, пока подрастет Шела, сын мой. Ибо он сказал: не умер бы и он подобно братьям его. Фамарь пошла и стала жить в доме отца своего.
GEN|38|12|Прошло много времени, и умерла дочь Шуи, жена Иудина. Иуда, утешившись, пошел в Фамну к стригущим скот его, сам и Хира, друг его, Одолламитянин.
GEN|38|13|И уведомили Фамарь, говоря: вот, свекор твой идет в Фамну стричь скот свой.
GEN|38|14|И сняла она с себя одежду вдовства своего, покрыла себя покрывалом и, закрывшись, села у ворот Енаима, что на дороге в Фамну. Ибо видела, что Шела вырос, и она не дана ему в жену.
GEN|38|15|И увидел ее Иуда и почел ее за блудницу, потому что она закрыла лице свое.
GEN|38|16|Он поворотил к ней и сказал: войду я к тебе. Ибо не знал, что это невестка его. Она сказала: что ты дашь мне, если войдешь ко мне?
GEN|38|17|Он сказал: я пришлю тебе козленка из стада. Она сказала: дашь ли ты мне залог, пока пришлешь?
GEN|38|18|Он сказал: какой дать тебе залог? Она сказала: печать твою, и перевязь твою, и трость твою, которая в руке твоей. И дал он ей и вошел к ней; и она зачала от него.
GEN|38|19|И, встав, пошла, сняла с себя покрывало свое и оделась в одежду вдовства своего.
GEN|38|20|Иуда же послал козленка чрез друга своего Одолламитянина, чтобы взять залог из руки женщины, но он не нашел ее.
GEN|38|21|И спросил жителей того места, говоря: где блудница, [которая] [была] в Енаиме при дороге? Но они сказали: здесь не было блудницы.
GEN|38|22|И возвратился он к Иуде и сказал: я не нашел ее; да и жители места того сказали: здесь не было блудницы.
GEN|38|23|Иуда сказал: пусть она возьмет себе, чтобы только не стали над нами смеяться; вот, я посылал этого козленка, но ты не нашел ее.
GEN|38|24|Прошло около трех месяцев, и сказали Иуде, говоря: Фамарь, невестка твоя, впала в блуд, и вот, она беременна от блуда. Иуда сказал: выведите ее, и пусть она будет сожжена.
GEN|38|25|Но когда повели ее, она послала сказать свекру своему: я беременна от того, чьи эти вещи. И сказала: узнавай, чья эта печать и перевязь и трость.
GEN|38|26|Иуда узнал и сказал: она правее меня, потому что я не дал ее Шеле, сыну моему. И не познавал ее более.
GEN|38|27|Во время родов ее оказалось, что близнецы в утробе ее.
GEN|38|28|И во время родов ее показалась рука; и взяла повивальная бабка и навязала ему на руку красную нить, сказав: этот вышел первый.
GEN|38|29|Но он возвратил руку свою; и вот, вышел брат его. И она сказала: как ты расторг себе преграду? И наречено ему имя: Фарес.
GEN|38|30|Потом вышел брат его с красной нитью на руке. И наречено ему имя: Зара.
GEN|39|1|Иосиф же отведен был в Египет, и купил его из рук Измаильтян, приведших его туда, Египтянин Потифар, царедворец фараонов, начальник телохранителей.
GEN|39|2|И был Господь с Иосифом: он был успешен в делах и жил в доме господина своего, Египтянина.
GEN|39|3|И увидел господин его, что Господь с ним и что всему, что он делает, Господь в руках его дает успех.
GEN|39|4|И снискал Иосиф благоволение в очах его и служил ему. И он поставил его над домом своим, и все, что имел, отдал на руки его.
GEN|39|5|И с того времени, как он поставил его над домом своим и над всем, что имел, Господь благословил дом Египтянина ради Иосифа, и было благословение Господне на всем, что имел он в доме и в поле.
GEN|39|6|И оставил он все, что имел, в руках Иосифа и не знал при нем ничего, кроме хлеба, который он ел. Иосиф же был красив станом и красив лицем.
GEN|39|7|И обратила взоры на Иосифа жена господина его и сказала: спи со мною.
GEN|39|8|Но он отказался и сказал жене господина своего: вот, господин мой не знает при мне ничего в доме, и все, что имеет, отдал в мои руки;
GEN|39|9|нет больше меня в доме сем; и он не запретил мне ничего, кроме тебя, потому что ты жена ему; как же сделаю я сие великое зло и согрешу пред Богом?
GEN|39|10|Когда так она ежедневно говорила Иосифу, а он не слушался ее, чтобы спать с нею и быть с нею,
GEN|39|11|случилось в один день, что он вошел в дом делать дело свое, а никого из домашних тут в доме не было;
GEN|39|12|она схватила его за одежду его и сказала: ложись со мной. Но он, оставив одежду свою в руках ее, побежал и выбежал вон.
GEN|39|13|Она же, увидев, что он оставил одежду свою в руках ее и побежал вон,
GEN|39|14|кликнула домашних своих и сказала им так: посмотрите, он привел к нам Еврея ругаться над нами. Он пришел ко мне, чтобы лечь со мною, но я закричала громким голосом,
GEN|39|15|и он, услышав, что я подняла вопль и закричала, оставил у меня одежду свою, и побежал, и выбежал вон.
GEN|39|16|И оставила одежду его у себя до прихода господина его в дом свой.
GEN|39|17|И пересказала ему те же слова, говоря: раб Еврей, которого ты привел к нам, приходил ко мне ругаться надо мною.
GEN|39|18|но, когда я подняла вопль и закричала, он оставил у меня одежду свою и убежал вон.
GEN|39|19|Когда господин его услышал слова жены своей, которые она сказала ему, говоря: так поступил со мною раб твой, то воспылал гневом;
GEN|39|20|и взял Иосифа господин его и отдал его в темницу, где заключены узники царя. И был он там в темнице.
GEN|39|21|И Господь был с Иосифом, и простер к нему милость, и даровал ему благоволение в очах начальника темницы.
GEN|39|22|И отдал начальник темницы в руки Иосифу всех узников, находившихся в темнице, и во всем, что они там ни делали, он был распорядителем.
GEN|39|23|Начальник темницы и не смотрел ни за чем, что было у него в руках, потому что Господь был с [Иосифом], и во всем, что он делал, Господь давал успех.
GEN|40|1|После сего виночерпий царя Египетского и хлебодар провинились пред господином своим, царем Египетским.
GEN|40|2|И прогневался фараон на двух царедворцев своих, на главного виночерпия и на главного хлебодара,
GEN|40|3|и отдал их под стражу в дом начальника телохранителей, в темницу, в место, где заключен был Иосиф.
GEN|40|4|Начальник телохранителей приставил к ним Иосифа, и он служил им. И пробыли они под стражею несколько времени.
GEN|40|5|Однажды виночерпию и хлебодару царя Египетского, заключенным в темнице, виделись сны, каждому свой сон, обоим в одну ночь, каждому сон особенного значения.
GEN|40|6|И пришел к ним Иосиф поутру, увидел их, и вот, они в смущении.
GEN|40|7|И спросил он царедворцев фараоновых, находившихся с ним в доме господина его под стражею, говоря: отчего у вас сегодня печальные лица?
GEN|40|8|Они сказали ему: нам виделись сны; а истолковать их некому. Иосиф сказал им: не от Бога ли истолкования? расскажите мне.
GEN|40|9|И рассказал главный виночерпий Иосифу сон свой и сказал ему: мне снилось, вот виноградная лоза предо мною;
GEN|40|10|на лозе три ветви; она развилась, показался на ней цвет, выросли и созрели на ней ягоды;
GEN|40|11|и чаша фараонова в руке у меня; я взял ягод, выжал их в чашу фараонову и подал чашу в руку фараону.
GEN|40|12|И сказал ему Иосиф: вот истолкование его: три ветви – это три дня;
GEN|40|13|через три дня фараон вознесет главу твою и возвратит тебя на место твое, и ты подашь чашу фараонову в руку его, по прежнему обыкновению, когда ты был у него виночерпием;
GEN|40|14|вспомни же меня, когда хорошо тебе будет, и сделай мне благодеяние, и упомяни обо мне фараону, и выведи меня из этого дома,
GEN|40|15|ибо я украден из земли Евреев; а также и здесь ничего не сделал, за что бы бросить меня в темницу.
GEN|40|16|Главный хлебодар увидел, что истолковал он хорошо, и сказал Иосифу: мне также снилось: вот на голове у меня три корзины решетчатых;
GEN|40|17|в верхней корзине всякая пища фараонова, изделие пекаря, и птицы клевали ее из корзины на голове моей.
GEN|40|18|И отвечал Иосиф и сказал: вот истолкование его: три корзины – это три дня;
GEN|40|19|через три дня фараон снимет с тебя голову твою и повесит тебя на дереве, и птицы будут клевать плоть твою с тебя.
GEN|40|20|На третий день, день рождения фараонова, сделал он пир для всех слуг своих и вспомнил о главном виночерпии и главном хлебодаре среди слуг своих;
GEN|40|21|и возвратил главного виночерпия на прежнее место, и он подал чашу в руку фараону,
GEN|40|22|а главного хлебодара повесил, как истолковал им Иосиф.
GEN|40|23|И не вспомнил главный виночерпий об Иосифе, но забыл его.
GEN|41|1|По прошествии двух лет фараону снилось: вот, он стоит у реки;
GEN|41|2|и вот, вышли из реки семь коров, хороших видом и тучных плотью, и паслись в тростнике;
GEN|41|3|но вот, после них вышли из реки семь коров других, худых видом и тощих плотью, и стали подле тех коров, на берегу реки;
GEN|41|4|и съели коровы худые видом и тощие плотью семь коров хороших видом и тучных. И проснулся фараон,
GEN|41|5|и заснул опять, и снилось ему в другой раз: вот, на одном стебле поднялось семь колосьев тучных и хороших;
GEN|41|6|но вот, после них выросло семь колосьев тощих и иссушенных восточным ветром;
GEN|41|7|и пожрали тощие колосья семь колосьев тучных и полных. И проснулся фараон и [понял, что] это сон.
GEN|41|8|Утром смутился дух его, и послал он, и призвал всех волхвов Египта и всех мудрецов его, и рассказал им фараон сон свой; но не было никого, кто бы истолковал его фараону.
GEN|41|9|И стал говорить главный виночерпий фараону и сказал: грехи мои вспоминаю я ныне;
GEN|41|10|фараон прогневался на рабов своих и отдал меня и главного хлебодара под стражу в дом начальника телохранителей;
GEN|41|11|и снился нам сон в одну ночь, мне и ему, каждому снился сон особенного значения;
GEN|41|12|там же был с нами молодой Еврей, раб начальника телохранителей; мы рассказали ему сны наши, и он истолковал нам каждому соответственно с его сновидением;
GEN|41|13|и как он истолковал нам, так и сбылось: я возвращен на место мое, а тот повешен.
GEN|41|14|И послал фараон и позвал Иосифа. И поспешно вывели его из темницы. Он остригся и переменил одежду свою и пришел к фараону.
GEN|41|15|Фараон сказал Иосифу: мне снился сон, и нет никого, кто бы истолковал его, а о тебе я слышал, что ты умеешь толковать сны.
GEN|41|16|И отвечал Иосиф фараону, говоря: это не мое; Бог даст ответ во благо фараону.
GEN|41|17|И сказал фараон Иосифу: мне снилось: вот, стою я на берегу реки;
GEN|41|18|и вот, вышли из реки семь коров тучных плотью и хороших видом и паслись в тростнике;
GEN|41|19|но вот, после них вышли семь коров других, худых, очень дурных видом и тощих плотью: я не видывал во всей земле Египетской таких худых, как они;
GEN|41|20|и съели тощие и худые коровы прежних семь коров тучных;
GEN|41|21|и вошли [тучные] в утробу их, но не приметно было, что они вошли в утробу их: они были так же худы видом, как и сначала. И я проснулся.
GEN|41|22|[Потом] снилось мне: вот, на одном стебле поднялись семь колосьев полных и хороших;
GEN|41|23|но вот, после них выросло семь колосьев тонких, тощих и иссушенных восточным ветром;
GEN|41|24|и пожрали тощие колосья семь колосьев хороших. Я рассказал это волхвам, но никто не изъяснил мне.
GEN|41|25|И сказал Иосиф фараону: сон фараонов один: что Бог сделает, то Он возвестил фараону.
GEN|41|26|Семь коров хороших, это семь лет; и семь колосьев хороших, это семь лет: сон один;
GEN|41|27|и семь коров тощих и худых, вышедших после тех, это семь лет, также и семь колосьев тощих и иссушенных восточным ветром, это семь лет голода.
GEN|41|28|Вот почему сказал я фараону: что Бог сделает, то Он показал фараону.
GEN|41|29|Вот, наступает семь лет великого изобилия во всей земле Египетской;
GEN|41|30|после них настанут семь лет голода, и забудется все то изобилие в земле Египетской, и истощит голод землю,
GEN|41|31|и неприметно будет прежнее изобилие на земле, по причине голода, который последует, ибо он будет очень тяжел.
GEN|41|32|А что сон повторился фараону дважды, [это значит], что сие истинно слово Божие, и что вскоре Бог исполнит сие.
GEN|41|33|И ныне да усмотрит фараон мужа разумного и мудрого и да поставит его над землею Египетскою.
GEN|41|34|Да повелит фараон поставить над землею надзирателей и собирать в семь лет изобилия пятую часть с земли Египетской;
GEN|41|35|пусть они берут всякий хлеб этих наступающих хороших годов и соберут в городах хлеб под ведение фараона в пищу, и пусть берегут;
GEN|41|36|и будет сия пища в запас для земли на семь лет голода, которые будут в земле Египетской, дабы земля не погибла от голода.
GEN|41|37|Сие понравилось фараону и всем слугам его.
GEN|41|38|И сказал фараон слугам своим: найдем ли мы такого, как он, человека, в котором был бы Дух Божий?
GEN|41|39|И сказал фараон Иосифу: так как Бог открыл тебе все сие, то нет столь разумного и мудрого, как ты;
GEN|41|40|ты будешь над домом моим, и твоего слова держаться будет весь народ мой; только престолом я буду больше тебя.
GEN|41|41|И сказал фараон Иосифу: вот, я поставляю тебя над всею землею Египетскою.
GEN|41|42|И снял фараон перстень свой с руки своей и надел его на руку Иосифа; одел его в виссонные одежды, возложил золотую цепь на шею ему;
GEN|41|43|велел везти его на второй из своих колесниц и провозглашать пред ним: преклоняйтесь! И поставил его над всею землею Египетскою.
GEN|41|44|И сказал фараон Иосифу: я фараон; без тебя никто не двинет ни руки своей, ни ноги своей во всей земле Египетской.
GEN|41|45|И нарек фараон Иосифу имя: Цафнаф–панеах, и дал ему в жену Асенефу, дочь Потифера, жреца Илиопольского. И пошел Иосиф по земле Египетской.
GEN|41|46|Иосифу было тридцать лет от рождения, когда он предстал пред лице фараона, царя Египетского. И вышел Иосиф от лица фараонова и прошел по всей земле Египетской.
GEN|41|47|Земля же в семь лет изобилия приносила [из зерна] по горсти.
GEN|41|48|И собрал он всякий хлеб семи лет, которые были [плодородны] в земле Египетской, и положил хлеб в городах; в [каждом] городе положил хлеб полей, окружающих его.
GEN|41|49|И скопил Иосиф хлеба весьма много, как песку морского, так что перестал и считать, ибо не стало счета.
GEN|41|50|До наступления годов голода, у Иосифа родились два сына, которых родила ему Асенефа, дочь Потифера, жреца Илиопольского.
GEN|41|51|И нарек Иосиф имя первенцу: Манассия, потому что [говорил он] Бог дал мне забыть все несчастья мои и весь дом отца моего.
GEN|41|52|А другому нарек имя: Ефрем, потому что [говорил он] Бог сделал меня плодовитым в земле страдания моего.
GEN|41|53|И прошли семь лет изобилия, которое было в земле Египетской,
GEN|41|54|и наступили семь лет голода, как сказал Иосиф. И был голод во всех землях, а во всей земле Египетской был хлеб.
GEN|41|55|Но когда и вся земля Египетская начала терпеть голод, то народ начал вопиять к фараону о хлебе. И сказал фараон всем Египтянам: пойдите к Иосифу и делайте, что он вам скажет.
GEN|41|56|И был голод по всей земле; и отворил Иосиф все житницы, и стал продавать хлеб Египтянам. Голод же усиливался в земле Египетской.
GEN|41|57|И из всех стран приходили в Египет покупать хлеб у Иосифа, ибо голод усилился по всей земле.
GEN|42|1|И узнал Иаков, что в Египте есть хлеб, и сказал Иаков сыновьям своим: что вы смотрите?
GEN|42|2|И сказал: вот, я слышал, что есть хлеб в Египте; пойдите туда и купите нам оттуда хлеба, чтобы нам жить и не умереть.
GEN|42|3|Десять братьев Иосифовых пошли купить хлеба в Египте,
GEN|42|4|а Вениамина, брата Иосифова, не послал Иаков с братьями его, ибо сказал: не случилось бы с ним беды.
GEN|42|5|И пришли сыны Израилевы покупать хлеб, вместе с другими пришедшими, ибо в земле Ханаанской был голод.
GEN|42|6|Иосиф же был начальником в земле той; он и продавал хлеб всему народу земли. Братья Иосифа пришли и поклонились ему лицем до земли.
GEN|42|7|И увидел Иосиф братьев своих и узнал их; но показал, будто не знает их, и говорил с ними сурово и сказал им: откуда вы пришли? Они сказали: из земли Ханаанской, купить пищи.
GEN|42|8|Иосиф узнал братьев своих, но они не узнали его.
GEN|42|9|И вспомнил Иосиф сны, которые снились ему о них; и сказал им: вы соглядатаи, вы пришли высмотреть наготу земли сей.
GEN|42|10|Они сказали ему: нет, господин наш; рабы твои пришли купить пищи;
GEN|42|11|мы все дети одного человека; мы люди честные; рабы твои не бывали соглядатаями.
GEN|42|12|Он сказал им: нет, вы пришли высмотреть наготу земли сей.
GEN|42|13|Они сказали: нас, рабов твоих, двенадцать братьев; мы сыновья одного человека в земле Ханаанской, и вот, меньший теперь с отцом нашим, а одного не стало.
GEN|42|14|И сказал им Иосиф: это самое я и говорил вам, сказав: вы соглядатаи;
GEN|42|15|вот как вы будете испытаны: [клянусь] жизнью фараона, вы не выйдете отсюда, если не придет сюда меньший брат ваш;
GEN|42|16|пошлите одного из вас, и пусть он приведет брата вашего, а вы будете задержаны; и откроется, правда ли у вас; и если нет, [то клянусь] жизнью фараона, что вы соглядатаи.
GEN|42|17|И отдал их под стражу на три дня.
GEN|42|18|И сказал им Иосиф в третий день: вот что сделайте, и останетесь живы, ибо я боюсь Бога:
GEN|42|19|если вы люди честные, то один брат из вас пусть содержится в доме, где вы заключены; а вы пойдите, отвезите хлеб, ради голода семейств ваших;
GEN|42|20|брата же вашего меньшого приведите ко мне, чтобы оправдались слова ваши и чтобы не умереть вам. Так они и сделали.
GEN|42|21|И говорили они друг другу: точно мы наказываемся за грех против брата нашего; мы видели страдание души его, когда он умолял нас, но не послушали; за то и постигло нас горе сие.
GEN|42|22|Рувим отвечал им и сказал: не говорил ли я вам: не грешите против отрока? но вы не послушались; вот, кровь его взыскивается.
GEN|42|23|А того не знали они, что Иосиф понимает; ибо между ними был переводчик.
GEN|42|24|И отошел от них, и заплакал. И возвратился к ним, и говорил с ними, и, взяв из них Симеона, связал его пред глазами их.
GEN|42|25|И приказал Иосиф наполнить мешки их хлебом, а серебро их возвратить каждому в мешок его, и дать им запасов на дорогу. Так и сделано с ними.
GEN|42|26|Они положили хлеб свой на ослов своих, и пошли оттуда.
GEN|42|27|И открыл один [из них] мешок свой, чтобы дать корму ослу своему на ночлеге, и увидел серебро свое в отверстии мешка его,
GEN|42|28|и сказал своим братьям: серебро мое возвращено; вот оно в мешке у меня. И смутилось сердце их, и они с трепетом друг другу говорили: что это Бог сделал с нами?
GEN|42|29|И пришли к Иакову, отцу своему, в землю Ханаанскую и рассказали ему все случившееся с ними, говоря:
GEN|42|30|начальствующий над тою землею говорил с нами сурово и принял нас за соглядатаев земли той.
GEN|42|31|И сказали мы ему: мы люди честные; мы не бывали соглядатаями;
GEN|42|32|нас двенадцать братьев, сыновей у отца нашего; одного не стало, а меньший теперь с отцом нашим в земле Ханаанской.
GEN|42|33|И сказал нам начальствующий над тою землею: вот как узнаю я, честные ли вы люди: оставьте у меня одного брата из вас, а вы возьмите хлеб ради голода семейств ваших и пойдите,
GEN|42|34|и приведите ко мне меньшого брата вашего; и узнаю я, что вы не соглядатаи, но люди честные; отдам вам брата вашего, и вы можете промышлять в этой земле.
GEN|42|35|Когда же они опорожняли мешки свои, вот, у каждого узел серебра его в мешке его. И увидели они узлы серебра своего, они и отец их, и испугались.
GEN|42|36|И сказал им Иаков, отец их: вы лишили меня детей: Иосифа нет, и Симеона нет, и Вениамина взять хотите, – все это на меня!
GEN|42|37|И сказал Рувим отцу своему, говоря: убей двух моих сыновей, если я не приведу его к тебе; отдай его на мои руки; я возвращу его тебе.
GEN|42|38|Он сказал: не пойдет сын мой с вами; потому что брат его умер, и он один остался; если случится с ним несчастье на пути, в который вы пойдете, то сведете вы седину мою с печалью во гроб.
GEN|43|1|Голод усилился на земле.
GEN|43|2|И когда они съели хлеб, который привезли из Египта, тогда отец их сказал им: пойдите опять, купите нам немного пищи.
GEN|43|3|И сказал ему Иуда, говоря: тот человек решительно объявил нам, сказав: не являйтесь ко мне на лице, если брата вашего не будет с вами.
GEN|43|4|Если пошлешь с нами брата нашего, то пойдем и купим тебе пищи,
GEN|43|5|а если не пошлешь, то не пойдем, ибо тот человек сказал нам: не являйтесь ко мне на лице, если брата вашего не будет с вами.
GEN|43|6|Израиль сказал: для чего вы сделали мне такое зло, сказав тому человеку, что у вас есть еще брат?
GEN|43|7|Они сказали: расспрашивал тот человек о нас и о родстве нашем, говоря: жив ли еще отец ваш? есть ли у вас брат? Мы и рассказали ему по этим расспросам. Могли ли мы знать, что он скажет: приведите брата вашего?
GEN|43|8|Иуда же сказал Израилю, отцу своему: отпусти отрока со мною, и мы встанем и пойдем, и живы будем и не умрем и мы, и ты, и дети наши;
GEN|43|9|я отвечаю за него, из моих рук потребуешь его; если я не приведу его к тебе и не поставлю его пред лицем твоим, то останусь я виновным пред тобою во все дни жизни;
GEN|43|10|если бы мы не медлили, то уже сходили бы два раза.
GEN|43|11|Израиль, отец их, сказал им: если так, то вот что сделайте: возьмите с собою плодов земли сей и отнесите в дар тому человеку несколько бальзама и несколько меду, стираксы и ладану, фисташков и миндальных орехов;
GEN|43|12|возьмите и другое серебро в руки ваши; а серебро, обратно положенное в отверстие мешков ваших, возвратите руками вашими: может быть, это недосмотр;
GEN|43|13|и брата вашего возьмите и, встав, пойдите опять к человеку тому;
GEN|43|14|Бог же Всемогущий да даст вам найти милость у человека того, чтобы он отпустил вам и другого брата вашего и Вениамина, а мне если уже быть бездетным, то пусть буду бездетным.
GEN|43|15|И взяли те люди дары эти, и серебра вдвое взяли в руки свои, и Вениамина, и встали, пошли в Египет и предстали пред лице Иосифа.
GEN|43|16|Иосиф, увидев между ними Вениамина, сказал начальнику дома своего: введи сих людей в дом и заколи что–нибудь из скота, и приготовь, потому что со мною будут есть эти люди в полдень.
GEN|43|17|И сделал человек тот, как сказал Иосиф, и ввел человек тот людей сих в дом Иосифов.
GEN|43|18|И испугались люди эти, что ввели их в дом Иосифов, и сказали: это за серебро, возвращенное прежде в мешки наши, ввели нас, чтобы придраться к нам и напасть на нас, и взять нас в рабство, и ослов наших.
GEN|43|19|И подошли они к начальнику дома Иосифова, и стали говорить ему у дверей дома,
GEN|43|20|и сказали: послушай, господин наш, мы приходили уже прежде покупать пищи,
GEN|43|21|и случилось, что, когда пришли мы на ночлег и открыли мешки наши, – вот серебро каждого в отверстии мешка его, серебро наше по весу его, и мы возвращаем его своими руками;
GEN|43|22|а для покупки пищи мы принесли другое серебро в руках наших, мы не знаем, кто положил серебро наше в мешки наши.
GEN|43|23|Он сказал: будьте спокойны, не бойтесь; Бог ваш и Бог отца вашего дал вам клад в мешках ваших; серебро ваше дошло до меня. И привел к ним Симеона.
GEN|43|24|И ввел тот человек людей сих в дом Иосифов и дал воды, и они омыли ноги свои; и дал корму ослам их.
GEN|43|25|И они приготовили дары к приходу Иосифа в полдень, ибо слышали, что там будут есть хлеб.
GEN|43|26|И пришел Иосиф домой; и они принесли ему в дом дары, которые были на руках их, и поклонились ему до земли.
GEN|43|27|Он спросил их о здоровье и сказал: здоров ли отец ваш старец, о котором вы говорили? жив ли еще он?
GEN|43|28|Они сказали: здоров раб твой, отец наш; еще жив. И преклонились они и поклонились.
GEN|43|29|И поднял глаза свои, и увидел Вениамина, брата своего, сына матери своей, и сказал: это брат ваш меньший, о котором вы сказывали мне? И сказал: да будет милость Божия с тобою, сын мой!
GEN|43|30|И поспешно удалился Иосиф, потому что воскипела любовь к брату его, и он готов был заплакать, и вошел он во внутреннюю комнату и плакал там.
GEN|43|31|И умыв лице свое, вышел, и скрепился и сказал: подавайте кушанье.
GEN|43|32|И подали ему особо, и им особо, и Египтянам, обедавшим с ним, особо, ибо Египтяне не могут есть с Евреями, потому что это мерзость для Египтян.
GEN|43|33|И сели они пред ним, первородный по первородству его, и младший по молодости его, и дивились эти люди друг пред другом.
GEN|43|34|И посылались им кушанья от него, и доля Вениамина была впятеро больше долей каждого из них. И пили, и довольно пили они с ним.
GEN|44|1|И приказал [Иосиф] начальнику дома своего, говоря: наполни мешки этих людей пищею, сколько они могут нести, и серебро каждого положи в отверстие мешка его,
GEN|44|2|а чашу мою, чашу серебряную, положи в отверстие мешка к младшему вместе с серебром за купленный им хлеб. И сделал тот по слову Иосифа, которое сказал он.
GEN|44|3|Утром, когда рассвело, эти люди были отпущены, они и ослы их.
GEN|44|4|Еще не далеко отошли они от города, как Иосиф сказал начальнику дома своего: ступай, догоняй этих людей и, когда догонишь, скажи им: для чего вы заплатили злом за добро?
GEN|44|5|Не та ли это, из которой пьет господин мой и он гадает на ней? Худо это вы сделали.
GEN|44|6|Он догнал их и сказал им эти слова.
GEN|44|7|Они сказали ему: для чего господин наш говорит такие слова? Нет, рабы твои не сделают такого дела.
GEN|44|8|Вот, серебро, найденное нами в отверстии мешков наших, мы обратно принесли тебе из земли Ханаанской: как же нам украсть из дома господина твоего серебро или золото?
GEN|44|9|У кого из рабов твоих найдется, тому смерть, и мы будем рабами господину нашему.
GEN|44|10|Он сказал: хорошо; как вы сказали, так пусть и будет: у кого найдется [чаша], тот будет мне рабом, а вы будете не виноваты.
GEN|44|11|Они поспешно спустили каждый свой мешок на землю и открыли каждый свой мешок.
GEN|44|12|Он обыскал, начал со старшего и окончил младшим; и нашлась чаша в мешке Вениаминовом.
GEN|44|13|И разодрали они одежды свои, и, возложив каждый на осла своего ношу, возвратились в город.
GEN|44|14|И пришли Иуда и братья его в дом Иосифа, который был еще дома, и пали пред ним на землю.
GEN|44|15|Иосиф сказал им: что это вы сделали? разве вы не знали, что такой человек, как я, конечно угадает?
GEN|44|16|Иуда сказал: что нам сказать господину нашему? что говорить? чем оправдываться? Бог нашел неправду рабов твоих; вот, мы рабы господину нашему, и мы, и тот, в чьих руках нашлась чаша.
GEN|44|17|Но [Иосиф] сказал: нет, я этого не сделаю; тот, в чьих руках нашлась чаша, будет мне рабом, а вы пойдите с миром к отцу вашему.
GEN|44|18|И подошел Иуда к нему и сказал: господин мой, позволь рабу твоему сказать слово в уши господина моего, и не прогневайся на раба твоего, ибо ты то же, что фараон.
GEN|44|19|Господин мой спрашивал рабов своих, говоря: есть ли у вас отец или брат?
GEN|44|20|Мы сказали господину нашему, что у нас есть отец престарелый, и младший сын, сын старости, которого брат умер, а он остался один [от] матери своей, и отец любит его.
GEN|44|21|Ты же сказал рабам твоим: приведите его ко мне, чтобы мне взглянуть на него.
GEN|44|22|Мы сказали господину нашему: отрок не может оставить отца своего, и если он оставит отца своего, то сей умрет.
GEN|44|23|Но ты сказал рабам твоим: если не придет с вами меньший брат ваш, то вы более не являйтесь ко мне на лице.
GEN|44|24|Когда мы пришли к рабу твоему, отцу нашему, то пересказали ему слова господина моего.
GEN|44|25|И сказал отец наш: пойдите опять, купите нам немного пищи.
GEN|44|26|Мы сказали: нельзя нам идти; а если будет с нами меньший брат наш, то пойдем; потому что нельзя нам видеть лица того человека, если не будет с нами меньшого брата нашего.
GEN|44|27|И сказал нам раб твой, отец наш: вы знаете, что жена моя родила мне двух [сынов];
GEN|44|28|один пошел от меня, и я сказал: верно он растерзан; и я не видал его доныне;
GEN|44|29|если и сего возьмете от глаз моих, и случится с ним несчастье, то сведете вы седину мою с горестью во гроб.
GEN|44|30|Теперь если я приду к рабу твоему, отцу нашему, и не будет с нами отрока, с душею которого связана душа его,
GEN|44|31|то он, увидев, что нет отрока, умрет; и сведут рабы твои седину раба твоего, отца нашего, с печалью во гроб.
GEN|44|32|Притом я, раб твой, взялся отвечать за отрока отцу моему, сказав: если не приведу его к тебе, то останусь я виновным пред отцом моим во все дни жизни.
GEN|44|33|Итак пусть я, раб твой, вместо отрока останусь рабом у господина моего, а отрок пусть идет с братьями своими:
GEN|44|34|ибо как пойду я к отцу моему, когда отрока не будет со мною? я увидел бы бедствие, которое постигло бы отца моего.
GEN|45|1|Иосиф не мог более удерживаться при всех стоявших около него и закричал: удалите от меня всех. И не оставалось при Иосифе никого, когда он открылся братьям своим.
GEN|45|2|И громко зарыдал он, и услышали Египтяне, и услышал дом фараонов.
GEN|45|3|И сказал Иосиф братьям своим: я – Иосиф, жив ли еще отец мой? Но братья его не могли отвечать ему, потому что они смутились пред ним.
GEN|45|4|И сказал Иосиф братьям своим: подойдите ко мне. Они подошли. Он сказал: я – Иосиф, брат ваш, которого вы продали в Египет;
GEN|45|5|но теперь не печальтесь и не жалейте о том, что вы продали меня сюда, потому что Бог послал меня перед вами для сохранения вашей жизни;
GEN|45|6|ибо теперь два года голода на земле: еще пять лет, в которые ни орать, ни жать не будут;
GEN|45|7|Бог послал меня перед вами, чтобы оставить вас на земле и сохранить вашу жизнь великим избавлением.
GEN|45|8|Итак не вы послали меня сюда, но Бог, Который и поставил меня отцом фараону и господином во всем доме его и владыкою во всей земле Египетской.
GEN|45|9|Идите скорее к отцу моему и скажите ему: так говорит сын твой Иосиф: Бог поставил меня господином над всем Египтом; приди ко мне, не медли;
GEN|45|10|ты будешь жить в земле Гесем; и будешь близ меня, ты, и сыны твои, и сыны сынов твоих, и мелкий и крупный скот твой, и все твое;
GEN|45|11|и прокормлю тебя там, ибо голод будет еще пять лет, чтобы не обнищал ты и дом твой и все твое.
GEN|45|12|И вот, очи ваши и очи брата моего Вениамина видят, что это мои уста говорят с вами;
GEN|45|13|скажите же отцу моему о всей славе моей в Египте и о всем, что вы видели, и приведите скорее отца моего сюда.
GEN|45|14|И пал он на шею Вениамину, брату своему, и плакал; и Вениамин плакал на шее его.
GEN|45|15|И целовал всех братьев своих и плакал, обнимая их. Потом говорили с ним братья его.
GEN|45|16|Дошел в дом фараона слух, что пришли братья Иосифа; и приятно было фараону и рабам его.
GEN|45|17|И сказал фараон Иосифу: скажи братьям твоим: вот что сделайте: навьючьте скот ваш, и ступайте в землю Ханаанскую;
GEN|45|18|и возьмите отца вашего и семейства ваши и придите ко мне; я дам вам лучшее в земле Египетской, и вы будете есть тук земли.
GEN|45|19|Тебе же повелеваю сказать им: сделайте сие: возьмите себе из земли Египетской колесниц для детей ваших и для жен ваших, и привезите отца вашего и придите;
GEN|45|20|и не жалейте вещей ваших, ибо лучшее из всей земли Египетской [дам] вам.
GEN|45|21|Так и сделали сыны Израилевы. И дал им Иосиф колесницы по приказанию фараона, и дал им путевой запас,
GEN|45|22|каждому из них он дал перемену одежд, а Вениамину дал триста сребренников и пять перемен одежд;
GEN|45|23|также и отцу своему послал десять ослов, навьюченных лучшими [произведениями] Египетскими, и десять ослиц, навьюченных зерном, хлебом и припасами отцу своему на путь.
GEN|45|24|И отпустил братьев своих, и они пошли. И сказал им: не ссорьтесь на дороге.
GEN|45|25|И пошли они из Египта, и пришли в землю Ханаанскую к Иакову, отцу своему,
GEN|45|26|и известили его, сказав: Иосиф жив, и теперь владычествует над всею землею Египетскою. Но сердце его смутилось, ибо он не верил им.
GEN|45|27|Когда же они пересказали ему все слова Иосифа, которые он говорил им, и когда увидел колесницы, которые прислал Иосиф, чтобы везти его, тогда ожил дух Иакова, отца их,
GEN|45|28|и сказал Израиль: довольно, еще жив сын мой Иосиф; пойду и увижу его, пока не умру.
GEN|46|1|И отправился Израиль со всем, что у него было, и пришел в Вирсавию, и принес жертвы Богу отца своего Исаака.
GEN|46|2|И сказал Бог Израилю в видении ночном: Иаков! Иаков! Он сказал: вот я.
GEN|46|3|[Бог] сказал: Я Бог, Бог отца твоего; не бойся идти в Египет, ибо там произведу от тебя народ великий;
GEN|46|4|Я пойду с тобою в Египет, Я и выведу тебя обратно. Иосиф своею рукою закроет глаза [твои].
GEN|46|5|Иаков отправился из Вирсавии; и повезли сыны Израилевы Иакова отца своего, и детей своих, и жен своих на колесницах, которые послал фараон, чтобы привезти его.
GEN|46|6|И взяли они скот свой и имущество свое, которое приобрели в земле Ханаанской, и пришли в Египет, – Иаков и весь род его с ним.
GEN|46|7|Сынов своих и внуков своих с собою, дочерей своих и внучек своих и весь род свой привел он с собою в Египет.
GEN|46|8|Вот имена сынов Израилевых, пришедших в Египет: Иаков и сыновья его. Первенец Иакова Рувим.
GEN|46|9|Сыны Рувима: Ханох и Фаллу, Хецрон и Харми.
GEN|46|10|Сыны Симеона: Иемуил и Иамин, и Огад, и Иахин, и Цохар, и Саул, сын Хананеянки.
GEN|46|11|Сыны Левия: Гирсон, Кааф и Мерари.
GEN|46|12|Сыны Иуды: Ир и Онан, и Шела, и Фарес, и Зара; но Ир и Онан умерли в земле Ханаанской. Сыны Фареса были: Есром и Хамул.
GEN|46|13|Сыны Иссахара: Фола и Фува, Иов и Шимрон.
GEN|46|14|Сыны Завулона: Серед и Елон, и Иахлеил.
GEN|46|15|Это сыны Лии, которых она родила Иакову в Месопотамии, и Дину, дочь его. Всех душ сынов его и дочерей его – тридцать три.
GEN|46|16|Сыны Гада: Цифион и Хагги, Шуни и Эцбон, Ери и Ароди и Арели.
GEN|46|17|Сыны Асира: Имна и Ишва, и Ишви, и Бриа, и Серах, сестра их. Сыны Брии: Хевер и Малхиил.
GEN|46|18|Это сыны Зелфы, которую Лаван дал Лии, дочери своей; она родила их Иакову шестнадцать душ.
GEN|46|19|Сыны Рахили, жены Иакова: Иосиф и Вениамин.
GEN|46|20|И родились у Иосифа в земле Египетской Манассия и Ефрем, которых родила ему Асенефа, дочь Потифера, жреца Илиопольского.
GEN|46|21|Сыны Вениамина: Бела и Бехер и Ашбел; Гера и Нааман, Эхи и Рош, Муппим и Хуппим и Ард.
GEN|46|22|Это сыны Рахили, которые родились у Иакова, всего четырнадцать душ.
GEN|46|23|Сын Дана: Хушим.
GEN|46|24|Сыны Неффалима: Иахцеил и Гуни, и Иецер, и Шиллем.
GEN|46|25|Это сыны Валлы, которую дал Лаван дочери своей Рахили; она родила их Иакову всего семь душ.
GEN|46|26|Всех душ, пришедших с Иаковом в Египет, которые произошли из чресл его, кроме жен сынов Иаковлевых, всего шестьдесят шесть душ.
GEN|46|27|Сынов Иосифа, которые родились у него в Египте, две души. Всех душ дома Иаковлева, перешедших в Египет, семьдесят.
GEN|46|28|Иуду послал он пред собою к Иосифу, чтобы он указал [путь] в Гесем. И пришли в землю Гесем.
GEN|46|29|Иосиф запряг колесницу свою и выехал навстречу Израилю, отцу своему, в Гесем, и, увидев его, пал на шею его, и долго плакал на шее его.
GEN|46|30|И сказал Израиль Иосифу: умру я теперь, увидев лице твое, ибо ты еще жив.
GEN|46|31|И сказал Иосиф братьям своим и дому отца своего: я пойду, извещу фараона и скажу ему: братья мои и дом отца моего, которые были в земле Ханаанской, пришли ко мне;
GEN|46|32|эти люди пастухи овец, ибо скотоводы они; и мелкий и крупный скот свой, и все, что у них, привели они.
GEN|46|33|Если фараон призовет вас и скажет: какое занятие ваше?
GEN|46|34|то вы скажите: [мы], рабы твои, скотоводами были от юности нашей доныне, и мы и отцы наши, чтобы вас поселили в земле Гесем. Ибо мерзость для Египтян всякий пастух овец.
GEN|47|1|И пришел Иосиф и известил фараона и сказал: отец мой и братья мои, с мелким и крупным скотом своим и со всем, что у них, пришли из земли Ханаанской; и вот, они в земле Гесем.
GEN|47|2|И из братьев своих он взял пять человек и представил их фараону.
GEN|47|3|И сказал фараон братьям его: какое ваше занятие? Они сказали фараону: пастухи овец рабы твои, и мы и отцы наши.
GEN|47|4|И сказали они фараону: мы пришли пожить в этой земле, потому что нет пажити для скота рабов твоих, ибо в земле Ханаанской сильный голод; итак позволь поселиться рабам твоим в земле Гесем.
GEN|47|5|И сказал фараон Иосифу: отец твой и братья твои пришли к тебе;
GEN|47|6|земля Египетская пред тобою; на лучшем месте земли посели отца твоего и братьев твоих; пусть живут они в земле Гесем; и если знаешь, что между ними есть способные люди, поставь их смотрителями над моим скотом.
GEN|47|7|И привел Иосиф Иакова, отца своего, и представил его фараону; и благословил Иаков фараона.
GEN|47|8|Фараон сказал Иакову: сколько лет жизни твоей?
GEN|47|9|Иаков сказал фараону: дней странствования моего сто тридцать лет; малы и несчастны дни жизни моей и не достигли до лет жизни отцов моих во днях странствования их.
GEN|47|10|И благословил фараона Иаков и вышел от фараона.
GEN|47|11|И поселил Иосиф отца своего и братьев своих, и дал им владение в земле Египетской, в лучшей части земли, в земле Раамсес, как повелел фараон.
GEN|47|12|И снабжал Иосиф отца своего и братьев своих и весь дом отца своего хлебом, по потребностям каждого семейства.
GEN|47|13|И не было хлеба по всей земле, потому что голод весьма усилился, и изнурены были от голода земля Египетская и земля Ханаанская.
GEN|47|14|Иосиф собрал все серебро, какое было в земле Египетской и в земле Ханаанской, за хлеб, который покупали, и внес Иосиф серебро в дом фараонов.
GEN|47|15|И серебро истощилось в земле Египетской и в земле Ханаанской. Все Египтяне пришли к Иосифу и говорили: дай нам хлеба; зачем нам умирать пред тобою, потому что серебро вышло у нас?
GEN|47|16|Иосиф сказал: пригоняйте скот ваш, и я буду давать вам за скот ваш, если серебро вышло у вас.
GEN|47|17|И пригоняли они к Иосифу скот свой; и давал им Иосиф хлеб за лошадей, и за стада мелкого скота, и за стада крупного скота, и за ослов; и снабжал их хлебом в тот год за весь скот их.
GEN|47|18|И прошел этот год; и пришли к нему на другой год и сказали ему: не скроем от господина нашего, что серебро истощилось и стада скота нашего у господина нашего; ничего не осталось у нас пред господином нашим, кроме тел наших и земель наших;
GEN|47|19|для чего нам погибать в глазах твоих, и нам и землям нашим? купи нас и земли наши за хлеб, и мы с землями нашими будем рабами фараону, а ты дай нам семян, чтобы нам быть живыми и не умереть, и чтобы не опустела земля.
GEN|47|20|И купил Иосиф всю землю Египетскую для фараона, потому что продали Египтяне каждый свое поле, ибо голод одолевал их. И досталась земля фараону.
GEN|47|21|И народ сделал он рабами от одного конца Египта до другого.
GEN|47|22|Только земли жрецов не купил, ибо жрецам от фараона положен был участок, и они питались своим участком, который дал им фараон; посему и не продали земли своей.
GEN|47|23|И сказал Иосиф народу: вот, я купил теперь для фараона вас и землю вашу; вот вам семена, и засевайте землю;
GEN|47|24|когда будет жатва, давайте пятую часть фараону, а четыре части останутся вам на засеяние полей, на пропитание вам и тем, кто в домах ваших, и на пропитание детям вашим.
GEN|47|25|Они сказали: ты спас нам жизнь; да обретем милость в очах господина нашего и да будем рабами фараону.
GEN|47|26|И поставил Иосиф в закон земле Египетской, даже до сего дня: пятую часть давать фараону, исключая только землю жрецов, которая не принадлежала фараону.
GEN|47|27|И жил Израиль в земле Египетской, в земле Гесем, и владели они ею, и плодились, и весьма умножились.
GEN|47|28|И жил Иаков в земле Египетской семнадцать лет; и было дней Иакова, годов жизни его, сто сорок семь лет.
GEN|47|29|И пришло время Израилю умереть, и призвал он сына своего Иосифа и сказал ему: если я нашел благоволение в очах твоих, положи руку твою под стегно мое и [клянись], что ты окажешь мне милость и правду, не похоронишь меня в Египте,
GEN|47|30|дабы мне лечь с отцами моими; вынесешь меня из Египта и похоронишь меня в их гробнице. [Иосиф] сказал: сделаю по слову твоему.
GEN|47|31|И сказал: клянись мне. И клялся ему. И поклонился Израиль на возглавие постели.
GEN|48|1|После того Иосифу сказали: вот, отец твой болен. И он взял с собою двух сынов своих, Манассию и Ефрема.
GEN|48|2|Иакова известили и сказали: вот, сын твой Иосиф идет к тебе. Израиль собрал силы свои и сел на постели.
GEN|48|3|И сказал Иаков Иосифу: Бог Всемогущий явился мне в Лузе, в земле Ханаанской, и благословил меня,
GEN|48|4|и сказал мне: вот, Я распложу тебя, и размножу тебя, и произведу от тебя множество народов, и дам землю сию потомству твоему после тебя, в вечное владение.
GEN|48|5|И ныне два сына твои, родившиеся тебе в земле Египетской, до моего прибытия к тебе в Египет, мои они; Ефрем и Манассия, как Рувим и Симеон, будут мои;
GEN|48|6|дети же твои, которые родятся от тебя после них, будут твои; они под именем братьев своих будут именоваться в их уделе.
GEN|48|7|Когда я шел из Месопотамии, умерла у меня Рахиль в земле Ханаанской, по дороге, не доходя несколько до Ефрафы, и я похоронил ее там на дороге к Ефрафе, что [ныне] Вифлеем.
GEN|48|8|И увидел Израиль сыновей Иосифа и сказал: кто это?
GEN|48|9|И сказал Иосиф отцу своему: это сыновья мои, которых Бог дал мне здесь. Иаков сказал: подведи их ко мне, и я благословлю их.
GEN|48|10|Глаза же Израилевы притупились от старости; не мог он видеть [ясно. Иосиф] подвел их к нему, и он поцеловал их и обнял их.
GEN|48|11|И сказал Израиль Иосифу: не надеялся я видеть твое лице; но вот, Бог показал мне и детей твоих.
GEN|48|12|И отвел их Иосиф от колен его и поклонился ему лицем своим до земли.
GEN|48|13|И взял Иосиф обоих, Ефрема в правую свою руку против левой Израиля, а Манассию в левую против правой Израиля, и подвел к нему.
GEN|48|14|Но Израиль простер правую руку свою и положил на голову Ефрему, хотя сей был меньший, а левую на голову Манассии. С намерением положил он так руки свои, хотя Манассия был первенец.
GEN|48|15|И благословил Иосифа и сказал: Бог, пред Которым ходили отцы мои Авраам и Исаак, Бог, пасущий меня с тех пор, как я существую, до сего дня,
GEN|48|16|Ангел, избавляющий меня от всякого зла, да благословит отроков сих; да будет на них наречено имя мое и имя отцов моих Авраама и Исаака, и да возрастут они во множество посреди земли.
GEN|48|17|И увидел Иосиф, что отец его положил правую руку свою на голову Ефрема; и прискорбно было ему это. И взял он руку отца своего, чтобы переложить ее с головы Ефрема на голову Манассии,
GEN|48|18|и сказал Иосиф отцу своему: не так, отец мой, ибо это – первенец; положи на его голову правую руку твою.
GEN|48|19|Но отец его не согласился и сказал: знаю, сын мой, знаю; и от него произойдет народ, и он будет велик; но меньший его брат будет больше его, и от семени его произойдет многочисленный народ.
GEN|48|20|И благословил их в тот день, говоря: тобою будет благословлять Израиль, говоря: Бог да сотворит тебе, как Ефрему и Манассии. И поставил Ефрема выше Манассии.
GEN|48|21|И сказал Израиль Иосифу: вот, я умираю; и Бог будет с вами и возвратит вас в землю отцов ваших;
GEN|48|22|я даю тебе, преимущественно пред братьями твоими, один участок, который я взял из рук Аморреев мечом моим и луком моим.
GEN|49|1|И призвал Иаков сыновей своих и сказал: соберитесь, и я возвещу вам, что будет с вами в грядущие дни;
GEN|49|2|сойдитесь и послушайте, сыны Иакова, послушайте Израиля, отца вашего.
GEN|49|3|Рувим, первенец мой! ты – крепость моя и начаток силы моей, верх достоинства и верх могущества;
GEN|49|4|но ты бушевал, как вода, – не будешь преимуществовать, ибо ты взошел на ложе отца твоего, ты осквернил постель мою, взошел.
GEN|49|5|Симеон и Левий братья, орудия жестокости мечи их;
GEN|49|6|в совет их да не внидет душа моя, и к собранию их да не приобщится слава моя, ибо они во гневе своем убили мужа и по прихоти своей перерезали жилы тельца;
GEN|49|7|проклят гнев их, ибо жесток, и ярость их, ибо свирепа; разделю их в Иакове и рассею их в Израиле.
GEN|49|8|Иуда! тебя восхвалят братья твои. Рука твоя на хребте врагов твоих; поклонятся тебе сыны отца твоего.
GEN|49|9|Молодой лев Иуда, с добычи, сын мой, поднимается. Преклонился он, лег, как лев и как львица: кто поднимет его?
GEN|49|10|Не отойдет скипетр от Иуды и законодатель от чресл его, доколе не приидет Примиритель, и Ему покорность народов.
GEN|49|11|Он привязывает к виноградной лозе осленка своего и к лозе лучшего винограда сына ослицы своей; моет в вине одежду свою и в крови гроздов одеяние свое;
GEN|49|12|блестящи очи [его] от вина, и белы зубы от молока.
GEN|49|13|Завулон при береге морском будет жить и у пристани корабельной, и предел его до Сидона.
GEN|49|14|Иссахар осел крепкий, лежащий между протоками вод;
GEN|49|15|и увидел он, что покой хорош, и что земля приятна: и преклонил плечи свои для ношения бремени и стал работать в уплату дани.
GEN|49|16|Дан будет судить народ свой, как одно из колен Израиля;
GEN|49|17|Дан будет змеем на дороге, аспидом на пути, уязвляющим ногу коня, так что всадник его упадет назад.
GEN|49|18|На помощь твою надеюсь, Господи!
GEN|49|19|Гад, – толпа будет теснить его, но он оттеснит ее по пятам.
GEN|49|20|Для Асира – слишком тучен хлеб его, и он будет доставлять царские яства.
GEN|49|21|Неффалим – теревинф рослый, распускающий прекрасные ветви.
GEN|49|22|Иосиф – отрасль плодоносного [дерева], отрасль плодоносного [дерева] над источником; ветви его простираются над стеною;
GEN|49|23|огорчали его, и стреляли и враждовали на него стрельцы,
GEN|49|24|но тверд остался лук его, и крепки мышцы рук его, от рук мощного [Бога] Иаковлева. Оттуда Пастырь и твердыня Израилева,
GEN|49|25|от Бога отца твоего, [Который] и да поможет тебе, и от Всемогущего, Который и да благословит тебя благословениями небесными свыше, благословениями бездны, лежащей долу, благословениями сосцов и утробы,
GEN|49|26|благословениями отца твоего, которые превышают благословения гор древних и приятности холмов вечных; да будут они на голове Иосифа и на темени избранного между братьями своими.
GEN|49|27|Вениамин, хищный волк, утром будет есть ловитву и вечером будет делить добычу.
GEN|49|28|Вот все двенадцать колен Израилевых; и вот что сказал им отец их; и благословил их, и дал им благословение, каждому свое.
GEN|49|29|И заповедал он им и сказал им: я прилагаюсь к народу моему; похороните меня с отцами моими в пещере, которая на поле Ефрона Хеттеянина,
GEN|49|30|в пещере, которая на поле Махпела, что пред Мамре, в земле Ханаанской, которую купил Авраам с полем у Ефрона Хеттеянина в собственность для погребения;
GEN|49|31|там похоронили Авраама и Сарру, жену его; там похоронили Исаака и Ревекку, жену его; и там похоронил я Лию;
GEN|49|32|это поле и пещера, которая на нем, куплена у сынов Хеттеевых.
GEN|49|33|И окончил Иаков завещание сыновьям своим, и положил ноги свои на постель, и скончался, и приложился к народу своему.
GEN|50|1|Иосиф пал на лице отца своего, и плакал над ним, и целовал его.
GEN|50|2|И повелел Иосиф слугам своим – врачам, бальзамировать отца его; и врачи набальзамировали Израиля.
GEN|50|3|И исполнилось ему сорок дней, ибо столько дней употребляется на бальзамирование, и оплакивали его Египтяне семьдесят дней.
GEN|50|4|Когда же прошли дни плача по нем, Иосиф сказал придворным фараона, говоря: если я обрел благоволение в очах ваших, то скажите фараону так:
GEN|50|5|отец мой заклял меня, сказав: вот, я умираю; во гробе моем, который я выкопал себе в земле Ханаанской, там похорони меня. И теперь хотел бы я пойти и похоронить отца моего и возвратиться.
GEN|50|6|И сказал фараон: пойди и похорони отца твоего, как он заклял тебя.
GEN|50|7|И пошел Иосиф хоронить отца своего. И пошли с ним все слуги фараона, старейшины дома его и все старейшины земли Египетской,
GEN|50|8|и весь дом Иосифа, и братья его, и дом отца его. Только детей своих и мелкий и крупный скот свой оставили в земле Гесем.
GEN|50|9|С ним отправились также колесницы и всадники, так что сонм был весьма велик.
GEN|50|10|И дошли они до Горен–гаатада при Иордане и плакали там плачем великим и весьма сильным; и сделал [Иосиф] плач по отце своем семь дней.
GEN|50|11|И видели жители земли той, Хананеи, плач в Горен–гаатаде, и сказали: велик плач этот у Египтян! Посему наречено имя [месту] тому: плач Египтян, что при Иордане.
GEN|50|12|И сделали сыновья [Иакова] с ним, как он заповедал им;
GEN|50|13|и отнесли его сыновья его в землю Ханаанскую и похоронили его в пещере на поле Махпела, которую купил Авраам с полем в собственность для погребения у Ефрона Хеттеянина, пред Мамре.
GEN|50|14|И возвратился Иосиф в Египет, сам и братья его и все ходившие с ним хоронить отца его, после погребения им отца своего.
GEN|50|15|И увидели братья Иосифовы, что умер отец их, и сказали: что, если Иосиф возненавидит нас и захочет отмстить нам за все зло, которое мы ему сделали?
GEN|50|16|И послали они сказать Иосифу: отец твой пред смертью своею завещал, говоря:
GEN|50|17|так скажите Иосифу: прости братьям твоим вину и грех их, так как они сделали тебе зло. И ныне прости вины рабов Бога отца твоего. Иосиф плакал, когда ему говорили это.
GEN|50|18|Пришли и сами братья его, и пали пред лицем его, и сказали: вот, мы рабы тебе.
GEN|50|19|И сказал Иосиф: не бойтесь, ибо я боюсь Бога;
GEN|50|20|вот, вы умышляли против меня зло; но Бог обратил это в добро, чтобы сделать то, что теперь есть: сохранить жизнь великому числу людей;
GEN|50|21|итак не бойтесь: я буду питать вас и детей ваших. И успокоил их и говорил по сердцу их.
GEN|50|22|И жил Иосиф в Египте сам и дом отца его; жил же Иосиф всего сто десять лет.
GEN|50|23|И видел Иосиф детей у Ефрема до третьего рода, также и сыновья Махира, сына Манассиина, родились на колени Иосифа.
GEN|50|24|И сказал Иосиф братьям своим: я умираю, но Бог посетит вас и выведет вас из земли сей в землю, о которой клялся Аврааму, Исааку и Иакову.
GEN|50|25|И заклял Иосиф сынов Израилевых, говоря: Бог посетит вас, и вынесите кости мои отсюда.
GEN|50|26|И умер Иосиф ста десяти лет. И набальзамировали его и положили в ковчег в Египте.
