SONG|1|1|所罗门 的雅歌 。
SONG|1|2|愿他用口与我亲吻。 你的爱情比酒更美，
SONG|1|3|你的膏油馨香， 你的名如倾泻而出的香膏， 所以童女都爱你。
SONG|1|4|愿你吸引我跟随你；让我们快跑吧！ 王领我进入他的内室。 我们必因你欢喜快乐， 我们要思念你的爱情， 胜似思念美酒。 她们爱你是理所当然的。
SONG|1|5|耶路撒冷 的女子啊， 我虽然黑，却是秀美， 如同 基达 的帐棚， 好像 所罗门 的幔子，
SONG|1|6|不要因太阳把我晒黑了就瞪着我。 我母亲的儿子向我发怒， 他们使我看守葡萄园； 我自己的葡萄园我却没有看守。
SONG|1|7|我心所爱的啊，请告诉我， 你在何处牧羊？ 正午在何处使羊歇卧？ 我何必像蒙着脸的女子 在你同伴的羊群旁边呢？
SONG|1|8|你这女子中最美丽的， 你若不知道， 只管跟随羊群的脚踪行， 在牧人的帐棚边，牧放你的小山羊。
SONG|1|9|我的佳偶， 你好比法老战车上的骏马。
SONG|1|10|你的两颊因发辫而秀美， 你的颈项因珠串而华丽。
SONG|1|11|我们要为你编上金链，镶上银饰。
SONG|1|12|王正坐席的时候， 我的哪哒香膏散发香味。
SONG|1|13|我的良人好像一袋没药， 在我胸怀中。
SONG|1|14|我的良人好像一束凤仙花， 在 隐．基底 的葡萄园中。
SONG|1|15|看哪，我的佳偶，你真美丽！ 看哪，你真美丽！你的眼睛是鸽子。
SONG|1|16|看哪，我的良人，你多英俊可爱！ 让我们以青草为床榻，
SONG|1|17|以香柏树为房子的栋梁， 以松树作屋顶的椽木。
SONG|2|1|我是 沙仑 的玫瑰花， 是谷中的百合花。
SONG|2|2|我的佳偶在女子中， 好像荆棘里的百合花。
SONG|2|3|我的良人在男子中， 如同苹果树在树林里。 我欢欢喜喜坐在他的荫下， 尝他果子的滋味，觉得甘甜。
SONG|2|4|他领我进入宴会厅， 为我插上爱的旗帜。
SONG|2|5|请你们用葡萄饼增补我力， 以苹果畅快我的心， 因我为爱而生病。
SONG|2|6|他的左手在我头下， 他的右手将我环抱。
SONG|2|7|耶路撒冷 的女子啊， 我指着羚羊或田野的母鹿嘱咐你们， 不要唤醒，不要挑动爱情，等它自发。
SONG|2|8|听啊！我良人的声音， 看哪！他穿山越岭而来。
SONG|2|9|我的良人像羚羊，像小鹿。 看哪，他站在我们的墙壁边， 从窗户往里观看， 从窗格子往里窥探。
SONG|2|10|我的良人对我说： “我的佳偶，起来！ 我的美人，与我同去！
SONG|2|11|看哪，因为冬天已逝， 雨水止住，已经过去了。
SONG|2|12|地上百花开放， 歌唱的时候到了， 斑鸠的声音在我们境内也听见了。
SONG|2|13|无花果树的果子渐渐成熟， 葡萄树开花，散发香气。 我的佳偶，起来！ 我的美人，与我同去！
SONG|2|14|我的鸽子啊，你在磐石穴中， 在陡岩的隐密处。 求你容我得见你的面貌， 求你容我得听你的声音； 因你的声音悦耳， 你的容貌秀美。
SONG|2|15|请为我们擒拿狐狸， 就是毁坏葡萄园的小狐狸， 我们的葡萄正在开花。”
SONG|2|16|我的良人属我，我也属他， 他在百合花中放牧。
SONG|2|17|我的良人哪， 等到天起凉风、 日影飞去的时候， 愿你归回，像羚羊， 像小鹿，在崎岖的山 上。
SONG|3|1|我夜间躺卧在床上， 寻找我心所爱的； 我寻找他，却寻不着。
SONG|3|2|“我要起来，绕行城中， 在街市上，在广场上， 寻找我心所爱的。” 我寻找他，却寻不着。
SONG|3|3|城中巡逻的守卫遇见我， “你们看见我心所爱的没有？”
SONG|3|4|我刚离开他们，就遇见我心所爱的。 我拉住他，不放他走， 领他进入我母亲的家， 到怀我者的内室。
SONG|3|5|耶路撒冷 的女子啊， 我指着羚羊或田野的母鹿嘱咐你们， 不要唤醒，不要挑动爱情，等它自发。
SONG|3|6|那如烟柱从旷野上来， 薰了没药、乳香，扑上商人各样香粉的是谁呢？
SONG|3|7|看哪，是 所罗门 的轿， 周围有六十个勇士， 都是 以色列 中的勇士。
SONG|3|8|他们的手都持刀，善于争战， 各人腰间佩刀，防备夜间恐怖的攻击。
SONG|3|9|所罗门 王用 黎巴嫩 木 为自己制作轿子。
SONG|3|10|轿柱是用银做的， 轿底是用金做的， 坐垫是紫色的， 其中所铺的是 耶路撒冷 女子的爱情。
SONG|3|11|锡安的女子啊， 你们要出去观看 所罗门 王！ 他头戴冠冕，就是在他结婚当天 心中喜乐的时候，他母亲给他戴上的。
SONG|4|1|看哪，我的佳偶，你真美丽！看哪，你真美丽！ 你的眼睛在面纱后好像鸽子。 你的头发如同一群山羊，从 基列山 下来。
SONG|4|2|你的牙齿如新剪毛的一群母羊，洗净之后走上来， 它们成对，没有一颗是单独的。
SONG|4|3|你的唇好像一条朱红线， 你的嘴秀美。 你的鬓角在面纱后， 如同迸开的石榴。
SONG|4|4|你的颈项犹如 大卫 为收藏军器而造的高塔， 其上悬挂一千个盾牌， 都是勇士的盾牌。
SONG|4|5|你的两乳好像百合花中吃草的一对小鹿， 是母鹿双生的。
SONG|4|6|我要往没药山和乳香冈去， 直到天起凉风、 日影飞去的时候。
SONG|4|7|我的佳偶，你全然美丽， 毫无瑕疵！
SONG|4|8|我的新娘，请你与我一同离开 黎巴嫩 ， 与我一同离开 黎巴嫩 。 从 亚玛拿 山巅， 从 示尼珥 ，就是 黑门山 顶， 从狮子的洞， 从豹子的山往下观看。
SONG|4|9|我的妹子，我的新娘， 你夺了我的心。 你明眸一瞥， 你颈项的链子， 夺了我的心！
SONG|4|10|我的妹子，我的新娘， 你的爱情 何其美！ 你的爱情比酒甜美！ 你膏油的馨香胜过一切香料！
SONG|4|11|我的新娘，你的唇滴下蜂蜜， 你的舌下有蜜，有奶。 你衣服的香气宛如 黎巴嫩 的芬芳。
SONG|4|12|我的妹子，我的新娘 是上锁的园子， 是禁闭的园子 ， 是封闭的泉源。
SONG|4|13|你园内所种的结了石榴， 有佳美的果子， 并凤仙花与哪哒树。
SONG|4|14|有哪哒和番红花， 香菖蒲和桂树， 并各样乳香木、没药、沉香， 与一切上等的香料。
SONG|4|15|你是园中的泉，活水的井， 是从 黎巴嫩 涌流而下的溪水。
SONG|4|16|北风啊，兴起！ 南风啊，吹来！ 吹在我的园内， 使其中的香气散发出来。 愿我的良人进入自己园里， 吃他佳美的果子。
SONG|5|1|我的妹子，我的新娘， 我进入我的园中， 采了我的没药和香料， 吃了我的蜂房和蜂蜜， 喝了我的酒和奶。 我的朋友，请吃！ 我亲爱的，请喝，多多地喝！
SONG|5|2|我身躺卧，我心却醒。 这是我良人的声音； 他敲门： “我的妹子，我的佳偶， 我的鸽子，我完美的人儿， 请你为我开门； 因我的头沾满露水， 我的发被夜露滴湿。”
SONG|5|3|我脱了衣裳，怎能再穿上呢？ 我洗了脚，怎可再弄脏呢？
SONG|5|4|我的良人从门缝里伸进他的手， 我便因他动了心。
SONG|5|5|我起来，要为我的良人开门。 我的两手滴下没药， 我的指头有没药汁滴在门闩上。
SONG|5|6|我为我的良人开了门， 我的良人却已转身走了。 他说话的时候，我魂不守舍。 我寻找他，竟寻不着， 我呼叫他，他却不回答。
SONG|5|7|城中巡逻的守卫遇见我， 打了我，伤了我， 看守城墙的人夺去我的披肩。
SONG|5|8|耶路撒冷 的女子啊，我嘱咐你们： 若遇见我的良人， 要告诉他，我为爱而生病。
SONG|5|9|你这女子中最美丽的， 你的良人有什么胜过别的良人呢？ 你的良人有什么胜过别的良人， 使你这样嘱咐我们？
SONG|5|10|我的良人红润发亮， 超乎万人之上。
SONG|5|11|他的头像千足的纯金， 他的发绺卷曲，黑如乌鸦。
SONG|5|12|他的眼如溪水旁的鸽子， 沐浴在奶中，安得合式 。
SONG|5|13|他的两颊如香花园， 如香草台 ； 他的嘴唇像百合花， 滴下没药汁。
SONG|5|14|他的双手宛如金条， 镶嵌水苍玉； 他的身体如同雕刻的象牙， 周围镶嵌蓝宝石。
SONG|5|15|他的腿好比白玉石柱， 安在精金座上； 他的容貌如 黎巴嫩 ， 佳美如香柏树。
SONG|5|16|他的口甘甜， 他全然可爱。 耶路撒冷 的女子啊， 这是我的良人， 这是我的朋友。
SONG|6|1|你这女子中最美丽的， 你的良人往何处去？ 你的良人转向何处去了？ 我们好与你同去寻找他。
SONG|6|2|我的良人进入自己园中， 到香花园， 在园内放牧， 采百合花。
SONG|6|3|我属我的良人， 我的良人属我； 他在百合花中放牧。
SONG|6|4|我的佳偶啊，你美丽如 得撒 ， 秀美如 耶路撒冷 ， 威武如展开旌旗的军队。
SONG|6|5|求你转开眼睛不要看我， 因你的眼睛使我慌乱。 你的头发如同一群山羊，从 基列山 下来。
SONG|6|6|你的牙齿如一群母羊，洗净之后走上来， 它们成对，没有一颗是单独的。
SONG|6|7|你的鬓角在面纱后， 如同迸开的石榴。
SONG|6|8|虽有六十王后、八十妃嫔， 并有无数的童女。
SONG|6|9|她是我独一的鸽子、我完美的人儿， 是她母亲独生的， 是生养她的所宠爱的。 女子见了都称她有福， 王后妃嫔见了也赞美她。
SONG|6|10|那俯视如晨曦、 美丽如月亮、皎洁如太阳、 威武如展开旌旗军队的是谁呢？
SONG|6|11|我下到坚果园， 要看谷中青翠的植物， 要看葡萄可曾发芽， 石榴可曾放蕊；
SONG|6|12|不知不觉， 我仿佛坐在我百姓高官 的战车中。
SONG|6|13|回来，回来， 书拉密 的女子； 回来，回来，我们要看你。 你们为何要观看 书拉密 的女子， 像观看两队人马在跳舞 呢？
SONG|7|1|尊贵的女子啊，你的脚在鞋中何等秀美！ 你的大腿圆润，好像美玉， 是巧匠的手做成的。
SONG|7|2|你的肚脐如圆杯， 不缺调和的酒。 你的肚子如一堆麦子， 周围有百合花。
SONG|7|3|你的两乳好像一对小鹿， 是母鹿双生的。
SONG|7|4|你的颈项如象牙塔， 你的眼睛像 希实本 、 巴特．拉并 门旁的水池， 你的鼻子仿佛朝向 大马士革 的 黎巴嫩 塔。
SONG|7|5|你的头在你身上好像 迦密山 ， 你头上的发呈紫色， 王被这发绺系住了。
SONG|7|6|我亲爱的，喜乐的女子啊， 你何等美丽！何等令人喜悦！
SONG|7|7|你的身材好像棕树， 你的两乳如同累累的果实。
SONG|7|8|我说：我要爬上棕树，抓住枝子。 愿你的两乳好像葡萄累累， 愿你鼻子的香气如苹果；
SONG|7|9|你的上颚如美酒， 直流入我良人的口里， 流入沉睡者的口中 。
SONG|7|10|我属我的良人， 他也恋慕我。
SONG|7|11|来吧！我的良人， 让我们往田间去， 在村庄住宿。
SONG|7|12|早晨让我们起来往葡萄园去， 看葡萄树发芽没有， 花开了没有， 石榴放蕊没有， 在那里我要将我的爱情给你。
SONG|7|13|曼陀罗草 散发香味， 在我们的门内有各样新陈佳美的果子； 我的良人，这都是我为你保存的。
SONG|8|1|惟愿你像我的兄弟， 像吃我母亲奶的兄弟。 我在外头遇见你就与你亲吻， 谁也不轻看我。
SONG|8|2|我必引导你， 领你进入我母亲的家， 她必教导我， 我必使你喝石榴汁酿的香酒。
SONG|8|3|他的左手在我头下， 他的右手将我环抱。
SONG|8|4|耶路撒冷 的女子啊， 我嘱咐你们， 不要唤醒、不要挑动爱情，等它自发。
SONG|8|5|那靠着良人从旷野上来的是谁呢？ 在苹果树下，我叫醒了你； 在那里，你母亲曾为了生你而阵痛， 在那里，生你的为你阵痛。
SONG|8|6|求你将我放在你心上如印记， 带在你臂上如戳记。 因为爱情如死之坚强， 热恋如阴间之牢固， 所发的光是火焰的光， 是极其猛烈的火焰 。
SONG|8|7|爱情，众水不能熄灭， 江河也不能淹没。 若有人拿家中所有的财宝要换爱情， 就全被藐视。
SONG|8|8|我们有一小妹， 她还没有乳房， 人来提亲的日子， 我们当为她怎么办呢？
SONG|8|9|她若是墙， 我们要在其上建造银塔； 她若是门， 我们要用香柏木板围护她。
SONG|8|10|我是墙， 我的两乳像塔。 那时，我在他眼中是找到平安的人。
SONG|8|11|所罗门 在 巴力．哈们 有一葡萄园， 他将这葡萄园租给看守的人， 每人为其中的果子要交一千银子。
SONG|8|12|我有属自己的葡萄园。 所罗门 哪，一千归你， 两百归看守果子的人。
SONG|8|13|你这住在园中的， 同伴都要听你的声音， 求你使我也得以听见。
SONG|8|14|我的良人哪，求你快来！ 像羚羊，像小鹿，在香草山上。
