3JOHN|1|1|我作長老的寫信給親愛的 該猶 ，就是我真心所愛的。
3JOHN|1|2|親愛的，我願你事事安寧，身體健康，正如你的心神安寧一樣。
3JOHN|1|3|我非常歡喜，有弟兄到這裏來，證實你對真理的忠誠，就是你按著真理而行。
3JOHN|1|4|我聽見我的兒女按真理而行，我的歡喜沒有比這個更大的。
3JOHN|1|5|親愛的，你對弟兄，特別是對作客旅的弟兄所做的都是忠誠的。
3JOHN|1|6|他們在教會面前證實了你的愛；你若以對得起上帝的方式，為他們送行就好了；
3JOHN|1|7|因為他們是為基督的名 出外，並沒有從未信的人接受甚麼。
3JOHN|1|8|所以，我們應當接待這樣的人，好讓我們與他們在真理上成為同工。
3JOHN|1|9|我曾寫過一些東西給教會，但他們中間那好作領袖的 丟特腓 不接納我們。
3JOHN|1|10|為此，我若去，要提起他所做的事，就是他用惡言攻擊我們，還不滿足，他自己不接納弟兄，有人願意接納，他還阻止，並且把接納弟兄的人趕出教會。
3JOHN|1|11|親愛的，不要效法惡，只要效法善。行善的人屬乎上帝；行惡的人未曾見過上帝。
3JOHN|1|12|低米丟 行善，有眾人給他作見證，又有真理給他作見證，就是我們也給他作見證，你知道我們的見證是真的。
3JOHN|1|13|我還有許多事要寫給你，卻不願意用筆墨來寫給你，
3JOHN|1|14|但盼望很快見到你，我們好面對面談論。
3JOHN|1|15|願你平安！朋友們都向你問安。請你替我按著名字一一向朋友們問安。
