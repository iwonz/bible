AMOS|1|1|verba Amos qui fuit in pastoralibus de Thecuae quae vidit super Israhel in diebus Oziae regis Iuda et in diebus Hieroboam filii Ioas regis Israhel ante duos annos terraemotus
AMOS|1|2|et dixit Dominus de Sion rugiet et de Hierusalem dabit vocem suam et luxerunt speciosa pastorum et exsiccatus est vertex Carmeli
AMOS|1|3|haec dicit Dominus super tribus sceleribus Damasci et super quattuor non convertam eum eo quod trituraverint in plaustris ferreis Galaad
AMOS|1|4|et mittam ignem in domum Azahel et devorabit domos Benadad
AMOS|1|5|et conteram vectem Damasci et disperdam habitatorem de campo Idoli et tenentem sceptrum de domo Voluptatis et transferetur populus Syriae Cyrenen dicit Dominus
AMOS|1|6|haec dicit Dominus super tribus sceleribus Gazae et super quattuor non convertam eum eo quod transtulerit captivitatem perfectam ut concluderet eam in Idumea
AMOS|1|7|et mittam ignem in murum Gazae et devorabit aedes eius
AMOS|1|8|et disperdam habitatorem de Azoto et tenentem sceptrum de Ascalone et convertam manum meam super Accaron et peribunt reliqui Philisthinorum dicit Dominus Deus
AMOS|1|9|haec dicit Dominus super tribus sceleribus Tyri et super quattuor non convertam eum eo quod concluserint captivitatem perfectam in Idumea et non sint recordati foederis fratrum
AMOS|1|10|et emittam ignem in murum Tyri et devorabit aedes eius
AMOS|1|11|haec dicit Dominus super tribus sceleribus Edom et super quattuor non convertam eum eo quod persecutus sit in gladio fratrem suum et violaverit misericordiam eius et tenuerit ultra furorem suum et indignationem suam servaverit usque in finem
AMOS|1|12|mittam ignem in Theman et devorabit aedes Bosrae
AMOS|1|13|haec dicit Dominus super tribus sceleribus filiorum Ammon et super quattuor non convertam eum eo quod dissecuerit praegnantes Galaad ad dilatandum terminum suum
AMOS|1|14|et succendam ignem in muro Rabbae et devorabit aedes eius in ululatu in die belli et in turbine in die commotionis
AMOS|1|15|et ibit Melchom in captivitatem ipse et principes eius simul dicit Dominus
AMOS|2|1|haec dicit Dominus super tribus sceleribus Moab et super quattuor non convertam eum eo quod incenderit ossa regis Idumeae usque ad cinerem
AMOS|2|2|et mittam ignem in Moab et devorabit aedes Carioth et morietur in sonitu Moab in clangore tubae
AMOS|2|3|et disperdam iudicem de medio eius et omnes principes eius interficiam cum eo dicit Dominus
AMOS|2|4|haec dicit Dominus super tribus sceleribus Iuda et super quattuor non convertam eum eo quod abiecerint legem Domini et mandata eius non custodierint deceperunt enim eos idola sua post quae abierant patres eorum
AMOS|2|5|et mittam ignem in Iuda et devorabit aedes Hierusalem
AMOS|2|6|haec dicit Dominus super tribus sceleribus Israhel et super quattuor non convertam eum pro eo quod vendiderit argento iustum et pauperem pro calciamentis
AMOS|2|7|qui conterunt super pulverem terrae capita pauperum et viam humilium declinant et filius ac pater eius ierunt ad puellam ut violarent nomen sanctum meum
AMOS|2|8|et super vestimentis pigneratis accubuerunt iuxta omne altare et vinum damnatorum bibebant in domo Dei sui
AMOS|2|9|ego autem exterminavi Amorreum a facie eorum cuius altitudo cedrorum altitudo eius et fortis ipse quasi quercus et contrivi fructum eius desuper et radices eius subter
AMOS|2|10|ego sum qui ascendere vos feci de terra Aegypti et eduxi vos in deserto quadraginta annis ut possideretis terram Amorrei
AMOS|2|11|et suscitavi de filiis vestris in prophetas et de iuvenibus vestris nazarenos numquid non ita est filii Israhel dicit Dominus
AMOS|2|12|et propinabatis nazarenis vino et prophetis mandabatis dicentes ne prophetetis
AMOS|2|13|ecce ego stridebo super vos sicut stridet plaustrum onustum faeno
AMOS|2|14|et peribit fuga a veloce et fortis non obtinebit virtutem suam et robustus non salvabit animam suam
AMOS|2|15|et tenens arcum non stabit et velox pedibus suis non salvabitur et ascensor equi non salvabit animam suam
AMOS|2|16|et robustus corde inter fortes nudus fugiet in die illa dicit Dominus
AMOS|3|1|audite verbum quod locutus est Dominus super vos filii Israhel super omni cognatione quam eduxi de terra Aegypti dicens
AMOS|3|2|tantummodo vos cognovi ex omnibus cognationibus terrae idcirco visitabo super vos omnes iniquitates vestras
AMOS|3|3|numquid ambulabunt duo pariter nisi convenerit eis
AMOS|3|4|numquid rugiet leo in saltu nisi habuerit praedam numquid dabit catulus leonis vocem de cubili suo nisi aliquid adprehenderit
AMOS|3|5|numquid cadet avis in laqueum terrae absque aucupe numquid auferetur laqueus de terra antequam quid ceperit
AMOS|3|6|si clanget tuba in civitate et populus non expavescet si erit malum in civitate quod Dominus non fecit
AMOS|3|7|quia non faciet Dominus Deus verbum nisi revelaverit secretum suum ad servos suos prophetas
AMOS|3|8|leo rugiet quis non timebit Dominus Deus locutus est quis non prophetabit
AMOS|3|9|auditum facite in aedibus Azoti et in aedibus terrae Aegypti et dicite congregamini super montes Samariae et videte insanias multas in medio eius et calumniam patientes in penetrabilibus eius
AMOS|3|10|et nescierunt facere rectum dicit Dominus thesaurizantes iniquitatem et rapinas in aedibus suis
AMOS|3|11|propterea haec dicit Dominus Deus tribulabitur et circumietur terra et detrahetur ex te fortitudo tua et diripientur aedes tuae
AMOS|3|12|haec dicit Dominus quomodo si eruat pastor de ore leonis duo crura aut extremum auriculae sic eruentur filii Israhel qui habitant in Samaria in plaga lectuli et in Damasco grabatti
AMOS|3|13|audite et contestamini in domo Iacob dicit Dominus Deus exercituum
AMOS|3|14|quia in die cum visitare coepero praevaricationes Israhel super eum visitabo et super altaria Bethel et amputabuntur cornua altaris et cadent in terram
AMOS|3|15|et percutiam domum hiemalem cum domo aestiva et peribunt domus eburneae et dissipabuntur aedes multae dicit Dominus
AMOS|4|1|audite verbum hoc vaccae pingues quae estis in monte Samariae quae calumniam facitis egenis et confringitis pauperes quae dicitis dominis vestris adferte et bibemus
AMOS|4|2|iuravit Dominus Deus in sancto suo quia ecce dies venient super vos et levabunt vos in contis et reliquias vestras in ollis ferventibus
AMOS|4|3|et per aperturas exibitis altera contra alteram et proiciemini in Armon dicit Dominus
AMOS|4|4|venite ad Bethel et impie agite ad Galgalam et multiplicate praevaricationem et offerte mane victimas vestras tribus diebus decimas vestras
AMOS|4|5|et sacrificate de fermentato laudem et vocate voluntarias oblationes et adnuntiate sic enim voluistis filii Israhel dicit Dominus Deus
AMOS|4|6|unde et ego dedi vobis stuporem dentium in cunctis urbibus vestris et indigentiam panum in omnibus locis vestris et non estis reversi ad me dicit Dominus
AMOS|4|7|ego quoque prohibui a vobis imbrem cum adhuc tres menses superessent usque ad messem et plui super civitatem unam et super civitatem alteram non plui pars una conpluta est et pars super quam non plui aruit
AMOS|4|8|et venerunt duae et tres civitates ad civitatem unam ut biberent aquam et non sunt satiatae et non redistis ad me dicit Dominus
AMOS|4|9|percussi vos in vento urente et in aurugine multitudinem hortorum vestrorum et vinearum vestrarum oliveta vestra et ficeta vestra comedit eruca et non redistis ad me dicit Dominus
AMOS|4|10|misi in vos mortem in via Aegypti percussi in gladio iuvenes vestros usque ad captivitatem equorum vestrorum et ascendere feci putredinem castrorum vestrorum in nares vestras et non redistis ad me dicit Dominus
AMOS|4|11|subverti vos sicut subvertit Deus Sodomam et Gomorram et facti estis quasi torris raptus de incendio et non redistis ad me dicit Dominus
AMOS|4|12|quapropter haec faciam tibi Israhel postquam autem haec fecero tibi praeparare in occursum Dei tui Israhel
AMOS|4|13|quia ecce formans montes et creans ventum et adnuntians homini eloquium suum faciens matutinam nebulam et gradiens super excelsa terrae Dominus Deus exercituum nomen eius
AMOS|5|1|audite verbum istud quod ego levo super vos planctum domus Israhel cecidit non adiciet ut resurgat
AMOS|5|2|virgo Israhel proiecta est in terram suam non est qui suscitet eam
AMOS|5|3|quia haec dicit Dominus Deus urbs de qua egrediebantur mille relinquentur in ea centum et de qua egrediebantur centum relinquentur in ea decem in domo Israhel
AMOS|5|4|quia haec dicit Dominus domui Israhel quaerite me et vivetis
AMOS|5|5|et nolite quaerere Bethel et in Galgala nolite intrare et in Bersabee non transibitis quia Galgala captiva ducetur et Bethel erit inutilis
AMOS|5|6|quaerite Dominum et vivite ne forte conburatur ut ignis domus Ioseph et devorabit et non erit qui extinguat Bethel
AMOS|5|7|qui convertitis in absinthium iudicium et iustitiam in terra relinquitis
AMOS|5|8|facientem Arcturum et Orionem et convertentem in mane tenebras et diem nocte mutantem qui vocat aquas maris et effundit eas super faciem terrae Dominus nomen eius
AMOS|5|9|qui subridet vastitatem super robustum et depopulationem super potentem adfert
AMOS|5|10|odio habuerunt in porta corripientem et loquentem perfecte abominati sunt
AMOS|5|11|idcirco pro eo quod diripiebatis pauperem et praedam electam tollebatis ab eo domos quadro lapide aedificabitis et non habitabitis in eis vineas amantissimas plantabitis et non bibetis vinum earum
AMOS|5|12|quia cognovi multa scelera vestra et fortia peccata vestra hostes iusti accipientes munus et pauperes in porta deprimentes
AMOS|5|13|ideo prudens in tempore illo tacebit quia tempus malum est
AMOS|5|14|quaerite bonum et non malum ut vivatis et erit Dominus Deus exercituum vobiscum sicut dixistis
AMOS|5|15|odite malum et diligite bonum et constituite in porta iudicium si forte misereatur Dominus Deus exercituum reliquiis Ioseph
AMOS|5|16|propterea haec dicit Dominus Deus exercituum Dominator in omnibus plateis planctus et in cunctis quae foris sunt dicetur vae vae et vocabunt agricolam ad luctum et ad planctum eos qui sciunt plangere
AMOS|5|17|et in omnibus vineis erit planctus quia pertransibo in medio tui dicit Dominus
AMOS|5|18|vae desiderantibus diem Domini ad quid eam vobis dies Domini ista tenebrae et non lux
AMOS|5|19|quomodo si fugiat vir a facie leonis et occurrat ei ursus et ingrediatur domum et innitatur manu sua super parietem et mordeat eum coluber
AMOS|5|20|numquid non tenebrae dies Domini et non lux et caligo et non splendor in ea
AMOS|5|21|odi et proieci festivitates vestras et non capiam odorem coetuum vestrorum
AMOS|5|22|quod si adtuleritis mihi holocaustomata et munera vestra non suscipiam et vota pinguium vestrorum non respiciam
AMOS|5|23|aufer a me tumultum carminum tuorum et cantica lyrae tuae non audiam
AMOS|5|24|et revelabitur quasi aqua iudicium et iustitia quasi torrens fortis
AMOS|5|25|numquid hostias et sacrificium obtulistis mihi in deserto quadraginta annis domus Israhel
AMOS|5|26|et portastis tabernaculum Moloch vestro et imaginem idolorum vestrorum sidus dei vestri quae fecistis vobis
AMOS|5|27|et migrare vos faciam trans Damascum dixit Dominus Deus exercituum nomen eius
AMOS|6|1|vae qui opulenti estis in Sion et confiditis in monte Samariae optimates capita populorum ingredientes pompatice domum Israhel
AMOS|6|2|transite in Chalanne et videte et ite inde in Emath magnam et descendite in Geth Palestinorum et ad optima quaeque regna horum si latior terminus eorum termino vestro est
AMOS|6|3|qui separati estis in diem malum et adpropinquatis solio iniquitatis
AMOS|6|4|qui dormitis in lectis eburneis et lascivitis in stratis vestris qui comeditis agnum de grege et vitulos de medio armenti
AMOS|6|5|qui canitis ad vocem psalterii sicut David putaverunt se habere vasa cantici
AMOS|6|6|bibentes in fialis vinum et optimo unguento delibuti et nihil patiebantur super contritione Ioseph
AMOS|6|7|quapropter nunc migrabunt in capite transmigrantium et auferetur factio lascivientium
AMOS|6|8|iuravit Dominus Deus in anima sua dicit Dominus Deus exercituum detestor ego superbiam Iacob et domos eius odi et tradam civitatem cum habitatoribus suis
AMOS|6|9|quod si reliqui fuerint decem viri in domo una et ipsi morientur
AMOS|6|10|et tollet eum propinquus suus et conburet eum ut efferat ossa de domo et dicet ei qui in penetrabilibus domus est numquid adhuc est apud te
AMOS|6|11|et respondebit finis est et dicet ei tace et non recorderis nominis Domini
AMOS|6|12|quia ecce Dominus mandabit et percutiet domum maiorem ruinis et domum minorem scissionibus
AMOS|6|13|numquid currere queunt in petris equi aut arari potest in bubalis quoniam convertistis in amaritudinem iudicium et fructum iustitiae in absinthium
AMOS|6|14|qui laetamini in nihili qui dicitis numquid non in fortitudine nostra adsumpsimus nobis cornua
AMOS|6|15|ecce enim suscitabo super vos domus Israhel dicit Dominus Deus exercituum gentem et conterent vos ab introitu Emath usque ad torrentem Deserti
AMOS|7|1|haec ostendit mihi Dominus Deus et ecce fictor lucustae in principio germinantium serotini imbris et ecce serotinus post tonsorem regis
AMOS|7|2|et factum est cum consummasset comedere herbam terrae et dixi Domine Deus propitius esto obsecro quis suscitabit Iacob quia parvulus est
AMOS|7|3|misertus est Dominus super hoc non erit dixit Dominus
AMOS|7|4|haec ostendit mihi Dominus Deus et ecce vocabat iudicium ad ignem Dominus Deus et devoravit abyssum multam et comedit simul partem
AMOS|7|5|et dixi Domine Deus quiesce obsecro quis suscitabit Iacob quia parvulus est
AMOS|7|6|misertus est Dominus super hoc sed et istud non erit dixit Dominus Deus
AMOS|7|7|haec ostendit mihi et ecce Dominus stans super murum litum et in manu eius trulla cementarii
AMOS|7|8|et dixit Dominus ad me quid tu vides Amos et dixi trullam cementarii et dixit Dominus ecce ego ponam trullam in medio populi mei Israhel non adiciam ultra superinducere eum
AMOS|7|9|et demolientur excelsa idoli et sanctificationes Israhel desolabuntur et consurgam super domum Hieroboam in gladio
AMOS|7|10|et misit Amasias sacerdos Bethel ad Hieroboam regem Israhel dicens rebellavit contra te Amos in medio domus Israhel non poterit terra sustinere universos sermones eius
AMOS|7|11|haec enim dicit Amos in gladio morietur Hieroboam et Israhel captivus migrabit de terra sua
AMOS|7|12|et dixit Amasias ad Amos qui vides gradere fuge in terram Iuda et comede ibi panem et ibi prophetabis
AMOS|7|13|et in Bethel non adicies ultra ut prophetes quia sanctificatio regis est et domus regni est
AMOS|7|14|et respondit Amos et dixit ad Amasiam non sum propheta et non sum filius prophetae sed armentarius ego sum vellicans sycomoros
AMOS|7|15|et tulit me Dominus cum sequerer gregem et dixit ad me Dominus vade propheta ad populum meum Israhel
AMOS|7|16|et nunc audi verbum Domini tu dicis non prophetabis super Israhel et non stillabis super domum idoli
AMOS|7|17|propter hoc haec dicit Dominus uxor tua in civitate fornicabitur et filii tui et filiae tuae in gladio cadent et humus tua funiculo metietur et tu in terra polluta morieris et Israhel captivus migrabit de terra sua
AMOS|8|1|haec ostendit mihi Dominus Deus et ecce uncinus pomorum
AMOS|8|2|et dixit quid tu vides Amos et dixi uncinum pomorum et dixit Dominus ad me venit finis super populum meum Israhel non adiciam ultra ut pertranseam eum
AMOS|8|3|et stridebunt cardines templi in die illa dicit Dominus Deus multi morientur in omni loco proicietur silentium
AMOS|8|4|audite hoc qui conteritis pauperem et deficere facitis egenos terrae
AMOS|8|5|dicentes quando transibit mensis et venundabimus merces et sabbatum et aperiemus frumentum ut inminuamus mensuram et augeamus siclum et subponamus stateras dolosas
AMOS|8|6|ut possideamus in argento egenos et pauperes pro calciamentis et quisquilias frumenti vendamus
AMOS|8|7|iuravit Dominus in superbia Iacob si oblitus fuero usque ad finem omnia opera eorum
AMOS|8|8|numquid super isto non commovebitur terra et lugebit omnis habitator eius et ascendet quasi fluvius universus et eicietur et defluet quasi rivus Aegypti
AMOS|8|9|et erit in die illa dicit Dominus occidet sol meridie et tenebrescere faciam terram in die luminis
AMOS|8|10|et convertam festivitates vestras in luctum et omnia cantica vestra in planctum et inducam super omne dorsum vestrum saccum et super omne caput calvitium et ponam eam quasi luctum unigeniti et novissima eius quasi diem amarum
AMOS|8|11|ecce dies veniunt dicit Dominus et mittam famem in terram non famem panis neque sitim aquae sed audiendi verbum Domini
AMOS|8|12|et commovebuntur a mari usque ad mare et ab aquilone usque ad orientem circumibunt quaerentes verbum Domini et non invenient
AMOS|8|13|in die illa deficient virgines pulchrae et adulescentes in siti
AMOS|8|14|qui iurant in delicto Samariae et dicunt vivit deus tuus Dan et vivit via Bersabee et cadent et non resurgent ultra
AMOS|9|1|vidi Dominum stantem super altare et dixit percute cardinem et commoveantur superliminaria avaritia enim in capite omnium et novissimum eorum in gladio interficiam non erit fuga eis fugiet et non salvabitur ex eis qui fugerit
AMOS|9|2|si descenderint usque ad infernum inde manus mea educet eos et si ascenderint usque ad caelum inde detraham eos
AMOS|9|3|et si absconditi fuerint in vertice Carmeli inde scrutans auferam eos et si celaverint se ab oculis meis in fundo maris ibi mandabo serpenti et mordebit eos
AMOS|9|4|et si abierint in captivitatem coram inimicis suis ibi mandabo gladio et occidet eos et ponam oculos meos super eos in malum et non in bonum
AMOS|9|5|et Dominus Deus exercituum qui tangit terram et tabescet et lugebunt omnes habitantes in ea et ascendet sicut rivus omnis et defluet sicut fluvius Aegypti
AMOS|9|6|qui aedificat in caelo ascensionem suam et fasciculum suum super terram fundavit qui vocat aquas maris et effundit eas super faciem terrae Dominus nomen eius
AMOS|9|7|numquid non ut filii Aethiopum vos estis mihi filii Israhel ait Dominus numquid non Israhel ascendere feci de terra Aegypti et Palestinos de Cappadocia et Syros de Cyrene
AMOS|9|8|ecce oculi Domini Dei super regnum peccans et conteram illud a facie terrae verumtamen conterens non conteram domum Iacob dicit Dominus
AMOS|9|9|ecce enim ego mandabo et concutiam in omnibus gentibus domum Israhel sicut concutitur in cribro et non cadet lapillus super terram
AMOS|9|10|in gladio morientur omnes peccatores populi mei qui dicunt non adpropinquabit et non veniet super nos malum
AMOS|9|11|in die illo suscitabo tabernaculum David quod cecidit et reaedificabo aperturas murorum eius et ea quae corruerant instaurabo et reaedificabo eum sicut diebus antiquis
AMOS|9|12|ut possideant reliquias Idumeae et omnes nationes eo quod invocatum sit nomen meum super eos dicit Dominus faciens haec
AMOS|9|13|ecce dies veniunt dicit Dominus et conprehendet arator messorem et calcator uvae mittentem semen et stillabunt montes dulcedinem et omnes colles culti erunt
AMOS|9|14|et convertam captivitatem populi mei Israhel et aedificabunt civitates desertas et habitabunt et plantabunt vineas et bibent vinum earum et facient hortos et comedent fructus eorum
