NAH|1|1|论 尼尼微 的默示， 伊勒歌斯 人 那鸿 所见异象的书。
NAH|1|2|耶和华是忌邪 、报应的上帝。 耶和华施报应，大有愤怒； 耶和华向他的敌人报应， 向他的仇敌怀怒。
NAH|1|3|耶和华不轻易发怒，大有能力， 但耶和华万不以有罪的为无罪。 他的道路在旋风和暴风之中， 云彩为他脚下的尘土。
NAH|1|4|他斥责海，使海枯干， 使一切江河干涸。 巴珊 和 迦密 衰残， 黎巴嫩 的花草也衰残了。
NAH|1|5|大山因他震动， 小山也都融化； 大地在他面前突起， 世界和住在其间的也都如此。
NAH|1|6|他发愤恨，谁能立得住呢？ 他发烈怒，谁能当得起呢？ 他的愤怒如火倾泄而出， 磐石因他崩裂。
NAH|1|7|耶和华本为善， 在患难的日子为人的保障， 并且认识那些投靠他的人；
NAH|1|8|但他必以涨溢的洪水淹没其地方 ， 又驱逐仇敌进入黑暗。
NAH|1|9|你们筹划何种计谋攻击耶和华呢？ 他必终结一切， 仇敌 不会再度兴起。
NAH|1|10|你们像杂乱的荆棘， 像喝醉了的人， 又如枯干的碎秸，全然烧灭。
NAH|1|11|有一人从你那里出来， 图谋邪恶，设恶计攻击耶和华。
NAH|1|12|耶和华如此说： “他们虽然势力强大，人数众多， 也要被剪除，归于无有。 我虽曾使你受苦， 却不再使你受苦。
NAH|1|13|现在，我要从你身上折断他的轭， 解开捆绑你的绳索。”
NAH|1|14|耶和华已经发命令，指着你说： “你的名下必不再留后； 我要从你神明的庙中除灭雕刻的偶像和铸造的偶像， 我必因你的卑贱，为你预备坟墓。”
NAH|1|15|看哪，山上有报佳音、传平安之人的脚踪。 犹大 啊，守你的节期， 还你的愿吧！ 因为恶人不再侵犯你， 他已灭绝净尽了。
NAH|2|1|那打碎你的人 上到你面前。 要看守堡垒，把守道路， 要挺起腰来，大大使力。
NAH|2|2|耶和华复兴 雅各 的荣华， 像复兴 以色列 的荣华； 因为蹂躏者曾经蹂躏他们， 毁坏了他们的葡萄枝。
NAH|2|3|他勇士的盾牌是红的， 精兵都穿朱红衣服。 在预备打仗的日子， 战车上的铁闪烁如火 ， 柏木的枪杆也已举起 ；
NAH|2|4|战车在街上疾行， 在广场上来往奔驰， 形状如火把， 飞驰如闪电。
NAH|2|5|他 招聚他的贵族； 他们前行时绊跌， 速上城墙， 预备屏障。
NAH|2|6|河闸开放， 宫殿冲没。
NAH|2|7|这是命定之事： 王后赤身被掳 ， 宫女捶胸， 哀鸣如鸽子。
NAH|2|8|尼尼微 自古以来 如同聚水的池子； 现在居民都在逃跑 。 “站住！站住！” 却无人回转。
NAH|2|9|你们抢夺金子吧！ 你们抢夺银子吧！ 因为所积蓄的无穷， 华美的宝器无数。
NAH|2|10|荒芜，荒凉，全然荒废， 人心害怕，双膝颤抖， 腰部疼痛，脸都变色。
NAH|2|11|狮子的洞， 幼狮喂养之处在哪里呢？ 公狮、母狮、小狮出入， 无人使它们惊吓之地在哪里呢？
NAH|2|12|公狮撕碎的足够给幼狮吃， 又为母狮掐死猎物， 把猎物塞满它的洞穴， 把撕碎的装满它的窝。
NAH|2|13|看哪，我与你为敌，将它的战车 焚烧成烟，刀剑必吞灭你的少壮狮子；我必从地上除灭你的猎物，你使者的声音必不再听见。这是万军之耶和华说的。
NAH|3|1|祸哉！这流人血的城， 欺诈连连，抢夺充斥， 掳掠的事总不止息。
NAH|3|2|鞭声响亮，车轮轰轰， 马匹跳跃，战车奔腾；
NAH|3|3|骑兵争先，刀剑发光， 枪矛闪烁，被杀的甚多， 尸首成堆，尸骸无数， 人因尸骸而绊跌，
NAH|3|4|都因那美貌的妓女多有淫行， 惯行邪术， 藉淫行诱惑 列国， 用邪术诱惑万族。
NAH|3|5|看哪，我与你为敌， 掀开你的下摆，蒙在你脸上， 使列邦看见你的赤体， 使列国观看你的羞辱。 这是万军之耶和华说的。
NAH|3|6|我必将可憎污秽之物抛在你身上， 使你被藐视，为众人所观看。
NAH|3|7|凡看见你的，都必逃离你，说： “ 尼尼微 荒凉了！有谁为你悲伤呢？ 我何处找到安慰你的人呢？”
NAH|3|8|你能胜过 挪亚们 吗？ 它坐落在众河之间， 周围有水， 海 作它的城郭， 海 作它的城墙。
NAH|3|9|古实 和 埃及 是它的力量， 没有穷尽， 弗 人和 路比 人是它的帮手。
NAH|3|10|但它被流放，被人掳去， 它的婴孩也被摔碎在各街头； 人为它的贵族抽签， 它的权贵都被锁链锁住。
NAH|3|11|你也必喝醉，昏迷错乱， 并因仇敌的缘故寻求庇护。
NAH|3|12|你一切的堡垒必如无花果树上初熟的果子， 一经摇动，就落在想吃的人口中。
NAH|3|13|看哪，你中间的士兵是妇女， 你国中的关口向仇敌敞开， 你的门闩被火焚烧。
NAH|3|14|你要打水预备受困； 要加强防御， 取土踹泥， 做成砖模。
NAH|3|15|在那里，火要吞灭你， 刀必杀戮你， 如蝻子般吞灭你。 你人数增多如蝻子， 增多如蝗虫吧！
NAH|3|16|你增添商贾，多过天上的星宿； 如蝻子蜕皮飞去。
NAH|3|17|你的领袖多如蝗虫， 你的将军仿佛成群的蝗虫； 天凉时齐落在篱笆上， 太阳一出就飞去， 人不知道落在何处。
NAH|3|18|亚述 王啊， 你的牧人睡觉， 你的贵族躺卧 ， 你的百姓散在山间， 无人招聚。
NAH|3|19|你的损伤并未减轻， 你的伤痕极其重大。 凡听见这消息的人都因你拍掌。 有谁没有时常遭受你的暴行呢？
