ZECH|1|1|Восьмого місяця другого року Дарія було Господнє слово до пророка Захарія, сина Берехії, сина Іддового, таке:
ZECH|1|2|Розгнівався Господь на батьків ваших палючим гнівом.
ZECH|1|3|І скажи їм: Так говорить Господь Саваот: Верніться до Мене, говорить Господь Саваот, і вернуся до вас, говорить Господь Саваот.
ZECH|1|4|Не будьте, як ваші батьки, що до них кликали стародавні пророки, говорячи: Так говорить Господь Саваот: Верніться з доріг ваших злих і з чинів ваших лихих! Та не слухали ви й не прислухались до Мене, говорить Господь.
ZECH|1|5|Де вони, батьки ваші? А пророки чи ж навіки живуть?
ZECH|1|6|Та слова Мої й постанови Мої, що Я наказав рабам Моїм пророкам, чи ж не досягли вони до ваших батьків? І вернулись вони та й сказали: Як задумав Господь Саваот зробити нам за нашими дорогами й за нашими чинами, так зробив Він із нами.
ZECH|1|7|Двадцятого й четвертого дня, одинадцятого місяця, це місяць шеват, за другого року Дарія було слово Господнє до пророка Захарія, сина Берехії, сина Іддового, таке:
ZECH|1|8|Бачив я цієї ночі, аж ось на червоному коні їде муж, і він стоїть між миртами, що в глибині, а за ним коні червоні, руді та білі.
ZECH|1|9|І сказав я: Що це, мій пане? І відказав мені той Ангол, що говорив зо мною: Я тобі покажу, що це таке.
ZECH|1|10|І відповів той муж, що стояв між миртами, та й сказав: Це ті, що Господь їх послав обійти землю.
ZECH|1|11|І відповіли вони Господньому Анголові, що стояв між миртами, та й сказали: Перейшли ми землю, і ось уся земля сидить спокійно.
ZECH|1|12|І відповів Ангол Господній та й сказав: Господи Саваоте, аж доки Ти не змилосердишся над Єрусалимом та над Юдиними містами, на які Ти гніваєшся оце сімдесят літ?
ZECH|1|13|І відповів Господь Анголові, що говорив зо мною, слова добрі, слова втішливі.
ZECH|1|14|І сказав до мене той Ангол, що говорив зо мною: Клич, говорячи: Так говорить Господь Саваот: Піклуюся Я про Єрусалим та про Сіон великим піклуванням.
ZECH|1|15|І гнівом великим Я гніваюся на ті спокійні народи, на яких Я мало гнівався, а вони допомогли злому.
ZECH|1|16|Тому так промовляє Господь: Вернуся Я до Єрусалиму з милосердям, храм Мій буде збудований у ньому, говорить Господь Саваот, а мірничий шнур буде розтягнений над Єрусалимом.
ZECH|1|17|Ще клич та й скажи: Так говорить Господь Саваот: Знов добром переповняться міста Мої, і Господь ще потішить Сіона, і ще вибере Єрусалима!
ZECH|1|18|(2-1) І звів я очі свої, та й побачив, аж ось чотири роги.
ZECH|1|19|(2-2) І запитав я Ангола, що говорив зо мною: Що це? А він відказав мені: Це ті роги, що розпорошили Юду й Ізраїля та Єрусалим.
ZECH|1|20|(2-3) І Господь показав мені чотирьох майстрів.
ZECH|1|21|(2-4) І запитав я: Що вони приходять зробити? А Він відказав, говорячи: Це ті роги, що розпорошили Юду, так що ніхто не підвів голови. А ці прийшли настрашити їх, щоб скинути роги тих народів, що підносять рога проти Юдиного краю, щоб його розпорошити.
ZECH|2|1|(2-5) І звів Я очі свої та й побачив, аж ось муж, а в його руці мірничий шнур.
ZECH|2|2|(2-6) І сказав я: Куди ти йдеш? А він відказав мені: Щоб зміряти Єрусалим, щоб побачити, яка ширина його та яка довжина його.
ZECH|2|3|(2-7) Аж ось Ангол, що говорив зо мною, виходить, а навпроти нього виходить Ангол інший.
ZECH|2|4|(2-8) І сказав він до нього: Біжи, говори цьому юнакові, кажучи: Невкріплений буде Єрусалим через многість людей та худоби в середині його.
ZECH|2|5|(2-9) А Я стану для нього, говорить Господь, огняним муром навколо, і стану славою в середині його.
ZECH|2|6|(2-10) Горе, горе, втікайте з північного краю, говорить Господь, бо на чотири небесні вітри розпорошу Я вас, промовляє Господь.
ZECH|2|7|(2-11) Горе, втікай до Сіону, мешканко дочки Вавилону!
ZECH|2|8|(2-12) Бо так промовляє Господь Саваот: Для слави послав Він мене до народів, що вас грабували, бо хто вас доторкується, той доторкується до зірця Його ока.
ZECH|2|9|(2-13) Бо ось тільки махну Я своєю рукою на них, і для їхніх рабів вони здобиччю стануть, і пізнаєте ви, що Господь Саваот мене вислав.
ZECH|2|10|(2-14) Співай же та тішся, о дочко Сіону, бо ось Я приходжу та перебуватиму посеред тебе, говорить Господь!
ZECH|2|11|(2-15) І дня того прилучаться люди численні до Господа, і стануть народом Мені, а Я перебуватиму посеред тебе, і довідаєшся, що Господь Саваот мене вислав до тебе.
ZECH|2|12|(2-16) І Юду, спадок Свій, посяде Господь на святій землі, і вибере Єрусалима Він ще!
ZECH|2|13|(2-17) Замовчи ж, всяке тіло, перед Господнім лицем, бо Він пробудився з мешкання святого Свого!
ZECH|3|1|І показав Він мені Ісуса, великого священика, що стояв перед лицем Господнього Ангола, а сатана стояв по правиці його, щоб противитися йому.
ZECH|3|2|І сказав Господь сатані: Господь буде картати тебе, сатано, і буде картати тебе Господь, Який вибрав Собі Єрусалима! Чи ж він не головешка, що вціліла від огню?
ZECH|3|3|А Ісус одягнений був у брудну одежу, і стояв перед лицем Ангола.
ZECH|3|4|І він заговорив та й сказав до тих, що стояли перед його лицем, говорячи: Здійміть з нього цю брудну одежу! І сказав він йому: Я зняв з тебе провину твою, і зодягну тебе в шати коштовні.
ZECH|3|5|І він сказав: Нехай покладуть чистого завоя на його голову! І поклали чистого завоя на його голову, і зодягли його в шати, а Ангол Господній стояв.
ZECH|3|6|І освідчив Ангол Господній Ісусові, промовляючи:
ZECH|3|7|Так говорить Господь Саваот: Якщо ти будеш ходити Моїми дорогами, і якщо стерегтимеш сторожу Мою, тоді й ти будеш судити Мій дім, і також будеш стерегти Мої подвір'я, і дам тобі ходити поміж тими, що стоять тут.
ZECH|3|8|Послухай но, Ісусе, великий священику, ти та ближні твої, що сидять перед тобою, бо вони мужі знаменні, бо ось Я приведу Свого раба Пагінця.
ZECH|3|9|Бо оце той камінь, що його Я поклав перед Ісусом. На одному камені сім очей. Ось Я вирізьблю на ньому різьбу його, говорить Господь Саваот, і відкину вину цієї землі за один день.
ZECH|3|10|Того дня, говорить Господь Саваот, ви будете кликати один одного під виноград і під фіґове дерево.
ZECH|4|1|І вернувся той Ангол, що говорив зо мною, і збудив мене, як чоловіка, якого будять зо сну його.
ZECH|4|2|І сказав він до мене: Що ти бачиш? А я відказав: Бачу я, ось світильник, увесь із золота, і чаша на верху його, і сім лямпад його на ньому, і по сім рурочок для лямпад, що на верху його.
ZECH|4|3|І дві оливки на ньому, одна з правиці чаші, а одна на лівиці її.
ZECH|4|4|І говорив я й сказав до Ангола, що говорив зо мною, кажучи: Що це, мій пане?
ZECH|4|5|І відповів Ангол, що говорив зо мною, та й сказав мені: Чи ж ти не знаєш, що це таке? А я відказав: Ні, пане!
ZECH|4|6|І відповів він, і сказав мені, говорячи: Оце таке Господнє слово до Зоровавеля: Не силою й не міццю, але тільки Моїм Духом, говорить Господь Саваот.
ZECH|4|7|Хто ти, горо велика? Перед Зоровавелем ти станеш рівниною. І він винесе наріжного каменя при криках: Милість, милість йому!
ZECH|4|8|І було мені слово Господнє таке:
ZECH|4|9|Зоровавелеві руки заклали цей дім, і руки його викінчать, і ти пізнаєш, що Господь Саваот послав мене до вас.
ZECH|4|10|Бо хто буде погорджувати днем малих речей? Але будуть тішитися, і будуть дивитись на теслярського виска в руці Зоровавеля ті семеро, Господні очі, що ходять по всій землі.
ZECH|4|11|І заговорив я та й до нього сказав: Що це за дві оливки праворуч свічника й ліворуч його?
ZECH|4|12|І заговорив я вдруге, та й до нього сказав: Що це за дві галузки оливок, що через дві золоті рурки виливають з себе золото?
ZECH|4|13|І сказав він до мене, говорячи: Хіба ти не знаєш, що це? А я відказав: Ні, пане!
ZECH|4|14|І він сказав: Це два Помазанці, що стоять перед Господом всієї землі.
ZECH|5|1|І знову підніс я свої очі, та й побачив, аж ось летить звій.
ZECH|5|2|І сказав він до мене: Що ти бачиш? А я відказав: Я бачу летючого звоя. Довжина його двадцять мірою ліктем, а ширина його десять ліктів.
ZECH|5|3|І сказав він мені: Це те прокляття, що виходить на поверхню всієї землі. Бо кожен злодій буде безкарний згідно з тим, що з цього боку звою написане, і кожен, хто присягає ложно, буде безкарний згідно з тим, що з того боку звою написане.
ZECH|5|4|І привів Я його, прокляття, говорить Господь Саваот, і прийде воно до дому злодія, і до дому того, хто ложно присягає Йменням Моїм, і воно міцно осядеться в середині дому його, і вигубить його, і дерева його та каміння його.
ZECH|5|5|І вийшов той Ангол, що говорив зо мною, та й до мене сказав: Зведи но свої очі й побач, що це виходить?
ZECH|5|6|І сказав я: Що це таке? А він відказав: Це ефа, що виходить. І ще він сказав: Це їхнє око в усьому Краї.
ZECH|5|7|Аж ось піднялася олив'яна покришка, а це була одна жінка, що сиділа посеред ефи.
ZECH|5|8|І він сказав: Це та несправедливість. І кинув її до середини ефи, і кинув олив'яного куска до її отвору.
ZECH|5|9|І звів я очі свої та й побачив, аж ось дві жінки виходять, і вітер гудів в їхніх крилах, а їхні крила як крила чорногуза. І підняли вони ефу між землею та між небом.
ZECH|5|10|І сказав я до Ангола, що зо мною говорив: Куди вони несуть цю ефу?
ZECH|5|11|І сказав він до мене: Щоб збудувати їй дім у краю Шін'ар. А коли він буде поставлений, то буде покладена там на місці своєму.
ZECH|6|1|І знову звів я очі свої та й побачив, аж ось чотири колесниці виходять з-між двох гір, а ті гори гори з міді.
ZECH|6|2|В колесниці першій коні червоні, а в колесниці другій коні чорні,
ZECH|6|3|а в колесниці третій коні білі, а в колесниці четвертій коні пасасті, міцні.
ZECH|6|4|І відповів я та й сказав до Ангола, що говорив зо мною: Що це таке, мій пане?
ZECH|6|5|І Ангол відповів та й сказав до мене: Це чотири небесні вітри, що виходять після стояння перед Господом усієї землі.
ZECH|6|6|У котрім коні чорні, ті виходять до північного краю, а ті білі вийшли за ними, а ті пасасті вийшли до південного краю,
ZECH|6|7|а ті сильні вийшли й шукали ходи, щоб перейти по землі. І він сказав: Ідіть, ходіть по землі! І ходили вони по землі.
ZECH|6|8|І кликнув він до мене й казав мені, говорячи: Побач, ті, що вийшли до північного краю, заспокоїли духа мого в північному краї.
ZECH|6|9|І було мені слово Господнє таке:
ZECH|6|10|Візьми від вигнання, від Хелдая, і від Товійї, і від Єдаї, і прийдеш ти того дня, і ввійдеш до дому Йошійї, Цефанієвого сина, що прийшли з Вавилону.
ZECH|6|11|І візьмеш срібло та золото, і зробиш корону, і покладеш на голову Ісуса, Єгосадакового сина, великого священика.
ZECH|6|12|І скажеш до нього, говорячи: Так говорить Господь Саваот, промовляючи: Оце муж, Цема ім'я йому, і зо свого місця виросте він, і збудує храма Господнього.
ZECH|6|13|І він збудує храма Господнього, і він буде носити величність, і сяде, і буде панувати на троні своєму, і він стане священиком на троні своєму, і рада миру буде поміж ними обома.
ZECH|6|14|А ті корони будуть Хелдаєві, і Товійї, і Єдаї, і Хенові, сину Цефанії, на пам'ятку в храмі Господньому.
ZECH|6|15|І далекі прийдуть, і побудують у храмі Господньому, і ви пізнаєте, що Господь Саваот послав мене до вас. І це станеться, якщо ви конче будете слухати голосу Господа, вашого Бога!
ZECH|7|1|І сталося, у четвертому році царя Дарія було Господнє слово до Захарія четвертого дня дев'ятого місяця, кіслева.
ZECH|7|2|І послав Бет-Ел Сар'ецера й Реґем-Мелеха та людей його, щоб Господа вблагати,
ZECH|7|3|щоб сказати священикам, які в домі Господа Саваота, та пророкам, говорячи: Чи я маю плакати п'ятого місяця та постити, як я робив це багато років?
ZECH|7|4|І було слово Господа Саваота таке:
ZECH|7|5|Говори до всього народу землі й до священиків, кажучи: Якщо ви постили та лементували п'ятого й сьомого місяця, і то сімдесят років чи то ви постили для Мене?
ZECH|7|6|А коли ви їсте та коли ви п'єте, чи ж то не собі ви їсте й не собі ви п'єте?
ZECH|7|7|Чи ж це не ті слова, які Господь виголошував через давніх пророків, коли Єрусалим був населений та спокійний, і його міста навколо нього, і південь, і рівнина були населені?
ZECH|7|8|І було до Захарія слово Господнє таке:
ZECH|7|9|Так говорить Господь Саваот, промовляючи: Судіть суд по правді, і чиніть один одному милосердя та милість.
ZECH|7|10|А вдови й сироти, чужинця та вбогого не гнобіть, і не думайте зла один одному в серці своєму!
ZECH|7|11|Та вони не хотіли слухати, і відвернули своє рамено від Мене, а вуха свої вчинили тяжкими, щоб не слухати,
ZECH|7|12|і серце своє зробили кременем, щоб не слухати Закону, та тих слів, що послав Господь Саваот Своїм Духом через давніх пророків. І був великий гнів від Господа Саваота.
ZECH|7|13|І сталося, як Я кликав, то вони не слухалися, так вони будуть кликати, та не буду Я слухати, каже Господь Саваот.
ZECH|7|14|І розвіяв Я їх по всіх народах, які не знали їх, а Край був спустошений по них, так що не було такого, хто б переходив чи вертався, і вони зробили улюблений Край спустошенням.
ZECH|8|1|І було мені слово Господнє таке:
ZECH|8|2|Так говорить Господь Саваот: Заздрю Я за Сіон великою заздрістю, і великою ревністю Я заздрю за нього.
ZECH|8|3|Так говорить Господь: Вернуся Я до Сіону, і буду пробувати в середині Єрусалиму, і буде зватися Єрусалим Містом Правди, а гора Господа Саваота горою святою.
ZECH|8|4|Так говорить Господь Саваот: Ще будуть сидіти на єрусалимських майданах діди та баби, і кожен з палицею в своїй руці через довгий вік.
ZECH|8|5|А міські майдани будуть переповнені хлопцями та дівчатами, що будуть бавитися на майданах його.
ZECH|8|6|Так говорить Господь Саваот: Коли дивне це в очах останку народу цього за цих днів, чи ж воно буде дивне в очах Моїх? промовляє Господь Саваот.
ZECH|8|7|Так говорить Господь Саваот: Ото Я спасу Свій народ із східнього краю та з краю заходу сонця.
ZECH|8|8|І спроваджу Я їх, і вони будуть пробувати в середині Єрусалиму, і стануть народом Моїм, а Я стану їм Богом у правді та в праведності.
ZECH|8|9|Так говорить Господь Саваот: Нехай стануть сильними ваші руки, ви, що слухаєте цими днями слова ці з уст пророків, що були в день закладин дому Господа Саваота, храму, щоб був побудований.
ZECH|8|10|Бо перед цими днями не було нагороди для людини, ані нагороди для худоби, і для того, хто виходив, і для того, хто входив не було спокою від ворога, і пускав Я всіх людей одного проти одного.
ZECH|8|11|Тому Я тепер для останку оцього народу не буду такий, як за тих давніх днів, промовляє Господь Саваот.
ZECH|8|12|Бо буде насіння миру: виноград дасть свій плід, а земля урожай свій подасть, а небо дасть росу свою, і вчиню Я, що решта оцього народу це все посяде.
ZECH|8|13|І станеться, як були ви прокляттям серед народів, доме Юдин та доме Ізраїлів, так Я вас спасу, і ви станете благословенням. Не бійтесь, хай зміцніють ваші руки!
ZECH|8|14|Бо так промовляє Господь Саваот: Як Я думав зробити вам зле, коли ваші батьки прогнівляли Мене, промовляє Господь Саваот, і не жалував Я,
ZECH|8|15|так знову задумав Я днями оцими вчинити добро Єрусалимові та Юдиному домові. Не бійтесь!
ZECH|8|16|Оце речі, які будете робити: Говоріть правду один одному, правду та суд миру судіть у ваших брамах.
ZECH|8|17|І не думайте зла в своїм серці один проти одного, і не любіть неправдивої присяги, бо це все оте, що зненавидив Я, промовляє Господь.
ZECH|8|18|І було мені слово Господнє таке:
ZECH|8|19|Так говорить Господь Саваот: Піст четвертого, і піст п'ятого, і піст сьомого, і піст десятого місяця стане для Юдиного дому на радість і на втіху, та на веселі свята, але правду та мир кохайте!
ZECH|8|20|Так говорить Господь Саваот: Ще прийдуть народи та мешканці численних міст.
ZECH|8|21|І прийдуть мешканці одного міста до другого, кажучи: Ходімо, ходімо вблагати Господа, шукати Господа Саваота! Піду також я.
ZECH|8|22|І поприходять численні народи та сильні люди шукати Господа Саваота в Єрусалимі, і благати Господа.
ZECH|8|23|Так говорить Господь Саваот: І станеться тими днями, що схоплять десять мужів з усіх язиків тих народів, і схоплять за полу юдея, говорячи: Ходімо з вами, бо ми чули: Бог з вами!
ZECH|9|1|Пророцтво Господнього слова на землю Хадрах та Дамаск, місця спочинку його, бо око Господнє на Арам та на всі Ізраїлеві племена,
ZECH|9|2|а також на Гамат, що межує із ним, на Тир та Сидон, бо він став дуже мудрий.
ZECH|9|3|І Тир твердиню собі збудував, і срібла нагромадив, як пороху, а щирого золота як багна на вулицях.
ZECH|9|4|Ось Господь зробить бідним його, і на морі поб'є його потугу, і він сам буде пожертий огнем.
ZECH|9|5|Побачить це Ашкелон, та й злякається, і Азза, і дуже настрашиться, і Екрон, бо надія його засоромиться. І згине цар із Аззи, а Ашкелон не буде заселений.
ZECH|9|6|І буде в Ашдоді сидіти байстрюк, і Я вигублю гордість филистимлян.
ZECH|9|7|І викину кров його з його уст, а гидоту його з-між зубів його, і для нашого Бога достанеться й він, і він буде, як князь той у Юді, а Екрон як євусей.
ZECH|9|8|І стану табором біля Свого дому проти війська, проти того, хто переходить і хто вертається; і вже не перейде гнобитель повз них, бо тепер Я це бачив Своїми очима.
ZECH|9|9|Радій вельми, о дочко Сіону, веселись, дочко Єрусалиму! Ось Цар твій до тебе гряде, справедливий і повний спасіння, покірний, і їде на ослі, і на молодім віслюкові, сині ослиці.
ZECH|9|10|І вигублю Я колесниці з Єфрема, і коня з Єрусалиму, і військовий лук знищений буде. І народам Він мир сповістить, а Його панування від моря до моря, і від Ріки аж до кінців землі.
ZECH|9|11|Також ти, за кров заповіту твого Я пустив твоїх в'язнів із ями, в якій немає води.
ZECH|9|12|До твердині верніться, о в'язні надії! І сьогодні звіщаю: Подвійно тобі поверну!
ZECH|9|13|Бо Юду собі натягну, немов лука, наповню Єфремом його, і збуджу твоїх синів, Сіоне, на синів твоїх, Яване, і вчиню Я тебе за меча для лицарства.
ZECH|9|14|А Господь з'явиться над ними, і стріла Його вийде, як блискавка, і Господь Бог засурмить у сурму, і піде південними бурями.
ZECH|9|15|І Господь Саваот берегтиме всіх їх, і вони поїдять та потопчуть каміння, що кидається, і вони будуть пити та будуть шуміти, немов те вино, і будуть повні, як чаша жертовна, неначе ті роги жертівника.
ZECH|9|16|І спасе їх Господь, їхній Бог, того дня, Свій народ, як отару, бо вони, як каміння корони, засяють у Краї Його.
ZECH|9|17|і що за добро Його буде, і що за краса Його! Збіжжя поможе рости юнакам, а дівчатам вино молоде.
ZECH|10|1|Просіть від Господа дощу часу весняного пізнього дощу, Господь чинить блискавки, і зливний дощ посилає їм, кожному траву на полі.
ZECH|10|2|Бо говорять марноту домові божки, і віщуни бачать лжу, і розказують сни неправдиві, потішають марнотою. Тому вони бродять, немов та отара, мандрують вони, бо без пастиря.
ZECH|10|3|На пастирів гнів Мій палає, а козлів навіщу, бо стадо Своє, Юдин дім покарає Господь Саваот, і вчинить Він їх, немов Своїм славним конем на війні.
ZECH|10|4|З нього буде наріжник, із нього кілок, з нього лук бойовий, з нього вийдуть керманичі разом усі,
ZECH|10|5|І будуть, немов те лицарство, що топче воно на війні, як болото на вулицях, і будуть вони воювати, бо з ними Господь, і кіннотних їздців засоромляться.
ZECH|10|6|І вчиню Я лицарським дім Юдин, а дім Йосипів спасу, і верну їх, бо змилосердивсь над ними, і стануть вони, ніби Я їх не кидав, Бо Я Господь Бог їхній, і буду Я їх вислуховувати.
ZECH|10|7|І стане лицарським Єфрем, і звеселіє їхнє серце, немов від вина, а їхні сини це побачать та будуть радіти, потішиться серце їхнє Господом.
ZECH|10|8|Я їм дам знака та їх позбираю, бо Я викупив їх, і множитись будуть, як множились.
ZECH|10|9|І розсію Я їх між народами, і в далеких краях вони будуть Мене згадувати, і житимуть з дітьми своїми, і вернуться.
ZECH|10|10|І верну їх із краю єгипетського, і позгромаджую їх із Ашшуру, і введу їх до краю Ґілеаду й Лівану, і місця не вистачить їм.
ZECH|10|11|І прийде по морі нещастя, і хвилі на морі ударить, і повисихають усі глибини Ріки, і буде понижена гордість Ашшуру, і від Єгипту відійметься берло.
ZECH|10|12|І зміцню їх у Господі, і Йменням Його вони будуть ходити, говорить Господь!
ZECH|11|1|Ліване, відкрий свої двері, і огонь пожере з твоїх кедрів!
ZECH|11|2|Голоси, кипарисе, бо кедр он упав, пограбовані пишні! Голосіте, башанські дуби, бо ліс неприступний звалився!
ZECH|11|3|Чути голос виття пастухів, бо гордощі їхні пограбовані! Чути рик левчуків, бо йорданська краса попустошена...
ZECH|11|4|Так говорить Господь, мій Бог: Паси ти отару, яка на заріз,
ZECH|11|5|що ріжуть їх їхні купці і не винні, а їхні продавці промовляють: Благословенний Господь, що я збагатів! А їхні пастухи не помилують їх!...
ZECH|11|6|Бо Я не помилую більше вже мешканців цеї землі, промовляє Господь. І ось передам Я людину, одного одному до рук, та до рук царя їхнього, і землю вони потовчуть, і Я з їхніх рук не врятую нікого!
ZECH|11|7|І пас Я отару, яка на заріз тим, хто торгує отарою. І взяв Я Собі два киї, і одного назвав: Милість, а одного назвав: Згода, і пас Я отару.
ZECH|11|8|І знищив Я трьох пастухів за один місяць. І Я втратив терпіння до них, бо душа їхня обридила Мене.
ZECH|11|9|Тому Я сказав: Не пастиму вас! Та вівця, що має померти, нехай умре, а що має погублена бути хай буде погублена, а позосталі хай тіло одна однієї з'їдять!
ZECH|11|10|І Я взяв Свого кия Милість, і його поламав, щоб зламати Свого заповіта, якого Я склав був зо всіма народами.
ZECH|11|11|І він зламаний був того дня, і пізнали покупці отари, які на Мене вважають, що це слово Господнє.
ZECH|11|12|І сказав Я до них: Якщо добре це в ваших очах, дайте платню Мою, а як ні, перестаньте! І вони Мою платню відважили тридцять срібняків.
ZECH|11|13|І промовив до мене Господь: Кинь її ганчареві, ту славну ціну, що вони оцінили Мене! І Я взяв оті тридцять срібняків, і те кинув до дому Господнього, до ганчаря.
ZECH|11|14|І зламав Я Свого кия другого, Згоду, щоб зламати братерство між Юдою та між Ізраїлем.
ZECH|11|15|І промовив до мене Господь: Ще візьми собі знаряддя пастуха нерозумного.
ZECH|11|16|Бо ось Я настановлю пастиря на землі, він загублених не відвідає, розпорошеного не буде шукати, і зламаної не вилікує, стоячої не годуватиме, а м'ясо ситої їстиме, і ратиці їхні поламає.
ZECH|11|17|Горе негідному пастиреві, який покидає отару! Меч на рамено його та в його праве око: конче всохне рамено йому, і конче стемніє його праве око!
ZECH|12|1|Пророцтво Господнього слова на Ізраїля. Говорить Господь, що небо напнув та землю заклав, і вформував дух людині у нутрі її:
ZECH|12|2|Ось Я Єрусалим учиню за келіха оп'яніння всім народам навколо, і на Юду також, коли буде в облозі на Єрусалим.
ZECH|12|3|І буде в той день, Я зроблю Єрусалима за камінь тяжкий всім народам: усі, хто буде його порушати, будуть конче поранені, і зберуться на нього всі народи землі.
ZECH|12|4|Того дня, промовляє Господь, ударю всіх коней сполошенням, і шаленством його верхівця, а над Юдиним домом відкрию Я очі Свої, і всіх коней народів поб'ю сліпотою.
ZECH|12|5|І скажуть тоді князі Юдині в серці своєму: Моя потуга то мешканці Єрусалиму у Господі Саваоті, їхньому Бозі!
ZECH|12|6|Того дня Я вчиню князів Юди, немов ту жаровню з огнем між дровами, і як палаючий смолоскип між снопами, і будуть вони пожирати праворуч і ліворуч всі довкільні народи. І знову осяде на місці своєму Єрусалим, у Єрусалимі.
ZECH|12|7|І Господь допоможе найперше Юдиним наметам, щоб не збільшилась слава Давидового дому та єрусалимського мешканця понад Юду.
ZECH|12|8|Того дня оборонить Господь єрусалимського мешканця, і буде того дня той, хто спотикається серед них, як Давид, а дім Давидів як Бог, як Ангол Господній перед ними.
ZECH|12|9|І станеться в день той, і Я буду шукати, щоб понищити всі ті народи, що приходять на Єрусалим.
ZECH|12|10|А на Давидів дім та на єрусалимського мешканця Я виллю Духа милости та молитви. І будуть дивитись на Мене, Кого прокололи, і будуть за Ним голосити, як голоситься за одинцем, і гірко заплачуть за Ним, як плачуть за первенцем.
ZECH|12|11|Того дня здійметься велике голосіння в Єрусалимі, як голосіння Гададріммона в Меґіддонській долині.
ZECH|12|12|І буде земля голосити, кожен рід окремо: окремо рід дому Давида, і окремо жінки їх, окремо рід дому Натана, й окремо жінки їх,
ZECH|12|13|окремо рід дому Левія, і окремо жінки їх, окремо рід Шім'ї, і окремо жінки їх.
ZECH|12|14|Усі роди, які позостали, кожен рід окремо, і окремо жінки їх.
ZECH|13|1|Того дня відкриється джерело для Давидового дому та для єрусалимських мешканців для жертви за гріх і за нечистоту.
ZECH|13|2|І станеться в день той, говорить Господь Саваот, повигублюю ймення бовванів з землі, і не будуть вони більше згадуватись, бо й пророків та духа нечистого виведу Я із землі!
ZECH|13|3|І станеться, коли буде хто пророкувати ще, то скажуть йому його батько та мати його, що його породили: Не будеш ти жити, бо ложне говориш Господнім Ім'ям! І заколють його його батько та мати його, що його породили, за те, що неправду він пророкував.
ZECH|13|4|І станеться в день той, посоромлені будуть пророки оті, кожен видінням своїм, коли пророкував він, і волосяниці не будуть вони зодягати, щоб обманювати.
ZECH|13|5|І скаже він: Я не пророк, я людина, що порає землю, бо земля мій набуток з юнацтва мого.
ZECH|13|6|А коли йому скаже хто: Що це за рани на твоїх руках? то відкаже: Побито мене в домі тих, хто кохає мене...
ZECH|13|7|О мечу, збудися на Мого пастиря та на мужа, Мого товариша, каже Господь Саваот! Удар пастиря і розпорошаться вівці, і Я оберну на малих Свою руку.
ZECH|13|8|І станеться в цілому Краї, говорить Господь, дві частині в нім витяті будуть, помруть, а третя частина зоставлена буде у ньому.
ZECH|13|9|І цю третю частину введу на огонь, і очищу їх, як очищається срібло, і їх випробую, як випробовується оте золото. Він кликати буде Ймення Моє, і Я йому відповім і скажу: Це народ Мій, а він скаже: Господь то мій Бог!
ZECH|14|1|Ось день настає для Господа, і серед тебе поділена буде здобич.
ZECH|14|2|І зберу всі народи до Єрусалиму на бій, і буде здобуте це місто, і пограбовані будуть доми, а жінки побезчещені. І вийде півміста в полон на вигнання, а решта народу не буде погублена з міста.
ZECH|14|3|І вийде Господь, і стане на прю із народами цими, як дня боротьби Його, за дня бою.
ZECH|14|4|І того дня стануть ноги Його на Оливній горі, що перед Єрусалимом зо сходу, а Оливна гора на свої половини роздвоїться, на схід і на захід, на дуже велику долину. І на північ осунеться половина гори, а половина її на південь.
ZECH|14|5|І втікати ви будете в долину Моїх гір, бо долина гірська сягатиме по Ацал. І втікати ви будете, як утікали перед землетрусом за днів Уззійї, царя Юдиного. І прийде Господь, Бог мій, і з Ним усі святі.
ZECH|14|6|І станеться в день той, світла не буде, і буде холод та замерзання.
ZECH|14|7|І буде єдиний то день, Господу знаний, то буде не день, і не ніч, і буде, на час вечора станеться світло.
ZECH|14|8|І станеться в день той, вийде з Єрусалиму живая вода, половина її до східнього моря, а половина її до моря західнього. Літом і зимою це буде.
ZECH|14|9|І стане Господь за царя над землею всією, Господь буде один того дня, і одне Ймення Його.
ZECH|14|10|Уся ця земля стане степом від Ґеви до Ріммону, на південь Єрусалиму, який стане високим, і пробуватиме на місці своєму від брами Веніямина аж до місця Першої брами, аж до брами Наріжинків, і від башти Хананеїла аж до царського чавила.
ZECH|14|11|І осядуть у ньому, і закляття вже більше не буде, і безпечно сидітиме Єрусалим.
ZECH|14|12|А оце буде рана, що нею поранить Господь всі народи, хто піде війною на Єрусалим: згниє тіло його, хоч він на ногах своїх буде стояти, і очі йому погниють в своїх ямках, і язик його погниє в своїх устах.
ZECH|14|13|І станеться в день той, між ними настане велике збентеження, і схопить один руку одного, і підійметься рука його понад руку свого ближнього.
ZECH|14|14|І навіть Юда воюватиме в Єрусалимі, і буде згромаджений маєток всіх навкільних народів, золото й срібло та одіж, дуже багато.
ZECH|14|15|І буде такий самий удар на коня, мула, верблюда й осла, та на всяку худобу, що буде в таборах у них, як пораза оця.
ZECH|14|16|І станеться, що позосталі з усіх тих народів, що приходили на Єрусалим, то будуть приходити з року на рік, щоб вклонятись Цареві, Господу Саваоту, і щоб святкувати свято Кучок.
ZECH|14|17|І станеться, хто від земних племен до Єрусалиму не прийде, щоб вклонятись Цареві, Господу Саваоту, то не буде дощу в них.
ZECH|14|18|А якщо не прийде племено єгипетське, і не ввійде всередину, то буде на них та пораза, якою народи ударить Господь, хто святкувати свято Кучок не прийде.
ZECH|14|19|Оце гріх Єгиптові буде, і гріх всім народам, хто святкувати свято Кучок не прийде.
ZECH|14|20|Буде того дня на кінських дзвінках: Святе Господеві, і будуть горнята в Господньому домі, немов ті кропильниці перед жертовником.
ZECH|14|21|І буде усяке горня в Єрусалимі та в Юді святістю для Господа Саваота, і будуть приходити всі, хто жертву приносить, і будуть з них брати й варитимуть в них. І того дня не буде вже більше купця в домі Господа Саваота.
