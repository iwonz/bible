EZRA|1|1|Now in the first year of Cyrus king of Persia, that the word of the LORD by the mouth of Jeremiah might be fulfilled, the LORD stirred up the spirit of Cyrus king of Persia, that he made a proclamation throughout all his kingdom, and put it also in writing, saying,
EZRA|1|2|Thus saith Cyrus king of Persia, The LORD God of heaven hath given me all the kingdoms of the earth; and he hath charged me to build him an house at Jerusalem, which is in Judah.
EZRA|1|3|Who is there among you of all his people? his God be with him, and let him go up to Jerusalem, which is in Judah, and build the house of the LORD God of Israel, (he is the God,) which is in Jerusalem.
EZRA|1|4|And whosoever remaineth in any place where he sojourneth, let the men of his place help him with silver, and with gold, and with goods, and with beasts, beside the freewill offering for the house of God that is in Jerusalem.
EZRA|1|5|Then rose up the chief of the fathers of Judah and Benjamin, and the priests, and the Levites, with all them whose spirit God had raised, to go up to build the house of the LORD which is in Jerusalem.
EZRA|1|6|And all they that were about them strengthened their hands with vessels of silver, with gold, with goods, and with beasts, and with precious things, beside all that was willingly offered.
EZRA|1|7|Also Cyrus the king brought forth the vessels of the house of the LORD, which Nebuchadnezzar had brought forth out of Jerusalem, and had put them in the house of his gods;
EZRA|1|8|Even those did Cyrus king of Persia bring forth by the hand of Mithredath the treasurer, and numbered them unto Sheshbazzar, the prince of Judah.
EZRA|1|9|And this is the number of them: thirty chargers of gold, a thousand chargers of silver, nine and twenty knives,
EZRA|1|10|Thirty basins of gold, silver basins of a second sort four hundred and ten, and other vessels a thousand.
EZRA|1|11|All the vessels of gold and of silver were five thousand and four hundred. All these did Sheshbazzar bring up with them of the captivity that were brought up from Babylon unto Jerusalem.
EZRA|2|1|Now these are the children of the province that went up out of the captivity, of those which had been carried away, whom Nebuchadnezzar the king of Babylon had carried away unto Babylon, and came again unto Jerusalem and Judah, every one unto his city;
EZRA|2|2|Which came with Zerubbabel: Jeshua, Nehemiah, Seraiah, Reelaiah, Mordecai, Bilshan, Mizpar, Bigvai, Rehum, Baanah. The number of the men of the people of Israel:
EZRA|2|3|The children of Parosh, two thousand an hundred seventy and two.
EZRA|2|4|The children of Shephatiah, three hundred seventy and two.
EZRA|2|5|The children of Arah, seven hundred seventy and five.
EZRA|2|6|The children of Pahathmoab, of the children of Jeshua and Joab, two thousand eight hundred and twelve.
EZRA|2|7|The children of Elam, a thousand two hundred fifty and four.
EZRA|2|8|The children of Zattu, nine hundred forty and five.
EZRA|2|9|The children of Zaccai, seven hundred and threescore.
EZRA|2|10|The children of Bani, six hundred forty and two.
EZRA|2|11|The children of Bebai, six hundred twenty and three.
EZRA|2|12|The children of Azgad, a thousand two hundred twenty and two.
EZRA|2|13|The children of Adonikam, six hundred sixty and six.
EZRA|2|14|The children of Bigvai, two thousand fifty and six.
EZRA|2|15|The children of Adin, four hundred fifty and four.
EZRA|2|16|The children of Ater of Hezekiah, ninety and eight.
EZRA|2|17|The children of Bezai, three hundred twenty and three.
EZRA|2|18|The children of Jorah, an hundred and twelve.
EZRA|2|19|The children of Hashum, two hundred twenty and three.
EZRA|2|20|The children of Gibbar, ninety and five.
EZRA|2|21|The children of Bethlehem, an hundred twenty and three.
EZRA|2|22|The men of Netophah, fifty and six.
EZRA|2|23|The men of Anathoth, an hundred twenty and eight.
EZRA|2|24|The children of Azmaveth, forty and two.
EZRA|2|25|The children of Kirjatharim, Chephirah, and Beeroth, seven hundred and forty and three.
EZRA|2|26|The children of Ramah and Gaba, six hundred twenty and one.
EZRA|2|27|The men of Michmas, an hundred twenty and two.
EZRA|2|28|The men of Bethel and Ai, two hundred twenty and three.
EZRA|2|29|The children of Nebo, fifty and two.
EZRA|2|30|The children of Magbish, an hundred fifty and six.
EZRA|2|31|The children of the other Elam, a thousand two hundred fifty and four.
EZRA|2|32|The children of Harim, three hundred and twenty.
EZRA|2|33|The children of Lod, Hadid, and Ono, seven hundred twenty and five.
EZRA|2|34|The children of Jericho, three hundred forty and five.
EZRA|2|35|The children of Senaah, three thousand and six hundred and thirty.
EZRA|2|36|The priests: the children of Jedaiah, of the house of Jeshua, nine hundred seventy and three.
EZRA|2|37|The children of Immer, a thousand fifty and two.
EZRA|2|38|The children of Pashur, a thousand two hundred forty and seven.
EZRA|2|39|The children of Harim, a thousand and seventeen.
EZRA|2|40|The Levites: the children of Jeshua and Kadmiel, of the children of Hodaviah, seventy and four.
EZRA|2|41|The singers: the children of Asaph, an hundred twenty and eight.
EZRA|2|42|The children of the porters: the children of Shallum, the children of Ater, the children of Talmon, the children of Akkub, the children of Hatita, the children of Shobai, in all an hundred thirty and nine.
EZRA|2|43|The Nethinims: the children of Ziha, the children of Hasupha, the children of Tabbaoth,
EZRA|2|44|The children of Keros, the children of Siaha, the children of Padon,
EZRA|2|45|The children of Lebanah, the children of Hagabah, the children of Akkub,
EZRA|2|46|The children of Hagab, the children of Shalmai, the children of Hanan,
EZRA|2|47|The children of Giddel, the children of Gahar, the children of Reaiah,
EZRA|2|48|The children of Rezin, the children of Nekoda, the children of Gazzam,
EZRA|2|49|The children of Uzza, the children of Paseah, the children of Besai,
EZRA|2|50|The children of Asnah, the children of Mehunim, the children of Nephusim,
EZRA|2|51|The children of Bakbuk, the children of Hakupha, the children of Harhur,
EZRA|2|52|The children of Bazluth, the children of Mehida, the children of Harsha,
EZRA|2|53|The children of Barkos, the children of Sisera, the children of Thamah,
EZRA|2|54|The children of Neziah, the children of Hatipha.
EZRA|2|55|The children of Solomon's servants: the children of Sotai, the children of Sophereth, the children of Peruda,
EZRA|2|56|The children of Jaalah, the children of Darkon, the children of Giddel,
EZRA|2|57|The children of Shephatiah, the children of Hattil, the children of Pochereth of Zebaim, the children of Ami.
EZRA|2|58|All the Nethinims, and the children of Solomon's servants, were three hundred ninety and two.
EZRA|2|59|And these were they which went up from Telmelah, Telharsa, Cherub, Addan, and Immer: but they could not shew their father's house, and their seed, whether they were of Israel:
EZRA|2|60|The children of Delaiah, the children of Tobiah, the children of Nekoda, six hundred fifty and two.
EZRA|2|61|And of the children of the priests: the children of Habaiah, the children of Koz, the children of Barzillai; which took a wife of the daughters of Barzillai the Gileadite, and was called after their name:
EZRA|2|62|These sought their register among those that were reckoned by genealogy, but they were not found: therefore were they, as polluted, put from the priesthood.
EZRA|2|63|And the Tirshatha said unto them, that they should not eat of the most holy things, till there stood up a priest with Urim and with Thummim.
EZRA|2|64|The whole congregation together was forty and two thousand three hundred and threescore,
EZRA|2|65|Beside their servants and their maids, of whom there were seven thousand three hundred thirty and seven: and there were among them two hundred singing men and singing women.
EZRA|2|66|Their horses were seven hundred thirty and six; their mules, two hundred forty and five;
EZRA|2|67|Their camels, four hundred thirty and five; their asses, six thousand seven hundred and twenty.
EZRA|2|68|And some of the chief of the fathers, when they came to the house of the LORD which is at Jerusalem, offered freely for the house of God to set it up in his place:
EZRA|2|69|They gave after their ability unto the treasure of the work threescore and one thousand drams of gold, and five thousand pound of silver, and one hundred priests' garments.
EZRA|2|70|So the priests, and the Levites, and some of the people, and the singers, and the porters, and the Nethinims, dwelt in their cities, and all Israel in their cities.
EZRA|3|1|And when the seventh month was come, and the children of Israel were in the cities, the people gathered themselves together as one man to Jerusalem.
EZRA|3|2|Then stood up Jeshua the son of Jozadak, and his brethren the priests, and Zerubbabel the son of Shealtiel, and his brethren, and builded the altar of the God of Israel, to offer burnt offerings thereon, as it is written in the law of Moses the man of God.
EZRA|3|3|And they set the altar upon his bases; for fear was upon them because of the people of those countries: and they offered burnt offerings thereon unto the LORD, even burnt offerings morning and evening.
EZRA|3|4|They kept also the feast of tabernacles, as it is written, and offered the daily burnt offerings by number, according to the custom, as the duty of every day required;
EZRA|3|5|And afterward offered the continual burnt offering, both of the new moons, and of all the set feasts of the LORD that were consecrated, and of every one that willingly offered a freewill offering unto the LORD.
EZRA|3|6|From the first day of the seventh month began they to offer burnt offerings unto the LORD. But the foundation of the temple of the LORD was not yet laid.
EZRA|3|7|They gave money also unto the masons, and to the carpenters; and meat, and drink, and oil, unto them of Zidon, and to them of Tyre, to bring cedar trees from Lebanon to the sea of Joppa, according to the grant that they had of Cyrus king of Persia.
EZRA|3|8|Now in the second year of their coming unto the house of God at Jerusalem, in the second month, began Zerubbabel the son of Shealtiel, and Jeshua the son of Jozadak, and the remnant of their brethren the priests and the Levites, and all they that were come out of the captivity unto Jerusalem; and appointed the Levites, from twenty years old and upward, to set forward the work of the house of the LORD.
EZRA|3|9|Then stood Jeshua with his sons and his brethren, Kadmiel and his sons, the sons of Judah, together, to set forward the workmen in the house of God: the sons of Henadad, with their sons and their brethren the Levites.
EZRA|3|10|And when the builders laid the foundation of the temple of the LORD, they set the priests in their apparel with trumpets, and the Levites the sons of Asaph with cymbals, to praise the LORD, after the ordinance of David king of Israel.
EZRA|3|11|And they sang together by course in praising and giving thanks unto the LORD; because he is good, for his mercy endureth for ever toward Israel. And all the people shouted with a great shout, when they praised the LORD, because the foundation of the house of the LORD was laid.
EZRA|3|12|But many of the priests and Levites and chief of the fathers, who were ancient men, that had seen the first house, when the foundation of this house was laid before their eyes, wept with a loud voice; and many shouted aloud for joy:
EZRA|3|13|So that the people could not discern the noise of the shout of joy from the noise of the weeping of the people: for the people shouted with a loud shout, and the noise was heard afar off.
EZRA|4|1|Now when the adversaries of Judah and Benjamin heard that the children of the captivity builded the temple unto the LORD God of Israel;
EZRA|4|2|Then they came to Zerubbabel, and to the chief of the fathers, and said unto them, Let us build with you: for we seek your God, as ye do; and we do sacrifice unto him since the days of Esarhaddon king of Assur, which brought us up hither.
EZRA|4|3|But Zerubbabel, and Jeshua, and the rest of the chief of the fathers of Israel, said unto them, Ye have nothing to do with us to build an house unto our God; but we ourselves together will build unto the LORD God of Israel, as king Cyrus the king of Persia hath commanded us.
EZRA|4|4|Then the people of the land weakened the hands of the people of Judah, and troubled them in building,
EZRA|4|5|And hired counsellors against them, to frustrate their purpose, all the days of Cyrus king of Persia, even until the reign of Darius king of Persia.
EZRA|4|6|And in the reign of Ahasuerus, in the beginning of his reign, wrote they unto him an accusation against the inhabitants of Judah and Jerusalem.
EZRA|4|7|And in the days of Artaxerxes wrote Bishlam, Mithredath, Tabeel, and the rest of their companions, unto Artaxerxes king of Persia; and the writing of the letter was written in the Syrian tongue, and interpreted in the Syrian tongue.
EZRA|4|8|Rehum the chancellor and Shimshai the scribe wrote a letter against Jerusalem to Artaxerxes the king in this sort:
EZRA|4|9|Then wrote Rehum the chancellor, and Shimshai the scribe, and the rest of their companions; the Dinaites, the Apharsathchites, the Tarpelites, the Apharsites, the Archevites, the Babylonians, the Susanchites, the Dehavites, and the Elamites,
EZRA|4|10|And the rest of the nations whom the great and noble Asnapper brought over, and set in the cities of Samaria, and the rest that are on this side the river, and at such a time.
EZRA|4|11|This is the copy of the letter that they sent unto him, even unto Artaxerxes the king; Thy servants the men on this side the river, and at such a time.
EZRA|4|12|Be it known unto the king, that the Jews which came up from thee to us are come unto Jerusalem, building the rebellious and the bad city, and have set up the walls thereof, and joined the foundations.
EZRA|4|13|Be it known now unto the king, that, if this city be builded, and the walls set up again, then will they not pay toll, tribute, and custom, and so thou shalt endamage the revenue of the kings.
EZRA|4|14|Now because we have maintenance from the king's palace, and it was not meet for us to see the king's dishonour, therefore have we sent and certified the king;
EZRA|4|15|That search may be made in the book of the records of thy fathers: so shalt thou find in the book of the records, and know that this city is a rebellious city, and hurtful unto kings and provinces, and that they have moved sedition within the same of old time: for which cause was this city destroyed.
EZRA|4|16|We certify the king that, if this city be builded again, and the walls thereof set up, by this means thou shalt have no portion on this side the river.
EZRA|4|17|Then sent the king an answer unto Rehum the chancellor, and to Shimshai the scribe, and to the rest of their companions that dwell in Samaria, and unto the rest beyond the river, Peace, and at such a time.
EZRA|4|18|The letter which ye sent unto us hath been plainly read before me.
EZRA|4|19|And I commanded, and search hath been made, and it is found that this city of old time hath made insurrection against kings, and that rebellion and sedition have been made therein.
EZRA|4|20|There have been mighty kings also over Jerusalem, which have ruled over all countries beyond the river; and toll, tribute, and custom, was paid unto them.
EZRA|4|21|Give ye now commandment to cause these men to cease, and that this city be not builded, until another commandment shall be given from me.
EZRA|4|22|Take heed now that ye fail not to do this: why should damage grow to the hurt of the kings?
EZRA|4|23|Now when the copy of king Artaxerxes' letter was read before Rehum, and Shimshai the scribe, and their companions, they went up in haste to Jerusalem unto the Jews, and made them to cease by force and power.
EZRA|4|24|Then ceased the work of the house of God which is at Jerusalem. So it ceased unto the second year of the reign of Darius king of Persia.
EZRA|5|1|Then the prophets, Haggai the prophet, and Zechariah the son of Iddo, prophesied unto the Jews that were in Judah and Jerusalem in the name of the God of Israel, even unto them.
EZRA|5|2|Then rose up Zerubbabel the son of Shealtiel, and Jeshua the son of Jozadak, and began to build the house of God which is at Jerusalem: and with them were the prophets of God helping them.
EZRA|5|3|At the same time came to them Tatnai, governor on this side the river, and Shetharboznai and their companions, and said thus unto them, Who hath commanded you to build this house, and to make up this wall?
EZRA|5|4|Then said we unto them after this manner, What are the names of the men that make this building?
EZRA|5|5|But the eye of their God was upon the elders of the Jews, that they could not cause them to cease, till the matter came to Darius: and then they returned answer by letter concerning this matter.
EZRA|5|6|The copy of the letter that Tatnai, governor on this side the river, and Shetharboznai and his companions the Apharsachites, which were on this side the river, sent unto Darius the king:
EZRA|5|7|They sent a letter unto him, wherein was written thus; Unto Darius the king, all peace.
EZRA|5|8|Be it known unto the king, that we went into the province of Judea, to the house of the great God, which is builded with great stones, and timber is laid in the walls, and this work goeth fast on, and prospereth in their hands.
EZRA|5|9|Then asked we those elders, and said unto them thus, Who commanded you to build this house, and to make up these walls?
EZRA|5|10|We asked their names also, to certify thee, that we might write the names of the men that were the chief of them.
EZRA|5|11|And thus they returned us answer, saying, We are the servants of the God of heaven and earth, and build the house that was builded these many years ago, which a great king of Israel builded and set up.
EZRA|5|12|But after that our fathers had provoked the God of heaven unto wrath, he gave them into the hand of Nebuchadnezzar the king of Babylon, the Chaldean, who destroyed this house, and carried the people away into Babylon.
EZRA|5|13|But in the first year of Cyrus the king of Babylon the same king Cyrus made a decree to build this house of God.
EZRA|5|14|And the vessels also of gold and silver of the house of God, which Nebuchadnezzar took out of the temple that was in Jerusalem, and brought them into the temple of Babylon, those did Cyrus the king take out of the temple of Babylon, and they were delivered unto one, whose name was Sheshbazzar, whom he had made governor;
EZRA|5|15|And said unto him, Take these vessels, go, carry them into the temple that is in Jerusalem, and let the house of God be builded in his place.
EZRA|5|16|Then came the same Sheshbazzar, and laid the foundation of the house of God which is in Jerusalem: and since that time even until now hath it been in building, and yet it is not finished.
EZRA|5|17|Now therefore, if it seem good to the king, let there be search made in the king's treasure house, which is there at Babylon, whether it be so, that a decree was made of Cyrus the king to build this house of God at Jerusalem, and let the king send his pleasure to us concerning this matter.
EZRA|6|1|Then Darius the king made a decree, and search was made in the house of the rolls, where the treasures were laid up in Babylon.
EZRA|6|2|And there was found at Achmetha, in the palace that is in the province of the Medes, a roll, and therein was a record thus written:
EZRA|6|3|In the first year of Cyrus the king the same Cyrus the king made a decree concerning the house of God at Jerusalem, Let the house be builded, the place where they offered sacrifices, and let the foundations thereof be strongly laid; the height thereof threescore cubits, and the breadth thereof threescore cubits;
EZRA|6|4|With three rows of great stones, and a row of new timber: and let the expenses be given out of the king's house:
EZRA|6|5|And also let the golden and silver vessels of the house of God, which Nebuchadnezzar took forth out of the temple which is at Jerusalem, and brought unto Babylon, be restored, and brought again unto the temple which is at Jerusalem, every one to his place, and place them in the house of God.
EZRA|6|6|Now therefore, Tatnai, governor beyond the river, Shetharboznai, and your companions the Apharsachites, which are beyond the river, be ye far from thence:
EZRA|6|7|Let the work of this house of God alone; let the governor of the Jews and the elders of the Jews build this house of God in his place.
EZRA|6|8|Moreover I make a decree what ye shall do to the elders of these Jews for the building of this house of God: that of the king's goods, even of the tribute beyond the river, forthwith expenses be given unto these men, that they be not hindered.
EZRA|6|9|And that which they have need of, both young bullocks, and rams, and lambs, for the burnt offerings of the God of heaven, wheat, salt, wine, and oil, according to the appointment of the priests which are at Jerusalem, let it be given them day by day without fail:
EZRA|6|10|That they may offer sacrifices of sweet savours unto the God of heaven, and pray for the life of the king, and of his sons.
EZRA|6|11|Also I have made a decree, that whosoever shall alter this word, let timber be pulled down from his house, and being set up, let him be hanged thereon; and let his house be made a dunghill for this.
EZRA|6|12|And the God that hath caused his name to dwell there destroy all kings and people, that shall put to their hand to alter and to destroy this house of God which is at Jerusalem. I Darius have made a decree; let it be done with speed.
EZRA|6|13|Then Tatnai, governor on this side the river, Shetharboznai, and their companions, according to that which Darius the king had sent, so they did speedily.
EZRA|6|14|And the elders of the Jews builded, and they prospered through the prophesying of Haggai the prophet and Zechariah the son of Iddo. And they builded, and finished it, according to the commandment of the God of Israel, and according to the commandment of Cyrus, and Darius, and Artaxerxes king of Persia.
EZRA|6|15|And this house was finished on the third day of the month Adar, which was in the sixth year of the reign of Darius the king.
EZRA|6|16|And the children of Israel, the priests, and the Levites, and the rest of the children of the captivity, kept the dedication of this house of God with joy.
EZRA|6|17|And offered at the dedication of this house of God an hundred bullocks, two hundred rams, four hundred lambs; and for a sin offering for all Israel, twelve he goats, according to the number of the tribes of Israel.
EZRA|6|18|And they set the priests in their divisions, and the Levites in their courses, for the service of God, which is at Jerusalem; as it is written in the book of Moses.
EZRA|6|19|And the children of the captivity kept the passover upon the fourteenth day of the first month.
EZRA|6|20|For the priests and the Levites were purified together, all of them were pure, and killed the passover for all the children of the captivity, and for their brethren the priests, and for themselves.
EZRA|6|21|And the children of Israel, which were come again out of captivity, and all such as had separated themselves unto them from the filthiness of the heathen of the land, to seek the LORD God of Israel, did eat,
EZRA|6|22|And kept the feast of unleavened bread seven days with joy: for the LORD had made them joyful, and turned the heart of the king of Assyria unto them, to strengthen their hands in the work of the house of God, the God of Israel.
EZRA|7|1|Now after these things, in the reign of Artaxerxes king of Persia, Ezra the son of Seraiah, the son of Azariah, the son of Hilkiah,
EZRA|7|2|The son of Shallum, the son of Zadok, the son of Ahitub,
EZRA|7|3|The son of Amariah, the son of Azariah, the son of Meraioth,
EZRA|7|4|The son of Zerahiah, the son of Uzzi, the son of Bukki,
EZRA|7|5|The son of Abishua, the son of Phinehas, the son of Eleazar, the son of Aaron the chief priest:
EZRA|7|6|This Ezra went up from Babylon; and he was a ready scribe in the law of Moses, which the LORD God of Israel had given: and the king granted him all his request, according to the hand of the LORD his God upon him.
EZRA|7|7|And there went up some of the children of Israel, and of the priests, and the Levites, and the singers, and the porters, and the Nethinims, unto Jerusalem, in the seventh year of Artaxerxes the king.
EZRA|7|8|And he came to Jerusalem in the fifth month, which was in the seventh year of the king.
EZRA|7|9|For upon the first day of the first month began he to go up from Babylon, and on the first day of the fifth month came he to Jerusalem, according to the good hand of his God upon him.
EZRA|7|10|For Ezra had prepared his heart to seek the law of the LORD, and to do it, and to teach in Israel statutes and judgments.
EZRA|7|11|Now this is the copy of the letter that the king Artaxerxes gave unto Ezra the priest, the scribe, even a scribe of the words of the commandments of the LORD, and of his statutes to Israel.
EZRA|7|12|Artaxerxes, king of kings, unto Ezra the priest, a scribe of the law of the God of heaven, perfect peace, and at such a time.
EZRA|7|13|I make a decree, that all they of the people of Israel, and of his priests and Levites, in my realm, which are minded of their own freewill to go up to Jerusalem, go with thee.
EZRA|7|14|Forasmuch as thou art sent of the king, and of his seven counsellors, to enquire concerning Judah and Jerusalem, according to the law of thy God which is in thine hand;
EZRA|7|15|And to carry the silver and gold, which the king and his counsellors have freely offered unto the God of Israel, whose habitation is in Jerusalem,
EZRA|7|16|And all the silver and gold that thou canst find in all the province of Babylon, with the freewill offering of the people, and of the priests, offering willingly for the house of their God which is in Jerusalem:
EZRA|7|17|That thou mayest buy speedily with this money bullocks, rams, lambs, with their meat offerings and their drink offerings, and offer them upon the altar of the house of your God which is in Jerusalem.
EZRA|7|18|And whatsoever shall seem good to thee, and to thy brethren, to do with the rest of the silver and the gold, that do after the will of your God.
EZRA|7|19|The vessels also that are given thee for the service of the house of thy God, those deliver thou before the God of Jerusalem.
EZRA|7|20|And whatsoever more shall be needful for the house of thy God, which thou shalt have occasion to bestow, bestow it out of the king's treasure house.
EZRA|7|21|And I, even I Artaxerxes the king, do make a decree to all the treasurers which are beyond the river, that whatsoever Ezra the priest, the scribe of the law of the God of heaven, shall require of you, it be done speedily,
EZRA|7|22|Unto an hundred talents of silver, and to an hundred measures of wheat, and to an hundred baths of wine, and to an hundred baths of oil, and salt without prescribing how much.
EZRA|7|23|Whatsoever is commanded by the God of heaven, let it be diligently done for the house of the God of heaven: for why should there be wrath against the realm of the king and his sons?
EZRA|7|24|Also we certify you, that touching any of the priests and Levites, singers, porters, Nethinims, or ministers of this house of God, it shall not be lawful to impose toll, tribute, or custom, upon them.
EZRA|7|25|And thou, Ezra, after the wisdom of thy God, that is in thine hand, set magistrates and judges, which may judge all the people that are beyond the river, all such as know the laws of thy God; and teach ye them that know them not.
EZRA|7|26|And whosoever will not do the law of thy God, and the law of the king, let judgment be executed speedily upon him, whether it be unto death, or to banishment, or to confiscation of goods, or to imprisonment.
EZRA|7|27|Blessed be the LORD God of our fathers, which hath put such a thing as this in the king's heart, to beautify the house of the LORD which is in Jerusalem:
EZRA|7|28|And hath extended mercy unto me before the king, and his counsellors, and before all the king's mighty princes. And I was strengthened as the hand of the LORD my God was upon me, and I gathered together out of Israel chief men to go up with me.
EZRA|8|1|These are now the chief of their fathers, and this is the genealogy of them that went up with me from Babylon, in the reign of Artaxerxes the king.
EZRA|8|2|Of the sons of Phinehas; Gershom: of the sons of Ithamar; Daniel: of the sons of David; Hattush.
EZRA|8|3|Of the sons of Shechaniah, of the sons of Pharosh; Zechariah: and with him were reckoned by genealogy of the males an hundred and fifty.
EZRA|8|4|Of the sons of Pahathmoab; Elihoenai the son of Zerahiah, and with him two hundred males.
EZRA|8|5|Of the sons of Shechaniah; the son of Jahaziel, and with him three hundred males.
EZRA|8|6|Of the sons also of Adin; Ebed the son of Jonathan, and with him fifty males.
EZRA|8|7|And of the sons of Elam; Jeshaiah the son of Athaliah, and with him seventy males.
EZRA|8|8|And of the sons of Shephatiah; Zebadiah the son of Michael, and with him fourscore males.
EZRA|8|9|Of the sons of Joab; Obadiah the son of Jehiel, and with him two hundred and eighteen males.
EZRA|8|10|And of the sons of Shelomith; the son of Josiphiah, and with him an hundred and threescore males.
EZRA|8|11|And of the sons of Bebai; Zechariah the son of Bebai, and with him twenty and eight males.
EZRA|8|12|And of the sons of Azgad; Johanan the son of Hakkatan, and with him an hundred and ten males.
EZRA|8|13|And of the last sons of Adonikam, whose names are these, Eliphelet, Jeiel, and Shemaiah, and with them threescore males.
EZRA|8|14|Of the sons also of Bigvai; Uthai, and Zabbud, and with them seventy males.
EZRA|8|15|And I gathered them together to the river that runneth to Ahava; and there abode we in tents three days: and I viewed the people, and the priests, and found there none of the sons of Levi.
EZRA|8|16|Then sent I for Eliezer, for Ariel, for Shemaiah, and for Elnathan, and for Jarib, and for Elnathan, and for Nathan, and for Zechariah, and for Meshullam, chief men; also for Joiarib, and for Elnathan, men of understanding.
EZRA|8|17|And I sent them with commandment unto Iddo the chief at the place Casiphia, and I told them what they should say unto Iddo, and to his brethren the Nethinims, at the place Casiphia, that they should bring unto us ministers for the house of our God.
EZRA|8|18|And by the good hand of our God upon us they brought us a man of understanding, of the sons of Mahli, the son of Levi, the son of Israel; and Sherebiah, with his sons and his brethren, eighteen;
EZRA|8|19|And Hashabiah, and with him Jeshaiah of the sons of Merari, his brethren and their sons, twenty;
EZRA|8|20|Also of the Nethinims, whom David and the princes had appointed for the service of the Levites, two hundred and twenty Nethinims: all of them were expressed by name.
EZRA|8|21|Then I proclaimed a fast there, at the river of Ahava, that we might afflict ourselves before our God, to seek of him a right way for us, and for our little ones, and for all our substance.
EZRA|8|22|For I was ashamed to require of the king a band of soldiers and horsemen to help us against the enemy in the way: because we had spoken unto the king, saying, The hand of our God is upon all them for good that seek him; but his power and his wrath is against all them that forsake him.
EZRA|8|23|So we fasted and besought our God for this: and he was intreated of us.
EZRA|8|24|Then I separated twelve of the chief of the priests, Sherebiah, Hashabiah, and ten of their brethren with them,
EZRA|8|25|And weighed unto them the silver, and the gold, and the vessels, even the offering of the house of our God, which the king, and his counsellors, and his lords, and all Israel there present, had offered:
EZRA|8|26|I even weighed unto their hand six hundred and fifty talents of silver, and silver vessels an hundred talents, and of gold an hundred talents;
EZRA|8|27|Also twenty basons of gold, of a thousand drams; and two vessels of fine copper, precious as gold.
EZRA|8|28|And I said unto them, Ye are holy unto the LORD; the vessels are holy also; and the silver and the gold are a freewill offering unto the LORD God of your fathers.
EZRA|8|29|Watch ye, and keep them, until ye weigh them before the chief of the priests and the Levites, and chief of the fathers of Israel, at Jerusalem, in the chambers of the house of the LORD.
EZRA|8|30|So took the priests and the Levites the weight of the silver, and the gold, and the vessels, to bring them to Jerusalem unto the house of our God.
EZRA|8|31|Then we departed from the river of Ahava on the twelfth day of the first month, to go unto Jerusalem: and the hand of our God was upon us, and he delivered us from the hand of the enemy, and of such as lay in wait by the way.
EZRA|8|32|And we came to Jerusalem, and abode there three days.
EZRA|8|33|Now on the fourth day was the silver and the gold and the vessels weighed in the house of our God by the hand of Meremoth the son of Uriah the priest; and with him was Eleazar the son of Phinehas; and with them was Jozabad the son of Jeshua, and Noadiah the son of Binnui, Levites;
EZRA|8|34|By number and by weight of every one: and all the weight was written at that time.
EZRA|8|35|Also the children of those that had been carried away, which were come out of the captivity, offered burnt offerings unto the God of Israel, twelve bullocks for all Israel, ninety and six rams, seventy and seven lambs, twelve he goats for a sin offering: all this was a burnt offering unto the LORD.
EZRA|8|36|And they delivered the king's commissions unto the king's lieutenants, and to the governors on this side the river: and they furthered the people, and the house of God.
EZRA|9|1|Now when these things were done, the princes came to me, saying, The people of Israel, and the priests, and the Levites, have not separated themselves from the people of the lands, doing according to their abominations, even of the Canaanites, the Hittites, the Perizzites, the Jebusites, the Ammonites, the Moabites, the Egyptians, and the Amorites.
EZRA|9|2|For they have taken of their daughters for themselves, and for their sons: so that the holy seed have mingled themselves with the people of those lands: yea, the hand of the princes and rulers hath been chief in this trespass.
EZRA|9|3|And when I heard this thing, I rent my garment and my mantle, and plucked off the hair of my head and of my beard, and sat down astonied.
EZRA|9|4|Then were assembled unto me every one that trembled at the words of the God of Israel, because of the transgression of those that had been carried away; and I sat astonied until the evening sacrifice.
EZRA|9|5|And at the evening sacrifice I arose up from my heaviness; and having rent my garment and my mantle, I fell upon my knees, and spread out my hands unto the LORD my God,
EZRA|9|6|And said, O my God, I am ashamed and blush to lift up my face to thee, my God: for our iniquities are increased over our head, and our trespass is grown up unto the heavens.
EZRA|9|7|Since the days of our fathers have we been in a great trespass unto this day; and for our iniquities have we, our kings, and our priests, been delivered into the hand of the kings of the lands, to the sword, to captivity, and to a spoil, and to confusion of face, as it is this day.
EZRA|9|8|And now for a little space grace hath been shewed from the LORD our God, to leave us a remnant to escape, and to give us a nail in his holy place, that our God may lighten our eyes, and give us a little reviving in our bondage.
EZRA|9|9|For we were bondmen; yet our God hath not forsaken us in our bondage, but hath extended mercy unto us in the sight of the kings of Persia, to give us a reviving, to set up the house of our God, and to repair the desolations thereof, and to give us a wall in Judah and in Jerusalem.
EZRA|9|10|And now, O our God, what shall we say after this? for we have forsaken thy commandments,
EZRA|9|11|Which thou hast commanded by thy servants the prophets, saying, The land, unto which ye go to possess it, is an unclean land with the filthiness of the people of the lands, with their abominations, which have filled it from one end to another with their uncleanness.
EZRA|9|12|Now therefore give not your daughters unto their sons, neither take their daughters unto your sons, nor seek their peace or their wealth for ever: that ye may be strong, and eat the good of the land, and leave it for an inheritance to your children for ever.
EZRA|9|13|And after all that is come upon us for our evil deeds, and for our great trespass, seeing that thou our God hast punished us less than our iniquities deserve, and hast given us such deliverance as this;
EZRA|9|14|Should we again break thy commandments, and join in affinity with the people of these abominations? wouldest not thou be angry with us till thou hadst consumed us, so that there should be no remnant nor escaping?
EZRA|9|15|O LORD God of Israel, thou art righteous: for we remain yet escaped, as it is this day: behold, we are before thee in our trespasses: for we cannot stand before thee because of this.
EZRA|10|1|Now when Ezra had prayed, and when he had confessed, weeping and casting himself down before the house of God, there assembled unto him out of Israel a very great congregation of men and women and children: for the people wept very sore.
EZRA|10|2|And Shechaniah the son of Jehiel, one of the sons of Elam, answered and said unto Ezra, We have trespassed against our God, and have taken strange wives of the people of the land: yet now there is hope in Israel concerning this thing.
EZRA|10|3|Now therefore let us make a covenant with our God to put away all the wives, and such as are born of them, according to the counsel of my lord, and of those that tremble at the commandment of our God; and let it be done according to the law.
EZRA|10|4|Arise; for this matter belongeth unto thee: we also will be with thee: be of good courage, and do it.
EZRA|10|5|Then arose Ezra, and made the chief priests, the Levites, and all Israel, to swear that they should do according to this word. And they sware.
EZRA|10|6|Then Ezra rose up from before the house of God, and went into the chamber of Johanan the son of Eliashib: and when he came thither, he did eat no bread, nor drink water: for he mourned because of the transgression of them that had been carried away.
EZRA|10|7|And they made proclamation throughout Judah and Jerusalem unto all the children of the captivity, that they should gather themselves together unto Jerusalem;
EZRA|10|8|And that whosoever would not come within three days, according to the counsel of the princes and the elders, all his substance should be forfeited, and himself separated from the congregation of those that had been carried away.
EZRA|10|9|Then all the men of Judah and Benjamin gathered themselves together unto Jerusalem within three days. It was the ninth month, on the twentieth day of the month; and all the people sat in the street of the house of God, trembling because of this matter, and for the great rain.
EZRA|10|10|And Ezra the priest stood up, and said unto them, Ye have transgressed, and have taken strange wives, to increase the trespass of Israel.
EZRA|10|11|Now therefore make confession unto the LORD God of your fathers, and do his pleasure: and separate yourselves from the people of the land, and from the strange wives.
EZRA|10|12|Then all the congregation answered and said with a loud voice, As thou hast said, so must we do.
EZRA|10|13|But the people are many, and it is a time of much rain, and we are not able to stand without, neither is this a work of one day or two: for we are many that have transgressed in this thing.
EZRA|10|14|Let now our rulers of all the congregation stand, and let all them which have taken strange wives in our cities come at appointed times, and with them the elders of every city, and the judges thereof, until the fierce wrath of our God for this matter be turned from us.
EZRA|10|15|Only Jonathan the son of Asahel and Jahaziah the son of Tikvah were employed about this matter: and Meshullam and Shabbethai the Levite helped them.
EZRA|10|16|And the children of the captivity did so. And Ezra the priest, with certain chief of the fathers, after the house of their fathers, and all of them by their names, were separated, and sat down in the first day of the tenth month to examine the matter.
EZRA|10|17|And they made an end with all the men that had taken strange wives by the first day of the first month.
EZRA|10|18|And among the sons of the priests there were found that had taken strange wives: namely, of the sons of Jeshua the son of Jozadak, and his brethren; Maaseiah, and Eliezer, and Jarib, and Gedaliah.
EZRA|10|19|And they gave their hands that they would put away their wives; and being guilty, they offered a ram of the flock for their trespass.
EZRA|10|20|And of the sons of Immer; Hanani, and Zebadiah.
EZRA|10|21|And of the sons of Harim; Maaseiah, and Elijah, and Shemaiah, and Jehiel, and Uzziah.
EZRA|10|22|And of the sons of Pashur; Elioenai, Maaseiah, Ishmael, Nethaneel, Jozabad, and Elasah.
EZRA|10|23|Also of the Levites; Jozabad, and Shimei, and Kelaiah, (the same is Kelita,) Pethahiah, Judah, and Eliezer.
EZRA|10|24|Of the singers also; Eliashib: and of the porters; Shallum, and Telem, and Uri.
EZRA|10|25|Moreover of Israel: of the sons of Parosh; Ramiah, and Jeziah, and Malchiah, and Miamin, and Eleazar, and Malchijah, and Benaiah.
EZRA|10|26|And of the sons of Elam; Mattaniah, Zechariah, and Jehiel, and Abdi, and Jeremoth, and Eliah.
EZRA|10|27|And of the sons of Zattu; Elioenai, Eliashib, Mattaniah, and Jeremoth, and Zabad, and Aziza.
EZRA|10|28|Of the sons also of Bebai; Jehohanan, Hananiah, Zabbai, and Athlai.
EZRA|10|29|And of the sons of Bani; Meshullam, Malluch, and Adaiah, Jashub, and Sheal, and Ramoth.
EZRA|10|30|And of the sons of Pahathmoab; Adna, and Chelal, Benaiah, Maaseiah, Mattaniah, Bezaleel, and Binnui, and Manasseh.
EZRA|10|31|And of the sons of Harim; Eliezer, Ishijah, Malchiah, Shemaiah, Shimeon,
EZRA|10|32|Benjamin, Malluch, and Shemariah.
EZRA|10|33|Of the sons of Hashum; Mattenai, Mattathah, Zabad, Eliphelet, Jeremai, Manasseh, and Shimei.
EZRA|10|34|Of the sons of Bani; Maadai, Amram, and Uel,
EZRA|10|35|Benaiah, Bedeiah, Chelluh,
EZRA|10|36|Vaniah, Meremoth, Eliashib,
EZRA|10|37|Mattaniah, Mattenai, and Jaasau,
EZRA|10|38|And Bani, and Binnui, Shimei,
EZRA|10|39|And Shelemiah, and Nathan, and Adaiah,
EZRA|10|40|Machnadebai, Shashai, Sharai,
EZRA|10|41|Azareel, and Shelemiah, Shemariah,
EZRA|10|42|Shallum, Amariah, and Joseph.
EZRA|10|43|Of the sons of Nebo; Jeiel, Mattithiah, Zabad, Zebina, Jadau, and Joel, Benaiah.
EZRA|10|44|All these had taken strange wives: and some of them had wives by whom they had children.
