1CHR|1|1|Adam, Sheth, Enosh,
1CHR|1|2|Kenan, Mahalaleel, Jered,
1CHR|1|3|Henoch, Methuselah, Lamech,
1CHR|1|4|Noah, Shem, Ham, and Japheth.
1CHR|1|5|The sons of Japheth; Gomer, and Magog, and Madai, and Javan, and Tubal, and Meshech, and Tiras.
1CHR|1|6|And the sons of Gomer; Ashchenaz, and Riphath, and Togarmah.
1CHR|1|7|And the sons of Javan; Elishah, and Tarshish, Kittim, and Dodanim.
1CHR|1|8|The sons of Ham; Cush, and Mizraim, Put, and Canaan.
1CHR|1|9|And the sons of Cush; Seba, and Havilah, and Sabta, and Raamah, and Sabtecha. And the sons of Raamah; Sheba, and Dedan.
1CHR|1|10|And Cush begat Nimrod: he began to be mighty upon the earth.
1CHR|1|11|And Mizraim begat Ludim, and Anamim, and Lehabim, and Naphtuhim,
1CHR|1|12|And Pathrusim, and Casluhim, (of whom came the Philistines,) and Caphthorim.
1CHR|1|13|And Canaan begat Zidon his firstborn, and Heth,
1CHR|1|14|The Jebusite also, and the Amorite, and the Girgashite,
1CHR|1|15|And the Hivite, and the Arkite, and the Sinite,
1CHR|1|16|And the Arvadite, and the Zemarite, and the Hamathite.
1CHR|1|17|The sons of Shem; Elam, and Asshur, and Arphaxad, and Lud, and Aram, and Uz, and Hul, and Gether, and Meshech.
1CHR|1|18|And Arphaxad begat Shelah, and Shelah begat Eber.
1CHR|1|19|And unto Eber were born two sons: the name of the one was Peleg; because in his days the earth was divided: and his brother's name was Joktan.
1CHR|1|20|And Joktan begat Almodad, and Sheleph, and Hazarmaveth, and Jerah,
1CHR|1|21|Hadoram also, and Uzal, and Diklah,
1CHR|1|22|And Ebal, and Abimael, and Sheba,
1CHR|1|23|And Ophir, and Havilah, and Jobab. All these were the sons of Joktan.
1CHR|1|24|Shem, Arphaxad, Shelah,
1CHR|1|25|Eber, Peleg, Reu,
1CHR|1|26|Serug, Nahor, Terah,
1CHR|1|27|Abram; the same is Abraham.
1CHR|1|28|The sons of Abraham; Isaac, and Ishmael.
1CHR|1|29|These are their generations: The firstborn of Ishmael, Nebaioth; then Kedar, and Adbeel, and Mibsam,
1CHR|1|30|Mishma, and Dumah, Massa, Hadad, and Tema,
1CHR|1|31|Jetur, Naphish, and Kedemah. These are the sons of Ishmael.
1CHR|1|32|Now the sons of Keturah, Abraham's concubine: she bare Zimran, and Jokshan, and Medan, and Midian, and Ishbak, and Shuah. And the sons of Jokshan; Sheba, and Dedan.
1CHR|1|33|And the sons of Midian; Ephah, and Epher, and Henoch, and Abida, and Eldaah. All these are the sons of Keturah.
1CHR|1|34|And Abraham begat Isaac. The sons of Isaac; Esau and Israel.
1CHR|1|35|The sons of Esau; Eliphaz, Reuel, and Jeush, and Jaalam, and Korah.
1CHR|1|36|The sons of Eliphaz; Teman, and Omar, Zephi, and Gatam, Kenaz, and Timna, and Amalek.
1CHR|1|37|The sons of Reuel; Nahath, Zerah, Shammah, and Mizzah.
1CHR|1|38|And the sons of Seir; Lotan, and Shobal, and Zibeon, and Anah, and Dishon, and Ezar, and Dishan.
1CHR|1|39|And the sons of Lotan; Hori, and Homam: and Timna was Lotan's sister.
1CHR|1|40|The sons of Shobal; Alian, and Manahath, and Ebal, Shephi, and Onam. and the sons of Zibeon; Aiah, and Anah.
1CHR|1|41|The sons of Anah; Dishon. And the sons of Dishon; Amram, and Eshban, and Ithran, and Cheran.
1CHR|1|42|The sons of Ezer; Bilhan, and Zavan, and Jakan. The sons of Dishan; Uz, and Aran.
1CHR|1|43|Now these are the kings that reigned in the land of Edom before any king reigned over the children of Israel; Bela the son of Beor: and the name of his city was Dinhabah.
1CHR|1|44|And when Bela was dead, Jobab the son of Zerah of Bozrah reigned in his stead.
1CHR|1|45|And when Jobab was dead, Husham of the land of the Temanites reigned in his stead.
1CHR|1|46|And when Husham was dead, Hadad the son of Bedad, which smote Midian in the field of Moab, reigned in his stead: and the name of his city was Avith.
1CHR|1|47|And when Hadad was dead, Samlah of Masrekah reigned in his stead.
1CHR|1|48|And when Samlah was dead, Shaul of Rehoboth by the river reigned in his stead.
1CHR|1|49|And when Shaul was dead, Baalhanan the son of Achbor reigned in his stead.
1CHR|1|50|And when Baalhanan was dead, Hadad reigned in his stead: and the name of his city was Pai; and his wife's name was Mehetabel, the daughter of Matred, the daughter of Mezahab.
1CHR|1|51|Hadad died also. And the dukes of Edom were; duke Timnah, duke Aliah, duke Jetheth,
1CHR|1|52|Duke Aholibamah, duke Elah, duke Pinon,
1CHR|1|53|Duke Kenaz, duke Teman, duke Mibzar,
1CHR|1|54|Duke Magdiel, duke Iram. These are the dukes of Edom.
1CHR|2|1|These are the sons of Israel; Reuben, Simeon, Levi, and Judah, Issachar, and Zebulun,
1CHR|2|2|Dan, Joseph, and Benjamin, Naphtali, Gad, and Asher.
1CHR|2|3|The sons of Judah; Er, and Onan, and Shelah: which three were born unto him of the daughter of Shua the Canaanitess. And Er, the firstborn of Judah, was evil in the sight of the LORD; and he slew him.
1CHR|2|4|And Tamar his daughter in law bore him Pharez and Zerah. All the sons of Judah were five.
1CHR|2|5|The sons of Pharez; Hezron, and Hamul.
1CHR|2|6|And the sons of Zerah; Zimri, and Ethan, and Heman, and Calcol, and Dara: five of them in all.
1CHR|2|7|And the sons of Carmi; Achar, the troubler of Israel, who transgressed in the thing accursed.
1CHR|2|8|And the sons of Ethan; Azariah.
1CHR|2|9|The sons also of Hezron, that were born unto him; Jerahmeel, and Ram, and Chelubai.
1CHR|2|10|And Ram begat Amminadab; and Amminadab begat Nahshon, prince of the children of Judah;
1CHR|2|11|And Nahshon begat Salma, and Salma begat Boaz,
1CHR|2|12|And Boaz begat Obed, and Obed begat Jesse,
1CHR|2|13|And Jesse begat his firstborn Eliab, and Abinadab the second, and Shimma the third,
1CHR|2|14|Nethaneel the fourth, Raddai the fifth,
1CHR|2|15|Ozem the sixth, David the seventh:
1CHR|2|16|Whose sisters were Zeruiah, and Abigail. And the sons of Zeruiah; Abishai, and Joab, and Asahel, three.
1CHR|2|17|And Abigail bare Amasa: and the father of Amasa was Jether the Ishmeelite.
1CHR|2|18|And Caleb the son of Hezron begat children of Azubah his wife, and of Jerioth: her sons are these; Jesher, and Shobab, and Ardon.
1CHR|2|19|And when Azubah was dead, Caleb took unto him Ephrath, which bare him Hur.
1CHR|2|20|And Hur begat Uri, and Uri begat Bezaleel.
1CHR|2|21|And afterward Hezron went in to the daughter of Machir the father of Gilead, whom he married when he was threescore years old; and she bare him Segub.
1CHR|2|22|And Segub begat Jair, who had three and twenty cities in the land of Gilead.
1CHR|2|23|And he took Geshur, and Aram, with the towns of Jair, from them, with Kenath, and the towns thereof, even threescore cities. All these belonged to the sons of Machir the father of Gilead.
1CHR|2|24|And after that Hezron was dead in Calebephratah, then Abiah Hezron's wife bare him Ashur the father of Tekoa.
1CHR|2|25|And the sons of Jerahmeel the firstborn of Hezron were, Ram the firstborn, and Bunah, and Oren, and Ozem, and Ahijah.
1CHR|2|26|Jerahmeel had also another wife, whose name was Atarah; she was the mother of Onam.
1CHR|2|27|And the sons of Ram the firstborn of Jerahmeel were, Maaz, and Jamin, and Eker.
1CHR|2|28|And the sons of Onam were, Shammai, and Jada. And the sons of Shammai; Nadab and Abishur.
1CHR|2|29|And the name of the wife of Abishur was Abihail, and she bare him Ahban, and Molid.
1CHR|2|30|And the sons of Nadab; Seled, and Appaim: but Seled died without children.
1CHR|2|31|And the sons of Appaim; Ishi. And the sons of Ishi; Sheshan. And the children of Sheshan; Ahlai.
1CHR|2|32|And the sons of Jada the brother of Shammai; Jether, and Jonathan: and Jether died without children.
1CHR|2|33|And the sons of Jonathan; Peleth, and Zaza. These were the sons of Jerahmeel.
1CHR|2|34|Now Sheshan had no sons, but daughters. And Sheshan had a servant, an Egyptian, whose name was Jarha.
1CHR|2|35|And Sheshan gave his daughter to Jarha his servant to wife; and she bare him Attai.
1CHR|2|36|And Attai begat Nathan, and Nathan begat Zabad,
1CHR|2|37|And Zabad begat Ephlal, and Ephlal begat Obed,
1CHR|2|38|And Obed begat Jehu, and Jehu begat Azariah,
1CHR|2|39|And Azariah begat Helez, and Helez begat Eleasah,
1CHR|2|40|And Eleasah begat Sisamai, and Sisamai begat Shallum,
1CHR|2|41|And Shallum begat Jekamiah, and Jekamiah begat Elishama.
1CHR|2|42|Now the sons of Caleb the brother of Jerahmeel were, Mesha his firstborn, which was the father of Ziph; and the sons of Mareshah the father of Hebron.
1CHR|2|43|And the sons of Hebron; Korah, and Tappuah, and Rekem, and Shema.
1CHR|2|44|And Shema begat Raham, the father of Jorkoam: and Rekem begat Shammai.
1CHR|2|45|And the son of Shammai was Maon: and Maon was the father of Bethzur.
1CHR|2|46|And Ephah, Caleb's concubine, bare Haran, and Moza, and Gazez: and Haran begat Gazez.
1CHR|2|47|And the sons of Jahdai; Regem, and Jotham, and Gesham, and Pelet, and Ephah, and Shaaph.
1CHR|2|48|Maachah, Caleb's concubine, bare Sheber, and Tirhanah.
1CHR|2|49|She bare also Shaaph the father of Madmannah, Sheva the father of Machbenah, and the father of Gibea: and the daughter of Caleb was Achsa.
1CHR|2|50|These were the sons of Caleb the son of Hur, the firstborn of Ephratah; Shobal the father of Kirjathjearim.
1CHR|2|51|Salma the father of Bethlehem, Hareph the father of Bethgader.
1CHR|2|52|And Shobal the father of Kirjathjearim had sons; Haroeh, and half of the Manahethites.
1CHR|2|53|And the families of Kirjathjearim; the Ithrites, and the Puhites, and the Shumathites, and the Mishraites; of them came the Zareathites, and the Eshtaulites,
1CHR|2|54|The sons of Salma; Bethlehem, and the Netophathites, Ataroth, the house of Joab, and half of the Manahethites, the Zorites.
1CHR|2|55|And the families of the scribes which dwelt at Jabez; the Tirathites, the Shimeathites, and Suchathites. These are the Kenites that came of Hemath, the father of the house of Rechab.
1CHR|3|1|Now these were the sons of David, which were born unto him in Hebron; the firstborn Amnon, of Ahinoam the Jezreelitess; the second Daniel, of Abigail the Carmelitess:
1CHR|3|2|The third, Absalom the son of Maachah the daughter of Talmai king of Geshur: the fourth, Adonijah the son of Haggith:
1CHR|3|3|The fifth, Shephatiah of Abital: the sixth, Ithream by Eglah his wife.
1CHR|3|4|These six were born unto him in Hebron; and there he reigned seven years and six months: and in Jerusalem he reigned thirty and three years.
1CHR|3|5|And these were born unto him in Jerusalem; Shimea, and Shobab, and Nathan, and Solomon, four, of Bathshua the daughter of Ammiel:
1CHR|3|6|Ibhar also, and Elishama, and Eliphelet,
1CHR|3|7|And Nogah, and Nepheg, and Japhia,
1CHR|3|8|And Elishama, and Eliada, and Eliphelet, nine.
1CHR|3|9|These were all the sons of David, beside the sons of the concubines, and Tamar their sister.
1CHR|3|10|And Solomon's son was Rehoboam, Abia his son, Asa his son, Jehoshaphat his son,
1CHR|3|11|Joram his son, Ahaziah his son, Joash his son,
1CHR|3|12|Amaziah his son, Azariah his son, Jotham his son,
1CHR|3|13|Ahaz his son, Hezekiah his son, Manasseh his son,
1CHR|3|14|Amon his son, Josiah his son.
1CHR|3|15|And the sons of Josiah were, the firstborn Johanan, the second Jehoiakim, the third Zedekiah, the fourth Shallum.
1CHR|3|16|And the sons of Jehoiakim: Jeconiah his son, Zedekiah his son.
1CHR|3|17|And the sons of Jeconiah; Assir, Salathiel his son,
1CHR|3|18|Malchiram also, and Pedaiah, and Shenazar, Jecamiah, Hoshama, and Nedabiah.
1CHR|3|19|And the sons of Pedaiah were, Zerubbabel, and Shimei: and the sons of Zerubbabel; Meshullam, and Hananiah, and Shelomith their sister:
1CHR|3|20|And Hashubah, and Ohel, and Berechiah, and Hasadiah, Jushabhesed, five.
1CHR|3|21|And the sons of Hananiah; Pelatiah, and Jesaiah: the sons of Rephaiah, the sons of Arnan, the sons of Obadiah, the sons of Shechaniah.
1CHR|3|22|And the sons of Shechaniah; Shemaiah: and the sons of Shemaiah; Hattush, and Igeal, and Bariah, and Neariah, and Shaphat, six.
1CHR|3|23|And the sons of Neariah; Elioenai, and Hezekiah, and Azrikam, three.
1CHR|3|24|And the sons of Elioenai were, Hodaiah, and Eliashib, and Pelaiah, and Akkub, and Johanan, and Dalaiah, and Anani, seven.
1CHR|4|1|The sons of Judah; Pharez, Hezron, and Carmi, and Hur, and Shobal.
1CHR|4|2|And Reaiah the son of Shobal begat Jahath; and Jahath begat Ahumai, and Lahad. These are the families of the Zorathites.
1CHR|4|3|And these were of the father of Etam; Jezreel, and Ishma, and Idbash: and the name of their sister was Hazelelponi:
1CHR|4|4|And Penuel the father of Gedor, and Ezer the father of Hushah. These are the sons of Hur, the firstborn of Ephratah, the father of Bethlehem.
1CHR|4|5|And Ashur the father of Tekoa had two wives, Helah and Naarah.
1CHR|4|6|And Naarah bare him Ahuzam, and Hepher, and Temeni, and Haahashtari. These were the sons of Naarah.
1CHR|4|7|And the sons of Helah were, Zereth, and Jezoar, and Ethnan.
1CHR|4|8|And Coz begat Anub, and Zobebah, and the families of Aharhel the son of Harum.
1CHR|4|9|And Jabez was more honorable than his brethren: and his mother called his name Jabez, saying, Because I bare him with sorrow.
1CHR|4|10|And Jabez called on the God of Israel, saying, Oh that thou wouldest bless me indeed, and enlarge my coast, and that thine hand might be with me, and that thou wouldest keep me from evil, that it may not grieve me! And God granted him that which he requested.
1CHR|4|11|And Chelub the brother of Shuah begat Mehir, which was the father of Eshton.
1CHR|4|12|And Eshton begat Bethrapha, and Paseah, and Tehinnah the father of Irnahash. These are the men of Rechah.
1CHR|4|13|And the sons of Kenaz; Othniel, and Seraiah: and the sons of Othniel; Hathath.
1CHR|4|14|And Meonothai begat Ophrah: and Seraiah begat Joab, the father of the valley of Charashim; for they were craftsmen.
1CHR|4|15|And the sons of Caleb the son of Jephunneh; Iru, Elah, and Naam: and the sons of Elah, even Kenaz.
1CHR|4|16|And the sons of Jehaleleel; Ziph, and Ziphah, Tiria, and Asareel.
1CHR|4|17|And the sons of Ezra were, Jether, and Mered, and Epher, and Jalon: and she bare Miriam, and Shammai, and Ishbah the father of Eshtemoa.
1CHR|4|18|And his wife Jehudijah bare Jered the father of Gedor, and Heber the father of Socho, and Jekuthiel the father of Zanoah. And these are the sons of Bithiah the daughter of Pharaoh, which Mered took.
1CHR|4|19|And the sons of his wife Hodiah the sister of Naham, the father of Keilah the Garmite, and Eshtemoa the Maachathite.
1CHR|4|20|And the sons of Shimon were, Amnon, and Rinnah, Benhanan, and Tilon. And the sons of Ishi were, Zoheth, and Benzoheth.
1CHR|4|21|The sons of Shelah the son of Judah were, Er the father of Lecah, and Laadah the father of Mareshah, and the families of the house of them that wrought fine linen, of the house of Ashbea,
1CHR|4|22|And Jokim, and the men of Chozeba, and Joash, and Saraph, who had the dominion in Moab, and Jashubilehem. And these are ancient things.
1CHR|4|23|These were the potters, and those that dwelt among plants and hedges: there they dwelt with the king for his work.
1CHR|4|24|The sons of Simeon were, Nemuel, and Jamin, Jarib, Zerah, and Shaul:
1CHR|4|25|Shallum his son, Mibsam his son, Mishma his son.
1CHR|4|26|And the sons of Mishma; Hamuel his son, Zacchur his son, Shimei his son.
1CHR|4|27|And Shimei had sixteen sons and six daughters: but his brethren had not many children, neither did all their family multiply, like to the children of Judah.
1CHR|4|28|And they dwelt at Beersheba, and Moladah, and Hazarshual,
1CHR|4|29|And at Bilhah, and at Ezem, and at Tolad,
1CHR|4|30|And at Bethuel, and at Hormah, and at Ziklag,
1CHR|4|31|And at Bethmarcaboth, and Hazarsusim, and at Bethbirei, and at Shaaraim. These were their cities unto the reign of David.
1CHR|4|32|And their villages were, Etam, and Ain, Rimmon, and Tochen, and Ashan, five cities:
1CHR|4|33|And all their villages that were round about the same cities, unto Baal. These were their habitations, and their genealogy.
1CHR|4|34|And Meshobab, and Jamlech, and Joshah, the son of Amaziah,
1CHR|4|35|And Joel, and Jehu the son of Josibiah, the son of Seraiah, the son of Asiel,
1CHR|4|36|And Elioenai, and Jaakobah, and Jeshohaiah, and Asaiah, and Adiel, and Jesimiel, and Benaiah,
1CHR|4|37|And Ziza the son of Shiphi, the son of Allon, the son of Jedaiah, the son of Shimri, the son of Shemaiah;
1CHR|4|38|These mentioned by their names were princes in their families: and the house of their fathers increased greatly.
1CHR|4|39|And they went to the entrance of Gedor, even unto the east side of the valley, to seek pasture for their flocks.
1CHR|4|40|And they found fat pasture and good, and the land was wide, and quiet, and peaceable; for they of Ham had dwelt there of old.
1CHR|4|41|And these written by name came in the days of Hezekiah king of Judah, and smote their tents, and the habitations that were found there, and destroyed them utterly unto this day, and dwelt in their rooms: because there was pasture there for their flocks.
1CHR|4|42|And some of them, even of the sons of Simeon, five hundred men, went to mount Seir, having for their captains Pelatiah, and Neariah, and Rephaiah, and Uzziel, the sons of Ishi.
1CHR|4|43|And they smote the rest of the Amalekites that were escaped, and dwelt there unto this day.
1CHR|5|1|Now the sons of Reuben the firstborn of Israel, (for he was the firstborn; but forasmuch as he defiled his father's bed, his birthright was given unto the sons of Joseph the son of Israel: and the genealogy is not to be reckoned after the birthright.
1CHR|5|2|For Judah prevailed above his brethren, and of him came the chief ruler; but the birthright was Joseph's:)
1CHR|5|3|The sons, I say, of Reuben the firstborn of Israel were, Hanoch, and Pallu, Hezron, and Carmi.
1CHR|5|4|The sons of Joel; Shemaiah his son, Gog his son, Shimei his son,
1CHR|5|5|Micah his son, Reaia his son, Baal his son,
1CHR|5|6|Beerah his son, whom Tilgathpilneser king of Assyria carried away captive: he was prince of the Reubenites.
1CHR|5|7|And his brethren by their families, when the genealogy of their generations was reckoned, were the chief, Jeiel, and Zechariah,
1CHR|5|8|And Bela the son of Azaz, the son of Shema, the son of Joel, who dwelt in Aroer, even unto Nebo and Baalmeon:
1CHR|5|9|And eastward he inhabited unto the entering in of the wilderness from the river Euphrates: because their cattle were multiplied in the land of Gilead.
1CHR|5|10|And in the days of Saul they made war with the Hagarites, who fell by their hand: and they dwelt in their tents throughout all the east land of Gilead.
1CHR|5|11|And the children of Gad dwelt over against them, in the land of Bashan unto Salcah:
1CHR|5|12|Joel the chief, and Shapham the next, and Jaanai, and Shaphat in Bashan.
1CHR|5|13|And their brethren of the house of their fathers were, Michael, and Meshullam, and Sheba, and Jorai, and Jachan, and Zia, and Heber, seven.
1CHR|5|14|These are the children of Abihail the son of Huri, the son of Jaroah, the son of Gilead, the son of Michael, the son of Jeshishai, the son of Jahdo, the son of Buz;
1CHR|5|15|Ahi the son of Abdiel, the son of Guni, chief of the house of their fathers.
1CHR|5|16|And they dwelt in Gilead in Bashan, and in her towns, and in all the suburbs of Sharon, upon their borders.
1CHR|5|17|All these were reckoned by genealogies in the days of Jotham king of Judah, and in the days of Jeroboam king of Israel.
1CHR|5|18|The sons of Reuben, and the Gadites, and half the tribe of Manasseh, of valiant men, men able to bear buckler and sword, and to shoot with bow, and skillful in war, were four and forty thousand seven hundred and threescore, that went out to the war.
1CHR|5|19|And they made war with the Hagarites, with Jetur, and Nephish, and Nodab.
1CHR|5|20|And they were helped against them, and the Hagarites were delivered into their hand, and all that were with them: for they cried to God in the battle, and he was intreated of them; because they put their trust in him.
1CHR|5|21|And they took away their cattle; of their camels fifty thousand, and of sheep two hundred and fifty thousand, and of asses two thousand, and of men an hundred thousand.
1CHR|5|22|For there fell down many slain, because the war was of God. And they dwelt in their steads until the captivity.
1CHR|5|23|And the children of the half tribe of Manasseh dwelt in the land: they increased from Bashan unto Baalhermon and Senir, and unto mount Hermon.
1CHR|5|24|And these were the heads of the house of their fathers, even Epher, and Ishi, and Eliel, and Azriel, and Jeremiah, and Hodaviah, and Jahdiel, mighty men of valor, famous men, and heads of the house of their fathers.
1CHR|5|25|And they transgressed against the God of their fathers, and went a whoring after the gods of the people of the land, whom God destroyed before them.
1CHR|5|26|And the God of Israel stirred up the spirit of Pul king of Assyria, and the spirit of Tilgathpilneser king of Assyria, and he carried them away, even the Reubenites, and the Gadites, and the half tribe of Manasseh, and brought them unto Halah, and Habor, and Hara, and to the river Gozan, unto this day.
1CHR|6|1|The sons of Levi; Gershon, Kohath, and Merari.
1CHR|6|2|And the sons of Kohath; Amram, Izhar, and Hebron, and Uzziel.
1CHR|6|3|And the children of Amram; Aaron, and Moses, and Miriam. The sons also of Aaron; Nadab, and Abihu, Eleazar, and Ithamar.
1CHR|6|4|Eleazar begat Phinehas, Phinehas begat Abishua,
1CHR|6|5|And Abishua begat Bukki, and Bukki begat Uzzi,
1CHR|6|6|And Uzzi begat Zerahiah, and Zerahiah begat Meraioth,
1CHR|6|7|Meraioth begat Amariah, and Amariah begat Ahitub,
1CHR|6|8|And Ahitub begat Zadok, and Zadok begat Ahimaaz,
1CHR|6|9|And Ahimaaz begat Azariah, and Azariah begat Johanan,
1CHR|6|10|And Johanan begat Azariah, (he it is that executed the priest's office in the temple that Solomon built in Jerusalem:)
1CHR|6|11|And Azariah begat Amariah, and Amariah begat Ahitub,
1CHR|6|12|And Ahitub begat Zadok, and Zadok begat Shallum,
1CHR|6|13|And Shallum begat Hilkiah, and Hilkiah begat Azariah,
1CHR|6|14|And Azariah begat Seraiah, and Seraiah begat Jehozadak,
1CHR|6|15|And Jehozadak went into captivity, when the LORD carried away Judah and Jerusalem by the hand of Nebuchadnezzar.
1CHR|6|16|The sons of Levi; Gershom, Kohath, and Merari.
1CHR|6|17|And these be the names of the sons of Gershom; Libni, and Shimei.
1CHR|6|18|And the sons of Kohath were, Amram, and Izhar, and Hebron, and Uzziel.
1CHR|6|19|The sons of Merari; Mahli, and Mushi. And these are the families of the Levites according to their fathers.
1CHR|6|20|Of Gershom; Libni his son, Jahath his son, Zimmah his son,
1CHR|6|21|Joah his son, Iddo his son, Zerah his son, Jeaterai his son.
1CHR|6|22|The sons of Kohath; Amminadab his son, Korah his son, Assir his son,
1CHR|6|23|Elkanah his son, and Ebiasaph his son, and Assir his son,
1CHR|6|24|Tahath his son, Uriel his son, Uzziah his son, and Shaul his son.
1CHR|6|25|And the sons of Elkanah; Amasai, and Ahimoth.
1CHR|6|26|As for Elkanah: the sons of Elkanah; Zophai his son, and Nahath his son,
1CHR|6|27|Eliab his son, Jeroham his son, Elkanah his son.
1CHR|6|28|And the sons of Samuel; the firstborn Vashni, and Abiah.
1CHR|6|29|The sons of Merari; Mahli, Libni his son, Shimei his son, Uzza his son,
1CHR|6|30|Shimea his son, Haggiah his son, Asaiah his son.
1CHR|6|31|And these are they whom David set over the service of song in the house of the LORD, after that the ark had rest.
1CHR|6|32|And they ministered before the dwelling place of the tabernacle of the congregation with singing, until Solomon had built the house of the LORD in Jerusalem: and then they waited on their office according to their order.
1CHR|6|33|And these are they that waited with their children. Of the sons of the Kohathites: Heman a singer, the son of Joel, the son of Shemuel,
1CHR|6|34|The son of Elkanah, the son of Jeroham, the son of Eliel, the son of Toah,
1CHR|6|35|The son of Zuph, the son of Elkanah, the son of Mahath, the son of Amasai,
1CHR|6|36|The son of Elkanah, the son of Joel, the son of Azariah, the son of Zephaniah,
1CHR|6|37|The son of Tahath, the son of Assir, the son of Ebiasaph, the son of Korah,
1CHR|6|38|The son of Izhar, the son of Kohath, the son of Levi, the son of Israel.
1CHR|6|39|And his brother Asaph, who stood on his right hand, even Asaph the son of Berachiah, the son of Shimea,
1CHR|6|40|The son of Michael, the son of Baaseiah, the son of Malchiah,
1CHR|6|41|The son of Ethni, the son of Zerah, the son of Adaiah,
1CHR|6|42|The son of Ethan, the son of Zimmah, the son of Shimei,
1CHR|6|43|The son of Jahath, the son of Gershom, the son of Levi.
1CHR|6|44|And their brethren the sons of Merari stood on the left hand: Ethan the son of Kishi, the son of Abdi, the son of Malluch,
1CHR|6|45|The son of Hashabiah, the son of Amaziah, the son of Hilkiah,
1CHR|6|46|The son of Amzi, the son of Bani, the son of Shamer,
1CHR|6|47|The son of Mahli, the son of Mushi, the son of Merari, the son of Levi.
1CHR|6|48|Their brethren also the Levites were appointed unto all manner of service of the tabernacle of the house of God.
1CHR|6|49|But Aaron and his sons offered upon the altar of the burnt offering, and on the altar of incense, and were appointed for all the work of the place most holy, and to make an atonement for Israel, according to all that Moses the servant of God had commanded.
1CHR|6|50|And these are the sons of Aaron; Eleazar his son, Phinehas his son, Abishua his son,
1CHR|6|51|Bukki his son, Uzzi his son, Zerahiah his son,
1CHR|6|52|Meraioth his son, Amariah his son, Ahitub his son,
1CHR|6|53|Zadok his son, Ahimaaz his son.
1CHR|6|54|Now these are their dwelling places throughout their castles in their coasts, of the sons of Aaron, of the families of the Kohathites: for theirs was the lot.
1CHR|6|55|And they gave them Hebron in the land of Judah, and the suburbs thereof round about it.
1CHR|6|56|But the fields of the city, and the villages thereof, they gave to Caleb the son of Jephunneh.
1CHR|6|57|And to the sons of Aaron they gave the cities of Judah, namely, Hebron, the city of refuge, and Libnah with her suburbs, and Jattir, and Eshtemoa, with their suburbs,
1CHR|6|58|And Hilen with her suburbs, Debir with her suburbs,
1CHR|6|59|And Ashan with her suburbs, and Bethshemesh with her suburbs:
1CHR|6|60|And out of the tribe of Benjamin; Geba with her suburbs, and Alemeth with her suburbs, and Anathoth with her suburbs. All their cities throughout their families were thirteen cities.
1CHR|6|61|And unto the sons of Kohath, which were left of the family of that tribe, were cities given out of the half tribe, namely, out of the half tribe of Manasseh, by lot, ten cities.
1CHR|6|62|And to the sons of Gershom throughout their families out of the tribe of Issachar, and out of the tribe of Asher, and out of the tribe of Naphtali, and out of the tribe of Manasseh in Bashan, thirteen cities.
1CHR|6|63|Unto the sons of Merari were given by lot, throughout their families, out of the tribe of Reuben, and out of the tribe of Gad, and out of the tribe of Zebulun, twelve cities.
1CHR|6|64|And the children of Israel gave to the Levites these cities with their suburbs.
1CHR|6|65|And they gave by lot out of the tribe of the children of Judah, and out of the tribe of the children of Simeon, and out of the tribe of the children of Benjamin, these cities, which are called by their names.
1CHR|6|66|And the residue of the families of the sons of Kohath had cities of their coasts out of the tribe of Ephraim.
1CHR|6|67|And they gave unto them, of the cities of refuge, Shechem in mount Ephraim with her suburbs; they gave also Gezer with her suburbs,
1CHR|6|68|And Jokmeam with her suburbs, and Bethhoron with her suburbs,
1CHR|6|69|And Aijalon with her suburbs, and Gathrimmon with her suburbs:
1CHR|6|70|And out of the half tribe of Manasseh; Aner with her suburbs, and Bileam with her suburbs, for the family of the remnant of the sons of Kohath.
1CHR|6|71|Unto the sons of Gershom were given out of the family of the half tribe of Manasseh, Golan in Bashan with her suburbs, and Ashtaroth with her suburbs:
1CHR|6|72|And out of the tribe of Issachar; Kedesh with her suburbs, Daberath with her suburbs,
1CHR|6|73|And Ramoth with her suburbs, and Anem with her suburbs:
1CHR|6|74|And out of the tribe of Asher; Mashal with her suburbs, and Abdon with her suburbs,
1CHR|6|75|And Hukok with her suburbs, and Rehob with her suburbs:
1CHR|6|76|And out of the tribe of Naphtali; Kedesh in Galilee with her suburbs, and Hammon with her suburbs, and Kirjathaim with her suburbs.
1CHR|6|77|Unto the rest of the children of Merari were given out of the tribe of Zebulun, Rimmon with her suburbs, Tabor with her suburbs:
1CHR|6|78|And on the other side Jordan by Jericho, on the east side of Jordan, were given them out of the tribe of Reuben, Bezer in the wilderness with her suburbs, and Jahzah with her suburbs,
1CHR|6|79|Kedemoth also with her suburbs, and Mephaath with her suburbs:
1CHR|6|80|And out of the tribe of Gad; Ramoth in Gilead with her suburbs, and Mahanaim with her suburbs,
1CHR|6|81|And Heshbon with her suburbs, and Jazer with her suburbs.
1CHR|7|1|Now the sons of Issachar were, Tola, and Puah, Jashub, and Shimrom, four.
1CHR|7|2|And the sons of Tola; Uzzi, and Rephaiah, and Jeriel, and Jahmai, and Jibsam, and Shemuel, heads of their father's house, to wit, of Tola: they were valiant men of might in their generations; whose number was in the days of David two and twenty thousand and six hundred.
1CHR|7|3|And the sons of Uzzi; Izrahiah: and the sons of Izrahiah; Michael, and Obadiah, and Joel, Ishiah, five: all of them chief men.
1CHR|7|4|And with them, by their generations, after the house of their fathers, were bands of soldiers for war, six and thirty thousand men: for they had many wives and sons.
1CHR|7|5|And their brethren among all the families of Issachar were valiant men of might, reckoned in all by their genealogies fourscore and seven thousand.
1CHR|7|6|The sons of Benjamin; Bela, and Becher, and Jediael, three.
1CHR|7|7|And the sons of Bela; Ezbon, and Uzzi, and Uzziel, and Jerimoth, and Iri, five; heads of the house of their fathers, mighty men of valor; and were reckoned by their genealogies twenty and two thousand and thirty and four.
1CHR|7|8|And the sons of Becher; Zemira, and Joash, and Eliezer, and Elioenai, and Omri, and Jerimoth, and Abiah, and Anathoth, and Alameth. All these are the sons of Becher.
1CHR|7|9|And the number of them, after their genealogy by their generations, heads of the house of their fathers, mighty men of valor, was twenty thousand and two hundred.
1CHR|7|10|The sons also of Jediael; Bilhan: and the sons of Bilhan; Jeush, and Benjamin, and Ehud, and Chenaanah, and Zethan, and Tharshish, and Ahishahar.
1CHR|7|11|All these the sons of Jediael, by the heads of their fathers, mighty men of valor, were seventeen thousand and two hundred soldiers, fit to go out for war and battle.
1CHR|7|12|Shuppim also, and Huppim, the children of Ir, and Hushim, the sons of Aher.
1CHR|7|13|The sons of Naphtali; Jahziel, and Guni, and Jezer, and Shallum, the sons of Bilhah.
1CHR|7|14|The sons of Manasseh; Ashriel, whom she bare: (but his concubine the Aramitess bare Machir the father of Gilead:
1CHR|7|15|And Machir took to wife the sister of Huppim and Shuppim, whose sister's name was Maachah;) and the name of the second was Zelophehad: and Zelophehad had daughters.
1CHR|7|16|And Maachah the wife of Machir bare a son, and she called his name Peresh; and the name of his brother was Sheresh; and his sons were Ulam and Rakem.
1CHR|7|17|And the sons of Ulam; Bedan. These were the sons of Gilead, the son of Machir, the son of Manasseh.
1CHR|7|18|And his sister Hammoleketh bare Ishod, and Abiezer, and Mahalah.
1CHR|7|19|And the sons of Shemidah were, Ahian, and Shechem, and Likhi, and Aniam.
1CHR|7|20|And the sons of Ephraim; Shuthelah, and Bered his son, and Tahath his son, and Eladah his son, and Tahath his son,
1CHR|7|21|And Zabad his son, and Shuthelah his son, and Ezer, and Elead, whom the men of Gath that were born in that land slew, because they came down to take away their cattle.
1CHR|7|22|And Ephraim their father mourned many days, and his brethren came to comfort him.
1CHR|7|23|And when he went in to his wife, she conceived, and bare a son, and he called his name Beriah, because it went evil with his house.
1CHR|7|24|(And his daughter was Sherah, who built Bethhoron the nether, and the upper, and Uzzensherah.)
1CHR|7|25|And Rephah was his son, also Resheph, and Telah his son, and Tahan his son.
1CHR|7|26|Laadan his son, Ammihud his son, Elishama his son.
1CHR|7|27|Non his son, Jehoshuah his son.
1CHR|7|28|And their possessions and habitations were, Bethel and the towns thereof, and eastward Naaran, and westward Gezer, with the towns thereof; Shechem also and the towns thereof, unto Gaza and the towns thereof:
1CHR|7|29|And by the borders of the children of Manasseh, Bethshean and her towns, Taanach and her towns, Megiddo and her towns, Dor and her towns. In these dwelt the children of Joseph the son of Israel.
1CHR|7|30|The sons of Asher; Imnah, and Isuah, and Ishuai, and Beriah, and Serah their sister.
1CHR|7|31|And the sons of Beriah; Heber, and Malchiel, who is the father of Birzavith.
1CHR|7|32|And Heber begat Japhlet, and Shomer, and Hotham, and Shua their sister.
1CHR|7|33|And the sons of Japhlet; Pasach, and Bimhal, and Ashvath. These are the children of Japhlet.
1CHR|7|34|And the sons of Shamer; Ahi, and Rohgah, Jehubbah, and Aram.
1CHR|7|35|And the sons of his brother Helem; Zophah, and Imna, and Shelesh, and Amal.
1CHR|7|36|The sons of Zophah; Suah, and Harnepher, and Shual, and Beri, and Imrah,
1CHR|7|37|Bezer, and Hod, and Shamma, and Shilshah, and Ithran, and Beera.
1CHR|7|38|And the sons of Jether; Jephunneh, and Pispah, and Ara.
1CHR|7|39|And the sons of Ulla; Arah, and Haniel, and Rezia.
1CHR|7|40|All these were the children of Asher, heads of their father's house, choice and mighty men of valor, chief of the princes. And the number throughout the genealogy of them that were apt to the war and to battle was twenty and six thousand men.
1CHR|8|1|Now Benjamin begat Bela his firstborn, Ashbel the second, and Aharah the third,
1CHR|8|2|Nohah the fourth, and Rapha the fifth.
1CHR|8|3|And the sons of Bela were, Addar, and Gera, and Abihud,
1CHR|8|4|And Abishua, and Naaman, and Ahoah,
1CHR|8|5|And Gera, and Shephuphan, and Huram.
1CHR|8|6|And these are the sons of Ehud: these are the heads of the fathers of the inhabitants of Geba, and they removed them to Manahath:
1CHR|8|7|And Naaman, and Ahiah, and Gera, he removed them, and begat Uzza, and Ahihud.
1CHR|8|8|And Shaharaim begat children in the country of Moab, after he had sent them away; Hushim and Baara were his wives.
1CHR|8|9|And he begat of Hodesh his wife, Jobab, and Zibia, and Mesha, and Malcham,
1CHR|8|10|And Jeuz, and Shachia, and Mirma. These were his sons, heads of the fathers.
1CHR|8|11|And of Hushim he begat Abitub, and Elpaal.
1CHR|8|12|The sons of Elpaal; Eber, and Misham, and Shamed, who built Ono, and Lod, with the towns thereof:
1CHR|8|13|Beriah also, and Shema, who were heads of the fathers of the inhabitants of Aijalon, who drove away the inhabitants of Gath:
1CHR|8|14|And Ahio, Shashak, and Jeremoth,
1CHR|8|15|And Zebadiah, and Arad, and Ader,
1CHR|8|16|And Michael, and Ispah, and Joha, the sons of Beriah;
1CHR|8|17|And Zebadiah, and Meshullam, and Hezeki, and Heber,
1CHR|8|18|Ishmerai also, and Jezliah, and Jobab, the sons of Elpaal;
1CHR|8|19|And Jakim, and Zichri, and Zabdi,
1CHR|8|20|And Elienai, and Zilthai, and Eliel,
1CHR|8|21|And Adaiah, and Beraiah, and Shimrath, the sons of Shimhi;
1CHR|8|22|And Ishpan, and Heber, and Eliel,
1CHR|8|23|And Abdon, and Zichri, and Hanan,
1CHR|8|24|And Hananiah, and Elam, and Antothijah,
1CHR|8|25|And Iphedeiah, and Penuel, the sons of Shashak;
1CHR|8|26|And Shamsherai, and Shehariah, and Athaliah,
1CHR|8|27|And Jaresiah, and Eliah, and Zichri, the sons of Jeroham.
1CHR|8|28|These were heads of the fathers, by their generations, chief men. These dwelt in Jerusalem.
1CHR|8|29|And at Gibeon dwelt the father of Gibeon; whose wife's name was Maachah:
1CHR|8|30|And his firstborn son Abdon, and Zur, and Kish, and Baal, and Nadab,
1CHR|8|31|And Gedor, and Ahio, and Zacher.
1CHR|8|32|And Mikloth begat Shimeah. And these also dwelt with their brethren in Jerusalem, over against them.
1CHR|8|33|And Ner begat Kish, and Kish begat Saul, and Saul begat Jonathan, and Malchishua, and Abinadab, and Eshbaal.
1CHR|8|34|And the son of Jonathan was Meribbaal; and Meribbaal begat Micah.
1CHR|8|35|And the sons of Micah were, Pithon, and Melech, and Tarea, and Ahaz.
1CHR|8|36|And Ahaz begat Jehoadah; and Jehoadah begat Alemeth, and Azmaveth, and Zimri; and Zimri begat Moza,
1CHR|8|37|And Moza begat Binea: Rapha was his son, Eleasah his son, Azel his son:
1CHR|8|38|And Azel had six sons, whose names are these, Azrikam, Bocheru, and Ishmael, and Sheariah, and Obadiah, and Hanan. All these were the sons of Azel.
1CHR|8|39|And the sons of Eshek his brother were, Ulam his firstborn, Jehush the second, and Eliphelet the third.
1CHR|8|40|And the sons of Ulam were mighty men of valor, archers, and had many sons, and sons' sons, an hundred and fifty. All these are of the sons of Benjamin.
1CHR|9|1|So all Israel were reckoned by genealogies; and, behold, they were written in the book of the kings of Israel and Judah, who were carried away to Babylon for their transgression.
1CHR|9|2|Now the first inhabitants that dwelt in their possessions in their cities were, the Israelites, the priests, Levites, and the Nethinims.
1CHR|9|3|And in Jerusalem dwelt of the children of Judah, and of the children of Benjamin, and of the children of Ephraim, and Manasseh;
1CHR|9|4|Uthai the son of Ammihud, the son of Omri, the son of Imri, the son of Bani, of the children of Pharez the son of Judah.
1CHR|9|5|And of the Shilonites; Asaiah the firstborn, and his sons.
1CHR|9|6|And of the sons of Zerah; Jeuel, and their brethren, six hundred and ninety.
1CHR|9|7|And of the sons of Benjamin; Sallu the son of Meshullam, the son of Hodaviah, the son of Hasenuah,
1CHR|9|8|And Ibneiah the son of Jeroham, and Elah the son of Uzzi, the son of Michri, and Meshullam the son of Shephathiah, the son of Reuel, the son of Ibnijah;
1CHR|9|9|And their brethren, according to their generations, nine hundred and fifty and six. All these men were chief of the fathers in the house of their fathers.
1CHR|9|10|And of the priests; Jedaiah, and Jehoiarib, and Jachin,
1CHR|9|11|And Azariah the son of Hilkiah, the son of Meshullam, the son of Zadok, the son of Meraioth, the son of Ahitub, the ruler of the house of God;
1CHR|9|12|And Adaiah the son of Jeroham, the son of Pashur, the son of Malchijah, and Maasiai the son of Adiel, the son of Jahzerah, the son of Meshullam, the son of Meshillemith, the son of Immer;
1CHR|9|13|And their brethren, heads of the house of their fathers, a thousand and seven hundred and threescore; very able men for the work of the service of the house of God.
1CHR|9|14|And of the Levites; Shemaiah the son of Hasshub, the son of Azrikam, the son of Hashabiah, of the sons of Merari;
1CHR|9|15|And Bakbakkar, Heresh, and Galal, and Mattaniah the son of Micah, the son of Zichri, the son of Asaph;
1CHR|9|16|And Obadiah the son of Shemaiah, the son of Galal, the son of Jeduthun, and Berechiah the son of Asa, the son of Elkanah, that dwelt in the villages of the Netophathites.
1CHR|9|17|And the porters were, Shallum, and Akkub, and Talmon, and Ahiman, and their brethren: Shallum was the chief;
1CHR|9|18|Who hitherto waited in the king's gate eastward: they were porters in the companies of the children of Levi.
1CHR|9|19|And Shallum the son of Kore, the son of Ebiasaph, the son of Korah, and his brethren, of the house of his father, the Korahites, were over the work of the service, keepers of the gates of the tabernacle: and their fathers, being over the host of the LORD, were keepers of the entry.
1CHR|9|20|And Phinehas the son of Eleazar was the ruler over them in time past, and the LORD was with him.
1CHR|9|21|And Zechariah the son of Meshelemiah was porter of the door of the tabernacle of the congregation.
1CHR|9|22|All these which were chosen to be porters in the gates were two hundred and twelve. These were reckoned by their genealogy in their villages, whom David and Samuel the seer did ordain in their set office.
1CHR|9|23|So they and their children had the oversight of the gates of the house of the LORD, namely, the house of the tabernacle, by wards.
1CHR|9|24|In four quarters were the porters, toward the east, west, north, and south.
1CHR|9|25|And their brethren, which were in their villages, were to come after seven days from time to time with them.
1CHR|9|26|For these Levites, the four chief porters, were in their set office, and were over the chambers and treasuries of the house of God.
1CHR|9|27|And they lodged round about the house of God, because the charge was upon them, and the opening thereof every morning pertained to them.
1CHR|9|28|And certain of them had the charge of the ministering vessels, that they should bring them in and out by tale.
1CHR|9|29|Some of them also were appointed to oversee the vessels, and all the instruments of the sanctuary, and the fine flour, and the wine, and the oil, and the frankincense, and the spices.
1CHR|9|30|And some of the sons of the priests made the ointment of the spices.
1CHR|9|31|And Mattithiah, one of the Levites, who was the firstborn of Shallum the Korahite, had the set office over the things that were made in the pans.
1CHR|9|32|And other of their brethren, of the sons of the Kohathites, were over the shewbread, to prepare it every sabbath.
1CHR|9|33|And these are the singers, chief of the fathers of the Levites, who remaining in the chambers were free: for they were employed in that work day and night.
1CHR|9|34|These chief fathers of the Levites were chief throughout their generations; these dwelt at Jerusalem.
1CHR|9|35|And in Gibeon dwelt the father of Gibeon, Jehiel, whose wife's name was Maachah:
1CHR|9|36|And his firstborn son Abdon, then Zur, and Kish, and Baal, and Ner, and Nadab.
1CHR|9|37|And Gedor, and Ahio, and Zechariah, and Mikloth.
1CHR|9|38|And Mikloth begat Shimeam. And they also dwelt with their brethren at Jerusalem, over against their brethren.
1CHR|9|39|And Ner begat Kish; and Kish begat Saul; and Saul begat Jonathan, and Malchishua, and Abinadab, and Eshbaal.
1CHR|9|40|And the son of Jonathan was Meribbaal: and Meribbaal begat Micah.
1CHR|9|41|And the sons of Micah were, Pithon, and Melech, and Tahrea, and Ahaz.
1CHR|9|42|And Ahaz begat Jarah; and Jarah begat Alemeth, and Azmaveth, and Zimri; and Zimri begat Moza;
1CHR|9|43|And Moza begat Binea; and Rephaiah his son, Eleasah his son, Azel his son.
1CHR|9|44|And Azel had six sons, whose names are these, Azrikam, Bocheru, and Ishmael, and Sheariah, and Obadiah, and Hanan: these were the sons of Azel.
1CHR|10|1|Now the Philistines fought against Israel; and the men of Israel fled from before the Philistines, and fell down slain in mount Gilboa.
1CHR|10|2|And the Philistines followed hard after Saul, and after his sons; and the Philistines slew Jonathan, and Abinadab, and Malchishua, the sons of Saul.
1CHR|10|3|And the battle went sore against Saul, and the archers hit him, and he was wounded of the archers.
1CHR|10|4|Then said Saul to his armourbearer, Draw thy sword, and thrust me through therewith; lest these uncircumcised come and abuse me. But his armourbearer would not; for he was sore afraid. So Saul took a sword, and fell upon it.
1CHR|10|5|And when his armourbearer saw that Saul was dead, he fell likewise on the sword, and died.
1CHR|10|6|So Saul died, and his three sons, and all his house died together.
1CHR|10|7|And when all the men of Israel that were in the valley saw that they fled, and that Saul and his sons were dead, then they forsook their cities, and fled: and the Philistines came and dwelt in them.
1CHR|10|8|And it came to pass on the morrow, when the Philistines came to strip the slain, that they found Saul and his sons fallen in mount Gilboa.
1CHR|10|9|And when they had stripped him, they took his head, and his armor, and sent into the land of the Philistines round about, to carry tidings unto their idols, and to the people.
1CHR|10|10|And they put his armor in the house of their gods, and fastened his head in the temple of Dagon.
1CHR|10|11|And when all Jabeshgilead heard all that the Philistines had done to Saul,
1CHR|10|12|They arose, all the valiant men, and took away the body of Saul, and the bodies of his sons, and brought them to Jabesh, and buried their bones under the oak in Jabesh, and fasted seven days.
1CHR|10|13|So Saul died for his transgression which he committed against the LORD, even against the word of the LORD, which he kept not, and also for asking counsel of one that had a familiar spirit, to enquire of it;
1CHR|10|14|And inquired not of the LORD: therefore he slew him, and turned the kingdom unto David the son of Jesse.
1CHR|11|1|Then all Israel gathered themselves to David unto Hebron, saying, Behold, we are thy bone and thy flesh.
1CHR|11|2|And moreover in time past, even when Saul was king, thou wast he that leddest out and broughtest in Israel: and the LORD thy God said unto thee, Thou shalt feed my people Israel, and thou shalt be ruler over my people Israel.
1CHR|11|3|Therefore came all the elders of Israel to the king to Hebron; and David made a covenant with them in Hebron before the LORD; and they anointed David king over Israel, according to the word of the LORD by Samuel.
1CHR|11|4|And David and all Israel went to Jerusalem, which is Jebus; where the Jebusites were, the inhabitants of the land.
1CHR|11|5|And the inhabitants of Jebus said to David, Thou shalt not come hither. Nevertheless David took the castle of Zion, which is the city of David.
1CHR|11|6|And David said, Whosoever smiteth the Jebusites first shall be chief and captain. So Joab the son of Zeruiah went first up, and was chief.
1CHR|11|7|And David dwelt in the castle; therefore they called it the city of David.
1CHR|11|8|And he built the city round about, even from Millo round about: and Joab repaired the rest of the city.
1CHR|11|9|So David waxed greater and greater: for the LORD of hosts was with him.
1CHR|11|10|These also are the chief of the mighty men whom David had, who strengthened themselves with him in his kingdom, and with all Israel, to make him king, according to the word of the LORD concerning Israel.
1CHR|11|11|And this is the number of the mighty men whom David had; Jashobeam, an Hachmonite, the chief of the captains: he lifted up his spear against three hundred slain by him at one time.
1CHR|11|12|And after him was Eleazar the son of Dodo, the Ahohite, who was one of the three mighties.
1CHR|11|13|He was with David at Pasdammim, and there the Philistines were gathered together to battle, where was a parcel of ground full of barley; and the people fled from before the Philistines.
1CHR|11|14|And they set themselves in the midst of that parcel, and delivered it, and slew the Philistines; and the LORD saved them by a great deliverance.
1CHR|11|15|Now three of the thirty captains went down to the rock to David, into the cave of Adullam; and the host of the Philistines encamped in the valley of Rephaim.
1CHR|11|16|And David was then in the hold, and the Philistines' garrison was then at Bethlehem.
1CHR|11|17|And David longed, and said, Oh that one would give me drink of the water of the well of Bethlehem, that is at the gate!
1CHR|11|18|And the three brake through the host of the Philistines, and drew water out of the well of Bethlehem, that was by the gate, and took it, and brought it to David: but David would not drink of it, but poured it out to the LORD.
1CHR|11|19|And said, My God forbid it me, that I should do this thing: shall I drink the blood of these men that have put their lives in jeopardy? for with the jeopardy of their lives they brought it. Therefore he would not drink it. These things did these three mightiest.
1CHR|11|20|And Abishai the brother of Joab, he was chief of the three: for lifting up his spear against three hundred, he slew them, and had a name among the three.
1CHR|11|21|Of the three, he was more honorable than the two; for he was their captain: howbeit he attained not to the first three.
1CHR|11|22|Benaiah the son of Jehoiada, the son of a valiant man of Kabzeel, who had done many acts; he slew two lionlike men of Moab: also he went down and slew a lion in a pit in a snowy day.
1CHR|11|23|And he slew an Egyptian, a man of great stature, five cubits high; and in the Egyptian's hand was a spear like a weaver's beam; and he went down to him with a staff, and plucked the spear out of the Egyptian's hand, and slew him with his own spear.
1CHR|11|24|These things did Benaiah the son of Jehoiada, and had the name among the three mighties.
1CHR|11|25|Behold, he was honorable among the thirty, but attained not to the first three: and David set him over his guard.
1CHR|11|26|Also the valiant men of the armies were, Asahel the brother of Joab, Elhanan the son of Dodo of Bethlehem,
1CHR|11|27|Shammoth the Harorite, Helez the Pelonite,
1CHR|11|28|Ira the son of Ikkesh the Tekoite, Abiezer the Antothite,
1CHR|11|29|Sibbecai the Hushathite, Ilai the Ahohite,
1CHR|11|30|Maharai the Netophathite, Heled the son of Baanah the Netophathite,
1CHR|11|31|Ithai the son of Ribai of Gibeah, that pertained to the children of Benjamin, Benaiah the Pirathonite,
1CHR|11|32|Hurai of the brooks of Gaash, Abiel the Arbathite,
1CHR|11|33|Azmaveth the Baharumite, Eliahba the Shaalbonite,
1CHR|11|34|The sons of Hashem the Gizonite, Jonathan the son of Shage the Hararite,
1CHR|11|35|Ahiam the son of Sacar the Hararite, Eliphal the son of Ur,
1CHR|11|36|Hepher the Mecherathite, Ahijah the Pelonite,
1CHR|11|37|Hezro the Carmelite, Naarai the son of Ezbai,
1CHR|11|38|Joel the brother of Nathan, Mibhar the son of Haggeri,
1CHR|11|39|Zelek the Ammonite, Naharai the Berothite, the armourbearer of Joab the son of Zeruiah,
1CHR|11|40|Ira the Ithrite, Gareb the Ithrite,
1CHR|11|41|Uriah the Hittite, Zabad the son of Ahlai,
1CHR|11|42|Adina the son of Shiza the Reubenite, a captain of the Reubenites, and thirty with him,
1CHR|11|43|Hanan the son of Maachah, and Joshaphat the Mithnite,
1CHR|11|44|Uzzia the Ashterathite, Shama and Jehiel the sons of Hothan the Aroerite,
1CHR|11|45|Jediael the son of Shimri, and Joha his brother, the Tizite,
1CHR|11|46|Eliel the Mahavite, and Jeribai, and Joshaviah, the sons of Elnaam, and Ithmah the Moabite,
1CHR|11|47|Eliel, and Obed, and Jasiel the Mesobaite.
1CHR|12|1|Now these are they that came to David to Ziklag, while he yet kept himself close because of Saul the son of Kish: and they were among the mighty men, helpers of the war.
1CHR|12|2|They were armed with bows, and could use both the right hand and the left in hurling stones and shooting arrows out of a bow, even of Saul's brethren of Benjamin.
1CHR|12|3|The chief was Ahiezer, then Joash, the sons of Shemaah the Gibeathite; and Jeziel, and Pelet, the sons of Azmaveth; and Berachah, and Jehu the Antothite.
1CHR|12|4|And Ismaiah the Gibeonite, a mighty man among the thirty, and over the thirty; and Jeremiah, and Jahaziel, and Johanan, and Josabad the Gederathite,
1CHR|12|5|Eluzai, and Jerimoth, and Bealiah, and Shemariah, and Shephatiah the Haruphite,
1CHR|12|6|Elkanah, and Jesiah, and Azareel, and Joezer, and Jashobeam, the Korhites,
1CHR|12|7|And Joelah, and Zebadiah, the sons of Jeroham of Gedor.
1CHR|12|8|And of the Gadites there separated themselves unto David into the hold to the wilderness men of might, and men of war fit for the battle, that could handle shield and buckler, whose faces were like the faces of lions, and were as swift as the roes upon the mountains;
1CHR|12|9|Ezer the first, Obadiah the second, Eliab the third,
1CHR|12|10|Mishmannah the fourth, Jeremiah the fifth,
1CHR|12|11|Attai the sixth, Eliel the seventh,
1CHR|12|12|Johanan the eighth, Elzabad the ninth,
1CHR|12|13|Jeremiah the tenth, Machbanai the eleventh.
1CHR|12|14|These were of the sons of Gad, captains of the host: one of the least was over an hundred, and the greatest over a thousand.
1CHR|12|15|These are they that went over Jordan in the first month, when it had overflown all his banks; and they put to flight all them of the valleys, both toward the east, and toward the west.
1CHR|12|16|And there came of the children of Benjamin and Judah to the hold unto David.
1CHR|12|17|And David went out to meet them, and answered and said unto them, If ye be come peaceably unto me to help me, mine heart shall be knit unto you: but if ye be come to betray me to mine enemies, seeing there is no wrong in mine hands, the God of our fathers look thereon, and rebuke it.
1CHR|12|18|Then the spirit came upon Amasai, who was chief of the captains, and he said, Thine are we, David, and on thy side, thou son of Jesse: peace, peace be unto thee, and peace be to thine helpers; for thy God helpeth thee. Then David received them, and made them captains of the band.
1CHR|12|19|And there fell some of Manasseh to David, when he came with the Philistines against Saul to battle: but they helped them not: for the lords of the Philistines upon advisement sent him away, saying, He will fall to his master Saul to the jeopardy of our heads.
1CHR|12|20|As he went to Ziklag, there fell to him of Manasseh, Adnah, and Jozabad, and Jediael, and Michael, and Jozabad, and Elihu, and Zilthai, captains of the thousands that were of Manasseh.
1CHR|12|21|And they helped David against the band of the rovers: for they were all mighty men of valor, and were captains in the host.
1CHR|12|22|For at that time day by day there came to David to help him, until it was a great host, like the host of God.
1CHR|12|23|And these are the numbers of the bands that were ready armed to the war, and came to David to Hebron, to turn the kingdom of Saul to him, according to the word of the LORD.
1CHR|12|24|The children of Judah that bare shield and spear were six thousand and eight hundred, ready armed to the war.
1CHR|12|25|Of the children of Simeon, mighty men of valor for the war, seven thousand and one hundred.
1CHR|12|26|Of the children of Levi four thousand and six hundred.
1CHR|12|27|And Jehoiada was the leader of the Aaronites, and with him were three thousand and seven hundred;
1CHR|12|28|And Zadok, a young man mighty of valor, and of his father's house twenty and two captains.
1CHR|12|29|And of the children of Benjamin, the kindred of Saul, three thousand: for hitherto the greatest part of them had kept the ward of the house of Saul.
1CHR|12|30|And of the children of Ephraim twenty thousand and eight hundred, mighty men of valor, famous throughout the house of their fathers.
1CHR|12|31|And of the half tribe of Manasseh eighteen thousand, which were expressed by name, to come and make David king.
1CHR|12|32|And of the children of Issachar, which were men that had understanding of the times, to know what Israel ought to do; the heads of them were two hundred; and all their brethren were at their commandment.
1CHR|12|33|Of Zebulun, such as went forth to battle, expert in war, with all instruments of war, fifty thousand, which could keep rank: they were not of double heart.
1CHR|12|34|And of Naphtali a thousand captains, and with them with shield and spear thirty and seven thousand.
1CHR|12|35|And of the Danites expert in war twenty and eight thousand and six hundred.
1CHR|12|36|And of Asher, such as went forth to battle, expert in war, forty thousand.
1CHR|12|37|And on the other side of Jordan, of the Reubenites, and the Gadites, and of the half tribe of Manasseh, with all manner of instruments of war for the battle, an hundred and twenty thousand.
1CHR|12|38|All these men of war, that could keep rank, came with a perfect heart to Hebron, to make David king over all Israel: and all the rest also of Israel were of one heart to make David king.
1CHR|12|39|And there they were with David three days, eating and drinking: for their brethren had prepared for them.
1CHR|12|40|Moreover they that were nigh them, even unto Issachar and Zebulun and Naphtali, brought bread on asses, and on camels, and on mules, and on oxen, and meat, meal, cakes of figs, and bunches of raisins, and wine, and oil, and oxen, and sheep abundantly: for there was joy in Israel.
1CHR|13|1|And David consulted with the captains of thousands and hundreds, and with every leader.
1CHR|13|2|And David said unto all the congregation of Israel, If it seem good unto you, and that it be of the LORD our God, let us send abroad unto our brethren every where, that are left in all the land of Israel, and with them also to the priests and Levites which are in their cities and suburbs, that they may gather themselves unto us:
1CHR|13|3|And let us bring again the ark of our God to us: for we inquired not at it in the days of Saul.
1CHR|13|4|And all the congregation said that they would do so: for the thing was right in the eyes of all the people.
1CHR|13|5|So David gathered all Israel together, from Shihor of Egypt even unto the entering of Hemath, to bring the ark of God from Kirjathjearim.
1CHR|13|6|And David went up, and all Israel, to Baalah, that is, to Kirjathjearim, which belonged to Judah, to bring up thence the ark of God the LORD, that dwelleth between the cherubim, whose name is called on it.
1CHR|13|7|And they carried the ark of God in a new cart out of the house of Abinadab: and Uzza and Ahio drave the cart.
1CHR|13|8|And David and all Israel played before God with all their might, and with singing, and with harps, and with psalteries, and with timbrels, and with cymbals, and with trumpets.
1CHR|13|9|And when they came unto the threshingfloor of Chidon, Uzza put forth his hand to hold the ark; for the oxen stumbled.
1CHR|13|10|And the anger of the LORD was kindled against Uzza, and he smote him, because he put his hand to the ark: and there he died before God.
1CHR|13|11|And David was displeased, because the LORD had made a breach upon Uzza: wherefore that place is called Perezuzza to this day.
1CHR|13|12|And David was afraid of God that day, saying, How shall I bring the ark of God home to me?
1CHR|13|13|So David brought not the ark home to himself to the city of David, but carried it aside into the house of Obededom the Gittite.
1CHR|13|14|And the ark of God remained with the family of Obededom in his house three months. And the LORD blessed the house of Obededom, and all that he had.
1CHR|14|1|Now Hiram king of Tyre sent messengers to David, and timber of cedars, with masons and carpenters, to build him an house.
1CHR|14|2|And David perceived that the LORD had confirmed him king over Israel, for his kingdom was lifted up on high, because of his people Israel.
1CHR|14|3|And David took more wives at Jerusalem: and David begat more sons and daughters.
1CHR|14|4|Now these are the names of his children which he had in Jerusalem; Shammua, and Shobab, Nathan, and Solomon,
1CHR|14|5|And Ibhar, and Elishua, and Elpalet,
1CHR|14|6|And Nogah, and Nepheg, and Japhia,
1CHR|14|7|And Elishama, and Beeliada, and Eliphalet.
1CHR|14|8|And when the Philistines heard that David was anointed king over all Israel, all the Philistines went up to seek David. And David heard of it, and went out against them.
1CHR|14|9|And the Philistines came and spread themselves in the valley of Rephaim.
1CHR|14|10|And David inquired of God, saying, Shall I go up against the Philistines? And wilt thou deliver them into mine hand? And the LORD said unto him, Go up; for I will deliver them into thine hand.
1CHR|14|11|So they came up to Baalperazim; and David smote them there. Then David said, God hath broken in upon mine enemies by mine hand like the breaking forth of waters: therefore they called the name of that place Baalperazim.
1CHR|14|12|And when they had left their gods there, David gave a commandment, and they were burned with fire.
1CHR|14|13|And the Philistines yet again spread themselves abroad in the valley.
1CHR|14|14|Therefore David inquired again of God; and God said unto him, Go not up after them; turn away from them, and come upon them over against the mulberry trees.
1CHR|14|15|And it shall be, when thou shalt hear a sound of going in the tops of the mulberry trees, that then thou shalt go out to battle: for God is gone forth before thee to smite the host of the Philistines.
1CHR|14|16|David therefore did as God commanded him: and they smote the host of the Philistines from Gibeon even to Gazer.
1CHR|14|17|And the fame of David went out into all lands; and the LORD brought the fear of him upon all nations.
1CHR|15|1|And David made him houses in the city of David, and prepared a place for the ark of God, and pitched for it a tent.
1CHR|15|2|Then David said, None ought to carry the ark of God but the Levites: for them hath the LORD chosen to carry the ark of God, and to minister unto him for ever.
1CHR|15|3|And David gathered all Israel together to Jerusalem, to bring up the ark of the LORD unto his place, which he had prepared for it.
1CHR|15|4|And David assembled the children of Aaron, and the Levites:
1CHR|15|5|Of the sons of Kohath; Uriel the chief, and his brethren an hundred and twenty:
1CHR|15|6|Of the sons of Merari; Asaiah the chief, and his brethren two hundred and twenty:
1CHR|15|7|Of the sons of Gershom; Joel the chief and his brethren an hundred and thirty:
1CHR|15|8|Of the sons of Elizaphan; Shemaiah the chief, and his brethren two hundred:
1CHR|15|9|Of the sons of Hebron; Eliel the chief, and his brethren fourscore:
1CHR|15|10|Of the sons of Uzziel; Amminadab the chief, and his brethren an hundred and twelve.
1CHR|15|11|And David called for Zadok and Abiathar the priests, and for the Levites, for Uriel, Asaiah, and Joel, Shemaiah, and Eliel, and Amminadab,
1CHR|15|12|And said unto them, Ye are the chief of the fathers of the Levites: sanctify yourselves, both ye and your brethren, that ye may bring up the ark of the LORD God of Israel unto the place that I have prepared for it.
1CHR|15|13|For because ye did it not at the first, the LORD our God made a breach upon us, for that we sought him not after the due order.
1CHR|15|14|So the priests and the Levites sanctified themselves to bring up the ark of the LORD God of Israel.
1CHR|15|15|And the children of the Levites bare the ark of God upon their shoulders with the staves thereon, as Moses commanded according to the word of the LORD.
1CHR|15|16|And David spake to the chief of the Levites to appoint their brethren to be the singers with instruments of music, psalteries and harps and cymbals, sounding, by lifting up the voice with joy.
1CHR|15|17|So the Levites appointed Heman the son of Joel; and of his brethren, Asaph the son of Berechiah; and of the sons of Merari their brethren, Ethan the son of Kushaiah;
1CHR|15|18|And with them their brethren of the second degree, Zechariah, Ben, and Jaaziel, and Shemiramoth, and Jehiel, and Unni, Eliab, and Benaiah, and Maaseiah, and Mattithiah, and Elipheleh, and Mikneiah, and Obededom, and Jeiel, the porters.
1CHR|15|19|So the singers, Heman, Asaph, and Ethan, were appointed to sound with cymbals of brass;
1CHR|15|20|And Zechariah, and Aziel, and Shemiramoth, and Jehiel, and Unni, and Eliab, and Maaseiah, and Benaiah, with psalteries on Alamoth;
1CHR|15|21|And Mattithiah, and Elipheleh, and Mikneiah, and Obededom, and Jeiel, and Azaziah, with harps on the Sheminith to excel.
1CHR|15|22|And Chenaniah, chief of the Levites, was for song: he instructed about the song, because he was skillful.
1CHR|15|23|And Berechiah and Elkanah were doorkeepers for the ark.
1CHR|15|24|And Shebaniah, and Jehoshaphat, and Nethaneel, and Amasai, and Zechariah, and Benaiah, and Eliezer, the priests, did blow with the trumpets before the ark of God: and Obededom and Jehiah were doorkeepers for the ark.
1CHR|15|25|So David, and the elders of Israel, and the captains over thousands, went to bring up the ark of the covenant of the LORD out of the house of Obededom with joy.
1CHR|15|26|And it came to pass, when God helped the Levites that bare the ark of the covenant of the LORD, that they offered seven bullocks and seven rams.
1CHR|15|27|And David was clothed with a robe of fine linen, and all the Levites that bare the ark, and the singers, and Chenaniah the master of the song with the singers: David also had upon him an ephod of linen.
1CHR|15|28|Thus all Israel brought up the ark of the covenant of the LORD with shouting, and with sound of the cornet, and with trumpets, and with cymbals, making a noise with psalteries and harps.
1CHR|15|29|And it came to pass, as the ark of the covenant of the LORD came to the city of David, that Michal, the daughter of Saul looking out at a window saw king David dancing and playing: and she despised him in her heart.
1CHR|16|1|So they brought the ark of God, and set it in the midst of the tent that David had pitched for it: and they offered burnt sacrifices and peace offerings before God.
1CHR|16|2|And when David had made an end of offering the burnt offerings and the peace offerings, he blessed the people in the name of the LORD.
1CHR|16|3|And he dealt to every one of Israel, both man and woman, to every one a loaf of bread, and a good piece of flesh, and a flagon of wine.
1CHR|16|4|And he appointed certain of the Levites to minister before the ark of the LORD, and to record, and to thank and praise the LORD God of Israel:
1CHR|16|5|Asaph the chief, and next to him Zechariah, Jeiel, and Shemiramoth, and Jehiel, and Mattithiah, and Eliab, and Benaiah, and Obededom: and Jeiel with psalteries and with harps; but Asaph made a sound with cymbals;
1CHR|16|6|Benaiah also and Jahaziel the priests with trumpets continually before the ark of the covenant of God.
1CHR|16|7|Then on that day David delivered first this psalm to thank the LORD into the hand of Asaph and his brethren.
1CHR|16|8|Give thanks unto the LORD, call upon his name, make known his deeds among the people.
1CHR|16|9|Sing unto him, sing psalms unto him, talk ye of all his wondrous works.
1CHR|16|10|Glory ye in his holy name: let the heart of them rejoice that seek the LORD.
1CHR|16|11|Seek the LORD and his strength, seek his face continually.
1CHR|16|12|Remember his marvelous works that he hath done, his wonders, and the judgments of his mouth;
1CHR|16|13|O ye seed of Israel his servant, ye children of Jacob, his chosen ones.
1CHR|16|14|He is the LORD our God; his judgments are in all the earth.
1CHR|16|15|Be ye mindful always of his covenant; the word which he commanded to a thousand generations;
1CHR|16|16|Even of the covenant which he made with Abraham, and of his oath unto Isaac;
1CHR|16|17|And hath confirmed the same to Jacob for a law, and to Israel for an everlasting covenant,
1CHR|16|18|Saying, Unto thee will I give the land of Canaan, the lot of your inheritance;
1CHR|16|19|When ye were but few, even a few, and strangers in it.
1CHR|16|20|And when they went from nation to nation, and from one kingdom to another people;
1CHR|16|21|He suffered no man to do them wrong: yea, he reproved kings for their sakes,
1CHR|16|22|Saying, Touch not mine anointed, and do my prophets no harm.
1CHR|16|23|Sing unto the LORD, all the earth; show forth from day to day his salvation.
1CHR|16|24|Declare his glory among the heathen; his marvelous works among all nations.
1CHR|16|25|For great is the LORD, and greatly to be praised: he also is to be feared above all gods.
1CHR|16|26|For all the gods of the people are idols: but the LORD made the heavens.
1CHR|16|27|Glory and honor are in his presence; strength and gladness are in his place.
1CHR|16|28|Give unto the LORD, ye kindred of the people, give unto the LORD glory and strength.
1CHR|16|29|Give unto the LORD the glory due unto his name: bring an offering, and come before him: worship the LORD in the beauty of holiness.
1CHR|16|30|Fear before him, all the earth: the world also shall be stable, that it be not moved.
1CHR|16|31|Let the heavens be glad, and let the earth rejoice: and let men say among the nations, The LORD reigneth.
1CHR|16|32|Let the sea roar, and the fulness thereof: let the fields rejoice, and all that is therein.
1CHR|16|33|Then shall the trees of the wood sing out at the presence of the LORD, because he cometh to judge the earth.
1CHR|16|34|O give thanks unto the LORD; for he is good; for his mercy endureth for ever.
1CHR|16|35|And say ye, Save us, O God of our salvation, and gather us together, and deliver us from the heathen, that we may give thanks to thy holy name, and glory in thy praise.
1CHR|16|36|Blessed be the LORD God of Israel for ever and ever. And all the people said, Amen, and praised the LORD.
1CHR|16|37|So he left there before the ark of the covenant of the LORD Asaph and his brethren, to minister before the ark continually, as every day's work required:
1CHR|16|38|And Obededom with their brethren, threescore and eight; Obededom also the son of Jeduthun and Hosah to be porters:
1CHR|16|39|And Zadok the priest, and his brethren the priests, before the tabernacle of the LORD in the high place that was at Gibeon,
1CHR|16|40|To offer burnt offerings unto the LORD upon the altar of the burnt offering continually morning and evening, and to do according to all that is written in the law of the LORD, which he commanded Israel;
1CHR|16|41|And with them Heman and Jeduthun, and the rest that were chosen, who were expressed by name, to give thanks to the LORD, because his mercy endureth for ever;
1CHR|16|42|And with them Heman and Jeduthun with trumpets and cymbals for those that should make a sound, and with musical instruments of God. And the sons of Jeduthun were porters.
1CHR|16|43|And all the people departed every man to his house: and David returned to bless his house.
1CHR|17|1|Now it came to pass, as David sat in his house, that David said to Nathan the prophet, Lo, I dwell in an house of cedars, but the ark of the covenant of the LORD remaineth under curtains.
1CHR|17|2|Then Nathan said unto David, Do all that is in thine heart; for God is with thee.
1CHR|17|3|And it came to pass the same night, that the word of God came to Nathan, saying,
1CHR|17|4|Go and tell David my servant, Thus saith the LORD, Thou shalt not build me an house to dwell in:
1CHR|17|5|For I have not dwelt in an house since the day that I brought up Israel unto this day; but have gone from tent to tent, and from one tabernacle to another.
1CHR|17|6|Wheresoever I have walked with all Israel, spake I a word to any of the judges of Israel, whom I commanded to feed my people, saying, Why have ye not built me an house of cedars?
1CHR|17|7|Now therefore thus shalt thou say unto my servant David, Thus saith the LORD of hosts, I took thee from the sheepcote, even from following the sheep, that thou shouldest be ruler over my people Israel:
1CHR|17|8|And I have been with thee whithersoever thou hast walked, and have cut off all thine enemies from before thee, and have made thee a name like the name of the great men that are in the earth.
1CHR|17|9|Also I will ordain a place for my people Israel, and will plant them, and they shall dwell in their place, and shall be moved no more; neither shall the children of wickedness waste them any more, as at the beginning,
1CHR|17|10|And since the time that I commanded judges to be over my people Israel. Moreover I will subdue all thine enemies. Furthermore I tell thee that the LORD will build thee an house.
1CHR|17|11|And it shall come to pass, when thy days be expired that thou must go to be with thy fathers, that I will raise up thy seed after thee, which shall be of thy sons; and I will establish his kingdom.
1CHR|17|12|He shall build me an house, and I will stablish his throne for ever.
1CHR|17|13|I will be his father, and he shall be my son: and I will not take my mercy away from him, as I took it from him that was before thee:
1CHR|17|14|But I will settle him in mine house and in my kingdom for ever: and his throne shall be established for evermore.
1CHR|17|15|According to all these words, and according to all this vision, so did Nathan speak unto David.
1CHR|17|16|And David the king came and sat before the LORD, and said, Who am I, O LORD God, and what is mine house, that thou hast brought me hitherto?
1CHR|17|17|And yet this was a small thing in thine eyes, O God; for thou hast also spoken of thy servant's house for a great while to come, and hast regarded me according to the estate of a man of high degree, O LORD God.
1CHR|17|18|What can David speak more to thee for the honor of thy servant? for thou knowest thy servant.
1CHR|17|19|O LORD, for thy servant's sake, and according to thine own heart, hast thou done all this greatness, in making known all these great things.
1CHR|17|20|O LORD, there is none like thee, neither is there any God beside thee, according to all that we have heard with our ears.
1CHR|17|21|And what one nation in the earth is like thy people Israel, whom God went to redeem to be his own people, to make thee a name of greatness and terribleness, by driving out nations from before thy people whom thou hast redeemed out of Egypt?
1CHR|17|22|For thy people Israel didst thou make thine own people for ever; and thou, LORD, becamest their God.
1CHR|17|23|Therefore now, LORD, let the thing that thou hast spoken concerning thy servant and concerning his house be established for ever, and do as thou hast said.
1CHR|17|24|Let it even be established, that thy name may be magnified for ever, saying, The LORD of hosts is the God of Israel, even a God to Israel: and let the house of David thy servant be established before thee.
1CHR|17|25|For thou, O my God, hast told thy servant that thou wilt build him an house: therefore thy servant hath found in his heart to pray before thee.
1CHR|17|26|And now, LORD, thou art God, and hast promised this goodness unto thy servant:
1CHR|17|27|Now therefore let it please thee to bless the house of thy servant, that it may be before thee for ever: for thou blessest, O LORD, and it shall be blessed for ever.
1CHR|18|1|Now after this it came to pass, that David smote the Philistines, and subdued them, and took Gath and her towns out of the hand of the Philistines.
1CHR|18|2|And he smote Moab; and the Moabites became David's servants, and brought gifts.
1CHR|18|3|And David smote Hadarezer king of Zobah unto Hamath, as he went to stablish his dominion by the river Euphrates.
1CHR|18|4|And David took from him a thousand chariots, and seven thousand horsemen, and twenty thousand footmen: David also houghed all the chariot horses, but reserved of them an hundred chariots.
1CHR|18|5|And when the Syrians of Damascus came to help Hadarezer king of Zobah, David slew of the Syrians two and twenty thousand men.
1CHR|18|6|Then David put garrisons in Syriadamascus; and the Syrians became David's servants, and brought gifts. Thus the LORD preserved David whithersoever he went.
1CHR|18|7|And David took the shields of gold that were on the servants of Hadarezer, and brought them to Jerusalem.
1CHR|18|8|Likewise from Tibhath, and from Chun, cities of Hadarezer, brought David very much brass, wherewith Solomon made the brazen sea, and the pillars, and the vessels of brass.
1CHR|18|9|Now when Tou king of Hamath heard how David had smitten all the host of Hadarezer king of Zobah;
1CHR|18|10|He sent Hadoram his son to king David, to enquire of his welfare, and to congratulate him, because he had fought against Hadarezer, and smitten him; (for Hadarezer had war with Tou;) and with him all manner of vessels of gold and silver and brass.
1CHR|18|11|Them also king David dedicated unto the LORD, with the silver and the gold that he brought from all these nations; from Edom, and from Moab, and from the children of Ammon, and from the Philistines, and from Amalek.
1CHR|18|12|Moreover Abishai the son of Zeruiah slew of the Edomites in the valley of salt eighteen thousand.
1CHR|18|13|And he put garrisons in Edom; and all the Edomites became David's servants. Thus the LORD preserved David whithersoever he went.
1CHR|18|14|So David reigned over all Israel, and executed judgment and justice among all his people.
1CHR|18|15|And Joab the son of Zeruiah was over the host; and Jehoshaphat the son of Ahilud, recorder.
1CHR|18|16|And Zadok the son of Ahitub, and Abimelech the son of Abiathar, were the priests; and Shavsha was scribe;
1CHR|18|17|And Benaiah the son of Jehoiada was over the Cherethites and the Pelethites; and the sons of David were chief about the king.
1CHR|19|1|Now it came to pass after this, that Nahash the king of the children of Ammon died, and his son reigned in his stead.
1CHR|19|2|And David said, I will show kindness unto Hanun the son of Nahash, because his father showed kindness to me. And David sent messengers to comfort him concerning his father. So the servants of David came into the land of the children of Ammon to Hanun, to comfort him.
1CHR|19|3|But the princes of the children of Ammon said to Hanun, Thinkest thou that David doth honor thy father, that he hath sent comforters unto thee? are not his servants come unto thee for to search, and to overthrow, and to spy out the land?
1CHR|19|4|Wherefore Hanun took David's servants, and shaved them, and cut off their garments in the midst hard by their buttocks, and sent them away.
1CHR|19|5|Then there went certain, and told David how the men were served. And he sent to meet them: for the men were greatly ashamed. And the king said, Tarry at Jericho until your beards be grown, and then return.
1CHR|19|6|And when the children of Ammon saw that they had made themselves odious to David, Hanun and the children of Ammon sent a thousand talents of silver to hire them chariots and horsemen out of Mesopotamia, and out of Syriamaachah, and out of Zobah.
1CHR|19|7|So they hired thirty and two thousand chariots, and the king of Maachah and his people; who came and pitched before Medeba. And the children of Ammon gathered themselves together from their cities, and came to battle.
1CHR|19|8|And when David heard of it, he sent Joab, and all the host of the mighty men.
1CHR|19|9|And the children of Ammon came out, and put the battle in array before the gate of the city: and the kings that were come were by themselves in the field.
1CHR|19|10|Now when Joab saw that the battle was set against him before and behind, he chose out of all the choice of Israel, and put them in array against the Syrians.
1CHR|19|11|And the rest of the people he delivered unto the hand of Abishai his brother, and they set themselves in array against the children of Ammon.
1CHR|19|12|And he said, If the Syrians be too strong for me, then thou shalt help me: but if the children of Ammon be too strong for thee, then I will help thee.
1CHR|19|13|Be of good courage, and let us behave ourselves valiantly for our people, and for the cities of our God: and let the LORD do that which is good in his sight.
1CHR|19|14|So Joab and the people that were with him drew nigh before the Syrians unto the battle; and they fled before him.
1CHR|19|15|And when the children of Ammon saw that the Syrians were fled, they likewise fled before Abishai his brother, and entered into the city. Then Joab came to Jerusalem.
1CHR|19|16|And when the Syrians saw that they were put to the worse before Israel, they sent messengers, and drew forth the Syrians that were beyond the river: and Shophach the captain of the host of Hadarezer went before them.
1CHR|19|17|And it was told David; and he gathered all Israel, and passed over Jordan, and came upon them, and set the battle in array against them. So when David had put the battle in array against the Syrians, they fought with him.
1CHR|19|18|But the Syrians fled before Israel; and David slew of the Syrians seven thousand men which fought in chariots, and forty thousand footmen, and killed Shophach the captain of the host.
1CHR|19|19|And when the servants of Hadarezer saw that they were put to the worse before Israel, they made peace with David, and became his servants: neither would the Syrians help the children of Ammon any more.
1CHR|20|1|And it came to pass, that after the year was expired, at the time that kings go out to battle, Joab led forth the power of the army, and wasted the country of the children of Ammon, and came and besieged Rabbah. But David tarried at Jerusalem. And Joab smote Rabbah, and destroyed it.
1CHR|20|2|And David took the crown of their king from off his head, and found it to weigh a talent of gold, and there were precious stones in it; and it was set upon David's head: and he brought also exceeding much spoil out of the city.
1CHR|20|3|And he brought out the people that were in it, and cut them with saws, and with harrows of iron, and with axes. Even so dealt David with all the cities of the children of Ammon. And David and all the people returned to Jerusalem.
1CHR|20|4|And it came to pass after this, that there arose war at Gezer with the Philistines; at which time Sibbechai the Hushathite slew Sippai, that was of the children of the giant: and they were subdued.
1CHR|20|5|And there was war again with the Philistines; and Elhanan the son of Jair slew Lahmi the brother of Goliath the Gittite, whose spear staff was like a weaver's beam.
1CHR|20|6|And yet again there was war at Gath, where was a man of great stature, whose fingers and toes were four and twenty, six on each hand, and six on each foot and he also was the son of the giant.
1CHR|20|7|But when he defied Israel, Jonathan the son of Shimea David's brother slew him.
1CHR|20|8|These were born unto the giant in Gath; and they fell by the hand of David, and by the hand of his servants.
1CHR|21|1|And Satan stood up against Israel, and provoked David to number Israel.
1CHR|21|2|And David said to Joab and to the rulers of the people, Go, number Israel from Beersheba even to Dan; and bring the number of them to me, that I may know it.
1CHR|21|3|And Joab answered, The LORD make his people an hundred times so many more as they be: but, my lord the king, are they not all my lord's servants? why then doth my lord require this thing? why will he be a cause of trespass to Israel?
1CHR|21|4|Nevertheless the king's word prevailed against Joab. Wherefore Joab departed, and went throughout all Israel, and came to Jerusalem.
1CHR|21|5|And Joab gave the sum of the number of the people unto David. And all they of Israel were a thousand thousand and an hundred thousand men that drew sword: and Judah was four hundred threescore and ten thousand men that drew sword.
1CHR|21|6|But Levi and Benjamin counted he not among them: for the king's word was abominable to Joab.
1CHR|21|7|And God was displeased with this thing; therefore he smote Israel.
1CHR|21|8|And David said unto God, I have sinned greatly, because I have done this thing: but now, I beseech thee, do away the iniquity of thy servant; for I have done very foolishly.
1CHR|21|9|And the LORD spake unto Gad, David's seer, saying,
1CHR|21|10|Go and tell David, saying, Thus saith the LORD, I offer thee three things: choose thee one of them, that I may do it unto thee.
1CHR|21|11|So Gad came to David, and said unto him, Thus saith the LORD, Choose thee
1CHR|21|12|Either three years' famine; or three months to be destroyed before thy foes, while that the sword of thine enemies overtaketh thee; or else three days the sword of the LORD, even the pestilence, in the land, and the angel of the LORD destroying throughout all the coasts of Israel. Now therefore advise thyself what word I shall bring again to him that sent me.
1CHR|21|13|And David said unto Gad, I am in a great strait: let me fall now into the hand of the LORD; for very great are his mercies: but let me not fall into the hand of man.
1CHR|21|14|So the LORD sent pestilence upon Israel: and there fell of Israel seventy thousand men.
1CHR|21|15|And God sent an angel unto Jerusalem to destroy it: and as he was destroying, the LORD beheld, and he repented him of the evil, and said to the angel that destroyed, It is enough, stay now thine hand. And the angel of the LORD stood by the threshingfloor of Ornan the Jebusite.
1CHR|21|16|And David lifted up his eyes, and saw the angel of the LORD stand between the earth and the heaven, having a drawn sword in his hand stretched out over Jerusalem. Then David and the elders of Israel, who were clothed in sackcloth, fell upon their faces.
1CHR|21|17|And David said unto God, Is it not I that commanded the people to be numbered? even I it is that have sinned and done evil indeed; but as for these sheep, what have they done? let thine hand, I pray thee, O LORD my God, be on me, and on my father's house; but not on thy people, that they should be plagued.
1CHR|21|18|Then the angel of the LORD commanded Gad to say to David, that David should go up, and set up an altar unto the LORD in the threshingfloor of Ornan the Jebusite.
1CHR|21|19|And David went up at the saying of Gad, which he spake in the name of the LORD.
1CHR|21|20|And Ornan turned back, and saw the angel; and his four sons with him hid themselves. Now Ornan was threshing wheat.
1CHR|21|21|And as David came to Ornan, Ornan looked and saw David, and went out of the threshingfloor, and bowed himself to David with his face to the ground.
1CHR|21|22|Then David said to Ornan, Grant me the place of this threshingfloor, that I may build an altar therein unto the LORD: thou shalt grant it me for the full price: that the plague may be stayed from the people.
1CHR|21|23|And Ornan said unto David, Take it to thee, and let my lord the king do that which is good in his eyes: lo, I give thee the oxen also for burnt offerings, and the threshing instruments for wood, and the wheat for the meat offering; I give it all.
1CHR|21|24|And king David said to Ornan, Nay; but I will verily buy it for the full price: for I will not take that which is thine for the LORD, nor offer burnt offerings without cost.
1CHR|21|25|So David gave to Ornan for the place six hundred shekels of gold by weight.
1CHR|21|26|And David built there an altar unto the LORD, and offered burnt offerings and peace offerings, and called upon the LORD; and he answered him from heaven by fire upon the altar of burnt offering.
1CHR|21|27|And the LORD commanded the angel; and he put up his sword again into the sheath thereof.
1CHR|21|28|At that time when David saw that the LORD had answered him in the threshingfloor of Ornan the Jebusite, then he sacrificed there.
1CHR|21|29|For the tabernacle of the LORD, which Moses made in the wilderness, and the altar of the burnt offering, were at that season in the high place at Gibeon.
1CHR|21|30|But David could not go before it to enquire of God: for he was afraid because of the sword of the angel of the LORD.
1CHR|22|1|Then David said, This is the house of the LORD God, and this is the altar of the burnt offering for Israel.
1CHR|22|2|And David commanded to gather together the strangers that were in the land of Israel; and he set masons to hew wrought stones to build the house of God.
1CHR|22|3|And David prepared iron in abundance for the nails for the doors of the gates, and for the joinings; and brass in abundance without weight;
1CHR|22|4|Also cedar trees in abundance: for the Zidonians and they of Tyre brought much cedar wood to David.
1CHR|22|5|And David said, Solomon my son is young and tender, and the house that is to be builded for the LORD must be exceeding magnificent, of fame and of glory throughout all countries: I will therefore now make preparation for it. So David prepared abundantly before his death.
1CHR|22|6|Then he called for Solomon his son, and charged him to build an house for the LORD God of Israel.
1CHR|22|7|And David said to Solomon, My son, as for me, it was in my mind to build an house unto the name of the LORD my God:
1CHR|22|8|But the word of the LORD came to me, saying, Thou hast shed blood abundantly, and hast made great wars: thou shalt not build an house unto my name, because thou hast shed much blood upon the earth in my sight.
1CHR|22|9|Behold, a son shall be born to thee, who shall be a man of rest; and I will give him rest from all his enemies round about: for his name shall be Solomon, and I will give peace and quietness unto Israel in his days.
1CHR|22|10|He shall build an house for my name; and he shall be my son, and I will be his father; and I will establish the throne of his kingdom over Israel for ever.
1CHR|22|11|Now, my son, the LORD be with thee; and prosper thou, and build the house of the LORD thy God, as he hath said of thee.
1CHR|22|12|Only the LORD give thee wisdom and understanding, and give thee charge concerning Israel, that thou mayest keep the law of the LORD thy God.
1CHR|22|13|Then shalt thou prosper, if thou takest heed to fulfil the statutes and judgments which the LORD charged Moses with concerning Israel: be strong, and of good courage; dread not, nor be dismayed.
1CHR|22|14|Now, behold, in my trouble I have prepared for the house of the LORD an hundred thousand talents of gold, and a thousand thousand talents of silver; and of brass and iron without weight; for it is in abundance: timber also and stone have I prepared; and thou mayest add thereto.
1CHR|22|15|Moreover there are workmen with thee in abundance, hewers and workers of stone and timber, and all manner of cunning men for every manner of work.
1CHR|22|16|Of the gold, the silver, and the brass, and the iron, there is no number. Arise therefore, and be doing, and the LORD be with thee.
1CHR|22|17|David also commanded all the princes of Israel to help Solomon his son, saying,
1CHR|22|18|Is not the LORD your God with you? and hath he not given you rest on every side? for he hath given the inhabitants of the land into mine hand; and the land is subdued before the LORD, and before his people.
1CHR|22|19|Now set your heart and your soul to seek the LORD your God; arise therefore, and build ye the sanctuary of the LORD God, to bring the ark of the covenant of the LORD, and the holy vessels of God, into the house that is to be built to the name of the LORD.
1CHR|23|1|So when David was old and full of days, he made Solomon his son king over Israel.
1CHR|23|2|And he gathered together all the princes of Israel, with the priests and the Levites.
1CHR|23|3|Now the Levites were numbered from the age of thirty years and upward: and their number by their polls, man by man, was thirty and eight thousand.
1CHR|23|4|Of which, twenty and four thousand were to set forward the work of the house of the LORD; and six thousand were officers and judges:
1CHR|23|5|Moreover four thousand were porters; and four thousand praised the LORD with the instruments which I made, said David, to praise therewith.
1CHR|23|6|And David divided them into courses among the sons of Levi, namely, Gershon, Kohath, and Merari.
1CHR|23|7|Of the Gershonites were, Laadan, and Shimei.
1CHR|23|8|The sons of Laadan; the chief was Jehiel, and Zetham, and Joel, three.
1CHR|23|9|The sons of Shimei; Shelomith, and Haziel, and Haran, three. These were the chief of the fathers of Laadan.
1CHR|23|10|And the sons of Shimei were, Jahath, Zina, and Jeush, and Beriah. These four were the sons of Shimei.
1CHR|23|11|And Jahath was the chief, and Zizah the second: but Jeush and Beriah had not many sons; therefore they were in one reckoning, according to their father's house.
1CHR|23|12|The sons of Kohath; Amram, Izhar, Hebron, and Uzziel, four.
1CHR|23|13|The sons of Amram; Aaron and Moses: and Aaron was separated, that he should sanctify the most holy things, he and his sons for ever, to burn incense before the LORD, to minister unto him, and to bless in his name for ever.
1CHR|23|14|Now concerning Moses the man of God, his sons were named of the tribe of Levi.
1CHR|23|15|The sons of Moses were, Gershom, and Eliezer.
1CHR|23|16|Of the sons of Gershom, Shebuel was the chief.
1CHR|23|17|And the sons of Eliezer were, Rehabiah the chief. And Eliezer had none other sons; but the sons of Rehabiah were very many.
1CHR|23|18|Of the sons of Izhar; Shelomith the chief.
1CHR|23|19|Of the sons of Hebron; Jeriah the first, Amariah the second, Jahaziel the third, and Jekameam the fourth.
1CHR|23|20|Of the sons of Uzziel; Micah the first and Jesiah the second.
1CHR|23|21|The sons of Merari; Mahli, and Mushi. The sons of Mahli; Eleazar, and Kish.
1CHR|23|22|And Eleazar died, and had no sons, but daughters: and their brethren the sons of Kish took them.
1CHR|23|23|The sons of Mushi; Mahli, and Eder, and Jeremoth, three.
1CHR|23|24|These were the sons of Levi after the house of their fathers; even the chief of the fathers, as they were counted by number of names by their polls, that did the work for the service of the house of the LORD, from the age of twenty years and upward.
1CHR|23|25|For David said, The LORD God of Israel hath given rest unto his people, that they may dwell in Jerusalem for ever:
1CHR|23|26|And also unto the Levites; they shall no more carry the tabernacle, nor any vessels of it for the service thereof.
1CHR|23|27|For by the last words of David the Levites were numbered from twenty years old and above:
1CHR|23|28|Because their office was to wait on the sons of Aaron for the service of the house of the LORD, in the courts, and in the chambers, and in the purifying of all holy things, and the work of the service of the house of God;
1CHR|23|29|Both for the shewbread, and for the fine flour for meat offering, and for the unleavened cakes, and for that which is baked in the pan, and for that which is fried, and for all manner of measure and size;
1CHR|23|30|And to stand every morning to thank and praise the LORD, and likewise at even:
1CHR|23|31|And to offer all burnt sacrifices unto the LORD in the sabbaths, in the new moons, and on the set feasts, by number, according to the order commanded unto them, continually before the LORD:
1CHR|23|32|And that they should keep the charge of the tabernacle of the congregation, and the charge of the holy place, and the charge of the sons of Aaron their brethren, in the service of the house of the LORD.
1CHR|24|1|Now these are the divisions of the sons of Aaron. The sons of Aaron; Nadab, and Abihu, Eleazar, and Ithamar.
1CHR|24|2|But Nadab and Abihu died before their father, and had no children: therefore Eleazar and Ithamar executed the priest's office.
1CHR|24|3|And David distributed them, both Zadok of the sons of Eleazar, and Ahimelech of the sons of Ithamar, according to their offices in their service.
1CHR|24|4|And there were more chief men found of the sons of Eleazar than of the sons of Ithamar, and thus were they divided. Among the sons of Eleazar there were sixteen chief men of the house of their fathers, and eight among the sons of Ithamar according to the house of their fathers.
1CHR|24|5|Thus were they divided by lot, one sort with another; for the governors of the sanctuary, and governors of the house of God, were of the sons of Eleazar, and of the sons of Ithamar.
1CHR|24|6|And Shemaiah the son of Nethaneel the scribe, one of the Levites, wrote them before the king, and the princes, and Zadok the priest, and Ahimelech the son of Abiathar, and before the chief of the fathers of the priests and Levites: one principal household being taken for Eleazar, and one taken for Ithamar.
1CHR|24|7|Now the first lot came forth to Jehoiarib, the second to Jedaiah,
1CHR|24|8|The third to Harim, the fourth to Seorim,
1CHR|24|9|The fifth to Malchijah, the sixth to Mijamin,
1CHR|24|10|The seventh to Hakkoz, the eighth to Abijah,
1CHR|24|11|The ninth to Jeshuah, the tenth to Shecaniah,
1CHR|24|12|The eleventh to Eliashib, the twelfth to Jakim,
1CHR|24|13|The thirteenth to Huppah, the fourteenth to Jeshebeab,
1CHR|24|14|The fifteenth to Bilgah, the sixteenth to Immer,
1CHR|24|15|The seventeenth to Hezir, the eighteenth to Aphses,
1CHR|24|16|The nineteenth to Pethahiah, the twentieth to Jehezekel,
1CHR|24|17|The one and twentieth to Jachin, the two and twentieth to Gamul,
1CHR|24|18|The three and twentieth to Delaiah, the four and twentieth to Maaziah.
1CHR|24|19|These were the orderings of them in their service to come into the house of the LORD, according to their manner, under Aaron their father, as the LORD God of Israel had commanded him.
1CHR|24|20|And the rest of the sons of Levi were these: Of the sons of Amram; Shubael: of the sons of Shubael; Jehdeiah.
1CHR|24|21|Concerning Rehabiah: of the sons of Rehabiah, the first was Isshiah.
1CHR|24|22|Of the Izharites; Shelomoth: of the sons of Shelomoth; Jahath.
1CHR|24|23|And the sons of Hebron; Jeriah the first, Amariah the second, Jahaziel the third, Jekameam the fourth.
1CHR|24|24|Of the sons of Uzziel; Michah: of the sons of Michah; Shamir.
1CHR|24|25|The brother of Michah was Isshiah: of the sons of Isshiah; Zechariah.
1CHR|24|26|The sons of Merari were Mahli and Mushi: the sons of Jaaziah; Beno.
1CHR|24|27|The sons of Merari by Jaaziah; Beno, and Shoham, and Zaccur, and Ibri.
1CHR|24|28|Of Mahli came Eleazar, who had no sons.
1CHR|24|29|Concerning Kish: the son of Kish was Jerahmeel.
1CHR|24|30|The sons also of Mushi; Mahli, and Eder, and Jerimoth. These were the sons of the Levites after the house of their fathers.
1CHR|24|31|These likewise cast lots over against their brethren the sons of Aaron in the presence of David the king, and Zadok, and Ahimelech, and the chief of the fathers of the priests and Levites, even the principal fathers over against their younger brethren.
1CHR|25|1|Moreover David and the captains of the host separated to the service of the sons of Asaph, and of Heman, and of Jeduthun, who should prophesy with harps, with psalteries, and with cymbals: and the number of the workmen according to their service was:
1CHR|25|2|Of the sons of Asaph; Zaccur, and Joseph, and Nethaniah, and Asarelah, the sons of Asaph under the hands of Asaph, which prophesied according to the order of the king.
1CHR|25|3|Of Jeduthun: the sons of Jeduthun; Gedaliah, and Zeri, and Jeshaiah, Hashabiah, and Mattithiah, six, under the hands of their father Jeduthun, who prophesied with a harp, to give thanks and to praise the LORD.
1CHR|25|4|Of Heman: the sons of Heman: Bukkiah, Mattaniah, Uzziel, Shebuel, and Jerimoth, Hananiah, Hanani, Eliathah, Giddalti, and Romamtiezer, Joshbekashah, Mallothi, Hothir, and Mahazioth:
1CHR|25|5|All these were the sons of Heman the king's seer in the words of God, to lift up the horn. And God gave to Heman fourteen sons and three daughters.
1CHR|25|6|All these were under the hands of their father for song in the house of the LORD, with cymbals, psalteries, and harps, for the service of the house of God, according to the king's order to Asaph, Jeduthun, and Heman.
1CHR|25|7|So the number of them, with their brethren that were instructed in the songs of the LORD, even all that were cunning, was two hundred fourscore and eight.
1CHR|25|8|And they cast lots, ward against ward, as well the small as the great, the teacher as the scholar.
1CHR|25|9|Now the first lot came forth for Asaph to Joseph: the second to Gedaliah, who with his brethren and sons were twelve:
1CHR|25|10|The third to Zaccur, he, his sons, and his brethren, were twelve:
1CHR|25|11|The fourth to Izri, he, his sons, and his brethren, were twelve:
1CHR|25|12|The fifth to Nethaniah, he, his sons, and his brethren, were twelve:
1CHR|25|13|The sixth to Bukkiah, he, his sons, and his brethren, were twelve:
1CHR|25|14|The seventh to Jesharelah, he, his sons, and his brethren, were twelve:
1CHR|25|15|The eighth to Jeshaiah, he, his sons, and his brethren, were twelve:
1CHR|25|16|The ninth to Mattaniah, he, his sons, and his brethren, were twelve:
1CHR|25|17|The tenth to Shimei, he, his sons, and his brethren, were twelve:
1CHR|25|18|The eleventh to Azareel, he, his sons, and his brethren, were twelve:
1CHR|25|19|The twelfth to Hashabiah, he, his sons, and his brethren, were twelve:
1CHR|25|20|The thirteenth to Shubael, he, his sons, and his brethren, were twelve:
1CHR|25|21|The fourteenth to Mattithiah, he, his sons, and his brethren, were twelve:
1CHR|25|22|The fifteenth to Jeremoth, he, his sons, and his brethren, were twelve:
1CHR|25|23|The sixteenth to Hananiah, he, his sons, and his brethren, were twelve:
1CHR|25|24|The seventeenth to Joshbekashah, he, his sons, and his brethren, were twelve:
1CHR|25|25|The eighteenth to Hanani, he, his sons, and his brethren, were twelve:
1CHR|25|26|The nineteenth to Mallothi, he, his sons, and his brethren, were twelve:
1CHR|25|27|The twentieth to Eliathah, he, his sons, and his brethren, were twelve:
1CHR|25|28|The one and twentieth to Hothir, he, his sons, and his brethren, were twelve:
1CHR|25|29|The two and twentieth to Giddalti, he, his sons, and his brethren, were twelve:
1CHR|25|30|The three and twentieth to Mahazioth, he, his sons, and his brethren, were twelve:
1CHR|25|31|The four and twentieth to Romamtiezer, he, his sons, and his brethren, were twelve.
1CHR|26|1|Concerning the divisions of the porters: Of the Korhites was Meshelemiah the son of Kore, of the sons of Asaph.
1CHR|26|2|And the sons of Meshelemiah were, Zechariah the firstborn, Jediael the second, Zebadiah the third, Jathniel the fourth,
1CHR|26|3|Elam the fifth, Jehohanan the sixth, Elioenai the seventh.
1CHR|26|4|Moreover the sons of Obededom were, Shemaiah the firstborn, Jehozabad the second, Joah the third, and Sacar the fourth, and Nethaneel the fifth.
1CHR|26|5|Ammiel the sixth, Issachar the seventh, Peulthai the eighth: for God blessed him.
1CHR|26|6|Also unto Shemaiah his son were sons born, that ruled throughout the house of their father: for they were mighty men of valor.
1CHR|26|7|The sons of Shemaiah; Othni, and Rephael, and Obed, Elzabad, whose brethren were strong men, Elihu, and Semachiah.
1CHR|26|8|All these of the sons of Obededom: they and their sons and their brethren, able men for strength for the service, were threescore and two of Obededom.
1CHR|26|9|And Meshelemiah had sons and brethren, strong men, eighteen.
1CHR|26|10|Also Hosah, of the children of Merari, had sons; Simri the chief, (for though he was not the firstborn, yet his father made him the chief;)
1CHR|26|11|Hilkiah the second, Tebaliah the third, Zechariah the fourth: all the sons and brethren of Hosah were thirteen.
1CHR|26|12|Among these were the divisions of the porters, even among the chief men, having wards one against another, to minister in the house of the LORD.
1CHR|26|13|And they cast lots, as well the small as the great, according to the house of their fathers, for every gate.
1CHR|26|14|And the lot eastward fell to Shelemiah. Then for Zechariah his son, a wise counselor, they cast lots; and his lot came out northward.
1CHR|26|15|To Obededom southward; and to his sons the house of Asuppim.
1CHR|26|16|To Shuppim and Hosah the lot came forth westward, with the gate Shallecheth, by the causeway of the going up, ward against ward.
1CHR|26|17|Eastward were six Levites, northward four a day, southward four a day, and toward Asuppim two and two.
1CHR|26|18|At Parbar westward, four at the causeway, and two at Parbar.
1CHR|26|19|These are the divisions of the porters among the sons of Kore, and among the sons of Merari.
1CHR|26|20|And of the Levites, Ahijah was over the treasures of the house of God, and over the treasures of the dedicated things.
1CHR|26|21|As concerning the sons of Laadan; the sons of the Gershonite Laadan, chief fathers, even of Laadan the Gershonite, were Jehieli.
1CHR|26|22|The sons of Jehieli; Zetham, and Joel his brother, which were over the treasures of the house of the LORD.
1CHR|26|23|Of the Amramites, and the Izharites, the Hebronites, and the Uzzielites:
1CHR|26|24|And Shebuel the son of Gershom, the son of Moses, was ruler of the treasures.
1CHR|26|25|And his brethren by Eliezer; Rehabiah his son, and Jeshaiah his son, and Joram his son, and Zichri his son, and Shelomith his son.
1CHR|26|26|Which Shelomith and his brethren were over all the treasures of the dedicated things, which David the king, and the chief fathers, the captains over thousands and hundreds, and the captains of the host, had dedicated.
1CHR|26|27|Out of the spoils won in battles did they dedicate to maintain the house of the LORD.
1CHR|26|28|And all that Samuel the seer, and Saul the son of Kish, and Abner the son of Ner, and Joab the son of Zeruiah, had dedicated; and whosoever had dedicated any thing, it was under the hand of Shelomith, and of his brethren.
1CHR|26|29|Of the Izharites, Chenaniah and his sons were for the outward business over Israel, for officers and judges.
1CHR|26|30|And of the Hebronites, Hashabiah and his brethren, men of valor, a thousand and seven hundred, were officers among them of Israel on this side Jordan westward in all the business of the LORD, and in the service of the king.
1CHR|26|31|Among the Hebronites was Jerijah the chief, even among the Hebronites, according to the generations of his fathers. In the fortieth year of the reign of David they were sought for, and there were found among them mighty men of valor at Jazer of Gilead.
1CHR|26|32|And his brethren, men of valor, were two thousand and seven hundred chief fathers, whom king David made rulers over the Reubenites, the Gadites, and the half tribe of Manasseh, for every matter pertaining to God, and affairs of the king.
1CHR|27|1|Now the children of Israel after their number, to wit, the chief fathers and captains of thousands and hundreds, and their officers that served the king in any matter of the courses, which came in and went out month by month throughout all the months of the year, of every course were twenty and four thousand.
1CHR|27|2|Over the first course for the first month was Jashobeam the son of Zabdiel: and in his course were twenty and four thousand.
1CHR|27|3|Of the children of Perez was the chief of all the captains of the host for the first month.
1CHR|27|4|And over the course of the second month was Dodai an Ahohite, and of his course was Mikloth also the ruler: in his course likewise were twenty and four thousand.
1CHR|27|5|The third captain of the host for the third month was Benaiah the son of Jehoiada, a chief priest: and in his course were twenty and four thousand.
1CHR|27|6|This is that Benaiah, who was mighty among the thirty, and above the thirty: and in his course was Ammizabad his son.
1CHR|27|7|The fourth captain for the fourth month was Asahel the brother of Joab, and Zebadiah his son after him: and in his course were twenty and four thousand.
1CHR|27|8|The fifth captain for the fifth month was Shamhuth the Izrahite: and in his course were twenty and four thousand.
1CHR|27|9|The sixth captain for the sixth month was Ira the son of Ikkesh the Tekoite: and in his course were twenty and four thousand.
1CHR|27|10|The seventh captain for the seventh month was Helez the Pelonite, of the children of Ephraim: and in his course were twenty and four thousand.
1CHR|27|11|The eighth captain for the eighth month was Sibbecai the Hushathite, of the Zarhites: and in his course were twenty and four thousand.
1CHR|27|12|The ninth captain for the ninth month was Abiezer the Anetothite, of the Benjamites: and in his course were twenty and four thousand.
1CHR|27|13|The tenth captain for the tenth month was Maharai the Netophathite, of the Zarhites: and in his course were twenty and four thousand.
1CHR|27|14|The eleventh captain for the eleventh month was Benaiah the Pirathonite, of the children of Ephraim: and in his course were twenty and four thousand.
1CHR|27|15|The twelfth captain for the twelfth month was Heldai the Netophathite, of Othniel: and in his course were twenty and four thousand.
1CHR|27|16|Furthermore over the tribes of Israel: the ruler of the Reubenites was Eliezer the son of Zichri: of the Simeonites, Shephatiah the son of Maachah:
1CHR|27|17|Of the Levites, Hashabiah the son of Kemuel: of the Aaronites, Zadok:
1CHR|27|18|Of Judah, Elihu, one of the brethren of David: of Issachar, Omri the son of Michael:
1CHR|27|19|Of Zebulun, Ishmaiah the son of Obadiah: of Naphtali, Jerimoth the son of Azriel:
1CHR|27|20|Of the children of Ephraim, Hoshea the son of Azaziah: of the half tribe of Manasseh, Joel the son of Pedaiah:
1CHR|27|21|Of the half tribe of Manasseh in Gilead, Iddo the son of Zechariah: of Benjamin, Jaasiel the son of Abner:
1CHR|27|22|Of Dan, Azareel the son of Jeroham. These were the princes of the tribes of Israel.
1CHR|27|23|But David took not the number of them from twenty years old and under: because the LORD had said he would increase Israel like to the stars of the heavens.
1CHR|27|24|Joab the son of Zeruiah began to number, but he finished not, because there fell wrath for it against Israel; neither was the number put in the account of the chronicles of king David.
1CHR|27|25|And over the king's treasures was Azmaveth the son of Adiel: and over the storehouses in the fields, in the cities, and in the villages, and in the castles, was Jehonathan the son of Uzziah:
1CHR|27|26|And over them that did the work of the field for tillage of the ground was Ezri the son of Chelub:
1CHR|27|27|And over the vineyards was Shimei the Ramathite: over the increase of the vineyards for the wine cellars was Zabdi the Shiphmite:
1CHR|27|28|And over the olive trees and the sycamore trees that were in the low plains was Baalhanan the Gederite: and over the cellars of oil was Joash:
1CHR|27|29|And over the herds that fed in Sharon was Shitrai the Sharonite: and over the herds that were in the valleys was Shaphat the son of Adlai:
1CHR|27|30|Over the camels also was Obil the Ishmaelite: and over the asses was Jehdeiah the Meronothite:
1CHR|27|31|And over the flocks was Jaziz the Hagerite. All these were the rulers of the substance which was king David's.
1CHR|27|32|Also Jonathan David's uncle was a counselor, a wise man, and a scribe: and Jehiel the son of Hachmoni was with the king's sons:
1CHR|27|33|And Ahithophel was the king's counselor: and Hushai the Archite was the king's companion:
1CHR|27|34|And after Ahithophel was Jehoiada the son of Benaiah, and Abiathar: and the general of the king's army was Joab.
1CHR|28|1|And David assembled all the princes of Israel, the princes of the tribes, and the captains of the companies that ministered to the king by course, and the captains over the thousands, and captains over the hundreds, and the stewards over all the substance and possession of the king, and of his sons, with the officers, and with the mighty men, and with all the valiant men, unto Jerusalem.
1CHR|28|2|Then David the king stood up upon his feet, and said, Hear me, my brethren, and my people: As for me, I had in mine heart to build an house of rest for the ark of the covenant of the LORD, and for the footstool of our God, and had made ready for the building:
1CHR|28|3|But God said unto me, Thou shalt not build an house for my name, because thou hast been a man of war, and hast shed blood.
1CHR|28|4|Howbeit the LORD God of Israel chose me before all the house of my father to be king over Israel for ever: for he hath chosen Judah to be the ruler; and of the house of Judah, the house of my father; and among the sons of my father he liked me to make me king over all Israel:
1CHR|28|5|And of all my sons, (for the LORD hath given me many sons,) he hath chosen Solomon my son to sit upon the throne of the kingdom of the LORD over Israel.
1CHR|28|6|And he said unto me, Solomon thy son, he shall build my house and my courts: for I have chosen him to be my son, and I will be his father.
1CHR|28|7|Moreover I will establish his kingdom for ever, if he be constant to do my commandments and my judgments, as at this day.
1CHR|28|8|Now therefore in the sight of all Israel the congregation of the LORD, and in the audience of our God, keep and seek for all the commandments of the LORD your God: that ye may possess this good land, and leave it for an inheritance for your children after you for ever.
1CHR|28|9|And thou, Solomon my son, know thou the God of thy father, and serve him with a perfect heart and with a willing mind: for the LORD searcheth all hearts, and understandeth all the imaginations of the thoughts: if thou seek him, he will be found of thee; but if thou forsake him, he will cast thee off for ever.
1CHR|28|10|Take heed now; for the LORD hath chosen thee to build an house for the sanctuary: be strong, and do it.
1CHR|28|11|Then David gave to Solomon his son the pattern of the porch, and of the houses thereof, and of the treasuries thereof, and of the upper chambers thereof, and of the inner parlors thereof, and of the place of the mercy seat,
1CHR|28|12|And the pattern of all that he had by the spirit, of the courts of the house of the LORD, and of all the chambers round about, of the treasuries of the house of God, and of the treasuries of the dedicated things:
1CHR|28|13|Also for the courses of the priests and the Levites, and for all the work of the service of the house of the LORD, and for all the vessels of service in the house of the LORD.
1CHR|28|14|He gave of gold by weight for things of gold, for all instruments of all manner of service; silver also for all instruments of silver by weight, for all instruments of every kind of service:
1CHR|28|15|Even the weight for the candlesticks of gold, and for their lamps of gold, by weight for every candlestick, and for the lamps thereof: and for the candlesticks of silver by weight, both for the candlestick, and also for the lamps thereof, according to the use of every candlestick.
1CHR|28|16|And by weight he gave gold for the tables of shewbread, for every table; and likewise silver for the tables of silver:
1CHR|28|17|Also pure gold for the fleshhooks, and the bowls, and the cups: and for the golden basins he gave gold by weight for every basin; and likewise silver by weight for every basin of silver:
1CHR|28|18|And for the altar of incense refined gold by weight; and gold for the pattern of the chariot of the cherubim, that spread out their wings, and covered the ark of the covenant of the LORD.
1CHR|28|19|All this, said David, the LORD made me understand in writing by his hand upon me, even all the works of this pattern.
1CHR|28|20|And David said to Solomon his son, Be strong and of good courage, and do it: fear not, nor be dismayed: for the LORD God, even my God, will be with thee; he will not fail thee, nor forsake thee, until thou hast finished all the work for the service of the house of the LORD.
1CHR|28|21|And, behold, the courses of the priests and the Levites, even they shall be with thee for all the service of the house of God: and there shall be with thee for all manner of workmanship every willing skillful man, for any manner of service: also the princes and all the people will be wholly at thy commandment.
1CHR|29|1|Furthermore David the king said unto all the congregation, Solomon my son, whom alone God hath chosen, is yet young and tender, and the work is great: for the palace is not for man, but for the LORD God.
1CHR|29|2|Now I have prepared with all my might for the house of my God the gold for things to be made of gold, and the silver for things of silver, and the brass for things of brass, the iron for things of iron, and wood for things of wood; onyx stones, and stones to be set, glistering stones, and of divers colors, and all manner of precious stones, and marble stones in abundance.
1CHR|29|3|Moreover, because I have set my affection to the house of my God, I have of mine own proper good, of gold and silver, which I have given to the house of my God, over and above all that I have prepared for the holy house.
1CHR|29|4|Even three thousand talents of gold, of the gold of Ophir, and seven thousand talents of refined silver, to overlay the walls of the houses withal:
1CHR|29|5|The gold for things of gold, and the silver for things of silver, and for all manner of work to be made by the hands of artificers. And who then is willing to consecrate his service this day unto the LORD?
1CHR|29|6|Then the chief of the fathers and princes of the tribes of Israel and the captains of thousands and of hundreds, with the rulers of the king's work, offered willingly,
1CHR|29|7|And gave for the service of the house of God of gold five thousand talents and ten thousand drams, and of silver ten thousand talents, and of brass eighteen thousand talents, and one hundred thousand talents of iron.
1CHR|29|8|And they with whom precious stones were found gave them to the treasure of the house of the LORD, by the hand of Jehiel the Gershonite.
1CHR|29|9|Then the people rejoiced, for that they offered willingly, because with perfect heart they offered willingly to the LORD: and David the king also rejoiced with great joy.
1CHR|29|10|Wherefore David blessed the LORD before all the congregation: and David said, Blessed be thou, LORD God of Israel our father, for ever and ever.
1CHR|29|11|Thine, O LORD is the greatness, and the power, and the glory, and the victory, and the majesty: for all that is in the heaven and in the earth is thine; thine is the kingdom, O LORD, and thou art exalted as head above all.
1CHR|29|12|Both riches and honor come of thee, and thou reignest over all; and in thine hand is power and might; and in thine hand it is to make great, and to give strength unto all.
1CHR|29|13|Now therefore, our God, we thank thee, and praise thy glorious name.
1CHR|29|14|But who am I, and what is my people, that we should be able to offer so willingly after this sort? for all things come of thee, and of thine own have we given thee.
1CHR|29|15|For we are strangers before thee, and sojourners, as were all our fathers: our days on the earth are as a shadow, and there is none abiding.
1CHR|29|16|O LORD our God, all this store that we have prepared to build thee an house for thine holy name cometh of thine hand, and is all thine own.
1CHR|29|17|I know also, my God, that thou triest the heart, and hast pleasure in uprightness. As for me, in the uprightness of mine heart I have willingly offered all these things: and now have I seen with joy thy people, which are present here, to offer willingly unto thee.
1CHR|29|18|O LORD God of Abraham, Isaac, and of Israel, our fathers, keep this for ever in the imagination of the thoughts of the heart of thy people, and prepare their heart unto thee:
1CHR|29|19|And give unto Solomon my son a perfect heart, to keep thy commandments, thy testimonies, and thy statutes, and to do all these things, and to build the palace, for the which I have made provision.
1CHR|29|20|And David said to all the congregation, Now bless the LORD your God. And all the congregation blessed the LORD God of their fathers, and bowed down their heads, and worshipped the LORD, and the king.
1CHR|29|21|And they sacrificed sacrifices unto the LORD, and offered burnt offerings unto the LORD, on the morrow after that day, even a thousand bullocks, a thousand rams, and a thousand lambs, with their drink offerings, and sacrifices in abundance for all Israel:
1CHR|29|22|And did eat and drink before the LORD on that day with great gladness. And they made Solomon the son of David king the second time, and anointed him unto the LORD to be the chief governor, and Zadok to be priest.
1CHR|29|23|Then Solomon sat on the throne of the LORD as king instead of David his father, and prospered; and all Israel obeyed him.
1CHR|29|24|And all the princes, and the mighty men, and all the sons likewise of king David, submitted themselves unto Solomon the king.
1CHR|29|25|And the LORD magnified Solomon exceedingly in the sight of all Israel, and bestowed upon him such royal majesty as had not been on any king before him in Israel.
1CHR|29|26|Thus David the son of Jesse reigned over all Israel.
1CHR|29|27|And the time that he reigned over Israel was forty years; seven years reigned he in Hebron, and thirty and three years reigned he in Jerusalem.
1CHR|29|28|And he died in a good old age, full of days, riches, and honor: and Solomon his son reigned in his stead.
1CHR|29|29|Now the acts of David the king, first and last, behold, they are written in the book of Samuel the seer, and in the book of Nathan the prophet, and in the book of Gad the seer,
1CHR|29|30|With all his reign and his might, and the times that went over him, and over Israel, and over all the kingdoms of the countries.
