NAH|1|1|Пророчество о Ниневии; книга видений Наума Елкосеянина.
NAH|1|2|Господь есть Бог ревнитель и мститель; мститель Господь и страшен в гневе: мстит Господь врагам Своим и не пощадит противников Своих.
NAH|1|3|Господь долготерпелив и велик могуществом, и не оставляет без наказания; в вихре и в буре шествие Господа, облако – пыль от ног Его.
NAH|1|4|Запретит Он морю, и оно высыхает, и все реки иссякают; вянет Васан и Кармил, и блекнет цвет на Ливане.
NAH|1|5|Горы трясутся пред Ним, и холмы тают, и земля колеблется пред лицем Его, и вселенная и все живущие в ней.
NAH|1|6|Пред негодованием Его кто устоит? И кто стерпит пламя гнева Его? Гнев Его разливается как огонь; скалы распадаются пред Ним.
NAH|1|7|Благ Господь, убежище в день скорби, и знает надеющихся на Него.
NAH|1|8|Но всепотопляющим наводнением разрушит до основания [Ниневию], и врагов Его постигнет мрак.
NAH|1|9|Что умышляете вы против Господа? Он совершит истребление, и бедствие уже не повторится,
NAH|1|10|ибо сплетшиеся между собою как терновник и упившиеся как пьяницы, они пожраны будут совершенно, как сухая солома.
NAH|1|11|Из тебя произошел умысливший злое против Господа, составивший совет нечестивый.
NAH|1|12|Так говорит Господь: хотя они безопасны и многочисленны, но они будут посечены и исчезнут; а тебя, хотя Я отягощал, более не буду отягощать.
NAH|1|13|И ныне Я сокрушу ярмо его, лежащее на тебе, и узы твои разорву.
NAH|1|14|А о тебе, [Ассур], Господь определил: не будет более семени с твоим именем; из дома бога твоего истреблю истуканов и кумиров; приготовлю тебе в нем могилу, потому что ты будешь в презрении.
NAH|1|15|Вот, на горах – стопы благовестника, возвещающего мир: празднуй, Иудея, праздники твои, исполняй обеты твои, ибо не будет более проходить по тебе нечестивый: он совсем уничтожен.
NAH|2|1|Поднимается на тебя разрушитель: охраняй твердыни, стереги дорогу, укрепи чресла, собирайся с силами.
NAH|2|2|Ибо восстановит Господь величие Иакова, как величие Израиля, потому что опустошили их опустошители и виноградные ветви их истребили.
NAH|2|3|Щит героев его красен; воины его в одеждах багряных; огнем сверкают колесницы в день приготовления к бою, и лес копьев волнуется.
NAH|2|4|По улицам несутся колесницы, гремят на площадях; блеск от них, как от огня; сверкают, как молния.
NAH|2|5|Он вызывает храбрых своих, но они спотыкаются на ходу своем; поспешают на стены города, но осада уже устроена.
NAH|2|6|Речные ворота отворяются, и дворец разрушается.
NAH|2|7|Решено: она будет обнажена и отведена в плен, и рабыни ее будут стонать как голуби, ударяя себя в грудь.
NAH|2|8|Ниневия со времени существования своего была как пруд, полный водою, а они бегут. "Стойте, стойте!" Но никто не оглядывается.
NAH|2|9|Расхищайте серебро, расхищайте золото! нет конца запасам всякой драгоценной утвари.
NAH|2|10|Разграблена, опустошена и разорена она, – и тает сердце, колени трясутся; у всех в чреслах сильная боль, и лица у всех потемнели.
NAH|2|11|Где теперь логовище львов и то пастбище для львенков, по которому ходил лев, львица и львенок, и никто не пугал их, –
NAH|2|12|лев, похищающий для насыщения щенков своих, и задушающий для львиц своих, и наполняющий добычею пещеры свои и логовища свои похищенным?
NAH|2|13|Вот, Я – на тебя! говорит Господь Саваоф. И сожгу в дыму колесницы твои, и меч пожрет львенков твоих, и истреблю с земли добычу твою, и не будет более слышим голос послов твоих.
NAH|3|1|Горе городу кровей! весь он полон обмана и убийства; не прекращается в нем грабительство.
NAH|3|2|Слышны хлопанье бича и стук крутящихся колес, ржание коня и грохот скачущей колесницы.
NAH|3|3|Несется конница, сверкает меч и блестят копья; убитых множество и груды трупов: нет конца трупам, спотыкаются о трупы их.
NAH|3|4|Это – за многие блудодеяния развратницы приятной наружности, искусной в чародеянии, которая блудодеяниями своими продает народы и чарованиями своими – племена.
NAH|3|5|Вот, Я – на тебя! говорит Господь Саваоф. И подниму на лице твое края одежды твоей и покажу народам наготу твою и царствам срамоту твою.
NAH|3|6|И забросаю тебя мерзостями, сделаю тебя презренною и выставлю тебя на позор.
NAH|3|7|И будет то, что всякий, увидев тебя, побежит от тебя и скажет: "разорена Ниневия! Кто пожалеет о ней? где найду я утешителей для тебя?"
NAH|3|8|Разве ты лучше Но–Аммона, находящегося между реками, окруженного водою, которого вал было море, и море служило стеною его?
NAH|3|9|Ефиопия и Египет с бесчисленным множеством других служили ему подкреплением; Копты и Ливийцы приходили на помощь тебе.
NAH|3|10|Но и он переселен, пошел в плен; даже и младенцы его разбиты на перекрестках всех улиц, а о знатных его бросали жребий, и все вельможи его окованы цепями.
NAH|3|11|Так и ты – опьянеешь и скроешься; так и ты будешь искать защиты от неприятеля.
NAH|3|12|Все укрепления твои подобны смоковнице со спелыми плодами: если тряхнуть их, то они упадут прямо в рот желающего есть.
NAH|3|13|Вот, и народ твой, как женщины у тебя: врагам твоим настежь отворятся ворота земли твоей, огонь пожрет запоры твои.
NAH|3|14|Начерпай воды на время осады; укрепляй крепости твои; пойди в грязь, топчи глину, исправь печь для обжигания кирпичей.
NAH|3|15|Там пожрет тебя огонь, посечет тебя меч, поест тебя как гусеница, хотя бы ты умножился как гусеница, умножился как саранча.
NAH|3|16|Купцов у тебя стало более, нежели звезд на небе; но эта саранча рассеется и улетит.
NAH|3|17|Князья твои – как саранча, и военачальники твои – как рои мошек, которые во время холода гнездятся в щелях [стен], и когда взойдет солнце, то разлетаются, и не узнаешь места, где они были.
NAH|3|18|Спят пастыри твои, царь Ассирийский, покоятся вельможи твои; народ твой рассеялся по горам, и некому собрать его.
NAH|3|19|Нет врачевства для раны твоей, болезненна язва твоя. Все, услышавшие весть о тебе, будут рукоплескать о тебе, ибо на кого не простиралась беспрестанно злоба твоя?
