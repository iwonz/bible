PHLM|1|1|Paul, a prisoner of Jesus Christ, and Timothy our brother, unto Philemon our dearly beloved, and fellowlabourer,
PHLM|1|2|And to our beloved Apphia, and Archippus our fellowsoldier, and to the church in thy house:
PHLM|1|3|Grace to you, and peace, from God our Father and the Lord Jesus Christ.
PHLM|1|4|I thank my God, making mention of thee always in my prayers,
PHLM|1|5|Hearing of thy love and faith, which thou hast toward the Lord Jesus, and toward all saints;
PHLM|1|6|That the communication of thy faith may become effectual by the acknowledging of every good thing which is in you in Christ Jesus.
PHLM|1|7|For we have great joy and consolation in thy love, because the bowels of the saints are refreshed by thee, brother.
PHLM|1|8|Wherefore, though I might be much bold in Christ to enjoin thee that which is convenient,
PHLM|1|9|Yet for love's sake I rather beseech thee, being such an one as Paul the aged, and now also a prisoner of Jesus Christ.
PHLM|1|10|I beseech thee for my son Onesimus, whom I have begotten in my bonds:
PHLM|1|11|Which in time past was to thee unprofitable, but now profitable to thee and to me:
PHLM|1|12|Whom I have sent again: thou therefore receive him, that is, mine own bowels:
PHLM|1|13|Whom I would have retained with me, that in thy stead he might have ministered unto me in the bonds of the gospel:
PHLM|1|14|But without thy mind would I do nothing; that thy benefit should not be as it were of necessity, but willingly.
PHLM|1|15|For perhaps he therefore departed for a season, that thou shouldest receive him for ever;
PHLM|1|16|Not now as a servant, but above a servant, a brother beloved, specially to me, but how much more unto thee, both in the flesh, and in the Lord?
PHLM|1|17|If thou count me therefore a partner, receive him as myself.
PHLM|1|18|If he hath wronged thee, or oweth thee ought, put that on mine account;
PHLM|1|19|I Paul have written it with mine own hand, I will repay it: albeit I do not say to thee how thou owest unto me even thine own self besides.
PHLM|1|20|Yea, brother, let me have joy of thee in the Lord: refresh my bowels in the Lord.
PHLM|1|21|Having confidence in thy obedience I wrote unto thee, knowing that thou wilt also do more than I say.
PHLM|1|22|But withal prepare me also a lodging: for I trust that through your prayers I shall be given unto you.
PHLM|1|23|There salute thee Epaphras, my fellowprisoner in Christ Jesus;
PHLM|1|24|Marcus, Aristarchus, Demas, Lucas, my fellowlabourers.
PHLM|1|25|The grace of our Lord Jesus Christ be with your spirit. Amen.
