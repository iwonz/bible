ECCL|1|1|在 耶路撒冷 作王、 大卫 的儿子、传道者的言语。
ECCL|1|2|传道者说：虚空的虚空， 虚空的虚空，全是虚空。
ECCL|1|3|人一切的劳碌， 就是他在日光之下的劳碌，有什么益处呢？
ECCL|1|4|一代过去，一代又来， 地却永远长存。
ECCL|1|5|太阳上升，太阳下落， 急归所出之地。
ECCL|1|6|风往南刮，又向北转， 不停旋转，绕回原路。
ECCL|1|7|江河都往海里流，海却不满； 江河从何处流，仍归回原处。
ECCL|1|8|万事令人厌倦， 人不能说尽。 眼看，看不饱； 耳听，听不足。
ECCL|1|9|已有的事，后必再有； 已行的事，后必再行。 日光之下并无新事。
ECCL|1|10|有一件事人指着说：“看，这是新的！” 它在我们以前的世代早已有了。
ECCL|1|11|已过的事，无人记念； 将来的事，后来的人也不记念。
ECCL|1|12|我传道者在 耶路撒冷 作过 以色列 的王。
ECCL|1|13|我用智慧专心探寻、考察天下所发生的一切事：上帝给世人何等沉重的担子，使他们在其中劳苦！
ECCL|1|14|我见日光之下所发生的一切事，看哪，全是虚空，全是捕风。
ECCL|1|15|弯曲的，不能变直； 缺乏的，不计其数。
ECCL|1|16|我心里说：“看哪，我大有智慧，胜过在我以前所有统治 耶路撒冷 的人；我的心也多经历智慧和知识的事。”
ECCL|1|17|我专心想要明白智慧，想要明白狂妄与愚昧，方知这也是捕风。
ECCL|1|18|因为多有智慧，就多有愁烦； 增加知识，就增加忧伤。
ECCL|2|1|我心里说：“来吧，让我用喜乐试试你，使你享福！”看哪，这也是虚空。
ECCL|2|2|论嬉笑，我说：“这是狂妄。”论享乐，“这有什么用呢？”
ECCL|2|3|我心以智慧引导我，我心里探究，如何用酒使身体舒畅，如何抓住愚昧，直等我看明世人在天下短暂一生中，当行何事为美。
ECCL|2|4|我大兴土木，为自己建造房屋，栽葡萄园，
ECCL|2|5|修造庭园和公园，在其中栽种各样果树，
ECCL|2|6|挖造水池，用以灌溉林中的幼树。
ECCL|2|7|我买了仆婢，也有生在家中的仆婢；又有许多牛群羊群，胜过我以前所有在 耶路撒冷 的人。
ECCL|2|8|我为自己积蓄金银，搜集各君王、各省份的财宝；又为自己得男女歌手和世人所喜爱的物，以及一个又一个的妃嫔。
ECCL|2|9|这样，我就日渐昌盛，胜过我以前所有在 耶路撒冷 的人。我的智慧仍然存留。
ECCL|2|10|凡我眼所求的，我没有克制它；我心所乐的，我没有不享受。因我的心要为一切的劳碌快乐，这是我从一切劳碌中所得的报偿 。
ECCL|2|11|后来，我回顾我手所经营的一切和我劳碌所做的工。看哪，全是虚空，全是捕风；在日光之下毫无益处。
ECCL|2|12|我转而回顾智慧、狂妄和愚昧。在王以后来的人又如何呢？不过做先前所做的就是了。
ECCL|2|13|于是我看出智慧胜过愚昧，如同光明胜过黑暗。
ECCL|2|14|智慧人的眼目光明 ，愚昧人却在黑暗里行。但我知道他们都有相同的遭遇。
ECCL|2|15|我心里就说：“愚昧人所遇见的，我也一样遇见，那么我何必更有智慧呢？”我心里说：“这也是虚空。”
ECCL|2|16|智慧人和愚昧人一样，不会长久被人记念，因为日后都被遗忘。可叹！智慧人和愚昧人都一样会死亡。
ECCL|2|17|于是我恨恶生命，因为在日光之下所发生的事我都以为烦恼，全是虚空，全是捕风。
ECCL|2|18|我恨恶一切的劳碌，就是我在日光之下所劳碌的，因为我所得的必须留给我以后的人。
ECCL|2|19|那人是智慧是愚昧，谁能知道呢？他竟要掌管我在日光之下用智慧劳碌所得的。这也是虚空。
ECCL|2|20|我转想我在日光之下所劳碌的一切工作，心就绝望。
ECCL|2|21|因为有人用智慧、知识、灵巧劳碌工作，所得来的却要遗留给未曾劳碌的人作产业。这也是虚空，大大不幸。
ECCL|2|22|人一切的劳碌操心，就是他在日光之下所劳碌的，又得着了什么呢？
ECCL|2|23|他日日忧虑，他的劳苦成为愁烦，连夜间心也不得休息。这也是虚空。
ECCL|2|24|难道一个人有吃有喝，且在劳碌中享福，不是福气吗？我看这也是出于上帝的手。
ECCL|2|25|论到吃用、享福，谁能胜过我呢？
ECCL|2|26|上帝喜爱谁，就给谁智慧、知识和喜乐；惟有罪人，上帝使他劳苦，将他所储藏、所堆积的归给上帝所喜爱的人。这也是虚空，也是捕风。
ECCL|3|1|凡事都有定期， 天下每一事务都有定时。
ECCL|3|2|生有时，死有时； 栽种有时，拔出 有时；
ECCL|3|3|杀戮有时，医治有时； 拆毁有时，建造有时；
ECCL|3|4|哭有时，笑有时； 哀恸有时，跳舞有时；
ECCL|3|5|丢石头有时，捡石头有时； 怀抱有时，不抱有时；
ECCL|3|6|寻找有时，失落有时； 保存有时，抛弃有时；
ECCL|3|7|撕裂有时，缝补有时； 沉默有时，说话有时；
ECCL|3|8|喜爱有时，恨恶有时； 战争有时，和平有时。
ECCL|3|9|这样，做事的人在他所劳碌的事上得到什么益处呢？
ECCL|3|10|我观看上帝给世人的担子，使他们在其中劳苦：
ECCL|3|11|上帝造万物，各按其时成为美好，又将永恒安放在世人心里；然而上帝从始至终的作为，人不能测透。
ECCL|3|12|我知道，人除了终身喜乐纳福，没有一件幸福的事。
ECCL|3|13|并且人人吃喝，在他的一切劳碌中享福，这也是上帝的赏赐。
ECCL|3|14|我知道上帝所做的都必存到永远；无所增添，无所减少。上帝这样做，是要人在他面前存敬畏的心。
ECCL|3|15|现今的事以前就有了，将来的事也早已有了，并且上帝使已过的事重新再来 。
ECCL|3|16|我又见日光之下，应有公平之处有奸恶，应有公义之处也有奸恶。
ECCL|3|17|我心里说：“上帝必审判义人和恶人，因为在那里，各样事务，一切工作，都有定时。”
ECCL|3|18|我心里说：“为世人的缘故，上帝考验他们，让他们看见自己不过像走兽一样。”
ECCL|3|19|因为世人遭遇的，走兽也遭遇，所遭遇的都一样：这个怎样死，那个也怎样死，他们都有一样的气息。人不能强于走兽，全是虚空；
ECCL|3|20|都归一处，都是出于尘土，也都归于尘土。
ECCL|3|21|谁知道人的气息是往上升，走兽的气息是下入地呢？
ECCL|3|22|总而言之，人能够在他经营的事上喜乐，是最好不过了，因为这是他应得的报偿。他身后的事谁能领他回来看呢？
ECCL|4|1|我转而观看日光之下所发生的一切欺压之事。看哪，受欺压的流泪，无人安慰；欺压他们的有权势，也无人安慰。
ECCL|4|2|因此，我赞叹那已死的死人，胜过那还活着的活人。
ECCL|4|3|但那尚未出生，就是未曾见过日光之下所发生之恶事的，比这两种人更幸福。
ECCL|4|4|我见人因彼此嫉妒而有一切的劳碌和各样工作的成就，这也是虚空，也是捕风。
ECCL|4|5|愚昧人抱着双臂， 自食其肉。
ECCL|4|6|一掌满满而得享安静， 胜过两掌满满而劳碌捕风。
ECCL|4|7|我转而观看日光之下有一件虚空的事：
ECCL|4|8|有人孤单无双，无子无兄弟，竟劳碌不息，眼目也不以财富为满足。他说：“我劳碌，自己却不享福，到底是为了谁呢？”这也是虚空，是极沉重的担子。
ECCL|4|9|两个人总比一个人好，他们劳碌同得美好的报偿。
ECCL|4|10|若是跌倒，这人可以扶起他的同伴；倘若孤身跌倒，没有别人扶起他来，这人就有祸了。
ECCL|4|11|再者，二人同睡就都暖和，一人独睡怎能暖和呢？
ECCL|4|12|若遇敌攻击，孤身难挡，二人就能抵挡他；三股合成的绳子不易折断。
ECCL|4|13|贫穷而有智慧的年轻人，胜过年老不再纳谏的愚昧王，
ECCL|4|14|那人从监牢里出来作王，在国中原是出身贫寒。
ECCL|4|15|我见日光之下所有行走的活人，都跟随那年轻人，就是接续作王的那位。
ECCL|4|16|他的百姓，就是他所治理的众人，多得无数；但后来的人还是不喜欢他。这也是虚空，也是捕风。
ECCL|5|1|你到上帝的殿要谨慎你的脚步；近前听，胜过愚昧人献祭，他们不知道自己在作恶。
ECCL|5|2|在上帝面前你不可冒失开口，也不可心急发言；因为上帝在天上，你在地上，所以你的话语要少。
ECCL|5|3|事务多，令人做梦；话语多，显出愚昧。
ECCL|5|4|你向上帝许愿，还愿不可迟延，因他不喜欢愚昧人，你许的愿应当偿还。
ECCL|5|5|你许愿不还，不如不许。
ECCL|5|6|不可放任你的口使肉体犯罪，也不可在使者 面前说是错许了。为何使上帝因你的声音发怒，败坏你手所做的呢？
ECCL|5|7|多梦多言，其中多有虚空，你只要敬畏上帝。
ECCL|5|8|你若在一个地区看见穷人受欺压，公义公平被掠夺，不要因此惊奇；有一位高过居高位的在鉴察，在他们之上还有更高的。
ECCL|5|9|况且地的益处归众人，就是君王也受田地的供应。
ECCL|5|10|喜爱银子的，不因得银子满足；喜爱财富的，也不因得利益知足。这也是虚空。
ECCL|5|11|货物增添，吃的人也增添，物主得什么益处呢？不过眼看而已！
ECCL|5|12|劳碌的人不拘吃多吃少，睡得香甜；富人的丰足却不容他睡觉。
ECCL|5|13|我见日光之下有一件令人忧伤的祸患，就是财主积存财富，反害自己。
ECCL|5|14|他因遭遇不幸 ，财产尽失；他生了儿子，手里却一无所有。
ECCL|5|15|他怎样从母胎赤身而来，也必照样赤身而去；他所劳碌得来的，手中分毫不能带去。
ECCL|5|16|这是一件令人忧伤的祸患。他来的时候怎样，去的时候也必怎样。他为风劳碌有什么益处呢？
ECCL|5|17|并且他终身在黑暗中吃喝 ，多有烦恼、病痛和怒气。
ECCL|5|18|看哪，我所见为善为美的，就是人在上帝赐他一生的日子吃喝，享受日光之下劳碌得来的好处，因为这是他应得的报偿。
ECCL|5|19|而且，一个人蒙上帝赏赐财富与资产，又使他能享用，能获取自己当有的报偿 ，在他的劳碌中喜乐，这是上帝的赏赐。
ECCL|5|20|他不多思念自己一生的日子，因为上帝使他的心充满喜乐。
ECCL|6|1|我见日光之下有一件祸患重压在人身上，
ECCL|6|2|就是人蒙上帝赐他财富、资产和尊荣，以致他心里所愿的一样都不缺，只是上帝使他不能享用，反被外人享用。这是虚空，也是祸患。
ECCL|6|3|人若生一百个儿子，活许多岁数；他即使寿命很长，心里却不因福乐而满足，又不得埋葬；我说，那流掉的胎比他倒好。
ECCL|6|4|因为这胎虚虚而来，暗暗而去，名字被黑暗遮蔽，
ECCL|6|5|而且没有见过天日，什么都不知道，这胎比那人倒享安息。
ECCL|6|6|那人虽然活千年，再活千年，却不能享福；众人岂不都归同一个地方去吗？
ECCL|6|7|人的劳碌都为口腹，心里却不知足。
ECCL|6|8|智慧人比愚昧人有什么益处呢？困苦人在众人面前知道如何行，有什么益处呢？
ECCL|6|9|眼睛所看的比心里妄想的倒好。这也是虚空，也是捕风。
ECCL|6|10|先前所有的，早已起了名，人早知道人是如何的，不能与比自己强壮的相争。
ECCL|6|11|话语多，虚空也增多，这对人有什么益处呢？
ECCL|6|12|人一生虚度的日子，如影儿经过，谁知道什么才是对他有益呢？谁能告诉他身后在日光之下会发生什么事呢？
ECCL|7|1|名誉强如美好的膏油， 人死去的日子胜过他出生的日子。
ECCL|7|2|往丧家去， 强如往宴乐的家， 因为死是众人的结局， 活人必将这事放在心上。
ECCL|7|3|忧愁强如喜笑， 因为面带愁容，终必使心喜乐。
ECCL|7|4|智慧人的心在遭丧之家； 愚昧人的心在快乐之家。
ECCL|7|5|听智慧人的责备， 强如听愚昧人歌唱；
ECCL|7|6|因为愚昧人的笑声， 好像锅子下面烧荆棘的爆声， 这也是虚空。
ECCL|7|7|勒索使智慧人变为愚妄， 贿赂能败坏人的心。
ECCL|7|8|事情的终局强如它的起头； 存心忍耐的，胜过居心骄傲的。
ECCL|7|9|你的心不要急躁恼怒， 因为恼怒存在愚昧人的怀中。
ECCL|7|10|不要说： 为什么先前的日子强过现今的日子呢？ 你这样问不是出于智慧。
ECCL|7|11|智慧加上产业是美好的， 对见天日的人都有益处。
ECCL|7|12|因为智慧庇护人， 好像金钱庇护人一样； 智慧能保全智慧者的生命， 这就是知识的益处。
ECCL|7|13|你要观看上帝的作为， 谁能使他所弯曲的变直呢？
ECCL|7|14|顺利时要喜乐；患难时当思考。上帝使这两样都发生，因此，人不知将会发生什么事。
ECCL|7|15|在虚度的日子里，我见过各样的事情，义人在他的义中灭亡，恶人在他的恶中倒享长寿。
ECCL|7|16|不要行义过分，也不要过于自逞智慧，何必自取败亡呢？
ECCL|7|17|不要行恶过分，也不要为人愚昧，何必未到期而死呢？
ECCL|7|18|你持守这个，那个也不要松手才好。敬畏上帝的人，这一切都能兼得。
ECCL|7|19|智慧使拥有智慧的人比城中十个官长更有能力。
ECCL|7|20|其实世上没有行善而不犯罪的义人。
ECCL|7|21|人所说的话，你不要都放在心上，免得听见你的仆人诅咒你。
ECCL|7|22|因为你心里知道，自己也曾屡次诅咒别人。
ECCL|7|23|我曾用智慧试验这一切事，我说：“要得智慧。”智慧却离我远。
ECCL|7|24|万事之理遥不可及，太深奥，谁能测透呢？
ECCL|7|25|我转念，一心要知道，要考察，要寻求智慧和万事的来由，要知道邪恶为愚昧，愚昧为狂妄。
ECCL|7|26|我发现有一种妇人比死还苦毒：她本身是陷阱，她的心是罗网，手是锁链。凡蒙上帝喜爱的人必能躲开她；有罪的人却被她缠住了。
ECCL|7|27|传道者说：“你看，我考察一件又一件，为要寻求万事的来由，这是我所寻得的：
ECCL|7|28|我继续寻找，却未找到；一千当中，我找到一个男的，但在这一切当中，却找不到一个女的。
ECCL|7|29|你看，我所找到的只有一件，就是上帝造的人是正直的，但他们却寻出许多诡计。”
ECCL|8|1|谁如 智慧人呢？ 谁知道事情的解释呢？ 人的智慧使他的脸发光， 改变他脸上的暴戾之气 。
ECCL|8|2|我劝你 因上帝誓言的缘故，当遵守王的命令。
ECCL|8|3|不要急躁离开王的面前，不要固执行恶，因为他凡事都随自己心意而行。
ECCL|8|4|王的话本有权力，谁能对他说：“你在做什么？”
ECCL|8|5|凡遵守命令的，必不经历祸患；智慧人的心知道适当的时机和必经的过程。
ECCL|8|6|各样事务都有时机和过程，但人有苦难重压在身。
ECCL|8|7|他不知道将来的事，其实将来如何，谁能告诉他呢？
ECCL|8|8|没有人能掌握生命，将生命留住；也没有人有权力掌管死期。这场争战无人能免；邪恶也不能救那行邪恶的人。
ECCL|8|9|这一切我都见过，我专心考察日光之下所发生的一切事，有时这人管辖那人，令他受害。
ECCL|8|10|我见恶人埋葬；从前他们进出圣地，他们在城中的作为被人忘记。这也是虚空。
ECCL|8|11|判罪之后不立刻执行，所以世人满怀作恶的心思。
ECCL|8|12|罪人虽然作恶百次，倒享长寿；然而我也知道，福乐必临到敬畏上帝的人，就是在他面前心存敬畏的人。
ECCL|8|13|恶人却不得福乐，他的日子好像影儿不得长久，因为他不敬畏上帝。
ECCL|8|14|世上有一件虚空的事，就是义人所遭遇的，反而照恶人所做的；恶人所遭遇的，反而照义人所做的。我说，这也是虚空。
ECCL|8|15|我就称赞快乐，原来人在日光之下，最大的福气莫过于吃喝快乐；他在日光之下，上帝赐他一生的日子，要从劳碌中享受所得。
ECCL|8|16|我专心想要明白智慧，要观看世上所发生的事。有人昼夜不得阖眼睡觉。
ECCL|8|17|我观看上帝一切的作为，知道人不能探求日光之下所发生的事；任凭他费多少力探索，都找不出来，智慧人虽说他明白，仍不能找出来。
ECCL|9|1|我将这一切事放在心上，详细研究这些，就知道义人和智慧人，并他们的作为都在上帝手中；或是爱，或是恨，都在他们面前，但人不能知道。
ECCL|9|2|凡临到众人的际遇都一样：义人和恶人，好人 ，洁净的人和不洁净的人，献祭的和不献祭的，都一样。好人如何，罪人也如何；起誓的如何，怕起誓的也如何。
ECCL|9|3|在日光之下发生的一切事中有一件祸患，就是众人的际遇都一样，并且世人的心充满了恶；活着的时候心里狂妄，后来就归死人那里去了。
ECCL|9|4|与一切活人相连的，那人还有指望，因为活着的狗胜过死了的狮子。
ECCL|9|5|活着的人知道必死；死了的人毫无所知，也不再得赏赐，因为他们的名 已被遗忘。
ECCL|9|6|他们的爱，他们的恨，他们的嫉妒，早就消灭了。在日光之下所发生的一切事，他们永不再有份了。
ECCL|9|7|你只管欢欢喜喜吃你的饭，心中快乐喝你的酒，因为上帝已经悦纳你的作为。
ECCL|9|8|你的衣服要时时洁白，你头上也不要缺少膏油。
ECCL|9|9|在你一生虚空的日子，就是上帝赐你在日光之下虚空 的日子，当与你所爱的妻快活度日，因为那是你一生中在日光之下劳碌所得的报偿。
ECCL|9|10|凡你手所当做的事，要尽力去做；因为在你所必须去的阴间没有工作，没有谋算，没有知识，也没有智慧。
ECCL|9|11|我转而回顾日光之下，快跑的未必能赢，强壮的未必战胜，智慧的未必得粮食，聪明的未必得财富，有学问的未必得人喜悦，全在乎各人遇上的时候和机会。
ECCL|9|12|人不知道自己的定期。鱼被险恶的网圈住，鸟被罗网捉住，祸患的时刻忽然临到，世人陷在其中也是如此。
ECCL|9|13|我见日光之下有一样智慧，在我看来是伟大的，
ECCL|9|14|就是有一人口稀少的小城，遇大君王前来攻击，修筑营垒，将城围困。
ECCL|9|15|城中有一个贫穷的智慧人，他用智慧救了那城，却没有人记念那穷人。
ECCL|9|16|我就说，智慧胜过勇力；然而那贫穷人的智慧被人藐视，他的话也无人听从。
ECCL|9|17|宁可听智慧人安静的话语，不听掌权者在愚昧人中的喊声。
ECCL|9|18|智慧胜过打仗的兵器；但一个罪人能败坏许多善事。
ECCL|10|1|死苍蝇使做香的膏油散发臭气； 同样，一点愚昧也能压倒智慧和尊荣。
ECCL|10|2|智慧人的心居右； 愚昧人的心居左。
ECCL|10|3|愚昧人的行径显出无知， 对众人说，他是愚昧人。
ECCL|10|4|掌权者的怒气若向你发作， 不要离开你的本位， 因为镇定能平息大过。
ECCL|10|5|我见日光之下有一件祸患， 似乎出于统治者的错误，
ECCL|10|6|就是愚昧人立在高位； 有钱人却坐在低位。
ECCL|10|7|我见仆人骑马， 王子像仆人在地上步行。
ECCL|10|8|挖陷坑的，自己必陷在其中； 拆城墙的，自己必被蛇咬。
ECCL|10|9|开凿石头的，会受损伤； 劈开木头的，必遭危险。
ECCL|10|10|铁器钝了，若不将刃磨快，就必多费力气； 但智慧的益处在于使人成功。
ECCL|10|11|尚未行法术，蛇若咬人， 行法术的人就得不到什么好处了。
ECCL|10|12|智慧人的口说出恩言； 愚昧人的嘴吞灭自己，
ECCL|10|13|他口中的话语起头是愚昧， 终局是邪恶的狂妄。
ECCL|10|14|愚昧人多有话语。 人不知将来会发生什么事， 他身后的事谁能告诉他呢？
ECCL|10|15|愚昧人的劳碌使自己困乏， 连进城的路他也不知道。
ECCL|10|16|邦国啊，你的君王若年少， 你的群臣早晨宴乐， 你就有祸了！
ECCL|10|17|邦国啊，你的君王若是贵族之子， 你的群臣按时吃喝， 是为强身，不为酒醉， 你就有福了！
ECCL|10|18|因人懒惰，房顶塌下； 因人手懒，房屋滴漏。
ECCL|10|19|摆设宴席是为欢乐。 酒能使人快活， 钱能叫万事应心。
ECCL|10|20|不可诅咒君王， 连起意也不可， 在卧室里也不可诅咒富人； 因为空中的飞鸟必传扬这声音， 有翅膀的必述说这事。
ECCL|11|1|当将你的粮食撒在水面上， 因为日子久了，你必能得着它。
ECCL|11|2|将你所拥有的分给七人，或八人， 因为你不知道会有什么灾祸临到地上。
ECCL|11|3|云若满了雨，就必倾倒在地上。 树向南倒，或向北倒， 树倒在何处，就留在何处。
ECCL|11|4|看风的，必不撒种； 望云的，必不收割。
ECCL|11|5|你不知道气息如何进入孕妇的骨头里 ；照样，造万物之上帝的作为，你也无从得知。
ECCL|11|6|早晨要撒种，晚上也不要歇手，因为你不知道哪一样发旺；前者或后者，或两者都一样好。
ECCL|11|7|光是甜美的，眼见日光是多么好啊！
ECCL|11|8|人活多少年，就当快乐多少年，然而也当想到黑暗的日子；因为这样的日子必多，所要来临的全是虚空。
ECCL|11|9|年轻人哪，你在年少时当快乐；在年轻时使你的心欢畅，做你心所愿做的，看你眼所爱看的；却要知道，为这一切，上帝必审问你。
ECCL|11|10|所以，当从心中除掉愁烦，从肉体除去痛苦；因为年少和年轻之时，全是虚空。
ECCL|12|1|你趁着年轻、衰老的日子尚未来到，就是你所说，我毫无喜悦的那些岁月来临之前，当记念造你的主。
ECCL|12|2|不要等到太阳、光明、月亮、星宿变为黑暗，雨后云又返回；
ECCL|12|3|看守房屋的发颤，强壮的屈身，推磨的妇女因人少而停工，从窗户往外看的眼光变为昏暗；
ECCL|12|4|街门关闭，推磨的声音微小，鸟一叫，就惊醒，唱歌女子的声音也都微弱；
ECCL|12|5|人怕高处，路上有惊慌；杏树开花，蚱蜢成为重担，欲望不再挑起；因为人归他永远的家，吊丧的在街上往来。
ECCL|12|6|不要等到银链折断 ，金罐破裂，瓶子在泉旁损坏，水轮在井口断裂，
ECCL|12|7|尘土仍归于地，像原来一样，气息仍归于赐气息的上帝。
ECCL|12|8|传道者说：“虚空的虚空，全是虚空。”
ECCL|12|9|再者，传道者因有智慧，将知识教导众人；他思量，考察，并列举出许多箴言。
ECCL|12|10|传道者专心寻求可喜悦的言语，是凭正直写的诚实话。
ECCL|12|11|智慧人的话语如同刺棒；这些嘉言好像钉稳的钉子，都是一个牧者所赐的。
ECCL|12|12|我儿，还有一点，你当受劝戒：著书多，没有穷尽；读书多，身体疲倦。
ECCL|12|13|这些事都已听见了，结论就是：敬畏上帝，谨守他的诫命，这是人当尽的本分。
ECCL|12|14|因为人所做的事，连一切隐藏的事，无论是善是恶，上帝都必审问。
