DEUT|1|1|Оце ті слова, що Мойсей говорив був до всього Ізраїля по тім боці Йордану в пустині, на степу, навпроти Червоного моря, між Параном, і між Тофелем, і Лаваном, і Гецеротом, і Ді-Загавом,
DEUT|1|2|одинадцять день дороги від Хориву, дорога до гори Сеїру, аж до Кадеш-Барнеа.
DEUT|1|3|І сталося сорокового року, одинадцятого місяця, першого дня місяця говорив Мойсей до Ізраїлевих синів усе, що Господь наказав був йому про них,
DEUT|1|4|по тому, як забив він Сигона, царя аморейського, що сидів у Хешбоні, і Оґа, царя башанського, що сидів в Аштароті в Едреї.
DEUT|1|5|На тім боці Йордану в моавському краї став Мойсей виясняти Закона, говорячи:
DEUT|1|6|Господь, Бог наш, промовляв до нас на Хориві, говорячи: Досить вам сидіти на цій горі!
DEUT|1|7|Оберніться й рушайте, і йдіть на гору амореянина, та до всіх сусідів його на степу, на горі, і в долині, і на півдні, і на побережжі моря, до Краю ханаанського та до Ливану, аж до Великої Річки, річки Ефрату.
DEUT|1|8|Ось Я дав вам цей Край! Увійдіть, і заволодійте цим Краєм, що за нього Господь був присяг вашим батькам, Авраамові, Ісакові та Якову, що дасть його їм та їхньому насінню по них.
DEUT|1|9|І сказав я того часу до вас, говорячи: Не можу я сам носити вас.
DEUT|1|10|Господь, Бог ваш, розмножив вас, і ось ви сьогодні, щодо численности, як зорі небесні!
DEUT|1|11|Господь, Бог ваших батьків, нехай додасть вам у тисячу раз, і нехай поблагословить вас, як Він говорив вам.
DEUT|1|12|Як я сам понесу тяготу вашу, і тягар ваш, і ваші суперечки?
DEUT|1|13|Візьміть собі мужів мудрих, і випробуваних, і знаних вашим племенам, і я поставлю їх на чолі вас.
DEUT|1|14|І ви відповіли мені та й сказали: Добра та річ, що ти кажеш зробити.
DEUT|1|15|І взяв я голів ваших племен, мужів мудрих та знаних, і поставив їх головами над вами, тисячниками, і сотниками, і п'ятдесятниками, і десятниками, та урядниками для ваших племен.
DEUT|1|16|І наказав я того часу вашим суддям, говорячи: Вислуховуйте суперечки між вашими братами, і розсуджуйте справедливо між чоловіком та між братом його, та між приходьком його.
DEUT|1|17|Не будете звертати уваги на обличчя в суді, як малого, так і великого вислухаєте, не будете боятися обличчя людини, бо суд Божий він! А ту справу, що буде занадто тяжка для вас, принесете мені, і я вислухаю її.
DEUT|1|18|І наказав я вам того часу про всі ті речі, що ви зробите.
DEUT|1|19|І ми рушили з Хориву, та й перейшли цю велику й страшну пустиню, що бачили ви, дорогою до гори амореянина, як наказав нам Господь, Бог наш, і ми прийшли аж до Кадеш-Барнеа.
DEUT|1|20|І сказав я до вас: Прийшли ви до Аморейської гори, що Господь, Бог наш, дає нам.
DEUT|1|21|Ось, Господь, Бог твій, віддає тобі цей Край. Увійди, заволодій, як говорив був тобі Господь, Бог батьків твоїх. Не бійся й не лякайся!
DEUT|1|22|А ви всі підійшли до мене та й сказали: Пошлімо мужів перед собою, і нехай вони вислідять нам той Край, та нехай принесуть нам відомість про дорогу, що нею підемо, та про міста, куди ввійдемо.
DEUT|1|23|І була та річ добра в моїх очах, і взяв я у вас дванадцять мужа, муж один для племени.
DEUT|1|24|І вони відійшли, і зійшли на гору, і прийшли аж до долини Ешкол, та й вислідили його, Край.
DEUT|1|25|І взяли вони в свою руку з плоду того Краю, і принесли до нас, і здали нам справу, і сказали: Добрий той Край, що Господь, Бог наш, дає нам!
DEUT|1|26|Та ви не хотіли йти, і були неслухняні наказам Господа, Бога вашого.
DEUT|1|27|І нарікали ви по ваших наметах і говорили: З ненависти до нас Господь вивів нас з єгипетського краю, щоб дати нас у руку амореянина на вигублення нас.
DEUT|1|28|Куди ми підемо? Брати наші розслабили наше серце, говорячи: Народ той більший та вищий від нас, міста великі й уміцнені аж до неба, і навіть велетнів ми бачили там.
DEUT|1|29|І сказав я до вас: Не лякайтеся й не бійтеся їх!
DEUT|1|30|Господь, Бог наш, що йде перед вами, Він буде воювати для вас, як зробив був з вами в Єгипті на ваших очах,
DEUT|1|31|і в пустині, де ти бачив, що Господь, Бог твій, носив тебе, як носить чоловік сина свого, у всій дорозі, якою ви йшли, аж до вашого приходу до цього місця.
DEUT|1|32|Та все таки ви не віруєте в Господа, вашого Бога,
DEUT|1|33|що йде перед вами в дорозі, щоб вишукати для вас місце на ваше таборування, вночі огнем, щоб ви бачили в дорозі, що будете нею ходити, а хмарою вдень.
DEUT|1|34|І Господь вислухав голос ваших слів, та й розгнівався, і заприсягнув, говорячи:
DEUT|1|35|Поправді кажу, ніхто серед цих людей, цього злого покоління, не побачить того доброго Краю, що присяг Я дати вашим батькам,
DEUT|1|36|окрім Калева, Єфуннеєвого сина, він побачить його, і йому Я дам той Край, по якому ступав він, та синам його, через те, що він виповняв наказа Господнього.
DEUT|1|37|Також на мене розгнівався був Господь через вас, говорячи: І ти не ввійдеш туди!
DEUT|1|38|Ісус, син Навинів, що стоїть перед тобою, він увійде туди; зміцни його, бо він зробить, що Ізраїль заволодіє ним.
DEUT|1|39|А діти ваші, про яких ви сказали: На здобич будуть вони, та сини ваші, що сьогодні не знають ні добра, ані зла, вони ввійдуть туди, і їм дам Я його, і вони заволодіють ним.
DEUT|1|40|А ви йдіть, та й рушайте в пустиню дорогою Червоного моря.
DEUT|1|41|А ви відповіли та й сказали мені: Згрішили ми Господеві! Ми вийдемо, і будемо воювати, цілком так, як наказав нам Господь, Бог наш. І приперезали ви кожен військову зброю свою, і відважилися вийти на гору.
DEUT|1|42|Але Господь до мене сказав: Скажи їм: Не вийдете, і не будете ви воювати, бо Я не серед вас, щоб не були ви побиті вашими ворогами.
DEUT|1|43|І промовляв я до вас, та ви не послухали, і були неслухняні наказам Господнім. І ви свавільно переступили наказа, і зійшли на гору.
DEUT|1|44|І вийшов навперейми вас амореянин, що сидить на тій горі, і гнали вас, як роблять то бджоли, і товкли вас в Сеїрі аж до Горми.
DEUT|1|45|І вернулися ви, і плакали перед Господнім лицем, та не слухав Господь вашого голосу, і не нахилив Свого вуха до вас.
DEUT|1|46|І сиділи ви в Кадешу багато днів, стільки днів, скільки там ви сиділи.
DEUT|2|1|І обернулися ми та й рушили в пустиню дорогою до Червоного моря, як Господь промовляв був до мене. І кружляли ми навколо гори Сеїр багато днів.
DEUT|2|2|І сказав Господь до мене, говорячи:
DEUT|2|3|Досить вам кружляти навколо цієї гори, оберніться на північ!
DEUT|2|4|А народові наказуй, говорячи: Ви переходите границі ваших братів, Ісавових синів, що мешкають у Сеїрі. І будуть вони боятися вас, та й ви пильно стережіться!
DEUT|2|5|Не дражніть їх, бо Я не дам вам з їхнього краю місця ані на стопу ноги, бо гору Сеїр Я дав Ісавові, як спадщину.
DEUT|2|6|Їжу купите від них за срібло і будете їсти, а також воду будете купувати в них за срібло і будете пити.
DEUT|2|7|Бо Господь, Бог твій, поблагословив тебе в кожному чині твоєї руки, знає Він ходу твою в цій великій пустині. Оце сорок літ Господь, Бог твій, з тобою, не відчув ти недостачі ні в чому.
DEUT|2|8|І перейшли ми від наших братів, Ісавових синів, що сидять у Сеїрі, від дороги степу, від Елату, і від Ецйон-Ґеверу. І обернулися ми, та й перейшли дорогою моавської пустині.
DEUT|2|9|І сказав Господь мені: Не ворогуй з Моавом, і не дратуй їх війною, бо Я не дам тобі з його краю спадщини, бо Лотовим синам дав Я Ар на спадок.
DEUT|2|10|Перед тим сиділи в ньому еми, народ великий, і численний, і високий, як велетні.
DEUT|2|11|Рефаями вважалися й вони, як велетні, а моавітяни кличуть їх: еми.
DEUT|2|12|А в Сеїрі перед тим сиділи були гореї, а Ісавові сини заволоділи ними та вигубили їх перед собою, та й осіли замість них, як зробив Ізраїль Краєві спадку свого, що дав їм Господь.
DEUT|2|13|Тепер устаньте, і перейдіть поток Зеред. І перейшли ми потік Зеред.
DEUT|2|14|А час, що ходили ми від Кадеш-Барнеа, аж перейшли потік Зеред, тридцять і вісім літ, аж вимерло все те покоління військових із табору, як Господь присягнув був їм.
DEUT|2|15|Також і Господня рука була на них, щоб вигубити їх із табору аж до решти.
DEUT|2|16|І сталося, коли вигинули всі військові і вимерли з-посеред народу,
DEUT|2|17|то Господь промовляв до мене, говорячи:
DEUT|2|18|Ти сьогодні проходиш моавську границю Ар.
DEUT|2|19|І прийдеш близько до Аммонових синів, не ненавидь їх і не дратуй їх, бо не дам тобі спадку з краю Аммонових синів, бо Лотовим синам Я дав його на спадщину.
DEUT|2|20|За край рефаїв вважався також він, рефаї сиділи в ньому перед тим, а аммонітяни кликали їх: замзуми,
DEUT|2|21|народ великий, і численний, і високий, як велетні. І вигубив їх Господь перед ними, і вигнали їх, і осіли замість них,
DEUT|2|22|як зробив Він Ісавовим синам, що сидять у Сеїрі, що заволоділи хореянами перед ними, і вигнали їх, і осіли замість них, і сидять аж до сьогодні.
DEUT|2|23|А аввеїв, що сидять по оселях аж до Ази, вигубили їх кафтори, що вийшли з Кафтору, та й осіли замість них.
DEUT|2|24|Уставайте, рушайте, та й перейдіть потік Арнон! Ось Я дав у твою руку Сигона, царя Хешбону, амореянина, а край його зачни забирати, та й воюй з ним.
DEUT|2|25|Того дня Я зачну наводити страх та жах перед тобою на народи під усім небом, які, коли почують чутку про тебе, то затремтять, і жахнуться перед тобою.
DEUT|2|26|І послав я послів з пустині Кедемот до Сигона, царя хешбонського, з мирними словами, говорячи:
DEUT|2|27|Нехай же я перейду в твоїм краї в дорозі, я піду дорогою, не збочу ні праворуч, ні ліворуч.
DEUT|2|28|Їжу за срібло продаси мені, і я їстиму, і воду даси мені за срібло, і я питиму. Нехай тільки перейду я ногами,
DEUT|2|29|як зробили мені Ісавові сини, що сидять у Сеїрі, і моави, що сидять ув Арі, аж перейду я Йордан до того Краю, що його нам дає Господь, Бог наш.
DEUT|2|30|Та не хотів Сигон, цар хешбонський, дати нам перейти через свою землю, бо Господь, Бог твій, зробив запеклим дух його, та ожорсточив його серце, щоб дати його в руку твою, як сьогодні це видко.
DEUT|2|31|І сказав Господь мені: Ось, Я зачав давати перед тобою Сигона та його край; зачни заволодівати, щоб успадкувати його край.
DEUT|2|32|І вийшов Сигон навпроти нас, він та ввесь народ його, на війну до Ягацу.
DEUT|2|33|І дав його нам Господь, Бог наш, і ми побили його й синів його та ввесь його народ.
DEUT|2|34|І того часу ми здобули всі його міста, і зробили закляттям кожне місто, чоловіків і жінок та дітей, нікого не позоставили ми.
DEUT|2|35|Тільки худобу забрали ми собі на здобич, та захоплене в містах, що ми їх здобули.
DEUT|2|36|Від Ароеру, що на березі арнонського потоку, і від міста, що в долині, і аж до Ґілеаду не було міста, яке було б сильніше від нас, усе віддав нам Господь, Бог наш.
DEUT|2|37|Тільки до краю Аммонових синів не наблизився ти, до всього побережжя потоку Яббоку, і до міст гори, та до всього, про що наказав був Господь, Бог наш.
DEUT|3|1|І обернулися ми, та й пішли дорогою до Башану. І вийшов навперейми нас Оґ, цар башанський, він та ввесь його народ, на війну до Едреї.
DEUT|3|2|І сказав Господь до мене: Не бійся його, бо в твою руку Я дав його, і ввесь народ його та край його, і зробиш йому, як зробив ти Сигонові, цареві амореян, що сидів у Хешбоні.
DEUT|3|3|І дав Господь, Бог наш, у нашу руку також Оґа, царя башанського, та ввесь його народ, і побили ми його, так що нікого не позосталося в нього.
DEUT|3|4|І здобули ми всі міста його, і того часу не було міста, що не взяли б ми від них, шістдесят міст, усю арґовську околицю, царство Оґа в Башані.
DEUT|3|5|Усі ці міста укріплені, мур високий, ворота й засув, окрім дуже багатьох відкритих міст.
DEUT|3|6|І вчинили ми їх закляттям, як зробили були Сигонові, цареві хешбонському, учинили закляттям усе місто, чоловіків, жінок та дітей.
DEUT|3|7|А всю худобу й захоплене з міст забрали ми собі на здобич.
DEUT|3|8|І взяли ми того часу той край з руки обох царів амореянина, що по другому боці Йордану, від Арнонського потоку аж до гори Гермон,
DEUT|3|9|сидоняни кличуть на Гермон Сірйон, а амореяни кличуть на нього Сенір,
DEUT|3|10|усі міста на рівнині, і ввесь Ґілеад, і ввесь Башан аж до Салхи й Едреї, міст царства Оґа в Башані.
DEUT|3|11|Бо тільки Оґ, цар башанський, позостав із решти рефаїв. Оце його ложе, ложе залізне; чи ж не воно в Раббі Аммонових синів, дев'ять ліктів довжина його, і чотири лікті ширина його, на міру ліктем чоловіка.
DEUT|3|12|А Край той того часу посіли ми. Від Ароеру, що над Арнонським потоком, і половину гори Ґілеад, і міста його я дав Рувимовим та Ґадовим.
DEUT|3|13|А решту Ґілеаду та ввесь Башан, царство Оґа, віддав я половині племени Манасіїного, усю околицю арґовську, на ввесь той Башан кличеться: Край рефаїв.
DEUT|3|14|Яір, син Манасіїн, узяв всю Арґову околицю аж до границі ґешурів та маахатів, і він назвав їх своїм іменем: Башан, села Яіра, і так їх кличуть аж до цього дня.
DEUT|3|15|А Махірові дав я Ґілеад.
DEUT|3|16|А Рувимовим та Ґадовим дав я від Ґілеаду й аж до Арнонського потоку, середину потоку та границю, і аж до потоку Яббоку, границі Аммонових синів,
DEUT|3|17|і степ, і Йордан, і границю його від Кіннерету аж до моря степу, моря Солоного, у узбіччя Пісґі на схід.
DEUT|3|18|І часу того наказав я вам, говорячи: Господь, Бог ваш, дав вам цей Край, щоб ви посіли його; узброєні перейдете перед вашими братами, Ізраїлевими синами, усі військові.
DEUT|3|19|Тільки ваші жінки, і ваші діти та ваша худоба, я знаю, що худоба ваша велика! будуть сидіти по ваших містах, що я дав вам,
DEUT|3|20|аж Господь дасть спочинок братам вашим, як вам, і посядуть також вони той Край, що Господь, Бог ваш, дає вам по той бік Йордану, і вернетесь кожен до спадку свого, що я дав вам.
DEUT|3|21|А Ісусові наказав я того часу, говорячи: Ото твої очі бачили все, що зробив був Господь, Бог ваш, обом тим царям, так зробить Господь усім царствам, куди ти переходиш.
DEUT|3|22|Не будеш боятися їх, бо Господь, Бог ваш, Він Той, що воює для вас.
DEUT|3|23|І благав я того часу Господа, говорячи:
DEUT|3|24|Владико Господи, Ти зачав показувати рабові Своєму велич Свою та міцну Свою руку! Бо хто інший Бог на небі та на землі, що зробить, як чини Твої, як великі діла Твої?
DEUT|3|25|Нехай перейду ж я та побачу той хороший Край, що по тім боці Йордану, ту гарну гірську землю та Ливан!
DEUT|3|26|Та Господь розгнівався на мене через вас, і не послухав мене. І сказав Господь до мене: Досить тобі, не говори більше до Мене в цій справі!
DEUT|3|27|Вийди на верхів'я Пісґі, і зведи свої очі на захід, і на північ, і на південь, і на схід, і побач своїми очима, бо ти не перейдеш цього Йордану!
DEUT|3|28|І напоуми Ісуса, і зміцни його, й укріпи його, бо він перейде перед цим народом, і він зробить, що вони посядуть той Край, який ти побачиш.
DEUT|3|29|І осіли ми в долині навпроти Бет-Пеору.
DEUT|4|1|А тепер, Ізраїлю, послухай постанов та законів, що я навчаю вас чинити, щоб жили ви, і ввійшли, й посіли цей Край, що Господь, Бог батьків ваших, дає вам.
DEUT|4|2|Не додавайте до того, що я вам наказую, і не зменшайте з того, щоб виконувати заповіді Господа, Бога вашого, що я наказав вам.
DEUT|4|3|Очі ваші бачили те, що Господь зробив був з Ваалом пеорським, бо кожного чоловіка, що пішов за пеорським Ваалом, вигубив його Господь, Бог твій, з-посеред тебе.
DEUT|4|4|А ви, що линули до Господа, Бога вашого, усі ви живі сьогодні.
DEUT|4|5|Дивіться, навчив я вас постанов та законів, як наказав мені Господь, Бог мій, чинити так серед того Краю, куди ви входите, щоб посісти його.
DEUT|4|6|Бережіть, і виконуйте їх, бо це мудрість ваша та ваш розум на очах народів, що вислухають усіх постанов тих та й скажуть: Тільки він мудрий та розумний народ, цей великий люд!
DEUT|4|7|Бо хто інший такий великий народ, що мав би богів, таких йому близьких, як Господь, Бог наш, кожного разу, як ми кличемо до Нього?
DEUT|4|8|І хто інший такий великий народ, що має постанови й закони такі справедливі, як увесь той Закон, що я даю перед вами сьогодні?
DEUT|4|9|Тільки стережися, і дуже пильнуй свою душу, щоб не забув ти тих речей, що бачили очі твої, і щоб вони не повиходили з серця твого по всі дні життя твого, а ти подаси їх до відома синам твоїм та синам твоїх синів,
DEUT|4|10|про день, коли стояв ти перед лицем Господа, Бога твого, на Хориві, як Господь говорив був до мене: Збери Мені той народ, і вони слухатимуть слів Моїх, із яких навчаться боятися Мене по всі дні, скільки вони житимуть на землі, та й синів своїх понавчають.
DEUT|4|11|І поприходили ви, та й поставали під горою, а гора та горіла огнем аж до самих небес, а при тому була темрява, хмара та мряка.
DEUT|4|12|І промовляв Господь до вас із середини огню, голос слів ви чули, та виду ви не бачили, окрім голосу.
DEUT|4|13|І Він оголосив перед вами заповіта Свого, що наказав вам чинити, Десять Заповідей, і написав їх на двох камінних таблицях.
DEUT|4|14|А мені Господь наказав того часу навчати вас постанов та законів, щоб виконували ви їх у Краю, куди ви переходите володіти ним.
DEUT|4|15|І будете ви сильно стерегти свої душі, бо не бачили ви того дня жодної постаті, коли говорив Господь до вас на Хориві з середини огню,
DEUT|4|16|щоб ви не зіпсулися, і не зробили собі ідола на подобу якогось боввана, зображення самця чи самиці,
DEUT|4|17|зображення всякої худобини, що на землі, зображення всякого крилатого птаха, що літає під небом,
DEUT|4|18|зображення всякого плазуючого по землі, зображення всякої риби, що в воді під землею,
DEUT|4|19|і щоб ти, звівши очі свої до неба, і побачивши сонце, і місяць, і зорі, усе військо небесне, щоб не був ти зведений і не вклонявся їм, і не служив їм; бо Господь, Бог твій, приділив їх усім народам під усім небом.
DEUT|4|20|А вас Господь узяв та й вивів вас із залізної гутничої печі, з Єгипту, щоб ви стали для Нього народом наділу, як сьогодні це видко.
DEUT|4|21|А Господь був розгнівався на мене за ваші діла, і поклявся, що не перейду я Йордану, і не ввійду до того хорошого Краю, що Господь, Бог твій, дає тобі на спадщину.
DEUT|4|22|Бо я умру в цьому краї, я не перейду Йордану, а ви перейдете й посядете той хороший Край.
DEUT|4|23|Стережіться, щоб не забули ви заповіту Господа, вашого Бога, якого склав з вами, щоб не зробили ви собі боввана на подобу всього, як наказав тобі Господь, Бог твій.
DEUT|4|24|Бо Господь, Бог твій, Він палючий огонь, Бог заздрісний.
DEUT|4|25|Коли ти породиш синів, і синів твоїх синів, і постарієте ви в Краю, і зіпсуєтеся, і зробите боввана на подобу чогось, і зробите зло в очах Господа, Бога свого, та Його розгнівите,
DEUT|4|26|то беру Я сьогодні за свідків проти вас небо й землю, що незабаром конче погинете в Краю, на вспадкування якого ви переходите туди Йордан. Не будуть довгі ваші дні в ньому, бо конче ви будете вигублені.
DEUT|4|27|І розпорошить вас Господь посеред народів, і будете ви нечисленні поміж людами, куди попровадить вас Господь.
DEUT|4|28|І будете служити там богам, ділу рук людських, дереву та каменеві, які не бачать, і не чують, і не їдять, і не нюхають.
DEUT|4|29|Та коли ви будете шукати звідти Господа, Бога свого, то знайдете, якщо будете шукати Його всім серцем своїм та всією душею своєю.
DEUT|4|30|Як будеш у біді своїй, і коли спіткають тебе в кінці днів усі оці речі, то вернешся ти до Господа, Бога свого, і послухаєш Його голосу.
DEUT|4|31|Бо Господь, Бог твій Бог милостивий: Він не залишить тебе й не знищить тебе, і не забуде заповіту батьків твоїх, яким їм присягнув був.
DEUT|4|32|Бо питай но про перші дні, що були перше тебе, від того дня, коли Бог створив людину на землі, і від кінця неба й аж до кінця неба, чи бувало щось таке, як ця велика річ, або чи чуте було щось таке, як вона:
DEUT|4|33|чи чув народ голос Бога, що говорив із середини огню, як чув ти і жив?
DEUT|4|34|Або чи намагався який бог піти взяти собі народ з-посеред іншого народу пробами, ознаками, і чудами, і війною, і сильною рукою, і раменом витягненим, і страхами великими, як усе те, що зробив був вам Господь, Бог ваш, в Єгипті на очах твоїх?
DEUT|4|35|Тобі було показане це, щоб ти пізнав, що Господь Він Бог, і нема іншого, окрім Нього.
DEUT|4|36|Він дав тобі з неба почути Його голос, щоб навчити тебе, а на землі показав тобі Свій великий огонь, і слова Його чув ти з середини огню.
DEUT|4|37|І тому, що кохав Він батьків твоїх, то вибрав їхнє насіння по них, і Сам Він вивів тебе Своєю великою силою з Єгипту,
DEUT|4|38|щоб прогнати перед тобою народи, більші й сильніші за тебе, щоб ввести тебе, та дати тобі їхній Край на спадок, як сьогодні це видко.
DEUT|4|39|І пізнаєш сьогодні, і візьмеш до серця свого, що Господь Він Бог на небі вгорі й на землі долі, іншого нема.
DEUT|4|40|І будеш пильнувати постанов Його та заповідей Його, що я наказую тобі сьогодні, щоб було добре тобі та синам твоїм по тобі, і щоб ти продовжив дні на землі, що Господь, Бог твій, дає тобі на всі дні.
DEUT|4|41|Тоді виділив Мойсей три місті по той бік Йордану на схід сонця,
DEUT|4|42|щоб утікав туди убійник, що замордує свого ближнього ненароком, а він не був йому ворогом ні вчора, ані позавчора. І втече він до одного з цих міст, і буде жити:
DEUT|4|43|Бецер у пустині, у краї рівниннім, Рувимовому, і Рамот у Ґілеаді Ґадовому, і Ґолан у Башані Манасіїному.
DEUT|4|44|І оце Закон, що Мойсей поклав перед Ізраїлевими синами,
DEUT|4|45|оце свідоцтва, і постанови, і закони, що Мойсей говорив їх до Ізраїлевих синів при виході їх із Єгипту,
DEUT|4|46|по той бік Йордану в долині навпроти Бет-Пеору в краю Сигона, царя аморейського, що сидів у Хешбоні, якого побив Мойсей та Ізраїлеві сини при виході їх із Єгипту.
DEUT|4|47|І вони оволоділи краєм його та краєм Оґа, башанського царя, обох аморейських царів, що по той бік Йордану на схід сонця,
DEUT|4|48|від Ароеру, що над берегом арнонського потоку, і аж до гори Сіон, цебто Гермон,
DEUT|4|49|і ввесь степ по тім боці Йордану на схід і аж до моря степу під узбіччям Пісґі.
DEUT|5|1|І скликав Мойсей усього Ізраїля, та й сказав до нього: Слухай, Ізраїлю, постанови й закони, які я говорю сьогодні в ваші уші, і навчіться їх, і будете пильнувати виконувати їх.
DEUT|5|2|Господь, Бог наш, склав з нами заповіта на Хориві.
DEUT|5|3|Не з батьками нашими склав Господь заповіта того, але з нами самими, що ми тут сьогодні всі живі.
DEUT|5|4|Обличчям в обличчя говорив Господь із вами на горі з середини огню.
DEUT|5|5|Я того часу стояв між Господом та між вами, щоб передавати вам Господні слова, бо ви боялися огню, і ви не зійшли на гору, коли Він говорив:
DEUT|5|6|Я Господь, Бог твій, що вивів тебе з єгипетського краю, з дому рабства.
DEUT|5|7|Хай не буде тобі інших богів при Мені!
DEUT|5|8|Не роби собі різьби й усякої подоби з того, що на небі вгорі, і що на землі долі, і що в воді під землею.
DEUT|5|9|Не вклоняйся їм, і не служи їм, бо Я Господь, Бог твій, Бог заздрісний, що карає провину батьків на синах, на третіх і на четвертих поколіннях тих, що ненавидять Мене,
DEUT|5|10|і що чинить милість тисячам поколінь тих, хто любить Мене, і хто виконує Мої заповіді.
DEUT|5|11|Не присягай Іменем Господа, Бога твого, надаремно, бо не помилує Господь того, хто присягає Його Ім'ям надаремно.
DEUT|5|12|Пильнуй дня суботнього, щоб святити його, як наказав тобі Господь, Бог твій.
DEUT|5|13|Шість день працюй, і роби всю працю свою,
DEUT|5|14|а день сьомий субота для Господа, Бога твого; не роби жодної праці ти й син твій та дочка твоя, і раб твій та невільниця твоя, і віл твій, і осел твій, і всяка худоба твоя, і приходько твій, що в брамах твоїх, щоб відпочив раб твій і невільниця твоя, як і ти.
DEUT|5|15|І будеш пам'ятати, що був ти рабом в єгипетському краї, і вивів тебе Господь, Бог твій, звідти сильною рукою та витягненим раменом, тому наказав тобі Господь, Бог твій, святкувати суботній день.
DEUT|5|16|Шануй свого батька та матір свою, як наказав був тобі Господь, Бог твій, щоб довгі були твої дні, і щоб було тобі добре на землі, яку Господь, Бог твій, дає тобі.
DEUT|5|17|Не вбивай!
DEUT|5|18|Не чини перелюбу!
DEUT|5|19|Не кради!
DEUT|5|20|Не свідчи неправдиво проти ближнього свого!
DEUT|5|21|І не бажай жони ближнього свого, і не бажай дому ближнього свого, ані поля його, ані раба його, ані невільниці його, ані вола його, ані осла його, ані всього, що є ближнього твого!
DEUT|5|22|Слова ці Господь промовляв до всього вашого зібрання, на горі з середини огню, хмари та мряки, сильним голосом. І більш не говорив, і написав їх на двох камінних таблицях, і дав їх мені.
DEUT|5|23|І сталося, коли ви слухали той голос з-посеред темряви, а гора горіла огнем, то прийшли до мене всі голови ваших племен та ваші старші,
DEUT|5|24|та й сказали: Тож Господь, Бог наш, показав нам славу Свою та велич Свою, і голос Його чули ми з середини огню. Цього дня ми бачили, що говорить Бог з людиною, і вона жива!
DEUT|5|25|А тепер нащо маємо вмирати? Бо спалить нас той великий огонь! Якщо ми будемо ще далі слухати голосу Господа Бога нашого, то помремо.
DEUT|5|26|Бо чи є таке тіло, щоб чуло, як ми, голос Бога Живого, що промовляє з середини огню, і жило б?
DEUT|5|27|Приступи сам, і слухай усе, що скаже Господь, Бог наш, і ти будеш говорити нам усе, що промовлятиме Господь, Бог наш, до тебе, а ми будемо слухати й виконаємо.
DEUT|5|28|І почув Господь голос ваших слів, коли ви промовляли до мене. І сказав до мене Господь: Чув Я голос цього народу, що промовляли до тебе. Добре все, що вони промовляли.
DEUT|5|29|О, коли б їхнє серце було їм на те, щоб боялись Мене й пильнували всіх Моїх заповідей по всі дні, щоб було добре їм та синам їхнім навіки!
DEUT|5|30|Іди, скажи їм: Вертайтесь собі до наметів своїх!
DEUT|5|31|А ти стій тут зо Мною, і Я буду промовляти до тебе кожну заповідь, і постанови, і закони, що будеш навчати їх, щоб вони виконували їх у Краї, що Я даю їм на спадщину його.
DEUT|5|32|І будеш пильнувати виконувати їх, як наказав вам Господь, Бог ваш, не збочите ні праворуч, ні ліворуч.
DEUT|5|33|Усією тією дорогою, що наказав вам Господь, Бог ваш, будете ходити, щоб жили ви й було вам добре, і щоб довгі були ваші дні в Краї, що ви оволодієте ним.
DEUT|6|1|А оце заповідь, постанови та закони, що наказав Господь, Бог ваш, щоб навчити вас виконувати їх у Краї, що ви переходите туди посісти його,
DEUT|6|2|щоб ти боявся Господа, Бога свого, щоб пильнувати всіх постанов Його та заповідей Його, що я наказую тобі, ти й син твій, та син твого сина по всі дні життя твого, і щоб були довгі твої дні.
DEUT|6|3|І слухай, Ізраїлю, і пильнуй виконувати це, щоб було добре тобі, і щоб ви сильно розмножились, як прирік був Господь, Бог батьків твоїх, дати Край, що тече молоком та медом.
DEUT|6|4|Слухай, Ізраїлю: Господь, Бог наш Господь один!
DEUT|6|5|І люби Господа, Бога твого, усім серцем своїм, і всією душею своєю, і всією силою своєю!
DEUT|6|6|І будуть ці слова, що Я сьогодні наказую, на серці твоїм.
DEUT|6|7|І пильно навчиш цього синів своїх, і будеш говорити про них, як сидітимеш удома, і як ходитимеш дорогою, і коли ти лежатимеш, і коли ти вставатимеш.
DEUT|6|8|І прив'яжеш їх на ознаку на руку свою, і будуть вони пов'язкою між очима твоїми.
DEUT|6|9|І напишеш їх на бічних одвірках дому свого та на брамах своїх.
DEUT|6|10|І станеться, коли Господь, Бог твій, уведе тебе до того Краю, якого присягнув був батькам твоїм, Авраамові, Ісакові та Якову, щоб дати тобі великі та гарні міста, яких ти не будував,
DEUT|6|11|та доми, повні всякого добра, яких ти не наповнював, і тесані колодязі, яких ти не тесав, і виноградники та оливки, яких ти не садив, і ти будеш їсти й наситишся,
DEUT|6|12|стережися тоді, щоб ти не забув Господа, що вивів тебе з єгипетського краю, з дому рабства!
DEUT|6|13|Бійся Господа, Бога свого, і Йому будеш служити, і Йменням Його будеш присягати.
DEUT|6|14|Не будеш ходити за іншими богами з богів тих народів, що в околицях ваших,
DEUT|6|15|бо Господь, Бог твій Бог заздрісний посеред тебе; щоб не запалився на тебе гнів Господа, Бога твого, і щоб Він не вигубив тебе з поверхні землі.
DEUT|6|16|Не будете спокушати Господа, Бога вашого, як спокушали ви в Массі.
DEUT|6|17|Будете конче пильнувати заповідей Господа, Бога вашого, і свідоцтва Його, і постанови Його, що наказав Він тобі.
DEUT|6|18|І будеш робити справедливе та добре в Господніх очах, щоб було тобі добре, і щоб увійшов ти та посів той хороший Край, що Господь присягнув був батькам твоїм,
DEUT|6|19|щоб вигнати всіх ворогів твоїх перед тобою, як говорив був Господь.
DEUT|6|20|Коли запитає тебе син твій колись, говорячи: Що це за свідоцтва й постанови та закони, що вам наказав Господь, Бог наш?
DEUT|6|21|то скажеш синові своєму: Ми були раби фараонові в Єгипті, а Господь вивів нас із Єгипту сильною рукою.
DEUT|6|22|І дав Господь ознаки та чуда великі та страшні на Єгипет, і на фараона та ввесь дім його на наших очах.
DEUT|6|23|А нас вивів звідти, щоб увести нас та дати той Край, що присягнув був Він нашим батькам.
DEUT|6|24|І наказав нам Господь чинити всі ті постанови, щоб боятися Господа, Бога нашого, щоб було добре нам усі дні, щоб утримати нас при житті, як дня цього.
DEUT|6|25|І буде нам праведність у тому, коли будемо пильнувати виконувати всі ці заповіді перед лицем Господа, Бога нашого, як Він наказав нам.
DEUT|7|1|Коли Господь, Бог твій, уведе тебе до того Краю, куди ти входиш, щоб заволодіти ним, то Він вижене численні поганські народи перед тобою: хіттеянина, і ґірґашеянина, і амореянина, і ханаанеянина, і періззеянина, і хіввеянина, і євусеянина, сім народів, численніших та міцніших за тебе.
DEUT|7|2|І коли дасть їх Господь, Бог твій, тобі, то ти їх понищиш: конче учиниш їх закляттям, не складеш із ними заповіту, і не будеш до них милосердний.
DEUT|7|3|І не споріднюйся з ними: дочки своєї не даси його синові, а його дочки не візьмеш для сина свого,
DEUT|7|4|бо він відверне сина твого від Мене, і вони служитимуть іншим богам, і запалиться Господній гнів на вас, і Він скоро тебе вигубить.
DEUT|7|5|Але тільки так будете їм робити: жертівники їхні порозбиваєте, а їхні стовпи поламаєте, святі їхні дерева постинаєте, а бовванів їхніх попалите в огні,
DEUT|7|6|бо ти святий народ для Господа, Бога свого, тебе вибрав Господь, Бог твій, щоб ти був Йому вибраним народом зо всіх народів, що на поверхні землі.
DEUT|7|7|Не через численність вашу понад усі народи Господь уподобав вас та вибрав вас, бож ви найменші зо всіх народів,
DEUT|7|8|але з Господньої любови до вас, і через додержання Його присяги, що присягнув був вашим батькам, Господь вивів вас сильною рукою, і викупив тебе з дому рабства, з руки фараона, царя єгипетського.
DEUT|7|9|І ти пізнаєш, що Господь, Бог твій, Він той Бог, той Бог вірний, що стереже заповіта та милість для тих, хто любить Його, та хто додержує Його заповіді на тисячу поколінь,
DEUT|7|10|і що надолужить ненависникам Своїм, їм самим, щоб вигубити їх; не загаїться Він щодо Свого ненависника, відплатить йому самому.
DEUT|7|11|А ти будеш виконувати заповіді й постанови та закони, що Я сьогодні наказую виконувати їх.
DEUT|7|12|І станеться, за те, що ви будете слухатися цих законів, і будете додержувати, і будете виконувати їх, то й Господь, Бог твій, буде додержувати для тебе заповіт та милість, що був присягнув батькам твоїм.
DEUT|7|13|І буде Він любити тебе, і поблагословить тебе, і розмножить тебе, і поблагословить плід твоєї, утроби та плід твоєї землі, збіжжя твоє, і сік твій виноградний, і сік твоїх оливок, порід биків твоїх і котіння отари твоєї на тій землі, яку присягнув батькам твоїм дати тобі.
DEUT|7|14|Ти будеш благословенний поміж усіма народами, не буде серед тебе безплідного та безплідної, також і між худобою твоєю.
DEUT|7|15|І Господь відхилить від тебе всяку хворобу, і жодних лютих єгипетських недуг, які ти знаєш, не наведе їх на тебе, а дасть їх на всіх твоїх ворогів.
DEUT|7|16|І ти винищиш всі ті народи, що Господь, Бог твій, дає тобі, не змилосердиться око твоє над ними, і не будеш служити їхнім богам, бо то пастка для тебе.
DEUT|7|17|Коли скажеш у серці своїм: Ті люди численніші від мене, як я зможу вигнати їх?
DEUT|7|18|не бійся їх! Пильно пам'ятай, що зробив був Господь, Бог твій, фараонові та всьому Єгиптові,
DEUT|7|19|ті великі випробовування, що бачили твої очі, і ознаки та чуда, і сильну руку та витягнене рамено, що ними вивів тебе Господь, Бог твій, так Господь, Бог твій, учинить усім тим народом, що ти їх боїшся.
DEUT|7|20|Також і шершнів пошле Господь, Бог твій, на нього, аж поки не вигинуть позосталі та ті, що поховалися перед тобою.
DEUT|7|21|Не бійся їх, бо серед тебе Господь, Бог твій, Бог великий та страшний.
DEUT|7|22|І викидатиме Господь, Бог твій, тих людей помалу з-перед тебе; не зможеш вигубити їх скоро, щоб не розмножилася над тобою польова звірина.
DEUT|7|23|І дасть їх Господь, Бог твій, перед тобою, і побентежить їх великим бентеженням, аж поки не будуть вигублені.
DEUT|7|24|І віддасть їхніх царів у руку твою, а ти вигубиш їхнє ім'я з-під неба, не встоїть ніхто перед тобою, аж поки ти не вигубиш їх.
DEUT|7|25|Бовванів їхніх богів попалите в огні, не будеш жадати срібла та золота, що на них, і не візьмеш його собі, щоб тим не впасти до пастки, бо то огида для Господа, Бога твого.
DEUT|7|26|І не внесеш цієї огиди до дому свого, і не станеш закляттям, як вона. Конче зогидиш її, і конче будеш бридитися нею, бо закляття вона.
DEUT|8|1|Усі заповіді, що я сьогодні наказав тобі, будете пильнувати виконувати, щоб ви жили, і множилися, і ввійшли й посіли той Край, що Господь присягнув вашим батькам.
DEUT|8|2|І будеш пам'ятати всю ту дорогу, що Господь, Бог твій, вів тебе нею по пустині ось уже сорок літ, щоб упокорити тебе, щоб випробувати тебе, щоб пізнати те, що в серці твоїм, чи будеш ти держати заповіді Його, чи ні.
DEUT|8|3|І впокорював Він тебе, і морив тебе голодом, і годував тебе манною, якої не знав ти й не знали батьки твої, щоб дати тобі знати, що не хлібом самим живе людина, але всім тим, що виходить із уст Господніх, живе людина.
DEUT|8|4|Одежа твоя не витиралася на тобі, а нога твоя не спухла от уже сорок літ.
DEUT|8|5|І пізнаєш ти в серці своїм, що, як навчає чоловік сина свого, так навчає тебе Господь, Бог твій.
DEUT|8|6|І будеш виконувати заповіді Господа, Бога свого, щоб ходити Його дорогами, та щоб боятися Його,
DEUT|8|7|бо Господь, Бог твій, уводить тебе до Краю хорошого, до Краю водних потоків, джерел та безодень, що виходять у долині й на горі,
DEUT|8|8|до Краю пшениці, й ячменю, і винограду, і фіґи, і гранату, до Краю оливкового дерева та меду,
DEUT|8|9|до Краю, де подостатком будеш їсти хліб, де не забракне нічого, до Краю, що каміння його залізо, а з його гір добуватимеш мідь.
DEUT|8|10|І будеш ти їсти й наситишся, і поблагословиш Господа, Бога свого, у тім добрім Краї, що дав Він тобі.
DEUT|8|11|Стережися, щоб не забув ти Господа, Бога свого, щоб не пильнувати Його заповідей, і законів Його, і постанов Його, що я сьогодні наказую тобі,
DEUT|8|12|щоб, коли ти будеш їсти й наситишся, і добрі доми будуватимеш, і осядеш у них,
DEUT|8|13|а худоба твоя велика та худоба твоя мала розмножиться, і срібло та золото розмножаться тобі, і все, що твоє, розмножиться,
DEUT|8|14|то щоб не загордилося серце твоє, і щоб не забув ти Господа, Бога свого, що вивів тебе з єгипетського краю, з дому рабства,
DEUT|8|15|що веде тебе цією великою пустинею, яка збуджує страх, де вуж, сараф, і скорпіон, і висохла земля, де немає води; що Він випроваджує тобі воду з крем'яної скелі,
DEUT|8|16|що в пустині годує тебе манною, якої не знали батьки твої, щоб упокоряти тебе, і щоб випробовувати тебе, щоб чинити тобі добро наостанку,
DEUT|8|17|щоб ти не сказав у серці своїм: Сила моя та міць моєї руки здобули мені цей добробут.
DEUT|8|18|І будеш ти пам'ятати Господа, Бога свого, бо Він Той, що дає тобі силу набути потугу, щоб виконати Свого заповіта, якого присягнув Він батькам твоїм, як дня цього.
DEUT|8|19|І станеться, якщо справді забудеш ти Господа, Бога свого, і підеш за іншими богами, і будеш їм служити, і будеш вклонятися їм, то врочисто свідчу вам сьогодні, ви конче погинете!
DEUT|8|20|Як ті люди, що Господь вигубляє з-перед вас, так ви погинете за те, що не будете слухатися голосу Господа, Бога вашого!
DEUT|9|1|Слухай, Ізраїлю: ти сьогодні переходиш Йордан, щоб увійти й заволодіти народами, більшими й міцнішими від тебе, містами великими й укріпленими аж до неба,
DEUT|9|2|народом великим та високим, велетнями, яких ти знаєш, і про яких ти чув: Хто стане перед велетнями?
DEUT|9|3|І познаєш сьогодні, що Господь, Бог твій, Він Той, що переходить перед тобою, як огонь поїдаючий, Він вигубить їх і Він понижуватиме їх перед тобою. І ти виженеш їх і вигубиш їх незабаром, як Господь говорив був тобі.
DEUT|9|4|Не скажи в серці своїм, коли Господь, Бог твій, буде їх виганяти з-перед тебе, говорячи: Через праведність мою ввів мене Господь посісти цей Край, і через неправедність цих людей Господь виганяє їх з-перед мене.
DEUT|9|5|Не через праведність твою, і не через простоту твого серця ти входиш володіти їхнім Краєм, але, через неправедність цих людей Господь, Бог твій, виганяє їх з-перед тебе, і щоб виконати те слово, що присягнув був Господь батькам твоїм, Авраамові, Ісакові та Якову.
DEUT|9|6|І пізнаєш, що не через праведність твою Господь, Бог твій, дає тобі посісти цей хороший Край, бо ти народ твердошиїй.
DEUT|9|7|Пам'ятай, не забудь, що ти гнівив Господа, Бога свого, у пустині від дня, коли вийшов ти з єгипетського краю аж до приходу вашого до цього місця, неслухняні були ви проти Господа.
DEUT|9|8|І на Хориві розгнівили були ви Господа, і Господь був розгнівався на вас, щоб вигубити вас.
DEUT|9|9|Коли я сходив на гору взяти кам'яні таблиці заповіту, що Господь склав був із вами, то сидів я на горі сорок день і сорок ночей, хліба не їв, і води не пив.
DEUT|9|10|І Господь дав мені обидві кам'яні таблиці, писані Божим перстом, а на них усі ті слова, що Господь говорив був із вами на горі з середини огню в дні зборів.
DEUT|9|11|І сталося, на кінці сорока день і сорока ночей дав мені Господь дві кам'яні таблиці, таблиці заповіту.
DEUT|9|12|І сказав мені Господь: Устань, швидко зійди звідси, бо зіпсувся народ твій, що ти вивів з Єгипту. Вони скоро збочили з дороги, яку Я наказав їм, зробили собі литого боввана.
DEUT|9|13|І сказав Господь до мене, говорячи: Бачив Я той народ, і ось він народ твердошиїй.
DEUT|9|14|Позостав Мене, і Я вигублю їх, і зітру їхнє ймення з-під неба, тебе зроблю народом міцнішим та численнішим від нього.
DEUT|9|15|І я обернувся, і зійшов із гори, а гора палає в огні, і обидві таблиці заповіту в обох руках моїх.
DEUT|9|16|І побачив я, а ось ви згрішили проти Господа, Бога вашого, зробили собі теля, литого боввана, зійшли скоро з дороги, яку Господь наказав був вам!
DEUT|9|17|І схопив я за обидві таблиці, та й кинув їх з обох своїх рук, і розторощив їх на ваших очах!...
DEUT|9|18|І впав я перед Господнім лицем, як перше, сорок день і сорок ночей хліба не їв і води не пив, за ввесь ваш гріх, що згрішили ви, як чинили зло в очах Господа, щоб Його розгнівити,
DEUT|9|19|бо боявся я гніву та люті, якими розгнівався був на вас Господь, щоб вигубити вас, та вислухав Господь мене й цього разу.
DEUT|9|20|А на Аарона Господь дуже розгнівався був, щоб погубити його. І молився я того часу також за Аарона.
DEUT|9|21|А гріх ваш, що вчинили ви, теля те я взяв та й спалив його в огні, і розторощив його, добре змолов, аж стало воно дрібним, немов порох. І кинув я порох його до потоку, що сходить з гори.
DEUT|9|22|І в Тав'ері, і в Массі, і в Ківрот-Гаттааві гнівили ви Господа.
DEUT|9|23|А коли Господь посилав вас з Кадеш-Барнеа, говорячи: Увійдіть, та й посядьте той Край, що Я дав вам, то були ви неслухняні наказу Господа, Бога вашого, і не повірили Йому, і не послухалися Його голосу.
DEUT|9|24|Неслухняні були ви Господеві від дня, як я вас пізнав.
DEUT|9|25|І впав я перед Господнім лицем на ті сорок день і сорок ночей, що я був упав, бо Господь сказав, що вигубить вас.
DEUT|9|26|І молився я до Господа й говорив: Владико Господи, не губи народу Свого та насліддя Свого, що Ти викупив Своєю величністю, що Ти вивів його з Єгипту сильною рукою!
DEUT|9|27|Згадай Своїх рабів Авраама, Ісака та Якова, не вважай на запеклість цього народу й на несправедливість та гріх його,
DEUT|9|28|щоб не сказав той край, звідки вивів ти нас: Не міг Господь увести їх до того Краю, що Ти говорив їм, та з Своєї ненависти до них Ти вивів їх, щоб побити їх у пустині.
DEUT|9|29|А вони народ Твій та насліддя Твоє, що Ти вивів Своєю великою силою та Своїм витягненим раменом.
DEUT|10|1|Того часу сказав був до мене Господь: Витеши собі дві камінні таблиці, як перші, та й вийде до Мене на гору, і зроби собі дерев'яного ковчега.
DEUT|10|2|А Я напишу на тих таблицях слова, що були на перших таблицях, які ти побив, і покладеш їх у ковчезі.
DEUT|10|3|І зробив я ковчега з акаційного дерева, і витесав я дві камінні таблиці, як перші, та й зійшов на гору, а обидві таблиці в руці моїй.
DEUT|10|4|І Він написав на тих таблицях, як перше письмо, Десять Заповідей, що Господь говорив був до вас на горі з середини огню в день зборів. І Господь дав їх мені.
DEUT|10|5|І обернувся я, та й зійшов із гори, і поклав ті таблиці, що зробив, до ковчегу. І були вони там, як наказав був Господь.
DEUT|10|6|А Ізраїлеві сини рушили з Беероту Яаканових синів до Мосери. Там помер Аарон, і був там похований, а священиком став замість нього його син Елеазар.
DEUT|10|7|А звідти рушили до Ґудґоди, а з Ґудґоди до Йотвати, до краю водних потоків.
DEUT|10|8|Того часу Господь відділив був Левієве плем'я, щоб носило ковчега Господнього заповіту, щоб стояло перед Господнім лицем, щоб служило Йому, і щоб благословляло Його Йменням аж до цього дня.
DEUT|10|9|Тому не було Левієві частки та спадку з братами. Господь Він спадщина його, як промовляв був Господь, Бог твій, йому.
DEUT|10|10|А я стояв на горі, як за тих перших днів, сорок день і сорок ночей. І вислухав Господь мене також цього разу, не захотів Господь погубити тебе.
DEUT|10|11|І сказав був до мене Господь: Устань, іди в похід перед народом. І ввійдуть вони, і посядуть той Край, що Я присягнув був їхнім батькам дати їм.
DEUT|10|12|А тепер, Ізраїлю, чого жадає від тебе Господь, Бог твій? Тільки того, щоб боятися Господа, Бога твого, ходити всіма Його дорогами, і любити Його, і служити Господеві, Богу твоєму, усім серцем своїм і всією душею своєю,
DEUT|10|13|виконувати заповіді Господа та постанови Його, що я наказую тобі сьогодні, щоб було тобі добре.
DEUT|10|14|Тож належить Господеві, Богу твоєму, небо, і небо небес, земля й усе, що на ній.
DEUT|10|15|Тільки батьків твоїх уподобав Господь, щоб любити їх, і вибрав вас, їхнє насіння по них, зо всіх народів, як бачиш цього дня.
DEUT|10|16|І ви обріжете крайню плоть свого серця, а шиї своєї не зробите більше твердою,
DEUT|10|17|бо Господь, Бог ваш Він Бог богів і Пан панів, Бог великий, сильний, та страшний, що не подивиться на обличчя, і підкупу не візьме.
DEUT|10|18|Він чинить суд сироті та вдові, і любить приходька, щоб дати йому хліба й одежу.
DEUT|10|19|І будете ви любити приходька, бо приходьками були ви самі в єгипетськім краї.
DEUT|10|20|Господа, Бога свого, будеш любити, Йому будеш служити, і до Нього будеш горнутись, а Йменням Його будеш присягати.
DEUT|10|21|Він хвала твоя, і Він Бог твій, що з тобою зробив був великі та страшні діла, які бачили очі твої.
DEUT|10|22|Сімдесятьма душами зійшли були твої батьки до Єгипту, а тепер, щодо численности, Господь, Бог твій, зробив тебе, як зорі на небі!
DEUT|11|1|І будеш ти любити Господа, Бога свого, і будеш додержувати постанови Його, і звичаї Його і закони Його, і заповіді Його по всі дні.
DEUT|11|2|І ви пізнаєте сьогодні, бо я навчаю не синів ваших, які не пізнали й не бачили карання Господа, Бога вашого, величність Його, руку Його сильну й рамено Його витягнене,
DEUT|11|3|і ознаки Його, і чини Його, що зробив був серед Єгипту фараонові, єгипетському цареві та всьому його краєві,
DEUT|11|4|і що Він зробив був війську Єгипта, коням його та колесницям його, що пустив над ними воду Червоного моря, коли вони гнались за вами, і вигубив їх Господь, і так є аж до дня цього,
DEUT|11|5|і що Він зробив був для вас у пустині аж до вашого приходу до цього місця,
DEUT|11|6|і що Він зробив був Датанові й Авіронові, синам Еліява, Рувимового сина, що земля відкрила була свої уста й поглинула їх, і їхні доми, і їхні намети, і всю власність, що була з ними, посеред усього Ізраїля.
DEUT|11|7|Бо очі ваші то ті, що бачили всякий великий чин Господа, що Він зробив.
DEUT|11|8|І будете ви виконувати всі заповіді Його, що я сьогодні наказую, щоб стали ви сильні, і ввійшли, і заволоділи тим Краєм, куди переходите ви, щоб посісти його,
DEUT|11|9|і щоб довго жили ви на тій землі, що Господь присягнув був вашим батькам дати їм та їхньому насінню Край, що тече молоком та медом.
DEUT|11|10|Бо цей Край, куди входиш ти заволодіти ним, він не такий, як єгипетський край, звідки вийшли ви, де ти засієш було насіння своє й поливаєш працею ніг своїх, як город варивний.
DEUT|11|11|А цей Край, куди ви переходите посісти його, то край гір та долин, із небесного дощу він напоюється.
DEUT|11|12|Край, що про нього дбає Господь, Бог твій, завжди на ньому очі Господа, Бога твого, від початку року аж до кінця року.
DEUT|11|13|І станеться, якщо справді ви будете слухати Моїх заповідей, що Я вам сьогодні наказую, любити Господа, Бога вашого, і служити Йому всім вашим серцем і всією вашою душею,
DEUT|11|14|то Я дам вам дощ вашого Краю своєчасно, дощ ранній і дощ пізній, і збереш ти своє збіжжя, і свій сік виноградний, і оливу свою.
DEUT|11|15|І дам Я траву на твоїм полі для твоєї худоби, і будеш ти їсти й наситишся.
DEUT|11|16|Стережіться, щоб не було зведене ваше серце, і щоб ви не відступили, і не служили іншим богам, і не вклонялися їм.
DEUT|11|17|А то запалиться гнів Господній на вас, і замкне небо, і не буде дощу, а земля не дасть свого урожаю, і ви скоро погинете з тієї доброї землі, що Господь дає вам.
DEUT|11|18|І покладете ви ці слова Мої на свої серця та на свої душі, і прив'яжете їх на знака на руці своїй, і вони будуть пов'язкою між вашими очима.
DEUT|11|19|І будете навчати про них синів своїх, говорячи про них, коли ти сидітимеш у домі своїм, і коли ходитимеш дорогою, і коли лежатимеш, і коли вставатимеш.
DEUT|11|20|І ти понаписуєш їх на бічних одвірках дому свого і на брамах своїх,
DEUT|11|21|щоб дні ваші та дні синів ваших на землі, яку Господь присягнув був батькам вашим дати їм, були такі довгі, як дні неба над землею.
DEUT|11|22|Бо якщо будете ви конче виконувати всі ті заповіді, що я наказав вам чинити їх, щоб любити Господа, Бога свого, щоб ходити всіма дорогами Його, і щоб горнутись до Нього,
DEUT|11|23|то Господь вижене всі ті народи перед вами, і ви посядете народи більші й міцніші від вас.
DEUT|11|24|Кожне місце, що на нього ступить ваша нога, буде ваше. Від пустині й Ливану, від Річки, річки Ефрату й аж до моря Останнього буде ваша границя.
DEUT|11|25|Не встоїть ніхто перед вами, ляк перед вами й страх перед вами дасть Господь, Бог ваш, на кожен той край, що ви ступите на нього, як Він говорив вам.
DEUT|11|26|Ось, сьогодні я даю перед вами благословення й прокляття:
DEUT|11|27|благословення, коли будете слухатися заповідей Господа, Бога вашого, які я наказую вам сьогодні,
DEUT|11|28|і прокляття, якщо не будете слухатися заповідей Господа, Бога свого, і збочите з дороги, яку я наказую вам сьогодні, щоб ходити за іншими богами, яких ви не знали.
DEUT|11|29|І станеться, коли Господь, Бог твій, уведе тебе до Краю, куди ти входиш посісти його, то даси благословення на горі Ґарізім, а прокляття на горі Евал.
DEUT|11|30|От вони на тому боці Йордану за дорогою заходу сонця, у краю ханаанеянина, що сидить у степу навпроти Ґілґалу при діброві Море.
DEUT|11|31|Бо ви переходите Йордан, щоб увійти посісти той Край, що дає вам Господь, Бог ваш. І посядете його, й осядете в ньому,
DEUT|11|32|і будете додержувати, щоб виконувати всі постанови й закони Його, які я сьогодні даю вам.
DEUT|12|1|Оце постанови та закони, які ви пильнуватимете виконувати в Краї, що дав Господь, Бог батьків твоїх, на насліддя його всі дні, які житимете на цій землі.
DEUT|12|2|Конче винищите всі ті місця, що служили там люди, яких ви виганяєте, своїм богам на високих горах і на пагірках, та під кожним зеленим деревом.
DEUT|12|3|І розвалите їхні жертівники, і поламаєте камінні стовпи для богів, і їхні святі дерева попалите в огні, а бовванів їхніх богів порубаєте, і вигубите їхнє ймення з того місця.
DEUT|12|4|Не робитимете так Господеві, вашому Богові,
DEUT|12|5|бо тільки на місці, яке вибере Господь, Бог ваш, зо всіх ваших племен, щоб покласти там Ім'я Своє, на місці перебування Його будете шукати, і ти прийдеш туди.
DEUT|12|6|І принесете туди свої цілопалення, і свої жертви, і свої десятини та приношення рук своїх, і обітниці свої, і дари свої, і перворідних худоби своєї великої та худоби своєї дрібної.
DEUT|12|7|І будете їсти там перед лицем Господа, Бога вашого, і будете тішитися всім, до чого доторкнеться ваша рука, ви та доми ваші, якими поблагословив тебе Господь, Бог твій.
DEUT|12|8|Там ви не зробите так, як ми робимо сьогодні тут, кожен усе, що йому здається справедливим в очах тільки його,
DEUT|12|9|бо ви дотепер не ввійшли до місця відпочинку й до спадщини, що Господь, Бог твій, дає тобі.
DEUT|12|10|А коли ви перейдете Йордан і осядете в Краї, що Господь, Бог ваш, дає вам на спадщину, і Він заспокоїть вас від усіх ворогів ваших навколо, і ви сидітимете безпечно,
DEUT|12|11|то станеться, на те місце, що його вибере Господь, Бог ваш, щоб Ім'я Його перебувало там, туди принесете все, що я вам наказую: свої цілопалення, і свої жертви, десятини свої та приношення рук своїх, і всі добірні жертви обітниць своїх, що обіцяєте Господеві.
DEUT|12|12|І будете тішитися перед лицем Господа, Бога вашого, ви й сини ваші, і дочки ваші, і раби ваші, і невільниці ваші, і Левит, що в ваших брамах, бо нема йому частки й спадку з вами.
DEUT|12|13|Стережися, щоб не приносив ти своїх цілопалень на кожному місці, яке побачиш,
DEUT|12|14|бо тільки на тому місці, яке вибере Господь в одному з племен твоїх, там принесеш свої цілопалення, і там зробиш усе, що я наказую тобі.
DEUT|12|15|Але скільки запрагне душа твоя, будеш різати й будеш їсти м'ясо, за благословенням Господа, Бога твого, що його дав тобі в усіх брамах твоїх; нечистий і чистий буде їсти його, як сарну й як оленя.
DEUT|12|16|Тільки крови не їстимеш, на землю виллєш її, як воду.
DEUT|12|17|Не зможеш ти їсти в брамах своїх десятини збіжжя свого, і соку виноградного свого, і оливи своєї, і перворідних худоби своєї великої й худоби своєї дрібної, і всіх обітниць своїх, що будеш обіцяти, і добровільних дарів своїх, і приношення своєї руки,
DEUT|12|18|бо тільки перед лицем Господа, Бога свого, будеш їсти його в місці, яке вибере Господь, Бог твій, ти, і син твій, і дочка твоя, і раб твій, і невільниця твоя, і Левит, що в брамах твоїх. І будеш ти радіти перед лицем Господа, Бога свого, усім, до чого доторкнеться рука твоя.
DEUT|12|19|Стережися, щоб не залишив ти Левита по всі дні на землі своїй.
DEUT|12|20|Коли Господь, Бог твій, поширить границю твою, як Він говорив тобі, і ти скажеш: Нехай я їм м'ясо, бо буде жадати душа твоя їсти м'ясо, то за всім жаданням душі своєї будеш ти їсти м'ясо.
DEUT|12|21|Коли буде далеке від тебе те місце, що вибере Господь, Бог твій, щоб перебувало там Ім'я Його, то заріжеш із худоби своєї великої та з худоби своєї дрібної, щоб дав Господь тобі, як наказав я тобі, і будеш їсти в брамах своїх усім жаданням своєї душі.
DEUT|12|22|Тільки як їсться сарну й оленя, так будеш їсти його, нечистий та чистий однаково можуть їсти його.
DEUT|12|23|Тільки будь обережним, щоб не їсти крови, бо кров вона душа, і ти не будеш їсти душі разом з м'ясом.
DEUT|12|24|Не будеш їсти її, на землю виллєш її, як воду.
DEUT|12|25|Не будеш їсти її, щоб було добре тобі та синам твоїм по тобі, коли робитимеш справедливе в Господніх очах.
DEUT|12|26|Тільки святощі свої, що будуть у тебе, та обітниці свої понесеш, і прийдеш до місця, яке вибере Господь.
DEUT|12|27|І принесеш своє цілопалення, м'ясо та кров, на жертівнику Господа, Бога свого, а кров твоїх інших жертов буде вилита на жертівнику Господа, Бога твого, а м'ясо будеш їсти.
DEUT|12|28|Виконуй і слухай усі ті слова, що я наказую тобі, щоб було добре тобі та синам твоїм по тобі навіки, коли будеш робити добре та справедливе в очах Господа, Бога свого.
DEUT|12|29|Коли Господь, Бог твій, вигубить народи, куди ти входиш, щоб посісти їх перед собою, і посядеш їх, і осядеш у їхньому Краї,
DEUT|12|30|то стережися, щоб не впасти до пастки за ними, коли вони будуть вигублені перед тобою, і щоб не шукав ти їхніх богів, говорячи: Як служать ті люди богам своїм, то зроблю так і я.
DEUT|12|31|Не зробиш так Господеві, Богу своєму; бо всяку гидоту, яку Господь зненавидів, робили вони богам своїм, бо навіть синів своїх та дочок своїх вони палять в огні для богів своїх.
DEUT|12|32|(13-1) Кожне слово, що я наказую його вам, будете додержувати виконувати, не додаси до нього, і не відіймеш від нього.
DEUT|13|1|(13-2) Якщо повстане серед тебе пророк або сновидець, і дасть тобі ознаку або чудо,
DEUT|13|2|(13-3) і збудеться та ознака й те чудо, що сказав він тобі, до того говорячи: Ходімо ж за іншими богами, яких ти не знав, і будемо їм служити,
DEUT|13|3|(13-4) то не слухайся слів того пророка або того сновидця, бо цим Господь, Бог ваш, випробовує вас, щоб пізнати, чи ви любите Господа, Бога вашого, усім своїм серцем і всією своєю душею.
DEUT|13|4|(13-5) За Господом, Богом вашим, будете ходити, і Його будете боятися, і заповіді його будете виконувати, і голосу Його будете слухатися, і Йому будете служити, і до Нього будете линути.
DEUT|13|5|(13-6) А пророк той або той сновидець нехай буде забитий, бо намовляв на відступство від Господа, Бога вашого, що вивів вас із єгипетського краю й викупив вас з дому рабства, щоб звести тебе з дороги, що наказав тобі Господь, Бог твій, ходити нею; і вигубиш зло з-посеред себе.
DEUT|13|6|(13-7) Коли намовить тебе брат твій, син твоєї матері, або син твій, або дочка твоя, або жінка твого лоня, або твій приятель, який тобі як душа твоя, таємно говорячи: Ходімо ж і служім іншим богам, яких не знав ти та батьки твої,
DEUT|13|7|(13-8) з богів тих народів, що навколо вас, близьких тобі або далеких від тебе, від кінця землі й аж до кінця землі,
DEUT|13|8|(13-9) то не будеш згоджуватися з ним і не будеш слухатися його, і не буде милосердитися око твоє над ним, і не змилосердишся й не сховаєш його,
DEUT|13|9|(13-10) бо конче заб'єш ти його, рука твоя буде на ньому найперше, щоб забити його, рука всього народу наостанку.
DEUT|13|10|(13-11) І закидаєш його камінням, і він помре, бо жадав відвернути тебе від Господа, Бога твого, що вивів тебе з єгипетського краю, з дому рабства.
DEUT|13|11|(13-12) А ввесь Ізраїль буде слухати і буде боятись, і більше не буде робити такої злої речі серед тебе.
DEUT|13|12|(13-13) Коли почуєш про одне з своїх міст, яке Господь, Бог твій, дає тобі, щоб сидіти там, що про нього кажуть:
DEUT|13|13|(13-14) вийшли люди, сини велійяалові, з-поміж тебе, і звели з правдивої дороги мешканців свого міста, кажучи: Ходімо ж, і служім іншим богам, яких ви не знали,
DEUT|13|14|(13-15) то будеш допитуватися, і будеш досліджувати, і будеш добре питати, а ось воно правда, дійсна та річ, була зроблена та гидота посеред тебе,
DEUT|13|15|(13-16) то конче вибий мешканців того міста вістрям меча, віддай на закляття його й усе, що в ньому, та худобу його вибий вістрям меча.
DEUT|13|16|(13-17) А всю здобич його збереш до середини майдану його, і спалиш огнем те місто та всю здобич його цілковито для Господа, Бога твого. І стане воно купою руїн навіки, не буде вже воно відбудоване.
DEUT|13|17|(13-18) І нічого з закляття нехай не прилипне до руки твоєї, щоб відвернувся Господь від палючого гніву Свого й дав тобі милосердя, і змилосердився над тобою, і розмножив тебе, як присягнув був батькам твоїм,
DEUT|13|18|(13-19) коли будеш слухатися голосу Господа, Бога свого, щоб виконувати всі заповіді Його, що я сьогодні наказую тобі, щоб виконувати те, що справедливе в очах Господа, Бога твого.
DEUT|14|1|Ви сини Господа, Бога вашого, не будете робити нарізів, і не вистригайте волосся над вашими очима за померлого,
DEUT|14|2|бо ти святий народ для Господа, Бога твого, і Господь тебе вибрав, щоб був ти Йому вибраним народом зо всіх народів, що на поверхні землі.
DEUT|14|3|Не будеш їсти жодної гидоти.
DEUT|14|4|Оце та худоба, що ви будете їсти: віл, кожне з овець і кожне з кіз,
DEUT|14|5|олень, і сарна, і буйвіл, і ланя, і зубр, і антилопа, і жирафа.
DEUT|14|6|Кожну з худоби, що має розділені копита та що має копита, роздвоєні розривом, що жує жуйку між худобою, те будете їсти.
DEUT|14|7|Тільки цього не будете їсти з тих, що жують жуйку й що мають розділені копита, розщіплені: верблюда, і зайця, і тушканчика, бо вони жують жуйку, та копит не розділили, нечисті вони для вас.
DEUT|14|8|І свині, бо має розділені ратиці, а жуйки не жує, нечиста вона для вас: їхнього м'яса не будете їсти, а до їхнього падла не доторкнетеся.
DEUT|14|9|Оце будете їсти зо всього, що в воді, усе, що має плавці та луску, будете їсти.
DEUT|14|10|А все, що не має плавців та луски, не будете їсти, нечисте воно для вас.
DEUT|14|11|Кожного чистого птаха будете їсти.
DEUT|14|12|А оце, чого з них ви не будете їсти: орла, і ґрифа, і морського орла,
DEUT|14|13|і коршака, і сокола за родом його,
DEUT|14|14|і всякого крука за родом його,
DEUT|14|15|і струся, і сови, і яструба за родом його,
DEUT|14|16|пугача, й ібіса, і лебедя,
DEUT|14|17|і пелікана, і сича, і рибалки,
DEUT|14|18|і бусла, і чаплі за родом її, і одуда, і кажана.
DEUT|14|19|І кожне плазуюче з птаства нечисте воно для вас, не будете їсти.
DEUT|14|20|Кожного чистого птаха будете їсти.
DEUT|14|21|Не будете їсти жодного падла, даси його приходькові, що в брамах твоїх, і він їстиме його, або продаси чужинцеві, бо ти народ святий для Господа, Бога свого. Не будеш варити ягняти в молоці матері його.
DEUT|14|22|Конче даси десятину з усього врожаю насіння твого, що рік-річно на полі зросте.
DEUT|14|23|І будеш ти їсти перед лицем Господа, Бога свого, у місці, яке Він вибере, щоб Ім'я Його перебувало там, десятину збіжжя свого, виноградного соку свого, і оливки своєї, і перворідних худоби своєї великої й худоби своєї дрібної, щоб навчився ти боятися Господа, Бога свого, по всі дні.
DEUT|14|24|А коли дорога буде занадто довга для тебе, так що не зможеш понести того, бо буде занадто далеке від тебе місце, яке вибере Господь, Бог твій, щоб покласти Ім'я Своє там, коли поблагословить тебе Господь, Бог твій,
DEUT|14|25|то даси в сріблі, і зав'яжеш те срібло в руці своїй, і підеш до місця, яке вибере Господь, Бог твій.
DEUT|14|26|І витратиш те срібло на все чого буде жадати душа твоя, на худобу велику й худобу дрібну, і на вино, і на п'янкий напій, і на все, чого зажадає від тебе душа твоя, і будеш ти їсти там перед лицем Господа, Бога свого, і будеш тішитися ти та дім твій.
DEUT|14|27|А Левит, що живе по брамах твоїх, не кидай його, бо нема йому частки й спадку з тобою.
DEUT|14|28|На кінці трьох років відділиш усю десятину свого врожаю в тім році, і покладеш у брамах своїх.
DEUT|14|29|І прийде Левит, бо нема йому частки й спадку з тобою, і приходько, і сирота, і вдова, що в брамах твоїх, і будуть їсти й наситяться, щоб поблагословив тебе Господь, Бог твій, у кожному чині твоєї руки, що будеш робити.
DEUT|15|1|У кінці семи літ зробиш відпущення.
DEUT|15|2|А оце те відпущення: кожен позикодавець, що позичає своєму ближньому, не буде натискати на свого ближнього та на брата свого, бо оголошено відпущення ради Господа.
DEUT|15|3|На чужинця будеш натискати, а що буде твоє в брата твого, те відпустить йому рука твоя,
DEUT|15|4|та тільки не буде серед тебе вбогого, бо конче поблагословить тебе Господь у Краї, якого Господь, Бог твій, дає тобі на спадок, щоб ти посів його,
DEUT|15|5|якщо тільки конче будеш ти слухатися голосу Господа, Бога свого, щоб додержувати виконувати кожну ту заповідь, що я наказую тобі сьогодні.
DEUT|15|6|Бо Господь, Бог твій, поблагословив тебе, як говорив був тобі, і ти зробиш, що багато людей даватимуть тобі позичку, а ти не даватимеш позички. І будеш ти панувати над багатьма народами, а над тобою не будуть панувати.
DEUT|15|7|Коли буде серед тебе вбогий, один із братів твоїх ув одній із брам твоїх у Краї твоїм, що Господь, Бог твій, дає тобі, то не зробиш запеклим свого серця, і не замкнеш своєї руки від убогого брата свого,
DEUT|15|8|бо конче відкриєш свою руку йому, і конче позичиш йому за його потребою, що буде бракувати йому.
DEUT|15|9|Стережися, щоб у серці твоїм не зродилася зла думка, щоб ти не сказав: Наблизився сьомий рік, рік відпущення, і буде зле твоє око на вбогого брата твого, і не даси ти йому, то він буде кликати на тебе до Господа, і буде на тобі гріх.
DEUT|15|10|Конче даси йому, і нехай не жаліє твоє серце, коли ти даватимеш йому, бо за ту річ поблагословить тебе Господь, Бог твій у кожнім чині твоїм, і в усьому, до чого доторкнеться рука твоя.
DEUT|15|11|Бо не передеться убогий з-посеред Краю, тому я наказую тобі, говорячи: Конче відкривай руку свою для брата свого, і вбогого свого, і для незаможного свого в Краї своїм.
DEUT|15|12|Коли буде проданий тобі брат твій єврей або єврейка, то буде служити тобі шість літ, а сьомого року відпустиш його вільним від себе.
DEUT|15|13|А коли відпустиш його вільним від себе, не відпустиш його порожньо,
DEUT|15|14|конче наділи його з худоби своєї дрібної, і з току свого, і з кадки чавила свого, чим поблагословив тебе Господь, Бог твій, те даси йому.
DEUT|15|15|І будеш пам'ятати, що рабом був ти сам у єгипетськім краї, та викупив тебе Господь, Бог твій, тому я наказую тобі про цю річ сьогодні.
DEUT|15|16|І станеться, коли він скаже тобі: Не вийду від тебе, бо полюбив я тебе та дім твій, бо добре йому з тобою,
DEUT|15|17|то візьмеш шило та й проколеш його вухо до дверей, і стане він тобі вічним рабом; і невільниці своїй зробиш так само.
DEUT|15|18|Нехай не буде тобі тяжким в очах твоїх те, що ти відпускаєш його вільним від себе, бо наємницьку платню він відробив тобі вдвоє за шість літ, і поблагословить тебе Господь, Бог твій, у всім, що ти робитимеш.
DEUT|15|19|Кожного перворідного самця, що народиться в худобі твоїй великій та в худобі твоїй дрібній, посвятиш Господеві, Богові своєму. Не будеш працювати перворідним вола свого, і не будеш стригти перворідного отари своєї.
DEUT|15|20|Перед лицем Господа, Бога свого, рік-річно будеш його їсти ти та дім твій у місці, яке вибере Господь.
DEUT|15|21|А коли буде в нім вада, кульгаве або сліпе, усяка зла вада, то не принесеш його в жертву для Господа, Бога свого,
DEUT|15|22|у брамах своїх будеш його їсти, нечистий і чистий разом, як сарну й як оленя.
DEUT|15|23|Тільки крови його не будеш їсти, на землю виллєш її, як воду.
DEUT|16|1|Додержуй місяця авіва, і справиш Пасху для Господа, Бога свого, бо в місяці авіві вивів тебе Господь, Бог твій, з Єгипту вночі.
DEUT|16|2|І заколи пасху для Господа, Бога свого, з худоби дрібної та з худоби великої в місці, яке вибере Господь, щоб там перебувало Ім'я Його.
DEUT|16|3|Не будеш їсти при тому квашеного, сім день будеш їсти при тому опрісноки, хліб бідування, бо в поспіху вийшов ти з єгипетського краю, щоб усі дні життя свого пам'ятати день свого виходу з єгипетського краю.
DEUT|16|4|І не буде бачене в тебе квашене сім день у всім краї твоїм. А з м'яса, що заколеш у жертву ввечері першого дня, ніщо не буде ночувати до ранку.
DEUT|16|5|Не будеш заколювати пасху в одному з тих твоїх міст, які Господь, Бог твій дає тобі.
DEUT|16|6|Але тільки на тому місці, яке вибере Господь, Бог твій, щоб там перебувало Ім'я Його, заколеш пасху ввечері, при заході сонця, у час твого виходу з Єгипту.
DEUT|16|7|І будеш варити, і будеш їсти на тому місці, яке вибере Господь, Бог твій. А рано обернешся, і підеш до наметів своїх.
DEUT|16|8|Шість день будеш їсти опрісноки, а сьомого дня віддання свята для Господа, Бога твого, не будеш робити зайняття.
DEUT|16|9|Сім тижнів відлічиш собі, від початку праці серпа на дозрілому збіжжі зачнеш лічити сім тижнів.
DEUT|16|10|І справиш свято Тижнів для Господа, Бога свого, у міру добровільного дару своєї руки, що нею даси, як поблагословить тебе Господь, Бог твій.
DEUT|16|11|І будеш радіти перед лицем Господа, Бога свого, ти, і син твій, і дочка твоя, і раб твій, і невільниця твоя, і Левит, що в брамах твоїх, і приходько, і сирота, і вдова, що серед тебе в місці, яке вибере Господь, Бог твій, щоб там перебувало Ім'я Його.
DEUT|16|12|І будеш пам'ятати, що ти сам був рабом в Єгипті, і будеш додержувати це, і будеш виконувати ці постанови.
DEUT|16|13|Свято Кучок будеш справляти собі сім день, коли збереш з току свого та з кадки чавила свого.
DEUT|16|14|І будеш радіти в святі своїм ти, і син твій, і дочка твоя, і раб твій, і невільниця твоя, і Левит, і приходько, і сирота, і вдова, що в брамах твоїх.
DEUT|16|15|Сім день будеш святкувати Господеві, Богові своєму, у місці, яке вибере Господь, бо поблагословить тебе Господь, Бог твій, у всім урожаї твоїм, і в усякім чині рук твоїх, і ти будеш тільки радісний.
DEUT|16|16|Три рази в році вся чоловіча стать буде з'являтися перед лице Господа, Бога твого, у місці, яке Він вибере: у свято Опрісноків, і в свято Тижнів, і в свято Кучок, і ніхто не буде бачений перед лицем Господнім упорожні,
DEUT|16|17|кожен принесе дар руки своєї, за благословенням Господа, Бога свого, що дав Він тобі.
DEUT|16|18|Суддів та урядників настановиш собі в усіх містах своїх, які Господь, Бог твій, дає тобі по племенах твоїх, і вони будуть судити народ справедливим судом.
DEUT|16|19|Не викривиш закону, не будеш дивитися на особу, і не візьмеш підкупу, бо підкуп осліплює очі мудрих і викривлює слова справедливих.
DEUT|16|20|За справедливістю, лише за справедливістю будеш гнатися, щоб жити й заволодіти Краєм, що Господь, Бог твій, дає тобі.
DEUT|16|21|Не посадиш собі святого дерева, усякого дерева при жертівнику Господа, Бога твого, що зробиш собі,
DEUT|16|22|і не поставиш собі стовпа, що ненавидить Господь, Бог твій.
DEUT|17|1|Не будеш приносити в жертву Господеві, Богові своєму вола або одне з дрібної худоби, що буде на ньому вада, усяка зла річ, бо це гидота для Господа, Бога твого.
DEUT|17|2|Коли буде знайдений серед тебе в одному з міст твоїх, які Господь, Бог твій, дає тобі, чоловік або жінка, що зробить зле в очах Господа, Бога твого, щоб недотримати заповіту,
DEUT|17|3|що пішов би й служив би іншим богам, і вклонявся б їм та сонцеві або місяцеві, або всім зорям небесним, чого я не наказав,
DEUT|17|4|і буде розказано тобі, і ти почуєш, і будеш добре допитуватися, а ото воно правда, дійсна та річ, була зроблена ота гидота серед Ізраїля,
DEUT|17|5|то випровадиш того чоловіка або ту жінку, що зробили ту злу річ, до брам своїх, того чоловіка або ту жінку, і вкаменуєш їх камінням, і вони погинуть.
DEUT|17|6|На слова двох свідків або трьох свідків буде забитий обвинувачений, що має померти; на слова одного свідка не буде забитий.
DEUT|17|7|Рука свідків буде на ньому найперше, щоб забити його, а рука всього народу наостанку. І вигубиш зло з-посеред себе.
DEUT|17|8|Коли б у суді була тобі неясна справа між кров'ю та кров'ю, між суперечкою та суперечкою, і між раною та раною справи суперечки в брамах твоїх, то встанеш, і підеш до місця, яке вибере його Господь, Бог твій.
DEUT|17|9|І прийдеш до священиків-Левитів і до судді, що буде в тих днях, і допитаєшся, і вони дадуть тобі слово присуду.
DEUT|17|10|І ти поступиш за тим словом, що подадуть тобі з того місця, яке вибере Господь, і будеш пильнувати робити все так, як навчать тебе.
DEUT|17|11|Ти поступиш за законом, що навчать тебе, і за вироком, що скажуть тобі, не відступиш ні праворуч ні ліворуч від слова, що подадуть тобі.
DEUT|17|12|А коли хто через зухвалість не послухається священика, що стоїть там на служенні Господеві, Богові твоєму, або судді, то помре той, і вигубиш те зло з Ізраїля.
DEUT|17|13|А ввесь народ буде слухати та буде боятися, і вже не буде поступати зухвало.
DEUT|17|14|Коли ти ввійдеш до того Краю, що Господь, Бог твій, дає тобі, і посядеш його, і осядеш у ньому, та й скажеш: Нехай я поставлю над собою царя, як усі народи, що в моїх околицях,
DEUT|17|15|то, ставлячи над собою царя, якого вибере Господь, Бог твій, конче з-посеред братів своїх поставиш над собою царя, не зможеш поставити над собою чоловіка чужинця, що він не брат твій.
DEUT|17|16|Тільки щоб він не примножував собі коней, і не вертав народу до Єгипту, щоб примножити коней, бож Господь сказав вам: Не вертайтеся вже більше тією дорогою.
DEUT|17|17|І хай не примножить він собі жінок, щоб не відступило його серце, і срібла та золота хай він не примножить собі дуже.
DEUT|17|18|І станеться, як буде він сидіти на троні царства свого, то напише собі відписа цього Закону з книги, що перед лицем священиків-Левитів.
DEUT|17|19|І буде вона з ним, і буде він читати в ній усі дні свого життя, щоб учився боятися Господа, Бога свого, щоб додержувати всіх слів цього Закону та тих постанов, щоб виконувати їх,
DEUT|17|20|щоб не гордувало серце його своїми братами, і щоб не збочував він ні праворуч, ні ліворуч від цієї заповіді, щоб продожив дні на своїм царстві він та сини його серед Ізраїля.
DEUT|18|1|Священикам-Левитам, усьому Левієвому племені не буде частки та спадку разом з Ізраїлем, огняні жертви Господа та частки Його будуть їм.
DEUT|18|2|А спадку не буде йому серед братів його: Господь Він спадок його, як Він говорив був йому.
DEUT|18|3|А оце буде належати священикам від народу, від тих, хто приносить жертву: коли це віл, коли це одне з дрібної худоби, то даси священикові плече, і щоки, і шлунок.
DEUT|18|4|Початок від збіжжя свого, від виноградного соку свого, і від оливки своєї, і початок стриження отари своєї даси ти йому.
DEUT|18|5|Бо його вибрав Господь, Бог твій, зо всіх племен твоїх, щоб ставав він служити в Господнє Ім'я, він та сини його по всі дні.
DEUT|18|6|А коли прийде Левит з одної з брам твоїх з усього Ізраїля, де він мешкає там, і прибуде за всім жаданням своєї душі до місця, яке вибере Господь,
DEUT|18|7|і буде він служити в Ім'я Господа, Бога свого, як усі його браття Левити, що стоять там перед Господнім лицем,
DEUT|18|8|то по рівній частці будуть вони їсти, опріч маєтку, проданого по батьках.
DEUT|18|9|Коли будеш входити до Краю, що дає тобі Господь, Бог твій, то не навчися чинити такого, як гидота цих народів.
DEUT|18|10|Нехай не знайдеться між тобою такий, хто переводить свого сина чи дочку свою через огонь, хто ворожить ворожбу, хто ворожить по хмарах, і хто ворожить по птахах, і хто чарівник,
DEUT|18|11|і хто чорнокнижник, і хто викликає духа померлого та духа віщого, і хто питає померлих.
DEUT|18|12|Бо гидота для Господа кожен, хто чинить таке, і через ті гидоти Господь, Бог твій, виганяє їх перед тобою.
DEUT|18|13|Бездоганний будеш ти перед Господом, Богом своїм,
DEUT|18|14|бо ці народи, що ти посядеш їх, слухають тих, хто ворожить по хмарах та ворожбитів, а ти не таке дав тобі Господь, Бог твій.
DEUT|18|15|Пророка з-посеред тебе, з братів твоїх, Такого, як я, поставить тобі Господь, Бог твій, Його будете слухати,
DEUT|18|16|згідно з усім, чого жадав ти від Господа, Бога свого, на Хориві в дні зборів, говорячи: Щоб більше не чути мені голосу Господа, Бога свого, а цього великого огню вже не побачити й не померти.
DEUT|18|17|І сказав до мене Господь: Добре сказали вони.
DEUT|18|18|Поставлю Пророка для них з-поміж їхніх братів, Такого, як ти, і дам Я слова Свої в уста Його, і Він їм говоритиме все, що Я накажу.
DEUT|18|19|І станеться, кожен, хто не слухатиме слів Моїх, що Той Пророк говоритиме Моїм Ім'ям, Я покараю того.
DEUT|18|20|А той пророк, що зухвало відважиться промовляти Моїм Ім'ям слова, яких Я не наказав був йому говорити, і що буде говорити, і що буде говорити ім'ям інших богів, хай помре той пророк.
DEUT|18|21|А коли ти скажеш у серці своєму: Як ми пізнаємо те слово, якого Господь не говорив?
DEUT|18|22|Що буде говорити той пророк Ім'ям Господа, і не станеться та річ, і не прийде, то це те слово, якого не сказав Господь. У зухвалості говорив його той пророк, і ти не будеш боятися його.
DEUT|19|1|Коли Господь, Бог твій, повигублює народи, що Господь, Бог твій, дає тобі їхній Край, і ти повиганяєш їх, і осядеш по їхніх містах та по їхніх домах,
DEUT|19|2|то три місті відділиш собі в середині свого Краю, що Господь, Бог твій, дає його тобі на володіння.
DEUT|19|3|Приготуєш собі дорогу, і поділиш натроє землю твого Краю, що Господь, Бог твій, дає тобі на спадок, і це буде на втікання туди кожного убійника.
DEUT|19|4|А оце справа убійника, що втече туди й буде жити: хто вб'є свого ближнього ненароком, а він не був ворогом його від учора й позавчора;
DEUT|19|5|або хто ввійде з своїм ближнім до лісу рубати дерева, і розмахнеться рука його з сокирою, щоб зрубати дерево, а залізо спаде з топорища й попаде в його ближнього, і той помре, то він утече до одного з тих міст, і буде жити,
DEUT|19|6|щоб не гнався месник за кров за убійником, коли розпалиться серце його, і щоб не догнав його, якщо буде довга та дорога, і не вбив його, хоч він не підлягає смерті, бо не був він ворогом його від учора й позавчора.
DEUT|19|7|Тому то я наказую тобі, говорячи: Три місті відділиш собі.
DEUT|19|8|А якщо Господь, Бог твій, розширить границю твою, як присягнув був батькам твоїм, і дасть тобі всю оцю землю, що говорив був дати батькам твоїм,
DEUT|19|9|коли ти будеш додержувати всі ці заповіді, щоб виконувати їх, що я наказую тобі сьогодні, щоб любити Господа, Бога свого, і щоб ходити дорогами Його всі дні, то додаси собі ще три місті понад ті три,
DEUT|19|10|щоб не була пролита неповинна кров серед твого Краю, що Господь, Бог твій, дає тобі на спадок, і не буде на тобі кров.
DEUT|19|11|А коли хто буде ненавидіти свого ближнього, і буде чатувати на нього, і повстане на нього та й уб'є його, і той помре, і втече він до одного з тих міст,
DEUT|19|12|то пошлють старші його міста, і візьмуть його звідти, і дадуть його в руку месника крови, і він помре.
DEUT|19|13|Не змилосердиться око твоє над ним, і ти усунеш кров неповинного з Ізраїля, і буде добре тобі.
DEUT|19|14|Не пересунеш межі свого ближнього, яку розмежували предки в наділі твоїм, яке посядеш ти в Краю, що Господь, Бог твій, дає його тобі на володіння.
DEUT|19|15|Не стане один свідок на кого для всякої провини і для всякого гріха, у кожнім гріху, що згрішить, на слова двох свідків або на слова трьох свідків відбудеться справа.
DEUT|19|16|Коли стане на кого неправдивий свідок, щоб свідчити проти нього підступно,
DEUT|19|17|то стануть двоє цих людей, що мають суперечку, перед лицем Господнім, перед священиками та суддями, що будуть у тих днях.
DEUT|19|18|І судді добре дослідять, а ось свідок неправдивий той свідок, неправду говорив на брата свого,
DEUT|19|19|то зробите йому так, як він замишляв був зробити своєму братові, і вигубиш зло з-посеред себе.
DEUT|19|20|А позосталі будуть слухати, і будуть боятися, і більш вже не будуть робити серед себе такого, як та річ зла.
DEUT|19|21|І не змилосердиться око твоє: життя за життя, око за око, зуб за зуба, рука за руку, нога за ногу.
DEUT|20|1|Коли ти вийдеш на війну проти свого ворога, та побачиш коні й вози, та народ, численніший від тебе, то не будеш боятися їх, бо з тобою Господь, Бог твій, що вивів тебе з єгипетського краю.
DEUT|20|2|І станеться, коли ви приступите до бою, то підійде священик і буде промовляти до народу,
DEUT|20|3|та й скаже до них: Слухай, Ізраїлю, ви приступаєте сьогодні до бою проти ваших ворогів. Нехай не зм'якне серце ваше, не бійтеся, і не страшіться, і не лякайтеся їх,
DEUT|20|4|бо Господь, Бог ваш, Він Той, що йде з вами воювати для вас з вашими ворогами, щоб спасти вас!
DEUT|20|5|А урядники будуть промовляти до народу, говорячи: Хто є тут такий, що збудував новий дім, та не справив обряду поновин? Нехай він іде й вертається до свого дому, щоб не померти на війні, і щоб інший хто не справив на ньому обряду поновин.
DEUT|20|6|І хто є тут такий, що засадив виноградника та не користався ним? Нехай він іде й вертається до свого дому, щоб не померти на війні, і щоб інший хто не скористався ним.
DEUT|20|7|А хто є тут такий, що засватав жінку, та не взяв її? Нехай він іде й вертається до свого дому, щоб не померти на війні, і щоб інший хто не взяв її.
DEUT|20|8|І далі промовлятимуть урядники до народу та й скажуть: Хто є тут такий, що лякливий та м'якосердий? Нехай він іде й вертається до свого дому, щоб не розслабив він серця братів своїх, як є серце його.
DEUT|20|9|І станеться, коли урядники закінчать промовляти до народу, то призначать зверхників для військових відділів на чоло народу.
DEUT|20|10|Коли ти приступиш до міста, щоб воювати з ним, то запропонуй йому перше мир.
DEUT|20|11|І станеться, якщо воно відповість тобі: Мир, і відчинить браму тобі, то ввесь той народ, що знаходиться в ньому, буде тобі на данину, і буде служити тобі.
DEUT|20|12|А якщо воно не замирить з тобою, і буде провадити з тобою війну, то обложиш його.
DEUT|20|13|І Господь, Бог твій, дасть його в руку твою, а ти повбиваєш усю чоловічу стать його вістрям меча.
DEUT|20|14|Тільки жінок, і дітей, і худобу, і все, що буде в тім місті, всю здобич його забереш собі, і будеш ти їсти здобич ворогів своїх, що дав тобі Господь, Бог твій.
DEUT|20|15|Так ти зробиш усім містам, дуже далеким від тебе, що вони не з міст цих народів.
DEUT|20|16|Тільки з міст тих народів, які Господь, Бог твій, дає тобі на володіння, не позоставиш при житті жодної душі,
DEUT|20|17|бо конче вчиниш їх закляттям: Хіттеянина, і Амореянина, і Ханаанеянина, і Періззеянина, і Хіввеянина, і Євусеянина, як наказав був тобі Господь, Бог твій,
DEUT|20|18|щоб вони не навчили вас робити такого, як усі їхні гидоти, що робили вони богам своїм, бо тоді згрішите ви перед Господом, Богом своїм.
DEUT|20|19|Коли будеш облягати місто багато днів, щоб воювати з ним та щоб здобути його, то не знищиш його дерева, і не піднесеш сокири на нього, бо з нього ти їстимеш, і його не будеш стинати, бо чи ж пільне дерево то чоловік, щоб увійти перед тобою до обложеного міста?
DEUT|20|20|Тільки дерево, що про нього ти знаєш, що воно не дерево на їжу, його знищиш та зітнеш, і будеш будувати з нього речі облягання проти того міста, яке провадить з тобою війну, аж до упадку його.
DEUT|21|1|Коли на землі, яку дає тобі Господь, Бог твій на володіння, буде знайдений забитий, що впав на полі, і не буде відомим, хто вбив його,
DEUT|21|2|то повиходять старші твої та судді твої, та й виміряють до тих міст, що навколо забитого.
DEUT|21|3|І станеться, коли довідаються про місто, найближче до забитого, то візьмуть старші того міста телицю з худоби великої, що нею не працьовано, що вона не тягана в ярмі.
DEUT|21|4|І старші того міста зведуть ту телицю до долини висихаючого потоку, що на ньому не орано, і що він не засіюваний, і там у долині висихаючого потоку переріжуть шию тій телиці.
DEUT|21|5|І підійдуть священики, Левієві сини, бо їх вибрав Господь, Бог твій, щоб служили Йому, і щоб благословляли Господнім Ім'ям, і за їхніми словами буде рішатися всяка суперечка та всяка пораза.
DEUT|21|6|І всі старші того міста, найближчі до забитого, умиють свої руки над телицею, що в долині висихаючого потоку їй перерізана шия.
DEUT|21|7|І освідчать вони та й скажуть: Руки наші не пролили цієї крови, а очі наші не бачили.
DEUT|21|8|Прости народові своєму, Ізраїлеві, якого Ти, Господи, викупив, і не дай неповинної крови посеред народу Свого, Ізраїля, І буде прощена їм та кров.
DEUT|21|9|А ти усунеш неповинну кров з-посеред себе, коли робитимеш справедливе в Господніх очах.
DEUT|21|10|Коли ти вийдеш на війну на ворогів своїх, і Господь, Бог твій, дасть їх у твою руку, і ти пополониш із них полонених,
DEUT|21|11|і побачиш серед полонених гарновиду жінку, і вподобаєш її собі, і візьмеш собі за жінку,
DEUT|21|12|то впровадиш її до середини свого дому, а вона оголить свою голову й обітне свої нігті.
DEUT|21|13|І здійме вона з себе одіж полону свого, і осяде в твоєму домі, та й буде оплакувати батька свого та матір свою місяць часу, а по тому ти ввійдеш до неї й станеш їй чоловіком, і вона стане тобі за жінку.
DEUT|21|14|І станеться, коли ти потім не полюбиш її, то відпустиш її за її волею, а продати не продаси її за срібло, і не будеш поводитися з нею як з невільницею, бо ти жив із нею.
DEUT|21|15|Коли хто матиме дві жінки, одна кохана, а одна зненавиджена, і вони вродять йому синів, та кохана й та зненавиджена, і буде перворідний син від зненавидженої,
DEUT|21|16|то станеться того дня, коли він робитиме синів своїх спадкоємцями того, що буде його, то не зможе він зробити перворідним сина тієї коханої за життя того перворідного сина зненавидженої,
DEUT|21|17|але за перворідного визнає сина зненавидженої, щоб дати йому подвійно з усього, що в нього знайдеться, бо він початок сили його, його право перворідства.
DEUT|21|18|Коли хто матиме неслухняного й непокірного сина, що не слухається голосу батька свого та голосу своєї матері, і докорятимуть йому, а він не буде їх слухатися,
DEUT|21|19|то батько його та мати його схоплять його, і приведуть його до старших його міста та до брами того місця.
DEUT|21|20|І скажуть вони до старших міста його: Оцей наш син неслухняний та непокірний, він не слухає голосу нашого, ласун та п'яниця.
DEUT|21|21|І всі люди його міста закидають його камінням, і він помре. І вигубиш те зло з-посеред себе, а ввесь Ізраїль буде слухатися й буде боятися.
DEUT|21|22|А коли буде на кому гріх смертного присуду, і буде він убитий, і ти повісиш його на дереві,
DEUT|21|23|то труп його не буде ночувати на дереві, але конче поховаєш його того дня, бо повішений Боже прокляття, і ти не занечистиш своєї землі, яку Господь, Бог твій, дає тобі на спадок.
DEUT|22|1|Коли побачиш вола свого брата або щось із отари, що заблудили, то ти не сховаєшся від них, а конче вернеш їх своєму братові.
DEUT|22|2|А якщо брат твій не близький до тебе, чи ти не знаєш його, то забереш те до дому свого, і воно буде з тобою, аж поки брат твій не буде шукати його, і повернеш його йому.
DEUT|22|3|І так зробиш ослові його, і так зробиш одежі його, і так зробиш усякій згубі брата свого, що згублена в нього, а ти знайдеш її, не зможеш ховати її.
DEUT|22|4|Коли побачиш осла свого брата або вола його, що впали на дорозі, то ти не сховаєшся від них, конче підіймеш їх разом із ним.
DEUT|22|5|Не буде чоловіча річ на жінці, а мужчина не зодягне жіночої одежі, бо кожен, хто чинить це, огида він для Господа, Бога свого.
DEUT|22|6|Коли спіткається на дорозі пташине кубло перед тобою на якомубудь дереві чи на землі з пташенятами або з яйцями, а мати сидить на пташенятах або на яйцях, то не візьмеш тієї матері з дітьми,
DEUT|22|7|конче відпустиш ту матір, а дітей візьмеш собі, щоб було добре тобі, і щоб ти продовжив свої дні.
DEUT|22|8|Коли збудуєш новий дім, то зробиш поруччя для даху свого, і не напровадиш крови на дім свій, коли спаде з нього хтось.
DEUT|22|9|Не будеш засівати свого виноградника подвійним насінням, щоб не зробити заклятим усе насіння: і що засієш, і врожай виноградника.
DEUT|22|10|Не будеш орати волом і ослом разом.
DEUT|22|11|Не одягнеш одежі з двійного матеріялу, з вовни й льону разом.
DEUT|22|12|Поробиш собі кутаси на чотирьох краях свого покриття, що ним покриваєшся.
DEUT|22|13|Коли хто візьме жінку, і ввійде до неї, але потім зненавидить її,
DEUT|22|14|і зводитиме на неї ганьбливі слова, і пустить про неї неславу та й скаже: Жінку цю взяв я, і зблизився з нею, та не знайшов у неї дівоцтва,
DEUT|22|15|то візьме батько тієї дівчини та мати її, і віднесуть доказа дівоцтва тієї дівчини до старших міста, до брами.
DEUT|22|16|І скаже батько тієї дівчини до старших: Я дав тому чоловікові дочку свою за жінку, та він зненавидів її.
DEUT|22|17|І ось він зводить на неї ганьбливі слова, говорячи: Я не знайшов у твоєї дочки дівоцтва, а оце знаки дівоцтва моєї дочки. І розтягнуть одежу перед старшими міста.
DEUT|22|18|А старші того міста візьмуть того чоловіка, та й покарають його,
DEUT|22|19|і накладуть на нього пеню, сто шеклів срібла, і дадуть батькові тієї дівчини, бо він пустив неславу на Ізраїлеву дівчину, а вона буде йому за жінку, він не зможе відпустити її по всі свої дні.
DEUT|22|20|А якщо правдою було це слово, не знайдене було дівоцтво в тієї дівчини,
DEUT|22|21|то приведуть ту дівчину до дверей дому батька її, і вкаменують її люди її міста камінням, і вона помре, бо зробила негідність між Ізраїлем на спроневірення дому батька свого, і вигубиш зло з-посеред себе.
DEUT|22|22|Коли буде знайдений хто, що лежить із заміжньою жінкою, то помруть вони обоє, той чоловік, що лежав із жінкою, і та жінка, і вигубиш зло з Ізраїля.
DEUT|22|23|Коли дівчина буде заручена чоловікові, і спіткає її хто в місті, і ляже з нею,
DEUT|22|24|то виведете їх обох до брами того міста, і вкаменуєте їх камінням, і вони помруть, ту дівчину за те, що не кричала в місті, а того чоловіка за те, що збезчестив жінку свого ближнього, і вигубиш зло серед себе.
DEUT|22|25|А як хто на полі спіткає заручену дівчину, і схопить її та й ляже з нею, то помре той чоловік, що ліг із нею, він сам,
DEUT|22|26|а тій дівчині не зробиш нічого, нема тій дівчині смертельного гріха, бо це таке, як повстане хто на свого ближнього й уб'є його, така це річ.
DEUT|22|27|Бо в полі він спіткав її, кричала та заручена дівчина, та не було кому врятувати її.
DEUT|22|28|Коли хто спіткає дівчину, що не була заручена, і схопить її, і ляже з нею, і застануть їх,
DEUT|22|29|то той чоловік, що лежав із нею, дасть батькові тієї дівчини п'ятдесят шеклів срібла, і вона стане йому за жінку, за те, що збезчестив її, не зможе він відпустити її по всі свої дні.
DEUT|22|30|(23-1) Ніхто не візьме жінки свого батька, і не відкриє подолка одежі батька свого.
DEUT|23|1|(23-2) Не ввійде на збори Господні ранений розчавленням ятер та з відрізаним членом.
DEUT|23|2|(23-3) Неправоложний не ввійде на збори Господні, також десяте покоління його не ввійде на збори Господні.
DEUT|23|3|(23-4) Не ввійде на збори Господні аммонітянин та моавітянин, також десяте їхнє покоління не ввійде на збори Господні, аж навіки,
DEUT|23|4|(23-5) за те, що вони не вийшли назустріч вас із хлібом та водою в дорозі, коли ви виходили з Єгипту, і що найняли були на тебе Валаама, Беорового сина з Петору Араму двох річок, щоб проклясти тебе.
DEUT|23|5|(23-6) Та не хотів Господь, Бог твій, слухати Валаама, і перемінив тобі Господь, Бог твій, те прокляття на благословення, бо любить тебе Господь, Бог твій.
DEUT|23|6|(23-7) Не будеш бажати для них миру й добра по всі свої дні навіки.
DEUT|23|7|(23-8) Не обридиш собі Ідумеянина, бо він твій брат; не обридиш собі Єгиптянина, бо був ти приходьком у краї його.
DEUT|23|8|(23-9) Сини, що народяться їм, покоління третє ввійде з них на збори Господні.
DEUT|23|9|(23-10) Коли табір вийде на ворогів твоїх, то будеш стерегтися всякої злої речі.
DEUT|23|10|(23-11) Коли поміж тебе буде хто, що буде нечистий з нічної пригоди, то він вийде поза табір, до середини табору не ввійде.
DEUT|23|11|(23-12) А коли наступатиме вечір, обмиється в воді, а по заході сонця ввійде до середини табору.
DEUT|23|12|(23-13) А місце на потребу буде тобі поза табором, щоб виходити тобі туди назовні.
DEUT|23|13|(23-14) А лопатка буде в тебе на поясі твоїм; і станеться, коли ти сидітимеш назовні, то будеш копати нею, і знову закриєш свою нечистість,
DEUT|23|14|(23-15) бо Господь, Бог твій, ходить у середині табору твого, щоб тебе спасати, і видавати ворогів твоїх тобі. І буде табір твій святий, і Він не побачить у тебе соромітної речі, і не відвернеться.
DEUT|23|15|(23-16) Не видавай панові раба його, який сховається до тебе від пана свого.
DEUT|23|16|(23-17) З тобою він сидітиме серед вас у місці, яке він вибере за добре собі в одній з твоїх брам, і ти не будеш гнобити його.
DEUT|23|17|(23-18) Блудниця не буде з Ізраїлевих дочок, і блудодій не буде з Ізраїлевих синів.
DEUT|23|18|(23-19) Не принесеш дару розпусниці й ціни пса до дому Господа, Бога твого, ні за яку обітницю, бо тож вони обоє гидота перед Господом, Богом твоїм.
DEUT|23|19|(23-20) Не будеш позичати братові своєму на відсоток срібла, на відсоток їжі та всякої речі, що позичається на відсоток.
DEUT|23|20|(23-21) Чужому позичиш на відсоток, а братові своєму не позичиш на відсоток, щоб поблагословив тебе Господь, Бог твій у всьому, до чого доторкнеться рука твоя на тій землі, куди ти входиш на володіння її.
DEUT|23|21|(23-22) Коли ти складеш обітницю Господеві, Богові твоєму, не загаюйся виконати її, бо конче буде жадати Господь, Бог твій, від тебе, і буде на тобі гріх.
DEUT|23|22|(23-23) А коли ти не складав обітниці, не буде на тобі гріха.
DEUT|23|23|(23-24) Що вийшло з уст твоїх, будеш додержувати й будеш виконувати, як обіцяв ти Господеві, Богові своєму, добровільну жертву, що промовляв ти своїми устами.
DEUT|23|24|(23-25) Коли ввійдеш до виноградника свого ближнього, то будеш їсти виноград, скільки схоче душа твоя, до свого насичення, а до посуду свого не візьмеш.
DEUT|23|25|(23-26) Коли ти ввійдеш на дозріле збіжжя свого ближнього, то будеш рвати колоски рукою своєю, а серпом не будеш жати на дозрілім збіжжі свого ближнього.
DEUT|24|1|Як хто візьме жінку, і стане їй чоловіком, і коли вона не знайде ласки в очах його, бо знайшов у ній яку ганебну річ, то напише їй листа розводового, і дасть в її руку, та й відпустить її з свого дому.
DEUT|24|2|І вийде вона з його дому, і піде, і вийде за іншого чоловіка,
DEUT|24|3|і коли зненавидить її той останній чоловік, то напише їй листа розводового, і дасть в її руку, та й відпустить її з свого дому. Або коли помре той останній чоловік, що взяв був її собі за жінку,
DEUT|24|4|не може перший її муж, що відпустив її, вернути й узяти її, щоб стала йому за жінку по тому, як була занечищена, бо це огида перед Господнім лицем, і ти не зробиш грішною тієї землі, яку Господь, Бог твій, дає тобі на спадок.
DEUT|24|5|Коли хто недавно одружився, не піде він до війська, і ніяка справа не покладеться на нього, вільний він буде один рік для свого дому, і порадує свою жінку, що взяв.
DEUT|24|6|Ніхто не візьме в заставу долішнього каменя жорен або горішнього каменя жорен, бо він душу взяв би в заставу.
DEUT|24|7|Коли буде хто знайдений, що вкрав кого з братів своїх, з Ізраїлевих синів, і буде поводитися з ним як із невільником, або й продасть його, то нехай помре той злодій, і ти вигубиш зло з-посеред себе.
DEUT|24|8|Стережися в хворобі прокази, щоб дуже пильнувати, і робити все те, як навчать вас священики-Левити; як наказав я їм, будете додержувати, щоб виконати те.
DEUT|24|9|Пам'ятайте те, що зробив був Господь, Бог твій, Маріямі в дорозі, коли ви виходили з Єгипту.
DEUT|24|10|Коли ти позичиш своєму ближньому позичку з чогось, не ввійдеш до дому його, щоб узяти заставу його,
DEUT|24|11|назовні будеш стояти, а той чоловік, що ти позичив йому, винесе до тебе заставу назовні.
DEUT|24|12|А якщо він чоловік убогий, не ляжеш спати, маючи заставу його,
DEUT|24|13|конче вернеш йому ту заставу при заході сонця, і буде він спати на одежі своїй, і буде благословляти тебе, а тобі буде це за праведність перед лицем Господа, Бога твого.
DEUT|24|14|Не будеш утискати наймита, убогого й незаможного з братів своїх та з приходька свого, що в Краї твоїм у брамах твоїх.
DEUT|24|15|Того ж дня даси йому заплату, і не зайде над нею незаплаченою сонце, бо вбогий він, і до неї лине душа його. І не буде він кликати на тебе до Господа, і не буде гріха на тобі.
DEUT|24|16|Не будуть забиті батьки за синів, а сини не будуть забиті за батьків, кожен за гріх свій смертю покараний буде.
DEUT|24|17|Не скривиш суду на приходька, на сироту, і не будеш брати в заставу вдовиної одежі.
DEUT|24|18|І будеш пам'ятати, що рабом був ти сам у Єгипті, і викупив тебе Господь, Бог твій, звідти, тому я наказую тобі робити цю річ.
DEUT|24|19|Коли будеш жати жниво своє на своїм полі, і забудеш на полі снопа, не вернешся взяти його, він буде приходькові, сироті та вдові, щоб поблагословив тебе Господь, Бог твій, у всім чині твоїх рук.
DEUT|24|20|Коли будеш оббивати оливку свою, не будеш переоббивати в галузках за собою: воно буде приходькові, сироті та вдові.
DEUT|24|21|Коли будеш збирати виноград свого виноградника, не будеш збирати полишеного за собою, воно буде приходькові, сироті та вдові.
DEUT|24|22|І будеш пам'ятати, що рабом був ти в єгипетськім краї, тому я наказую тобі робити цю річ.
DEUT|25|1|Коли буде суперечка між людьми, і вони прийдуть до суду, то розсудять їх, і оправдають справедливого, а несправедливого осудять.
DEUT|25|2|І станеться, якщо вартий биття той несправедливий, то покладе його суддя, і буде його бити перед собою, число ударів згідно з його несправедливістю.
DEUT|25|3|Сорока ударами буде його бити, не більше; щоб не бити його більше над те великим биттям, і щоб не був злегковажений брат твій на очах твоїх.
DEUT|25|4|Не зав'яжеш рота волові, коли він молотить.
DEUT|25|5|Коли браття сидітимуть разом, і один із них помре, а сина в нього нема, то жінка померлого не вийде заміж назовні за чужого, дівер її прийде до неї та й візьме її собі за жінку, і подіверує її.
DEUT|25|6|І буде перворідний, що вона породить, стане він ім'ям його брата, що помер, і не буде стерте ім'я його з Ізраїля.
DEUT|25|7|А якщо той чоловік не схоче взяти своєї братової, то братова його вийде до брами до старших та й скаже: Дівер мій відмовився відновити своєму братові ім'я в Ізраїлі, не хотів подіверувати мене.
DEUT|25|8|І покличуть його старші його міста, і промовлятимуть до нього, а він устане та й скаже: Не хочу взяти її,
DEUT|25|9|то підійде його братова до нього на очах старших, і здійме йому чобота з ноги його, і плюне в обличчя його, і заговорить, і скаже: Так робиться чоловікові, що не будує дому свого брата.
DEUT|25|10|І буде зване ім'я його в Ізраїлі: Дім роззутого.
DEUT|25|11|Коли чоловіки будуть сваритися разом один з одним, і підійде жінка одного, щоб оберегти свого чоловіка від руки того, що б'є, і простягне свою руку, і схопить за сором його,
DEUT|25|12|то відрубаєш руку її, нехай не змилосердиться око твоє!
DEUT|25|13|Не буде в тебе в торбі твоїй подвійного каменя до ваги, великого й малого,
DEUT|25|14|не буде тобі в твоїм домі подвійної ефи, великої й малої.
DEUT|25|15|Камінь до ваги буде в тебе повний і справедливий, ефа буде в тебе повна й справедлива, щоб продовжилися дні твої на землі, яку Господь, Бог твій, дає тобі.
DEUT|25|16|Бо огида перед Господом, Богом твоїм, кожен, хто чинить таке, хто чинить несправедливість.
DEUT|25|17|Пам'ятайте, що зробив був тобі Амалик у дорозі, коли ви виходили з Єгипту,
DEUT|25|18|що спіткав тебе в дорозі, і повбивав між тобою всіх задніх ослаблених, коли ти був змучений та струджений, а він не боявся Бога.
DEUT|25|19|І станеться, коли Господь, Бог твій, дасть тобі мир від усіх ворогів твоїх навколо в Краї, що Господь, Бог твій, дає тобі як спадок, щоб посісти його, то зітреш пам'ять Амалика з-під неба. Не забудь!
DEUT|26|1|І станеться, коли ти ввійдеш до того Краю, що Господь, Бог твій, дає тобі як спадок, і посядеш його, і осядеш у ньому,
DEUT|26|2|то візьмеш із початків усякого плоду землі, що збереш із Краю свого, що Господь, Бог твій, дає тобі, і покладеш їх у кіш, та й підеш до місця, яке вибере Господь, Бог твій, щоб там пробувало Ім'я Його.
DEUT|26|3|І прийдеш ти до священика, що буде тими днями, та й скажеш йому: Засвідчую це сьогодні Господеві, Богові твоєму, що я ввійшов до Краю, що Господь заприсягнув був батькам нашим, щоб дати нам.
DEUT|26|4|І візьме священик того коша з твоєї руки, і покладе його перед жертівником Господа, Бога твого.
DEUT|26|5|А ти відповіси та й скажеш перед лицем Господа, Бога свого: Мандрівний арамеянин був мій батько, і він зійшов до Єгипту, і часово замешкав там із небагатьма людьми, та й став там народом великим, сильним та численним.
DEUT|26|6|І чинили нам зло єгиптяни, і гнобили нас, і давали нас на роботу тяжку.
DEUT|26|7|І голосили ми до Господа, Бога батьків наших. І почув Господь голос наш, і побачив нашу біду, і труд наш, і утиск наш.
DEUT|26|8|І вивів нас Господь із Єгипту рукою сильною та раменом витягненим, і страхом великим, і ознаками та чудами.
DEUT|26|9|І привів нас до цього місця, і дав нам цей Край, Край, що тече молоком та медом.
DEUT|26|10|А тепер оце приніс я початок плоду тієї землі, яку Ти дав мені, Господи. І покладеш його перед лицем Господа, Бога свого, і поклонишся перед лицем Господа, Бога свого.
DEUT|26|11|І будеш радіти всім добром, що дав тобі Господь, Бог твій, тобі та домові твоєму, ти, і Левит, і приходько, що посеред тебе.
DEUT|26|12|А коли ти скінчиш десятинити всю десятину врожаю свого року третього, року десятини, і даси Левиту, приходькові, сироті та вдові, і будуть вони їсти в брамах твоїх і наситяться,
DEUT|26|13|то скажеш перед лицем Господа, Бога свого: Забрав я присвячене з дому, та й дав його Левиту та приходькові, сироті та вдові, за всіма Твоїми заповідями, що Ти наказав був мені, я не переступив котроїсь із заповідей Твоїх і не забув.
DEUT|26|14|Не їв я з нього в жалобі своїй, і не брав з нього в нечистості, і не дав з нього для померлого, я слухався голосу Господа, Бога свого, чинив усе, як наказав Ти мені.
DEUT|26|15|Споглянь же з святого мешкання Свого, із небес, і поблагослови народ Свій, Ізраїля, та землю, яку Ти дав нам, як присягнув був нашим батькам, Край, що тече молоком та медом.
DEUT|26|16|Цього дня Господь, Бог твій, наказує тобі виконувати ці постанови та закони, а ти будеш додержувати, та будеш виконувати їх усім серцем своїм та всією душею своєю.
DEUT|26|17|Ти сьогодні засвідчив Господеві, що Він буде тобі Богом, і що ти будеш ходити дорогами Його, і що будеш виконувати постанови Його, і заповіді Його, і закони Його, і що будеш слухатися голосу Його.
DEUT|26|18|А Господь сьогодні засвідчив тобі, що ти будеш Йому народом вибраним, як Він наказав був тобі, і що ти виконуватимеш усі заповіді Його,
DEUT|26|19|і що Він ставить тебе найвищим понад усі народи, яких Господь учинив, на хвалу, і на ім'я, і на славу, і що будеш ти для Господа, Бога свого, народом святим, як Він говорив вам.
DEUT|27|1|І наказав Мойсей та Ізраїлеві старші народові, говорячи: Додержуйте всіх заповідей, що я сьогодні наказую вам!
DEUT|27|2|І станеться того дня, коли ви перейдете Йордан до того Краю, що дає тобі Господь, Бог твій, то поставиш собі велике каміння, і повапниш їх вапном.
DEUT|27|3|І понаписуєш на них усі слова цього Закону, коли перейдеш, щоб увійшов ти до того Краю, що Господь, Бог твій, дає тобі, Край, що тече молоком та медом, як промовляв був Господь, Бог батьків твоїх, до тебе.
DEUT|27|4|І станеться, коли ви перейдете Йордан, поставите те каміння, що я наказую вам сьогодні, на горі Евал, і повапните їх вапном.
DEUT|27|5|І збудуєш там жертівника для Господа, Бога свого, жертівника з каміння, не піднесеш над ними заліза.
DEUT|27|6|З нетесаного каміння збудуєш жертівника Господа, Бога свого, і принесеш на ньому цілопалення Господеві, Богові своєму.
DEUT|27|7|І принесеш на жертву мирні жертви, і будеш там їсти, і будеш тішитися перед лицем Господа, Бога свого.
DEUT|27|8|І напишеш на тих каміннях усі слова цього Закону дуже виразно.
DEUT|27|9|І промовляв Мойсей та всі священики-Левити, до всього Ізраїля, говорячи: Уважай та слухай, Ізраїлю, ти цього дня став народом Господа, Бога свого.
DEUT|27|10|І будеш ти слухатися Господа, Бога свого, і будеш виконувати заповіді Його та постанови Його, що я наказую тобі сьогодні.
DEUT|27|11|І наказав Мойсей того дня народові, говорячи:
DEUT|27|12|Оці стануть на горі Ґарізім, щоб благословляти народ, коли ви перейдете Йордан: Симеон, і Левій, і Юда, і Іссахар, і Йосип, і Веніямин.
DEUT|27|13|А оці стануть для клятви на горі Евал: Рувим, Ґад, і Асир, і Завулон, Дан і Нефталим.
DEUT|27|14|І відповідять Левити, і скажуть до всіх Ізраїлевих мужів сильним голосом:
DEUT|27|15|Проклята людина, що зробить боввана різаного або литого, гидоту для Господа, чин різьбарських рук, і поставить таємно! І відповість увесь народ, та й скаже: амінь!
DEUT|27|16|Проклятий той, хто легковажить свого батька та свою матір! А ввесь народ скаже: амінь!
DEUT|27|17|Проклятий, хто пересуває межу свого ближнього!
DEUT|27|18|Проклятий, хто робить блудячим сліпого в дорозі! А ввесь народ скаже: амінь!
DEUT|27|19|Проклятий, хто перекручує право приходька, сироти та вдови! А ввесь народ скаже: амінь!
DEUT|27|20|Проклятий, хто лягає з жінкою батька свого, бо відкрив він подолка одежі свого батька! А ввесь народ скаже: амінь!
DEUT|27|21|Проклятий, хто лягає з усяким скотом! А ввесь народ скаже: амінь!
DEUT|27|22|Проклятий, хто лягає з сестрою своєю, дочкою свого батька або з дочкою своєї матері! А ввесь народ скаже: амінь!
DEUT|27|23|Проклятий, хто лягає з тещею своєю! А ввесь народ скаже: амінь!
DEUT|27|24|Проклятий, хто вбиває свого ближнього потаємно! А ввесь народ скаже: амінь!
DEUT|27|25|Проклятий, хто бере підкупа, щоб забити кого, пролляти кров неповинну! А ввесь народ скаже: амінь!
DEUT|27|26|Проклятий, хто не дотримає слів цього Закону, щоб виконувати їх! А ввесь народ скаже: амінь!
DEUT|28|1|І станеться, якщо дійсно будеш ти слухатися голосу Господа, Бога свого, щоб додержувати виконання всіх Його заповідей, що я наказую тобі сьогодні, то поставить тебе Господь, Бог твій, найвищим над усі народи землі.
DEUT|28|2|І прийдуть на тебе всі оці благословення, і досягнуть тебе, коли ти слухатимешся голосу Господа, Бога свого.
DEUT|28|3|Благословенний ти в місті, і благословенний ти на полі!
DEUT|28|4|Благословенний плід утроби твоєї, і плід твоєї землі, і плід худоби твоєї, порід биків твоїх і котіння отари твоєї!
DEUT|28|5|Благословенний твій кіш та діжа твоя!
DEUT|28|6|Благословенний ти у вході своїм, і благословенний ти в виході своїм!
DEUT|28|7|Господь учинить, що вороги твої, які повстають на тебе, будуть побиті перед тобою, вони однією дорогою вийдуть навперейми тебе, а сімома дорогами втікатимуть перед тобою.
DEUT|28|8|Господь накаже Своєму благословенню бути з тобою в коморах твоїх, та в усьому, чого доторкнеться рука твоя, і благословлятиме тебе в Краю, що Господь, Бог твій, дає тобі.
DEUT|28|9|Господь поставить тебе Собі за святий народ, як присягнув був тобі, коли ти будеш додержуватися заповідей Господа, Бога твого, і підеш дорогами Його.
DEUT|28|10|І побачать усі народи землі, що Господнє Ім'я кличеться на тобі, і будуть боятися тебе.
DEUT|28|11|І Господь дасть тобі добрий приріст у плоді утроби твоєї, і в плоді худоби твоєї, і в плоді поля твого на тій землі, що Господь заприсягнув був батькам твоїм, щоб дати тобі.
DEUT|28|12|Господь відчинить для тебе Свою добру скарбницю, небеса, щоб дати дощ для Краю твого в часі його, і щоб поблагословити всякий чин твоєї руки. І ти позичатимеш багатьом народам, а сам не позичатимеш ні в кого.
DEUT|28|13|І вчинить тебе Господь головою, а не хвостом, і ти будеш тільки верхом, а не будеш долом, коли будеш слухатися заповідей Господа, Бога свого, що я сьогодні наказую тобі, щоб додержувати й виконувати,
DEUT|28|14|і не відступиш від усіх тих слів, що я сьогодні наказую вам, ані праворуч, ані ліворуч, щоб ходити за іншими богами й служити їм.
DEUT|28|15|Та станеться, коли ти не будеш слухатися голосу Господа, Бога свого, щоб додержувати виконання всіх Його заповідей та постанов Його, що я сьогодні наказую тобі, то прийдуть на тебе всі оці прокляття, і досягнуть тебе:
DEUT|28|16|Проклятий ти в місті, і проклятий ти в полі!
DEUT|28|17|Проклятий кіш твій та діжа твоя!
DEUT|28|18|Проклятий плід утроби твоєї та плід твоєї землі, порід биків твоїх та котіння отари твоєї!
DEUT|28|19|Проклятий ти у вході своїм, і проклятий ти в виході своїм!
DEUT|28|20|Пошле Господь на тебе прокляття, і замішання, і нещастя на всякий почин твоєї руки, що ти зробиш, аж поки ти не будеш вигублений, і аж поки ти скоро не загинеш через зло твоїх чинів, що опустив ти Мене.
DEUT|28|21|Приліпить Господь до тебе моровицю, аж поки вона не вигубить тебе з-над землі, куди ти входиш посісти її.
DEUT|28|22|Ударить Господь тебе сухотами, і пропасницею, і запаленням, і гарячкою, і мечем, і посухою, і іржею, і вони будуть гнати тебе, аж поки ти не загинеш.
DEUT|28|23|І стане небо твоє, що над твоєю головою, міддю, а земля, що під тобою, залізом.
DEUT|28|24|Дасть Господь замість дощу Краєві твоєму куряву, а порох із неба буде сходити на тебе, аж поки не будеш ти вигублений.
DEUT|28|25|Віддасть тебе Господь на поразку твоїм ворогам. Однією дорогою ти вийдеш навперейми його, а сімома дорогами втікатимеш перед ним, і будеш розпорошений по всіх царствах землі.
DEUT|28|26|І буде твій труп на їжу для всякого птаства небесного та для худоби земної, і не буде нікого, хто б їх пополошив.
DEUT|28|27|Ударить тебе Господь єгипетським гнояком, ґудзами, лишаями, струпами такими, що не зможеш їх вилікувати.
DEUT|28|28|Ударить тебе Господь божевіллям, і сліпотою, і туподумством.
DEUT|28|29|І будеш ти мацати в південь, як мацає сліпий у темряві, і не матимеш поводження в дорогах своїх, і будеш ти по всі дні тільки утискуваний та грабований, та не буде кому боронити.
DEUT|28|30|Одружишся з жінкою, та хто інший лежатиме з нею. Хату збудуєш, та в ній не сидітимеш. Засадиш виноградника, та не будеш користатися ним.
DEUT|28|31|Заколений буде віл твій на очах твоїх, та їсти не будеш із нього. Твій осел буде заграбований перед тобою, і не вернеться до тебе. Отара твоя віддана буде ворогам твоїм, і не буде кому боронити тебе.
DEUT|28|32|Сини твої та дочки твої будуть віддані іншому народові, а очі твої будуть бачити й гинути за ними цілий день, а твоя рука не матиме сили.
DEUT|28|33|Плід твоєї землі та ввесь труд твій поїсть народ, якого ти не знав, а ти будеш тільки утискуваний та гноблений по всі дні.
DEUT|28|34|І ти збожеволієш від того, що бачитимуть очі твої.
DEUT|28|35|Ударить тебе Господь злим гнояком на колінах і на стегнах, від якого не зможеш вилікуватися, від стопи ніг твоїх і аж до черепа твого.
DEUT|28|36|Відведе Господь тебе та царя твого, якого поставиш над собою, до народу, якого не знав ти та батьки твої, і ти будеш служити там іншим богам, дереву та каменеві.
DEUT|28|37|І станеш ти страхіттям, поговором та посміховищем серед усіх народів, куди відведе тебе Господь.
DEUT|28|38|Багато насіння винесеш на поле, та мало збереш, бо пожере його сарана.
DEUT|28|39|Позасаджуєш виноградники й будеш обробляти, та не будеш пити вина й не будеш збирати, бо пожере його черва.
DEUT|28|40|Будуть у тебе оливки по всім краї твоїм, та оливою не будеш маститися, бо поспадає оливка твоя.
DEUT|28|41|Ти породиш синів і дочок, та не будуть для тебе вони, бо підуть у неволю.
DEUT|28|42|Усяке твоє дерево та плід твоєї землі обсяде черва.
DEUT|28|43|Приходько, що серед тебе, піднесеться понад тебе високо-високо, а ти зійдеш низько-низько.
DEUT|28|44|Він тобі позичатиме, а ти йому не позичатимеш, він стане головою, а ти станеш хвостом.
DEUT|28|45|І прийдуть на тебе всі оці прокляття, і будуть гнати тебе, і доженуть тебе, аж поки ти будеш вигублений, бо не слухав ти голосу Господа, Бога свого, щоб виконувати заповіді Його та постанови Його, що Він наказав був тобі.
DEUT|28|46|І будуть вони на тобі на ознаку та на доказ, та на насінні твоєму аж навіки.
DEUT|28|47|За те, що не служив ти Господеві, Богові своєму, у радості та в добрі серця, із рясноти всього,
DEUT|28|48|то будеш служити ворогові своєму, якого Господь пошле на тебе, у голоді, і в прагненні, і в наготі, і в недостатку всього, а він дасть залізне ярмо на твою шию, аж поки вигубить тебе.
DEUT|28|49|Господь нанесе на тебе народ іздалека, з кінця землі, так, як летить орел, народ, що мови його ти не розумієш,
DEUT|28|50|народ жорстокий, що не зважатиме на старого, а для юнака не буде милостивий.
DEUT|28|51|І він буде жерти плід твоєї худоби та плід твоєї землі, аж поки вигубить тебе, і він не позоставить тобі збіжжя, ані виноградного соку, ані оливи, ані породу биків твоїх, ані котіння отари твоєї, аж поки вигубить тебе.
DEUT|28|52|І він буде облягати тебе в усіх твоїх брамах, аж поки порозвалює по всім твоїм краї твої міцні і укріплені мури, на які ти надіявся, і буде гнобити тебе в усіх твоїх брамах по всім твоїм краї, що дав тобі Господь, Бог твій.
DEUT|28|53|І будеш ти їсти плід утроби своєї, тіло синів своїх та дочок своїх, що дав тобі Господь, Бог твій, в облозі та в утиску, яким буде гнобити тебе твій ворог.
DEUT|28|54|Кожен найлагідніший серед тебе й найбільше випещений, буде око його лихе на брата свого, і на жінку лоня свого, і на решту синів своїх, що позоставить їх ворог,
DEUT|28|55|щоб не дати ані одному з них тіла синів своїх, що буде він їсти, бо йому не позостанеться нічого в облозі та в утискові, яким буде утискати тебе твій ворог по всіх твоїх брамах.
DEUT|28|56|Найлагідніша між тобою й найбільше випещена, що через пещення та ніжність не пробувала ставити на землю стопи своєї ноги, зле буде око її на мужа лоня свого, і на сина свого, і на дочку свою,
DEUT|28|57|і на послід, що виходить з-поміж ніг її при породі, і на дітей своїх, що породить, бо поїсть їх таємно через недостаток усього в облозі та в утиску, яким буде гнобити тебе твій ворог у брамах твоїх.
DEUT|28|58|Якщо ти не будеш додержувати, щоб виконувати всі слова цього Закону, написані в цій книзі, щоб боятися того славного й страшного Ймення Господа, Бога твого,
DEUT|28|59|то Господь наведе надзвичайні порази на тебе, та порази на насіння твоє, порази великі та певні, і хвороби злі та постійні.
DEUT|28|60|І наведе Він на тебе всякий єгипетський біль, якого боявся ти, а він пристане до тебе.
DEUT|28|61|Також усяку хворобу та всяку поразу, що не написана в книзі цього Закону, наведе їх Господь на тебе, аж поки будеш ти вигублений.
DEUT|28|62|І позостане вас мало, замість того, що були ви, щодо численности, як зорі небесні, бо ти не слухався голосу Господа, Бога свого.
DEUT|28|63|І станеться, як Господь радів був вами, коли робив вам добро, і коли розмножував вас, так буде радіти Господь вами, коли вигублятиме вас та коли винищуватиме вас, і ви будете вирвані з-над цієї землі, куди ти входиш посісти її.
DEUT|28|64|І розпорошить тебе Господь серед усіх народів від кінця землі й аж до кінця землі, і ти служитимеш там іншим богам, яких не знав ані ти, ані батьки твої, дереву та каменеві.
DEUT|28|65|І поміж цими народами не будеш ти спокійний, і не буде місця спочинку для стопи твоїх ніг. І Господь дасть тобі там серце тремтяче, і ослаблення очей, і омлівання душі.
DEUT|28|66|І буде життя твоє висіти на волоску перед тобою і ти боятимешся вдень та вночі, і не будеш певний свого життя.
DEUT|28|67|Уранці ти скажеш: О, якби вечір!, а ввечері скажеш: О, якби ранок! зо страху серця свого, що будеш боятися, та з видіння очей своїх, що будеш бачити.
DEUT|28|68|І верне тебе Господь до Єгипту на кораблях тією дорогою, про яку я казав тобі, що вже більше не побачиш її, і там ви продаватиметеся ворогам своїм за рабів та за невільниць, та не буде покупця...
DEUT|29|1|(28-69) Оце слова заповіту, що наказав був Господь Мойсеєві скласти з Ізраїлевими синами в моавському краї, окрім того заповіту, що склав був із ними на Хориві.
DEUT|29|2|(29-1) І скликав Мойсей усього Ізраїля та й сказав їм: Ви бачили все, що зробив був Господь на ваших очах в єгипетськім краї фараонові, і всім рабам його та всьому його краєві,
DEUT|29|3|(29-2) ті великі випробування, що бачили очі твої, ті великі ознаки та чуда,
DEUT|29|4|(29-3) та не дав вам Господь серця, щоб пізнати, і очей, щоб бачити, і ушей, щоб слухати, аж до дня цього.
DEUT|29|5|(29-4) І провадив я вас сорок літ пустинею, не зужилися одежі ваші на вас, а чобіт твій не зужився на твоїй нозі.
DEUT|29|6|(29-5) Не їли ви хліба, і вина та п'янкого напою не пили ви, щоб пізнати, що Я Господь, Бог ваш.
DEUT|29|7|(29-6) А коли ви прийшли до цього місця, то вийшов був навперейми вас на війну Сигон, цар хешбонський, та Оґ, цар башанський, і побили ми їх,
DEUT|29|8|(29-7) і забрали ми їхній край, та й дали його на спадок Рувимовим та Ґадовим та половині племени Манасіїного.
DEUT|29|9|(29-8) Додержуй же слів цього заповіту, і виконуй їх, щоб мали ви поводження в усьому, що будете робити.
DEUT|29|10|(29-9) Ви стоїте сьогодні всі перед лицем Господа, Бога вашого: голови ваші, племена ваші, старші ваші та урядники ваші, усякий Ізраїлів муж,
DEUT|29|11|(29-10) діти ваші, ваші жінки та твій приходько, що посеред таборів твоїх від колія дров твоїх аж до черпача твоєї води,
DEUT|29|12|(29-11) щоб ти ввійшов у заповіт Господа, Бога свого, та в клятву Його, що Господь, Бог твій, сьогодні складає з тобою,
DEUT|29|13|(29-12) щоб поставити сьогодні тебе народом для Себе, а Він буде тобі Богом, як Він говорив був тобі, і як присягнув був батькам твоїм, Авраамові, Ісакові та Якову.
DEUT|29|14|(29-13) І не з вами самими я складаю цього заповіта та цю клятву,
DEUT|29|15|(29-14) але теж і з тим, хто тут з нами сьогодні стоїть перед лицем Господа, Бога нашого, так і з тим, хто сьогодні не з нами тут.
DEUT|29|16|(29-15) Бо ви знаєте, що ми сиділи були в єгипетськім краї, і що ми проходили серед тих народів, які ви перейшли,
DEUT|29|17|(29-16) І ви бачили їхні огиди та їхніх бовванів, дерево та камінь, срібло та золото, що з ними.
DEUT|29|18|(29-17) Стережіться, щоб не був серед вас чоловік або жінка, або рід, або плем'я, що серце його сьогодні відвертається від Господа, Бога нашого, щоб піти служити богам цих народів, щоб не був серед вас корінь, що вирощує їдь та полин,
DEUT|29|19|(29-18) щоб не було, що коли він почує слова цього прокляття, то поблагословиться в серці своїм, говорячи: Мир буде мені, хоч і ходитиму в сваволі свого серця. Тоді загине і напоєний, і спрагнений.
DEUT|29|20|(29-19) Не захоче Господь простити йому, бо тоді запалиться Господній гнів та лютість Його на цього чоловіка, і буде лежати на ньому все прокляття, написане в цій книзі, і Господь витре ім'я його з-під неба.
DEUT|29|21|(29-20) І відділить його Господь на зло від усіх Ізраїлевих племен, згідно з усіма прокляттями заповіту, написаного в цій книзі Закону.
DEUT|29|22|(29-21) І скаже останнє покоління, ваші сини, що постануть за вами, і чужий, що прийде з далекої країни, і побачить порази цього Краю та його хвороби, які пошле Господь на нього:
DEUT|29|23|(29-22) сірка та сіль, погорілище уся земля його, не буде вона засіювана, і не пустить рослин, і не зійде на ній жодна трава, як по знищенні Содому та Гомори, Адми та Цевоїму, що поруйнував був Господь у гніві Своїм та в люті Своїй.
DEUT|29|24|(29-23) І скажуть усі ті народи: Для чого Господь зробив так цьому Краєві? Що то за горіння цього великого гніву?
DEUT|29|25|(29-24) І скажуть: За те, що вони покинули заповіта Господа, Бога своїх батьків, якого Він склав був із ними, коли виводив їх з єгипетського краю.
DEUT|29|26|(29-25) І вони пішли, і служили іншим богам, і вклонялися їм, богам, що не знали їх, і що Він не приділив їм.
DEUT|29|27|(29-26) І запалився Господній гнів на цей Край, щоб навести на нього все прокляття, написане в цій книзі.
DEUT|29|28|(29-27) І вирвав їх Господь з-над цієї землі в гніві, і в люті, і в великім обуренні, та й кинув їх до іншого краю, як цього дня.
DEUT|29|29|(29-28) Закрите те, що є Господа, Бога нашого, а відкрите наше та наших синів аж навіки, щоб виконувати всі слова цього Закону.
DEUT|30|1|І станеться, коли прийдуть на тебе всі ці слова, благословення та прокляття, що я дав перед тобою, і ти візьмеш їх до свого серця серед усіх цих народів, куди закинув тебе Господь, Бог твій,
DEUT|30|2|і ти навернешся до Господа, Бога свого, і будеш слухатися Його голосу в усьому, що я сьогодні тобі наказую, ти та сини твої, усім своїм серцем та всією своєю душею,
DEUT|30|3|то поверне з неволі Господь, Бог твій, тебе, і змилосердиться над тобою, і знову позбирає тебе зо всіх народів, куди розпорошив тебе Господь, Бог твій.
DEUT|30|4|Якщо буде твій вигнанець на кінці неба, то й звідти позбирає тебе Господь, Бог твій, і звідти Він візьме тебе.
DEUT|30|5|І введе тебе Господь, Бог твій, до Краю, що посіли батьки твої, і ти посядеш його, і Він учинить добро тобі, і розмножить тебе більше за батьків твоїх.
DEUT|30|6|І обріже Господь, Бог твій, серце твоє та серце насіння твого, щоб ти любив Господа, Бога свого, усім своїм серцем та всією душею своєю, щоб жити тобі.
DEUT|30|7|І дасть Господь, Бог твій, усі ці прокляття на ворогів твоїх, та на тих, хто ненавидить тебе, хто гнав тебе.
DEUT|30|8|А ти вернешся, і будеш слухатися Господнього голосу, і будеш виконувати всі Його заповіді, які я сьогодні наказую тобі.
DEUT|30|9|І зробить Господь, Бог твій, що будеш ти мати надмір у кожному чині своєї руки, у плоді утроби своєї, і в плоді худоби своєї, і в плоді своєї землі на добре, бо Господь знову буде радіти тобою на добро, як радів був твоїми батьками,
DEUT|30|10|коли будеш слухатися голосу Господа, Бога свого, щоб дотримувати заповіді Його та постанови Його, написані в цій книзі Закону, коли навернешся до Господа, Бога свого, усім серцем своїм та всією душею своєю,
DEUT|30|11|бо ця заповідь, що я сьогодні наказую тобі, не тяжка вона для тебе, і не далека вона.
DEUT|30|12|Не на небі вона, щоб сказати: Хто зійде на небо для нас, та нам її візьме і нам оголосить, а ми будемо виконувати її?
DEUT|30|13|І не по тім боці моря вона, щоб сказати: Хто піде для нас на той бік моря, і візьме її нам, і оголосить її нам, а ми будемо виконувати її?
DEUT|30|14|Бож дуже близька до тебе та річ, вона в устах твоїх та в серці твоїм, щоб виконувати її.
DEUT|30|15|Дивися: я сьогодні дав перед тобою життя та добро, і смерть та зло.
DEUT|30|16|Бо я сьогодні наказую тобі любити Господа, Бога свого, ходити Його дорогами, та додержувати заповіді Його, і постанови Його, і закона Його, щоб ти жив, і розмножився, і поблагословить тебе Господь, Бог твій, у Краї, куди ти входиш на насліддя.
DEUT|30|17|А якщо серце твоє відвернеться, і не будеш ти слухатися, і даси себе звести, і станеш вклонятися іншим богам, і будеш їм служити,
DEUT|30|18|я сьогодні представив вам, що конче погинете ви, недовго житимете на цій землі, до якої ти переходиш Йордан, щоб увійти туди на оволодіння її.
DEUT|30|19|Сьогодні взяв я за свідків проти вас небо й землю, життя та смерть дав я перед вами, благословення та прокляття. І ти вибери життя, щоб жив ти та насіння твоє,
DEUT|30|20|щоб любити Господа, Бога свого, щоб слухатися голосу Його та щоб линути до Нього, бож Він життя твоє, і довгота днів твоїх, щоб сидіти на цій землі, яку заприсягнув Господь батькам твоїм Авраамові, Ісакові та Якову, дати їм.
DEUT|31|1|І пішов Мойсей, і промовляв до всього Ізраїля оці слова,
DEUT|31|2|та й сказав їм: Я сьогодні віку ста й двадцяти літ. Не можу вже виходити та входити, і Господь сказав мені: Не перейдеш ти цього Йордану.
DEUT|31|3|Господь, Бог твій, Він піде перед тобою, Він вигубить ці народи перед тобою, і ти заволодієш ними. Ісус перейде перед тобою, як говорив був Господь.
DEUT|31|4|І зробить їм Господь, як зробив був Сигонові та Оґові, аморейським царям та їхньому краєві, яких вигубив Він.
DEUT|31|5|І дасть їх Господь перед вас, а ви зробите їм згідно з усією заповіддю, що я вам наказав був.
DEUT|31|6|Будьте сильні та відважні, не бійтеся, не лякайтеся перед ними, бо Господь, Бог твій, Він Той хто ходить з тобою, не опустить Він тебе й не покине тебе.
DEUT|31|7|І покликав Мойсей Ісуса, та й до нього сказав на очах усього Ізраїля: Будь сильний та відважний, бо ти ввійдеш з цим народом до того Краю, якого Господь заприсягнув їхнім батькам, щоб їм дати, і ти даси їм його на спадок.
DEUT|31|8|А Господь, Він Той, що піде перед тобою, не опустить тебе й не покине тебе, не бійся й не лякайся.
DEUT|31|9|І написав Мойсей цього Закона, та й дав його до священиків, Левієвих синів, що носять ковчега Господнього заповіту, та до всіх Ізраїлевих старших.
DEUT|31|10|І наказав їм Мойсей, говорячи: У кінці семи літ, окресленого часу року відпущення, у свято Кучок,
DEUT|31|11|коли прийде ввесь Ізраїль з'явитися перед лицем Господа, Бога свого, у місці, яке вибере Він, будеш читати цього Закона перед усім Ізраїлем до їхніх ушей.
DEUT|31|12|Збери той народ, чоловіків, і жінок, і дітей, і приходька свого, що в твоїх брамах, щоб вони чули й щоб навчалися, і боялися Господа, Бога вашого, і додержували виконувати всі слова цього Закону.
DEUT|31|13|А їхні сини, що не знали, будуть чути та навчатися боятися Господа, Бога вашого, по всі дні, що ви житимете на цій землі, куди ви переходите Йордан, щоб посісти її.
DEUT|31|14|І сказав Господь до Мойсея: Оце наблизилися дні твої до смерти. Поклич Ісуса, і станьте в скинії заповіту, а Я йому накажу. І пішов Мойсей та Ісус, і стали в скинії заповіту.
DEUT|31|15|І появився Господь у скинії в стовпі хмари, і став той стовп хмари біля скинійного входу.
DEUT|31|16|І сказав Господь до Мойсея: Ось ти спочинеш з батьками своїми, а цей народ устане та й буде блудодіяти з богами того чужого Краю, куди він увіходить, щоб бути в середині його, і покине Мене, і зламає заповіта Мого, що склав був Я з ним.
DEUT|31|17|І того дня запалиться Мій гнів на нього, і Я покину їх, і сховаю Своє лице від них, а він буде знищений, і знайдуть його численні нещастя та утиски. І скаже він того дня: Хіба не через те, що нема в мене мого Бога, знайшли мене ці нещастя?
DEUT|31|18|А Я того дня конче сховаю лице Своє через усе те зло, що зробив він, бо звернувся до інших богів.
DEUT|31|19|А тепер запишіть собі оцю пісню, і навчи її Ізраїлевих синів. Вклади її в їхні уста, щоб була мені ця пісня за свідка на Ізраїлевих синів.
DEUT|31|20|Коли Я введу його до тієї землі, яку присягнув його батькам, що тече молоком та медом, і він буде їсти й насититься, і потовстіє, і звернеться до інших богів, і будуть служити їм, а Мене кинуть з образою, і зламає він заповіта Мого,
DEUT|31|21|то станеться, коли знайдуть його численні нещастя та утиски, що пісня ця стане проти нього за свідка, бо вона не забудеться з уст насіння його. Бо Я знаю наставлення серця його, що він чинить сьогодні, перше ніж введу його до того Краю, що Я присягнув.
DEUT|31|22|І написав Мойсей ту пісню того дня, і навчив її Ізраїлевих синів.
DEUT|31|23|І наказав він Ісусові, Навиновому синові, та й сказав: Будь сильний та відважний, бо ти впровадиш Ізраїлевих синів до того Краю, що Я присягнув їм, а Я буду з тобою.
DEUT|31|24|І сталося, як Мойсей скінчив писати слова цього Закону до книги аж до кінця їх,
DEUT|31|25|то Мойсей наказав Левитам, що носять ковчега Господнього заповіту, говорячи:
DEUT|31|26|Візьміть книгу цього Закону, і покладіть її збоку ковчега заповіту Господа, Бога вашого, і вона буде там на тебе за свідка.
DEUT|31|27|Бо я знаю неслухняність твою та тверду твою шию. Бо ще сьогодні, коли я живу з вами, ви були неслухняні Господеві, а тим більш будете по смерті моїй!
DEUT|31|28|Зберіть до мене всіх старших ваших племен та урядників ваших, а я буду промовляти до їхніх ушей ці слова, і покличу небо й землю на свідчення проти них.
DEUT|31|29|Бо я знаю, що по смерті моїй, псуючися, зіпсуєтеся ви, і відхилитесь з тієї дороги, яку я наказав вам, і в кінці днів спіткає вас нещастя, коли будете робити зло в Господніх очах, щоб гнівити Його чином своїх рук.
DEUT|31|30|І промовляв Мойсей до ушей всієї Ізраїлевої громади слова оцієї пісні аж до закінчення їх:
DEUT|32|1|Слухай, небо, а я говоритиму, і хай почує земля мову уст моїх!
DEUT|32|2|Нехай ллється наука моя, мов той дощ, хай тече, як роса, моя мова, як краплі дощу на траву, та як злива на зелень.
DEUT|32|3|Як буду я кликати Ймення Господнє, то славу віддайте ви нашому Богові!
DEUT|32|4|Він Скеля, а діло Його досконале, всі бо дороги Його справедливі, Бог вірний, і кривди немає в Ньому, справедливий і праведний Він.
DEUT|32|5|Зіпсулись вони, не Його то сини, покоління невірне й покручене.
DEUT|32|6|Чи тим віддасте Господеві, народе нікчемний й немудрий? Чи ж не Він Батько твій, твій Творець? Він тебе вчинив, і Він міцно поставив тебе.
DEUT|32|7|Пам'ятай про дні давні, розважайте про роки усіх поколінь, запитай свого батька, і покаже тобі твоїх тих старших, а вони тобі скажуть.
DEUT|32|8|Як Всевишній народам спадок давав, коли Він розділяв синів людських, Він поставив границі народам за числом Ізраїлевих синів.
DEUT|32|9|Бо частка Господня народ Його, Яків відміряний уділ спадщини Його.
DEUT|32|10|Знайшов Він його на пустинній землі та в степу завивання пустельних гієн, та й його оточив, уважав Він за ним, зберігав Він його, як зіницю оту свого ока.
DEUT|32|11|Як гніздо своє будить орел, як ширяє він понад своїми малятами, крила свої простягає, бере їх, та носить їх він на рамені крилатім своїм,
DEUT|32|12|так Господь Сам провадив його, а бога чужого при нім не було.
DEUT|32|13|Він його садовив на висотах землі, і він їв польові врожаї, Він медом із скелі його годував, і оливою з скельного кременя,
DEUT|32|14|маслом з худоби великої та молоком від худоби дрібної, разом із лоєм ягнят та баранів з Башану й козлів, разом з такою пшеницею, як лій на нирках, і кров виноградної ягоди пив ти вином.
DEUT|32|15|І потовстів Єшурун та й брикатися став. І ти потовстів, погрубів, став гладкий. І покинув він Бога, що його створив, і Скелю спасіння свого злегковажив.
DEUT|32|16|Чужими богами Його роздражнили, Його розгнівили своїми гидотами.
DEUT|32|17|Вони демонам жертви складали, не Богу, складали богам, що не відали їх, новим, що недавно прийшли, не лякалися їх батьки ваші!
DEUT|32|18|Забуваєш ти Скелю, Яка породила тебе, і забуваєш ти Бога, що тебе народив.
DEUT|32|19|І побачив Господь, та й зненавидів їх, через гнів на синів Своїх і на дочок Своїх,
DEUT|32|20|та й сказав: Лице Я Своє заховаю від них, побачу, який їх кінець, бо вони покоління розбещене, діти, що в них нема віри.
DEUT|32|21|Роздражнили Мене вони тим, хто не Бог, Мене розгнівили своїми марнотами, тому роздражню Я їх тим, хто не народ, нерозумним народом розгніваю їх.
DEUT|32|22|Бо був загорівся огонь Мого гніву, і палився він аж до шеолу найглибшого, і він землю поїв та її врожай, і спалив був підвалини гір.
DEUT|32|23|Я на них нагромаджу нещастя, зуживу Свої стріли на них.
DEUT|32|24|Будуть виснажені вони голодом, і поїджені будуть огнем та заразою лютою, і зуба звірини нашлю Я на них, з отрутою плазунів по землі.
DEUT|32|25|Надворі забиватиме меч, а в кімнатах страхіття, як юнака, так і дівчину, грудне немовля з чоловіком посивілим.
DEUT|32|26|Я сказав: Повигублюю їх, відірву від людей їхню пам'ять,
DEUT|32|27|та це Я відклав з-за ворожого гніву, щоб противники їх не згордилися, щоб вони не сказали: Піднеслася наша рука, і не Господь учинив усе це.
DEUT|32|28|Бо вони люд безрадний, і нема в них розумування.
DEUT|32|29|Коли б були мудрі вони, зрозуміли б оце, розсудили б були про кінець свій.
DEUT|32|30|Як може один гнати тисячу, а два проганять десять тисяч, коли то не те, що їх продала їхня Скеля, і Господь видав їх?
DEUT|32|31|Не така бо їх скеля, як наша та Скеля, хай судять самі вороги.
DEUT|32|32|Бо їх виноград з винограду содомського та з піль тих гоморських, винні ягоди їхні отруйні то ягоди, вони грона гіркоти для них,
DEUT|32|33|вино їхнє зміїна отрута і гадюча погибельна їдь!
DEUT|32|34|Чи замкнене в Мене не це, у скарбницях Моїх запечатане?
DEUT|32|35|Моя пімста й відплата на час, коли їхня нога посковзнеться, бо близький день погибелі їх, поспішає майбутнє для них.
DEUT|32|36|Бо розсудить Господь Свій народ, і змилосердиться Він над Своїми рабами, як побачить, що їхня рука ослабіла, і нема ні невільного, ані вільного.
DEUT|32|37|І Він скаже тоді: Де їх боги, де скеля, що в ній поховались вони,
DEUT|32|38|що їли вони лій кривавих їх жертов, пили вино жертов їх литих? Нехай встануть і вам допоможуть, і хай будуть покровом для вас.
DEUT|32|39|Побачте тепер, що Я Я є Той, і Бога немає крім Мене. Побиваю й оживлюю Я, і не врятує ніхто від Моєї руки.
DEUT|32|40|Бо до неба підношу Я руку Свою та й кажу: Я навіки Живий!
DEUT|32|41|Поправді кажу вам: Я вістря Свого меча нагострю, і рука Моя схопиться суду, тоді відімщу Я Своїм ворогам, і Своїм ненависникам Я відплачу.
DEUT|32|42|Я стріли Свої понапоюю кров'ю, а Мій меч поїдатиме м'ясо, кров'ю забитого й бранця, головами кучматими ворога.
DEUT|32|43|Радійте, погани, з народом Його, бо Він відімститься за кров Своїх всіх рабів, і пімсту поверне Своїм ворогам, і викупить землю Свою, Свій народ.
DEUT|32|44|І прийшов Мойсей, і промовляв всі слова цієї пісні до ушей народу, він та Ісус, син Навинів.
DEUT|32|45|А коли Мойсей скінчив промовляти всі ці слова до всього Ізраїля,
DEUT|32|46|то сказав він до них: Приложіть свої серця до всіх тих слів, які я сьогодні чинив свідками проти вас, що ви накажете їх своїм синам, щоб додержували виконувати всі слова цього Закону.
DEUT|32|47|Бо це для вас не слово порожнє, воно життя ваше, і цим словом ви продовжите дні на цій землі, куди ви переходите Йордан, щоб посісти її.
DEUT|32|48|І Господь промовляв до Мойсея того самого дня, говорячи:
DEUT|32|49|Вийди на ту гору Аварім, на гору Нево, що в моавському краї, що навпроти Єрихону, і побач ханаанський Край, що Я даю Ізраїлевим синам на володіння.
DEUT|32|50|І вмри на горі, куди ти вийдеш, і долучися до своєї рідні, як помер був твій брат Аарон на Гор-горі, і долучився до своєї рідні,
DEUT|32|51|за те, що ви спроневірилися були Мені серед Ізраїлевих синів при воді Меріви в Кадешу на пустині Цін, за те, що ви не освятили Мене серед Ізраїлевих синів.
DEUT|32|52|Бо знавпроти побачиш ти той Край, та не ввійдеш туди, до того Краю, що Я даю Ізраїлевим синам.
DEUT|33|1|А оце благословення, яким поблагословив Ізраїлевих синів Мойсей, чоловік Божий, перед своєю смертю,
DEUT|33|2|та й сказав: Господь від Сінаю прибув, і зійшов від Сеїру до них, появився у світлі з Парану гори, і прийшов із Меріви Кадешу. По правиці Його огонь Закону для них.
DEUT|33|3|Теж народи Він любить. Всі святії його у руці Твоїй, і вони припадають до ніг Твоїх, слухають мови Твоєї.
DEUT|33|4|Дав Мойсей нам Закона, спадщину зборові Якова.
DEUT|33|5|І був Він царем в Єшуруні, як народнії голови разом збирались, племена Ізраїлеві.
DEUT|33|6|Рувим хай живе, і нехай не помре, і число люду його нехай буде велике.
DEUT|33|7|А це про Юду. І він сказав: Почуй, Господи, голосу Юди, і до народу його Ти впровадиш його. Йому воюватимуть руки його, а Ти будеш поміч йому на його ворогів.
DEUT|33|8|А про Левія сказав: Твій туммім і твій урім для чоловіка святого Твого, що його Ти був випробував у Массі, що суперечку з ним мав над водою Меріви,
DEUT|33|9|що каже про батька свого та про матір свою: Не бачив тебе, що братів своїх не пізнає, і не знає синів своїх, бо додержують слова Твого, і вони заповіту Твого стережуть.
DEUT|33|10|Навчають вони про права Твої Якова, а про Закона Твойого Ізраїля, приносять кадило Тобі та на жертівник Твій цілопалення.
DEUT|33|11|Поблагослови його силу, о Господи, а чин його рук уподобай Собі. Поламай стегна тим, що стають проти нього, та ненависть мають на нього, щоб більш не повстали вони!
DEUT|33|12|Про Веніямина сказав: Він Господній улюбленець, перебуває безпечно при Ньому, а Він окриває його цілий день і в раменах Його спочиває.
DEUT|33|13|А про Йосипа він сказав: Благословенний від Господа Край Його дарами з неба, з роси та з безодні, що долі лежить,
DEUT|33|14|і з дару врожаїв від сонця, і з дару рослини від місяців,
DEUT|33|15|і з верхів'я гір сходу, і з дару відвічних пагірків,
DEUT|33|16|і з дару землі та її повноти. А милість Того, що в терновім кущі пробував, нехай прийде на голову Йосипа та на тім'я вирізненого між братами своїми.
DEUT|33|17|Величність його як вола його перворідного, а роги його роги буйвола, ними буде колоти народи всі разом, аж до кінців землі, а вони міріяди Єфремові, а вони Манасіїні тисячі.
DEUT|33|18|А про Завулона сказав: Радій, Завулоне, як будеш виходити, і ти, Іссахаре, у наметах своїх!
DEUT|33|19|Вони кличуть народи на гори, приносять там праведні жертви, бо будуть вони споживати достаток морський та скарби, зариті в піску.
DEUT|33|20|А про Ґада сказав: Благословенний, хто Ґада розширює! Він ліг, як левиця, і жере рам'я й череп.
DEUT|33|21|Забезпечив він частку для себе, бо там частка прихована від Праводавця, і прийшов із головами народу, виконав правду Господню і Його постанови з Ізраїлем.
DEUT|33|22|А на Дана сказав: Дан левів левчук, що з Башану вискакує.
DEUT|33|23|А на Нефталима сказав: Нефталим ситий милістю, і повен Господнього благословення, захід та південь посядь!
DEUT|33|24|А про Асира сказав: Асир благословенний найбільше з синів, уподобаний серед братів своїх, і в оливу вмочає він ногу свою.
DEUT|33|25|Залізо та мідь то запора твоя, а сила твоя як усі твої дні.
DEUT|33|26|Немає такого, як Бог, Єшуруне, що їде по небу на поміч тобі, а Своєю величністю їде на хмарах.
DEUT|33|27|Покрова твоя Бог Предвічний і ти в вічних раменах Його. І вигнав Він ворога перед тобою, і сказав: Повинищуй його!
DEUT|33|28|І перебуває Ізраїль безпечно, самотно, він Яковове джерело в Краї збіжжя й вина, а небо його сипле краплями росу.
DEUT|33|29|Ти блаженний, Ізраїлю! Який інший народ, якого спасає Господь, як тебе? Він Щит допомоги твоєї, і Меч Він твоєї величности. І будуть твої вороги при тобі упокорюватись, а ти по висотах їх будеш ступати.
DEUT|34|1|І вийшов Мойсей із моавських степів на гору Нево, на верхів'я Пісґі, що навпроти Єрихону, а Господь дав йому побачити ввесь Край: Ґілеад аж до Дану,
DEUT|34|2|і ввесь Нефталим, і край Єфрема та Манасії, і ввесь край Юди аж до Останнього моря,
DEUT|34|3|і південь, і рівнину долини Єрихону, пальмового міста аж до Цоару.
DEUT|34|4|І сказав Господь до нього: Оце той Край, що Я присягнув Авраамові, Ісакові та Якову, говорячи: Насінню твоєму Я дам його. Я вчинив, що ти бачиш його власними очима, та туди не перейдеш.
DEUT|34|5|І впокоївся там Мойсей, Господній раб, у моавському краї на приказ Господа.
DEUT|34|6|І похований він у долині в моавському краї навпроти Бет-Пеору, і ніхто не знає гробу його аж до цього дня.
DEUT|34|7|А Мойсей був віку ста й двадцяти літ, коли він помер, та не затемнилось око його, і вологість його не зменшилась.
DEUT|34|8|І оплакували Мойсея Ізраїлеві сини в моавських степах тридцять день, та й покінчилися дні оплакування жалоби за Мойсеєм.
DEUT|34|9|А Ісус, син Навинів, був повний духа мудрости, бо Мойсей поклав свої руки на нього. І слухали його Ізраїлеві сини, і робили, як Господь наказав був Мойсеєві.
DEUT|34|10|І не появився вже в Ізраїлі пророк, як Мойсей, що знав його Господь обличчя-в-обличчя,
DEUT|34|11|щодо всіх ознак та чуд, що Господь послав його чинити в єгипетськім краї фараонові й усім рабам його та всьому його краєві,
DEUT|34|12|і щодо всієї тієї сильної руки, і щодо всього того страху великого, що Мойсей чинив на очах усього Ізраїля.
