LEV|1|1|И воззвал Господь к Моисею и сказал ему из скинии собрания, говоря:
LEV|1|2|объяви сынам Израилевым и скажи им: когда кто из вас хочет принести жертву Господу, то, если из скота, приносите жертву вашу из скота крупного и мелкого.
LEV|1|3|Если жертва его есть всесожжение из крупного скота, пусть принесет ее мужеского пола, без порока; пусть приведет ее к дверям скинии собрания, чтобы приобрести ему благоволение пред Господом;
LEV|1|4|и возложит руку свою на голову [жертвы] всесожжения – и приобретет он благоволение, во очищение грехов его;
LEV|1|5|и заколет тельца пред Господом; сыны же Аароновы, священники, принесут кровь и покропят кровью со всех сторон на жертвенник, который у входа скинии собрания;
LEV|1|6|и снимет кожу с [жертвы] всесожжения и рассечет ее на части;
LEV|1|7|сыны же Аароновы, священники, положат на жертвенник огонь и на огне разложат дрова;
LEV|1|8|и разложат сыны Аароновы, священники, части, голову и тук на дровах, которые на огне, на жертвеннике;
LEV|1|9|а внутренности [жертвы] и ноги ее вымоет он водою, и сожжет священник все на жертвеннике: [это] всесожжение, жертва, благоухание, приятное Господу.
LEV|1|10|Если жертва всесожжения его из мелкого скота, из овец, или из коз, пусть принесет ее мужеского пола, без порока.
LEV|1|11|и заколет ее пред Господом на северной стороне жертвенника, и сыны Аароновы, священники, покропят кровью ее на жертвенник со всех сторон;
LEV|1|12|и рассекут ее на части, [отделив] голову ее и тук ее, и разложит их священник на дровах, которые на огне, на жертвеннике,
LEV|1|13|а внутренности и ноги вымоет водою, и принесет священник все и сожжет на жертвеннике: [это] всесожжение, жертва, благоухание, приятное Господу.
LEV|1|14|Если же из птиц приносит он Господу всесожжение, пусть принесет жертву свою из горлиц, или из молодых голубей;
LEV|1|15|священник принесет ее к жертвеннику, и свернет ей голову, и сожжет на жертвеннике, а кровь выцедит к стене жертвенника;
LEV|1|16|зоб ее с перьями ее отнимет и бросит его подле жертвенника на восточную сторону, где пепел;
LEV|1|17|и надломит ее в крыльях ее, не отделяя их, и сожжет ее священник на жертвеннике, на дровах, которые на огне: это всесожжение, жертва, благоухание, приятное Господу.
LEV|2|1|Если какая душа хочет принести Господу жертву приношения хлебного, пусть принесет пшеничной муки, и вольет на нее елея, и положит на нее ливана,
LEV|2|2|и принесет ее к сынам Аароновым, священникам, и возьмет полную горсть муки с елеем и со всем ливаном, и сожжет сие священник в память на жертвеннике; [это] жертва, благоухание, приятное Господу;
LEV|2|3|а остатки от приношения хлебного Аарону и сынам его: [это] великая святыня из жертв Господних.
LEV|2|4|Если же приносишь жертву приношения хлебного из печеного в печи, [то приноси] пшеничные хлебы пресные, смешанные с елеем, и лепешки пресные, помазанные елеем.
LEV|2|5|Если жертва твоя приношение хлебное со сковороды, то это должна быть пшеничная мука, смешанная с елеем, пресная;
LEV|2|6|разломи ее на куски и влей на нее елея: это приношение хлебное.
LEV|2|7|Если жертва твоя приношение хлебное из горшка, то должно сделать оное из пшеничной муки с елеем,
LEV|2|8|и принеси приношение, которое из сего составлено, Господу; представь оное священнику, а он принесет его к жертвеннику;
LEV|2|9|и возьмет священник из сей жертвы часть в память и сожжет на жертвеннике: [это] жертва, благоухание, приятное Господу;
LEV|2|10|а остатки приношения хлебного Аарону и сынам его: [это] великая святыня из жертв Господних.
LEV|2|11|Никакого приношения хлебного, которое приносите Господу, не делайте квасного, ибо ни квасного, ни меду не должны вы сожигать в жертву Господу;
LEV|2|12|как приношение начатков приносите их Господу, а на жертвенник не должно возносить их в приятное благоухание.
LEV|2|13|Всякое приношение твое хлебное соли солью, и не оставляй жертвы твоей без соли завета Бога твоего: при всяком приношении твоем приноси соль.
LEV|2|14|Если приносишь Господу приношение хлебное из первых плодов, приноси в дар от первых плодов твоих из колосьев, высушенных на огне, растолченные зерна,
LEV|2|15|и влей на них елея, и положи на них ливана: это приношение хлебное;
LEV|2|16|и сожжет священник в память часть зерен и елея со всем ливаном: [это] жертва Господу.
LEV|3|1|Если жертва его жертва мирная, и если он приносит из крупного скота, мужеского или женского пола, пусть принесет ее Господу, не имеющую порока,
LEV|3|2|и возложит руку свою на голову жертвы своей, и заколет ее у дверей скинии собрания; сыны же Аароновы, священники, покропят кровью на жертвенник со всех сторон;
LEV|3|3|и принесет он из мирной жертвы в жертву Господу тук, покрывающий внутренности, и весь тук, который на внутренностях,
LEV|3|4|и обе почки и тук, который на них, который на стегнах, и сальник, который на печени; с почками он отделит это;
LEV|3|5|и сыны Аароновы сожгут это на жертвеннике вместе со всесожжением, которое на дровах, на огне: [это] жертва, благоухание, приятное Господу.
LEV|3|6|А если из мелкого скота приносит он мирную жертву Господу, мужеского или женского пола, пусть принесет ее, не имеющую порока.
LEV|3|7|Если из овец приносит он жертву свою, пусть представит ее пред Господа,
LEV|3|8|и возложит руку свою на голову жертвы своей, и заколет ее пред скиниею собрания, и сыны Аароновы покропят кровью ее на жертвенник со всех сторон;
LEV|3|9|и пусть принесет из мирной жертвы в жертву Господу тук ее, весь курдюк, отрезав его по самую хребтовую кость, и тук, покрывающий внутренности, и весь тук, который на внутренностях,
LEV|3|10|и обе почки и тук, который на них, который на стегнах, и сальник, который на печени; с почками он отделит это;
LEV|3|11|священник сожжет это на жертвеннике; [это] пища огня – жертва Господу.
LEV|3|12|А если он приносит жертву из коз, пусть представит ее пред Господа,
LEV|3|13|и возложит руку свою на голову ее, и заколет ее перед скиниею собрания, и покропят сыны Аароновы кровью ее на жертвенник со всех сторон;
LEV|3|14|и принесет из нее в приношение, в жертву Господу тук, покрывающий внутренности, и весь тук, который на внутренностях,
LEV|3|15|и обе почки и тук, который на них, который на стегнах, и сальник, который на печени; с почками он отделит это
LEV|3|16|и сожжет их священник на жертвеннике: [это] пища огня – приятное благоухание [Господу]; весь тук Господу.
LEV|3|17|Это постановление вечное в роды ваши, во всех жилищах ваших; никакого тука и никакой крови не ешьте.
LEV|4|1|И сказал Господь Моисею, говоря:
LEV|4|2|скажи сынам Израилевым: если какая душа согрешит по ошибке против каких–либо заповедей Господних и сделает что–нибудь, чего не должно делать;
LEV|4|3|если священник помазанный согрешит и сделает виновным народ, – то за грех свой, которым согрешил, пусть представит из крупного скота тельца, без порока, Господу в жертву о грехе,
LEV|4|4|и приведет тельца к дверям скинии собрания пред Господа, и возложит руки свои на голову тельца, и заколет тельца пред Господом;
LEV|4|5|и возьмет священник помазанный, крови тельца и внесет ее в скинию собрания,
LEV|4|6|и омочит священник перст свой в кровь и покропит кровью семь раз пред Господом пред завесою святилища;
LEV|4|7|и возложит священник крови [тельца] пред Господом на роги жертвенника благовонных курений, который в скинии собрания, а остальную кровь тельца выльет к подножию жертвенника всесожжений, который у входа скинии собрания;
LEV|4|8|и вынет из тельца за грех весь тук его, тук, покрывающий внутренности, и весь тук, который на внутренностях,
LEV|4|9|и обе почки и тук, который на них, который на стегнах, и сальник на печени; с почками отделит он это,
LEV|4|10|как отделяется из тельца жертвы мирной; и сожжет их священник на жертвеннике всесожжения;
LEV|4|11|а кожу тельца и все мясо его с головою и с ногами его, и внутренности его и нечистоту его,
LEV|4|12|всего тельца пусть вынесет вне стана на чистое место, где высыпается пепел, и сожжет его огнем на дровах; где высыпается пепел, там пусть сожжен будет.
LEV|4|13|Если же все общество Израилево согрешит по ошибке и скрыто будет дело от глаз собрания, и сделает что–нибудь против заповедей Господних, чего не надлежало делать, и будет виновно,
LEV|4|14|то, когда узнан будет грех, которым они согрешили, пусть от всего общества представят они из крупного скота тельца в жертву за грех и приведут его пред скинию собрания;
LEV|4|15|и возложат старейшины общества руки свои на голову тельца пред Господом и заколют тельца пред Господом.
LEV|4|16|И внесет священник помазанный крови тельца в скинию собрания,
LEV|4|17|и омочит священник перст свой в кровь и покропит семь раз пред Господом пред завесою [святилища];
LEV|4|18|и возложит крови на роги жертвенника, который пред лицем Господним в скинии собрания, а остальную кровь выльет к подножию жертвенника всесожжений, который у входа скинии собрания;
LEV|4|19|и весь тук его вынет из него и сожжет на жертвеннике;
LEV|4|20|и сделает с тельцом то, что делается с тельцом за грех; так должен сделать с ним, и так очистит их священник, и прощено будет им;
LEV|4|21|и вынесет тельца вне стана, и сожжет его так, как сожег прежнего тельца. Это жертва за грех общества.
LEV|4|22|А если согрешит начальник, и сделает по ошибке что–нибудь против заповедей Господа, Бога своего, чего не надлежало делать, и будет виновен,
LEV|4|23|то, когда узнан будет им грех, которым он согрешил, пусть приведет он в жертву козла без порока,
LEV|4|24|и возложит руку свою на голову козла, и заколет его на месте, где заколаются всесожжения пред Господом: это жертва за грех;
LEV|4|25|и возьмет священник перстом своим крови от жертвы за грех и возложит на роги жертвенника всесожжения, а остальную кровь его выльет к подножию жертвенника всесожжения;
LEV|4|26|и весь тук его сожжет на жертвеннике, подобно как тук жертвы мирной, и так очистит его священник от греха его, и прощено будет ему.
LEV|4|27|Если же кто из народа земли согрешит по ошибке и сделает что–нибудь против заповедей Господних, чего не надлежало делать, и виновен будет,
LEV|4|28|то, когда узнан будет им грех, которым он согрешил, пусть приведет он в жертву козу без порока за грех свой, которым он согрешил,
LEV|4|29|и возложит руку свою на голову жертвы за грех, и заколют [козу] в жертву за грех на месте, [где заколают] жертву всесожжения;
LEV|4|30|и возьмет священник крови ее перстом своим, и возложит на роги жертвенника всесожжения, а остальную кровь ее выльет к подножию жертвенника;
LEV|4|31|и весь тук ее отделит, подобно как отделяется тук из жертвы мирной, и сожжет [его] священник на жертвеннике в приятное благоухание Господу; и так очистит его священник, и прощено будет ему.
LEV|4|32|А если из стада овец захочет он принести жертву за грех, пусть принесет женского пола, без порока,
LEV|4|33|и возложит руку свою на голову жертвы за грех, и заколет ее в жертву за грех на том месте, где заколают жертву всесожжения;
LEV|4|34|и возьмет священник перстом своим крови от сей жертвы за грех и возложит на роги жертвенника всесожжения, а остальную кровь ее выльет к подножию жертвенника;
LEV|4|35|и весь тук ее отделит, как отделяется тук овцы из жертвы мирной, и сожжет сие священник на жертвеннике в жертву Господу; и так очистит его священник от греха, которым он согрешил, и прощено будет ему.
LEV|5|1|Если кто согрешит тем, что слышал голос проклятия и был свидетелем, или видел, или знал, но не объявил, то он понесет на себе грех.
LEV|5|2|Или если прикоснется к чему–нибудь нечистому, или к трупу зверя нечистого, или к трупу скота нечистого, или к трупу гада нечистого, но не знал того, то он нечист и виновен.
LEV|5|3|Или если прикоснется к нечистоте человеческой, какая бы то ни была нечистота, от которой оскверняются, и он не знал того, но после узнает, то он виновен.
LEV|5|4|Или если кто безрассудно устами своими поклянется сделать что–нибудь худое или доброе, какое бы то ни было дело, в котором люди безрассудно клянутся, и он не знал того, но после узнает, то он виновен в том.
LEV|5|5|Если он виновен в чем–нибудь из сих, и исповедается, в чем он согрешил,
LEV|5|6|то пусть принесет Господу за грех свой, которым он согрешил, жертву повинности из мелкого скота, овцу или козу, за грех, и очистит его священник от греха его.
LEV|5|7|Если же он не в состоянии принести овцы, то в повинность за грех свой пусть принесет Господу двух горлиц или двух молодых голубей, одного в жертву за грех, а другого во всесожжение;
LEV|5|8|пусть принесет их к священнику, и [священник] представит прежде ту [из сих птиц], которая за грех, и надломит голову ее от шеи ее, но не отделит;
LEV|5|9|и покропит кровью сей жертвы за грех на стену жертвенника, а остальную кровь выцедит к подножию жертвенника: это жертва за грех;
LEV|5|10|а другую употребит во всесожжение по установлению; и так очистит его священник от греха его, которым он согрешил, и прощено будет ему.
LEV|5|11|Если же он не в состоянии принести двух горлиц или двух молодых голубей, пусть принесет за то, что согрешил, десятую часть ефы пшеничной муки в жертву за грех; пусть не льет на нее елея, и ливана пусть не кладет на нее, ибо это жертва за грех;
LEV|5|12|и принесет ее к священнику, а священник возьмет из нее полную горсть в память и сожжет на жертвеннике в жертву Господу: это жертва за грех;
LEV|5|13|и так очистит его священник от греха его, которым он согрешил в котором–нибудь из оных [случаев], и прощено будет ему; [остаток] же принадлежит священнику, как приношение хлебное.
LEV|5|14|И сказал Господь Моисею, говоря:
LEV|5|15|если кто сделает преступление и по ошибке согрешит против посвященного Господу, пусть за вину свою принесет Господу из стада овец овна без порока, по твоей оценке, серебряными сиклями по сиклю священному, в жертву повинности;
LEV|5|16|за ту святыню, против которой он согрешил, пусть воздаст и прибавит к тому пятую долю, и отдаст сие священнику, и священник очистит его овном жертвы повинности, и прощено будет ему.
LEV|5|17|Если кто согрешит и сделает что–нибудь против заповедей Господних, чего не надлежало делать, и по неведению сделается виновным и понесет на себе грех,
LEV|5|18|пусть принесет к священнику в жертву повинности овна без порока, по оценке твоей, и загладит священник проступок его, в чем он преступил по неведению, и прощено будет ему.
LEV|5|19|Это жертва повинности, [которою] он провинился пред Господом.
LEV|5|20|И сказал Господь Моисею, говоря:
LEV|5|21|если кто согрешит и сделает преступление пред Господом и запрется пред ближним своим в том, что ему поручено, или у него положено, или им похищено, или обманет ближнего своего,
LEV|5|22|или найдет потерянное и запрется в том, и поклянется ложно в чем–нибудь, что люди делают и тем грешат, –
LEV|5|23|то, согрешив и сделавшись виновным, он должен возвратить похищенное, что похитил, или отнятое, что отнял, или порученное, что ему поручено, или потерянное, что он нашел;
LEV|5|24|или если он в чем поклялся ложно, то должен отдать сполна, и приложить к тому пятую долю и отдать тому, кому принадлежит, в день приношения жертвы повинности;
LEV|5|25|и за вину свою пусть принесет Господу к священнику в жертву повинности из стада овец овна без порока, по оценке твоей;
LEV|5|26|и очистит его священник пред Господом, и прощено будет ему, что бы он ни сделал, все, в чем он сделался виновным.
LEV|6|1|И сказал Господь Моисею, говоря:
LEV|6|2|заповедай Аарону и сынам его: вот закон всесожжения: всесожжение пусть остается на месте сожигания на жертвеннике всю ночь до утра, и огонь жертвенника пусть горит на нем.
LEV|6|3|и пусть священник оденется в льняную одежду свою, и наденет на тело свое льняное нижнее платье, и снимет пепел от всесожжения, которое сжег огонь на жертвеннике, и положит его подле жертвенника;
LEV|6|4|и пусть снимет с себя одежды свои, и наденет другие одежды, и вынесет пепел вне стана на чистое место;
LEV|6|5|а огонь на жертвеннике пусть горит, не угасает; и пусть священник зажигает на нем дрова каждое утро, и раскладывает на нем всесожжение, и сожигает на нем тук мирной жертвы;
LEV|6|6|огонь непрестанно пусть горит на жертвеннике [и] не угасает.
LEV|6|7|Вот закон о приношении хлебном: сыны Аароновы должны приносить его пред Господа к жертвеннику;
LEV|6|8|и пусть возьмет [священник] горстью своею из приношения хлебного и пшеничной муки и елея и весь ливан, который на жертве, и сожжет на жертвеннике: [это] приятное благоухание, в память пред Господом;
LEV|6|9|а остальное из него пусть едят Аарон и сыны его; пресным должно есть его на святом месте, на дворе скинии собрания пусть едят его;
LEV|6|10|не должно печь его квасным. Сие даю Я им в долю из жертв Моих. Это великая святыня, подобно как жертва за грех и жертва повинности.
LEV|6|11|Все потомки Аароновы мужеского пола могут есть ее. Это вечный участок в роды ваши из жертв Господних. Все, прикасающееся к ним, освятится.
LEV|6|12|И сказал Господь Моисею, говоря:
LEV|6|13|вот приношение от Аарона и сынов его, которое принесут они Господу в день помазания его: десятая часть ефы пшеничной муки в жертву постоянную, половина сего для утра и половина для вечера;
LEV|6|14|на сковороде в елее она должна быть приготовлена; напитанную [елеем] приноси ее в кусках, как разламывается в куски приношение хлебное; приноси ее в приятное благоухание Господу;
LEV|6|15|и священник, помазанный на место его из сынов его, должен совершать сие: это вечный устав Господа. Вся она должна быть сожжена;
LEV|6|16|и всякое хлебное приношение от священника все да будет сожигаемо, а не съедаемо.
LEV|6|17|И сказал Господь Моисею, говоря:
LEV|6|18|скажи Аарону и сынам его: вот закон о жертве за грех: жертва за грех должна быть заколаема пред Господом на том месте, где заколается всесожжение; это великая святыня;
LEV|6|19|священник, совершающий жертву за грех, должен есть ее; она должна быть съедаема на святом месте, на дворе скинии собрания;
LEV|6|20|все, что прикоснется к мясу ее, освятится; и если кровью ее обрызгана будет одежда, то обрызганное омой на святом месте;
LEV|6|21|глиняный сосуд, в котором она варилась, должно разбить; если же она варилась в медном сосуде, то должно его вычистить и вымыть водою;
LEV|6|22|весь мужеский пол священнического рода может есть ее: это великая святыня.
LEV|6|23|а всякая жертва за грех, от которой кровь вносится в скинию собрания для очищения во святилище, не должна быть съедаема; ее должно сожигать на огне.
LEV|7|1|Вот закон о жертве повинности: это великая святыня;
LEV|7|2|жертву повинности должно заколать на том месте, где заколается всесожжение, и кровью ее кропить на жертвенник со всех сторон;
LEV|7|3|[приносящий] должен представить из нее весь тук, курдюк и тук, покрывающий внутренности,
LEV|7|4|и обе почки и тук, который на них, который на стегнах, и сальник, который на печени; с почками пусть он отделит сие;
LEV|7|5|и сожжет сие священник на жертвеннике в жертву Господу: это жертва повинности.
LEV|7|6|Весь мужеский пол священнического рода может есть ее; на святом месте должно есть ее: это великая святыня.
LEV|7|7|Как о жертве за грех, так и о жертве повинности закон один: она принадлежит священнику, который очищает посредством ее.
LEV|7|8|И когда священник приносит чью–нибудь жертву всесожжения, кожа от [жертвы] всесожжения, которое он приносит, принадлежит священнику;
LEV|7|9|и всякое приношение хлебное, которое печено в печи, и всякое приготовленное в горшке или на сковороде, принадлежит священнику, приносящему его;
LEV|7|10|и всякое приношение хлебное, смешанное с елеем и сухое, принадлежит всем сынам Аароновым, как одному, так и другому.
LEV|7|11|Вот закон о жертве мирной, которую приносят Господу:
LEV|7|12|если кто в благодарность приносит ее, то при жертве благодарности он должен принести пресные хлебы, смешанные с елеем, и пресные лепешки, помазанные елеем, и пшеничную муку, напитанную [елеем], хлебы, смешанные с елеем;
LEV|7|13|кроме лепешек пусть он приносит в приношение свое квасный хлеб, при мирной жертве благодарной;
LEV|7|14|одно что–нибудь из всего приношения своего пусть принесет он в возношение Господу: это принадлежит священнику, кропящему кровью мирной жертвы;
LEV|7|15|мясо мирной жертвы благодарности должно съесть в день приношения ее, не должно оставлять от него до утра.
LEV|7|16|Если же кто приносит жертву по обету, или от усердия, то жертву его должно есть в день приношения, и на другой день оставшееся от нее есть можно,
LEV|7|17|а оставшееся от жертвенного мяса к третьему дню должно сжечь на огне;
LEV|7|18|если же будут есть мясо мирной жертвы на третий день, то она не будет благоприятна; кто ее принесет, тому ни во что не вменится: это осквернение, и кто будет есть ее, тот понесет на себе грех;
LEV|7|19|мяса сего, если оно прикоснется к чему–либо нечистому, не должно есть, но должно сжечь его на огне; а мясо чистое может есть всякий чистый;
LEV|7|20|если же какая душа, имея на себе нечистоту, будет есть мясо мирной жертвы Господней, то истребится душа та из народа своего;
LEV|7|21|и если какая душа, прикоснувшись к чему–нибудь нечистому, к нечистоте человеческой, или к нечистому скоту, или какому–нибудь нечистому гаду, будет есть мясо мирной жертвы Господней, то истребится душа та из народа своего.
LEV|7|22|И сказал Господь Моисею, говоря:
LEV|7|23|скажи сынам Израилевым: никакого тука ни из вола, ни из овцы, ни из козла не ешьте.
LEV|7|24|Тук из мертвого и тук из растерзанного зверем можно употреблять на всякое дело; а есть не ешьте его;
LEV|7|25|ибо, кто будет есть тук из скота, который приносится в жертву Господу, истребится душа та из народа своего;
LEV|7|26|и никакой крови не ешьте во всех жилищах ваших ни из птиц, ни из скота;
LEV|7|27|а кто будет есть какую–нибудь кровь, истребится душа та из народа своего.
LEV|7|28|И сказал Господь Моисею, говоря:
LEV|7|29|скажи сынам Израилевым: кто представляет мирную жертву свою Господу, тот из мирной жертвы часть должен принести в приношение Господу;
LEV|7|30|своими руками должен он принести в жертву Господу: тук с грудью должен он принести, потрясая грудь пред лицем Господним;
LEV|7|31|тук сожжет священник на жертвеннике, а грудь принадлежит Аарону и сынам его;
LEV|7|32|и правое плечо, как возношение, из мирных жертв ваших отдавайте священнику:
LEV|7|33|кто из сынов Аароновых приносит кровь из мирной жертвы и тук, тому и правое плечо на долю;
LEV|7|34|ибо Я беру от сынов Израилевых из мирных жертв их грудь потрясания и плечо возношения, и отдаю их Аарону священнику и сынам его в вечный участок от сынов Израилевых.
LEV|7|35|Вот участок Аарону и участок сынам его из жертв Господних со дня, когда они предстанут пред Господа для священнодействия,
LEV|7|36|который повелел Господь давать им со дня помазания их от сынов Израилевых. [Это] вечное постановление в роды их. –
LEV|7|37|Вот закон о всесожжении, о приношении хлебном, о жертве за грех, о жертве повинности, о жертве посвящения и о жертве мирной,
LEV|7|38|который дал Господь Моисею на горе Синае, когда повелел сынам Израилевым, в пустыне Синайской, приносить Господу приношения их.
LEV|8|1|И сказал Господь Моисею, говоря:
LEV|8|2|возьми Аарона и сынов его с ним, и одежды и елей помазания, и тельца для жертвы за грех и двух овнов, и корзину опресноков,
LEV|8|3|и собери все общество ко входу скинии собрания.
LEV|8|4|Моисей сделал так, как повелел ему Господь, и собралось общество ко входу скинии собрания.
LEV|8|5|И сказал Моисей к обществу: вот что повелел Господь сделать.
LEV|8|6|И привел Моисей Аарона и сынов его и омыл их водою;
LEV|8|7|и возложил на него хитон, и опоясал его поясом, и надел на него верхнюю ризу, и возложил на него ефод, и опоясал его поясом ефода и прикрепил им ефод на нем,
LEV|8|8|и возложил на него наперсник, и на наперсник положил урим и туммим,
LEV|8|9|и возложил на голову его кидар, а на кидар с передней стороны его возложил полированную дощечку, диадиму святыни, как повелел Господь Моисею.
LEV|8|10|И взял Моисей елей помазания, и помазал скинию и все, что в ней, и освятил это;
LEV|8|11|и покропил им на жертвенник семь раз, и помазал жертвенник и все принадлежности его и умывальницу и подножие ее, чтобы освятить их;
LEV|8|12|и возлил елей помазания на голову Аарона и помазал его, чтоб освятить его.
LEV|8|13|И привел Моисей сынов Аароновых, и одел их в хитоны, и опоясал их поясом, и возложил на них кидары, как повелел Господь Моисею.
LEV|8|14|И привел тельца для жертвы за грех, и Аарон и сыны его возложили руки свои на голову тельца за грех;
LEV|8|15|и заколол [его] и взял крови, и перстом своим возложил на роги жертвенника со всех сторон, и очистил жертвенник, а [остальную] кровь вылил к подножию жертвенника, и освятил его, чтобы сделать его чистым.
LEV|8|16|И взял весь тук, который на внутренностях, и сальник на печени, и обе почки и тук их, и сжег Моисей на жертвеннике;
LEV|8|17|а тельца и кожу его, и мясо его, и нечистоту его сжег на огне вне стана, как повелел Господь Моисею.
LEV|8|18|И привел овна для всесожжения, и возложили Аарон и сыны его руки свои на голову овна;
LEV|8|19|и заколол [его] Моисей и покропил кровью на жертвенник со всех сторон;
LEV|8|20|и рассек овна на части, и сжег Моисей голову и части и тук,
LEV|8|21|а внутренности и ноги вымыл водою, и сжег Моисей всего овна на жертвеннике: это всесожжение в приятное благоухание, это жертва Господу, как повелел Господь Моисею.
LEV|8|22|И привел другого овна, овна посвящения, и возложили Аарон и сыны его руки свои на голову овна;
LEV|8|23|и заколол [его] Моисей, и взял крови его, и возложил на край правого уха Ааронова и на большой палец правой руки его и на большой палец правой ноги его.
LEV|8|24|И привел Моисей сынов Аароновых, и возложил крови на край правого уха их и на большой палец правой руки их и на большой палец правой ноги их, и покропил Моисей кровью на жертвенник со всех сторон.
LEV|8|25|И взял тук и курдюк и весь тук, который на внутренностях, и сальник на печени, и обе почки и тук их и правое плечо;
LEV|8|26|и из корзины с опресноками, которая пред Господом, взял один опреснок и один хлеб с елеем и одну лепешку, и возложил на тук и на правое плечо;
LEV|8|27|и положил все это на руки Аарону и на руки сынам его, и принес это, потрясая пред лицем Господним;
LEV|8|28|и взял это Моисей с рук их и сжег на жертвеннике со всесожжением: это жертва посвящения в приятное благоухание, это жертва Господу.
LEV|8|29|И взял Моисей грудь и принес ее, потрясая пред лицем Господним: это была доля Моисеева от овна посвящения, как повелел Господь Моисею.
LEV|8|30|И взял Моисей елея помазания и крови, которая на жертвеннике, и покропил Аарона и одежды его, и сынов его и одежды сынов его с ним; и так освятил Аарона и одежды его, и сынов его и одежды сынов его с ним.
LEV|8|31|И сказал Моисей Аарону и сынам его: сварите мясо у входа скинии собрания и там ешьте его с хлебом, который в корзине посвящения, как мне повелено и сказано: Аарон и сыны его должны есть его;
LEV|8|32|а остатки мяса и хлеба сожгите на огне.
LEV|8|33|Семь дней не отходите от дверей скинии собрания, пока не исполнятся дни посвящения вашего, ибо семь дней должно совершаться посвящение ваше;
LEV|8|34|как сегодня было сделано, так повелел Господь делать для очищения вас;
LEV|8|35|у входа скинии собрания будьте день и ночь в продолжение семи дней и будьте на страже у Господа, чтобы не умереть, ибо так мне повелено [от Господа Бога].
LEV|8|36|И исполнил Аарон и сыны его все, что повелел Господь чрез Моисея.
LEV|9|1|В восьмой день призвал Моисей Аарона и сынов его и старейшин Израилевых
LEV|9|2|и сказал Аарону: возьми себе из волов тельца в жертву за грех и овна во всесожжение, обоих без порока, и представь пред лице Господне;
LEV|9|3|и сынам Израилевым скажи: возьмите козла в жертву за грех, и тельца, и агнца, однолетних, без порока, во всесожжение,
LEV|9|4|и вола и овна в жертву мирную, чтобы совершить жертвоприношение пред лицем Господним, и приношение хлебное, смешанное с елеем, ибо сегодня Господь явится вам.
LEV|9|5|И принесли то, что приказал Моисей, пред скинию собрания, и пришло все общество и стало пред лицем Господним.
LEV|9|6|И сказал Моисей: вот что повелел Господь сделать, и явится вам слава Господня.
LEV|9|7|И сказал Моисей Аарону: приступи к жертвеннику и соверши жертву твою о грехе и всесожжение твое, и очисти себя и народ, и сделай приношение от народа, и очисти их, как повелел Господь.
LEV|9|8|И приступил Аарон к жертвеннику и заколол тельца, который за него, в жертву за грех:
LEV|9|9|сыны Аарона поднесли ему кровь, и он омочил перст свой в крови и возложил на роги жертвенника, а [остальную] кровь вылил к подножию жертвенника,
LEV|9|10|а тук и почки и сальник на печени от жертвы за грех сжег на жертвеннике, как повелел Господь Моисею;
LEV|9|11|мясо же и кожу сжег на огне вне стана.
LEV|9|12|И заколол всесожжение, и сыны Аарона поднесли ему кровь; он покропил ею на жертвенник со всех сторон;
LEV|9|13|и принесли ему всесожжение в кусках и голову, и он сжег на жертвеннике,
LEV|9|14|а внутренности и ноги омыл и сжег со всесожжением на жертвеннике.
LEV|9|15|И принес приношение от народа, и взял от народа козла за грех, и заколол его, и принес его в жертву за грех, как и прежнего.
LEV|9|16|И принес всесожжение и совершил его по уставу.
LEV|9|17|И принес приношение хлебное, и наполнил им руки свои, и сжег на жертвеннике сверх утреннего всесожжения.
LEV|9|18|И заколол вола и овна, которые от народа, в жертву мирную; и сыны Аарона поднесли ему кровь, и он покропил ею на жертвенник со всех сторон;
LEV|9|19|[поднесли] и тук из вола, и из овна курдюк, и [тук] покрывающий [внутренности], почки и сальник на печени,
LEV|9|20|и положили тук на грудь, и он сжег тук на жертвеннике;
LEV|9|21|грудь же и правое плечо принес Аарон, потрясая пред лицем Господним, как повелел Моисей.
LEV|9|22|И поднял Аарон руки свои, [обратившись] к народу, и благословил его, и сошел, совершив жертву за грех, всесожжение и жертву мирную.
LEV|9|23|И вошли Моисей и Аарон в скинию собрания, и вышли, и благословили народ. И явилась слава Господня всему народу:
LEV|9|24|и вышел огонь от Господа и сжег на жертвеннике всесожжение и тук; и видел весь народ, и воскликнул от радости, и пал на лице свое.
LEV|10|1|Надав и Авиуд, сыны Аароновы, взяли каждый свою кадильницу, и положили в них огня, и вложили в него курений, и принесли пред Господа огонь чуждый, которого Он не велел им;
LEV|10|2|и вышел огонь от Господа и сжег их, и умерли они пред лицем Господним.
LEV|10|3|И сказал Моисей Аарону: вот о чем говорил Господь, когда сказал: в приближающихся ко Мне освящусь и пред всем народом прославлюсь. Аарон молчал.
LEV|10|4|И позвал Моисей Мисаила и Елцафана, сынов Узиила, дяди Ааронова, и сказал им: пойдите, вынесите братьев ваших из святилища за стан.
LEV|10|5|И пошли и вынесли их в хитонах их за стан, как сказал Моисей.
LEV|10|6|Аарону же и Елеазару и Ифамару, сынам его, Моисей сказал: голов ваших не обнажайте и одежд ваших не раздирайте, чтобы вам не умереть и не навести гнева на все общество; но братья ваши, весь дом Израилев, могут плакать о сожженных, которых сожег Господь,
LEV|10|7|и из дверей скинии собрания не выходите, чтобы не умереть вам, ибо на вас елей помазания Господня. И сделали по слову Моисея.
LEV|10|8|И сказал Господь Аарону, говоря:
LEV|10|9|вина и крепких напитков не пей ты и сыны твои с тобою, когда входите в скинию собрания, чтобы не умереть. [Это] вечное постановление в роды ваши,
LEV|10|10|чтобы вы могли отличать священное от несвященного и нечистое от чистого,
LEV|10|11|и научать сынов Израилевых всем уставам, которые изрек им Господь чрез Моисея.
LEV|10|12|И сказал Моисей Аарону и Елеазару и Ифамару, оставшимся сынам его: возьмите приношение хлебное, оставшееся от жертв Господних, и ешьте его пресное у жертвенника, ибо это великая святыня;
LEV|10|13|и ешьте его на святом месте, ибо это участок твой и участок сынов твоих из жертв Господних: так мне повелено [от Господа];
LEV|10|14|и грудь потрясания и плечо возношения ешьте на чистом месте, ты и сыновья твои и дочери твои с тобою, ибо это дано в участок тебе и в участок сынам твоим из мирных жертв сынов Израилевых;
LEV|10|15|плечо возношения и грудь потрясания должны они приносить с жертвами тука, потрясая пред лицем Господним, и да будет это вечным участком тебе и сыновьям твоим с тобою, как повелел Господь.
LEV|10|16|И козла жертвы за грех искал Моисей, и вот, он сожжен. И разгневался на Елеазара и Ифамара, оставшихся сынов Аароновых, и сказал:
LEV|10|17|почему вы не ели жертвы за грех на святом месте? ибо она святыня великая, и она дана вам, чтобы снимать грехи с общества и очищать их пред Господом;
LEV|10|18|вот, кровь ее не внесена внутрь святилища, а вы должны были есть ее на святом месте, как повелено мне.
LEV|10|19|Аарон сказал Моисею: вот, сегодня принесли они жертву свою за грех и всесожжение свое пред Господом, и это случилось со мною; если я сегодня съем жертву за грех, будет ли это угодно Господу?
LEV|10|20|И услышал Моисей и одобрил.
LEV|11|1|И сказал Господь Моисею и Аарону, говоря им:
LEV|11|2|скажите сынам Израилевым: вот животные, которые можно вам есть из всего скота на земле:
LEV|11|3|всякий скот, у которого раздвоены копыта и на копытах глубокий разрез, и который жует жвачку, ешьте;
LEV|11|4|только сих не ешьте из жующих жвачку и имеющих раздвоенные копыта: верблюда, потому что он жует жвачку, но копыта у него не раздвоены, нечист он для вас;
LEV|11|5|и тушканчика, потому что он жует жвачку, но копыта у него не раздвоены, нечист он для вас,
LEV|11|6|и зайца, потому что он жует жвачку, но копыта у него не раздвоены, нечист он для вас;
LEV|11|7|и свиньи, потому что копыта у нее раздвоены и на копытах разрез глубокий, но она не жует жвачки, нечиста она для вас;
LEV|11|8|мяса их не ешьте и к трупам их не прикасайтесь; нечисты они для вас.
LEV|11|9|Из всех [животных], которые в воде, ешьте сих: у которых есть перья и чешуя в воде, в морях ли, или реках, тех ешьте;
LEV|11|10|а все те, у которых нет перьев и чешуи, в морях ли, или реках, из всех плавающих в водах и из всего живущего в водах, скверны для вас;
LEV|11|11|они должны быть скверны для вас: мяса их не ешьте и трупов их гнушайтесь;
LEV|11|12|все [животные], у которых нет перьев и чешуи в воде, скверны для вас.
LEV|11|13|Из птиц же гнушайтесь сих: орла, грифа и морского орла,
LEV|11|14|коршуна и сокола с породою его,
LEV|11|15|всякого ворона с породою его,
LEV|11|16|страуса, совы, чайки и ястреба с породою его,
LEV|11|17|филина, рыболова и ибиса,
LEV|11|18|лебедя, пеликана и сипа,
LEV|11|19|цапли, зуя с породою его, удода и нетопыря.
LEV|11|20|Все [животные] пресмыкающиеся, крылатые, ходящие на четырех [ногах], скверны для нас;
LEV|11|21|из всех пресмыкающихся, крылатых, ходящих на четырех [ногах], тех только ешьте, у которых есть голени выше ног, чтобы скакать ими по земле;
LEV|11|22|сих ешьте из них: саранчу с ее породою, солам с ее породою, харгол с ее породою и хагаб с ее породою.
LEV|11|23|Всякое [другое] пресмыкающееся, крылатое, у которого четыре ноги, скверно для вас;
LEV|11|24|от них вы будете нечисты: всякий, кто прикоснется к трупу их, нечист будет до вечера;
LEV|11|25|и всякий, кто возьмет труп их, должен омыть одежду свою и нечист будет до вечера.
LEV|11|26|Всякий скот, у которого копыта раздвоены, но нет глубокого разреза, и который не жует жвачки, нечист для вас: всякий, кто прикоснется к нему, будет нечист.
LEV|11|27|Из всех зверей четвероногих те, которые ходят на лапах, нечисты для вас: всякий, кто прикоснется к трупу их, нечист будет до вечера;
LEV|11|28|кто возьмет труп их, тот должен омыть одежды свои и нечист будет до вечера: нечисты они для вас.
LEV|11|29|Вот что нечисто для вас из животных, пресмыкающихся по земле: крот, мышь, ящерица с ее породою,
LEV|11|30|анака, хамелеон, летаа, хомет и тиншемет, –
LEV|11|31|сии нечисты для вас из всех пресмыкающихся: всякий, кто прикоснется к ним мертвым, нечист будет до вечера.
LEV|11|32|И все, на что упадет которое–нибудь из них мертвое, всякий деревянный сосуд, или одежда, или кожа, или мешок, и всякая вещь, которая употребляется на дело, будут нечисты: в воду должно положить их, и нечисты будут до вечера, потом будут чисты;
LEV|11|33|если же которое–нибудь из них упадет в какой–нибудь глиняный сосуд, то находящееся в нем будет нечисто, и самый [сосуд] разбейте.
LEV|11|34|Всякая пища, которую едят, на которой была вода [из такого] [сосуда], нечиста будет, и всякое питье, которое пьют, во всяком [таком] сосуде нечисто будет.
LEV|11|35|Все, на что упадет что–нибудь от трупа их, нечисто будет: печь и очаг должно разломать, они нечисты; и они должны быть нечисты для вас;
LEV|11|36|только источник и колодезь, вмещающий воду, остаются чистыми; а кто прикоснется к трупу их, тот нечист.
LEV|11|37|И если что–нибудь от трупа их упадет на какое–либо семя, которое сеют, то оно чисто;
LEV|11|38|если же тогда, как вода налита на семя, упадет на него что–нибудь от трупа их, то оно нечисто для вас.
LEV|11|39|И когда умрет какой–либо скот, который употребляется вами в пищу, то прикоснувшийся к трупу его нечист будет до вечера;
LEV|11|40|и тот, кто будет есть мертвечину его, должен омыть одежды свои и нечист будет до вечера; и тот, кто понесет труп его, должен омыть одежды свои и нечист будет до вечера.
LEV|11|41|Всякое животное, пресмыкающееся по земле, скверно для вас, не должно есть [его];
LEV|11|42|всего ползающего на чреве и всего ходящего на четырех ногах, и многоножных из животных пресмыкающихся по земле, не ешьте, ибо они скверны;
LEV|11|43|не оскверняйте душ ваших каким – либо животным пресмыкающимся и не делайте себя чрез них нечистыми, чтоб быть чрез них нечистыми,
LEV|11|44|ибо Я – Господь Бог ваш: освящайтесь и будьте святы, ибо Я свят; и не оскверняйте душ ваших каким–либо животным, ползающим по земле,
LEV|11|45|ибо Я – Господь, выведший вас из земли Египетской, чтобы быть вашим Богом. Итак будьте святы, потому что Я свят.
LEV|11|46|Вот закон о скоте, о птицах, о всех животных, живущих в водах, и о всех животных, пресмыкающихся по земле,
LEV|11|47|чтобы отличать нечистое от чистого, и животных, которых можно есть, от животных, которых есть не должно.
LEV|12|1|И сказал Господь Моисею, говоря:
LEV|12|2|скажи сынам Израилевым: если женщина зачнет и родит [младенца] мужеского пола, то она нечиста будет семь дней; как во дни страдания ее очищением, она будет нечиста;
LEV|12|3|в восьмой же день обрежется у него крайняя плоть его;
LEV|12|4|и тридцать три дня должна она сидеть, очищаясь от кровей своих; ни к чему священному не должна прикасаться и к святилищу не должна приходить, пока не исполнятся дни очищения ее.
LEV|12|5|Если же она родит [младенца] женского пола, то во время очищения своего она будет нечиста две недели, и шестьдесят шесть дней должна сидеть, очищаясь от кровей своих.
LEV|12|6|По окончании дней очищения своего за сына или за дочь она должна принести однолетнего агнца во всесожжение и молодого голубя или горлицу в жертву за грех, ко входу скинии собрания к священнику;
LEV|12|7|он принесет это пред Господа и очистит ее, и она будет чиста от течения кровей ее. Вот закон о родившей [младенца] мужеского или женского пола.
LEV|12|8|Если же она не в состоянии принести агнца, то пусть возьмет двух горлиц или двух молодых голубей, одного во всесожжение, а другого в жертву за грех, и очистит ее священник, и она будет чиста.
LEV|13|1|И сказал Господь Моисею и Аарону, говоря:
LEV|13|2|когда у кого появится на коже тела его опухоль, или лишаи, или пятно, и на коже тела его сделается как бы язва проказы, то должно привести его к Аарону священнику, или к одному из сынов его, священников;
LEV|13|3|священник осмотрит язву на коже тела, и если волосы на язве изменились в белые, и язва оказывается углубленною в кожу тела его, то это язва проказы; священник, осмотрев его, объявит его нечистым.
LEV|13|4|А если на коже тела его пятно белое, но оно не окажется углубленным в кожу, и волосы на нем не изменились в белые, то священник [имеющего] язву должен заключить на семь дней;
LEV|13|5|в седьмой день священник осмотрит его, и если язва остается в своем виде и не распространяется язва по коже, то священник должен заключить его на другие семь дней;
LEV|13|6|в седьмой день опять священник осмотрит его, и если язва менее приметна и не распространилась язва по коже, то священник должен объявить его чистым: это лишаи, и пусть он омоет одежды свои, и будет чист.
LEV|13|7|Если же лишаи станут распространяться по коже, после того как он являлся к священнику для очищения, то он вторично должен явиться к священнику;
LEV|13|8|священник, увидев, что лишаи распространяются по коже, объявит его нечистым: это проказа.
LEV|13|9|Если будет на ком язва проказы, то должно привести его к священнику;
LEV|13|10|священник осмотрит, и если опухоль на коже бела, и волос изменился в белый, и на опухоли живое мясо,
LEV|13|11|то это застарелая проказа на коже тела его; и священник объявит его нечистым и заключит его, ибо он нечист.
LEV|13|12|Если же проказа расцветет на коже, и покроет проказа всю кожу больного от головы его до ног, сколько могут видеть глаза священника,
LEV|13|13|и увидит священник, что проказа покрыла все тело его, то он объявит больного чистым, потому что все превратилось в белое: он чист.
LEV|13|14|Когда же окажется на нем живое мясо, то он нечист;
LEV|13|15|священник, увидев живое мясо, объявит его нечистым; живое мясо нечисто: это проказа.
LEV|13|16|Если же живое мясо изменится и обратится в белое, пусть он придет к священнику;
LEV|13|17|священник осмотрит его, и если язва обратилась в белое, священник объявит больного чистым; он чист.
LEV|13|18|Если у кого на коже тела был нарыв и зажил,
LEV|13|19|и на месте нарыва появилась белая опухоль, или пятно белое или красноватое, то он должен явиться к священнику;
LEV|13|20|священник осмотрит его, и если оно окажется ниже кожи, и волос его изменился в белый, то священник объявит его нечистым: это язва проказы, она расцвела на нарыве;
LEV|13|21|если же священник увидит, что волос на ней не бел, и она не ниже кожи, и притом мало приметна, то священник заключит его на семь дней;
LEV|13|22|если она станет очень распространяться по коже, то священник объявит его нечистым: это язва;
LEV|13|23|если же пятно остается на своем месте и не распространяется, то это воспаление нарыва, и священник объявит его чистым.
LEV|13|24|Или если у кого на коже тела будет ожог, и на зажившем ожоге окажется красноватое или белое пятно,
LEV|13|25|и священник увидит, что волос на пятне изменился в белый, и оно окажется углубленным в коже, то это проказа, она расцвела на ожоге; и священник объявит его нечистым: это язва проказы;
LEV|13|26|если же священник увидит, что волос на пятне не бел, и оно не ниже кожи, и притом мало приметно, то священник заключит его на семь дней;
LEV|13|27|в седьмой день священник осмотрит его, и если оно очень распространяется по коже, то священник объявит его нечистым: это язва проказы;
LEV|13|28|если же пятно остается на своем месте и не распространяется по коже, и притом мало приметно, то это опухоль от ожога; священник объявит его чистым, ибо это воспаление от ожога.
LEV|13|29|Если у мужчины или у женщины будет язва на голове или на бороде,
LEV|13|30|и осмотрит священник язву, и она окажется углубленною в коже, и волос на ней желтоватый тонкий, то священник объявит их нечистыми: это паршивость, это проказа на голове или на бороде;
LEV|13|31|если же священник осмотрит язву паршивости и она не окажется углубленною в коже, и волос на ней не черный, то священник [имеющего] язву паршивости заключит на семь дней;
LEV|13|32|в седьмой день священник осмотрит язву, и если паршивость не распространяется, и нет на ней желтоватого волоса, и паршивость не окажется углубленною в коже,
LEV|13|33|то [больного] должно остричь, но паршивого места не остригать, и священник должен паршивого вторично заключить на семь дней;
LEV|13|34|в седьмой день священник осмотрит паршивость, и если паршивость не распространяется по коже и не окажется углубленною в коже, то священник объявит его чистым; пусть он омоет одежды свои, и будет чист.
LEV|13|35|Если же после очищения его будет очень распространяться паршивость по коже,
LEV|13|36|и священник увидит, что паршивость распространяется по коже, то священник пусть не ищет желтоватого волоса: он нечист.
LEV|13|37|Если же паршивость остается в своем виде, и показывается на ней волос черный, то паршивость прошла, он чист; священник объявит его чистым.
LEV|13|38|Если у мужчины или у женщины на коже тела их будут пятна, пятна белые,
LEV|13|39|и священник увидит, что на коже тела их пятна бледно–белые, то это лишай, расцветший на коже: он чист.
LEV|13|40|Если у кого на голове вылезли [волосы], то это плешивый: он чист;
LEV|13|41|а если на передней стороне головы вылезли [волосы], то это лысый: он чист.
LEV|13|42|Если же на плеши или на лысине будет белое или красноватое пятно, то на плеши его или на лысине его расцвела проказа;
LEV|13|43|священник осмотрит его, и если увидит, что опухоль язвы бела [или] красновата на плеши его или на лысине его, видом похожа на проказу кожи тела,
LEV|13|44|то он прокаженный, нечист он; священник должен объявить его нечистым, у него на голове язва.
LEV|13|45|У прокаженного, на котором эта язва, должна быть разодрана одежда, и голова его должна быть не покрыта, и до уст он должен быть закрыт и кричать: нечист! нечист!
LEV|13|46|Во все дни, доколе на нем язва, он должен быть нечист, нечист он; он должен жить отдельно, вне стана жилище его.
LEV|13|47|Если язва проказы будет на одежде, на одежде шерстяной, или на одежде льняной,
LEV|13|48|или на основе, или на утоке из льна или шерсти, или на коже, или на каком–нибудь изделии кожаном,
LEV|13|49|и пятно будет зеленоватое или красноватое на одежде, или на коже, или на основе, или на утоке, или на какой–нибудь кожаной вещи, – то это язва проказы: должно показать ее священнику;
LEV|13|50|священник осмотрит язву и заключит зараженное язвою на семь дней;
LEV|13|51|в седьмой день осмотрит священник зараженное, и если язва распространилась по одежде, или по основе, или по утоку, или по коже, или по какому–либо изделию, сделанному из кожи, то это проказа едкая, язва нечистая;
LEV|13|52|он должен сжечь одежду, или основу, или уток шерстяной или льняной, или какую бы то ни было кожаную вещь, на которой будет язва, ибо это проказа едкая: должно сжечь на огне.
LEV|13|53|Если же священник увидит, что язва не распространилась по одежде, или по основе, или по утоку, или по какой бы то ни было кожаной вещи,
LEV|13|54|то священник прикажет омыть то, на чем язва, и вторично заключит на семь дней;
LEV|13|55|если по омытии зараженной [вещи] священник увидит, что язва не изменила вида своего и не распространилась язва, то она нечиста, сожги ее на огне; это выеденная ямина на лицевой стороне или на изнанке;
LEV|13|56|если же священник увидит, что язва по омытии ее сделалась менее приметна, то священник пусть оторвет ее от одежды, или от кожи, или от основы, или от утока.
LEV|13|57|Если же она опять покажется на одежде, или на основе, или на утоке, или на какой–нибудь кожаной вещи, то это расцветающая язва: сожги на огне то, на чем язва.
LEV|13|58|Если же одежду, или основу, или уток, или какую–нибудь кожаную вещь вымоешь, и сойдет с них язва, то должно вымыть их вторично, и они будут чисты.
LEV|13|59|Вот закон о язве проказы на одежде шерстяной или льняной, или на основе и на утоке, или на какой–нибудь кожаной вещи, как объявлять ее чистою или нечистою.
LEV|14|1|И сказал Господь Моисею, говоря:
LEV|14|2|вот закон о прокаженном, когда надобно его очистить: приведут его к священнику;
LEV|14|3|священник выйдет вон из стана, и если священник увидит, что прокаженный исцелился от болезни прокажения,
LEV|14|4|то священник прикажет взять для очищаемого двух птиц живых чистых, кедрового дерева, червленую нить и иссопа,
LEV|14|5|и прикажет священник заколоть одну птицу над глиняным сосудом, над живою водою;
LEV|14|6|а сам он возьмет живую птицу, кедровое дерево, червленую нить и иссоп, и омочит их и живую птицу в крови птицы заколотой над живою водою,
LEV|14|7|и покропит на очищаемого от проказы семь раз, и объявит его чистым, и пустит живую птицу в поле.
LEV|14|8|Очищаемый омоет одежды свои, острижет все волосы свои, омоется водою, и будет чист; потом войдет в стан и пробудет семь дней вне шатра своего;
LEV|14|9|в седьмой день обреет все волосы свои, голову свою, бороду свою, брови глаз своих, все волосы свои обреет, и омоет одежды свои, и омоет тело свое водою, и будет чист;
LEV|14|10|в восьмой день возьмет он двух овнов без порока, и одну овцу однолетнюю без порока, и три десятых части ефы пшеничной муки, смешанной с елеем, в приношение хлебное, и один лог елея;
LEV|14|11|священник очищающий поставит очищаемого человека с ними пред Господом у входа скинии собрания;
LEV|14|12|и возьмет священник одного овна, и представит его в жертву повинности, и лог елея, и принесет это, потрясая пред Господом;
LEV|14|13|и заколет овна на том месте, где заколают жертву за грех и всесожжение, на месте святом, ибо сия жертва повинности, подобно жертве за грех, принадлежит священнику: это великая святыня;
LEV|14|14|и возьмет священник крови жертвы повинности, и возложит священник на край правого уха очищаемого и на большой палец правой руки его и на большой палец правой ноги его;
LEV|14|15|и возьмет священник из лога елея и польет на левую свою ладонь;
LEV|14|16|и омочит священник правый перст свой в елей, который на левой ладони его, и покропит елеем с перста своего семь раз пред лицем Господа;
LEV|14|17|оставшийся же елей, который на ладони его, возложит священник на край правого уха очищаемого, на большой палец правой руки его и на большой палец правой ноги его, на [места, где] кровь жертвы повинности;
LEV|14|18|а остальной елей, который на ладони священника, возложит он на голову очищаемого, и очистит его священник пред лицем Господа.
LEV|14|19|И совершит священник жертву за грех, и очистит очищаемого от нечистоты его; после того заколет [жертву] всесожжения;
LEV|14|20|и возложит священник всесожжение и приношение хлебное на жертвенник; и очистит его священник, и он будет чист.
LEV|14|21|Если же он беден и не имеет достатка, то пусть возьмет одного овна в жертву повинности для потрясания, чтоб очистить себя, и одну десятую часть [ефы] пшеничной муки, смешанной с елеем, в приношение хлебное, и лог елея,
LEV|14|22|и двух горлиц или двух молодых голубей, что достанет рука его, одну [из птиц] в жертву за грех, а другую во всесожжение;
LEV|14|23|и принесет их в восьмой день очищения своего к священнику ко входу скинии собрания, пред лице Господа;
LEV|14|24|священник возьмет овна жертвы повинности и лог елея, и принесет это священник, потрясая пред Господом;
LEV|14|25|и заколет овна в жертву повинности, и возьмет священник крови жертвы повинности, и возложит на край правого уха очищаемого и на большой палец правой руки его и на большой палец правой ноги его;
LEV|14|26|и нальет священник елея на левую свою ладонь,
LEV|14|27|и елеем, который на левой ладони его, покропит священник с правого перста своего семь раз пред лицем Господним;
LEV|14|28|и возложит священник елея, который на ладони его, на край правого уха очищаемого, на большой палец правой руки его и на большой палец правой ноги его, на места, [где] кровь жертвы повинности;
LEV|14|29|а остальной елей, который на ладони священника, возложит он на голову очищаемого, чтоб очистить его пред лицем Господа;
LEV|14|30|и принесет одну из горлиц или одного из молодых голубей, что достанет рука [очищаемого],
LEV|14|31|из того, что достанет рука его, одну [птицу] в жертву за грех, а другую во всесожжение, вместе с приношением хлебным; и очистит священник очищаемого пред лицем Господа.
LEV|14|32|Вот закон о прокаженном, который во время очищения своего не имеет достатка.
LEV|14|33|И сказал Господь Моисею и Аарону, говоря:
LEV|14|34|когда войдете в землю Ханаанскую, которую Я даю вам во владение, и Я наведу язву проказы на домы в земле владения вашего,
LEV|14|35|тогда тот, чей дом, должен пойти и сказать священнику: у меня на доме показалась как бы язва.
LEV|14|36|Священник прикажет опорожнить дом, прежде нежели войдет священник осматривать язву, чтобы не сделалось нечистым все, что в доме; после сего придет священник осматривать дом.
LEV|14|37|Если он, осмотрев язву, увидит, что язва на стенах дома состоит из зеленоватых или красноватых ямин, которые окажутся углубленными в стене,
LEV|14|38|то священник выйдет из дома к дверям дома и запрет дом на семь дней.
LEV|14|39|В седьмой день опять придет священник, и если увидит, что язва распространилась по стенам дома,
LEV|14|40|то священник прикажет выломать камни, на которых язва, и бросить их вне города на место нечистое;
LEV|14|41|а дом внутри пусть весь оскоблят, и обмазку, которую отскоблят, высыпят вне города на место нечистое;
LEV|14|42|и возьмут другие камни, и вставят вместо тех камней, и возьмут другую обмазку, и обмажут дом.
LEV|14|43|Если язва опять появится и будет цвести на доме после того, как выломали камни и оскоблили дом и обмазали,
LEV|14|44|то священник придет и осмотрит, и если язва на доме распространилась, то это едкая проказа на доме, нечист он;
LEV|14|45|должно разломать сей дом, и камни его и дерево его и всю обмазку дома вынести вне города на место нечистое;
LEV|14|46|кто входит в дом во все время, когда он заперт, тот нечист до вечера;
LEV|14|47|и кто спит в доме том, тот должен вымыть одежды свои; и кто ест в доме том, тот должен вымыть одежды свои.
LEV|14|48|Если же священник придет и увидит, что язва на доме не распространилась после того, как обмазали дом, то священник объявит дом чистым, потому что язва прошла.
LEV|14|49|И чтобы очистить дом, возьмет он две птицы, кедрового дерева, червленую нить и иссопа,
LEV|14|50|и заколет одну птицу над глиняным сосудом, над живою водою;
LEV|14|51|и возьмет кедровое дерево и иссоп, и червленую нить и живую птицу, и омочит их в крови птицы заколотой и в живой воде, и покропит дом семь раз;
LEV|14|52|и очистит дом кровью птицы и живою водою, и живою птицею и кедровым деревом, и иссопом и червленою нитью;
LEV|14|53|и пустит живую птицу вне города в поле и очистит дом, и будет чист.
LEV|14|54|Вот закон о всякой язве проказы и о паршивости,
LEV|14|55|и о проказе на одежде и на доме,
LEV|14|56|и об опухоли, и о лишаях, и о пятнах, –
LEV|14|57|чтобы указать, когда это нечисто и когда чисто. Вот закон о проказе.
LEV|15|1|И сказал Господь Моисею и Аарону, говоря:
LEV|15|2|объявите сынам Израилевым и скажите им: если у кого будет истечение из тела его, то от истечения своего он нечист.
LEV|15|3|И вот [закон] о нечистоте его от истечения его: когда течет из тела его истечение его, и когда задерживается в теле его истечение его, это нечистота его;
LEV|15|4|всякая постель, на которой ляжет имеющий истечение, нечиста, и всякая вещь, на которую сядет, нечиста;
LEV|15|5|и кто прикоснется к постели его, тот должен вымыть одежды свои и омыться водою и нечист будет до вечера;
LEV|15|6|кто сядет на какую–либо вещь, на которой сидел имеющий истечение, тот должен вымыть одежды свои и омыться водою и нечист будет до вечера;
LEV|15|7|и кто прикоснется к телу имеющего истечение, тот должен вымыть одежды свои и омыться водою и нечист будет до вечера;
LEV|15|8|если имеющий истечение плюнет на чистого, то сей должен вымыть одежды свои и омыться водою, и нечист будет до вечера;
LEV|15|9|и всякая повозка, в которой ехал имеющий истечение, нечиста [будет до вечера];
LEV|15|10|и всякий, кто прикоснется к чему–нибудь, что было под ним, нечист будет до вечера; и кто понесет это, должен вымыть одежды свои и омыться водою, и нечист будет до вечера;
LEV|15|11|и всякий, к кому прикоснется имеющий истечение, не омыв рук своих водою, должен вымыть одежды свои и омыться водою, и нечист будет до вечера;
LEV|15|12|глиняный сосуд, к которому прикоснется имеющий истечение, должно разбить, а всякий деревянный сосуд должно вымыть водою.
LEV|15|13|А когда имеющий истечение освободится от истечения своего, тогда должен он отсчитать себе семь дней для очищения своего и вымыть одежды свои, и омыть тело свое живою водою, и будет чист;
LEV|15|14|и в восьмой день возьмет он себе двух горлиц или двух молодых голубей, и придет пред лице Господне ко входу скинии собрания, и отдаст их священнику;
LEV|15|15|и принесет священник из сих [птиц] одну в жертву за грех, а другую во всесожжение, и очистит его священник пред Господом от истечения его.
LEV|15|16|Если у кого случится излияние семени, то он должен омыть водою все тело свое, и нечист будет до вечера;
LEV|15|17|и всякая одежда и всякая кожа, на которую попадет семя, должна быть вымыта водою, и нечиста будет до вечера;
LEV|15|18|если мужчина ляжет с женщиной и [будет] у него излияние семени, то они должны омыться водою, и нечисты будут до вечера.
LEV|15|19|Если женщина имеет истечение крови, текущей из тела ее, то она должна сидеть семь дней во время очищения своего, и всякий, кто прикоснется к ней, нечист будет до вечера;
LEV|15|20|и все, на чем она ляжет в продолжение очищения своего, нечисто; и все, на чем сядет, нечисто;
LEV|15|21|и всякий, кто прикоснется к постели ее, должен вымыть одежды свои и омыться водою и нечист будет до вечера;
LEV|15|22|и всякий, кто прикоснется к какой–нибудь вещи, на которой она сидела, должен вымыть одежды свои и омыться водою, и нечист будет до вечера;
LEV|15|23|и если кто прикоснется к чему–нибудь на постели или на той вещи, на которой она сидела, нечист будет до вечера;
LEV|15|24|если переспит с нею муж, то нечистота ее будет на нем; он нечист будет семь дней, и всякая постель, на которой он ляжет, будет нечиста.
LEV|15|25|Если у женщины течет кровь многие дни не во время очищения ее, или если она имеет истечение долее [обыкновенного] очищения ее, то во все время истечения нечистоты ее, подобно как в продолжение очищения своего, она нечиста;
LEV|15|26|всякая постель, на которой она ляжет во все время истечения своего, будет [нечиста], подобно как постель в продолжение очищения ее; и всякая вещь, на которую она сядет, будет нечиста, как нечисто это во время очищения ее;
LEV|15|27|и всякий, кто прикоснется к ним, будет нечист, и должен вымыть одежды свои и омыться водою, и нечист будет до вечера.
LEV|15|28|А когда она освободится от истечения своего, тогда должна отсчитать себе семь дней, и потом будет чиста;
LEV|15|29|в восьмой день возьмет она себе двух горлиц или двух молодых голубей и принесет их к священнику ко входу скинии собрания;
LEV|15|30|и принесет священник одну [из птиц] в жертву за грех, а другую во всесожжение, и очистит ее священник пред Господом от истечения нечистоты ее.
LEV|15|31|Так предохраняйте сынов Израилевых от нечистоты их, чтоб они не умерли в нечистоте своей, оскверняя жилище Мое, которое среди них:
LEV|15|32|вот закон об имеющем истечение и о том, у кого случится излияние семени, делающее его нечистым,
LEV|15|33|и о страдающей очищением своим, и о имеющих истечение, мужчине или женщине, и о муже, который переспит с нечистою.
LEV|16|1|И говорил Господь Моисею по смерти двух сынов Аароновых, когда они, приступив пред лице Господне, умерли,
LEV|16|2|и сказал Господь Моисею: скажи Аарону, брату твоему, чтоб он не во всякое время входил во святилище за завесу пред крышку, что на ковчеге, дабы ему не умереть, ибо над крышкою Я буду являться в облаке.
LEV|16|3|Вот с чем должен входить Аарон во святилище: с тельцом в жертву за грех и с овном во всесожжение;
LEV|16|4|священный льняной хитон должен надевать он, нижнее платье льняное да будет на теле его, и льняным поясом пусть опоясывается, и льняной кидар надевает: это священные одежды; и пусть омывает он тело свое водою и надевает их;
LEV|16|5|и от общества сынов Израилевых пусть возьмет двух козлов в жертву за грех и одного овна во всесожжение.
LEV|16|6|И принесет Аарон тельца в жертву за грех за себя и очистит себя и дом свой.
LEV|16|7|И возьмет двух козлов и поставит их пред лицем Господним у входа скинии собрания;
LEV|16|8|и бросит Аарон об обоих козлах жребии: один жребий для Господа, а другой жребий для отпущения;
LEV|16|9|и приведет Аарон козла, на которого вышел жребий для Господа, и принесет его в жертву за грех,
LEV|16|10|а козла, на которого вышел жребий для отпущения, поставит живого пред Господом, чтобы совершить над ним очищение и отослать его в пустыню для отпущения.
LEV|16|11|И приведет Аарон тельца в жертву за грех за себя, и очистит себя и дом свой, и заколет тельца в жертву за грех за себя;
LEV|16|12|и возьмет горящих угольев полную кадильницу с жертвенника, который пред лицем Господним, и благовонного мелко–истолченного курения полные горсти, и внесет за завесу;
LEV|16|13|и положит курение на огонь пред лицем Господним, и облако курения покроет крышку, которая над [ковчегом] откровения, дабы ему не умереть;
LEV|16|14|и возьмет крови тельца и покропит перстом своим на крышку спереди и пред крышкою, семь раз покропит кровью с перста своего.
LEV|16|15|И заколет козла в жертву за грех за народ, и внесет кровь его за завесу, и сделает с кровью его то же, что делал с кровью тельца и покропит ею на крышку и пред крышкою, –
LEV|16|16|и очистит святилище от нечистот сынов Израилевых и от преступлений их, во всех грехах их. Так должен поступить он и со скиниею собрания, находящеюся у них, среди нечистот их.
LEV|16|17|Ни один человек не должен быть в скинии собрания, когда входит он для очищения святилища, до самого выхода его. И так очистит он себя, дом свой и все общество Израилево.
LEV|16|18|И выйдет он к жертвеннику, который пред лицем Господним, и очистит его, и возьмет крови тельца и крови козла, и возложит на роги жертвенника со всех сторон,
LEV|16|19|и покропит на него кровью с перста своего семь раз, и очистит его, и освятит его от нечистот сынов Израилевых.
LEV|16|20|И совершив очищение святилища, скинии собрания и жертвенника, приведет он живого козла,
LEV|16|21|и возложит Аарон обе руки свои на голову живого козла, и исповедает над ним все беззакония сынов Израилевых и все преступления их и все грехи их, и возложит их на голову козла, и отошлет с нарочным человеком в пустыню:
LEV|16|22|и понесет козел на себе все беззакония их в землю непроходимую, и пустит он козла в пустыню.
LEV|16|23|И войдет Аарон в скинию собрания, и снимет льняные одежды, которые надевал, входя во святилище, и оставит их там,
LEV|16|24|и омоет тело свое водою на святом месте, и наденет одежды свои, и выйдет и совершит всесожжение за себя и всесожжение за народ, и очистит себя и народ;
LEV|16|25|а тук жертвы за грех воскурит на жертвеннике.
LEV|16|26|И тот, кто отводил козла для отпущения, должен вымыть одежды свои, омыть тело свое водою, и потом может войти в стан.
LEV|16|27|А тельца за грех и козла за грех, которых кровь внесена была для очищения святилища, пусть вынесут вон из стана и сожгут на огне кожи их и мясо их и нечистоту их;
LEV|16|28|кто сожжет их, тот должен вымыть одежды свои и омыть тело свое водою, и после того может войти в стан.
LEV|16|29|И да будет сие для вас вечным постановлением: в седьмой месяц, в десятый [день] месяца смиряйте души ваши и никакого дела не делайте, ни туземец, ни пришлец, поселившийся между вами,
LEV|16|30|ибо в сей день очищают вас, чтобы сделать вас чистыми от всех грехов ваших, чтобы вы были чисты пред лицем Господним;
LEV|16|31|это суббота покоя для вас, смиряйте души ваши: это постановление вечное.
LEV|16|32|Очищать же должен священник, который помазан и который посвящен, чтобы священнодействовать ему вместо отца своего: и наденет он льняные одежды, одежды священные,
LEV|16|33|и очистит Святое–святых и скинию собрания, и жертвенник очистит, и священников и весь народ общества очистит.
LEV|16|34|И да будет сие для вас вечным постановлением: очищать сынов Израилевых от всех грехов их однажды в году. И сделал он так, как повелел Господь Моисею.
LEV|17|1|И сказал Господь Моисею, говоря:
LEV|17|2|объяви Аарону и сынам его и всем сынам Израилевым и скажи им: вот что повелевает Господь:
LEV|17|3|если кто из дома Израилева заколет тельца или овцу или козу в стане, или если кто заколет вне стана
LEV|17|4|и не приведет ко входу скинии собрания, чтобы представить в жертву Господу пред жилищем Господним, то человеку тому вменена будет кровь: он пролил кровь, и истребится человек тот из народа своего;
LEV|17|5|[это] для того, чтобы приводили сыны Израилевы жертвы свои, которые они заколают на поле, чтобы приводили их пред Господа ко входу скинии собрания, к священнику, и заколали их Господу в жертвы мирные;
LEV|17|6|и покропит священник кровью на жертвенник Господень у входа скинии собрания и воскурит тук в приятное благоухание Господу,
LEV|17|7|чтоб они впредь не приносили жертв своих идолам, за которыми блудно ходят они. Сие да будет для них постановлением вечным в роды их.
LEV|17|8|[Еще] скажи им: если кто из дома Израилева и из пришельцев, которые живут между вами, приносит всесожжение или жертву
LEV|17|9|и не приведет ко входу скинии собрания, чтобы совершить ее Господу, то истребится человек тот из народа своего.
LEV|17|10|Если кто из дома Израилева и из пришельцев, которые живут между вами, будет есть какую–нибудь кровь, то обращу лице Мое на душу того, кто будет есть кровь, и истреблю ее из народа ее,
LEV|17|11|потому что душа тела в крови, и Я назначил ее вам для жертвенника, чтобы очищать души ваши, ибо кровь сия душу очищает;
LEV|17|12|потому Я и сказал сынам Израилевым: ни одна душа из вас не должна есть крови, и пришлец, живущий между вами, не должен есть крови.
LEV|17|13|Если кто из сынов Израилевых и из пришельцев, живущих между вами, на ловле поймает зверя или птицу, которую можно есть, то он должен дать вытечь крови ее и покрыть ее землею,
LEV|17|14|ибо душа всякого тела [есть] кровь его, она душа его; потому Я сказал сынам Израилевым: не ешьте крови ни из какого тела, потому что душа всякого тела есть кровь его: всякий, кто будет есть ее, истребится.
LEV|17|15|И всякий, кто будет есть мертвечину или растерзанное зверем, туземец или пришлец, должен вымыть одежды свои и омыться водою, и нечист будет до вечера, а [потом] будет чист;
LEV|17|16|если же не вымоет [одежд своих] и не омоет тела своего, то понесет на себе беззаконие свое.
LEV|18|1|И сказал Господь Моисею, говоря:
LEV|18|2|объяви сынам Израилевым и скажи им: Я Господь, Бог ваш.
LEV|18|3|По делам земли Египетской, в которой вы жили, не поступайте, и по делам земли Ханаанской, в которую Я веду вас, не поступайте, и по установлениям их не ходите:
LEV|18|4|Мои законы исполняйте и Мои постановления соблюдайте, поступая по ним. Я Господь, Бог ваш.
LEV|18|5|Соблюдайте постановления Мои и законы Мои, которые исполняя, человек будет жив. Я Господь.
LEV|18|6|Никто ни к какой родственнице по плоти не должен приближаться с тем, чтобы открыть наготу. Я Господь.
LEV|18|7|Наготы отца твоего и наготы матери твоей не открывай: она мать твоя, не открывай наготы ее.
LEV|18|8|Наготы жены отца твоего не открывай: это нагота отца твоего.
LEV|18|9|Наготы сестры твоей, дочери отца твоего или дочери матери твоей, родившейся в доме или вне дома, не открывай наготы их.
LEV|18|10|Наготы дочери сына твоего или дочери дочери твоей, не открывай наготы их, ибо они твоя нагота.
LEV|18|11|Наготы дочери жены отца твоего, родившейся от отца твоего, она сестра твоя [по отцу], не открывай наготы ее.
LEV|18|12|Наготы сестры отца твоего не открывай, она единокровная отцу твоему.
LEV|18|13|Наготы сестры матери твоей не открывай, ибо она единокровная матери твоей.
LEV|18|14|Наготы брата отца твоего не открывай и к жене его не приближайся: она тетка твоя.
LEV|18|15|Наготы невестки твоей не открывай: она жена сына твоего, не открывай наготы ее.
LEV|18|16|Наготы жены брата твоего не открывай, это нагота брата твоего.
LEV|18|17|Наготы жены и дочери ее не открывай; дочери сына ее и дочери дочери ее не бери, чтоб открыть наготу их, они единокровные ее; это беззаконие.
LEV|18|18|Не бери жены вместе с сестрою ее, чтобы сделать ее соперницею, чтоб открыть наготу ее при ней, при жизни ее.
LEV|18|19|И к жене во время очищения нечистот ее не приближайся, чтоб открыть наготу ее.
LEV|18|20|И с женою ближнего твоего не ложись, чтобы излить семя и оскверниться с нею.
LEV|18|21|Из детей твоих не отдавай на служение Молоху и не бесчести имени Бога твоего. Я Господь.
LEV|18|22|Не ложись с мужчиною, как с женщиною: это мерзость.
LEV|18|23|И ни с каким скотом не ложись, чтоб излить [семя] и оскверниться от него; и женщина не должна становиться пред скотом для совокупления с ним: это гнусно.
LEV|18|24|Не оскверняйте себя ничем этим, ибо всем этим осквернили себя народы, которых Я прогоняю от вас:
LEV|18|25|и осквернилась земля, и Я воззрел на беззаконие ее, и свергнула с себя земля живущих на ней.
LEV|18|26|А вы соблюдайте постановления Мои и законы Мои и не делайте всех этих мерзостей, ни туземец, ни пришлец, живущий между вами,
LEV|18|27|ибо все эти мерзости делали люди сей земли, что пред вами, и осквернилась земля;
LEV|18|28|чтоб и вас не свергнула с себя земля, когда вы станете осквернять ее, как она свергнула народы, бывшие прежде вас;
LEV|18|29|ибо если кто будет делать все эти мерзости, то души делающих это истреблены будут из народа своего.
LEV|18|30|Итак соблюдайте повеления Мои, чтобы не поступать по гнусным обычаям, по которым поступали прежде вас, и чтобы не оскверняться ими. Я Господь, Бог ваш.
LEV|19|1|И сказал Господь Моисею, говоря:
LEV|19|2|объяви всему обществу сынов Израилевых и скажи им: святы будьте, ибо свят Я Господь, Бог ваш.
LEV|19|3|Бойтесь каждый матери своей и отца своего и субботы Мои храните. Я Господь, Бог ваш.
LEV|19|4|Не обращайтесь к идолам и богов литых не делайте себе. Я Господь, Бог ваш.
LEV|19|5|Когда будете приносить Господу жертву мирную, то приносите ее, чтобы приобрести себе благоволение:
LEV|19|6|в день жертвоприношения вашего и на другой день должно есть ее, а оставшееся к третьему дню должно сжечь на огне;
LEV|19|7|если же кто станет есть ее на третий день, это гнусно, это не будет благоприятно;
LEV|19|8|кто станет есть ее, тот понесет на себе грех, ибо он осквернил святыню Господню, и истребится душа та из народа своего.
LEV|19|9|Когда будете жать жатву на земле вашей, не дожинай до края поля твоего, и оставшегося от жатвы твоей не подбирай,
LEV|19|10|и виноградника твоего не обирай дочиста, и попадавших ягод в винограднике не подбирай; оставь это бедному и пришельцу. Я Господь, Бог ваш.
LEV|19|11|Не крадите, не лгите и не обманывайте друг друга.
LEV|19|12|Не клянитесь именем Моим во лжи, и не бесчести имени Бога твоего. Я Господь.
LEV|19|13|Не обижай ближнего твоего и не грабительствуй. Плата наемнику не должна оставаться у тебя до утра.
LEV|19|14|Не злословь глухого и пред слепым не клади ничего, чтобы преткнуться ему; бойся Бога твоего. Я Господь.
LEV|19|15|Не делайте неправды на суде; не будь лицеприятен к нищему и не угождай лицу великого; по правде суди ближнего твоего.
LEV|19|16|Не ходи переносчиком в народе твоем и не восставай на жизнь ближнего твоего. Я Господь.
LEV|19|17|Не враждуй на брата твоего в сердце твоем; обличи ближнего твоего, и не понесешь за него греха.
LEV|19|18|Не мсти и не имей злобы на сынов народа твоего, но люби ближнего твоего, как самого себя. Я Господь.
LEV|19|19|Уставы Мои соблюдайте; скота твоего не своди с иною породою; поля твоего не засевай двумя родами [семян]; в одежду из разнородных нитей, из шерсти и льна, не одевайся.
LEV|19|20|Если кто переспит с женщиною, а она раба, обрученная мужу, но еще не выкупленная, или свобода еще не дана ей, то должно наказать их, но не смертью, потому что она несвободная:
LEV|19|21|пусть приведет он Господу ко входу скинии собрания жертву повинности, овна в жертву повинности своей;
LEV|19|22|и очистит его священник овном повинности пред Господом от греха, которым он согрешил, и прощен будет ему грех, которым он согрешил.
LEV|19|23|Когда придете в землю, [которую Господь Бог даст вам], и посадите какое–либо плодовое дерево, то плоды его почитайте за необрезанные: три года должно почитать их за необрезанные, не должно есть их;
LEV|19|24|а в четвертый год все плоды его должны быть посвящены для празднеств Господних;
LEV|19|25|в пятый же год вы можете есть плоды его и собирать себе все произведения его. Я Господь, Бог ваш.
LEV|19|26|Не ешьте с кровью; не ворожите и не гадайте.
LEV|19|27|Не стригите головы вашей кругом, и не порти края бороды твоей.
LEV|19|28|Ради умершего не делайте нарезов на теле вашем и не накалывайте на себе письмен. Я Господь.
LEV|19|29|Не оскверняй дочери твоей, допуская ее до блуда, чтобы не блудодействовала земля и не наполнилась земля развратом.
LEV|19|30|Субботы Мои храните и святилище Мое чтите. Я Господь.
LEV|19|31|Не обращайтесь к вызывающим мертвых, и к волшебникам не ходите, и не доводите себя до осквернения от них. Я Господь, Бог ваш.
LEV|19|32|Пред лицем седого вставай и почитай лице старца, и бойся Бога твоего. Я Господь.
LEV|19|33|Когда поселится пришлец в земле вашей, не притесняйте его:
LEV|19|34|пришлец, поселившийся у вас, да будет для вас то же, что туземец ваш; люби его, как себя; ибо и вы были пришельцами в земле Египетской. Я Господь, Бог ваш.
LEV|19|35|Не делайте неправды в суде, в мере, в весе и в измерении:
LEV|19|36|да будут у вас весы верные, гири верные, ефа верная и гин верный. Я Господь, Бог ваш, Который вывел вас из земли Египетской.
LEV|19|37|Соблюдайте все уставы Мои и все законы Мои и исполняйте их. Я Господь.
LEV|20|1|И сказал Господь Моисею, говоря:
LEV|20|2|скажи сие сынам Израилевым: кто из сынов Израилевых и из пришельцев, живущих между Израильтянами, даст из детей своих Молоху, тот да будет предан смерти: народ земли да побьет его камнями;
LEV|20|3|и Я обращу лице Мое на человека того и истреблю его из народа его за то, что он дал из детей своих Молоху, чтоб осквернить святилище Мое и обесчестить святое имя Мое;
LEV|20|4|и если народ земли не обратит очей своих на человека того, когда он даст из детей своих Молоху, и не умертвит его,
LEV|20|5|то Я обращу лице Мое на человека того и на род его и истреблю его из народа его, и всех блудящих по следам его, чтобы блудно ходить вслед Молоха.
LEV|20|6|И если какая душа обратится к вызывающим мертвых и к волшебникам, чтобы блудно ходить вслед их, то Я обращу лице Мое на ту душу и истреблю ее из народа ее.
LEV|20|7|Освящайте себя и будьте святы, ибо Я Господь, Бог ваш, [свят].
LEV|20|8|Соблюдайте постановления Мои и исполняйте их, ибо Я Господь, освящающий вас.
LEV|20|9|Кто будет злословить отца своего или мать свою, тот да будет предан смерти; отца своего и мать свою он злословил: кровь его на нем.
LEV|20|10|Если кто будет прелюбодействовать с женой замужнею, если кто будет прелюбодействовать с женою ближнего своего, – да будут преданы смерти и прелюбодей и прелюбодейка.
LEV|20|11|Кто ляжет с женою отца своего, тот открыл наготу отца своего: оба они да будут преданы смерти, кровь их на них.
LEV|20|12|Если кто ляжет с невесткою своею, то оба они да будут преданы смерти: мерзость сделали они, кровь их на них.
LEV|20|13|Если кто ляжет с мужчиною, как с женщиною, то оба они сделали мерзость: да будут преданы смерти, кровь их на них.
LEV|20|14|Если кто возьмет себе жену и мать ее: это беззаконие; на огне должно сжечь его и их, чтобы не было беззакония между вами.
LEV|20|15|Кто смесится со скотиною, того предать смерти, и скотину убейте.
LEV|20|16|Если женщина пойдет к какой–нибудь скотине, чтобы совокупиться с нею, то убей женщину и скотину: да будут они преданы смерти, кровь их на них.
LEV|20|17|Если кто возьмет сестру свою, дочь отца своего или дочь матери своей, и увидит наготу ее, и она увидит наготу его: это срам, да будут они истреблены пред глазами сынов народа своего; он открыл наготу сестры своей: грех свой понесет он.
LEV|20|18|Если кто ляжет с женою во время болезни [кровоочищения] и откроет наготу ее, то он обнажил истечения ее, и она открыла течение кровей своих: оба они да будут истреблены из народа своего.
LEV|20|19|Наготы сестры матери твоей и сестры отца твоего не открывай, ибо таковой обнажает плоть свою: грех свой понесут они.
LEV|20|20|Кто ляжет с теткою своею, тот открыл наготу дяди своего; грех свой понесут они, бездетными умрут.
LEV|20|21|Если кто возьмет жену брата своего: это гнусно; он открыл наготу брата своего, бездетны будут они.
LEV|20|22|Соблюдайте все уставы Мои и все законы Мои и исполняйте их, – и не свергнет вас с себя земля, в которую Я веду вас жить.
LEV|20|23|Не поступайте по обычаям народа, который Я прогоняю от вас; ибо они все это делали, и Я вознегодовал на них,
LEV|20|24|и сказал Я вам: вы владейте землею их, и вам отдаю в наследие землю, в которой течет молоко и мед. Я Господь, Бог ваш, Который отделил вас от всех народов.
LEV|20|25|Отличайте скот чистый от нечистого и птицу чистую от нечистой и не оскверняйте душ ваших скотом и птицею и всем пресмыкающимся по земле, что отличил Я, как нечистое.
LEV|20|26|Будьте предо Мною святы, ибо Я свят Господь, и Я отделил вас от народов, чтобы вы были Мои.
LEV|20|27|Мужчина ли или женщина, если будут они вызывать мертвых или волхвовать, да будут преданы смерти: камнями должно побить их, кровь их на них.
LEV|21|1|И сказал Господь Моисею: объяви священникам, сынам Аароновым, и скажи им: да не оскверняют себя [прикосновением] к умершему из народа своего;
LEV|21|2|только к ближнему родственнику своему, к матери своей и к отцу своему, к сыну своему и дочери своей, к брату своему
LEV|21|3|и к сестре своей, девице, живущей при нем и не бывшей замужем, можно ему [прикасаться], не оскверняя себя;
LEV|21|4|и [прикосновением] к кому бы то ни было в народе своем не должен он осквернять себя, чтобы не сделаться нечистым.
LEV|21|5|Они не должны брить головы своей и подстригать края бороды своей и делать нарезы на теле своем.
LEV|21|6|Они должны быть святы Богу своему и не должны бесчестить имени Бога своего, ибо они приносят жертвы Господу, хлеб Богу своему, и потому должны быть святы.
LEV|21|7|Они не должны брать за себя блудницу и опороченную, не должны брать и жену, отверженную мужем своим, ибо они святы Богу своему.
LEV|21|8|Святи его, ибо он приносит хлеб Богу твоему: да будет он у тебя свят, ибо свят Я Господь, освящающий вас.
LEV|21|9|Если дочь священника осквернит себя блудодеянием, то она бесчестит отца своего; огнем должно сжечь ее.
LEV|21|10|Великий же священник из братьев своих, на голову которого возлит елей помазания, и который освящен, чтобы облачаться в [священные] одежды, не должен обнажать головы своей и раздирать одежд своих;
LEV|21|11|и ни к какому умершему не должен он приступать: даже [прикосновением к умершему] отцу своему и матери своей он не должен осквернять себя.
LEV|21|12|И от святилища он не должен отходить и бесчестить святилище Бога своего, ибо освящение елеем помазания Бога его на нем. Я Господь.
LEV|21|13|В жену он должен брать девицу.
LEV|21|14|вдову, или отверженную, или опороченную, [или] блудницу, не должен он брать, но девицу из народа своего должен он брать в жену;
LEV|21|15|он не должен порочить семени своего в народе своем, ибо Я Господь, освящающий его.
LEV|21|16|И сказал Господь Моисею, говоря:
LEV|21|17|скажи Аарону: никто из семени твоего во [все] роды их, у которого [на теле] будет недостаток, не должен приступать, чтобы приносить хлеб Богу своему;
LEV|21|18|никто, у кого на теле есть недостаток, не должен приступать, ни слепой, ни хромой, ни уродливый,
LEV|21|19|ни такой, у которого переломлена нога или переломлена рука,
LEV|21|20|ни горбатый, ни с сухим членом, ни с бельмом на глазу, ни коростовый, ни паршивый, ни с поврежденными ятрами;
LEV|21|21|ни один человек из семени Аарона священника, у которого [на] [теле] есть недостаток, не должен приступать, чтобы приносить жертвы Господу; недостаток [на нем], поэтому не должен он приступать, чтобы приносить хлеб Богу своему;
LEV|21|22|хлеб Бога своего из великих святынь и из святынь он может есть;
LEV|21|23|но к завесе не должен он приходить и к жертвеннику не должен приступать, потому что недостаток на нем: не должен он бесчестить святилища Моего, ибо Я Господь, освящающий их.
LEV|21|24|И объявил [это] Моисей Аарону и сынам его и всем сынам Израилевым.
LEV|22|1|И сказал Господь Моисею, говоря:
LEV|22|2|скажи Аарону и сынам его, чтоб они осторожно поступали со святынями сынов Израилевых и не бесчестили святаго имени Моего в том, что они посвящают Мне. Я Господь.
LEV|22|3|Скажи им: если кто из всего потомства вашего в роды ваши, имея на себе нечистоту, приступит к святыням, которые посвящают сыны Израилевы Господу, то истребится душа та от лица Моего. Я Господь.
LEV|22|4|Кто из семени Ааронова прокажен, или имеет истечение, тот не должен есть святынь, пока не очистится; и кто прикоснется к чему–нибудь нечистому от мертвого, или у кого случится излияние семени,
LEV|22|5|или кто прикоснется к какому–нибудь гаду, от которого он сделается нечист, или к человеку, от которого он сделается нечист какою бы то ни было нечистотою, –
LEV|22|6|тот, прикоснувшийся к сему, нечист будет до вечера и не должен есть святынь, прежде нежели омоет тело свое водою;
LEV|22|7|но когда зайдет солнце и он очистится, тогда может он есть святыни, ибо это его пища.
LEV|22|8|Мертвечины и звероядины он не должен есть, чтобы не оскверниться этим. Я Господь.
LEV|22|9|Да соблюдают они повеления Мои, чтобы не понести на себе греха и не умереть в нем, когда нарушат сие. Я Господь, освящающий их.
LEV|22|10|Никто посторонний не должен есть святыни; поселившийся у священника и наемник не должен есть святыни;
LEV|22|11|если же священник купит себе человека за серебро, то сей может есть оную; также и домочадцы его могут есть хлеб его.
LEV|22|12|Если дочь священника выйдет в замужество за постороннего, то она не должна есть приносимых святынь;
LEV|22|13|когда же дочь священника будет вдова, или разведенная, и детей нет у нее, и возвратится в дом отца своего, как [была] в юности своей, тогда она может есть хлеб отца своего; а посторонний никто не должен есть его.
LEV|22|14|Кто по ошибке съест [что–нибудь] из святыни, тот должен отдать священнику святыню и приложить к ней пятую ее долю.
LEV|22|15|[Священники] сами не должны порочить святыни сынов Израилевых, которые они приносят Господу,
LEV|22|16|и не должны навлекать на себя вину в преступлении, когда будут есть святыни свои, ибо Я Господь, освящающий их.
LEV|22|17|И сказал Господь Моисею, говоря:
LEV|22|18|объяви Аарону и сынам его и всем сынам Израилевым и скажи им: если кто из дома Израилева, или из пришельцев, [поселившихся] между Израильтянами, по обету ли какому, или по усердию приносит жертву свою, которую приносят Господу во всесожжение,
LEV|22|19|то, чтобы сим приобрести благоволение [от Бога, жертва] [должна быть] без порока, мужеского пола, из крупного скота, из овец и из коз;
LEV|22|20|никакого [животного], на котором есть порок, не приносите; ибо это не приобретет вам благоволения.
LEV|22|21|И если кто приносит мирную жертву Господу, исполняя обет, или по усердию, из крупного скота или из мелкого, то [жертва должна быть] без порока, чтоб быть угодною [Богу]: никакого порока не должно быть на ней;
LEV|22|22|[животного] слепого, или поврежденного, или уродливого, или больного, или коростового, или паршивого, таких не приносите Господу и в жертву не давайте их на жертвенник Господень;
LEV|22|23|тельца и агнца с членами, несоразмерно длинными или короткими, в жертву усердия принести можешь; а если по обету, то это не угодно будет [Богу];
LEV|22|24|[животного], у которого ятра раздавлены, разбиты, оторваны или вырезаны, не приносите Господу и в земле вашей не делайте [сего];
LEV|22|25|и из рук иноземцев не приносите всех таковых [животных] в дар Богу вашему, потому что на них повреждение, порок на них: не приобретут они вам благоволения.
LEV|22|26|И сказал Господь Моисею, говоря:
LEV|22|27|когда родится теленок, или ягненок, или козленок, то семь дней он должен пробыть при матери своей, а от восьмого дня и далее будет благоугоден для приношения в жертву Господу;
LEV|22|28|но ни коровы, ни овцы не заколайте в один день с порождением ее.
LEV|22|29|Если приносите Господу жертву благодарения, то приносите ее так, чтоб она приобрела вам благоволение;
LEV|22|30|в тот же день должно съесть ее, не оставляйте от нее до утра. Я Господь.
LEV|22|31|И соблюдайте заповеди Мои и исполняйте их. Я Господь.
LEV|22|32|Не бесчестите святого имени Моего, чтоб Я был святим среди сынов Израилевых. Я Господь, освящающий вас,
LEV|22|33|Который вывел вас из земли Египетской, чтоб быть вашим Богом. Я Господь.
LEV|23|1|И сказал Господь Моисею, говоря:
LEV|23|2|объяви сынам Израилевым и скажи им о праздниках Господних, в которые должно созывать священные собрания. Вот праздники Мои:
LEV|23|3|шесть дней можно делать дела, а в седьмой день суббота покоя, священное собрание; никакого дела не делайте; это суббота Господня во всех жилищах ваших.
LEV|23|4|Вот праздники Господни, священные собрания, которые вы должны созывать в свое время:
LEV|23|5|в первый месяц, в четырнадцатый [день] месяца вечером Пасха Господня;
LEV|23|6|и в пятнадцатый день того же месяца праздник опресноков Господу; семь дней ешьте опресноки;
LEV|23|7|в первый день да будет у вас священное собрание; никакой работы не работайте;
LEV|23|8|и в течение семи дней приносите жертвы Господу; в седьмой день также священное собрание; никакой работы не работайте.
LEV|23|9|И сказал Господь Моисею, говоря:
LEV|23|10|объяви сынам Израилевым и скажи им: когда придете в землю, которую Я даю вам, и будете жать на ней жатву, то принесите первый сноп жатвы вашей к священнику;
LEV|23|11|он вознесет этот сноп пред Господом, чтобы вам приобрести благоволение; на другой день праздника вознесет его священник;
LEV|23|12|и в день возношения снопа принесите во всесожжение Господу агнца однолетнего, без порока,
LEV|23|13|и с ним хлебного приношения две десятых части [ефы] пшеничной муки, смешанной с елеем, в жертву Господу, в приятное благоухание, и возлияния к нему четверть гина вина;
LEV|23|14|никакого [нового] хлеба, ни сушеных зерен, ни зерен сырых не ешьте до того дня, в который принесете приношения Богу вашему: это вечное постановление в роды ваши во всех жилищах ваших.
LEV|23|15|Отсчитайте себе от первого дня после праздника, от того дня, в который приносите сноп потрясания, семь полных недель,
LEV|23|16|до первого дня после седьмой недели отсчитайте пятьдесят дней, [и] [тогда] принесите новое хлебное приношение Господу:
LEV|23|17|от жилищ ваших приносите два хлеба возношения, которые должны состоять из двух десятых частей [ефы] пшеничной муки и должны быть испечены кислые, [как] первый плод Господу;
LEV|23|18|вместе с хлебами представьте семь агнцев без порока, однолетних, и из крупного скота одного тельца и двух овнов; да будет это во всесожжение Господу, и хлебное приношение и возлияние к ним, в жертву, в приятное благоухание Господу.
LEV|23|19|Приготовьте также из [стада] коз одного козла в жертву за грех и двух однолетних агнцев в жертву мирную.
LEV|23|20|священник должен принести это, потрясая пред Господом, вместе с потрясаемыми хлебами первого плода и с двумя агнцами, и это будет святынею Господу; священнику, [который приносит, это принадлежит];
LEV|23|21|и созывайте [народ] в сей день, священное собрание да будет у вас, никакой работы не работайте: это постановление вечное во всех жилищах ваших в роды ваши.
LEV|23|22|Когда будете жать жатву на земле вашей, не дожинай до края поля твоего, когда жнешь, и оставшегося от жатвы твоей не подбирай; бедному и пришельцу оставь это. Я Господь, Бог ваш.
LEV|23|23|И сказал Господь Моисею, говоря:
LEV|23|24|скажи сынам Израилевым: в седьмой месяц, в первый [день] месяца да будет у вас покой, праздник труб, священное собрание.
LEV|23|25|никакой работы не работайте и приносите жертву Господу.
LEV|23|26|И сказал Господь Моисею, говоря:
LEV|23|27|также в девятый [день] седьмого месяца сего, день очищения, да будет у вас священное собрание; смиряйте души ваши и приносите жертву Господу;
LEV|23|28|никакого дела не делайте в день сей, ибо это день очищения, дабы очистить вас пред лицем Господа, Бога вашего;
LEV|23|29|а всякая душа, которая не смирит себя в этот день, истребится из народа своего;
LEV|23|30|и если какая душа будет делать какое–нибудь дело в день сей, Я истреблю ту душу из народа ее;
LEV|23|31|никакого дела не делайте: это постановление вечное в роды ваши, во всех жилищах ваших;
LEV|23|32|это для вас суббота покоя, и смиряйте души ваши, с вечера девятого [дня] месяца; от вечера до вечера празднуйте субботу вашу.
LEV|23|33|И сказал Господь Моисею, говоря:
LEV|23|34|скажи сынам Израилевым: с пятнадцатого дня того же седьмого месяца праздник кущей, семь дней Господу;
LEV|23|35|в первый день священное собрание, никакой работы не работайте;
LEV|23|36|в [течение] семи дней приносите жертву Господу; в восьмой день священное собрание да будет у вас, и приносите жертву Господу: это отдание праздника, никакой работы не работайте.
LEV|23|37|Вот праздники Господни, в которые должно созывать священные собрания, чтобы приносить в жертву Господу всесожжение, хлебное приношение, заколаемые жертвы и возлияния, каждое в свой день,
LEV|23|38|кроме суббот Господних и кроме даров ваших, и кроме всех обетов ваших и кроме всего [приносимого] по усердию вашему, что вы даете Господу.
LEV|23|39|А в пятнадцатый день седьмого месяца, когда вы собираете произведения земли, празднуйте праздник Господень семь дней: в первый день покой и в восьмой день покой;
LEV|23|40|в первый день возьмите себе ветви красивых дерев, ветви пальмовые и ветви дерев широколиственных и верб речных, и веселитесь пред Господом Богом вашим семь дней;
LEV|23|41|и празднуйте этот праздник Господень семь дней в году: это постановление вечное в роды ваши; в седьмой месяц празднуйте его;
LEV|23|42|в кущах живите семь дней; всякий туземец Израильтянин должен жить в кущах,
LEV|23|43|чтобы знали роды ваши, что в кущах поселил Я сынов Израилевых, когда вывел их из земли Египетской. Я Господь, Бог ваш.
LEV|23|44|И объявил Моисей сынам Израилевым о праздниках Господних.
LEV|24|1|И сказал Господь Моисею, говоря:
LEV|24|2|прикажи сынам Израилевым, чтоб они принесли тебе елея чистого, выбитого, для освещения, чтобы непрестанно горел светильник;
LEV|24|3|вне завесы [ковчега] откровения в скинии собрания Аарон [и сыны его] должны ставить оный пред Господом от вечера до утра всегда: это вечное постановление в роды ваши;
LEV|24|4|на подсвечнике чистом должны они ставить светильник пред Господом всегда.
LEV|24|5|И возьми пшеничной муки и испеки из нее двенадцать хлебов; в каждом хлебе должны быть две десятых [ефы];
LEV|24|6|и положи их в два ряда, по шести в ряд, на чистом столе пред Господом;
LEV|24|7|и положи на [каждый] ряд чистого ливана, и будет это при хлебе, в память, в жертву Господу;
LEV|24|8|в каждый день субботы постоянно должно полагать их пред Господом от сынов Израилевых: это завет вечный;
LEV|24|9|они будут принадлежать Аарону и сынам его, которые будут есть их на святом месте, ибо это великая святыня для них из жертв Господних: [это] постановление вечное.
LEV|24|10|И вышел сын одной Израильтянки, родившейся от Египтянина, к сынам Израилевым, и поссорился в стане сын Израильтянки с Израильтянином;
LEV|24|11|хулил сын Израильтянки имя [Господне] и злословил. И привели его к Моисею;
LEV|24|12|и посадили его под стражу, доколе не будет объявлена им воля Господня.
LEV|24|13|И сказал Господь Моисею, говоря:
LEV|24|14|выведи злословившего вон из стана, и все слышавшие пусть положат руки свои на голову его, и все общество побьет его камнями;
LEV|24|15|и сынам Израилевым скажи: кто будет злословить Бога своего, тот понесет грех свой;
LEV|24|16|и хулитель имени Господня должен умереть, камнями побьет его все общество: пришлец ли, туземец ли станет хулить имя [Господне], предан будет смерти.
LEV|24|17|Кто убьет какого–либо человека, тот предан будет смерти.
LEV|24|18|Кто убьет скотину, должен заплатить за нее, скотину за скотину.
LEV|24|19|Кто сделает повреждение на теле ближнего своего, тому должно сделать то же, что он сделал:
LEV|24|20|перелом за перелом, око за око, зуб за зуб; как он сделал повреждение на [теле] человека, так и ему должно сделать.
LEV|24|21|Кто убьет скотину, должен заплатить за нее; а кто убьет человека, того должно предать смерти.
LEV|24|22|Один суд должен быть у вас, как для пришельца, так и для туземца; ибо Я Господь, Бог ваш.
LEV|24|23|И сказал Моисей сынам Израилевым; и вывели злословившего вон из стана, и побили его камнями, и сделали сыны Израилевы, как повелел Господь Моисею.
LEV|25|1|И сказал Господь Моисею на горе Синае, говоря:
LEV|25|2|объяви сынам Израилевым и скажи им: когда придете в землю, которую Я даю вам, тогда земля должна покоиться в субботу Господню;
LEV|25|3|шесть лет засевай поле твое и шесть лет обрезывай виноградник твой, и собирай произведения их,
LEV|25|4|а в седьмой год да будет суббота покоя земли, суббота Господня: поля твоего не засевай и виноградника твоего не обрезывай;
LEV|25|5|что само вырастет на жатве твоей, не сжинай, и гроздов с необрезанных лоз твоих не снимай; да будет это год покоя земли;
LEV|25|6|и будет это в продолжение субботы земли [всем] вам в пищу, тебе и рабу твоему, и рабе твоей, и наемнику твоему, и поселенцу твоему, поселившемуся у тебя;
LEV|25|7|и скоту твоему и зверям, которые на земле твоей, да будут все произведения ее в пищу.
LEV|25|8|И насчитай себе семь субботних лет, семь раз по семи лет, чтоб было у тебя в семи субботних годах сорок девять лет;
LEV|25|9|и воструби трубою в седьмой месяц, в десятый [день] месяца, в день очищения вострубите трубою по всей земле вашей;
LEV|25|10|и освятите пятидесятый год и объявите свободу на земле всем жителям ее: да будет это у вас юбилей; и возвратитесь каждый во владение свое, и каждый возвратитесь в свое племя.
LEV|25|11|Пятидесятый год да будет у вас юбилей: не сейте и не жните, что само вырастет на земле, и не снимайте ягод с необрезанных [лоз] ее,
LEV|25|12|ибо это юбилей: священным да будет он для вас; с поля ешьте произведения ее.
LEV|25|13|В юбилейный год возвратитесь каждый во владение свое.
LEV|25|14|Если будешь продавать что ближнему твоему, или будешь покупать что у ближнего твоего, не обижайте друг друга;
LEV|25|15|по расчислению лет после юбилея ты должен покупать у ближнего твоего, и по расчислению лет дохода он должен продавать тебе;
LEV|25|16|если много [остается] лет, умножь цену; а если мало лет [остается], уменьши цену, ибо известное число [лет] жатв он продает тебе.
LEV|25|17|Не обижайте один другого; бойся Бога твоего, ибо Я Господь, Бог ваш.
LEV|25|18|Исполняйте постановления Мои, и храните законы Мои и исполняйте их, и будете жить спокойно на земле;
LEV|25|19|и будет земля давать плод свой, и будете есть досыта, и будете жить спокойно на ней.
LEV|25|20|Если скажете: что же нам есть в седьмой год, когда мы не будем ни сеять, ни собирать произведений наших?
LEV|25|21|Я пошлю благословение Мое на вас в шестой год, и он принесет произведений на три года;
LEV|25|22|и будете сеять в восьмой год, но есть будете произведения старые до девятого года; доколе не поспеют произведения его, будете есть старое.
LEV|25|23|Землю не должно продавать навсегда, ибо Моя земля: вы пришельцы и поселенцы у Меня;
LEV|25|24|по всей земле владения вашего дозволяйте выкуп земли.
LEV|25|25|Если брат твой обеднеет и продаст от владения своего, то придет близкий его родственник и выкупит проданное братом его;
LEV|25|26|если же некому за него выкупить, но сам он будет иметь достаток и найдет, сколько нужно на выкуп,
LEV|25|27|то пусть он расчислит годы продажи своей и возвратит остальное тому, кому он продал, и вступит опять во владение свое;
LEV|25|28|если же не найдет рука его, сколько нужно возвратить ему, то проданное им останется в руках покупщика до юбилейного года, а в юбилейный год отойдет оно, и он опять вступит во владение свое.
LEV|25|29|Если кто продаст жилой дом в городе, [огражденном] стеною, то выкупить его можно до истечения года от продажи его: в течение года выкупить его можно;
LEV|25|30|если же не будет он выкуплен до истечения целого года, то дом, который в городе, имеющем стену, останется навсегда у купившего его в роды его, и в юбилей не отойдет [от него].
LEV|25|31|А домы в селениях, вокруг которых нет стены, должно считать наравне с полем земли: выкупать их можно, и в юбилей они отходят.
LEV|25|32|А города левитов, домы в городах владения их, левитам всегда можно выкупать;
LEV|25|33|а кто из левитов не выкупит, то проданный дом в городе владения их в юбилей отойдет, потому что домы в городах левитских составляют их владение среди сынов Израилевых;
LEV|25|34|и полей вокруг городов их продавать нельзя, потому что это вечное владение их.
LEV|25|35|Если брат твой обеднеет и придет в упадок у тебя, то поддержи его, пришлец ли он, или поселенец, чтоб он жил с тобою;
LEV|25|36|не бери от него роста и прибыли и бойся Бога твоего; чтоб жил брат твой с тобою;
LEV|25|37|серебра твоего не отдавай ему в рост и хлеба твоего не отдавай ему для [получения] прибыли.
LEV|25|38|Я Господь, Бог ваш, Который вывел вас из земли Египетской, чтобы дать вам землю Ханаанскую, чтоб быть вашим Богом.
LEV|25|39|Когда обеднеет у тебя брат твой и продан будет тебе, то не налагай на него работы рабской:
LEV|25|40|он должен быть у тебя как наемник, как поселенец; до юбилейного года пусть работает у тебя,
LEV|25|41|а [тогда] пусть отойдет он от тебя, сам и дети его с ним, и возвратится в племя свое, и вступит опять во владение отцов своих,
LEV|25|42|потому что они – Мои рабы, которых Я вывел из земли Египетской: не должно продавать их, как продают рабов;
LEV|25|43|не господствуй над ним с жестокостью и бойся Бога твоего.
LEV|25|44|А чтобы раб твой и рабыня твоя были у тебя, то покупайте себе раба и рабыню у народов, которые вокруг вас;
LEV|25|45|также и из детей поселенцев, поселившихся у вас, можете покупать, и из племени их, которое у вас, которое у них родилось в земле вашей, и они могут быть вашей собственностью;
LEV|25|46|можете передавать их в наследство и сынам вашим по себе, как имение; вечно владейте ими, как рабами. А над братьями вашими, сынами Израилевыми, друг над другом, не господствуйте с жестокостью.
LEV|25|47|Если пришлец или поселенец твой будет иметь достаток, а брат твой пред ним обеднеет и продастся пришельцу, поселившемуся у тебя, или кому–нибудь из племени пришельца,
LEV|25|48|то после продажи можно выкупить его; кто–нибудь из братьев его должен выкупить его,
LEV|25|49|или дядя его, или сын дяди его должен выкупить его, или кто–нибудь из родства его, из племени его, должен выкупить его; или если будет иметь достаток, сам выкупится.
LEV|25|50|И он должен рассчитаться с купившим его, [начиная] от того года, когда он продал себя, до года юбилейного, и серебро, за которое он продал себя, должно отдать ему по числу лет; как временный наемник он должен быть у него;
LEV|25|51|и если еще много [остается] лет, то по мере их он должен отдать в выкуп за себя серебро, за которое он куплен;
LEV|25|52|если же мало остается лет до юбилейного года, то он должен сосчитать и по мере лет отдать за себя выкуп.
LEV|25|53|Он должен быть у него, как наемник, во все годы; он не должен господствовать над ним с жестокостью в глазах твоих.
LEV|25|54|Если же он не выкупится таким образом, то в юбилейный год отойдет сам и дети его с ним,
LEV|25|55|потому что сыны Израилевы Мои рабы; они Мои рабы, которых Я вывел из земли Египетской. Я Господь, Бог ваш.
LEV|26|1|Не делайте себе кумиров и изваяний, и столбов не ставьте у себя, и камней с изображениями не кладите в земле вашей, чтобы кланяться пред ними, ибо Я Господь Бог ваш.
LEV|26|2|Субботы Мои соблюдайте и святилище Мое чтите: Я Господь.
LEV|26|3|Если вы будете поступать по уставам Моим и заповеди Мои будете хранить и исполнять их,
LEV|26|4|то Я дам вам дожди в свое время, и земля даст произрастения свои, и дерева полевые дадут плод свой;
LEV|26|5|и молотьба [хлеба] будет достигать у вас собирания винограда, собирание винограда будет достигать посева, и будете есть хлеб свой досыта, и будете жить на земле [вашей] безопасно;
LEV|26|6|пошлю мир на землю [вашу], ляжете, и никто вас не обеспокоит, сгоню лютых зверей с земли [вашей], и меч не пройдет по земле вашей;
LEV|26|7|и будете прогонять врагов ваших, и падут они пред вами от меча;
LEV|26|8|пятеро из вас прогонят сто, и сто из вас прогонят тьму, и падут враги ваши пред вами от меча;
LEV|26|9|призрю на вас, и плодородными сделаю вас, и размножу вас, и буду тверд в завете Моем с вами;
LEV|26|10|и будете есть старое прошлогоднее, и выбросите старое ради нового;
LEV|26|11|и поставлю жилище Мое среди вас, и душа Моя не возгнушается вами;
LEV|26|12|и буду ходить среди вас и буду вашим Богом, а вы будете Моим народом.
LEV|26|13|Я Господь Бог ваш, Который вывел вас из земли Египетской, чтоб вы не были там рабами, и сокрушил узы ярма вашего, и повел вас с поднятою головою.
LEV|26|14|Если же не послушаете Меня и не будете исполнять всех заповедей сих,
LEV|26|15|и если презрите Мои постановления, и если душа ваша возгнушается Моими законами, так что вы не будете исполнять всех заповедей Моих, нарушив завет Мой, –
LEV|26|16|то и Я поступлю с вами так: пошлю на вас ужас, чахлость и горячку, от которых истомятся глаза и измучится душа, и будете сеять семена ваши напрасно, и враги ваши съедят их;
LEV|26|17|обращу лице Мое на вас, и падете пред врагами вашими, и будут господствовать над вами неприятели ваши, и побежите, когда никто не гонится за вами.
LEV|26|18|Если и при всем том не послушаете Меня, то Я всемеро увеличу наказание за грехи ваши,
LEV|26|19|и сломлю гордое упорство ваше, и небо ваше сделаю, как железо, и землю вашу, как медь;
LEV|26|20|и напрасно будет истощаться сила ваша, и земля ваша не даст произрастений своих, и дерева земли не дадут плодов своих.
LEV|26|21|Если же [после сего] пойдете против Меня и не захотите слушать Меня, то Я прибавлю вам ударов всемеро за грехи ваши:
LEV|26|22|пошлю на вас зверей полевых, которые лишат вас детей, истребят скот ваш и вас уменьшат, так что опустеют дороги ваши.
LEV|26|23|Если и после сего не исправитесь и пойдете против Меня,
LEV|26|24|то и Я пойду против вас и поражу вас всемеро за грехи ваши,
LEV|26|25|и наведу на вас мстительный меч в отмщение за завет; если же вы укроетесь в города ваши, то пошлю на вас язву, и преданы будете в руки врага;
LEV|26|26|хлеб, подкрепляющий [человека], истреблю у вас; десять женщин будут печь хлеб ваш в одной печи и будут отдавать хлеб ваш весом; вы будете есть и не будете сыты.
LEV|26|27|Если же и после сего не послушаете Меня и пойдете против Меня,
LEV|26|28|то и Я в ярости пойду против вас и накажу вас всемеро за грехи ваши,
LEV|26|29|и будете есть плоть сынов ваших, и плоть дочерей ваших будете есть;
LEV|26|30|разорю высоты ваши и разрушу столбы ваши, и повергну трупы ваши на обломки идолов ваших, и возгнушается душа Моя вами;
LEV|26|31|города ваши сделаю пустынею, и опустошу святилища ваши, и не буду обонять приятного благоухания [жертв] ваших;
LEV|26|32|опустошу землю [вашу], так что изумятся о ней враги ваши, поселившиеся на ней;
LEV|26|33|а вас рассею между народами и обнажу вслед вас меч, и будет земля ваша пуста и города ваши разрушены.
LEV|26|34|Тогда удовлетворит себя земля за субботы свои во все дни запустения [своего]; когда вы будете в земле врагов ваших, тогда будет покоиться земля и удовлетворит себя за субботы свои;
LEV|26|35|во все дни запустения [своего] будет она покоиться, сколько ни покоилась в субботы ваши, когда вы жили на ней.
LEV|26|36|Оставшимся из вас пошлю в сердца робость в земле врагов их, и шум колеблющегося листа погонит их, и побегут, как от меча, и падут, когда никто не преследует,
LEV|26|37|и споткнутся друг на друга, как от меча, между тем как никто не преследует, и не будет у вас силы противостоять врагам вашим;
LEV|26|38|и погибнете между народами, и пожрет вас земля врагов ваших;
LEV|26|39|а оставшиеся из вас исчахнут за свои беззакония в землях врагов ваших и за беззакония отцов своих исчахнут;
LEV|26|40|тогда признаются они в беззаконии своем и в беззаконии отцов своих, как они совершали преступления против Меня и шли против Меня,
LEV|26|41|[за что] и Я шел против них и ввел их в землю врагов их; тогда покорится необрезанное сердце их, и тогда потерпят они за беззакония свои.
LEV|26|42|И Я вспомню завет Мой с Иаковом и завет Мой с Исааком, и завет Мой с Авраамом вспомню, и землю вспомню;
LEV|26|43|тогда как земля оставлена будет ими и будет удовлетворять себя за субботы свои, опустев от них, и они будут терпеть за свое беззаконие, за то, что презирали законы Мои и душа их гнушалась постановлениями Моими,
LEV|26|44|и тогда как они будут в земле врагов их, – Я не презрю их и не возгнушаюсь ими до того, чтоб истребить их, чтоб разрушить завет Мой с ними, ибо Я Господь, Бог их;
LEV|26|45|вспомню для них завет с предками, которых вывел Я из земли Египетской пред глазами народов, чтоб быть их Богом. Я Господь.
LEV|26|46|Вот постановления и определения и законы, которые постановил Господь между Собою и между сынами Израилевыми на горе Синае, чрез Моисея.
LEV|27|1|И сказал Господь Моисею, говоря:
LEV|27|2|объяви сынам Израилевым и скажи им: если кто дает обет посвятить душу Господу по оценке твоей,
LEV|27|3|то оценка твоя мужчине от двадцати лет до шестидесяти должна быть пятьдесят сиклей серебряных, по сиклю священному;
LEV|27|4|если же это женщина, то оценка твоя должна быть тридцать сиклей;
LEV|27|5|от пяти лет до двадцати оценка твоя мужчине должна быть двадцать сиклей, а женщине десять сиклей;
LEV|27|6|а от месяца до пяти лет оценка твоя мужчине должна быть пять сиклей серебра, а женщине оценка твоя три сикля серебра;
LEV|27|7|от шестидесяти лет и выше мужчине оценка твоя должна быть пятнадцать сиклей серебра, а женщине десять сиклей.
LEV|27|8|Если же он беден и не в силах [отдать] по оценке твоей, то пусть представят его священнику, и священник пусть оценит его: соразмерно с состоянием давшего обет пусть оценит его священник.
LEV|27|9|Если же то будет скот, который приносят в жертву Господу, то все, что дано Господу, должно быть свято:
LEV|27|10|не должно выменивать его и заменять хорошее худым, или худое хорошим; если же станет кто заменять скотину скотиною, то и она и замен ее будет святынею.
LEV|27|11|Если же то будет какая–нибудь скотина нечистая, которую не приносят в жертву Господу, то должно представить скотину священнику,
LEV|27|12|и священник оценит ее, хороша ли она, или худа, и как оценит священник, так и должно быть;
LEV|27|13|если же кто хочет выкупить ее, то пусть прибавит пятую долю к оценке твоей.
LEV|27|14|Если кто посвящает дом свой в святыню Господу, то священник должен оценить его, хорош ли он, или худ, и как оценит его священник, так и состоится;
LEV|27|15|если же посвятивший захочет выкупить дом свой, то пусть прибавит пятую часть серебра оценки твоей, и [тогда] будет его.
LEV|27|16|Если поле из своего владения посвятит кто Господу, то оценка твоя должна быть по мере посева: за посев хомера ячменя пятьдесят сиклей серебра;
LEV|27|17|если от юбилейного года посвящает кто поле свое, – должно состояться по оценке твоей;
LEV|27|18|если же после юбилея посвящает кто поле свое, то священник должен рассчитать серебро по мере лет, оставшихся до юбилейного года, и должно убавить из оценки твоей;
LEV|27|19|если же захочет выкупить поле посвятивший его, то пусть он прибавит пятую часть серебра оценки твоей, и оно останется за ним;
LEV|27|20|если же он не выкупит поля, и будет продано поле другому человеку, то уже нельзя выкупить:
LEV|27|21|поле то, когда оно в юбилей отойдет, будет святынею Господу, как бы поле заклятое; священнику достанется оно во владение.
LEV|27|22|А если кто посвятит Господу поле купленное, которое не из полей его владения,
LEV|27|23|то священник должен рассчитать ему количество оценки до юбилейного года, и должен он отдать по расчету в тот же день, [как] святыню Господню;
LEV|27|24|поле же в юбилейный год перейдет опять к тому, у кого куплено, кому принадлежит владение той земли.
LEV|27|25|Всякая оценка твоя должна быть по сиклю священному, двадцать гер должно быть в сикле.
LEV|27|26|Только первенцев из скота, которые по первенству принадлежат Господу, не должен никто посвящать: вол ли то, или мелкий скот, – Господни они.
LEV|27|27|Если же скот нечистый, то должно выкупить по оценке твоей и приложить к тому пятую часть; если не выкупят, то должно продать по оценке твоей.
LEV|27|28|Только все заклятое, что под заклятием отдает человек Господу из своей собственности, – человека ли, скотину ли, поле ли своего владения, – не продается и не выкупается: все заклятое есть великая святыня Господня;
LEV|27|29|все заклятое, что заклято от людей, не выкупается: оно должно быть предано смерти.
LEV|27|30|И всякая десятина на земле из семян земли и из плодов дерева принадлежит Господу: это святыня Господня;
LEV|27|31|если же кто захочет выкупить десятину свою, то пусть приложит к [цене] ее пятую долю.
LEV|27|32|И всякую десятину из крупного и мелкого скота, из всего, что проходит под жезлом десятое, должно посвящать Господу;
LEV|27|33|не должно разбирать, хорошее ли то, или худое, и не должно заменять его; если же кто заменит его, то и само оно и замен его будет святынею и не может быть выкуплено.
LEV|27|34|Вот заповеди, которые заповедал Господь Моисею для сынов Израилевых на горе Синае.
