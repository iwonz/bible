DEUT|1|1|These be the words which Moses spake unto all Israel on this side Jordan in the wilderness, in the plain over against the Red sea, between Paran, and Tophel, and Laban, and Hazeroth, and Dizahab.
DEUT|1|2|(There are eleven days' journey from Horeb by the way of mount Seir unto Kadeshbarnea.)
DEUT|1|3|And it came to pass in the fortieth year, in the eleventh month, on the first day of the month, that Moses spake unto the children of Israel, according unto all that the LORD had given him in commandment unto them;
DEUT|1|4|After he had slain Sihon the king of the Amorites, which dwelt in Heshbon, and Og the king of Bashan, which dwelt at Astaroth in Edrei:
DEUT|1|5|On this side Jordan, in the land of Moab, began Moses to declare this law, saying,
DEUT|1|6|The LORD our God spake unto us in Horeb, saying, Ye have dwelt long enough in this mount:
DEUT|1|7|Turn you, and take your journey, and go to the mount of the Amorites, and unto all the places nigh thereunto, in the plain, in the hills, and in the vale, and in the south, and by the sea side, to the land of the Canaanites, and unto Lebanon, unto the great river, the river Euphrates.
DEUT|1|8|Behold, I have set the land before you: go in and possess the land which the LORD sware unto your fathers, Abraham, Isaac, and Jacob, to give unto them and to their seed after them.
DEUT|1|9|And I spake unto you at that time, saying, I am not able to bear you myself alone:
DEUT|1|10|The LORD your God hath multiplied you, and, behold, ye are this day as the stars of heaven for multitude.
DEUT|1|11|(The LORD God of your fathers make you a thousand times so many more as ye are, and bless you, as he hath promised you!)
DEUT|1|12|How can I myself alone bear your cumbrance, and your burden, and your strife?
DEUT|1|13|Take you wise men, and understanding, and known among your tribes, and I will make them rulers over you.
DEUT|1|14|And ye answered me, and said, The thing which thou hast spoken is good for us to do.
DEUT|1|15|So I took the chief of your tribes, wise men, and known, and made them heads over you, captains over thousands, and captains over hundreds, and captains over fifties, and captains over tens, and officers among your tribes.
DEUT|1|16|And I charged your judges at that time, saying, Hear the causes between your brethren, and judge righteously between every man and his brother, and the stranger that is with him.
DEUT|1|17|Ye shall not respect persons in judgment; but ye shall hear the small as well as the great; ye shall not be afraid of the face of man; for the judgment is God's: and the cause that is too hard for you, bring it unto me, and I will hear it.
DEUT|1|18|And I commanded you at that time all the things which ye should do.
DEUT|1|19|And when we departed from Horeb, we went through all that great and terrible wilderness, which ye saw by the way of the mountain of the Amorites, as the LORD our God commanded us; and we came to Kadeshbarnea.
DEUT|1|20|And I said unto you, Ye are come unto the mountain of the Amorites, which the LORD our God doth give unto us.
DEUT|1|21|Behold, the LORD thy God hath set the land before thee: go up and possess it, as the LORD God of thy fathers hath said unto thee; fear not, neither be discouraged.
DEUT|1|22|And ye came near unto me every one of you, and said, We will send men before us, and they shall search us out the land, and bring us word again by what way we must go up, and into what cities we shall come.
DEUT|1|23|And the saying pleased me well: and I took twelve men of you, one of a tribe:
DEUT|1|24|And they turned and went up into the mountain, and came unto the valley of Eshcol, and searched it out.
DEUT|1|25|And they took of the fruit of the land in their hands, and brought it down unto us, and brought us word again, and said, It is a good land which the LORD our God doth give us.
DEUT|1|26|Notwithstanding ye would not go up, but rebelled against the commandment of the LORD your God:
DEUT|1|27|And ye murmured in your tents, and said, Because the LORD hated us, he hath brought us forth out of the land of Egypt, to deliver us into the hand of the Amorites, to destroy us.
DEUT|1|28|Whither shall we go up? our brethren have discouraged our heart, saying, The people is greater and taller than we; the cities are great and walled up to heaven; and moreover we have seen the sons of the Anakims there.
DEUT|1|29|Then I said unto you, Dread not, neither be afraid of them.
DEUT|1|30|The LORD your God which goeth before you, he shall fight for you, according to all that he did for you in Egypt before your eyes;
DEUT|1|31|And in the wilderness, where thou hast seen how that the LORD thy God bare thee, as a man doth bear his son, in all the way that ye went, until ye came into this place.
DEUT|1|32|Yet in this thing ye did not believe the LORD your God,
DEUT|1|33|Who went in the way before you, to search you out a place to pitch your tents in, in fire by night, to show you by what way ye should go, and in a cloud by day.
DEUT|1|34|And the LORD heard the voice of your words, and was wroth, and sware, saying,
DEUT|1|35|Surely there shall not one of these men of this evil generation see that good land, which I sware to give unto your fathers.
DEUT|1|36|Save Caleb the son of Jephunneh; he shall see it, and to him will I give the land that he hath trodden upon, and to his children, because he hath wholly followed the LORD.
DEUT|1|37|Also the LORD was angry with me for your sakes, saying, Thou also shalt not go in thither.
DEUT|1|38|But Joshua the son of Nun, which standeth before thee, he shall go in thither: encourage him: for he shall cause Israel to inherit it.
DEUT|1|39|Moreover your little ones, which ye said should be a prey, and your children, which in that day had no knowledge between good and evil, they shall go in thither, and unto them will I give it, and they shall possess it.
DEUT|1|40|But as for you, turn you, and take your journey into the wilderness by the way of the Red sea.
DEUT|1|41|Then ye answered and said unto me, We have sinned against the LORD, we will go up and fight, according to all that the LORD our God commanded us. And when ye had girded on every man his weapons of war, ye were ready to go up into the hill.
DEUT|1|42|And the LORD said unto me, Say unto them. Go not up, neither fight; for I am not among you; lest ye be smitten before your enemies.
DEUT|1|43|So I spake unto you; and ye would not hear, but rebelled against the commandment of the LORD, and went presumptuously up into the hill.
DEUT|1|44|And the Amorites, which dwelt in that mountain, came out against you, and chased you, as bees do, and destroyed you in Seir, even unto Hormah.
DEUT|1|45|And ye returned and wept before the LORD; but the LORD would not hearken to your voice, nor give ear unto you.
DEUT|1|46|So ye abode in Kadesh many days, according unto the days that ye abode there.
DEUT|2|1|Then we turned, and took our journey into the wilderness by the way of the Red sea, as the LORD spake unto me: and we compassed mount Seir many days.
DEUT|2|2|And the LORD spake unto me, saying,
DEUT|2|3|Ye have compassed this mountain long enough: turn you northward.
DEUT|2|4|And command thou the people, saying, Ye are to pass through the coast of your brethren the children of Esau, which dwell in Seir; and they shall be afraid of you: take ye good heed unto yourselves therefore:
DEUT|2|5|Meddle not with them; for I will not give you of their land, no, not so much as a foot breadth; because I have given mount Seir unto Esau for a possession.
DEUT|2|6|Ye shall buy meat of them for money, that ye may eat; and ye shall also buy water of them for money, that ye may drink.
DEUT|2|7|For the LORD thy God hath blessed thee in all the works of thy hand: he knoweth thy walking through this great wilderness: these forty years the LORD thy God hath been with thee; thou hast lacked nothing.
DEUT|2|8|And when we passed by from our brethren the children of Esau, which dwelt in Seir, through the way of the plain from Elath, and from Eziongaber, we turned and passed by the way of the wilderness of Moab.
DEUT|2|9|And the LORD said unto me, Distress not the Moabites, neither contend with them in battle: for I will not give thee of their land for a possession; because I have given Ar unto the children of Lot for a possession.
DEUT|2|10|The Emims dwelt therein in times past, a people great, and many, and tall, as the Anakims;
DEUT|2|11|Which also were accounted giants, as the Anakims; but the Moabites called them Emims.
DEUT|2|12|The Horims also dwelt in Seir beforetime; but the children of Esau succeeded them, when they had destroyed them from before them, and dwelt in their stead; as Israel did unto the land of his possession, which the LORD gave unto them.
DEUT|2|13|Now rise up, said I, and get you over the brook Zered. And we went over the brook Zered.
DEUT|2|14|And the space in which we came from Kadeshbarnea, until we were come over the brook Zered, was thirty and eight years; until all the generation of the men of war were wasted out from among the host, as the LORD sware unto them.
DEUT|2|15|For indeed the hand of the LORD was against them, to destroy them from among the host, until they were consumed.
DEUT|2|16|So it came to pass, when all the men of war were consumed and dead from among the people,
DEUT|2|17|That the LORD spake unto me, saying,
DEUT|2|18|Thou art to pass over through Ar, the coast of Moab, this day:
DEUT|2|19|And when thou comest nigh over against the children of Ammon, distress them not, nor meddle with them: for I will not give thee of the land of the children of Ammon any possession; because I have given it unto the children of Lot for a possession.
DEUT|2|20|(That also was accounted a land of giants: giants dwelt therein in old time; and the Ammonites call them Zamzummims;
DEUT|2|21|A people great, and many, and tall, as the Anakims; but the LORD destroyed them before them; and they succeeded them, and dwelt in their stead:
DEUT|2|22|As he did to the children of Esau, which dwelt in Seir, when he destroyed the Horims from before them; and they succeeded them, and dwelt in their stead even unto this day:
DEUT|2|23|And the Avims which dwelt in Hazerim, even unto Azzah, the Caphtorims, which came forth out of Caphtor, destroyed them, and dwelt in their stead.)
DEUT|2|24|Rise ye up, take your journey, and pass over the river Arnon: behold, I have given into thine hand Sihon the Amorite, king of Heshbon, and his land: begin to possess it, and contend with him in battle.
DEUT|2|25|This day will I begin to put the dread of thee and the fear of thee upon the nations that are under the whole heaven, who shall hear report of thee, and shall tremble, and be in anguish because of thee.
DEUT|2|26|And I sent messengers out of the wilderness of Kedemoth unto Sihon king of Heshbon with words of peace, saying,
DEUT|2|27|Let me pass through thy land: I will go along by the high way, I will neither turn unto the right hand nor to the left.
DEUT|2|28|Thou shalt sell me meat for money, that I may eat; and give me water for money, that I may drink: only I will pass through on my feet;
DEUT|2|29|(As the children of Esau which dwell in Seir, and the Moabites which dwell in Ar, did unto me;) until I shall pass over Jordan into the land which the LORD our God giveth us.
DEUT|2|30|But Sihon king of Heshbon would not let us pass by him: for the LORD thy God hardened his spirit, and made his heart obstinate, that he might deliver him into thy hand, as appeareth this day.
DEUT|2|31|And the LORD said unto me, Behold, I have begun to give Sihon and his land before thee: begin to possess, that thou mayest inherit his land.
DEUT|2|32|Then Sihon came out against us, he and all his people, to fight at Jahaz.
DEUT|2|33|And the LORD our God delivered him before us; and we smote him, and his sons, and all his people.
DEUT|2|34|And we took all his cities at that time, and utterly destroyed the men, and the women, and the little ones, of every city, we left none to remain:
DEUT|2|35|Only the cattle we took for a prey unto ourselves, and the spoil of the cities which we took.
DEUT|2|36|From Aroer, which is by the brink of the river of Arnon, and from the city that is by the river, even unto Gilead, there was not one city too strong for us: the LORD our God delivered all unto us:
DEUT|2|37|Only unto the land of the children of Ammon thou camest not, nor unto any place of the river Jabbok, nor unto the cities in the mountains, nor unto whatsoever the LORD our God forbade us.
DEUT|3|1|Then we turned, and went up the way to Bashan: and Og the king of Bashan came out against us, he and all his people, to battle at Edrei.
DEUT|3|2|And the LORD said unto me, Fear him not: for I will deliver him, and all his people, and his land, into thy hand; and thou shalt do unto him as thou didst unto Sihon king of the Amorites, which dwelt at Heshbon.
DEUT|3|3|So the LORD our God delivered into our hands Og also, the king of Bashan, and all his people: and we smote him until none was left to him remaining.
DEUT|3|4|And we took all his cities at that time, there was not a city which we took not from them, threescore cities, all the region of Argob, the kingdom of Og in Bashan.
DEUT|3|5|All these cities were fenced with high walls, gates, and bars; beside unwalled towns a great many.
DEUT|3|6|And we utterly destroyed them, as we did unto Sihon king of Heshbon, utterly destroying the men, women, and children, of every city.
DEUT|3|7|But all the cattle, and the spoil of the cities, we took for a prey to ourselves.
DEUT|3|8|And we took at that time out of the hand of the two kings of the Amorites the land that was on this side Jordan, from the river of Arnon unto mount Hermon;
DEUT|3|9|(Which Hermon the Sidonians call Sirion; and the Amorites call it Shenir;)
DEUT|3|10|All the cities of the plain, and all Gilead, and all Bashan, unto Salchah and Edrei, cities of the kingdom of Og in Bashan.
DEUT|3|11|For only Og king of Bashan remained of the remnant of giants; behold his bedstead was a bedstead of iron; is it not in Rabbath of the children of Ammon? nine cubits was the length thereof, and four cubits the breadth of it, after the cubit of a man.
DEUT|3|12|And this land, which we possessed at that time, from Aroer, which is by the river Arnon, and half mount Gilead, and the cities thereof, gave I unto the Reubenites and to the Gadites.
DEUT|3|13|And the rest of Gilead, and all Bashan, being the kingdom of Og, gave I unto the half tribe of Manasseh; all the region of Argob, with all Bashan, which was called the land of giants.
DEUT|3|14|Jair the son of Manasseh took all the country of Argob unto the coasts of Geshuri and Maachathi; and called them after his own name, Bashanhavothjair, unto this day.
DEUT|3|15|And I gave Gilead unto Machir.
DEUT|3|16|And unto the Reubenites and unto the Gadites I gave from Gilead even unto the river Arnon half the valley, and the border even unto the river Jabbok, which is the border of the children of Ammon;
DEUT|3|17|The plain also, and Jordan, and the coast thereof, from Chinnereth even unto the sea of the plain, even the salt sea, under Ashdothpisgah eastward.
DEUT|3|18|And I commanded you at that time, saying, The LORD your God hath given you this land to possess it: ye shall pass over armed before your brethren the children of Israel, all that are meet for the war.
DEUT|3|19|But your wives, and your little ones, and your cattle, (for I know that ye have much cattle,) shall abide in your cities which I have given you;
DEUT|3|20|Until the LORD have given rest unto your brethren, as well as unto you, and until they also possess the land which the LORD your God hath given them beyond Jordan: and then shall ye return every man unto his possession, which I have given you.
DEUT|3|21|And I commanded Joshua at that time, saying, Thine eyes have seen all that the LORD your God hath done unto these two kings: so shall the LORD do unto all the kingdoms whither thou passest.
DEUT|3|22|Ye shall not fear them: for the LORD your God he shall fight for you.
DEUT|3|23|And I besought the LORD at that time, saying,
DEUT|3|24|O Lord GOD, thou hast begun to show thy servant thy greatness, and thy mighty hand: for what God is there in heaven or in earth, that can do according to thy works, and according to thy might?
DEUT|3|25|I pray thee, let me go over, and see the good land that is beyond Jordan, that goodly mountain, and Lebanon.
DEUT|3|26|But the LORD was wroth with me for your sakes, and would not hear me: and the LORD said unto me, Let it suffice thee; speak no more unto me of this matter.
DEUT|3|27|Get thee up into the top of Pisgah, and lift up thine eyes westward, and northward, and southward, and eastward, and behold it with thine eyes: for thou shalt not go over this Jordan.
DEUT|3|28|But charge Joshua, and encourage him, and strengthen him: for he shall go over before this people, and he shall cause them to inherit the land which thou shalt see.
DEUT|3|29|So we abode in the valley over against Bethpeor.
DEUT|4|1|Now therefore hearken, O Israel, unto the statutes and unto the judgments, which I teach you, for to do them, that ye may live, and go in and possess the land which the LORD God of your fathers giveth you.
DEUT|4|2|Ye shall not add unto the word which I command you, neither shall ye diminish ought from it, that ye may keep the commandments of the LORD your God which I command you.
DEUT|4|3|Your eyes have seen what the LORD did because of Baalpeor: for all the men that followed Baalpeor, the LORD thy God hath destroyed them from among you.
DEUT|4|4|But ye that did cleave unto the LORD your God are alive every one of you this day.
DEUT|4|5|Behold, I have taught you statutes and judgments, even as the LORD my God commanded me, that ye should do so in the land whither ye go to possess it.
DEUT|4|6|Keep therefore and do them; for this is your wisdom and your understanding in the sight of the nations, which shall hear all these statutes, and say, Surely this great nation is a wise and understanding people.
DEUT|4|7|For what nation is there so great, who hath God so nigh unto them, as the LORD our God is in all things that we call upon him for?
DEUT|4|8|And what nation is there so great, that hath statutes and judgments so righteous as all this law, which I set before you this day?
DEUT|4|9|Only take heed to thyself, and keep thy soul diligently, lest thou forget the things which thine eyes have seen, and lest they depart from thy heart all the days of thy life: but teach them thy sons, and thy sons' sons;
DEUT|4|10|Specially the day that thou stoodest before the LORD thy God in Horeb, when the LORD said unto me, Gather me the people together, and I will make them hear my words, that they may learn to fear me all the days that they shall live upon the earth, and that they may teach their children.
DEUT|4|11|And ye came near and stood under the mountain; and the mountain burned with fire unto the midst of heaven, with darkness, clouds, and thick darkness.
DEUT|4|12|And the LORD spake unto you out of the midst of the fire: ye heard the voice of the words, but saw no similitude; only ye heard a voice.
DEUT|4|13|And he declared unto you his covenant, which he commanded you to perform, even ten commandments; and he wrote them upon two tables of stone.
DEUT|4|14|And the LORD commanded me at that time to teach you statutes and judgments, that ye might do them in the land whither ye go over to possess it.
DEUT|4|15|Take ye therefore good heed unto yourselves; for ye saw no manner of similitude on the day that the LORD spake unto you in Horeb out of the midst of the fire:
DEUT|4|16|Lest ye corrupt yourselves, and make you a graven image, the similitude of any figure, the likeness of male or female,
DEUT|4|17|The likeness of any beast that is on the earth, the likeness of any winged fowl that flieth in the air,
DEUT|4|18|The likeness of any thing that creepeth on the ground, the likeness of any fish that is in the waters beneath the earth:
DEUT|4|19|And lest thou lift up thine eyes unto heaven, and when thou seest the sun, and the moon, and the stars, even all the host of heaven, shouldest be driven to worship them, and serve them, which the LORD thy God hath divided unto all nations under the whole heaven.
DEUT|4|20|But the LORD hath taken you, and brought you forth out of the iron furnace, even out of Egypt, to be unto him a people of inheritance, as ye are this day.
DEUT|4|21|Furthermore the LORD was angry with me for your sakes, and sware that I should not go over Jordan, and that I should not go in unto that good land, which the LORD thy God giveth thee for an inheritance:
DEUT|4|22|But I must die in this land, I must not go over Jordan: but ye shall go over, and possess that good land.
DEUT|4|23|Take heed unto yourselves, lest ye forget the covenant of the LORD your God, which he made with you, and make you a graven image, or the likeness of any thing, which the LORD thy God hath forbidden thee.
DEUT|4|24|For the LORD thy God is a consuming fire, even a jealous God.
DEUT|4|25|When thou shalt beget children, and children's children, and ye shall have remained long in the land, and shall corrupt yourselves, and make a graven image, or the likeness of any thing, and shall do evil in the sight of the LORD thy God, to provoke him to anger:
DEUT|4|26|I call heaven and earth to witness against you this day, that ye shall soon utterly perish from off the land whereunto ye go over Jordan to possess it; ye shall not prolong your days upon it, but shall utterly be destroyed.
DEUT|4|27|And the LORD shall scatter you among the nations, and ye shall be left few in number among the heathen, whither the LORD shall lead you.
DEUT|4|28|And there ye shall serve gods, the work of men's hands, wood and stone, which neither see, nor hear, nor eat, nor smell.
DEUT|4|29|But if from thence thou shalt seek the LORD thy God, thou shalt find him, if thou seek him with all thy heart and with all thy soul.
DEUT|4|30|When thou art in tribulation, and all these things are come upon thee, even in the latter days, if thou turn to the LORD thy God, and shalt be obedient unto his voice;
DEUT|4|31|(For the LORD thy God is a merciful God;) he will not forsake thee, neither destroy thee, nor forget the covenant of thy fathers which he sware unto them.
DEUT|4|32|For ask now of the days that are past, which were before thee, since the day that God created man upon the earth, and ask from the one side of heaven unto the other, whether there hath been any such thing as this great thing is, or hath been heard like it?
DEUT|4|33|Did ever people hear the voice of God speaking out of the midst of the fire, as thou hast heard, and live?
DEUT|4|34|Or hath God assayed to go and take him a nation from the midst of another nation, by temptations, by signs, and by wonders, and by war, and by a mighty hand, and by a stretched out arm, and by great terrors, according to all that the LORD your God did for you in Egypt before your eyes?
DEUT|4|35|Unto thee it was showed, that thou mightest know that the LORD he is God; there is none else beside him.
DEUT|4|36|Out of heaven he made thee to hear his voice, that he might instruct thee: and upon earth he showed thee his great fire; and thou heardest his words out of the midst of the fire.
DEUT|4|37|And because he loved thy fathers, therefore he chose their seed after them, and brought thee out in his sight with his mighty power out of Egypt;
DEUT|4|38|To drive out nations from before thee greater and mightier than thou art, to bring thee in, to give thee their land for an inheritance, as it is this day.
DEUT|4|39|Know therefore this day, and consider it in thine heart, that the LORD he is God in heaven above, and upon the earth beneath: there is none else.
DEUT|4|40|Thou shalt keep therefore his statutes, and his commandments, which I command thee this day, that it may go well with thee, and with thy children after thee, and that thou mayest prolong thy days upon the earth, which the LORD thy God giveth thee, for ever.
DEUT|4|41|Then Moses severed three cities on this side Jordan toward the sunrising;
DEUT|4|42|That the slayer might flee thither, which should kill his neighbor unawares, and hated him not in times past; and that fleeing unto one of these cities he might live:
DEUT|4|43|Namely, Bezer in the wilderness, in the plain country, of the Reubenites; and Ramoth in Gilead, of the Gadites; and Golan in Bashan, of the Manassites.
DEUT|4|44|And this is the law which Moses set before the children of Israel:
DEUT|4|45|These are the testimonies, and the statutes, and the judgments, which Moses spake unto the children of Israel, after they came forth out of Egypt.
DEUT|4|46|On this side Jordan, in the valley over against Bethpeor, in the land of Sihon king of the Amorites, who dwelt at Heshbon, whom Moses and the children of Israel smote, after they were come forth out of Egypt:
DEUT|4|47|And they possessed his land, and the land of Og king of Bashan, two kings of the Amorites, which were on this side Jordan toward the sunrising;
DEUT|4|48|From Aroer, which is by the bank of the river Arnon, even unto mount Sion, which is Hermon,
DEUT|4|49|And all the plain on this side Jordan eastward, even unto the sea of the plain, under the springs of Pisgah.
DEUT|5|1|And Moses called all Israel, and said unto them, Hear, O Israel, the statutes and judgments which I speak in your ears this day, that ye may learn them, and keep, and do them.
DEUT|5|2|The LORD our God made a covenant with us in Horeb.
DEUT|5|3|The LORD made not this covenant with our fathers, but with us, even us, who are all of us here alive this day.
DEUT|5|4|The LORD talked with you face to face in the mount out of the midst of the fire,
DEUT|5|5|(I stood between the LORD and you at that time, to show you the word of the LORD: for ye were afraid by reason of the fire, and went not up into the mount;) saying,
DEUT|5|6|I am the LORD thy God, which brought thee out of the land of Egypt, from the house of bondage.
DEUT|5|7|Thou shalt have none other gods before me.
DEUT|5|8|Thou shalt not make thee any graven image, or any likeness of any thing that is in heaven above, or that is in the earth beneath, or that is in the waters beneath the earth:
DEUT|5|9|Thou shalt not bow down thyself unto them, nor serve them: for I the LORD thy God am a jealous God, visiting the iniquity of the fathers upon the children unto the third and fourth generation of them that hate me,
DEUT|5|10|And showing mercy unto thousands of them that love me and keep my commandments.
DEUT|5|11|Thou shalt not take the name of the LORD thy God in vain: for the LORD will not hold him guiltless that taketh his name in vain.
DEUT|5|12|Keep the sabbath day to sanctify it, as the LORD thy God hath commanded thee.
DEUT|5|13|Six days thou shalt labor, and do all thy work:
DEUT|5|14|But the seventh day is the sabbath of the LORD thy God: in it thou shalt not do any work, thou, nor thy son, nor thy daughter, nor thy manservant, nor thy maidservant, nor thine ox, nor thine ass, nor any of thy cattle, nor thy stranger that is within thy gates; that thy manservant and thy maidservant may rest as well as thou.
DEUT|5|15|And remember that thou wast a servant in the land of Egypt, and that the LORD thy God brought thee out thence through a mighty hand and by a stretched out arm: therefore the LORD thy God commanded thee to keep the sabbath day.
DEUT|5|16|Honor thy father and thy mother, as the LORD thy God hath commanded thee; that thy days may be prolonged, and that it may go well with thee, in the land which the LORD thy God giveth thee.
DEUT|5|17|Thou shalt not kill.
DEUT|5|18|Neither shalt thou commit adultery.
DEUT|5|19|Neither shalt thou steal.
DEUT|5|20|Neither shalt thou bear false witness against thy neighbor.
DEUT|5|21|Neither shalt thou desire thy neighbor's wife, neither shalt thou covet thy neighbor's house, his field, or his manservant, or his maidservant, his ox, or his ass, or any thing that is thy neighbor's.
DEUT|5|22|These words the LORD spake unto all your assembly in the mount out of the midst of the fire, of the cloud, and of the thick darkness, with a great voice: and he added no more. And he wrote them in two tables of stone, and delivered them unto me.
DEUT|5|23|And it came to pass, when ye heard the voice out of the midst of the darkness, (for the mountain did burn with fire,) that ye came near unto me, even all the heads of your tribes, and your elders;
DEUT|5|24|And ye said, Behold, the LORD our God hath showed us his glory and his greatness, and we have heard his voice out of the midst of the fire: we have seen this day that God doth talk with man, and he liveth.
DEUT|5|25|Now therefore why should we die? for this great fire will consume us: if we hear the voice of the LORD our God any more, then we shall die.
DEUT|5|26|For who is there of all flesh, that hath heard the voice of the living God speaking out of the midst of the fire, as we have, and lived?
DEUT|5|27|Go thou near, and hear all that the LORD our God shall say: and speak thou unto us all that the LORD our God shall speak unto thee; and we will hear it, and do it.
DEUT|5|28|And the LORD heard the voice of your words, when ye spake unto me; and the LORD said unto me, I have heard the voice of the words of this people, which they have spoken unto thee: they have well said all that they have spoken.
DEUT|5|29|O that there were such an heart in them, that they would fear me, and keep all my commandments always, that it might be well with them, and with their children for ever!
DEUT|5|30|Go say to them, Get you into your tents again.
DEUT|5|31|But as for thee, stand thou here by me, and I will speak unto thee all the commandments, and the statutes, and the judgments, which thou shalt teach them, that they may do them in the land which I give them to possess it.
DEUT|5|32|Ye shall observe to do therefore as the LORD your God hath commanded you: ye shall not turn aside to the right hand or to the left.
DEUT|5|33|Ye shall walk in all the ways which the LORD your God hath commanded you, that ye may live, and that it may be well with you, and that ye may prolong your days in the land which ye shall possess.
DEUT|6|1|Now these are the commandments, the statutes, and the judgments, which the LORD your God commanded to teach you, that ye might do them in the land whither ye go to possess it:
DEUT|6|2|That thou mightest fear the LORD thy God, to keep all his statutes and his commandments, which I command thee, thou, and thy son, and thy son's son, all the days of thy life; and that thy days may be prolonged.
DEUT|6|3|Hear therefore, O Israel, and observe to do it; that it may be well with thee, and that ye may increase mightily, as the LORD God of thy fathers hath promised thee, in the land that floweth with milk and honey.
DEUT|6|4|Hear, O Israel: The LORD our God is one LORD:
DEUT|6|5|And thou shalt love the LORD thy God with all thine heart, and with all thy soul, and with all thy might.
DEUT|6|6|And these words, which I command thee this day, shall be in thine heart:
DEUT|6|7|And thou shalt teach them diligently unto thy children, and shalt talk of them when thou sittest in thine house, and when thou walkest by the way, and when thou liest down, and when thou risest up.
DEUT|6|8|And thou shalt bind them for a sign upon thine hand, and they shall be as frontlets between thine eyes.
DEUT|6|9|And thou shalt write them upon the posts of thy house, and on thy gates.
DEUT|6|10|And it shall be, when the LORD thy God shall have brought thee into the land which he sware unto thy fathers, to Abraham, to Isaac, and to Jacob, to give thee great and goodly cities, which thou buildedst not,
DEUT|6|11|And houses full of all good things, which thou filledst not, and wells digged, which thou diggedst not, vineyards and olive trees, which thou plantedst not; when thou shalt have eaten and be full;
DEUT|6|12|Then beware lest thou forget the LORD, which brought thee forth out of the land of Egypt, from the house of bondage.
DEUT|6|13|Thou shalt fear the LORD thy God, and serve him, and shalt swear by his name.
DEUT|6|14|Ye shall not go after other gods, of the gods of the people which are round about you;
DEUT|6|15|(For the LORD thy God is a jealous God among you) lest the anger of the LORD thy God be kindled against thee, and destroy thee from off the face of the earth.
DEUT|6|16|Ye shall not tempt the LORD your God, as ye tempted him in Massah.
DEUT|6|17|Ye shall diligently keep the commandments of the LORD your God, and his testimonies, and his statutes, which he hath commanded thee.
DEUT|6|18|And thou shalt do that which is right and good in the sight of the LORD: that it may be well with thee, and that thou mayest go in and possess the good land which the LORD sware unto thy fathers.
DEUT|6|19|To cast out all thine enemies from before thee, as the LORD hath spoken.
DEUT|6|20|And when thy son asketh thee in time to come, saying, What mean the testimonies, and the statutes, and the judgments, which the LORD our God hath commanded you?
DEUT|6|21|Then thou shalt say unto thy son, We were Pharaoh's bondmen in Egypt; and the LORD brought us out of Egypt with a mighty hand:
DEUT|6|22|And the LORD showed signs and wonders, great and sore, upon Egypt, upon Pharaoh, and upon all his household, before our eyes:
DEUT|6|23|And he brought us out from thence, that he might bring us in, to give us the land which he sware unto our fathers.
DEUT|6|24|And the LORD commanded us to do all these statutes, to fear the LORD our God, for our good always, that he might preserve us alive, as it is at this day.
DEUT|6|25|And it shall be our righteousness, if we observe to do all these commandments before the LORD our God, as he hath commanded us.
DEUT|7|1|When the LORD thy God shall bring thee into the land whither thou goest to possess it, and hath cast out many nations before thee, the Hittites, and the Girgashites, and the Amorites, and the Canaanites, and the Perizzites, and the Hivites, and the Jebusites, seven nations greater and mightier than thou;
DEUT|7|2|And when the LORD thy God shall deliver them before thee; thou shalt smite them, and utterly destroy them; thou shalt make no covenant with them, nor show mercy unto them:
DEUT|7|3|Neither shalt thou make marriages with them; thy daughter thou shalt not give unto his son, nor his daughter shalt thou take unto thy son.
DEUT|7|4|For they will turn away thy son from following me, that they may serve other gods: so will the anger of the LORD be kindled against you, and destroy thee suddenly.
DEUT|7|5|But thus shall ye deal with them; ye shall destroy their altars, and break down their images, and cut down their groves, and burn their graven images with fire.
DEUT|7|6|For thou art an holy people unto the LORD thy God: the LORD thy God hath chosen thee to be a special people unto himself, above all people that are upon the face of the earth.
DEUT|7|7|The LORD did not set his love upon you, nor choose you, because ye were more in number than any people; for ye were the fewest of all people:
DEUT|7|8|But because the LORD loved you, and because he would keep the oath which he had sworn unto your fathers, hath the LORD brought you out with a mighty hand, and redeemed you out of the house of bondmen, from the hand of Pharaoh king of Egypt.
DEUT|7|9|Know therefore that the LORD thy God, he is God, the faithful God, which keepeth covenant and mercy with them that love him and keep his commandments to a thousand generations;
DEUT|7|10|And repayeth them that hate him to their face, to destroy them: he will not be slack to him that hateth him, he will repay him to his face.
DEUT|7|11|Thou shalt therefore keep the commandments, and the statutes, and the judgments, which I command thee this day, to do them.
DEUT|7|12|Wherefore it shall come to pass, if ye hearken to these judgments, and keep, and do them, that the LORD thy God shall keep unto thee the covenant and the mercy which he sware unto thy fathers:
DEUT|7|13|And he will love thee, and bless thee, and multiply thee: he will also bless the fruit of thy womb, and the fruit of thy land, thy corn, and thy wine, and thine oil, the increase of thy kine, and the flocks of thy sheep, in the land which he sware unto thy fathers to give thee.
DEUT|7|14|Thou shalt be blessed above all people: there shall not be male or female barren among you, or among your cattle.
DEUT|7|15|And the LORD will take away from thee all sickness, and will put none of the evil diseases of Egypt, which thou knowest, upon thee; but will lay them upon all them that hate thee.
DEUT|7|16|And thou shalt consume all the people which the LORD thy God shall deliver thee; thine eye shall have no pity upon them: neither shalt thou serve their gods; for that will be a snare unto thee.
DEUT|7|17|If thou shalt say in thine heart, These nations are more than I; how can I dispossess them?
DEUT|7|18|Thou shalt not be afraid of them: but shalt well remember what the LORD thy God did unto Pharaoh, and unto all Egypt;
DEUT|7|19|The great temptations which thine eyes saw, and the signs, and the wonders, and the mighty hand, and the stretched out arm, whereby the LORD thy God brought thee out: so shall the LORD thy God do unto all the people of whom thou art afraid.
DEUT|7|20|Moreover the LORD thy God will send the hornet among them, until they that are left, and hide themselves from thee, be destroyed.
DEUT|7|21|Thou shalt not be affrighted at them: for the LORD thy God is among you, a mighty God and terrible.
DEUT|7|22|And the LORD thy God will put out those nations before thee by little and little: thou mayest not consume them at once, lest the beasts of the field increase upon thee.
DEUT|7|23|But the LORD thy God shall deliver them unto thee, and shall destroy them with a mighty destruction, until they be destroyed.
DEUT|7|24|And he shall deliver their kings into thine hand, and thou shalt destroy their name from under heaven: there shall no man be able to stand before thee, until thou have destroyed them.
DEUT|7|25|The graven images of their gods shall ye burn with fire: thou shalt not desire the silver or gold that is on them, nor take it unto thee, lest thou be snared therein: for it is an abomination to the LORD thy God.
DEUT|7|26|Neither shalt thou bring an abomination into thine house, lest thou be a cursed thing like it: but thou shalt utterly detest it, and thou shalt utterly abhor it; for it is a cursed thing.
DEUT|8|1|All the commandments which I command thee this day shall ye observe to do, that ye may live, and multiply, and go in and possess the land which the LORD sware unto your fathers.
DEUT|8|2|And thou shalt remember all the way which the LORD thy God led thee these forty years in the wilderness, to humble thee, and to prove thee, to know what was in thine heart, whether thou wouldest keep his commandments, or no.
DEUT|8|3|And he humbled thee, and suffered thee to hunger, and fed thee with manna, which thou knewest not, neither did thy fathers know; that he might make thee know that man doth not live by bread only, but by every word that proceedeth out of the mouth of the LORD doth man live.
DEUT|8|4|Thy raiment waxed not old upon thee, neither did thy foot swell, these forty years.
DEUT|8|5|Thou shalt also consider in thine heart, that, as a man chasteneth his son, so the LORD thy God chasteneth thee.
DEUT|8|6|Therefore thou shalt keep the commandments of the LORD thy God, to walk in his ways, and to fear him.
DEUT|8|7|For the LORD thy God bringeth thee into a good land, a land of brooks of water, of fountains and depths that spring out of valleys and hills;
DEUT|8|8|A land of wheat, and barley, and vines, and fig trees, and pomegranates; a land of oil olive, and honey;
DEUT|8|9|A land wherein thou shalt eat bread without scarceness, thou shalt not lack any thing in it; a land whose stones are iron, and out of whose hills thou mayest dig brass.
DEUT|8|10|When thou hast eaten and art full, then thou shalt bless the LORD thy God for the good land which he hath given thee.
DEUT|8|11|Beware that thou forget not the LORD thy God, in not keeping his commandments, and his judgments, and his statutes, which I command thee this day:
DEUT|8|12|Lest when thou hast eaten and art full, and hast built goodly houses, and dwelt therein;
DEUT|8|13|And when thy herds and thy flocks multiply, and thy silver and thy gold is multiplied, and all that thou hast is multiplied;
DEUT|8|14|Then thine heart be lifted up, and thou forget the LORD thy God, which brought thee forth out of the land of Egypt, from the house of bondage;
DEUT|8|15|Who led thee through that great and terrible wilderness, wherein were fiery serpents, and scorpions, and drought, where there was no water; who brought thee forth water out of the rock of flint;
DEUT|8|16|Who fed thee in the wilderness with manna, which thy fathers knew not, that he might humble thee, and that he might prove thee, to do thee good at thy latter end;
DEUT|8|17|And thou say in thine heart, My power and the might of mine hand hath gotten me this wealth.
DEUT|8|18|But thou shalt remember the LORD thy God: for it is he that giveth thee power to get wealth, that he may establish his covenant which he sware unto thy fathers, as it is this day.
DEUT|8|19|And it shall be, if thou do at all forget the LORD thy God, and walk after other gods, and serve them, and worship them, I testify against you this day that ye shall surely perish.
DEUT|8|20|As the nations which the LORD destroyeth before your face, so shall ye perish; because ye would not be obedient unto the voice of the LORD your God.
DEUT|9|1|Hear, O Israel: Thou art to pass over Jordan this day, to go in to possess nations greater and mightier than thyself, cities great and fenced up to heaven,
DEUT|9|2|A people great and tall, the children of the Anakims, whom thou knowest, and of whom thou hast heard say, Who can stand before the children of Anak!
DEUT|9|3|Understand therefore this day, that the LORD thy God is he which goeth over before thee; as a consuming fire he shall destroy them, and he shall bring them down before thy face: so shalt thou drive them out, and destroy them quickly, as the LORD hath said unto thee.
DEUT|9|4|Speak not thou in thine heart, after that the LORD thy God hath cast them out from before thee, saying, For my righteousness the LORD hath brought me in to possess this land: but for the wickedness of these nations the LORD doth drive them out from before thee.
DEUT|9|5|Not for thy righteousness, or for the uprightness of thine heart, dost thou go to possess their land: but for the wickedness of these nations the LORD thy God doth drive them out from before thee, and that he may perform the word which the LORD sware unto thy fathers, Abraham, Isaac, and Jacob.
DEUT|9|6|Understand therefore, that the LORD thy God giveth thee not this good land to possess it for thy righteousness; for thou art a stiffnecked people.
DEUT|9|7|Remember, and forget not, how thou provokedst the LORD thy God to wrath in the wilderness: from the day that thou didst depart out of the land of Egypt, until ye came unto this place, ye have been rebellious against the LORD.
DEUT|9|8|Also in Horeb ye provoked the LORD to wrath, so that the LORD was angry with you to have destroyed you.
DEUT|9|9|When I was gone up into the mount to receive the tables of stone, even the tables of the covenant which the LORD made with you, then I abode in the mount forty days and forty nights, I neither did eat bread nor drink water:
DEUT|9|10|And the LORD delivered unto me two tables of stone written with the finger of God; and on them was written according to all the words, which the LORD spake with you in the mount out of the midst of the fire in the day of the assembly.
DEUT|9|11|And it came to pass at the end of forty days and forty nights, that the LORD gave me the two tables of stone, even the tables of the covenant.
DEUT|9|12|And the LORD said unto me, Arise, get thee down quickly from hence; for thy people which thou hast brought forth out of Egypt have corrupted themselves; they are quickly turned aside out of the way which I commanded them; they have made them a molten image.
DEUT|9|13|Furthermore the LORD spake unto me, saying, I have seen this people, and, behold, it is a stiffnecked people:
DEUT|9|14|Let me alone, that I may destroy them, and blot out their name from under heaven: and I will make of thee a nation mightier and greater than they.
DEUT|9|15|So I turned and came down from the mount, and the mount burned with fire: and the two tables of the covenant were in my two hands.
DEUT|9|16|And I looked, and, behold, ye had sinned against the LORD your God, and had made you a molten calf: ye had turned aside quickly out of the way which the LORD had commanded you.
DEUT|9|17|And I took the two tables, and cast them out of my two hands, and brake them before your eyes.
DEUT|9|18|And I fell down before the LORD, as at the first, forty days and forty nights: I did neither eat bread, nor drink water, because of all your sins which ye sinned, in doing wickedly in the sight of the LORD, to provoke him to anger.
DEUT|9|19|For I was afraid of the anger and hot displeasure, wherewith the LORD was wroth against you to destroy you. But the LORD hearkened unto me at that time also.
DEUT|9|20|And the LORD was very angry with Aaron to have destroyed him: and I prayed for Aaron also the same time.
DEUT|9|21|And I took your sin, the calf which ye had made, and burnt it with fire, and stamped it, and ground it very small, even until it was as small as dust: and I cast the dust thereof into the brook that descended out of the mount.
DEUT|9|22|And at Taberah, and at Massah, and at Kibrothhattaavah, ye provoked the LORD to wrath.
DEUT|9|23|Likewise when the LORD sent you from Kadeshbarnea, saying, Go up and possess the land which I have given you; then ye rebelled against the commandment of the LORD your God, and ye believed him not, nor hearkened to his voice.
DEUT|9|24|Ye have been rebellious against the LORD from the day that I knew you.
DEUT|9|25|Thus I fell down before the LORD forty days and forty nights, as I fell down at the first; because the LORD had said he would destroy you.
DEUT|9|26|I prayed therefore unto the LORD, and said, O Lord GOD, destroy not thy people and thine inheritance, which thou hast redeemed through thy greatness, which thou hast brought forth out of Egypt with a mighty hand.
DEUT|9|27|Remember thy servants, Abraham, Isaac, and Jacob; look not unto the stubbornness of this people, nor to their wickedness, nor to their sin:
DEUT|9|28|Lest the land whence thou broughtest us out say, Because the LORD was not able to bring them into the land which he promised them, and because he hated them, he hath brought them out to slay them in the wilderness.
DEUT|9|29|Yet they are thy people and thine inheritance, which thou broughtest out by thy mighty power and by thy stretched out arm.
DEUT|10|1|At that time the LORD said unto me, Hew thee two tables of stone like unto the first, and come up unto me into the mount, and make thee an ark of wood.
DEUT|10|2|And I will write on the tables the words that were in the first tables which thou brakest, and thou shalt put them in the ark.
DEUT|10|3|And I made an ark of shittim wood, and hewed two tables of stone like unto the first, and went up into the mount, having the two tables in mine hand.
DEUT|10|4|And he wrote on the tables, according to the first writing, the ten commandments, which the LORD spake unto you in the mount out of the midst of the fire in the day of the assembly: and the LORD gave them unto me.
DEUT|10|5|And I turned myself and came down from the mount, and put the tables in the ark which I had made; and there they be, as the LORD commanded me.
DEUT|10|6|And the children of Israel took their journey from Beeroth of the children of Jaakan to Mosera: there Aaron died, and there he was buried; and Eleazar his son ministered in the priest's office in his stead.
DEUT|10|7|From thence they journeyed unto Gudgodah; and from Gudgodah to Jotbath, a land of rivers of waters.
DEUT|10|8|At that time the LORD separated the tribe of Levi, to bear the ark of the covenant of the LORD, to stand before the LORD to minister unto him, and to bless in his name, unto this day.
DEUT|10|9|Wherefore Levi hath no part nor inheritance with his brethren; the LORD is his inheritance, according as the LORD thy God promised him.
DEUT|10|10|And I stayed in the mount, according to the first time, forty days and forty nights; and the LORD hearkened unto me at that time also, and the LORD would not destroy thee.
DEUT|10|11|And the LORD said unto me, Arise, take thy journey before the people, that they may go in and possess the land, which I sware unto their fathers to give unto them.
DEUT|10|12|And now, Israel, what doth the LORD thy God require of thee, but to fear the LORD thy God, to walk in all his ways, and to love him, and to serve the LORD thy God with all thy heart and with all thy soul,
DEUT|10|13|To keep the commandments of the LORD, and his statutes, which I command thee this day for thy good?
DEUT|10|14|Behold, the heaven and the heaven of heavens is the LORD's thy God, the earth also, with all that therein is.
DEUT|10|15|Only the LORD had a delight in thy fathers to love them, and he chose their seed after them, even you above all people, as it is this day.
DEUT|10|16|Circumcise therefore the foreskin of your heart, and be no more stiffnecked.
DEUT|10|17|For the LORD your God is God of gods, and Lord of lords, a great God, a mighty, and a terrible, which regardeth not persons, nor taketh reward:
DEUT|10|18|He doth execute the judgment of the fatherless and widow, and loveth the stranger, in giving him food and raiment.
DEUT|10|19|Love ye therefore the stranger: for ye were strangers in the land of Egypt.
DEUT|10|20|Thou shalt fear the LORD thy God; him shalt thou serve, and to him shalt thou cleave, and swear by his name.
DEUT|10|21|He is thy praise, and he is thy God, that hath done for thee these great and terrible things, which thine eyes have seen.
DEUT|10|22|Thy fathers went down into Egypt with threescore and ten persons; and now the LORD thy God hath made thee as the stars of heaven for multitude.
DEUT|11|1|Therefore thou shalt love the LORD thy God, and keep his charge, and his statutes, and his judgments, and his commandments, alway.
DEUT|11|2|And know ye this day: for I speak not with your children which have not known, and which have not seen the chastisement of the LORD your God, his greatness, his mighty hand, and his stretched out arm,
DEUT|11|3|And his miracles, and his acts, which he did in the midst of Egypt unto Pharaoh the king of Egypt, and unto all his land;
DEUT|11|4|And what he did unto the army of Egypt, unto their horses, and to their chariots; how he made the water of the Red sea to overflow them as they pursued after you, and how the LORD hath destroyed them unto this day;
DEUT|11|5|And what he did unto you in the wilderness, until ye came into this place;
DEUT|11|6|And what he did unto Dathan and Abiram, the sons of Eliab, the son of Reuben: how the earth opened her mouth, and swallowed them up, and their households, and their tents, and all the substance that was in their possession, in the midst of all Israel:
DEUT|11|7|But your eyes have seen all the great acts of the LORD which he did.
DEUT|11|8|Therefore shall ye keep all the commandments which I command you this day, that ye may be strong, and go in and possess the land, whither ye go to possess it;
DEUT|11|9|And that ye may prolong your days in the land, which the LORD sware unto your fathers to give unto them and to their seed, a land that floweth with milk and honey.
DEUT|11|10|For the land, whither thou goest in to possess it, is not as the land of Egypt, from whence ye came out, where thou sowedst thy seed, and wateredst it with thy foot, as a garden of herbs:
DEUT|11|11|But the land, whither ye go to possess it, is a land of hills and valleys, and drinketh water of the rain of heaven:
DEUT|11|12|A land which the LORD thy God careth for: the eyes of the LORD thy God are always upon it, from the beginning of the year even unto the end of the year.
DEUT|11|13|And it shall come to pass, if ye shall hearken diligently unto my commandments which I command you this day, to love the LORD your God, and to serve him with all your heart and with all your soul,
DEUT|11|14|That I will give you the rain of your land in his due season, the first rain and the latter rain, that thou mayest gather in thy corn, and thy wine, and thine oil.
DEUT|11|15|And I will send grass in thy fields for thy cattle, that thou mayest eat and be full.
DEUT|11|16|Take heed to yourselves, that your heart be not deceived, and ye turn aside, and serve other gods, and worship them;
DEUT|11|17|And then the LORD's wrath be kindled against you, and he shut up the heaven, that there be no rain, and that the land yield not her fruit; and lest ye perish quickly from off the good land which the LORD giveth you.
DEUT|11|18|Therefore shall ye lay up these my words in your heart and in your soul, and bind them for a sign upon your hand, that they may be as frontlets between your eyes.
DEUT|11|19|And ye shall teach them your children, speaking of them when thou sittest in thine house, and when thou walkest by the way, when thou liest down, and when thou risest up.
DEUT|11|20|And thou shalt write them upon the door posts of thine house, and upon thy gates:
DEUT|11|21|That your days may be multiplied, and the days of your children, in the land which the LORD sware unto your fathers to give them, as the days of heaven upon the earth.
DEUT|11|22|For if ye shall diligently keep all these commandments which I command you, to do them, to love the LORD your God, to walk in all his ways, and to cleave unto him;
DEUT|11|23|Then will the LORD drive out all these nations from before you, and ye shall possess greater nations and mightier than yourselves.
DEUT|11|24|Every place whereon the soles of your feet shall tread shall be yours: from the wilderness and Lebanon, from the river, the river Euphrates, even unto the uttermost sea shall your coast be.
DEUT|11|25|There shall no man be able to stand before you: for the LORD your God shall lay the fear of you and the dread of you upon all the land that ye shall tread upon, as he hath said unto you.
DEUT|11|26|Behold, I set before you this day a blessing and a curse;
DEUT|11|27|A blessing, if ye obey the commandments of the LORD your God, which I command you this day:
DEUT|11|28|And a curse, if ye will not obey the commandments of the LORD your God, but turn aside out of the way which I command you this day, to go after other gods, which ye have not known.
DEUT|11|29|And it shall come to pass, when the LORD thy God hath brought thee in unto the land whither thou goest to possess it, that thou shalt put the blessing upon mount Gerizim, and the curse upon mount Ebal.
DEUT|11|30|Are they not on the other side Jordan, by the way where the sun goeth down, in the land of the Canaanites, which dwell in the champaign over against Gilgal, beside the plains of Moreh?
DEUT|11|31|For ye shall pass over Jordan to go in to possess the land which the LORD your God giveth you, and ye shall possess it, and dwell therein.
DEUT|11|32|And ye shall observe to do all the statutes and judgments which I set before you this day.
DEUT|12|1|These are the statutes and judgments, which ye shall observe to do in the land, which the LORD God of thy fathers giveth thee to possess it, all the days that ye live upon the earth.
DEUT|12|2|Ye shall utterly destroy all the places, wherein the nations which ye shall possess served their gods, upon the high mountains, and upon the hills, and under every green tree:
DEUT|12|3|And ye shall overthrow their altars, and break their pillars, and burn their groves with fire; and ye shall hew down the graven images of their gods, and destroy the names of them out of that place.
DEUT|12|4|Ye shall not do so unto the LORD your God.
DEUT|12|5|But unto the place which the LORD your God shall choose out of all your tribes to put his name there, even unto his habitation shall ye seek, and thither thou shalt come:
DEUT|12|6|And thither ye shall bring your burnt offerings, and your sacrifices, and your tithes, and heave offerings of your hand, and your vows, and your freewill offerings, and the firstlings of your herds and of your flocks:
DEUT|12|7|And there ye shall eat before the LORD your God, and ye shall rejoice in all that ye put your hand unto, ye and your households, wherein the LORD thy God hath blessed thee.
DEUT|12|8|Ye shall not do after all the things that we do here this day, every man whatsoever is right in his own eyes.
DEUT|12|9|For ye are not as yet come to the rest and to the inheritance, which the LORD your God giveth you.
DEUT|12|10|But when ye go over Jordan, and dwell in the land which the LORD your God giveth you to inherit, and when he giveth you rest from all your enemies round about, so that ye dwell in safety;
DEUT|12|11|Then there shall be a place which the LORD your God shall choose to cause his name to dwell there; thither shall ye bring all that I command you; your burnt offerings, and your sacrifices, your tithes, and the heave offering of your hand, and all your choice vows which ye vow unto the LORD:
DEUT|12|12|And ye shall rejoice before the LORD your God, ye, and your sons, and your daughters, and your menservants, and your maidservants, and the Levite that is within your gates; forasmuch as he hath no part nor inheritance with you.
DEUT|12|13|Take heed to thyself that thou offer not thy burnt offerings in every place that thou seest:
DEUT|12|14|But in the place which the LORD shall choose in one of thy tribes, there thou shalt offer thy burnt offerings, and there thou shalt do all that I command thee.
DEUT|12|15|Notwithstanding thou mayest kill and eat flesh in all thy gates, whatsoever thy soul lusteth after, according to the blessing of the LORD thy God which he hath given thee: the unclean and the clean may eat thereof, as of the roebuck, and as of the hart.
DEUT|12|16|Only ye shall not eat the blood; ye shall pour it upon the earth as water.
DEUT|12|17|Thou mayest not eat within thy gates the tithe of thy corn, or of thy wine, or of thy oil, or the firstlings of thy herds or of thy flock, nor any of thy vows which thou vowest, nor thy freewill offerings, or heave offering of thine hand:
DEUT|12|18|But thou must eat them before the LORD thy God in the place which the LORD thy God shall choose, thou, and thy son, and thy daughter, and thy manservant, and thy maidservant, and the Levite that is within thy gates: and thou shalt rejoice before the LORD thy God in all that thou puttest thine hands unto.
DEUT|12|19|Take heed to thyself that thou forsake not the Levite as long as thou livest upon the earth.
DEUT|12|20|When the LORD thy God shall enlarge thy border, as he hath promised thee, and thou shalt say, I will eat flesh, because thy soul longeth to eat flesh; thou mayest eat flesh, whatsoever thy soul lusteth after.
DEUT|12|21|If the place which the LORD thy God hath chosen to put his name there be too far from thee, then thou shalt kill of thy herd and of thy flock, which the LORD hath given thee, as I have commanded thee, and thou shalt eat in thy gates whatsoever thy soul lusteth after.
DEUT|12|22|Even as the roebuck and the hart is eaten, so thou shalt eat them: the unclean and the clean shall eat of them alike.
DEUT|12|23|Only be sure that thou eat not the blood: for the blood is the life; and thou mayest not eat the life with the flesh.
DEUT|12|24|Thou shalt not eat it; thou shalt pour it upon the earth as water.
DEUT|12|25|Thou shalt not eat it; that it may go well with thee, and with thy children after thee, when thou shalt do that which is right in the sight of the LORD.
DEUT|12|26|Only thy holy things which thou hast, and thy vows, thou shalt take, and go unto the place which the LORD shall choose:
DEUT|12|27|And thou shalt offer thy burnt offerings, the flesh and the blood, upon the altar of the LORD thy God: and the blood of thy sacrifices shall be poured out upon the altar of the LORD thy God, and thou shalt eat the flesh.
DEUT|12|28|Observe and hear all these words which I command thee, that it may go well with thee, and with thy children after thee for ever, when thou doest that which is good and right in the sight of the LORD thy God.
DEUT|12|29|When the LORD thy God shall cut off the nations from before thee, whither thou goest to possess them, and thou succeedest them, and dwellest in their land;
DEUT|12|30|Take heed to thyself that thou be not snared by following them, after that they be destroyed from before thee; and that thou inquire not after their gods, saying, How did these nations serve their gods? even so will I do likewise.
DEUT|12|31|Thou shalt not do so unto the LORD thy God: for every abomination to the LORD, which he hateth, have they done unto their gods; for even their sons and their daughters they have burnt in the fire to their gods.
DEUT|12|32|What thing soever I command you, observe to do it: thou shalt not add thereto, nor diminish from it.
DEUT|13|1|If there arise among you a prophet, or a dreamer of dreams, and giveth thee a sign or a wonder,
DEUT|13|2|And the sign or the wonder come to pass, whereof he spake unto thee, saying, Let us go after other gods, which thou hast not known, and let us serve them;
DEUT|13|3|Thou shalt not hearken unto the words of that prophet, or that dreamer of dreams: for the LORD your God proveth you, to know whether ye love the LORD your God with all your heart and with all your soul.
DEUT|13|4|Ye shall walk after the LORD your God, and fear him, and keep his commandments, and obey his voice, and ye shall serve him, and cleave unto him.
DEUT|13|5|And that prophet, or that dreamer of dreams, shall be put to death; because he hath spoken to turn you away from the LORD your God, which brought you out of the land of Egypt, and redeemed you out of the house of bondage, to thrust thee out of the way which the LORD thy God commanded thee to walk in. So shalt thou put the evil away from the midst of thee.
DEUT|13|6|If thy brother, the son of thy mother, or thy son, or thy daughter, or the wife of thy bosom, or thy friend, which is as thine own soul, entice thee secretly, saying, Let us go and serve other gods, which thou hast not known, thou, nor thy fathers;
DEUT|13|7|Namely, of the gods of the people which are round about you, nigh unto thee, or far off from thee, from the one end of the earth even unto the other end of the earth;
DEUT|13|8|Thou shalt not consent unto him, nor hearken unto him; neither shall thine eye pity him, neither shalt thou spare, neither shalt thou conceal him:
DEUT|13|9|But thou shalt surely kill him; thine hand shall be first upon him to put him to death, and afterwards the hand of all the people.
DEUT|13|10|And thou shalt stone him with stones, that he die; because he hath sought to thrust thee away from the LORD thy God, which brought thee out of the land of Egypt, from the house of bondage.
DEUT|13|11|And all Israel shall hear, and fear, and shall do no more any such wickedness as this is among you.
DEUT|13|12|If thou shalt hear say in one of thy cities, which the LORD thy God hath given thee to dwell there, saying,
DEUT|13|13|Certain men, the children of Belial, are gone out from among you, and have withdrawn the inhabitants of their city, saying, Let us go and serve other gods, which ye have not known;
DEUT|13|14|Then shalt thou inquire, and make search, and ask diligently; and, behold, if it be truth, and the thing certain, that such abomination is wrought among you;
DEUT|13|15|Thou shalt surely smite the inhabitants of that city with the edge of the sword, destroying it utterly, and all that is therein, and the cattle thereof, with the edge of the sword.
DEUT|13|16|And thou shalt gather all the spoil of it into the midst of the street thereof, and shalt burn with fire the city, and all the spoil thereof every whit, for the LORD thy God: and it shall be an heap for ever; it shall not be built again.
DEUT|13|17|And there shall cleave nought of the cursed thing to thine hand: that the LORD may turn from the fierceness of his anger, and show thee mercy, and have compassion upon thee, and multiply thee, as he hath sworn unto thy fathers;
DEUT|13|18|When thou shalt hearken to the voice of the LORD thy God, to keep all his commandments which I command thee this day, to do that which is right in the eyes of the LORD thy God.
DEUT|14|1|Ye are the children of the LORD your God: ye shall not cut yourselves, nor make any baldness between your eyes for the dead.
DEUT|14|2|For thou art an holy people unto the LORD thy God, and the LORD hath chosen thee to be a peculiar people unto himself, above all the nations that are upon the earth.
DEUT|14|3|Thou shalt not eat any abominable thing.
DEUT|14|4|These are the beasts which ye shall eat: the ox, the sheep, and the goat,
DEUT|14|5|The hart, and the roebuck, and the fallow deer, and the wild goat, and the pygarg, and the wild ox, and the chamois.
DEUT|14|6|And every beast that parteth the hoof, and cleaveth the cleft into two claws, and cheweth the cud among the beasts, that ye shall eat.
DEUT|14|7|Nevertheless these ye shall not eat of them that chew the cud, or of them that divide the cloven hoof; as the camel, and the hare, and the coney: for they chew the cud, but divide not the hoof; therefore they are unclean unto you.
DEUT|14|8|And the swine, because it divideth the hoof, yet cheweth not the cud, it is unclean unto you: ye shall not eat of their flesh, nor touch their dead carcass.
DEUT|14|9|These ye shall eat of all that are in the waters: all that have fins and scales shall ye eat:
DEUT|14|10|And whatsoever hath not fins and scales ye may not eat; it is unclean unto you.
DEUT|14|11|Of all clean birds ye shall eat.
DEUT|14|12|But these are they of which ye shall not eat: the eagle, and the ossifrage, and the ospray,
DEUT|14|13|And the glede, and the kite, and the vulture after his kind,
DEUT|14|14|And every raven after his kind,
DEUT|14|15|And the owl, and the night hawk, and the cuckoo, and the hawk after his kind,
DEUT|14|16|The little owl, and the great owl, and the swan,
DEUT|14|17|And the pelican, and the gier eagle, and the cormorant,
DEUT|14|18|And the stork, and the heron after her kind, and the lapwing, and the bat.
DEUT|14|19|And every creeping thing that flieth is unclean unto you: they shall not be eaten.
DEUT|14|20|But of all clean fowls ye may eat.
DEUT|14|21|Ye shall not eat of anything that dieth of itself: thou shalt give it unto the stranger that is in thy gates, that he may eat it; or thou mayest sell it unto an alien: for thou art an holy people unto the LORD thy God. Thou shalt not seethe a kid in his mother's milk.
DEUT|14|22|Thou shalt truly tithe all the increase of thy seed, that the field bringeth forth year by year.
DEUT|14|23|And thou shalt eat before the LORD thy God, in the place which he shall choose to place his name there, the tithe of thy corn, of thy wine, and of thine oil, and the firstlings of thy herds and of thy flocks; that thou mayest learn to fear the LORD thy God always.
DEUT|14|24|And if the way be too long for thee, so that thou art not able to carry it; or if the place be too far from thee, which the LORD thy God shall choose to set his name there, when the LORD thy God hath blessed thee:
DEUT|14|25|Then shalt thou turn it into money, and bind up the money in thine hand, and shalt go unto the place which the LORD thy God shall choose:
DEUT|14|26|And thou shalt bestow that money for whatsoever thy soul lusteth after, for oxen, or for sheep, or for wine, or for strong drink, or for whatsoever thy soul desireth: and thou shalt eat there before the LORD thy God, and thou shalt rejoice, thou, and thine household,
DEUT|14|27|And the Levite that is within thy gates; thou shalt not forsake him; for he hath no part nor inheritance with thee.
DEUT|14|28|At the end of three years thou shalt bring forth all the tithe of thine increase the same year, and shalt lay it up within thy gates:
DEUT|14|29|And the Levite, (because he hath no part nor inheritance with thee,) and the stranger, and the fatherless, and the widow, which are within thy gates, shall come, and shall eat and be satisfied; that the LORD thy God may bless thee in all the work of thine hand which thou doest.
DEUT|15|1|At the end of every seven years thou shalt make a release.
DEUT|15|2|And this is the manner of the release: Every creditor that lendeth ought unto his neighbor shall release it; he shall not exact it of his neighbor, or of his brother; because it is called the LORD's release.
DEUT|15|3|Of a foreigner thou mayest exact it again: but that which is thine with thy brother thine hand shall release;
DEUT|15|4|Save when there shall be no poor among you; for the LORD shall greatly bless thee in the land which the LORD thy God giveth thee for an inheritance to possess it:
DEUT|15|5|Only if thou carefully hearken unto the voice of the LORD thy God, to observe to do all these commandments which I command thee this day.
DEUT|15|6|For the LORD thy God blesseth thee, as he promised thee: and thou shalt lend unto many nations, but thou shalt not borrow; and thou shalt reign over many nations, but they shall not reign over thee.
DEUT|15|7|If there be among you a poor man of one of thy brethren within any of thy gates in thy land which the LORD thy God giveth thee, thou shalt not harden thine heart, nor shut thine hand from thy poor brother:
DEUT|15|8|But thou shalt open thine hand wide unto him, and shalt surely lend him sufficient for his need, in that which he wanteth.
DEUT|15|9|Beware that there be not a thought in thy wicked heart, saying, The seventh year, the year of release, is at hand; and thine eye be evil against thy poor brother, and thou givest him nought; and he cry unto the LORD against thee, and it be sin unto thee.
DEUT|15|10|Thou shalt surely give him, and thine heart shall not be grieved when thou givest unto him: because that for this thing the LORD thy God shall bless thee in all thy works, and in all that thou puttest thine hand unto.
DEUT|15|11|For the poor shall never cease out of the land: therefore I command thee, saying, Thou shalt open thine hand wide unto thy brother, to thy poor, and to thy needy, in thy land.
DEUT|15|12|And if thy brother, an Hebrew man, or an Hebrew woman, be sold unto thee, and serve thee six years; then in the seventh year thou shalt let him go free from thee.
DEUT|15|13|And when thou sendest him out free from thee, thou shalt not let him go away empty:
DEUT|15|14|Thou shalt furnish him liberally out of thy flock, and out of thy floor, and out of thy winepress: of that wherewith the LORD thy God hath blessed thee thou shalt give unto him.
DEUT|15|15|And thou shalt remember that thou wast a bondman in the land of Egypt, and the LORD thy God redeemed thee: therefore I command thee this thing to day.
DEUT|15|16|And it shall be, if he say unto thee, I will not go away from thee; because he loveth thee and thine house, because he is well with thee;
DEUT|15|17|Then thou shalt take an awl, and thrust it through his ear unto the door, and he shall be thy servant for ever. And also unto thy maidservant thou shalt do likewise.
DEUT|15|18|It shall not seem hard unto thee, when thou sendest him away free from thee; for he hath been worth a double hired servant to thee, in serving thee six years: and the LORD thy God shall bless thee in all that thou doest.
DEUT|15|19|All the firstling males that come of thy herd and of thy flock thou shalt sanctify unto the LORD thy God: thou shalt do no work with the firstling of thy bullock, nor shear the firstling of thy sheep.
DEUT|15|20|Thou shalt eat it before the LORD thy God year by year in the place which the LORD shall choose, thou and thy household.
DEUT|15|21|And if there be any blemish therein, as if it be lame, or blind, or have any ill blemish, thou shalt not sacrifice it unto the LORD thy God.
DEUT|15|22|Thou shalt eat it within thy gates: the unclean and the clean person shall eat it alike, as the roebuck, and as the hart.
DEUT|15|23|Only thou shalt not eat the blood thereof; thou shalt pour it upon the ground as water.
DEUT|16|1|Observe the month of Abib, and keep the passover unto the LORD thy God: for in the month of Abib the LORD thy God brought thee forth out of Egypt by night.
DEUT|16|2|Thou shalt therefore sacrifice the passover unto the LORD thy God, of the flock and the herd, in the place which the LORD shall choose to place his name there.
DEUT|16|3|Thou shalt eat no leavened bread with it; seven days shalt thou eat unleavened bread therewith, even the bread of affliction; for thou camest forth out of the land of Egypt in haste: that thou mayest remember the day when thou camest forth out of the land of Egypt all the days of thy life.
DEUT|16|4|And there shall be no leavened bread seen with thee in all thy coast seven days; neither shall there any thing of the flesh, which thou sacrificedst the first day at even, remain all night until the morning.
DEUT|16|5|Thou mayest not sacrifice the passover within any of thy gates, which the LORD thy God giveth thee:
DEUT|16|6|But at the place which the LORD thy God shall choose to place his name in, there thou shalt sacrifice the passover at even, at the going down of the sun, at the season that thou camest forth out of Egypt.
DEUT|16|7|And thou shalt roast and eat it in the place which the LORD thy God shall choose: and thou shalt turn in the morning, and go unto thy tents.
DEUT|16|8|Six days thou shalt eat unleavened bread: and on the seventh day shall be a solemn assembly to the LORD thy God: thou shalt do no work therein.
DEUT|16|9|Seven weeks shalt thou number unto thee: begin to number the seven weeks from such time as thou beginnest to put the sickle to the corn.
DEUT|16|10|And thou shalt keep the feast of weeks unto the LORD thy God with a tribute of a freewill offering of thine hand, which thou shalt give unto the LORD thy God, according as the LORD thy God hath blessed thee:
DEUT|16|11|And thou shalt rejoice before the LORD thy God, thou, and thy son, and thy daughter, and thy manservant, and thy maidservant, and the Levite that is within thy gates, and the stranger, and the fatherless, and the widow, that are among you, in the place which the LORD thy God hath chosen to place his name there.
DEUT|16|12|And thou shalt remember that thou wast a bondman in Egypt: and thou shalt observe and do these statutes.
DEUT|16|13|Thou shalt observe the feast of tabernacles seven days, after that thou hast gathered in thy corn and thy wine:
DEUT|16|14|And thou shalt rejoice in thy feast, thou, and thy son, and thy daughter, and thy manservant, and thy maidservant, and the Levite, the stranger, and the fatherless, and the widow, that are within thy gates.
DEUT|16|15|Seven days shalt thou keep a solemn feast unto the LORD thy God in the place which the LORD shall choose: because the LORD thy God shall bless thee in all thine increase, and in all the works of thine hands, therefore thou shalt surely rejoice.
DEUT|16|16|Three times in a year shall all thy males appear before the LORD thy God in the place which he shall choose; in the feast of unleavened bread, and in the feast of weeks, and in the feast of tabernacles: and they shall not appear before the LORD empty:
DEUT|16|17|Every man shall give as he is able, according to the blessing of the LORD thy God which he hath given thee.
DEUT|16|18|Judges and officers shalt thou make thee in all thy gates, which the LORD thy God giveth thee, throughout thy tribes: and they shall judge the people with just judgment.
DEUT|16|19|Thou shalt not wrest judgment; thou shalt not respect persons, neither take a gift: for a gift doth blind the eyes of the wise, and pervert the words of the righteous.
DEUT|16|20|That which is altogether just shalt thou follow, that thou mayest live, and inherit the land which the LORD thy God giveth thee.
DEUT|16|21|Thou shalt not plant thee a grove of any trees near unto the altar of the LORD thy God, which thou shalt make thee.
DEUT|16|22|Neither shalt thou set thee up any image; which the LORD thy God hateth.
DEUT|17|1|Thou shalt not sacrifice unto the LORD thy God any bullock, or sheep, wherein is blemish, or any evilfavouredness: for that is an abomination unto the LORD thy God.
DEUT|17|2|If there be found among you, within any of thy gates which the LORD thy God giveth thee, man or woman, that hath wrought wickedness in the sight of the LORD thy God, in transgressing his covenant,
DEUT|17|3|And hath gone and served other gods, and worshipped them, either the sun, or moon, or any of the host of heaven, which I have not commanded;
DEUT|17|4|And it be told thee, and thou hast heard of it, and inquired diligently, and, behold, it be true, and the thing certain, that such abomination is wrought in Israel:
DEUT|17|5|Then shalt thou bring forth that man or that woman, which have committed that wicked thing, unto thy gates, even that man or that woman, and shalt stone them with stones, till they die.
DEUT|17|6|At the mouth of two witnesses, or three witnesses, shall he that is worthy of death be put to death; but at the mouth of one witness he shall not be put to death.
DEUT|17|7|The hands of the witnesses shall be first upon him to put him to death, and afterward the hands of all the people. So thou shalt put the evil away from among you.
DEUT|17|8|If there arise a matter too hard for thee in judgment, between blood and blood, between plea and plea, and between stroke and stroke, being matters of controversy within thy gates: then shalt thou arise, and get thee up into the place which the LORD thy God shall choose;
DEUT|17|9|And thou shalt come unto the priests the Levites, and unto the judge that shall be in those days, and inquire; and they shall show thee the sentence of judgment:
DEUT|17|10|And thou shalt do according to the sentence, which they of that place which the LORD shall choose shall show thee; and thou shalt observe to do according to all that they inform thee:
DEUT|17|11|According to the sentence of the law which they shall teach thee, and according to the judgment which they shall tell thee, thou shalt do: thou shalt not decline from the sentence which they shall show thee, to the right hand, nor to the left.
DEUT|17|12|And the man that will do presumptuously, and will not hearken unto the priest that standeth to minister there before the LORD thy God, or unto the judge, even that man shall die: and thou shalt put away the evil from Israel.
DEUT|17|13|And all the people shall hear, and fear, and do no more presumptuously.
DEUT|17|14|When thou art come unto the land which the LORD thy God giveth thee, and shalt possess it, and shalt dwell therein, and shalt say, I will set a king over me, like as all the nations that are about me;
DEUT|17|15|Thou shalt in any wise set him king over thee, whom the LORD thy God shall choose: one from among thy brethren shalt thou set king over thee: thou mayest not set a stranger over thee, which is not thy brother.
DEUT|17|16|But he shall not multiply horses to himself, nor cause the people to return to Egypt, to the end that he should multiply horses: forasmuch as the LORD hath said unto you, Ye shall henceforth return no more that way.
DEUT|17|17|Neither shall he multiply wives to himself, that his heart turn not away: neither shall he greatly multiply to himself silver and gold.
DEUT|17|18|And it shall be, when he sitteth upon the throne of his kingdom, that he shall write him a copy of this law in a book out of that which is before the priests the Levites:
DEUT|17|19|And it shall be with him, and he shall read therein all the days of his life: that he may learn to fear the LORD his God, to keep all the words of this law and these statutes, to do them:
DEUT|17|20|That his heart be not lifted up above his brethren, and that he turn not aside from the commandment, to the right hand, or to the left: to the end that he may prolong his days in his kingdom, he, and his children, in the midst of Israel.
DEUT|18|1|The priests the Levites, and all the tribe of Levi, shall have no part nor inheritance with Israel: they shall eat the offerings of the LORD made by fire, and his inheritance.
DEUT|18|2|Therefore shall they have no inheritance among their brethren: the LORD is their inheritance, as he hath said unto them.
DEUT|18|3|And this shall be the priest's due from the people, from them that offer a sacrifice, whether it be ox or sheep; and they shall give unto the priest the shoulder, and the two cheeks, and the maw.
DEUT|18|4|The firstfruit also of thy corn, of thy wine, and of thine oil, and the first of the fleece of thy sheep, shalt thou give him.
DEUT|18|5|For the LORD thy God hath chosen him out of all thy tribes, to stand to minister in the name of the LORD, him and his sons for ever.
DEUT|18|6|And if a Levite come from any of thy gates out of all Israel, where he sojourned, and come with all the desire of his mind unto the place which the LORD shall choose;
DEUT|18|7|Then he shall minister in the name of the LORD his God, as all his brethren the Levites do, which stand there before the LORD.
DEUT|18|8|They shall have like portions to eat, beside that which cometh of the sale of his patrimony.
DEUT|18|9|When thou art come into the land which the LORD thy God giveth thee, thou shalt not learn to do after the abominations of those nations.
DEUT|18|10|There shall not be found among you any one that maketh his son or his daughter to pass through the fire, or that useth divination, or an observer of times, or an enchanter, or a witch.
DEUT|18|11|Or a charmer, or a consulter with familiar spirits, or a wizard, or a necromancer.
DEUT|18|12|For all that do these things are an abomination unto the LORD: and because of these abominations the LORD thy God doth drive them out from before thee.
DEUT|18|13|Thou shalt be perfect with the LORD thy God.
DEUT|18|14|For these nations, which thou shalt possess, hearkened unto observers of times, and unto diviners: but as for thee, the LORD thy God hath not suffered thee so to do.
DEUT|18|15|The LORD thy God will raise up unto thee a Prophet from the midst of thee, of thy brethren, like unto me; unto him ye shall hearken;
DEUT|18|16|According to all that thou desiredst of the LORD thy God in Horeb in the day of the assembly, saying, Let me not hear again the voice of the LORD my God, neither let me see this great fire any more, that I die not.
DEUT|18|17|And the LORD said unto me, They have well spoken that which they have spoken.
DEUT|18|18|I will raise them up a Prophet from among their brethren, like unto thee, and will put my words in his mouth; and he shall speak unto them all that I shall command him.
DEUT|18|19|And it shall come to pass, that whosoever will not hearken unto my words which he shall speak in my name, I will require it of him.
DEUT|18|20|But the prophet, which shall presume to speak a word in my name, which I have not commanded him to speak, or that shall speak in the name of other gods, even that prophet shall die.
DEUT|18|21|And if thou say in thine heart, How shall we know the word which the LORD hath not spoken?
DEUT|18|22|When a prophet speaketh in the name of the LORD, if the thing follow not, nor come to pass, that is the thing which the LORD hath not spoken, but the prophet hath spoken it presumptuously: thou shalt not be afraid of him.
DEUT|19|1|When the LORD thy God hath cut off the nations, whose land the LORD thy God giveth thee, and thou succeedest them, and dwellest in their cities, and in their houses;
DEUT|19|2|Thou shalt separate three cities for thee in the midst of thy land, which the LORD thy God giveth thee to possess it.
DEUT|19|3|Thou shalt prepare thee a way, and divide the coasts of thy land, which the LORD thy God giveth thee to inherit, into three parts, that every slayer may flee thither.
DEUT|19|4|And this is the case of the slayer, which shall flee thither, that he may live: Whoso killeth his neighbor ignorantly, whom he hated not in time past;
DEUT|19|5|As when a man goeth into the wood with his neighbor to hew wood, and his hand fetcheth a stroke with the axe to cut down the tree, and the head slippeth from the helve, and lighteth upon his neighbor, that he die; he shall flee unto one of those cities, and live:
DEUT|19|6|Lest the avenger of the blood pursue the slayer, while his heart is hot, and overtake him, because the way is long, and slay him; whereas he was not worthy of death, inasmuch as he hated him not in time past.
DEUT|19|7|Wherefore I command thee, saying, Thou shalt separate three cities for thee.
DEUT|19|8|And if the LORD thy God enlarge thy coast, as he hath sworn unto thy fathers, and give thee all the land which he promised to give unto thy fathers;
DEUT|19|9|If thou shalt keep all these commandments to do them, which I command thee this day, to love the LORD thy God, and to walk ever in his ways; then shalt thou add three cities more for thee, beside these three:
DEUT|19|10|That innocent blood be not shed in thy land, which the LORD thy God giveth thee for an inheritance, and so blood be upon thee.
DEUT|19|11|But if any man hate his neighbor, and lie in wait for him, and rise up against him, and smite him mortally that he die, and fleeth into one of these cities:
DEUT|19|12|Then the elders of his city shall send and fetch him thence, and deliver him into the hand of the avenger of blood, that he may die.
DEUT|19|13|Thine eye shall not pity him, but thou shalt put away the guilt of innocent blood from Israel, that it may go well with thee.
DEUT|19|14|Thou shalt not remove thy neighbor's landmark, which they of old time have set in thine inheritance, which thou shalt inherit in the land that the LORD thy God giveth thee to possess it.
DEUT|19|15|One witness shall not rise up against a man for any iniquity, or for any sin, in any sin that he sinneth: at the mouth of two witnesses, or at the mouth of three witnesses, shall the matter be established.
DEUT|19|16|If a false witness rise up against any man to testify against him that which is wrong;
DEUT|19|17|Then both the men, between whom the controversy is, shall stand before the LORD, before the priests and the judges, which shall be in those days;
DEUT|19|18|And the judges shall make diligent inquisition: and, behold, if the witness be a false witness, and hath testified falsely against his brother;
DEUT|19|19|Then shall ye do unto him, as he had thought to have done unto his brother: so shalt thou put the evil away from among you.
DEUT|19|20|And those which remain shall hear, and fear, and shall henceforth commit no more any such evil among you.
DEUT|19|21|And thine eye shall not pity; but life shall go for life, eye for eye, tooth for tooth, hand for hand, foot for foot.
DEUT|20|1|When thou goest out to battle against thine enemies, and seest horses, and chariots, and a people more than thou, be not afraid of them: for the LORD thy God is with thee, which brought thee up out of the land of Egypt.
DEUT|20|2|And it shall be, when ye are come nigh unto the battle, that the priest shall approach and speak unto the people,
DEUT|20|3|And shall say unto them, Hear, O Israel, ye approach this day unto battle against your enemies: let not your hearts faint, fear not, and do not tremble, neither be ye terrified because of them;
DEUT|20|4|For the LORD your God is he that goeth with you, to fight for you against your enemies, to save you.
DEUT|20|5|And the officers shall speak unto the people, saying, What man is there that hath built a new house, and hath not dedicated it? let him go and return to his house, lest he die in the battle, and another man dedicate it.
DEUT|20|6|And what man is he that hath planted a vineyard, and hath not yet eaten of it? let him also go and return unto his house, lest he die in the battle, and another man eat of it.
DEUT|20|7|And what man is there that hath betrothed a wife, and hath not taken her? let him go and return unto his house, lest he die in the battle, and another man take her.
DEUT|20|8|And the officers shall speak further unto the people, and they shall say, What man is there that is fearful and fainthearted? let him go and return unto his house, lest his brethren's heart faint as well as his heart.
DEUT|20|9|And it shall be, when the officers have made an end of speaking unto the people that they shall make captains of the armies to lead the people.
DEUT|20|10|When thou comest nigh unto a city to fight against it, then proclaim peace unto it.
DEUT|20|11|And it shall be, if it make thee answer of peace, and open unto thee, then it shall be, that all the people that is found therein shall be tributaries unto thee, and they shall serve thee.
DEUT|20|12|And if it will make no peace with thee, but will make war against thee, then thou shalt besiege it:
DEUT|20|13|And when the LORD thy God hath delivered it into thine hands, thou shalt smite every male thereof with the edge of the sword:
DEUT|20|14|But the women, and the little ones, and the cattle, and all that is in the city, even all the spoil thereof, shalt thou take unto thyself; and thou shalt eat the spoil of thine enemies, which the LORD thy God hath given thee.
DEUT|20|15|Thus shalt thou do unto all the cities which are very far off from thee, which are not of the cities of these nations.
DEUT|20|16|But of the cities of these people, which the LORD thy God doth give thee for an inheritance, thou shalt save alive nothing that breatheth:
DEUT|20|17|But thou shalt utterly destroy them; namely, the Hittites, and the Amorites, the Canaanites, and the Perizzites, the Hivites, and the Jebusites; as the LORD thy God hath commanded thee:
DEUT|20|18|That they teach you not to do after all their abominations, which they have done unto their gods; so should ye sin against the LORD your God.
DEUT|20|19|When thou shalt besiege a city a long time, in making war against it to take it, thou shalt not destroy the trees thereof by forcing an axe against them: for thou mayest eat of them, and thou shalt not cut them down (for the tree of the field is man's life) to employ them in the siege:
DEUT|20|20|Only the trees which thou knowest that they be not trees for meat, thou shalt destroy and cut them down; and thou shalt build bulwarks against the city that maketh war with thee, until it be subdued.
DEUT|21|1|If one be found slain in the land which the LORD thy God giveth thee to possess it, lying in the field, and it be not known who hath slain him:
DEUT|21|2|Then thy elders and thy judges shall come forth, and they shall measure unto the cities which are round about him that is slain:
DEUT|21|3|And it shall be, that the city which is next unto the slain man, even the elders of that city shall take an heifer, which hath not been wrought with, and which hath not drawn in the yoke;
DEUT|21|4|And the elders of that city shall bring down the heifer unto a rough valley, which is neither eared nor sown, and shall strike off the heifer's neck there in the valley:
DEUT|21|5|And the priests the sons of Levi shall come near; for them the LORD thy God hath chosen to minister unto him, and to bless in the name of the LORD; and by their word shall every controversy and every stroke be tried:
DEUT|21|6|And all the elders of that city, that are next unto the slain man, shall wash their hands over the heifer that is beheaded in the valley:
DEUT|21|7|And they shall answer and say, Our hands have not shed this blood, neither have our eyes seen it.
DEUT|21|8|Be merciful, O LORD, unto thy people Israel, whom thou hast redeemed, and lay not innocent blood unto thy people of Israel's charge. And the blood shall be forgiven them.
DEUT|21|9|So shalt thou put away the guilt of innocent blood from among you, when thou shalt do that which is right in the sight of the LORD.
DEUT|21|10|When thou goest forth to war against thine enemies, and the LORD thy God hath delivered them into thine hands, and thou hast taken them captive,
DEUT|21|11|And seest among the captives a beautiful woman, and hast a desire unto her, that thou wouldest have her to thy wife;
DEUT|21|12|Then thou shalt bring her home to thine house, and she shall shave her head, and pare her nails;
DEUT|21|13|And she shall put the raiment of her captivity from off her, and shall remain in thine house, and bewail her father and her mother a full month: and after that thou shalt go in unto her, and be her husband, and she shall be thy wife.
DEUT|21|14|And it shall be, if thou have no delight in her, then thou shalt let her go whither she will; but thou shalt not sell her at all for money, thou shalt not make merchandise of her, because thou hast humbled her.
DEUT|21|15|If a man have two wives, one beloved, and another hated, and they have born him children, both the beloved and the hated; and if the firstborn son be hers that was hated:
DEUT|21|16|Then it shall be, when he maketh his sons to inherit that which he hath, that he may not make the son of the beloved firstborn before the son of the hated, which is indeed the firstborn:
DEUT|21|17|But he shall acknowledge the son of the hated for the firstborn, by giving him a double portion of all that he hath: for he is the beginning of his strength; the right of the firstborn is his.
DEUT|21|18|If a man have a stubborn and rebellious son, which will not obey the voice of his father, or the voice of his mother, and that, when they have chastened him, will not hearken unto them:
DEUT|21|19|Then shall his father and his mother lay hold on him, and bring him out unto the elders of his city, and unto the gate of his place;
DEUT|21|20|And they shall say unto the elders of his city, This our son is stubborn and rebellious, he will not obey our voice; he is a glutton, and a drunkard.
DEUT|21|21|And all the men of his city shall stone him with stones, that he die: so shalt thou put evil away from among you; and all Israel shall hear, and fear.
DEUT|21|22|And if a man have committed a sin worthy of death, and he be to be put to death, and thou hang him on a tree:
DEUT|21|23|His body shall not remain all night upon the tree, but thou shalt in any wise bury him that day; (for he that is hanged is accursed of God;) that thy land be not defiled, which the LORD thy God giveth thee for an inheritance.
DEUT|22|1|Thou shalt not see thy brother's ox or his sheep go astray, and hide thyself from them: thou shalt in any case bring them again unto thy brother.
DEUT|22|2|And if thy brother be not nigh unto thee, or if thou know him not, then thou shalt bring it unto thine own house, and it shall be with thee until thy brother seek after it, and thou shalt restore it to him again.
DEUT|22|3|In like manner shalt thou do with his ass; and so shalt thou do with his raiment; and with all lost thing of thy brother's, which he hath lost, and thou hast found, shalt thou do likewise: thou mayest not hide thyself.
DEUT|22|4|Thou shalt not see thy brother's ass or his ox fall down by the way, and hide thyself from them: thou shalt surely help him to lift them up again.
DEUT|22|5|The woman shall not wear that which pertaineth unto a man, neither shall a man put on a woman's garment: for all that do so are abomination unto the LORD thy God.
DEUT|22|6|If a bird's nest chance to be before thee in the way in any tree, or on the ground, whether they be young ones, or eggs, and the dam sitting upon the young, or upon the eggs, thou shalt not take the dam with the young:
DEUT|22|7|But thou shalt in any wise let the dam go, and take the young to thee; that it may be well with thee, and that thou mayest prolong thy days.
DEUT|22|8|When thou buildest a new house, then thou shalt make a battlement for thy roof, that thou bring not blood upon thine house, if any man fall from thence.
DEUT|22|9|Thou shalt not sow thy vineyard with divers seeds: lest the fruit of thy seed which thou hast sown, and the fruit of thy vineyard, be defiled.
DEUT|22|10|Thou shalt not plow with an ox and an ass together.
DEUT|22|11|Thou shalt not wear a garment of divers sorts, as of woolen and linen together.
DEUT|22|12|Thou shalt make thee fringes upon the four quarters of thy vesture, wherewith thou coverest thyself.
DEUT|22|13|If any man take a wife, and go in unto her, and hate her,
DEUT|22|14|And give occasions of speech against her, and bring up an evil name upon her, and say, I took this woman, and when I came to her, I found her not a maid:
DEUT|22|15|Then shall the father of the damsel, and her mother, take and bring forth the tokens of the damsel's virginity unto the elders of the city in the gate:
DEUT|22|16|And the damsel's father shall say unto the elders, I gave my daughter unto this man to wife, and he hateth her;
DEUT|22|17|And, lo, he hath given occasions of speech against her, saying, I found not thy daughter a maid; and yet these are the tokens of my daughter's virginity. And they shall spread the cloth before the elders of the city.
DEUT|22|18|And the elders of that city shall take that man and chastise him;
DEUT|22|19|And they shall amerce him in an hundred shekels of silver, and give them unto the father of the damsel, because he hath brought up an evil name upon a virgin of Israel: and she shall be his wife; he may not put her away all his days.
DEUT|22|20|But if this thing be true, and the tokens of virginity be not found for the damsel:
DEUT|22|21|Then they shall bring out the damsel to the door of her father's house, and the men of her city shall stone her with stones that she die: because she hath wrought folly in Israel, to play the whore in her father's house: so shalt thou put evil away from among you.
DEUT|22|22|If a man be found lying with a woman married to an husband, then they shall both of them die, both the man that lay with the woman, and the woman: so shalt thou put away evil from Israel.
DEUT|22|23|If a damsel that is a virgin be betrothed unto an husband, and a man find her in the city, and lie with her;
DEUT|22|24|Then ye shall bring them both out unto the gate of that city, and ye shall stone them with stones that they die; the damsel, because she cried not, being in the city; and the man, because he hath humbled his neighbor's wife: so thou shalt put away evil from among you.
DEUT|22|25|But if a man find a betrothed damsel in the field, and the man force her, and lie with her: then the man only that lay with her shall die.
DEUT|22|26|But unto the damsel thou shalt do nothing; there is in the damsel no sin worthy of death: for as when a man riseth against his neighbor, and slayeth him, even so is this matter:
DEUT|22|27|For he found her in the field, and the betrothed damsel cried, and there was none to save her.
DEUT|22|28|If a man find a damsel that is a virgin, which is not betrothed, and lay hold on her, and lie with her, and they be found;
DEUT|22|29|Then the man that lay with her shall give unto the damsel's father fifty shekels of silver, and she shall be his wife; because he hath humbled her, he may not put her away all his days.
DEUT|22|30|A man shall not take his father's wife, nor discover his father's skirt.
DEUT|23|1|He that is wounded in the stones, or hath his privy member cut off, shall not enter into the congregation of the LORD.
DEUT|23|2|A bastard shall not enter into the congregation of the LORD; even to his tenth generation shall he not enter into the congregation of the LORD.
DEUT|23|3|An Ammonite or Moabite shall not enter into the congregation of the LORD; even to their tenth generation shall they not enter into the congregation of the LORD for ever:
DEUT|23|4|Because they met you not with bread and with water in the way, when ye came forth out of Egypt; and because they hired against thee Balaam the son of Beor of Pethor of Mesopotamia, to curse thee.
DEUT|23|5|Nevertheless the LORD thy God would not hearken unto Balaam; but the LORD thy God turned the curse into a blessing unto thee, because the LORD thy God loved thee.
DEUT|23|6|Thou shalt not seek their peace nor their prosperity all thy days for ever.
DEUT|23|7|Thou shalt not abhor an Edomite; for he is thy brother: thou shalt not abhor an Egyptian; because thou wast a stranger in his land.
DEUT|23|8|The children that are begotten of them shall enter into the congregation of the LORD in their third generation.
DEUT|23|9|When the host goeth forth against thine enemies, then keep thee from every wicked thing.
DEUT|23|10|If there be among you any man, that is not clean by reason of uncleanness that chanceth him by night, then shall he go abroad out of the camp, he shall not come within the camp:
DEUT|23|11|But it shall be, when evening cometh on, he shall wash himself with water: and when the sun is down, he shall come into the camp again.
DEUT|23|12|Thou shalt have a place also without the camp, whither thou shalt go forth abroad:
DEUT|23|13|And thou shalt have a paddle upon thy weapon; and it shall be, when thou wilt ease thyself abroad, thou shalt dig therewith, and shalt turn back and cover that which cometh from thee:
DEUT|23|14|For the LORD thy God walketh in the midst of thy camp, to deliver thee, and to give up thine enemies before thee; therefore shall thy camp be holy: that he see no unclean thing in thee, and turn away from thee.
DEUT|23|15|Thou shalt not deliver unto his master the servant which is escaped from his master unto thee:
DEUT|23|16|He shall dwell with thee, even among you, in that place which he shall choose in one of thy gates, where it liketh him best: thou shalt not oppress him.
DEUT|23|17|There shall be no whore of the daughters of Israel, nor a sodomite of the sons of Israel.
DEUT|23|18|Thou shalt not bring the hire of a whore, or the price of a dog, into the house of the LORD thy God for any vow: for even both these are abomination unto the LORD thy God.
DEUT|23|19|Thou shalt not lend upon usury to thy brother; usury of money, usury of victuals, usury of any thing that is lent upon usury:
DEUT|23|20|Unto a stranger thou mayest lend upon usury; but unto thy brother thou shalt not lend upon usury: that the LORD thy God may bless thee in all that thou settest thine hand to in the land whither thou goest to possess it.
DEUT|23|21|When thou shalt vow a vow unto the LORD thy God, thou shalt not slack to pay it: for the LORD thy God will surely require it of thee; and it would be sin in thee.
DEUT|23|22|But if thou shalt forbear to vow, it shall be no sin in thee.
DEUT|23|23|That which is gone out of thy lips thou shalt keep and perform; even a freewill offering, according as thou hast vowed unto the LORD thy God, which thou hast promised with thy mouth.
DEUT|23|24|When thou comest into thy neighbor's vineyard, then thou mayest eat grapes thy fill at thine own pleasure; but thou shalt not put any in thy vessel.
DEUT|23|25|When thou comest into the standing corn of thy neighbor, then thou mayest pluck the ears with thine hand; but thou shalt not move a sickle unto thy neighbor's standing corn.
DEUT|24|1|When a man hath taken a wife, and married her, and it come to pass that she find no favor in his eyes, because he hath found some uncleanness in her: then let him write her a bill of divorcement, and give it in her hand, and send her out of his house.
DEUT|24|2|And when she is departed out of his house, she may go and be another man's wife.
DEUT|24|3|And if the latter husband hate her, and write her a bill of divorcement, and giveth it in her hand, and sendeth her out of his house; or if the latter husband die, which took her to be his wife;
DEUT|24|4|Her former husband, which sent her away, may not take her again to be his wife, after that she is defiled; for that is abomination before the LORD: and thou shalt not cause the land to sin, which the LORD thy God giveth thee for an inheritance.
DEUT|24|5|When a man hath taken a new wife, he shall not go out to war, neither shall he be charged with any business: but he shall be free at home one year, and shall cheer up his wife which he hath taken.
DEUT|24|6|No man shall take the nether or the upper millstone to pledge: for he taketh a man's life to pledge.
DEUT|24|7|If a man be found stealing any of his brethren of the children of Israel, and maketh merchandise of him, or selleth him; then that thief shall die; and thou shalt put evil away from among you.
DEUT|24|8|Take heed in the plague of leprosy, that thou observe diligently, and do according to all that the priests the Levites shall teach you: as I commanded them, so ye shall observe to do.
DEUT|24|9|Remember what the LORD thy God did unto Miriam by the way, after that ye were come forth out of Egypt.
DEUT|24|10|When thou dost lend thy brother any thing, thou shalt not go into his house to fetch his pledge.
DEUT|24|11|Thou shalt stand abroad, and the man to whom thou dost lend shall bring out the pledge abroad unto thee.
DEUT|24|12|And if the man be poor, thou shalt not sleep with his pledge:
DEUT|24|13|In any case thou shalt deliver him the pledge again when the sun goeth down, that he may sleep in his own raiment, and bless thee: and it shall be righteousness unto thee before the LORD thy God.
DEUT|24|14|Thou shalt not oppress an hired servant that is poor and needy, whether he be of thy brethren, or of thy strangers that are in thy land within thy gates:
DEUT|24|15|At his day thou shalt give him his hire, neither shall the sun go down upon it; for he is poor, and setteth his heart upon it: lest he cry against thee unto the LORD, and it be sin unto thee.
DEUT|24|16|The fathers shall not be put to death for the children, neither shall the children be put to death for the fathers: every man shall be put to death for his own sin.
DEUT|24|17|Thou shalt not pervert the judgment of the stranger, nor of the fatherless; nor take a widow's raiment to pledge:
DEUT|24|18|But thou shalt remember that thou wast a bondman in Egypt, and the LORD thy God redeemed thee thence: therefore I command thee to do this thing.
DEUT|24|19|When thou cuttest down thine harvest in thy field, and hast forgot a sheaf in the field, thou shalt not go again to fetch it: it shall be for the stranger, for the fatherless, and for the widow: that the LORD thy God may bless thee in all the work of thine hands.
DEUT|24|20|When thou beatest thine olive tree, thou shalt not go over the boughs again: it shall be for the stranger, for the fatherless, and for the widow.
DEUT|24|21|When thou gatherest the grapes of thy vineyard, thou shalt not glean it afterward: it shall be for the stranger, for the fatherless, and for the widow.
DEUT|24|22|And thou shalt remember that thou wast a bondman in the land of Egypt: therefore I command thee to do this thing.
DEUT|25|1|If there be a controversy between men, and they come unto judgment, that the judges may judge them; then they shall justify the righteous, and condemn the wicked.
DEUT|25|2|And it shall be, if the wicked man be worthy to be beaten, that the judge shall cause him to lie down, and to be beaten before his face, according to his fault, by a certain number.
DEUT|25|3|Forty stripes he may give him, and not exceed: lest, if he should exceed, and beat him above these with many stripes, then thy brother should seem vile unto thee.
DEUT|25|4|Thou shalt not muzzle the ox when he treadeth out the corn.
DEUT|25|5|If brethren dwell together, and one of them die, and have no child, the wife of the dead shall not marry without unto a stranger: her husband's brother shall go in unto her, and take her to him to wife, and perform the duty of an husband's brother unto her.
DEUT|25|6|And it shall be, that the firstborn which she beareth shall succeed in the name of his brother which is dead, that his name be not put out of Israel.
DEUT|25|7|And if the man like not to take his brother's wife, then let his brother's wife go up to the gate unto the elders, and say, My husband's brother refuseth to raise up unto his brother a name in Israel, he will not perform the duty of my husband's brother.
DEUT|25|8|Then the elders of his city shall call him, and speak unto him: and if he stand to it, and say, I like not to take her;
DEUT|25|9|Then shall his brother's wife come unto him in the presence of the elders, and loose his shoe from off his foot, and spit in his face, and shall answer and say, So shall it be done unto that man that will not build up his brother's house.
DEUT|25|10|And his name shall be called in Israel, The house of him that hath his shoe loosed.
DEUT|25|11|When men strive together one with another, and the wife of the one draweth near for to deliver her husband out of the hand of him that smiteth him, and putteth forth her hand, and taketh him by the secrets:
DEUT|25|12|Then thou shalt cut off her hand, thine eye shall not pity her.
DEUT|25|13|Thou shalt not have in thy bag divers weights, a great and a small.
DEUT|25|14|Thou shalt not have in thine house divers measures, a great and a small.
DEUT|25|15|But thou shalt have a perfect and just weight, a perfect and just measure shalt thou have: that thy days may be lengthened in the land which the LORD thy God giveth thee.
DEUT|25|16|For all that do such things, and all that do unrighteously, are an abomination unto the LORD thy God.
DEUT|25|17|Remember what Amalek did unto thee by the way, when ye were come forth out of Egypt;
DEUT|25|18|How he met thee by the way, and smote the hindmost of thee, even all that were feeble behind thee, when thou wast faint and weary; and he feared not God.
DEUT|25|19|Therefore it shall be, when the LORD thy God hath given thee rest from all thine enemies round about, in the land which the LORD thy God giveth thee for an inheritance to possess it, that thou shalt blot out the remembrance of Amalek from under heaven; thou shalt not forget it.
DEUT|26|1|And it shall be, when thou art come in unto the land which the LORD thy God giveth thee for an inheritance, and possessest it, and dwellest therein;
DEUT|26|2|That thou shalt take of the first of all the fruit of the earth, which thou shalt bring of thy land that the LORD thy God giveth thee, and shalt put it in a basket, and shalt go unto the place which the LORD thy God shall choose to place his name there.
DEUT|26|3|And thou shalt go unto the priest that shall be in those days, and say unto him, I profess this day unto the LORD thy God, that I am come unto the country which the LORD sware unto our fathers for to give us.
DEUT|26|4|And the priest shall take the basket out of thine hand, and set it down before the altar of the LORD thy God.
DEUT|26|5|And thou shalt speak and say before the LORD thy God, A Syrian ready to perish was my father, and he went down into Egypt, and sojourned there with a few, and became there a nation, great, mighty, and populous:
DEUT|26|6|And the Egyptians evil entreated us, and afflicted us, and laid upon us hard bondage:
DEUT|26|7|And when we cried unto the LORD God of our fathers, the LORD heard our voice, and looked on our affliction, and our labor, and our oppression:
DEUT|26|8|And the LORD brought us forth out of Egypt with a mighty hand, and with an outstretched arm, and with great terribleness, and with signs, and with wonders:
DEUT|26|9|And he hath brought us into this place, and hath given us this land, even a land that floweth with milk and honey.
DEUT|26|10|And now, behold, I have brought the firstfruits of the land, which thou, O LORD, hast given me. And thou shalt set it before the LORD thy God, and worship before the LORD thy God:
DEUT|26|11|And thou shalt rejoice in every good thing which the LORD thy God hath given unto thee, and unto thine house, thou, and the Levite, and the stranger that is among you.
DEUT|26|12|When thou hast made an end of tithing all the tithes of thine increase the third year, which is the year of tithing, and hast given it unto the Levite, the stranger, the fatherless, and the widow, that they may eat within thy gates, and be filled;
DEUT|26|13|Then thou shalt say before the LORD thy God, I have brought away the hallowed things out of mine house, and also have given them unto the Levite, and unto the stranger, to the fatherless, and to the widow, according to all thy commandments which thou hast commanded me: I have not transgressed thy commandments, neither have I forgotten them.
DEUT|26|14|I have not eaten thereof in my mourning, neither have I taken away ought thereof for any unclean use, nor given ought thereof for the dead: but I have hearkened to the voice of the LORD my God, and have done according to all that thou hast commanded me.
DEUT|26|15|Look down from thy holy habitation, from heaven, and bless thy people Israel, and the land which thou hast given us, as thou swarest unto our fathers, a land that floweth with milk and honey.
DEUT|26|16|This day the LORD thy God hath commanded thee to do these statutes and judgments: thou shalt therefore keep and do them with all thine heart, and with all thy soul.
DEUT|26|17|Thou hast avouched the LORD this day to be thy God, and to walk in his ways, and to keep his statutes, and his commandments, and his judgments, and to hearken unto his voice:
DEUT|26|18|And the LORD hath avouched thee this day to be his peculiar people, as he hath promised thee, and that thou shouldest keep all his commandments;
DEUT|26|19|And to make thee high above all nations which he hath made, in praise, and in name, and in honor; and that thou mayest be an holy people unto the LORD thy God, as he hath spoken.
DEUT|27|1|And Moses with the elders of Israel commanded the people, saying, Keep all the commandments which I command you this day.
DEUT|27|2|And it shall be on the day when ye shall pass over Jordan unto the land which the LORD thy God giveth thee, that thou shalt set thee up great stones, and plaster them with plaster:
DEUT|27|3|And thou shalt write upon them all the words of this law, when thou art passed over, that thou mayest go in unto the land which the LORD thy God giveth thee, a land that floweth with milk and honey; as the LORD God of thy fathers hath promised thee.
DEUT|27|4|Therefore it shall be when ye be gone over Jordan, that ye shall set up these stones, which I command you this day, in mount Ebal, and thou shalt plaster them with plaster.
DEUT|27|5|And there shalt thou build an altar unto the LORD thy God, an altar of stones: thou shalt not lift up any iron tool upon them.
DEUT|27|6|Thou shalt build the altar of the LORD thy God of whole stones: and thou shalt offer burnt offerings thereon unto the LORD thy God:
DEUT|27|7|And thou shalt offer peace offerings, and shalt eat there, and rejoice before the LORD thy God.
DEUT|27|8|And thou shalt write upon the stones all the words of this law very plainly.
DEUT|27|9|And Moses and the priests the Levites spake unto all Israel, saying, Take heed, and hearken, O Israel; this day thou art become the people of the LORD thy God.
DEUT|27|10|Thou shalt therefore obey the voice of the LORD thy God, and do his commandments and his statutes, which I command thee this day.
DEUT|27|11|And Moses charged the people the same day, saying,
DEUT|27|12|These shall stand upon mount Gerizim to bless the people, when ye are come over Jordan; Simeon, and Levi, and Judah, and Issachar, and Joseph, and Benjamin:
DEUT|27|13|And these shall stand upon mount Ebal to curse; Reuben, Gad, and Asher, and Zebulun, Dan, and Naphtali.
DEUT|27|14|And the Levites shall speak, and say unto all the men of Israel with a loud voice,
DEUT|27|15|Cursed be the man that maketh any graven or molten image, an abomination unto the LORD, the work of the hands of the craftsman, and putteth it in a secret place. And all the people shall answer and say, Amen.
DEUT|27|16|Cursed be he that setteth light by his father or his mother. And all the people shall say, Amen.
DEUT|27|17|Cursed be he that removeth his neighbor's landmark. And all the people shall say, Amen.
DEUT|27|18|Cursed be he that maketh the blind to wander out of the way. And all the people shall say, Amen.
DEUT|27|19|Cursed be he that perverteth the judgment of the stranger, fatherless, and widow. And all the people shall say, Amen.
DEUT|27|20|Cursed be he that lieth with his father's wife; because he uncovereth his father's skirt. And all the people shall say, Amen.
DEUT|27|21|Cursed be he that lieth with any manner of beast. And all the people shall say, Amen.
DEUT|27|22|Cursed be he that lieth with his sister, the daughter of his father, or the daughter of his mother. And all the people shall say, Amen.
DEUT|27|23|Cursed be he that lieth with his mother in law. And all the people shall say, Amen.
DEUT|27|24|Cursed be he that smiteth his neighbor secretly. And all the people shall say, Amen.
DEUT|27|25|Cursed be he that taketh reward to slay an innocent person. And all the people shall say, Amen.
DEUT|27|26|Cursed be he that confirmeth not all the words of this law to do them. And all the people shall say, Amen.
DEUT|28|1|And it shall come to pass, if thou shalt hearken diligently unto the voice of the LORD thy God, to observe and to do all his commandments which I command thee this day, that the LORD thy God will set thee on high above all nations of the earth:
DEUT|28|2|And all these blessings shall come on thee, and overtake thee, if thou shalt hearken unto the voice of the LORD thy God.
DEUT|28|3|Blessed shalt thou be in the city, and blessed shalt thou be in the field.
DEUT|28|4|Blessed shall be the fruit of thy body, and the fruit of thy ground, and the fruit of thy cattle, the increase of thy kine, and the flocks of thy sheep.
DEUT|28|5|Blessed shall be thy basket and thy store.
DEUT|28|6|Blessed shalt thou be when thou comest in, and blessed shalt thou be when thou goest out.
DEUT|28|7|The LORD shall cause thine enemies that rise up against thee to be smitten before thy face: they shall come out against thee one way, and flee before thee seven ways.
DEUT|28|8|The LORD shall command the blessing upon thee in thy storehouses, and in all that thou settest thine hand unto; and he shall bless thee in the land which the LORD thy God giveth thee.
DEUT|28|9|The LORD shall establish thee an holy people unto himself, as he hath sworn unto thee, if thou shalt keep the commandments of the LORD thy God, and walk in his ways.
DEUT|28|10|And all people of the earth shall see that thou art called by the name of the LORD; and they shall be afraid of thee.
DEUT|28|11|And the LORD shall make thee plenteous in goods, in the fruit of thy body, and in the fruit of thy cattle, and in the fruit of thy ground, in the land which the LORD sware unto thy fathers to give thee.
DEUT|28|12|The LORD shall open unto thee his good treasure, the heaven to give the rain unto thy land in his season, and to bless all the work of thine hand: and thou shalt lend unto many nations, and thou shalt not borrow.
DEUT|28|13|And the LORD shall make thee the head, and not the tail; and thou shalt be above only, and thou shalt not be beneath; if that thou hearken unto the commandments of the LORD thy God, which I command thee this day, to observe and to do them:
DEUT|28|14|And thou shalt not go aside from any of the words which I command thee this day, to the right hand, or to the left, to go after other gods to serve them.
DEUT|28|15|But it shall come to pass, if thou wilt not hearken unto the voice of the LORD thy God, to observe to do all his commandments and his statutes which I command thee this day; that all these curses shall come upon thee, and overtake thee:
DEUT|28|16|Cursed shalt thou be in the city, and cursed shalt thou be in the field.
DEUT|28|17|Cursed shall be thy basket and thy store.
DEUT|28|18|Cursed shall be the fruit of thy body, and the fruit of thy land, the increase of thy kine, and the flocks of thy sheep.
DEUT|28|19|Cursed shalt thou be when thou comest in, and cursed shalt thou be when thou goest out.
DEUT|28|20|The LORD shall send upon thee cursing, vexation, and rebuke, in all that thou settest thine hand unto for to do, until thou be destroyed, and until thou perish quickly; because of the wickedness of thy doings, whereby thou hast forsaken me.
DEUT|28|21|The LORD shall make the pestilence cleave unto thee, until he have consumed thee from off the land, whither thou goest to possess it.
DEUT|28|22|The LORD shall smite thee with a consumption, and with a fever, and with an inflammation, and with an extreme burning, and with the sword, and with blasting, and with mildew; and they shall pursue thee until thou perish.
DEUT|28|23|And thy heaven that is over thy head shall be brass, and the earth that is under thee shall be iron.
DEUT|28|24|The LORD shall make the rain of thy land powder and dust: from heaven shall it come down upon thee, until thou be destroyed.
DEUT|28|25|The LORD shall cause thee to be smitten before thine enemies: thou shalt go out one way against them, and flee seven ways before them: and shalt be removed into all the kingdoms of the earth.
DEUT|28|26|And thy carcass shall be meat unto all fowls of the air, and unto the beasts of the earth, and no man shall fray them away.
DEUT|28|27|The LORD will smite thee with the botch of Egypt, and with the emerods, and with the scab, and with the itch, whereof thou canst not be healed.
DEUT|28|28|The LORD shall smite thee with madness, and blindness, and astonishment of heart:
DEUT|28|29|And thou shalt grope at noonday, as the blind gropeth in darkness, and thou shalt not prosper in thy ways: and thou shalt be only oppressed and spoiled evermore, and no man shall save thee.
DEUT|28|30|Thou shalt betroth a wife, and another man shall lie with her: thou shalt build an house, and thou shalt not dwell therein: thou shalt plant a vineyard, and shalt not gather the grapes thereof.
DEUT|28|31|Thine ox shall be slain before thine eyes, and thou shalt not eat thereof: thine ass shall be violently taken away from before thy face, and shall not be restored to thee: thy sheep shall be given unto thine enemies, and thou shalt have none to rescue them.
DEUT|28|32|Thy sons and thy daughters shall be given unto another people, and thine eyes shall look, and fail with longing for them all the day long; and there shall be no might in thine hand.
DEUT|28|33|The fruit of thy land, and all thy labors, shall a nation which thou knowest not eat up; and thou shalt be only oppressed and crushed alway:
DEUT|28|34|So that thou shalt be mad for the sight of thine eyes which thou shalt see.
DEUT|28|35|The LORD shall smite thee in the knees, and in the legs, with a sore botch that cannot be healed, from the sole of thy foot unto the top of thy head.
DEUT|28|36|The LORD shall bring thee, and thy king which thou shalt set over thee, unto a nation which neither thou nor thy fathers have known; and there shalt thou serve other gods, wood and stone.
DEUT|28|37|And thou shalt become an astonishment, a proverb, and a byword, among all nations whither the LORD shall lead thee.
DEUT|28|38|Thou shalt carry much seed out into the field, and shalt gather but little in; for the locust shall consume it.
DEUT|28|39|Thou shalt plant vineyards, and dress them, but shalt neither drink of the wine, nor gather the grapes; for the worms shall eat them.
DEUT|28|40|Thou shalt have olive trees throughout all thy coasts, but thou shalt not anoint thyself with the oil; for thine olive shall cast his fruit.
DEUT|28|41|Thou shalt beget sons and daughters, but thou shalt not enjoy them; for they shall go into captivity.
DEUT|28|42|All thy trees and fruit of thy land shall the locust consume.
DEUT|28|43|The stranger that is within thee shall get up above thee very high; and thou shalt come down very low.
DEUT|28|44|He shall lend to thee, and thou shalt not lend to him: he shall be the head, and thou shalt be the tail.
DEUT|28|45|Moreover all these curses shall come upon thee, and shall pursue thee, and overtake thee, till thou be destroyed; because thou hearkenedst not unto the voice of the LORD thy God, to keep his commandments and his statutes which he commanded thee:
DEUT|28|46|And they shall be upon thee for a sign and for a wonder, and upon thy seed for ever.
DEUT|28|47|Because thou servedst not the LORD thy God with joyfulness, and with gladness of heart, for the abundance of all things;
DEUT|28|48|Therefore shalt thou serve thine enemies which the LORD shall send against thee, in hunger, and in thirst, and in nakedness, and in want of all things: and he shall put a yoke of iron upon thy neck, until he have destroyed thee.
DEUT|28|49|The LORD shall bring a nation against thee from far, from the end of the earth, as swift as the eagle flieth; a nation whose tongue thou shalt not understand;
DEUT|28|50|A nation of fierce countenance, which shall not regard the person of the old, nor show favor to the young:
DEUT|28|51|And he shall eat the fruit of thy cattle, and the fruit of thy land, until thou be destroyed: which also shall not leave thee either corn, wine, or oil, or the increase of thy kine, or flocks of thy sheep, until he have destroyed thee.
DEUT|28|52|And he shall besiege thee in all thy gates, until thy high and fenced walls come down, wherein thou trustedst, throughout all thy land: and he shall besiege thee in all thy gates throughout all thy land, which the LORD thy God hath given thee.
DEUT|28|53|And thou shalt eat the fruit of thine own body, the flesh of thy sons and of thy daughters, which the LORD thy God hath given thee, in the siege, and in the straitness, wherewith thine enemies shall distress thee:
DEUT|28|54|So that the man that is tender among you, and very delicate, his eye shall be evil toward his brother, and toward the wife of his bosom, and toward the remnant of his children which he shall leave:
DEUT|28|55|So that he will not give to any of them of the flesh of his children whom he shall eat: because he hath nothing left him in the siege, and in the straitness, wherewith thine enemies shall distress thee in all thy gates.
DEUT|28|56|The tender and delicate woman among you, which would not adventure to set the sole of her foot upon the ground for delicateness and tenderness, her eye shall be evil toward the husband of her bosom, and toward her son, and toward her daughter,
DEUT|28|57|And toward her young one that cometh out from between her feet, and toward her children which she shall bear: for she shall eat them for want of all things secretly in the siege and straitness, wherewith thine enemy shall distress thee in thy gates.
DEUT|28|58|If thou wilt not observe to do all the words of this law that are written in this book, that thou mayest fear this glorious and fearful name, THE LORD THY GOD;
DEUT|28|59|Then the LORD will make thy plagues wonderful, and the plagues of thy seed, even great plagues, and of long continuance, and sore sicknesses, and of long continuance.
DEUT|28|60|Moreover he will bring upon thee all the diseases of Egypt, which thou wast afraid of; and they shall cleave unto thee.
DEUT|28|61|Also every sickness, and every plague, which is not written in the book of this law, them will the LORD bring upon thee, until thou be destroyed.
DEUT|28|62|And ye shall be left few in number, whereas ye were as the stars of heaven for multitude; because thou wouldest not obey the voice of the LORD thy God.
DEUT|28|63|And it shall come to pass, that as the LORD rejoiced over you to do you good, and to multiply you; so the LORD will rejoice over you to destroy you, and to bring you to nought; and ye shall be plucked from off the land whither thou goest to possess it.
DEUT|28|64|And the LORD shall scatter thee among all people, from the one end of the earth even unto the other; and there thou shalt serve other gods, which neither thou nor thy fathers have known, even wood and stone.
DEUT|28|65|And among these nations shalt thou find no ease, neither shall the sole of thy foot have rest: but the LORD shall give thee there a trembling heart, and failing of eyes, and sorrow of mind:
DEUT|28|66|And thy life shall hang in doubt before thee; and thou shalt fear day and night, and shalt have none assurance of thy life:
DEUT|28|67|In the morning thou shalt say, Would God it were even! and at even thou shalt say, Would God it were morning! for the fear of thine heart wherewith thou shalt fear, and for the sight of thine eyes which thou shalt see.
DEUT|28|68|And the LORD shall bring thee into Egypt again with ships, by the way whereof I spake unto thee, Thou shalt see it no more again: and there ye shall be sold unto your enemies for bondmen and bondwomen, and no man shall buy you.
DEUT|29|1|These are the words of the covenant, which the LORD commanded Moses to make with the children of Israel in the land of Moab, beside the covenant which he made with them in Horeb.
DEUT|29|2|And Moses called unto all Israel, and said unto them, Ye have seen all that the LORD did before your eyes in the land of Egypt unto Pharaoh, and unto all his servants, and unto all his land;
DEUT|29|3|The great temptations which thine eyes have seen, the signs, and those great miracles:
DEUT|29|4|Yet the LORD hath not given you an heart to perceive, and eyes to see, and ears to hear, unto this day.
DEUT|29|5|And I have led you forty years in the wilderness: your clothes are not waxen old upon you, and thy shoe is not waxen old upon thy foot.
DEUT|29|6|Ye have not eaten bread, neither have ye drunk wine or strong drink: that ye might know that I am the LORD your God.
DEUT|29|7|And when ye came unto this place, Sihon the king of Heshbon, and Og the king of Bashan, came out against us unto battle, and we smote them:
DEUT|29|8|And we took their land, and gave it for an inheritance unto the Reubenites, and to the Gadites, and to the half tribe of Manasseh.
DEUT|29|9|Keep therefore the words of this covenant, and do them, that ye may prosper in all that ye do.
DEUT|29|10|Ye stand this day all of you before the LORD your God; your captains of your tribes, your elders, and your officers, with all the men of Israel,
DEUT|29|11|Your little ones, your wives, and thy stranger that is in thy camp, from the hewer of thy wood unto the drawer of thy water:
DEUT|29|12|That thou shouldest enter into covenant with the LORD thy God, and into his oath, which the LORD thy God maketh with thee this day:
DEUT|29|13|That he may establish thee to day for a people unto himself, and that he may be unto thee a God, as he hath said unto thee, and as he hath sworn unto thy fathers, to Abraham, to Isaac, and to Jacob.
DEUT|29|14|Neither with you only do I make this covenant and this oath;
DEUT|29|15|But with him that standeth here with us this day before the LORD our God, and also with him that is not here with us this day:
DEUT|29|16|(For ye know how we have dwelt in the land of Egypt; and how we came through the nations which ye passed by;
DEUT|29|17|And ye have seen their abominations, and their idols, wood and stone, silver and gold, which were among them:)
DEUT|29|18|Lest there should be among you man, or woman, or family, or tribe, whose heart turneth away this day from the LORD our God, to go and serve the gods of these nations; lest there should be among you a root that beareth gall and wormwood;
DEUT|29|19|And it come to pass, when he heareth the words of this curse, that he bless himself in his heart, saying, I shall have peace, though I walk in the imagination of mine heart, to add drunkenness to thirst:
DEUT|29|20|The LORD will not spare him, but then the anger of the LORD and his jealousy shall smoke against that man, and all the curses that are written in this book shall lie upon him, and the LORD shall blot out his name from under heaven.
DEUT|29|21|And the LORD shall separate him unto evil out of all the tribes of Israel, according to all the curses of the covenant that are written in this book of the law:
DEUT|29|22|So that the generation to come of your children that shall rise up after you, and the stranger that shall come from a far land, shall say, when they see the plagues of that land, and the sicknesses which the LORD hath laid upon it;
DEUT|29|23|And that the whole land thereof is brimstone, and salt, and burning, that it is not sown, nor beareth, nor any grass groweth therein, like the overthrow of Sodom, and Gomorrah, Admah, and Zeboim, which the LORD overthrew in his anger, and in his wrath:
DEUT|29|24|Even all nations shall say, Wherefore hath the LORD done thus unto this land? what meaneth the heat of this great anger?
DEUT|29|25|Then men shall say, Because they have forsaken the covenant of the LORD God of their fathers, which he made with them when he brought them forth out of the land of Egypt:
DEUT|29|26|For they went and served other gods, and worshipped them, gods whom they knew not, and whom he had not given unto them:
DEUT|29|27|And the anger of the LORD was kindled against this land, to bring upon it all the curses that are written in this book:
DEUT|29|28|And the LORD rooted them out of their land in anger, and in wrath, and in great indignation, and cast them into another land, as it is this day.
DEUT|29|29|The secret things belong unto the LORD our God: but those things which are revealed belong unto us and to our children for ever, that we may do all the words of this law.
DEUT|30|1|And it shall come to pass, when all these things are come upon thee, the blessing and the curse, which I have set before thee, and thou shalt call them to mind among all the nations, whither the LORD thy God hath driven thee,
DEUT|30|2|And shalt return unto the LORD thy God, and shalt obey his voice according to all that I command thee this day, thou and thy children, with all thine heart, and with all thy soul;
DEUT|30|3|That then the LORD thy God will turn thy captivity, and have compassion upon thee, and will return and gather thee from all the nations, whither the LORD thy God hath scattered thee.
DEUT|30|4|If any of thine be driven out unto the outmost parts of heaven, from thence will the LORD thy God gather thee, and from thence will he fetch thee:
DEUT|30|5|And the LORD thy God will bring thee into the land which thy fathers possessed, and thou shalt possess it; and he will do thee good, and multiply thee above thy fathers.
DEUT|30|6|And the LORD thy God will circumcise thine heart, and the heart of thy seed, to love the LORD thy God with all thine heart, and with all thy soul, that thou mayest live.
DEUT|30|7|And the LORD thy God will put all these curses upon thine enemies, and on them that hate thee, which persecuted thee.
DEUT|30|8|And thou shalt return and obey the voice of the LORD, and do all his commandments which I command thee this day.
DEUT|30|9|And the LORD thy God will make thee plenteous in every work of thine hand, in the fruit of thy body, and in the fruit of thy cattle, and in the fruit of thy land, for good: for the LORD will again rejoice over thee for good, as he rejoiced over thy fathers:
DEUT|30|10|If thou shalt hearken unto the voice of the LORD thy God, to keep his commandments and his statutes which are written in this book of the law, and if thou turn unto the LORD thy God with all thine heart, and with all thy soul.
DEUT|30|11|For this commandment which I command thee this day, it is not hidden from thee, neither is it far off.
DEUT|30|12|It is not in heaven, that thou shouldest say, Who shall go up for us to heaven, and bring it unto us, that we may hear it, and do it?
DEUT|30|13|Neither is it beyond the sea, that thou shouldest say, Who shall go over the sea for us, and bring it unto us, that we may hear it, and do it?
DEUT|30|14|But the word is very nigh unto thee, in thy mouth, and in thy heart, that thou mayest do it.
DEUT|30|15|See, I have set before thee this day life and good, and death and evil;
DEUT|30|16|In that I command thee this day to love the LORD thy God, to walk in his ways, and to keep his commandments and his statutes and his judgments, that thou mayest live and multiply: and the LORD thy God shall bless thee in the land whither thou goest to possess it.
DEUT|30|17|But if thine heart turn away, so that thou wilt not hear, but shalt be drawn away, and worship other gods, and serve them;
DEUT|30|18|I denounce unto you this day, that ye shall surely perish, and that ye shall not prolong your days upon the land, whither thou passest over Jordan to go to possess it.
DEUT|30|19|I call heaven and earth to record this day against you, that I have set before you life and death, blessing and cursing: therefore choose life, that both thou and thy seed may live:
DEUT|30|20|That thou mayest love the LORD thy God, and that thou mayest obey his voice, and that thou mayest cleave unto him: for he is thy life, and the length of thy days: that thou mayest dwell in the land which the LORD sware unto thy fathers, to Abraham, to Isaac, and to Jacob, to give them.
DEUT|31|1|And Moses went and spake these words unto all Israel.
DEUT|31|2|And he said unto them, I am an hundred and twenty years old this day; I can no more go out and come in: also the LORD hath said unto me, Thou shalt not go over this Jordan.
DEUT|31|3|The LORD thy God, he will go over before thee, and he will destroy these nations from before thee, and thou shalt possess them: and Joshua, he shall go over before thee, as the LORD hath said.
DEUT|31|4|And the LORD shall do unto them as he did to Sihon and to Og, kings of the Amorites, and unto the land of them, whom he destroyed.
DEUT|31|5|And the LORD shall give them up before your face, that ye may do unto them according unto all the commandments which I have commanded you.
DEUT|31|6|Be strong and of a good courage, fear not, nor be afraid of them: for the LORD thy God, he it is that doth go with thee; he will not fail thee, nor forsake thee.
DEUT|31|7|And Moses called unto Joshua, and said unto him in the sight of all Israel, Be strong and of a good courage: for thou must go with this people unto the land which the LORD hath sworn unto their fathers to give them; and thou shalt cause them to inherit it.
DEUT|31|8|And the LORD, he it is that doth go before thee; he will be with thee, he will not fail thee, neither forsake thee: fear not, neither be dismayed.
DEUT|31|9|And Moses wrote this law, and delivered it unto the priests the sons of Levi, which bare the ark of the covenant of the LORD, and unto all the elders of Israel.
DEUT|31|10|And Moses commanded them, saying, At the end of every seven years, in the solemnity of the year of release, in the feast of tabernacles,
DEUT|31|11|When all Israel is come to appear before the LORD thy God in the place which he shall choose, thou shalt read this law before all Israel in their hearing.
DEUT|31|12|Gather the people together, men and women, and children, and thy stranger that is within thy gates, that they may hear, and that they may learn, and fear the LORD your God, and observe to do all the words of this law:
DEUT|31|13|And that their children, which have not known any thing, may hear, and learn to fear the LORD your God, as long as ye live in the land whither ye go over Jordan to possess it.
DEUT|31|14|And the LORD said unto Moses, Behold, thy days approach that thou must die: call Joshua, and present yourselves in the tabernacle of the congregation, that I may give him a charge. And Moses and Joshua went, and presented themselves in the tabernacle of the congregation.
DEUT|31|15|And the LORD appeared in the tabernacle in a pillar of a cloud: and the pillar of the cloud stood over the door of the tabernacle.
DEUT|31|16|And the LORD said unto Moses, Behold, thou shalt sleep with thy fathers; and this people will rise up, and go a whoring after the gods of the strangers of the land, whither they go to be among them, and will forsake me, and break my covenant which I have made with them.
DEUT|31|17|Then my anger shall be kindled against them in that day, and I will forsake them, and I will hide my face from them, and they shall be devoured, and many evils and troubles shall befall them; so that they will say in that day, Are not these evils come upon us, because our God is not among us?
DEUT|31|18|And I will surely hide my face in that day for all the evils which they shall have wrought, in that they are turned unto other gods.
DEUT|31|19|Now therefore write ye this song for you, and teach it the children of Israel: put it in their mouths, that this song may be a witness for me against the children of Israel.
DEUT|31|20|For when I shall have brought them into the land which I sware unto their fathers, that floweth with milk and honey; and they shall have eaten and filled themselves, and waxen fat; then will they turn unto other gods, and serve them, and provoke me, and break my covenant.
DEUT|31|21|And it shall come to pass, when many evils and troubles are befallen them, that this song shall testify against them as a witness; for it shall not be forgotten out of the mouths of their seed: for I know their imagination which they go about, even now, before I have brought them into the land which I sware.
DEUT|31|22|Moses therefore wrote this song the same day, and taught it the children of Israel.
DEUT|31|23|And he gave Joshua the son of Nun a charge, and said, Be strong and of a good courage: for thou shalt bring the children of Israel into the land which I sware unto them: and I will be with thee.
DEUT|31|24|And it came to pass, when Moses had made an end of writing the words of this law in a book, until they were finished,
DEUT|31|25|That Moses commanded the Levites, which bare the ark of the covenant of the LORD, saying,
DEUT|31|26|Take this book of the law, and put it in the side of the ark of the covenant of the LORD your God, that it may be there for a witness against thee.
DEUT|31|27|For I know thy rebellion, and thy stiff neck: behold, while I am yet alive with you this day, ye have been rebellious against the LORD; and how much more after my death?
DEUT|31|28|Gather unto me all the elders of your tribes, and your officers, that I may speak these words in their ears, and call heaven and earth to record against them.
DEUT|31|29|For I know that after my death ye will utterly corrupt yourselves, and turn aside from the way which I have commanded you; and evil will befall you in the latter days; because ye will do evil in the sight of the LORD, to provoke him to anger through the work of your hands.
DEUT|31|30|And Moses spake in the ears of all the congregation of Israel the words of this song, until they were ended.
DEUT|32|1|Give ear, O ye heavens, and I will speak; and hear, O earth, the words of my mouth.
DEUT|32|2|My doctrine shall drop as the rain, my speech shall distil as the dew, as the small rain upon the tender herb, and as the showers upon the grass:
DEUT|32|3|Because I will publish the name of the LORD: ascribe ye greatness unto our God.
DEUT|32|4|He is the Rock, his work is perfect: for all his ways are judgment: a God of truth and without iniquity, just and right is he.
DEUT|32|5|They have corrupted themselves, their spot is not the spot of his children: they are a perverse and crooked generation.
DEUT|32|6|Do ye thus requite the LORD, O foolish people and unwise? is not he thy father that hath bought thee? hath he not made thee, and established thee?
DEUT|32|7|Remember the days of old, consider the years of many generations: ask thy father, and he will show thee; thy elders, and they will tell thee.
DEUT|32|8|When the Most High divided to the nations their inheritance, when he separated the sons of Adam, he set the bounds of the people according to the number of the children of Israel.
DEUT|32|9|For the LORD's portion is his people; Jacob is the lot of his inheritance.
DEUT|32|10|He found him in a desert land, and in the waste howling wilderness; he led him about, he instructed him, he kept him as the apple of his eye.
DEUT|32|11|As an eagle stirreth up her nest, fluttereth over her young, spreadeth abroad her wings, taketh them, beareth them on her wings:
DEUT|32|12|So the LORD alone did lead him, and there was no strange god with him.
DEUT|32|13|He made him ride on the high places of the earth, that he might eat the increase of the fields; and he made him to suck honey out of the rock, and oil out of the flinty rock;
DEUT|32|14|Butter of kine, and milk of sheep, with fat of lambs, and rams of the breed of Bashan, and goats, with the fat of kidneys of wheat; and thou didst drink the pure blood of the grape.
DEUT|32|15|But Jeshurun waxed fat, and kicked: thou art waxen fat, thou art grown thick, thou art covered with fatness; then he forsook God which made him, and lightly esteemed the Rock of his salvation.
DEUT|32|16|They provoked him to jealousy with strange gods, with abominations provoked they him to anger.
DEUT|32|17|They sacrificed unto devils, not to God; to gods whom they knew not, to new gods that came newly up, whom your fathers feared not.
DEUT|32|18|Of the Rock that begat thee thou art unmindful, and hast forgotten God that formed thee.
DEUT|32|19|And when the LORD saw it, he abhorred them, because of the provoking of his sons, and of his daughters.
DEUT|32|20|And he said, I will hide my face from them, I will see what their end shall be: for they are a very froward generation, children in whom is no faith.
DEUT|32|21|They have moved me to jealousy with that which is not God; they have provoked me to anger with their vanities: and I will move them to jealousy with those which are not a people; I will provoke them to anger with a foolish nation.
DEUT|32|22|For a fire is kindled in mine anger, and shall burn unto the lowest hell, and shall consume the earth with her increase, and set on fire the foundations of the mountains.
DEUT|32|23|I will heap mischiefs upon them; I will spend mine arrows upon them.
DEUT|32|24|They shall be burnt with hunger, and devoured with burning heat, and with bitter destruction: I will also send the teeth of beasts upon them, with the poison of serpents of the dust.
DEUT|32|25|The sword without, and terror within, shall destroy both the young man and the virgin, the suckling also with the man of gray hairs.
DEUT|32|26|I said, I would scatter them into corners, I would make the remembrance of them to cease from among men:
DEUT|32|27|Were it not that I feared the wrath of the enemy, lest their adversaries should behave themselves strangely, and lest they should say, Our hand is high, and the LORD hath not done all this.
DEUT|32|28|For they are a nation void of counsel, neither is there any understanding in them.
DEUT|32|29|O that they were wise, that they understood this, that they would consider their latter end!
DEUT|32|30|How should one chase a thousand, and two put ten thousand to flight, except their Rock had sold them, and the LORD had shut them up?
DEUT|32|31|For their rock is not as our Rock, even our enemies themselves being judges.
DEUT|32|32|For their vine is of the vine of Sodom, and of the fields of Gomorrah: their grapes are grapes of gall, their clusters are bitter:
DEUT|32|33|Their wine is the poison of dragons, and the cruel venom of asps.
DEUT|32|34|Is not this laid up in store with me, and sealed up among my treasures?
DEUT|32|35|To me belongeth vengeance and recompence; their foot shall slide in due time: for the day of their calamity is at hand, and the things that shall come upon them make haste.
DEUT|32|36|For the LORD shall judge his people, and repent himself for his servants, when he seeth that their power is gone, and there is none shut up, or left.
DEUT|32|37|And he shall say, Where are their gods, their rock in whom they trusted,
DEUT|32|38|Which did eat the fat of their sacrifices, and drank the wine of their drink offerings? let them rise up and help you, and be your protection.
DEUT|32|39|See now that I, even I, am he, and there is no god with me: I kill, and I make alive; I wound, and I heal: neither is there any that can deliver out of my hand.
DEUT|32|40|For I lift up my hand to heaven, and say, I live for ever.
DEUT|32|41|If I whet my glittering sword, and mine hand take hold on judgment; I will render vengeance to mine enemies, and will reward them that hate me.
DEUT|32|42|I will make mine arrows drunk with blood, and my sword shall devour flesh; and that with the blood of the slain and of the captives, from the beginning of revenges upon the enemy.
DEUT|32|43|Rejoice, O ye nations, with his people: for he will avenge the blood of his servants, and will render vengeance to his adversaries, and will be merciful unto his land, and to his people.
DEUT|32|44|And Moses came and spake all the words of this song in the ears of the people, he, and Hoshea the son of Nun.
DEUT|32|45|And Moses made an end of speaking all these words to all Israel:
DEUT|32|46|And he said unto them, Set your hearts unto all the words which I testify among you this day, which ye shall command your children to observe to do, all the words of this law.
DEUT|32|47|For it is not a vain thing for you; because it is your life: and through this thing ye shall prolong your days in the land, whither ye go over Jordan to possess it.
DEUT|32|48|And the LORD spake unto Moses that selfsame day, saying,
DEUT|32|49|Get thee up into this mountain Abarim, unto mount Nebo, which is in the land of Moab, that is over against Jericho; and behold the land of Canaan, which I give unto the children of Israel for a possession:
DEUT|32|50|And die in the mount whither thou goest up, and be gathered unto thy people; as Aaron thy brother died in mount Hor, and was gathered unto his people:
DEUT|32|51|Because ye trespassed against me among the children of Israel at the waters of MeribahKadesh, in the wilderness of Zin; because ye sanctified me not in the midst of the children of Israel.
DEUT|32|52|Yet thou shalt see the land before thee; but thou shalt not go thither unto the land which I give the children of Israel.
DEUT|33|1|And this is the blessing, wherewith Moses the man of God blessed the children of Israel before his death.
DEUT|33|2|And he said, The LORD came from Sinai, and rose up from Seir unto them; he shined forth from mount Paran, and he came with ten thousands of saints: from his right hand went a fiery law for them.
DEUT|33|3|Yea, he loved the people; all his saints are in thy hand: and they sat down at thy feet; every one shall receive of thy words.
DEUT|33|4|Moses commanded us a law, even the inheritance of the congregation of Jacob.
DEUT|33|5|And he was king in Jeshurun, when the heads of the people and the tribes of Israel were gathered together.
DEUT|33|6|Let Reuben live, and not die; and let not his men be few.
DEUT|33|7|And this is the blessing of Judah: and he said, Hear, LORD, the voice of Judah, and bring him unto his people: let his hands be sufficient for him; and be thou an help to him from his enemies.
DEUT|33|8|And of Levi he said, Let thy Thummim and thy Urim be with thy holy one, whom thou didst prove at Massah, and with whom thou didst strive at the waters of Meribah;
DEUT|33|9|Who said unto his father and to his mother, I have not seen him; neither did he acknowledge his brethren, nor knew his own children: for they have observed thy word, and kept thy covenant.
DEUT|33|10|They shall teach Jacob thy judgments, and Israel thy law: they shall put incense before thee, and whole burnt sacrifice upon thine altar.
DEUT|33|11|Bless, LORD, his substance, and accept the work of his hands; smite through the loins of them that rise against him, and of them that hate him, that they rise not again.
DEUT|33|12|And of Benjamin he said, The beloved of the LORD shall dwell in safety by him; and the Lord shall cover him all the day long, and he shall dwell between his shoulders.
DEUT|33|13|And of Joseph he said, Blessed of the LORD be his land, for the precious things of heaven, for the dew, and for the deep that coucheth beneath,
DEUT|33|14|And for the precious fruits brought forth by the sun, and for the precious things put forth by the moon,
DEUT|33|15|And for the chief things of the ancient mountains, and for the precious things of the lasting hills,
DEUT|33|16|And for the precious things of the earth and fulness thereof, and for the good will of him that dwelt in the bush: let the blessing come upon the head of Joseph, and upon the top of the head of him that was separated from his brethren.
DEUT|33|17|His glory is like the firstling of his bullock, and his horns are like the horns of unicorns: with them he shall push the people together to the ends of the earth: and they are the ten thousands of Ephraim, and they are the thousands of Manasseh.
DEUT|33|18|And of Zebulun he said, Rejoice, Zebulun, in thy going out; and, Issachar, in thy tents.
DEUT|33|19|They shall call the people unto the mountain; there they shall offer sacrifices of righteousness: for they shall suck of the abundance of the seas, and of treasures hid in the sand.
DEUT|33|20|And of Gad he said, Blessed be he that enlargeth Gad: he dwelleth as a lion, and teareth the arm with the crown of the head.
DEUT|33|21|And he provided the first part for himself, because there, in a portion of the lawgiver, was he seated; and he came with the heads of the people, he executed the justice of the LORD, and his judgments with Israel.
DEUT|33|22|And of Dan he said, Dan is a lion's whelp: he shall leap from Bashan.
DEUT|33|23|And of Naphtali he said, O Naphtali, satisfied with favor, and full with the blessing of the LORD: possess thou the west and the south.
DEUT|33|24|And of Asher he said, Let Asher be blessed with children; let him be acceptable to his brethren, and let him dip his foot in oil.
DEUT|33|25|Thy shoes shall be iron and brass; and as thy days, so shall thy strength be.
DEUT|33|26|There is none like unto the God of Jeshurun, who rideth upon the heaven in thy help, and in his excellency on the sky.
DEUT|33|27|The eternal God is thy refuge, and underneath are the everlasting arms: and he shall thrust out the enemy from before thee; and shall say, Destroy them.
DEUT|33|28|Israel then shall dwell in safety alone: the fountain of Jacob shall be upon a land of corn and wine; also his heavens shall drop down dew.
DEUT|33|29|Happy art thou, O Israel: who is like unto thee, O people saved by the LORD, the shield of thy help, and who is the sword of thy excellency! and thine enemies shall be found liars unto thee; and thou shalt tread upon their high places.
DEUT|34|1|And Moses went up from the plains of Moab unto the mountain of Nebo, to the top of Pisgah, that is over against Jericho. And the LORD showed him all the land of Gilead, unto Dan,
DEUT|34|2|And all Naphtali, and the land of Ephraim, and Manasseh, and all the land of Judah, unto the utmost sea,
DEUT|34|3|And the south, and the plain of the valley of Jericho, the city of palm trees, unto Zoar.
DEUT|34|4|And the LORD said unto him, This is the land which I sware unto Abraham, unto Isaac, and unto Jacob, saying, I will give it unto thy seed: I have caused thee to see it with thine eyes, but thou shalt not go over thither.
DEUT|34|5|So Moses the servant of the LORD died there in the land of Moab, according to the word of the LORD.
DEUT|34|6|And he buried him in a valley in the land of Moab, over against Bethpeor: but no man knoweth of his sepulchre unto this day.
DEUT|34|7|And Moses was an hundred and twenty years old when he died: his eye was not dim, nor his natural force abated.
DEUT|34|8|And the children of Israel wept for Moses in the plains of Moab thirty days: so the days of weeping and mourning for Moses were ended.
DEUT|34|9|And Joshua the son of Nun was full of the spirit of wisdom; for Moses had laid his hands upon him: and the children of Israel hearkened unto him, and did as the LORD commanded Moses.
DEUT|34|10|And there arose not a prophet since in Israel like unto Moses, whom the LORD knew face to face,
DEUT|34|11|In all the signs and the wonders, which the LORD sent him to do in the land of Egypt to Pharaoh, and to all his servants, and to all his land,
DEUT|34|12|And in all that mighty hand, and in all the great terror which Moses showed in the sight of all Israel.
