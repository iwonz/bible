1PET|1|1|Peter, an apostle of Jesus Christ, To God's elect, strangers in the world, scattered throughout Pontus, Galatia, Cappadocia, Asia and Bithynia,
1PET|1|2|who have been chosen according to the foreknowledge of God the Father, through the sanctifying work of the Spirit, for obedience to Jesus Christ and sprinkling by his blood: Grace and peace be yours in abundance.
1PET|1|3|Praise be to the God and Father of our Lord Jesus Christ! In his great mercy he has given us new birth into a living hope through the resurrection of Jesus Christ from the dead,
1PET|1|4|and into an inheritance that can never perish, spoil or fade--kept in heaven for you,
1PET|1|5|who through faith are shielded by God's power until the coming of the salvation that is ready to be revealed in the last time.
1PET|1|6|In this you greatly rejoice, though now for a little while you may have had to suffer grief in all kinds of trials.
1PET|1|7|These have come so that your faith--of greater worth than gold, which perishes even though refined by fire--may be proved genuine and may result in praise, glory and honor when Jesus Christ is revealed.
1PET|1|8|Though you have not seen him, you love him; and even though you do not see him now, you believe in him and are filled with an inexpressible and glorious joy,
1PET|1|9|for you are receiving the goal of your faith, the salvation of your souls.
1PET|1|10|Concerning this salvation, the prophets, who spoke of the grace that was to come to you, searched intently and with the greatest care,
1PET|1|11|trying to find out the time and circumstances to which the Spirit of Christ in them was pointing when he predicted the sufferings of Christ and the glories that would follow.
1PET|1|12|It was revealed to them that they were not serving themselves but you, when they spoke of the things that have now been told you by those who have preached the gospel to you by the Holy Spirit sent from heaven. Even angels long to look into these things.
1PET|1|13|Therefore, prepare your minds for action; be self-controlled; set your hope fully on the grace to be given you when Jesus Christ is revealed.
1PET|1|14|As obedient children, do not conform to the evil desires you had when you lived in ignorance.
1PET|1|15|But just as he who called you is holy, so be holy in all you do;
1PET|1|16|for it is written: "Be holy, because I am holy."
1PET|1|17|Since you call on a Father who judges each man's work impartially, live your lives as strangers here in reverent fear.
1PET|1|18|For you know that it was not with perishable things such as silver or gold that you were redeemed from the empty way of life handed down to you from your forefathers,
1PET|1|19|but with the precious blood of Christ, a lamb without blemish or defect.
1PET|1|20|He was chosen before the creation of the world, but was revealed in these last times for your sake.
1PET|1|21|Through him you believe in God, who raised him from the dead and glorified him, and so your faith and hope are in God.
1PET|1|22|Now that you have purified yourselves by obeying the truth so that you have sincere love for your brothers, love one another deeply, from the heart.
1PET|1|23|For you have been born again, not of perishable seed, but of imperishable, through the living and enduring word of God.
1PET|1|24|For, "All men are like grass, and all their glory is like the flowers of the field; the grass withers and the flowers fall,
1PET|1|25|but the word of the Lord stands forever." And this is the word that was preached to you.
1PET|2|1|Therefore, rid yourselves of all malice and all deceit, hypocrisy, envy, and slander of every kind.
1PET|2|2|Like newborn babies, crave pure spiritual milk, so that by it you may grow up in your salvation,
1PET|2|3|now that you have tasted that the Lord is good.
1PET|2|4|As you come to him, the living Stone--rejected by men but chosen by God and precious to him--
1PET|2|5|you also, like living stones, are being built into a spiritual house to be a holy priesthood, offering spiritual sacrifices acceptable to God through Jesus Christ.
1PET|2|6|For in Scripture it says: "See, I lay a stone in Zion, a chosen and precious cornerstone, and the one who trusts in him will never be put to shame."
1PET|2|7|Now to you who believe, this stone is precious. But to those who do not believe, "The stone the builders rejected has become the capstone, "
1PET|2|8|and, "A stone that causes men to stumble and a rock that makes them fall." They stumble because they disobey the message--which is also what they were destined for.
1PET|2|9|But you are a chosen people, a royal priesthood, a holy nation, a people belonging to God, that you may declare the praises of him who called you out of darkness into his wonderful light.
1PET|2|10|Once you were not a people, but now you are the people of God; once you had not received mercy, but now you have received mercy.
1PET|2|11|Dear friends, I urge you, as aliens and strangers in the world, to abstain from sinful desires, which war against your soul.
1PET|2|12|Live such good lives among the pagans that, though they accuse you of doing wrong, they may see your good deeds and glorify God on the day he visits us.
1PET|2|13|Submit yourselves for the Lord's sake to every authority instituted among men: whether to the king, as the supreme authority,
1PET|2|14|or to governors, who are sent by him to punish those who do wrong and to commend those who do right.
1PET|2|15|For it is God's will that by doing good you should silence the ignorant talk of foolish men.
1PET|2|16|Live as free men, but do not use your freedom as a cover-up for evil; live as servants of God.
1PET|2|17|Show proper respect to everyone: Love the brotherhood of believers, fear God, honor the king.
1PET|2|18|Slaves, submit yourselves to your masters with all respect, not only to those who are good and considerate, but also to those who are harsh.
1PET|2|19|For it is commendable if a man bears up under the pain of unjust suffering because he is conscious of God.
1PET|2|20|But how is it to your credit if you receive a beating for doing wrong and endure it? But if you suffer for doing good and you endure it, this is commendable before God.
1PET|2|21|To this you were called, because Christ suffered for you, leaving you an example, that you should follow in his steps.
1PET|2|22|"He committed no sin, and no deceit was found in his mouth."
1PET|2|23|When they hurled their insults at him, he did not retaliate; when he suffered, he made no threats. Instead, he entrusted himself to him who judges justly.
1PET|2|24|He himself bore our sins in his body on the tree, so that we might die to sins and live for righteousness; by his wounds you have been healed.
1PET|2|25|For you were like sheep going astray, but now you have returned to the Shepherd and Overseer of your souls.
1PET|3|1|Wives, in the same way be submissive to your husbands so that, if any of them do not believe the word, they may be won over without words by the behavior of their wives,
1PET|3|2|when they see the purity and reverence of your lives.
1PET|3|3|Your beauty should not come from outward adornment, such as braided hair and the wearing of gold jewelry and fine clothes.
1PET|3|4|Instead, it should be that of your inner self, the unfading beauty of a gentle and quiet spirit, which is of great worth in God's sight.
1PET|3|5|For this is the way the holy women of the past who put their hope in God used to make themselves beautiful. They were submissive to their own husbands,
1PET|3|6|like Sarah, who obeyed Abraham and called him her master. You are her daughters if you do what is right and do not give way to fear.
1PET|3|7|Husbands, in the same way be considerate as you live with your wives, and treat them with respect as the weaker partner and as heirs with you of the gracious gift of life, so that nothing will hinder your prayers.
1PET|3|8|Finally, all of you, live in harmony with one another; be sympathetic, love as brothers, be compassionate and humble.
1PET|3|9|Do not repay evil with evil or insult with insult, but with blessing, because to this you were called so that you may inherit a blessing.
1PET|3|10|For, "Whoever would love life and see good days must keep his tongue from evil and his lips from deceitful speech.
1PET|3|11|He must turn from evil and do good; he must seek peace and pursue it.
1PET|3|12|For the eyes of the Lord are on the righteous and his ears are attentive to their prayer, but the face of the Lord is against those who do evil."
1PET|3|13|Who is going to harm you if you are eager to do good?
1PET|3|14|But even if you should suffer for what is right, you are blessed. "Do not fear what they fear; do not be frightened."
1PET|3|15|But in your hearts set apart Christ as Lord. Always be prepared to give an answer to everyone who asks you to give the reason for the hope that you have. But do this with gentleness and respect,
1PET|3|16|keeping a clear conscience, so that those who speak maliciously against your good behavior in Christ may be ashamed of their slander.
1PET|3|17|It is better, if it is God's will, to suffer for doing good than for doing evil.
1PET|3|18|For Christ died for sins once for all, the righteous for the unrighteous, to bring you to God. He was put to death in the body but made alive by the Spirit,
1PET|3|19|through whom also he went and preached to the spirits in prison
1PET|3|20|who disobeyed long ago when God waited patiently in the days of Noah while the ark was being built. In it only a few people, eight in all, were saved through water,
1PET|3|21|and this water symbolizes baptism that now saves you also--not the removal of dirt from the body but the pledge of a good conscience toward God. It saves you by the resurrection of Jesus Christ,
1PET|3|22|who has gone into heaven and is at God's right hand--with angels, authorities and powers in submission to him.
1PET|4|1|Therefore, since Christ suffered in his body, arm yourselves also with the same attitude, because he who has suffered in his body is done with sin.
1PET|4|2|As a result, he does not live the rest of his earthly life for evil human desires, but rather for the will of God.
1PET|4|3|For you have spent enough time in the past doing what pagans choose to do--living in debauchery, lust, drunkenness, orgies, carousing and detestable idolatry.
1PET|4|4|They think it strange that you do not plunge with them into the same flood of dissipation, and they heap abuse on you.
1PET|4|5|But they will have to give account to him who is ready to judge the living and the dead.
1PET|4|6|For this is the reason the gospel was preached even to those who are now dead, so that they might be judged according to men in regard to the body, but live according to God in regard to the spirit.
1PET|4|7|The end of all things is near. Therefore be clear minded and self-controlled so that you can pray.
1PET|4|8|Above all, love each other deeply, because love covers over a multitude of sins.
1PET|4|9|Offer hospitality to one another without grumbling.
1PET|4|10|Each one should use whatever gift he has received to serve others, faithfully administering God's grace in its various forms.
1PET|4|11|If anyone speaks, he should do it as one speaking the very words of God. If anyone serves, he should do it with the strength God provides, so that in all things God may be praised through Jesus Christ. To him be the glory and the power for ever and ever. Amen.
1PET|4|12|Dear friends, do not be surprised at the painful trial you are suffering, as though something strange were happening to you.
1PET|4|13|But rejoice that you participate in the sufferings of Christ, so that you may be overjoyed when his glory is revealed.
1PET|4|14|If you are insulted because of the name of Christ, you are blessed, for the Spirit of glory and of God rests on you.
1PET|4|15|If you suffer, it should not be as a murderer or thief or any other kind of criminal, or even as a meddler.
1PET|4|16|However, if you suffer as a Christian, do not be ashamed, but praise God that you bear that name.
1PET|4|17|For it is time for judgment to begin with the family of God; and if it begins with us, what will the outcome be for those who do not obey the gospel of God?
1PET|4|18|And, "If it is hard for the righteous to be saved, what will become of the ungodly and the sinner?"
1PET|4|19|So then, those who suffer according to God's will should commit themselves to their faithful Creator and continue to do good.
1PET|5|1|To the elders among you, I appeal as a fellow elder, a witness of Christ's sufferings and one who also will share in the glory to be revealed:
1PET|5|2|Be shepherds of God's flock that is under your care, serving as overseers--not because you must, but because you are willing, as God wants you to be; not greedy for money, but eager to serve;
1PET|5|3|not lording it over those entrusted to you, but being examples to the flock.
1PET|5|4|And when the Chief Shepherd appears, you will receive the crown of glory that will never fade away.
1PET|5|5|Young men, in the same way be submissive to those who are older. All of you, clothe yourselves with humility toward one another, because, "God opposes the proud but gives grace to the humble."
1PET|5|6|Humble yourselves, therefore, under God's mighty hand, that he may lift you up in due time.
1PET|5|7|Cast all your anxiety on him because he cares for you.
1PET|5|8|Be self-controlled and alert. Your enemy the devil prowls around like a roaring lion looking for someone to devour.
1PET|5|9|Resist him, standing firm in the faith, because you know that your brothers throughout the world are undergoing the same kind of sufferings.
1PET|5|10|And the God of all grace, who called you to his eternal glory in Christ, after you have suffered a little while, will himself restore you and make you strong, firm and steadfast.
1PET|5|11|To him be the power for ever and ever. Amen.
1PET|5|12|With the help of Silas, whom I regard as a faithful brother, I have written to you briefly, encouraging you and testifying that this is the true grace of God. Stand fast in it.
1PET|5|13|She who is in Babylon, chosen together with you, sends you her greetings, and so does my son Mark.
1PET|5|14|Greet one another with a kiss of love. Peace to all of you who are in Christ.
