DEUT|1|1|haec sunt verba quae locutus est Moses ad omnem Israhel trans Iordanem in solitudine campestri contra mare Rubrum inter Pharan et Thophel et Laban et Aseroth ubi auri est plurimum
DEUT|1|2|undecim diebus de Horeb per viam montis Seir usque Cadesbarne
DEUT|1|3|quadragesimo anno undecimo mense prima die mensis locutus est Moses ad filios Israhel omnia quae praeceperat illi Dominus ut diceret eis
DEUT|1|4|postquam percussit Seon regem Amorreorum qui habitavit in Esebon et Og regem Basan qui mansit in Aseroth et in Edrai
DEUT|1|5|trans Iordanem in terra Moab coepitque Moses explanare legem et dicere
DEUT|1|6|Dominus Deus noster locutus est ad nos in Horeb dicens sufficit vobis quod in hoc monte mansistis
DEUT|1|7|revertimini et venite ad montem Amorreorum et ad cetera quae ei proxima sunt campestria atque montana et humiliora loca contra meridiem et iuxta litus maris terram Chananeorum et Libani usque ad flumen magnum Eufraten
DEUT|1|8|en inquit tradidi vobis ingredimini et possidete eam super qua iuravit Dominus patribus vestris Abraham et Isaac et Iacob ut daret illam eis et semini eorum post eos
DEUT|1|9|dixique vobis illo in tempore
DEUT|1|10|non possum solus sustinere vos quia Dominus Deus vester multiplicavit vos et estis hodie sicut stellae caeli plurimae
DEUT|1|11|Dominus Deus patrum vestrorum addat ad hunc numerum multa milia et benedicat vobis sicut locutus est
DEUT|1|12|non valeo solus vestra negotia sustinere et pondus ac iurgia
DEUT|1|13|date e vobis viros sapientes et gnaros et quorum conversatio sit probata in tribubus vestris ut ponam eos vobis principes
DEUT|1|14|tunc respondistis mihi bona res est quam vis facere
DEUT|1|15|tulique de tribubus vestris viros sapientes et nobiles et constitui eos principes tribunos et centuriones et quinquagenarios ac decanos qui docerent vos singula
DEUT|1|16|praecepique eis dicens audite illos et quod iustum est iudicate sive civis sit ille sive peregrinus
DEUT|1|17|nulla erit distantia personarum ita parvum audietis ut magnum nec accipietis cuiusquam personam quia Dei iudicium est quod si difficile vobis aliquid visum fuerit referte ad me et ego audiam
DEUT|1|18|praecepique omnia quae facere deberetis
DEUT|1|19|profecti autem de Horeb transivimus per heremum terribilem et maximam quam vidistis per viam montis Amorrei sicut praeceperat Dominus Deus noster nobis cumque venissemus in Cadesbarne
DEUT|1|20|dixi vobis venistis ad montem Amorrei quem Dominus Deus noster daturus est nobis
DEUT|1|21|vide terram quam Dominus Deus tuus dat tibi ascende et posside eam sicut locutus est Dominus Deus patribus tuis noli metuere nec quicquam paveas
DEUT|1|22|et accessistis ad me omnes atque dixistis mittamus viros qui considerent terram et renuntient per quod iter debeamus ascendere et ad quas pergere civitates
DEUT|1|23|cumque mihi sermo placuisset misi e vobis duodecim viros singulos de tribubus suis
DEUT|1|24|qui cum perrexissent et ascendissent in montana venerunt usque ad vallem Botri et considerata terra
DEUT|1|25|sumentes de fructibus eius ut ostenderent ubertatem adtulerunt ad nos atque dixerunt bona est terra quam Dominus Deus noster daturus est nobis
DEUT|1|26|et noluistis ascendere sed increduli ad sermonem Domini Dei nostri
DEUT|1|27|murmurati estis in tabernaculis vestris atque dixistis odit nos Dominus et idcirco eduxit nos de terra Aegypti ut traderet in manu Amorrei atque deleret
DEUT|1|28|quo ascendemus nuntii terruerunt cor nostrum dicentes maxima multitudo est et nobis in statura procerior urbes magnae et ad caelum usque munitae filios Enacim vidimus ibi
DEUT|1|29|et dixi vobis nolite metuere nec timeatis eos
DEUT|1|30|Dominus Deus qui ductor est vester pro vobis ipse pugnabit sicut fecit in Aegypto videntibus cunctis
DEUT|1|31|et in solitudine ipse vidisti portavit te Dominus Deus tuus ut solet homo gestare parvulum filium suum in omni via per quam ambulasti donec veniretis ad locum istum
DEUT|1|32|et nec sic quidem credidistis Domino Deo vestro
DEUT|1|33|qui praecessit vos in via et metatus est locum in quo tentoria figere deberetis nocte ostendens vobis iter per ignem et die per columnam nubis
DEUT|1|34|cumque audisset Dominus vocem sermonum vestrorum iratus iuravit et ait
DEUT|1|35|non videbit quispiam de hominibus generationis huius pessimae terram bonam quam sub iuramento pollicitus sum patribus vestris
DEUT|1|36|praeter Chaleb filium Iepphonne ipse enim videbit eam et ipsi dabo terram quam calcavit et filiis eius quia secutus est Dominum
DEUT|1|37|nec miranda indignatio in populum cum mihi quoque iratus Dominus propter vos dixerit nec tu ingredieris illuc
DEUT|1|38|sed Iosue filius Nun minister tuus ipse intrabit pro te hunc exhortare et robora et ipse terram sorte dividat Israheli
DEUT|1|39|parvuli vestri de quibus dixistis quod captivi ducerentur et filii qui hodie boni ac mali ignorant distantiam ipsi ingredientur et ipsis dabo terram et possidebunt eam
DEUT|1|40|vos autem revertimini et abite in solitudinem per viam maris Rubri
DEUT|1|41|et respondistis mihi peccavimus Domino ascendemus atque pugnabimus sicut praecepit Dominus Deus noster cumque instructi armis pergeretis in montem
DEUT|1|42|ait mihi Dominus dic ad eos nolite ascendere neque pugnetis non enim sum vobiscum ne cadatis coram inimicis vestris
DEUT|1|43|locutus sum et non audistis sed adversantes imperio Domini et tumentes superbia ascendistis in montem
DEUT|1|44|itaque egressus Amorreus qui habitabat in montibus et obviam veniens persecutus est vos sicut solent apes persequi et cecidit de Seir usque Horma
DEUT|1|45|cumque reversi ploraretis coram Domino non audivit vos nec voci vestrae voluit adquiescere
DEUT|1|46|sedistis ergo in Cadesbarne multo tempore
DEUT|2|1|profectique inde venimus in solitudinem quae ducit ad mare Rubrum sicut mihi dixerat Dominus et circumivimus montem Seir longo tempore
DEUT|2|2|dixitque Dominus ad me
DEUT|2|3|sufficit vobis circumire montem istum ite contra aquilonem
DEUT|2|4|et populo praecipe dicens transibitis per terminos fratrum vestrorum filiorum Esau qui habitant in Seir et timebunt vos
DEUT|2|5|videte ergo diligenter ne moveamini contra eos neque enim dabo vobis de terra eorum quantum potest unius pedis calcare vestigium quia in possessionem Esau dedi montem Seir
DEUT|2|6|cibos emetis ab eis pecunia et comedetis aquam emptam haurietis et bibetis
DEUT|2|7|Dominus Deus tuus benedixit tibi in omni opere manuum tuarum novit iter tuum quomodo transieris solitudinem hanc magnam per quadraginta annos habitans tecum Dominus Deus tuus et nihil tibi defuit
DEUT|2|8|cumque transissemus fratres nostros filios Esau qui habitabant in Seir per viam campestrem de Helath et de Asiongaber venimus ad iter quod ducit in desertum Moab
DEUT|2|9|dixitque Dominus ad me non pugnes contra Moabitas nec ineas adversum eos proelium non enim dabo tibi quicquam de terra eorum quia filiis Loth tradidi Ar in possessionem
DEUT|2|10|Emim primi fuerunt habitatores eius populus magnus et validus et tam excelsus ut de Enacim stirpe
DEUT|2|11|quasi gigantes crederentur et essent similes filiorum Enacim denique Moabitae appellant eos Emim
DEUT|2|12|in Seir autem prius habitaverunt Horim quibus expulsis atque deletis habitaverunt filii Esau sicut fecit Israhel in terra possessionis suae quam dedit ei Dominus
DEUT|2|13|surgentes ergo ut transiremus torrentem Zared venimus ad eum
DEUT|2|14|tempus autem quo ambulavimus de Cadesbarne usque ad transitum torrentis Zared triginta octo annorum fuit donec consumeretur omnis generatio hominum bellatorum de castris sicut iuraverat Dominus
DEUT|2|15|cuius manus fuit adversum eos ut interirent de castrorum medio
DEUT|2|16|postquam autem universi ceciderunt pugnatores
DEUT|2|17|locutus est Dominus ad me dicens
DEUT|2|18|tu transibis hodie terminos Moab urbem nomine Ar
DEUT|2|19|et accedens in vicina filiorum Ammon cave ne pugnes contra eos nec movearis ad proelium non enim dabo tibi de terra filiorum Ammon quia filiis Loth dedi eam in possessionem
DEUT|2|20|terra gigantum reputata est et in ipsa olim habitaverunt gigantes quos Ammanitae vocant Zomzommim
DEUT|2|21|populus magnus et multus et procerae longitudinis sicut Enacim quos delevit Dominus a facie eorum et fecit illos habitare pro eis
DEUT|2|22|sicut fecerat filiis Esau qui habitant in Seir delens Horreos et terram eorum illis tradens quam possident usque in praesens
DEUT|2|23|Eveos quoque qui habitabant in Aserim usque Gazam Cappadoces expulerunt qui egressi de Cappadocia deleverunt eos et habitaverunt pro illis
DEUT|2|24|surgite et transite torrentem Arnon ecce tradidi in manu tua Seon regem Esebon Amorreum et terram eius incipe possidere et committe adversum eum proelium
DEUT|2|25|hodie incipiam mittere terrorem atque formidinem tuam in populos qui habitant sub omni caelo ut audito nomine tuo paveant et in morem parturientium contremescant et dolore teneantur
DEUT|2|26|misi ergo nuntios de solitudine Cademoth ad Seon regem Esebon verbis pacificis dicens
DEUT|2|27|transibimus per terram tuam publica gradiemur via non declinabimus neque ad dextram neque ad sinistram
DEUT|2|28|alimenta pretio vende nobis ut vescamur aquam pecunia tribue et sic bibemus tantum est ut nobis concedas transitum
DEUT|2|29|sicut fecerunt filii Esau qui habitant in Seir et Moabitae qui morantur in Ar donec veniamus ad Iordanem et transeamus in terram quam Dominus Deus noster daturus est nobis
DEUT|2|30|noluitque Seon rex Esebon dare nobis transitum quia induraverat Dominus Deus tuus spiritum eius et obfirmaverat cor illius ut traderetur in manus tuas sicut nunc vides
DEUT|2|31|dixitque Dominus ad me ecce coepi tradere tibi Seon et terram eius incipe possidere eam
DEUT|2|32|egressusque est Seon obviam nobis cum omni populo suo ad proelium in Iesa
DEUT|2|33|et tradidit eum Dominus Deus noster nobis percussimusque eum cum filiis et omni populo suo
DEUT|2|34|cunctasque urbes in tempore illo cepimus interfectis habitatoribus earum viris ac mulieribus et parvulis non reliquimus in eis quicquam
DEUT|2|35|absque iumentis quae in partem venere praedantium et spoliis urbium quas cepimus
DEUT|2|36|ab Aroer quae est super ripam torrentis Arnon oppido quod in valle situm est usque Galaad non fuit vicus et civitas quae nostras effugeret manus omnes tradidit Dominus Deus noster nobis
DEUT|2|37|absque terra filiorum Ammon ad quam non accessimus et cunctis quae adiacent torrenti Ieboc et urbibus montanis universisque locis a quibus nos prohibuit Dominus Deus noster
DEUT|3|1|itaque conversi ascendimus per iter Basan egressusque est Og rex Basan in occursum nobis cum populo suo ad bellandum in Edrai
DEUT|3|2|dixitque Dominus ad me ne timeas eum quia in manu tua traditus est cum omni populo ac terra sua faciesque ei sicut fecisti Seon regi Amorreorum qui habitavit in Esebon
DEUT|3|3|tradidit ergo Dominus Deus noster in manibus nostris etiam Og regem Basan et universum populum eius percussimusque eos usque ad internicionem
DEUT|3|4|vastantes cunctas civitates illius uno tempore non fuit oppidum quod nos effugeret sexaginta urbes omnem regionem Argob regni Og in Basan
DEUT|3|5|cunctae urbes erant munitae muris altissimis portisque et vectibus absque oppidis innumeris quae non habebant muros
DEUT|3|6|et delevimus eos sicut feceramus Seon regi Esebon disperdentes omnem civitatem virosque ac mulieres et parvulos
DEUT|3|7|iumenta autem et spolia urbium diripuimus
DEUT|3|8|tulimusque illo in tempore terram de manu duorum regum Amorreorum qui erant trans Iordanem a torrente Arnon usque ad montem Hermon
DEUT|3|9|quem Sidonii Sarion vocant et Amorrei Sanir
DEUT|3|10|omnes civitates quae sitae sunt in planitie et universam terram Galaad et Basan usque Selcha et Edrai civitates regni Og in Basan
DEUT|3|11|solus quippe Og rex Basan restiterat de stirpe gigantum monstratur lectus eius ferreus qui est in Rabbath filiorum Ammon novem cubitos habens longitudinis et quattuor latitudinis ad mensuram cubiti virilis manus
DEUT|3|12|terramque possedimus in tempore illo ab Aroer quae est super ripam torrentis Arnon usque ad mediam partem montis Galaad et civitates illius dedi Ruben et Gad
DEUT|3|13|reliquam autem partem Galaad et omnem Basan regni Og tradidi mediae tribui Manasse omnem regionem Argob cuncta Basan vocatur terra gigantum
DEUT|3|14|Iair filius Manasse possedit omnem regionem Argob usque ad terminos Gesuri et Machathi vocavitque ex nomine suo Basan Avothiair id est villas Iair usque in praesentem diem
DEUT|3|15|Machir quoque dedi Galaad
DEUT|3|16|et tribubus Ruben et Gad dedi terram Galaad usque ad torrentem Arnon medium torrentis et finium usque ad torrentem Ieboc qui est terminus filiorum Ammon
DEUT|3|17|et planitiem solitudinis atque Iordanem et terminos Chenereth usque ad mare Deserti quod est Salsissimum ad radices montis Phasga contra orientem
DEUT|3|18|praecepique vobis in tempore illo dicens Dominus Deus vester dat vobis terram hanc in hereditatem expediti praecedite fratres vestros filios Israhel omnes viri robusti
DEUT|3|19|absque uxoribus et parvulis ac iumentis novi enim quod plura habeatis pecora et in urbibus remanere debebunt quas tradidi vobis
DEUT|3|20|donec requiem tribuat Dominus fratribus vestris sicut vobis tribuit et possideant etiam ipsi terram quam daturus est eis trans Iordanem tunc revertetur unusquisque in possessionem suam quam dedi vobis
DEUT|3|21|Iosue quoque in tempore illo praecepi dicens oculi tui viderunt quae fecit Dominus Deus vester duobus his regibus sic faciet omnibus regnis ad quae transiturus es
DEUT|3|22|ne timeas eos Dominus enim Deus vester pugnabit pro vobis
DEUT|3|23|precatusque sum Dominum in tempore illo dicens
DEUT|3|24|Domine Deus tu coepisti ostendere servo tuo magnitudinem tuam manumque fortissimam neque enim est alius Deus vel in caelo vel in terra qui possit facere opera tua et conparari fortitudini tuae
DEUT|3|25|transibo igitur et videbo terram hanc optimam trans Iordanem et montem istum egregium et Libanum
DEUT|3|26|iratusque est Dominus mihi propter vos nec exaudivit me sed dixit mihi sufficit tibi nequaquam ultra loquaris de hac re ad me
DEUT|3|27|ascende cacumen Phasgae et oculos tuos circumfer ad occidentem et aquilonem austrumque et orientem et aspice nec enim transibis Iordanem istum
DEUT|3|28|praecipe Iosue et corrobora eum atque conforta quia ipse praecedet populum istum et dividet eis terram quam visurus es
DEUT|3|29|mansimusque in valle contra fanum Phogor
DEUT|4|1|et nunc Israhel audi praecepta et iudicia quae ego doceo te ut faciens ea vivas et ingrediens possideas terram quam Dominus Deus patrum vestrorum daturus est vobis
DEUT|4|2|non addetis ad verbum quod vobis loquor neque auferetis ex eo custodite mandata Domini Dei vestri quae ego praecipio vobis
DEUT|4|3|oculi vestri viderunt omnia quae fecit Dominus contra Beelphegor quomodo contriverit omnes cultores eius de medio vestri
DEUT|4|4|vos autem qui adheretis Domino Deo vestro vivitis universi usque in praesentem diem
DEUT|4|5|scitis quod docuerim vos praecepta atque iustitias sicut mandavit mihi Dominus Deus meus sic facietis ea in terra quam possessuri estis
DEUT|4|6|et observabitis et implebitis opere haec est enim vestra sapientia et intellectus coram populis ut audientes universa praecepta haec dicant en populus sapiens et intellegens gens magna
DEUT|4|7|nec est alia natio tam grandis quae habeat deos adpropinquantes sibi sicut Dominus Deus noster adest cunctis obsecrationibus nostris
DEUT|4|8|quae est enim alia gens sic inclita ut habeat caerimonias iustaque iudicia et universam legem quam ego proponam hodie ante oculos vestros
DEUT|4|9|custodi igitur temet ipsum et animam tuam sollicite ne obliviscaris verborum quae viderunt oculi tui et ne excedant de corde tuo cunctis diebus vitae tuae docebis ea filios ac nepotes tuos
DEUT|4|10|diem in quo stetisti coram Domino Deo tuo in Horeb quando Dominus locutus est mihi dicens congrega ad me populum ut audiat sermones meos et discat timere me omni tempore quo vivit in terra doceantque filios suos
DEUT|4|11|et accessistis ad radices montis qui ardebat usque ad caelum erantque in eo tenebrae nubes et caligo
DEUT|4|12|locutusque est Dominus ad vos de medio ignis vocem verborum eius audistis et formam penitus non vidistis
DEUT|4|13|et ostendit vobis pactum suum quod praecepit ut faceretis et decem verba quae scripsit in duabus tabulis lapideis
DEUT|4|14|mihique mandavit in illo tempore ut docerem vos caerimonias et iudicia quae facere deberetis in terra quam possessuri estis
DEUT|4|15|custodite igitur sollicite animas vestras non vidistis aliquam similitudinem in die qua locutus est Dominus vobis in Horeb de medio ignis
DEUT|4|16|ne forte decepti faciatis vobis sculptam similitudinem aut imaginem masculi vel feminae
DEUT|4|17|similitudinem omnium iumentorum quae sunt super terram vel avium sub caelo volantium
DEUT|4|18|atque reptilium quae moventur in terra sive piscium qui sub terra morantur in aquis
DEUT|4|19|ne forte oculis elevatis ad caelum videas solem et lunam et omnia astra caeli et errore deceptus adores ea et colas quae creavit Dominus Deus tuus in ministerium cunctis gentibus quae sub caelo sunt
DEUT|4|20|vos autem tulit Dominus et eduxit de fornace ferrea Aegypti ut haberet populum hereditarium sicut est in praesenti die
DEUT|4|21|iratusque est Dominus contra me propter sermones vestros et iuravit ut non transirem Iordanem nec ingrederer terram optimam quam daturus est vobis
DEUT|4|22|ecce morior in hac humo non transibo Iordanem vos transibitis et possidebitis terram egregiam
DEUT|4|23|cave nequando obliviscaris pacti Domini Dei tui quod pepigit tecum et facias tibi sculptam similitudinem eorum quae fieri Dominus prohibuit
DEUT|4|24|quia Dominus Deus tuus ignis consumens est Deus aemulator
DEUT|4|25|si genueritis filios ac nepotes et morati fueritis in terra deceptique feceritis vobis aliquam similitudinem patrantes malum coram Domino Deo vestro ut eum ad iracundiam provocetis
DEUT|4|26|testes invoco hodie caelum et terram cito perituros vos esse de terra quam transito Iordane possessuri estis non habitabitis in ea longo tempore sed delebit vos Dominus
DEUT|4|27|atque disperget in omnes gentes et remanebitis pauci in nationibus ad quas vos ducturus est Dominus
DEUT|4|28|ibique servietis diis qui hominum manu fabricati sunt ligno et lapidi qui non vident non audiunt non comedunt non odorantur
DEUT|4|29|cumque quaesieris ibi Dominum Deum tuum invenies eum si tamen toto corde quaesieris et tota tribulatione animae tuae
DEUT|4|30|postquam te invenerint omnia quae praedicta sunt novissimo tempore reverteris ad Dominum Deum tuum et audies vocem eius
DEUT|4|31|quia Deus misericors Dominus Deus tuus est non dimittet te nec omnino delebit neque obliviscetur pacti in quo iuravit patribus tuis
DEUT|4|32|interroga de diebus antiquis qui fuerunt ante te ex die quo creavit Deus hominem super terram a summo caeli usque ad summum eius si facta est aliquando huiuscemodi res aut umquam cognitum est
DEUT|4|33|ut audiret populus vocem Dei loquentis de medio ignis sicut tu audisti et vixisti
DEUT|4|34|si fecit Deus ut ingrederetur et tolleret sibi gentem de medio nationum per temptationes signa atque portenta per pugnam et robustam manum extentumque brachium et horribiles visiones iuxta omnia quae fecit pro vobis Dominus Deus vester in Aegypto videntibus oculis tuis
DEUT|4|35|ut scires quoniam Dominus ipse est Deus et non est alius praeter unum
DEUT|4|36|de caelo te fecit audire vocem suam ut doceret te et in terra ostendit tibi ignem suum maximum et audisti verba illius de medio ignis
DEUT|4|37|quia dilexit patres tuos et elegit semen eorum post eos eduxitque te praecedens in virtute sua magna ex Aegypto
DEUT|4|38|ut deleret nationes maximas et fortiores te in introitu tuo et introduceret te daretque tibi terram earum in possessionem sicut cernis in praesenti die
DEUT|4|39|scito ergo hodie et cogitato in corde tuo quod Dominus ipse sit Deus in caelo sursum et in terra deorsum et non sit alius
DEUT|4|40|custodi praecepta eius atque mandata quae ego praecipio tibi ut bene sit tibi et filiis tuis post te et permaneas multo tempore super terram quam Dominus Deus tuus daturus est tibi
DEUT|4|41|tunc separavit Moses tres civitates trans Iordanem ad orientalem plagam
DEUT|4|42|ut confugiat ad eas qui occiderit nolens proximum suum nec fuerit inimicus ante unum et alterum diem et ad harum aliquam urbium possit evadere
DEUT|4|43|Bosor in solitudine quae sita est in terra campestri de tribu Ruben et Ramoth in Galaad quae est in tribu Gad et Golam in Basan quae est in tribu Manasse
DEUT|4|44|ista est lex quam proposuit Moses coram filiis Israhel
DEUT|4|45|et haec testimonia et caerimoniae atque iudicia quae locutus est ad filios Israhel quando egressi sunt de Aegypto
DEUT|4|46|trans Iordanem in valle contra fanum Phogor in terra Seon regis Amorrei qui habitavit in Esebon quem percussit Moses filii quoque Israhel egressi ex Aegypto
DEUT|4|47|possederunt terram eius et terram Og regis Basan duorum regum Amorreorum qui erant trans Iordanem ad solis ortum
DEUT|4|48|ab Aroer quae sita est super ripam torrentis Arnon usque ad montem Sion qui est et Hermon
DEUT|4|49|omnem planitiem trans Iordanem ad orientalem plagam usque ad mare Solitudinis et usque ad radices montis Phasga
DEUT|5|1|vocavitque Moses omnem Israhelem et dixit ad eum audi Israhel caerimonias atque iudicia quae ego loquor in auribus vestris hodie discite ea et opere conplete
DEUT|5|2|Dominus Deus noster pepigit nobiscum foedus in Horeb
DEUT|5|3|non cum patribus nostris iniit pactum sed nobiscum qui inpraesentiarum sumus et vivimus
DEUT|5|4|facie ad faciem locutus est nobis in monte de medio ignis
DEUT|5|5|ego sequester et medius fui inter Dominum et vos in tempore illo ut adnuntiarem vobis verba eius timuistis enim ignem et non ascendistis in montem et ait
DEUT|5|6|ego Dominus Deus tuus qui eduxi te de terra Aegypti de domo servitutis
DEUT|5|7|non habebis deos alienos in conspectu meo
DEUT|5|8|non facies tibi sculptile nec similitudinem omnium quae in caelo sunt desuper et quae in terra deorsum et quae versantur in aquis sub terra
DEUT|5|9|non adorabis ea et non coles ego enim sum Dominus Deus tuus Deus aemulator reddens iniquitatem patrum super filios in tertiam et quartam generationem his qui oderunt me
DEUT|5|10|et faciens misericordiam in multa milia diligentibus me et custodientibus praecepta mea
DEUT|5|11|non usurpabis nomen Domini Dei tui frustra quia non erit inpunitus qui super re vana nomen eius adsumpserit
DEUT|5|12|observa diem sabbati ut sanctifices eum sicut praecepit tibi Dominus Deus tuus
DEUT|5|13|sex diebus operaberis et facies omnia opera tua
DEUT|5|14|septimus dies sabbati est id est requies Domini Dei tui non facies in eo quicquam operis tu et filius tuus et filia servus et ancilla et bos et asinus et omne iumentum tuum et peregrinus qui est intra portas tuas ut requiescat servus et ancilla tua sicut et tu
DEUT|5|15|memento quod et ipse servieris in Aegypto et eduxerit te inde Dominus Deus tuus in manu forti et brachio extento idcirco praecepit tibi ut observares diem sabbati
DEUT|5|16|honora patrem tuum et matrem sicut praecepit tibi Dominus Deus tuus ut longo vivas tempore et bene sit tibi in terra quam Dominus Deus tuus daturus est tibi
DEUT|5|17|non occides
DEUT|5|18|neque moechaberis
DEUT|5|19|furtumque non facies
DEUT|5|20|nec loqueris contra proximum tuum falsum testimonium
DEUT|5|21|non concupisces uxorem proximi tui non domum non agrum non servum non ancillam non bovem non asinum et universa quae illius sunt
DEUT|5|22|haec verba locutus est Dominus ad omnem multitudinem vestram in monte de medio ignis et nubis et caliginis voce magna nihil addens amplius et scripsit ea in duabus tabulis lapideis quas tradidit mihi
DEUT|5|23|vos autem postquam audistis vocem de medio tenebrarum et montem ardere vidistis accessistis ad me omnes principes tribuum et maiores natu atque dixistis
DEUT|5|24|ecce ostendit nobis Dominus Deus noster maiestatem et magnitudinem suam vocem eius audivimus de medio ignis et probavimus hodie quod loquente Deo cum homine vixerit homo
DEUT|5|25|cur ergo morimur et devorabit nos ignis hic maximus si enim audierimus ultra vocem Domini Dei nostri moriemur
DEUT|5|26|quid est omnis caro ut audiat vocem Dei viventis qui de medio ignis loquitur sicut nos audivimus et possit vivere
DEUT|5|27|tu magis accede et audi cuncta quae dixerit Dominus Deus noster tibi loquerisque ad nos et nos audientes faciemus ea
DEUT|5|28|quod cum audisset Dominus ait ad me audivi vocem verborum populi huius quae locuti sunt tibi bene omnia sunt locuti
DEUT|5|29|quis det talem eos habere mentem ut timeant me et custodiant universa mandata mea in omni tempore ut bene sit eis et filiis eorum in sempiternum
DEUT|5|30|vade et dic eis revertimini in tentoria vestra
DEUT|5|31|tu vero hic sta mecum et loquar tibi omnia mandata et caerimonias atque iudicia quae docebis eos ut faciant ea in terra quam dabo illis in possessionem
DEUT|5|32|custodite igitur et facite quae praecepit Dominus Deus vobis non declinabitis neque ad dextram neque ad sinistram
DEUT|5|33|sed per viam quam praecepit Dominus Deus vester ambulabitis ut vivatis et bene sit vobis et protelentur dies in terra possessionis vestrae
DEUT|6|1|haec sunt praecepta et caerimoniae atque iudicia quae mandavit Dominus Deus vester ut docerem vos et faciatis ea in terra ad quam transgredimini possidendam
DEUT|6|2|ut timeas Dominum Deum tuum et custodias omnia mandata et praecepta eius quae ego praecipio tibi et filiis ac nepotibus tuis cunctis diebus vitae tuae ut prolongentur dies tui
DEUT|6|3|audi Israhel et observa ut facias et bene sit tibi et multipliceris amplius sicut pollicitus est Dominus Deus patrum tuorum tibi terram lacte et melle manantem
DEUT|6|4|audi Israhel Dominus Deus noster Dominus unus est
DEUT|6|5|diliges Dominum Deum tuum ex toto corde tuo et ex tota anima tua et ex tota fortitudine tua
DEUT|6|6|eruntque verba haec quae ego praecipio tibi hodie in corde tuo
DEUT|6|7|et narrabis ea filiis tuis et meditaberis sedens in domo tua et ambulans in itinere dormiens atque consurgens
DEUT|6|8|et ligabis ea quasi signum in manu tua eruntque et movebuntur inter oculos tuos
DEUT|6|9|scribesque ea in limine et ostiis domus tuae
DEUT|6|10|cumque introduxerit te Dominus Deus tuus in terram pro qua iuravit patribus tuis Abraham Isaac et Iacob et dederit tibi civitates magnas et optimas quas non aedificasti
DEUT|6|11|domos plenas cunctarum opum quas non extruxisti cisternas quas non fodisti vineta et oliveta quae non plantasti
DEUT|6|12|et comederis et saturatus fueris
DEUT|6|13|cave diligenter ne obliviscaris Domini qui eduxit te de terra Aegypti de domo servitutis Dominum Deum tuum timebis et ipsi servies ac per nomen illius iurabis
DEUT|6|14|non ibitis post deos alienos cunctarum gentium quae in circuitu vestro sunt
DEUT|6|15|quoniam Deus aemulator Dominus Deus tuus in medio tui nequando irascatur furor Domini Dei tui contra te et auferat te de superficie terrae
DEUT|6|16|non temptabis Dominum Deum tuum sicut temptasti in loco temptationis
DEUT|6|17|custodi praecepta Domini Dei tui ac testimonia et caerimonias quas praecepit tibi
DEUT|6|18|et fac quod placitum est et bonum in conspectu Domini ut bene sit tibi et ingressus possideas terram optimam de qua iuravit Dominus patribus tuis
DEUT|6|19|ut deleret omnes inimicos tuos coram te sicut locutus est
DEUT|6|20|cum interrogaverit te filius tuus cras dicens quid sibi volunt testimonia haec et caerimoniae atque iudicia quae praecepit Dominus Deus noster nobis
DEUT|6|21|dices ei servi eramus Pharaonis in Aegypto et eduxit nos Dominus de Aegypto in manu forti
DEUT|6|22|fecitque signa atque prodigia magna et pessima in Aegypto contra Pharaonem et omnem domum illius in conspectu nostro
DEUT|6|23|et eduxit nos inde ut introductis daret terram super qua iuravit patribus nostris
DEUT|6|24|praecepitque nobis Dominus ut faciamus omnia legitima haec et timeamus Dominum Deum nostrum et bene sit nobis cunctis diebus vitae nostrae sicut est hodie
DEUT|6|25|eritque nostri misericors si custodierimus et fecerimus omnia praecepta eius coram Domino Deo nostro sicut mandavit nobis
DEUT|7|1|cum introduxerit te Dominus Deus tuus in terram quam possessurus ingredieris et deleverit gentes multas coram te Hettheum et Gergeseum et Amorreum Chananeum et Ferezeum et Eveum et Iebuseum septem gentes multo maioris numeri quam tu es et robustiores te
DEUT|7|2|tradideritque eas Dominus Deus tuus tibi percuties eas usque ad internicionem non inibis cum eis foedus nec misereberis earum
DEUT|7|3|neque sociabis cum eis coniugia filiam tuam non dabis filio eius nec filiam illius accipies filio tuo
DEUT|7|4|quia seducet filium tuum ne sequatur me et ut magis serviat diis alienis irasceturque furor Domini et delebit te cito
DEUT|7|5|quin potius haec facietis eis aras eorum subvertite confringite statuas lucosque succidite et sculptilia conburite
DEUT|7|6|quia populus sanctus es Domino Deo tuo te elegit Dominus Deus tuus ut sis ei populus peculiaris de cunctis populis qui sunt super terram
DEUT|7|7|non quia cunctas gentes numero vincebatis vobis iunctus est Dominus et elegit vos cum omnibus sitis populis pauciores
DEUT|7|8|sed quia dilexit vos Dominus et custodivit iuramentum quod iuravit patribus vestris eduxitque vos in manu forti et redemit de domo servitutis de manu Pharaonis regis Aegypti
DEUT|7|9|et scies quia Dominus Deus tuus ipse est Deus fortis et fidelis custodiens pactum et misericordiam diligentibus se et his qui custodiunt praecepta eius in mille generationes
DEUT|7|10|et reddens odientibus se statim ita ut disperdat eos et ultra non differat protinus eis restituens quod merentur
DEUT|7|11|custodi ergo praecepta et caerimonias atque iudicia quae ego mando tibi hodie ut facias
DEUT|7|12|si postquam audieris haec iudicia custodieris ea et feceris custodiet et Dominus Deus tuus tibi pactum et misericordiam quam iuravit patribus tuis
DEUT|7|13|et diliget te ac multiplicabit benedicetque fructui ventris tui et fructui terrae tuae frumento tuo atque vindemiae oleo et armentis gregibus ovium tuarum super terram pro qua iuravit patribus tuis ut daret eam tibi
DEUT|7|14|benedictus eris inter omnes populos non erit apud te sterilis utriusque sexus tam in hominibus quam in gregibus tuis
DEUT|7|15|auferet Dominus a te omnem languorem et infirmitates Aegypti pessimas quas novisti non inferet tibi sed cunctis hostibus tuis
DEUT|7|16|devorabis omnes populos quos Dominus Deus tuus daturus est tibi non parcet eis oculus tuus nec servies diis eorum ne sint in ruinam tui
DEUT|7|17|si dixeris in corde tuo plures sunt gentes istae quam ego quomodo potero delere eas
DEUT|7|18|noli metuere sed recordare quae fecerit Dominus Deus tuus Pharaoni et cunctis Aegyptiis
DEUT|7|19|plagas maximas quas viderunt oculi tui et signa atque portenta manumque robustam et extentum brachium ut educeret te Dominus Deus tuus sic faciet cunctis populis quos metuis
DEUT|7|20|insuper et crabrones mittet Dominus Deus tuus in eos donec deleat omnes atque disperdat qui te fugerint et latere potuerint
DEUT|7|21|non timebis eos quia Dominus Deus tuus in medio tui est Deus magnus et terribilis
DEUT|7|22|ipse consumet nationes has in conspectu tuo paulatim atque per partes non poteris delere eas pariter ne forte multiplicentur contra te bestiae terrae
DEUT|7|23|dabitque eos Dominus Deus tuus in conspectu tuo et interficiet illos donec penitus deleantur
DEUT|7|24|tradet reges eorum in manus tuas et disperdes nomina eorum sub caelo nullus poterit resistere tibi donec conteras eos
DEUT|7|25|sculptilia eorum igne conbures non concupisces argentum et aurum de quibus facta sunt neque adsumes ex eis tibi quicquam ne offendas propter ea quia abominatio est Domini Dei tui
DEUT|7|26|nec inferes quippiam ex idolo in domum tuam ne fias anathema sicut et illud est quasi spurcitiam detestaberis et velut inquinamentum ac sordes abominationi habebis quia anathema est
DEUT|8|1|omne mandatum quod ego praecipio tibi hodie cave diligenter ut facias ut possitis vivere et multiplicemini ingressique possideatis terram pro qua iuravit Dominus patribus vestris
DEUT|8|2|et recordaberis cuncti itineris per quod adduxit te Dominus Deus tuus quadraginta annis per desertum ut adfligeret te atque temptaret et nota fierent quae in tuo animo versabantur utrum custodires mandata illius an non
DEUT|8|3|adflixit te penuria et dedit tibi cibum manna quem ignorabas tu et patres tui ut ostenderet tibi quod non in solo pane vivat homo sed in omni verbo quod egreditur ex ore Domini
DEUT|8|4|vestimentum tuum quo operiebaris nequaquam vetustate defecit et pes tuus non est subtritus en quadragesimus annus est
DEUT|8|5|ut recogites in corde tuo quia sicut erudit homo filium suum sic Dominus Deus tuus erudivit te
DEUT|8|6|ut custodias mandata Domini Dei tui et ambules in viis eius et timeas eum
DEUT|8|7|Dominus enim Deus tuus introducet te in terram bonam terram rivorum aquarumque et fontium in cuius campis et montibus erumpunt fluviorum abyssi
DEUT|8|8|terram frumenti hordei vinearum in qua ficus et mala granata et oliveta nascuntur terram olei ac mellis
DEUT|8|9|ubi absque ulla penuria comedes panem tuum et rerum omnium abundantia perfrueris cuius lapides ferrum sunt et de montibus eius aeris metalla fodiuntur
DEUT|8|10|ut cum comederis et satiatus fueris benedicas Domino Deo tuo pro terra optima quam dedit tibi
DEUT|8|11|observa et cave nequando obliviscaris Domini Dei tui et neglegas mandata eius atque iudicia et caerimonias quas ego praecipio tibi hodie
DEUT|8|12|ne postquam comederis et satiatus domos pulchras aedificaveris et habitaveris in eis
DEUT|8|13|habuerisque armenta et ovium greges argenti et auri cunctarumque rerum copiam
DEUT|8|14|elevetur cor tuum et non reminiscaris Domini Dei tui qui eduxit te de terra Aegypti de domo servitutis
DEUT|8|15|et ductor tuus fuit in solitudine magna atque terribili in qua erat serpens flatu adurens et scorpio ac dipsas et nullae omnino aquae qui eduxit rivos de petra durissima
DEUT|8|16|et cibavit te manna in solitudine quod nescierunt patres tui et postquam adflixit ac probavit ad extremum misertus est tui
DEUT|8|17|ne diceres in corde tuo fortitudo mea et robur manus meae haec mihi omnia praestiterunt
DEUT|8|18|sed recorderis Domini Dei tui quod ipse tibi vires praebuerit ut impleret pactum suum super quo iuravit patribus tuis sicut praesens indicat dies
DEUT|8|19|sin autem oblitus Domini Dei tui secutus fueris alienos deos coluerisque illos et adoraveris ecce nunc praedico tibi quod omnino dispereas
DEUT|8|20|sicut gentes quas delevit Dominus in introitu tuo ita et vos peribitis si inoboedientes fueritis voci Domini Dei vestri
DEUT|9|1|audi Israhel tu transgredieris hodie Iordanem ut possideas nationes maximas et fortiores te civitates ingentes et ad caelum usque muratas
DEUT|9|2|populum magnum atque sublimem filios Enacim quos ipse vidisti et audisti quibus nullus potest ex adverso resistere
DEUT|9|3|scies ergo hodie quod Dominus Deus tuus ipse transibit ante te ignis devorans atque consumens qui conterat eos et deleat atque disperdat ante faciem tuam velociter sicut locutus est tibi
DEUT|9|4|ne dicas in corde tuo cum deleverit eos Dominus Deus tuus in conspectu tuo propter iustitiam meam introduxit me Dominus ut terram hanc possiderem cum propter impietates suas istae deletae sint nationes
DEUT|9|5|neque enim propter iustitias tuas et aequitatem cordis tui ingredieris ut possideas terras eorum sed quia illae egerunt impie te introeunte deletae sunt et ut conpleret verbum suum Dominus quod sub iuramento pollicitus est patribus tuis Abraham Isaac et Iacob
DEUT|9|6|scito igitur quod non propter iustitias tuas Dominus Deus tuus dederit tibi terram hanc optimam in possessionem cum durissimae cervicis sis populus
DEUT|9|7|memento et ne obliviscaris quomodo ad iracundiam provocaveris Dominum Deum tuum in solitudine ex eo die quo es egressus ex Aegypto usque ad locum istum semper adversum Dominum contendisti
DEUT|9|8|nam et in Horeb provocasti eum et iratus delere te voluit
DEUT|9|9|quando ascendi in montem ut acciperem tabulas lapideas tabulas pacti quod pepigit vobiscum Dominus et perseveravi in monte quadraginta diebus ac noctibus panem non comedens et aquam non bibens
DEUT|9|10|deditque mihi Dominus duas tabulas lapideas scriptas digito Dei et continentes omnia verba quae vobis in monte locutus est de medio ignis quando contio populi congregata est
DEUT|9|11|cumque transissent quadraginta dies et totidem noctes dedit mihi Dominus duas tabulas lapideas tabulas foederis
DEUT|9|12|dixitque mihi surge et descende hinc cito quia populus tuus quos eduxisti de Aegypto deseruerunt velociter viam quam demonstrasti eis feceruntque sibi conflatile
DEUT|9|13|rursumque ait Dominus ad me cerno quod populus iste durae cervicis sit
DEUT|9|14|dimitte me ut conteram eum et deleam nomen eius sub caelo et constituam te super gentem quae hac maior et fortior sit
DEUT|9|15|cumque de monte ardente descenderem et duas tabulas foederis utraque tenerem manu
DEUT|9|16|vidissemque vos peccasse Domino Deo vestro et fecisse vobis vitulum conflatilem ac deseruisse velociter viam eius quam vobis ostenderat
DEUT|9|17|proieci tabulas de manibus meis confregique eas in conspectu vestro
DEUT|9|18|et procidi ante Dominum sicut prius quadraginta diebus et noctibus panem non comedens et aquam non bibens propter omnia peccata vestra quae gessistis contra Dominum et eum ad iracundiam provocastis
DEUT|9|19|timui enim indignationem et iram illius qua adversum vos concitatus delere vos voluit et exaudivit me Dominus etiam hac vice
DEUT|9|20|adversum Aaron quoque vehementer iratus voluit eum conterere et pro illo similiter deprecatus sum
DEUT|9|21|peccatum autem vestrum quod feceratis id est vitulum arripiens igne conbusi et in frusta comminuens omninoque in pulverem redigens proieci in torrentem qui de monte descendit
DEUT|9|22|in Incendio quoque et in Temptatione et in sepulchris Concupiscentiae provocastis Dominum
DEUT|9|23|et quando misit vos de Cadesbarne dicens ascendite et possidete terram quam dedi vobis et contempsistis imperium Domini Dei vestri et non credidistis ei neque vocem eius audire voluistis
DEUT|9|24|sed semper fuistis rebelles a die qua nosse vos coepi
DEUT|9|25|et iacui coram Domino quadraginta diebus ac noctibus quibus eum suppliciter deprecabar ne deleret vos ut fuerat comminatus
DEUT|9|26|et orans dixi Domine Deus ne disperdas populum tuum et hereditatem tuam quam redemisti in magnitudine tua quos eduxisti de Aegypto in manu forti
DEUT|9|27|recordare servorum tuorum Abraham Isaac et Iacob ne aspicias duritiam populi huius et impietatem atque peccatum
DEUT|9|28|ne forte dicant habitatores terrae de qua eduxisti nos non poterat Dominus introducere eos in terram quam pollicitus est eis et oderat illos idcirco eduxit ut interficeret eos in solitudine
DEUT|9|29|qui sunt populus tuus et hereditas tua quos eduxisti in fortitudine tua magna et in brachio tuo extento
DEUT|10|1|in tempore illo dixit Dominus ad me dola tibi duas tabulas lapideas sicut priores fuerunt et ascende ad me in montem faciesque arcam ligneam
DEUT|10|2|et scribam in tabulis verba quae fuerunt in his quas ante confregisti ponesque eas in arca
DEUT|10|3|feci igitur arcam de lignis setthim cumque dolassem duas tabulas lapideas instar priorum ascendi in montem habens eas in manibus
DEUT|10|4|scripsitque in tabulis iuxta id quod prius scripserat verba decem quae locutus est Dominus ad vos in monte de medio ignis quando populus congregatus est et dedit eas mihi
DEUT|10|5|reversusque de monte descendi et posui tabulas in arcam quam feceram quae hucusque ibi sunt sicut mihi praecepit Dominus
DEUT|10|6|filii autem Israhel castra moverunt ex Beroth filiorum Iacan in Musera ubi Aaron mortuus ac sepultus est pro quo sacerdotio functus est filius eius Eleazar
DEUT|10|7|inde venerunt in Gadgad de quo loco profecti castrametati sunt in Ietabatha in terra aquarum atque torrentium
DEUT|10|8|eo tempore separavit tribum Levi ut portaret arcam foederis Domini et staret coram eo in ministerio ac benediceret in nomine illius usque in praesentem diem
DEUT|10|9|quam ob rem non habuit Levi partem neque possessionem cum fratribus suis quia ipse Dominus possessio eius est sicut promisit ei Dominus Deus tuus
DEUT|10|10|ego autem steti in monte sicut prius quadraginta diebus ac noctibus exaudivitque me Dominus etiam hac vice et te perdere noluit
DEUT|10|11|dixitque mihi vade et praecede populum ut ingrediatur et possideat terram quam iuravi patribus eorum ut traderem eis
DEUT|10|12|et nunc Israhel quid Dominus Deus tuus petit a te nisi ut timeas Dominum Deum tuum et ambules in viis eius et diligas eum ac servias Domino Deo tuo in toto corde tuo et in tota anima tua
DEUT|10|13|custodiasque mandata Domini et caerimonias eius quas ego hodie praecipio ut bene sit tibi
DEUT|10|14|en Domini Dei tui caelum est et caelum caeli terra et omnia quae in ea sunt
DEUT|10|15|et tamen patribus tuis conglutinatus est Dominus et amavit eos elegitque semen eorum post eos id est vos de cunctis gentibus sicut hodie conprobatur
DEUT|10|16|circumcidite igitur praeputium cordis vestri et cervicem vestram ne induretis amplius
DEUT|10|17|quia Dominus Deus vester ipse est Deus deorum et Dominus dominantium Deus magnus et potens et terribilis qui personam non accipit nec munera
DEUT|10|18|facit iudicium pupillo et viduae amat peregrinum et dat ei victum atque vestitum
DEUT|10|19|et vos ergo amate peregrinos quia et ipsi fuistis advenae in terra Aegypti
DEUT|10|20|Dominum Deum tuum timebis et ei servies ipsi adherebis iurabisque in nomine illius
DEUT|10|21|ipse est laus tua et Deus tuus qui fecit tibi haec magnalia et terribilia quae viderunt oculi tui
DEUT|10|22|in septuaginta animabus descenderunt patres tui in Aegyptum et ecce nunc multiplicavit te Dominus Deus tuus sicut astra caeli
DEUT|11|1|ama itaque Dominum Deum tuum et observa praecepta eius et caerimonias iudicia atque mandata omni tempore
DEUT|11|2|cognoscite hodie quae ignorant filii vestri qui non viderunt disciplinam Domini Dei vestri magnalia eius et robustam manum extentumque brachium
DEUT|11|3|signa et opera quae fecit in medio Aegypti Pharaoni regi et universae terrae eius
DEUT|11|4|omnique exercitui Aegyptiorum et equis ac curribus quomodo operuerint eos aquae Rubri maris cum vos persequerentur et deleverit eos Dominus usque in praesentem diem
DEUT|11|5|vobisque quae fecerit in solitudine donec veniretis ad hunc locum
DEUT|11|6|et Dathan atque Abiram filiis Heliab qui fuit filius Ruben quos aperto ore suo terra absorbuit cum domibus et tabernaculis et universa substantia eorum quam habebant in medio Israhelis
DEUT|11|7|oculi vestri viderunt omnia opera Domini magna quae fecit
DEUT|11|8|ut custodiatis universa mandata illius quae ego hodie praecipio vobis et possitis introire et possidere terram ad quam ingredimini
DEUT|11|9|multoque in ea vivatis tempore quam sub iuramento pollicitus est Dominus patribus vestris et semini eorum lacte et melle manantem
DEUT|11|10|terra enim ad quam ingredieris possidendam non est sicut terra Aegypti de qua existi ubi iacto semine in hortorum morem aquae ducuntur inriguae
DEUT|11|11|sed montuosa est et campestris de caelo expectans pluvias
DEUT|11|12|quam Dominus Deus tuus semper invisit et oculi illius in ea sunt a principio anni usque ad finem eius
DEUT|11|13|si ergo oboedieritis mandatis meis quae hodie praecipio vobis ut diligatis Dominum Deum vestrum et serviatis ei in toto corde vestro et in tota anima vestra
DEUT|11|14|dabo pluviam terrae vestrae temporivam et serotinam ut colligatis frumentum et vinum et oleum
DEUT|11|15|faenum ex agris ad pascenda iumenta et ut ipsi comedatis ac saturemini
DEUT|11|16|cavete ne forte decipiatur cor vestrum et recedatis a Domino serviatisque diis alienis et adoretis eos
DEUT|11|17|iratusque Dominus claudat caelum et pluviae non descendant nec terra det germen suum pereatisque velociter de terra optima quam Dominus daturus est vobis
DEUT|11|18|ponite haec verba mea in cordibus et in animis vestris et suspendite ea pro signo in manibus et inter vestros oculos conlocate
DEUT|11|19|docete filios vestros ut illa meditentur quando sederis in domo tua et ambulaveris in via et accubueris atque surrexeris
DEUT|11|20|scribes ea super postes et ianuas domus tuae
DEUT|11|21|ut multiplicentur dies tui et filiorum tuorum in terra quam iuravit Dominus patribus tuis ut daret eis quamdiu caelum inminet terrae
DEUT|11|22|si enim custodieritis mandata quae ego praecipio vobis et feceritis ea ut diligatis Dominum Deum vestrum et ambuletis in omnibus viis eius adherentes ei
DEUT|11|23|disperdet Dominus omnes gentes istas ante faciem vestram et possidebitis eas quae maiores et fortiores vobis sunt
DEUT|11|24|omnis locus quem calcaverit pes vester vester erit a deserto et Libano a flumine magno Eufraten usque ad mare occidentale erunt termini vestri
DEUT|11|25|nullus stabit contra vos terrorem vestrum et formidinem dabit Dominus Deus vester super omnem terram quam calcaturi estis sicut locutus est vobis
DEUT|11|26|en propono in conspectu vestro hodie benedictionem et maledictionem
DEUT|11|27|benedictionem si oboedieritis mandatis Domini Dei vestri quae ego praecipio vobis
DEUT|11|28|maledictionem si non audieritis mandata Domini Dei vestri sed recesseritis de via quam ego nunc ostendo vobis et ambulaveritis post deos alienos quos ignoratis
DEUT|11|29|cum introduxerit te Dominus Deus tuus in terram ad quam pergis habitandam pones benedictionem super montem Garizim maledictionem super montem Hebal
DEUT|11|30|qui sunt trans Iordanem post viam quae vergit ad solis occubitum in terra Chananei qui habitat in campestribus contra Galgalam quae est iuxta vallem tendentem et intrantem procul
DEUT|11|31|vos enim transibitis Iordanem ut possideatis terram quam Dominus Deus vester daturus est vobis et habeatis ac possideatis illam
DEUT|11|32|videte ergo ut impleatis caerimonias atque iudicia quae ego hodie ponam in conspectu vestro
DEUT|12|1|haec sunt praecepta atque iudicia quae facere debetis in terra quam Dominus Deus patrum tuorum daturus est tibi ut possideas eam cunctis diebus quibus super humum gradieris
DEUT|12|2|subvertite omnia loca in quibus coluerunt gentes quas possessuri estis deos suos super montes excelsos et colles et subter omne lignum frondosum
DEUT|12|3|dissipate aras earum et confringite statuas lucos igne conburite et idola comminuite disperdite nomina eorum de locis illis
DEUT|12|4|non facietis ita Domino Deo vestro
DEUT|12|5|sed ad locum quem elegerit Dominus Deus vester de cunctis tribubus vestris ut ponat nomen suum ibi et habitet in eo venietis
DEUT|12|6|et offeretis in illo loco holocausta et victimas vestras decimas et primitias manuum vestrarum et vota atque donaria primogenita boum et ovium
DEUT|12|7|et comedetis ibi in conspectu Domini Dei vestri ac laetabimini in cunctis ad quae miseritis manum vos et domus vestrae in quibus benedixerit vobis Dominus Deus vester
DEUT|12|8|non facietis ibi quae nos hic facimus hodie singuli quod sibi rectum videtur
DEUT|12|9|neque enim usque in praesens tempus venistis ad requiem et possessionem quam Dominus Deus daturus est vobis
DEUT|12|10|transibitis Iordanem et habitabitis in terram quam Dominus Deus vester daturus est vobis ut requiescatis a cunctis hostibus per circuitum et absque ullo timore habitetis
DEUT|12|11|in loco quem elegerit Dominus Deus vester ut sit nomen eius in eo illuc omnia quae praecipio conferetis holocausta et hostias ac decimas et primitias manuum vestrarum et quicquid praecipuum est in muneribus quae vovistis Domino
DEUT|12|12|ibi epulabimini coram Domino Deo vestro vos filii ac filiae vestrae famuli et famulae atque Levites qui in vestris urbibus commorantur neque enim habet aliam partem et possessionem inter vos
DEUT|12|13|cave ne offeras holocausta tua in omni loco quem videris
DEUT|12|14|sed in eo quem elegerit Dominus in una tribuum tuarum offeres hostias et facies quaecumque praecipio tibi
DEUT|12|15|sin autem comedere volueris et te esus carnium delectarit occide et comede iuxta benedictionem Domini Dei tui quam dedit tibi in urbibus tuis sive inmundum fuerit hoc est maculatum et debile sive mundum hoc est integrum et sine macula quod offerri licet sicut capream et cervum comedes
DEUT|12|16|absque esu dumtaxat sanguinis quod super terram quasi aquam effundes
DEUT|12|17|non poteris comedere in oppidis tuis decimam frumenti et vini et olei tui primogenita armentorum et pecorum et omnia quae voveris et sponte offerre volueris et primitias manuum tuarum
DEUT|12|18|sed coram Domino Deo tuo comedes ea in loco quem elegerit Dominus Deus tuus tu et filius tuus ac filia servus et famula atque Levites qui manet in urbibus tuis et laetaberis et reficieris coram Domino Deo tuo in cunctis ad quae extenderis manum tuam
DEUT|12|19|cave ne derelinquas Leviten omni tempore quo versaris in terra
DEUT|12|20|quando dilataverit Dominus Deus tuus terminos tuos sicut locutus est tibi et volueris vesci carnibus quas desiderat anima tua
DEUT|12|21|locus autem quem elegerit Dominus Deus tuus ut sit nomen eius ibi si procul fuerit occides de armentis et pecoribus quae habueris sicut praecepi tibi et comedes in oppidis tuis ut tibi placet
DEUT|12|22|sicut comeditur caprea et cervus ita vesceris eis et mundus et inmundus in commune vescentur
DEUT|12|23|hoc solum cave ne sanguinem comedas sanguis enim eorum pro anima est et idcirco non debes animam comedere cum carnibus
DEUT|12|24|sed super terram fundes quasi aquam
DEUT|12|25|ut sit tibi bene et filiis tuis post te cum feceris quod placet in conspectu Domini
DEUT|12|26|quae autem sanctificaveris et voveris Domino tolles et venies ad locum quem elegerit Dominus
DEUT|12|27|et offeres oblationes tuas carnem et sanguinem super altare Domini Dei tui sanguinem hostiarum fundes in altari carnibus autem ipse vesceris
DEUT|12|28|observa et audi omnia quae ego praecipio tibi ut bene sit tibi et filiis tuis post te in sempiternum cum feceris quod bonum est et placitum in conspectu Domini Dei tui
DEUT|12|29|quando disperderit Dominus Deus tuus ante faciem tuam gentes ad quas ingredieris possidendas et possederis eas atque habitaveris in terra earum
DEUT|12|30|cave ne imiteris eas postquam te fuerint introeunte subversae et requiras caerimonias earum dicens sicut coluerunt gentes istae deos suos ita et ego colam
DEUT|12|31|non facies similiter Domino Deo tuo omnes enim abominationes quas aversatur Dominus fecerunt diis suis offerentes filios et filias et conburentes igne
DEUT|12|32|quod praecipio tibi hoc tantum facito Domino nec addas quicquam nec minuas
DEUT|13|1|si surrexerit in medio tui prophetes aut qui somnium vidisse se dicat et praedixerit signum atque portentum
DEUT|13|2|et evenerit quod locutus est et dixerit tibi eamus et sequamur deos alienos quos ignoras et serviamus eis
DEUT|13|3|non audies verba prophetae illius aut somniatoris quia temptat vos Dominus Deus vester ut palam fiat utrum diligatis eum an non in toto corde et in tota anima vestra
DEUT|13|4|Dominum Deum vestrum sequimini et ipsum timete mandata illius custodite et audite vocem eius ipsi servietis et ipsi adherebitis
DEUT|13|5|propheta autem ille aut fictor somniorum interficietur quia locutus est ut vos averteret a Domino Deo vestro qui eduxit vos de terra Aegypti et redemit de domo servitutis ut errare te faceret de via quam tibi praecepit Dominus Deus tuus et auferes malum de medio tui
DEUT|13|6|si tibi voluerit persuadere frater tuus filius matris tuae aut filius tuus vel filia sive uxor quae est in sinu tuo aut amicus quem diligis ut animam tuam clam dicens eamus et serviamus diis alienis quos ignoras tu et patres tui
DEUT|13|7|cunctarum in circuitu gentium quae iuxta vel procul sunt ab initio usque ad finem terrae
DEUT|13|8|non adquiescas ei nec audias neque parcat ei oculus tuus ut miserearis et occultes eum
DEUT|13|9|sed statim interficies sit primum manus tua super eum et post te omnis populus mittat manum
DEUT|13|10|lapidibus obrutus necabitur quia voluit te abstrahere a Domino Deo tuo qui eduxit te de terra Aegypti de domo servitutis
DEUT|13|11|ut omnis Israhel audiens timeat et nequaquam ultra faciat quippiam huius rei simile
DEUT|13|12|si audieris in una urbium tuarum quas Dominus Deus tuus dabit tibi ad habitandum dicentes aliquos
DEUT|13|13|egressi sunt filii Belial de medio tui et averterunt habitatores urbis tuae atque dixerunt eamus et serviamus diis alienis quos ignoratis
DEUT|13|14|quaere sollicite et diligenter rei veritate perspecta si inveneris certum esse quod dicitur et abominationem hanc opere perpetratam
DEUT|13|15|statim percuties habitatores urbis illius in ore gladii et delebis eam omniaque quae in illa sunt usque ad pecora
DEUT|13|16|quicquid etiam supellectilis fuerit congregabis in medium platearum eius et cum ipsa civitate succendes ita ut universa consumas Domino Deo tuo et sit tumulus sempiternus non aedificabitur amplius
DEUT|13|17|et non adherebit de illo anathemate quicquam in manu tua ut avertatur Dominus ab ira furoris sui et misereatur tui multiplicetque te sicut iuravit patribus tuis
DEUT|13|18|quando audieris vocem Domini Dei tui custodiens omnia praecepta eius quae ego praecipio tibi hodie ut facias quod placitum est in conspectu Domini Dei tui
DEUT|13|19|
DEUT|14|1|filii estote Domini Dei vestri non vos incidetis nec facietis calvitium super mortuo
DEUT|14|2|quoniam populus sanctus es Domino Deo tuo et te elegit ut sis ei in populum peculiarem de cunctis gentibus quae sunt super terram
DEUT|14|3|ne comedatis quae inmunda sunt
DEUT|14|4|hoc est animal quod comedere debetis bovem et ovem et capram
DEUT|14|5|cervum capream bubalum tragelaphum pygargon orygem camelopardalum
DEUT|14|6|omne animal quod in duas partes ungulam findit et ruminat comedetis
DEUT|14|7|de his autem quae ruminant et ungulam non findunt haec comedere non debetis camelum leporem choerogyllium quia ruminant et non dividunt ungulam inmunda erunt vobis
DEUT|14|8|sus quoque quoniam dividit ungulam et non ruminat inmunda erit carnibus eorum non vescemini et cadavera non tangetis
DEUT|14|9|haec comedetis ex omnibus quae morantur in aquis quae habent pinnulas et squamas comedite
DEUT|14|10|quae absque pinnulis et squamis sunt ne comedatis quia inmunda sunt
DEUT|14|11|omnes aves mundas comedite
DEUT|14|12|inmundas ne comedatis aquilam scilicet et grypem et alietum
DEUT|14|13|ixon et vulturem ac milvum iuxta genus suum
DEUT|14|14|et omne corvini generis
DEUT|14|15|strutionem ac noctuam et larum atque accipitrem iuxta genus suum
DEUT|14|16|herodium et cycnum et ibin
DEUT|14|17|ac mergulum porphirionem et nycticoracem
DEUT|14|18|onocrotalum et charadrium singula in genere suo upupam quoque et vespertilionem
DEUT|14|19|et omne quod reptat et pinnulas habet inmundum erit nec comedetur
DEUT|14|20|omne quod mundum est comedite
DEUT|14|21|quicquid morticinum est ne vescamini ex eo peregrino qui intra portas tuas est da ut comedat aut vende ei quia tu populus sanctus Domini Dei tui es non coques hedum in lacte matris suae
DEUT|14|22|decimam partem separabis de cunctis frugibus tuis quae nascuntur in terra per annos singulos
DEUT|14|23|et comedes in conspectu Domini Dei tui in loco quem elegerit ut in eo nomen illius invocetur decimam frumenti tui et vini et olei et primogenita de armentis et ovibus tuis ut discas timere Dominum Deum tuum omni tempore
DEUT|14|24|cum autem longior fuerit via et locus quem elegerit Dominus Deus tuus tibique benedixerit nec potueris ad eum haec cuncta portare
DEUT|14|25|vendes omnia et in pretium rediges portabisque manu tua et proficisceris ad locum quem elegerit Dominus Deus tuus
DEUT|14|26|et emes ex eadem pecunia quicquid tibi placuerit sive ex armentis sive ex ovibus vinum quoque et siceram et omne quod desiderat anima tua et comedes coram Domino Deo tuo et epulaberis tu et domus tua
DEUT|14|27|et Levita qui intra portas tuas est cave ne derelinquas eum quia non habet aliam partem in possessione tua
DEUT|14|28|anno tertio separabis aliam decimam ex omnibus quae nascuntur tibi eo tempore et repones intra ianuas tuas
DEUT|14|29|venietque Levites qui aliam non habet partem nec possessionem tecum et peregrinus et pupillus ac vidua qui intra portas tuas sunt et comedent et saturabuntur ut benedicat tibi Dominus Deus tuus in cunctis operibus manuum tuarum quae feceris
DEUT|15|1|septimo anno facies remissionem
DEUT|15|2|quae hoc ordine celebrabitur cui debetur aliquid ab amico vel proximo ac fratre suo repetere non poterit quia annus remissionis est Domini
DEUT|15|3|a peregrino et advena exiges civem et propinquum repetendi non habes potestatem
DEUT|15|4|et omnino indigens et mendicus non erit inter vos ut benedicat tibi Dominus in terra quam traditurus est tibi in possessionem
DEUT|15|5|si tamen audieris vocem Domini Dei tui et custodieris universa quae iussit et quae ego hodie praecipio tibi benedicet tibi ut pollicitus est
DEUT|15|6|fenerabis gentibus multis et ipse a nullo accipies mutuum dominaberis nationibus plurimis et tui nemo dominabitur
DEUT|15|7|si unus de fratribus tuis qui morantur intra portas civitatis tuae in terra quam Dominus Deus tuus daturus est tibi ad paupertatem venerit non obdurabis cor tuum nec contrahes manum
DEUT|15|8|sed aperies eam pauperi et dabis mutuum quod eum indigere perspexeris
DEUT|15|9|cave ne forte subripiat tibi impia cogitatio et dicas in corde tuo adpropinquat septimus annus remissionis et avertas oculos a paupere fratre tuo nolens ei quod postulat mutuum commodare ne clamet contra te ad Dominum et fiat tibi in peccatum
DEUT|15|10|sed dabis ei nec ages quippiam callide in eius necessitatibus sublevandis ut benedicat tibi Dominus Deus tuus in omni tempore et in cunctis ad quae manum miseris
DEUT|15|11|non deerunt pauperes in terra habitationis tuae idcirco ego praecipio tibi ut aperias manum fratri tuo egeno et pauperi qui tecum versatur in terra
DEUT|15|12|cum tibi venditus fuerit frater tuus hebraeus aut hebraea et sex annis servierit tibi in septimo anno dimittes eum liberum
DEUT|15|13|et quem libertate donaveris nequaquam vacuum abire patieris
DEUT|15|14|sed dabis viaticum de gregibus et de area et torculari tuo quibus Dominus Deus tuus benedixerit tibi
DEUT|15|15|memento quod et ipse servieris in terra Aegypti et liberaverit te Dominus Deus tuus et idcirco ego nunc praecipiam tibi
DEUT|15|16|sin autem dixerit nolo egredi eo quod diligat te et domum tuam et bene sibi apud te esse sentiat
DEUT|15|17|adsumes subulam et perforabis aurem eius in ianua domus tuae et serviet tibi usque in aeternum ancillae quoque similiter facies
DEUT|15|18|non avertes ab eis oculos tuos quando dimiseris eos liberos quoniam iuxta mercedem mercennarii per sex annos servivit tibi ut benedicat tibi Dominus Deus tuus in cunctis operibus quae agis
DEUT|15|19|de primogenitis quae nascuntur in armentis et ovibus tuis quicquid sexus est masculini sanctificabis Domino Deo tuo non operaberis in primogenito bovis et non tondebis primogenita ovium
DEUT|15|20|in conspectu Domini Dei tui comedes ea per annos singulos in loco quem elegerit Dominus tu et domus tua
DEUT|15|21|sin autem habuerit maculam et vel claudum fuerit vel caecum aut in aliqua parte deforme vel debile non immolabitur Domino Deo tuo
DEUT|15|22|sed intra portas urbis tuae comedes illud tam mundus quam inmundus similiter vescentur eis quasi caprea et cervo
DEUT|15|23|hoc solum observabis ut sanguinem eorum non comedas sed effundas in terram quasi aquam
DEUT|16|1|observa mensem novarum frugum et verni primum temporis ut facias phase Domino Deo tuo quoniam in isto mense eduxit te Dominus Deus tuus de Aegypto nocte
DEUT|16|2|immolabisque phase Domino Deo tuo de ovibus et de bubus in loco quem elegerit Dominus Deus tuus ut habitet nomen eius ibi
DEUT|16|3|non comedes in eo panem fermentatum septem diebus comedes absque fermento adflictionis panem quoniam in pavore egressus es de Aegypto ut memineris diei egressionis tuae de Aegypto omnibus diebus vitae tuae
DEUT|16|4|non apparebit fermentum in omnibus terminis tuis septem diebus et non manebit de carnibus eius quod immolatum est vesperi in die primo mane
DEUT|16|5|non poteris immolare phase in qualibet urbium tuarum quas Dominus Deus tuus daturus est tibi
DEUT|16|6|sed in loco quem elegerit Dominus Deus tuus ut habitet nomen eius ibi immolabis phase vesperi ad solis occasum quando egressus es de Aegypto
DEUT|16|7|et coques et comedes in loco quem elegerit Dominus Deus tuus maneque consurgens vades in tabernacula tua
DEUT|16|8|sex diebus comedes azyma et in die septimo quia collecta est Domini Dei tui non facies opus
DEUT|16|9|septem ebdomadas numerabis tibi ab ea die qua falcem in segetem miseris
DEUT|16|10|et celebrabis diem festum ebdomadarum Domino Deo tuo oblationem spontaneam manus tuae quam offeres iuxta benedictionem Domini Dei tui
DEUT|16|11|et epulaberis coram Domino Deo tuo tu et filius tuus et filia tua et servus tuus et ancilla et Levites qui est intra portas tuas et advena ac pupillus et vidua qui morantur vobiscum in loco quem elegerit Dominus Deus tuus ut habitet nomen eius ibi
DEUT|16|12|et recordaberis quoniam servus fueris in Aegypto custodiesque ac facies quae praecepta sunt
DEUT|16|13|sollemnitatem quoque tabernaculorum celebrabis per septem dies quando collegeris de area et torculari fruges tuas
DEUT|16|14|et epulaberis in festivitate tua tu et filius tuus et filia et servus tuus et ancilla Levites quoque et advena et pupillus ac vidua qui intra portas tuas sunt
DEUT|16|15|septem diebus Domino Deo tuo festa celebrabis in loco quem elegerit Dominus benedicetque tibi Dominus Deus tuus in cunctis frugibus tuis et in omni opere manuum tuarum erisque in laetitia
DEUT|16|16|tribus vicibus per annum apparebit omne masculinum tuum in conspectu Domini Dei tui in loco quem elegerit in sollemnitate azymorum et in sollemnitate ebdomadarum et in sollemnitate tabernaculorum non apparebit ante Dominum vacuus
DEUT|16|17|sed offeret unusquisque secundum quod habuerit iuxta benedictionem Domini Dei sui quam dederit ei
DEUT|16|18|iudices et magistros constitues in omnibus portis tuis quas Dominus Deus tuus dederit tibi per singulas tribus tuas ut iudicent populum iusto iudicio
DEUT|16|19|nec in alteram partem declinent non accipies personam nec munera quia munera excaecant oculos sapientium et mutant verba iustorum
DEUT|16|20|iuste quod iustum est persequeris ut vivas et possideas terram quam Dominus Deus tuus dederit tibi
DEUT|16|21|non plantabis lucum et omnem arborem iuxta altare Domini Dei tui
DEUT|16|22|nec facies tibi atque constitues statuam quae odit Dominus Deus tuus
DEUT|17|1|non immolabis Domino Deo tuo bovem et ovem in quo est macula aut quippiam vitii quia abominatio est Domini Dei tui
DEUT|17|2|cum repperti fuerint apud te intra unam portarum tuarum quas Dominus Deus tuus dabit tibi vir aut mulier qui faciant malum in conspectu Domini Dei tui et transgrediantur pactum illius
DEUT|17|3|ut vadant et serviant diis alienis et adorent eos solem et lunam et omnem militiam caeli quae non praecepi
DEUT|17|4|et hoc tibi fuerit nuntiatum audiensque inquisieris diligenter et verum esse reppereris et abominatio facta est in Israhel
DEUT|17|5|educes virum ac mulierem qui rem sceleratissimam perpetrarunt ad portas civitatis tuae et lapidibus obruentur
DEUT|17|6|in ore duorum aut trium testium peribit qui interficietur nemo occidatur uno contra se dicente testimonium
DEUT|17|7|manus testium prima interficiet eum et manus reliqui populi extrema mittetur ut auferas malum de medio tui
DEUT|17|8|si difficile et ambiguum apud te iudicium esse perspexeris inter sanguinem et sanguinem causam et causam lepram et non lepram et iudicum intra portas tuas videris verba variari surge et ascende ad locum quem elegerit Dominus Deus tuus
DEUT|17|9|veniesque ad sacerdotes levitici generis et ad iudicem qui fuerit illo tempore quaeresque ab eis qui indicabunt tibi iudicii veritatem
DEUT|17|10|et facies quodcumque dixerint qui praesunt loco quem elegerit Dominus et docuerint te
DEUT|17|11|iuxta legem eius sequeris sententiam eorum nec declinabis ad dextram vel ad sinistram
DEUT|17|12|qui autem superbierit nolens oboedire sacerdotis imperio qui eo tempore ministrat Domino Deo tuo et decreto iudicis morietur homo ille et auferes malum de Israhel
DEUT|17|13|cunctusque populus audiens timebit ut nullus deinceps intumescat superbia
DEUT|17|14|cum ingressus fueris terram quam Dominus Deus tuus dabit tibi et possederis eam habitaverisque in illa et dixeris constituam super me regem sicut habent omnes per circuitum nationes
DEUT|17|15|eum constitues quem Dominus Deus tuus elegerit de numero fratrum tuorum non poteris alterius gentis hominem regem facere qui non sit frater tuus
DEUT|17|16|cumque fuerit constitutus non multiplicabit sibi equos nec reducet populum in Aegyptum equitatus numero sublevatus praesertim cum Dominus praeceperit vobis ut nequaquam amplius per eandem viam revertamini
DEUT|17|17|non habebit uxores plurimas quae inliciant animum eius neque argenti et auri inmensa pondera
DEUT|17|18|postquam autem sederit in solio regni sui describet sibi deuteronomium legis huius in volumine accipiens exemplar a sacerdotibus leviticae tribus
DEUT|17|19|et habebit secum legetque illud omnibus diebus vitae suae ut discat timere Dominum Deum suum et custodire verba et caerimonias eius quae lege praecepta sunt
DEUT|17|20|nec elevetur cor eius in superbiam super fratres suos neque declinet in partem dextram vel sinistram ut longo tempore regnet ipse et filii eius super Israhel
DEUT|18|1|non habebunt sacerdotes et Levitae et omnes qui de eadem tribu sunt partem et hereditatem cum reliquo Israhel quia sacrificia Domini et oblationes eius comedent
DEUT|18|2|et nihil aliud accipient de possessione fratrum suorum Dominus enim ipse est hereditas eorum sicut locutus est illis
DEUT|18|3|hoc erit iudicium sacerdotum a populo et ab his qui offerunt victimas sive bovem sive ovem immolaverint dabunt sacerdoti armum ac ventriculum
DEUT|18|4|primitias frumenti vini et olei et lanarum partem ex ovium tonsione
DEUT|18|5|ipsum enim elegit Dominus Deus tuus de cunctis tribubus tuis ut stet et ministret nomini Domini ipse et filii eius in sempiternum
DEUT|18|6|si exierit Levites de una urbium tuarum ex omni Israhel in qua habitat et voluerit venire desiderans locum quem elegerit Dominus
DEUT|18|7|ministrabit in nomine Dei sui sicut omnes fratres eius Levitae qui stabunt eo tempore coram Domino
DEUT|18|8|partem ciborum eandem accipiet quam et ceteri excepto eo quod in urbe sua ex paterna ei successione debetur
DEUT|18|9|quando ingressus fueris terram quam Dominus Deus tuus dabit tibi cave ne imitari velis abominationes illarum gentium
DEUT|18|10|nec inveniatur in te qui lustret filium suum aut filiam ducens per ignem aut qui ariolos sciscitetur et observet somnia atque auguria ne sit maleficus
DEUT|18|11|ne incantator ne pythones consulat ne divinos et quaerat a mortuis veritatem
DEUT|18|12|omnia enim haec abominatur Dominus et propter istiusmodi scelera delebit eos in introitu tuo
DEUT|18|13|perfectus eris et absque macula cum Domino Deo tuo
DEUT|18|14|gentes istae quarum possidebis terram augures et divinos audiunt tu autem a Domino Deo tuo aliter institutus es
DEUT|18|15|prophetam de gente tua et de fratribus tuis sicut me suscitabit tibi Dominus Deus tuus ipsum audies
DEUT|18|16|ut petisti a Domino Deo tuo in Horeb quando contio congregata est atque dixisti ultra non audiam vocem Domini Dei mei et ignem hunc maximum amplius non videbo ne moriar
DEUT|18|17|et ait Dominus mihi bene omnia sunt locuti
DEUT|18|18|prophetam suscitabo eis de medio fratrum suorum similem tui et ponam verba mea in ore eius loqueturque ad eos omnia quae praecepero illi
DEUT|18|19|qui autem verba eius quae loquetur in nomine meo audire noluerit ego ultor existam
DEUT|18|20|propheta autem qui arrogantia depravatus voluerit loqui in nomine meo quae ego non praecepi illi ut diceret aut ex nomine alienorum deorum interficietur
DEUT|18|21|quod si tacita cogitatione responderis quomodo possum intellegere verbum quod non est locutus Dominus
DEUT|18|22|hoc habebis signum quod in nomine Domini propheta ille praedixerit et non evenerit hoc Dominus non locutus est sed per tumorem animi sui propheta confinxit et idcirco non timebis eum
DEUT|19|1|cum disperderit Dominus Deus tuus gentes quarum tibi traditurus est terram et possederis eam habitaverisque in urbibus eius et in aedibus
DEUT|19|2|tres civitates separabis tibi in medio terrae quam Dominus Deus tuus dabit tibi in possessionem
DEUT|19|3|sternens diligenter viam et in tres aequaliter partes totam terrae tuae provinciam divides ut habeat e vicino qui propter homicidium profugus est quo possit evadere
DEUT|19|4|haec erit lex homicidae fugientis cuius vita servanda est qui percusserit proximum suum nesciens et qui heri et nudius tertius nullum contra eum habuisse odium conprobatur
DEUT|19|5|sed abisse simpliciter cum eo in silvam ad ligna caedenda et in succisione lignorum securis fugerit manu ferrumque lapsum de manubrio amicum eius percusserit et occiderit hic ad unam supradictarum urbium confugiet et vivet
DEUT|19|6|ne forsitan proximus eius cuius effusus est sanguis dolore stimulatus persequatur et adprehendat eum si longior via fuerit et percutiat animam eius qui non est reus mortis quia nullum contra eum qui occisus est odium prius habuisse monstratur
DEUT|19|7|idcirco praecipio tibi ut tres civitates aequalis inter se spatii dividas
DEUT|19|8|cum autem dilataverit Dominus Deus tuus terminos tuos sicut iuravit patribus tuis et dederit tibi cunctam terram quam eis pollicitus est
DEUT|19|9|si tamen custodieris mandata eius et feceris quae hodie praecipio tibi ut diligas Dominum Deum tuum et ambules in viis eius omni tempore addes tibi tres alias civitates et supradictarum trium urbium numerum duplicabis
DEUT|19|10|ut non effundatur sanguis innoxius in medio terrae quam Dominus Deus tuus dabit tibi possidendam nec sis sanguinis reus
DEUT|19|11|si quis autem odio habens proximum suum insidiatus fuerit vitae eius surgensque percusserit illum et mortuus fuerit fugeritque ad unam de supradictis urbibus
DEUT|19|12|mittent seniores civitatis illius et arripient eum de loco effugii tradentque in manu proximi cuius sanguis effusus est et morietur
DEUT|19|13|nec misereberis eius et auferes innoxium sanguinem de Israhel ut bene sit tibi
DEUT|19|14|non adsumes et transferes terminos proximi tui quos fixerunt priores in possessione tua quam Dominus Deus tuus dabit tibi in terra quam acceperis possidendam
DEUT|19|15|non stabit testis unus contra aliquem quicquid illud peccati et facinoris fuerit sed in ore duorum aut trium testium stabit omne verbum
DEUT|19|16|si steterit testis mendax contra hominem accusans eum praevaricationis
DEUT|19|17|stabunt ambo quorum causa est ante Dominum in conspectu sacerdotum et iudicum qui fuerint in diebus illis
DEUT|19|18|cumque diligentissime perscrutantes invenerint falsum testem dixisse contra fratrem suum mendacium
DEUT|19|19|reddent ei sicut fratri suo facere cogitavit et auferes malum de medio tui
DEUT|19|20|ut audientes ceteri timorem habeant et nequaquam talia audeant facere
DEUT|19|21|non misereberis eius sed animam pro anima oculum pro oculo dentem pro dente manum pro manu pedem pro pede exiges
DEUT|20|1|si exieris ad bellum contra hostes tuos et videris equitatum et currus et maiorem quam tu habes adversarii exercitus multitudinem non timebis eos quia Dominus Deus tuus tecum est qui eduxit te de terra Aegypti
DEUT|20|2|adpropinquante autem iam proelio stabit sacerdos ante aciem et sic loquetur ad populum
DEUT|20|3|audi Israhel vos hodie contra inimicos vestros pugnam committitis non pertimescat cor vestrum nolite metuere nolite cedere nec formidetis eos
DEUT|20|4|quia Dominus Deus vester in medio vestri est et pro vobis contra adversarios dimicabit ut eruat vos de periculo
DEUT|20|5|duces quoque per singulas turmas audiente exercitu proclamabunt quis est homo qui aedificavit domum novam et non dedicavit eam vadat et revertatur in domum suam ne forte moriatur in bello et alius dedicet illam
DEUT|20|6|quis est homo qui plantavit vineam et necdum eam fecit esse communem et de qua vesci omnibus liceat vadat et revertatur in domum suam ne forte moriatur in bello et alius homo eius fungatur officio
DEUT|20|7|quis est homo qui despondit uxorem et non accepit eam vadat et revertatur in domum suam ne forte moriatur in bello et alius homo accipiat eam
DEUT|20|8|his dictis addent reliqua et loquentur ad populum quis est homo formidolosus et corde pavido vadat et revertatur in domum suam ne pavere faciat corda fratrum suorum sicut ipse timore perterritus est
DEUT|20|9|cumque siluerint exercitus duces et finem loquendi fecerint unusquisque suos ad bellandum cuneos praeparabit
DEUT|20|10|si quando accesseris ad expugnandam civitatem offeres ei primum pacem
DEUT|20|11|si receperit et aperuerit tibi portas cunctus populus qui in ea est salvabitur et serviet tibi sub tributo
DEUT|20|12|sin autem foedus inire noluerint et receperint contra te bellum obpugnabis eam
DEUT|20|13|cumque tradiderit Dominus Deus tuus illam in manu tua percuties omne quod in ea generis masculini est in ore gladii
DEUT|20|14|absque mulieribus et infantibus iumentis et ceteris quae in civitate sunt omnem praedam exercitui divides et comedes de spoliis hostium tuorum quae Dominus Deus tuus dederit tibi
DEUT|20|15|sic facies cunctis civitatibus quae a te procul valde sunt et non sunt de his urbibus quas in possessionem accepturus es
DEUT|20|16|de his autem civitatibus quae dabuntur tibi nullum omnino permittes vivere
DEUT|20|17|sed interficies in ore gladii Hettheum videlicet et Amorreum et Chananeum Ferezeum et Eveum et Iebuseum sicut praecepit tibi Dominus Deus tuus
DEUT|20|18|ne forte doceant vos facere cunctas abominationes quas ipsi operati sunt diis suis et peccetis in Dominum Deum vestrum
DEUT|20|19|quando obsederis civitatem multo tempore et munitionibus circumdederis ut expugnes eam non succides arbores de quibus vesci potest nec securibus per circuitum debes vastare regionem quoniam lignum est et non homo nec potest bellantium contra te augere numerum
DEUT|20|20|si qua autem ligna non sunt pomifera sed agrestia et in ceteros apta usus succide et extrue machinas donec capias civitatem quae contra te dimicat
DEUT|21|1|quando inventum fuerit in terra quam Dominus Deus tuus daturus est tibi hominis cadaver occisi et ignoratur caedis reus
DEUT|21|2|egredientur maiores natu et iudices tui et metientur a loco cadaveris singularum per circuitum spatia civitatum
DEUT|21|3|et quam viciniorem ceteris esse perspexerint seniores civitatis eius tollent vitulam de armento quae non traxit iugum nec terram scidit vomere
DEUT|21|4|et ducent eam ad vallem asperam atque saxosam quae numquam arata est nec sementem recepit et caedent in ea cervices vitulae
DEUT|21|5|accedentque sacerdotes filii Levi quos elegerit Dominus Deus tuus ut ministrent ei et benedicant in nomine eius et ad verbum eorum omne negotium et quicquid mundum vel inmundum est iudicetur
DEUT|21|6|et maiores natu civitatis illius ad interfectum lavabuntque manus suas super vitulam quae in valle percussa est
DEUT|21|7|et dicent manus nostrae non effuderunt hunc sanguinem nec oculi viderunt
DEUT|21|8|propitius esto populo tuo Israhel quem redemisti Domine et non reputes sanguinem innocentem in medio populi tui Israhel et auferetur ab eis reatus sanguinis
DEUT|21|9|tu autem alienus eris ab innocentis cruore qui fusus est cum feceris quod praecepit Dominus
DEUT|21|10|si egressus fueris ad pugnam contra inimicos tuos et tradiderit eos Dominus Deus tuus in manu tua captivosque duxeris
DEUT|21|11|et videris in numero captivorum mulierem pulchram et adamaveris eam voluerisque habere uxorem
DEUT|21|12|introduces in domum tuam quae radet caesariem et circumcidet ungues
DEUT|21|13|et deponet vestem in qua capta est sedensque in domo tua flebit patrem et matrem suam uno mense et postea intrabis ad eam dormiesque cum illa et erit uxor tua
DEUT|21|14|sin autem postea non sederit animo tuo dimittes eam liberam nec vendere poteris pecunia nec opprimere per potentiam quia humiliasti eam
DEUT|21|15|si habuerit homo uxores duas unam dilectam et alteram odiosam genuerintque ex eo liberos et fuerit filius odiosae primogenitus
DEUT|21|16|volueritque substantiam inter filios suos dividere non poterit filium dilectae facere primogenitum et praeferre filio odiosae
DEUT|21|17|sed filium odiosae agnoscet primogenitum dabitque ei de his quae habuerit cuncta duplicia iste est enim principium liberorum eius et huic debentur primogenita
DEUT|21|18|si genuerit homo filium contumacem et protervum qui non audiat patris aut matris imperium et coercitus oboedire contempserit
DEUT|21|19|adprehendent eum et ducent ad seniores civitatis illius et ad portam iudicii
DEUT|21|20|dicentque ad eos filius noster iste protervus et contumax est monita nostra audire contemnit comesationibus vacat et luxuriae atque conviviis
DEUT|21|21|lapidibus eum obruet populus civitatis et morietur ut auferatis malum de medio vestri et universus Israhel audiens pertimescat
DEUT|21|22|quando peccaverit homo quod morte plectendum est et adiudicatus morti adpensus fuerit in patibulo
DEUT|21|23|non permanebit cadaver eius in ligno sed in eadem die sepelietur quia maledictus a Deo est qui pendet in ligno et nequaquam contaminabis terram tuam quam Dominus Deus tuus dederit tibi in possessionem
DEUT|22|1|non videbis bovem fratris tui aut ovem errantem et praeteribis sed reduces fratri tuo
DEUT|22|2|etiam si non est propinquus tuus frater nec nosti eum duces in domum tuam et erunt apud te quamdiu quaerat ea frater tuus et recipiat
DEUT|22|3|similiter facies de asino et de vestimento et de omni re fratris tui quae perierit si inveneris eam ne neglegas quasi alienam
DEUT|22|4|si videris asinum fratris tui aut bovem cecidisse in via non despicies sed sublevabis cum eo
DEUT|22|5|non induetur mulier veste virili nec vir utetur veste feminea abominabilis enim apud Deum est qui facit haec
DEUT|22|6|si ambulans per viam in arbore vel in terra nidum avis inveneris et matrem pullis vel ovis desuper incubantem non tenebis eam cum filiis
DEUT|22|7|sed abire patieris captos tenens filios ut bene sit tibi et longo vivas tempore
DEUT|22|8|cum aedificaveris domum novam facies murum tecti per circuitum ne effundatur sanguis in domo tua et sis reus labente alio et in praeceps ruente
DEUT|22|9|non seres vineam tuam altero semine ne et sementis quam sevisti et quae nascuntur ex vinea pariter sanctificentur
DEUT|22|10|non arabis in bove simul et asino
DEUT|22|11|non indueris vestimento quod ex lana linoque contextum est
DEUT|22|12|funiculos in fimbriis facies per quattuor angulos pallii tui quo operieris
DEUT|22|13|si duxerit vir uxorem et postea eam odio habuerit
DEUT|22|14|quaesieritque occasiones quibus dimittat eam obiciens ei nomen pessimum et dixerit uxorem hanc accepi et ingressus ad eam non inveni virginem
DEUT|22|15|tollent eam pater et mater eius et ferent secum signa virginitatis eius ad seniores urbis qui in porta sunt
DEUT|22|16|et dicet pater filiam meam dedi huic uxorem quam quia odit
DEUT|22|17|inponet ei nomen pessimum ut dicat non inveni filiam tuam virginem et ecce haec sunt signa virginitatis filiae meae expandent vestimentum coram senibus civitatis
DEUT|22|18|adprehendentque senes urbis illius virum et verberabunt illum
DEUT|22|19|condemnantes insuper centum siclis argenti quos dabit patri puellae quoniam diffamavit nomen pessimum super virginem Israhel habebitque eam uxorem et non poterit dimittere omni tempore vitae suae
DEUT|22|20|quod si verum est quod obicit et non est in puella inventa virginitas
DEUT|22|21|eicient eam extra fores domus patris sui et lapidibus obruent viri civitatis eius et morietur quoniam fecit nefas in Israhel ut fornicaretur in domo patris sui et auferes malum de medio tui
DEUT|22|22|si dormierit vir cum uxore alterius uterque morientur id est adulter et adultera et auferes malum de Israhel
DEUT|22|23|si puellam virginem desponderit vir et invenerit eam aliquis in civitate et concubuerit cum illa
DEUT|22|24|educes utrumque ad portam civitatis illius et lapidibus obruentur puella quia non clamavit cum esset in civitate vir quia humiliavit uxorem proximi sui et auferes malum de medio tui
DEUT|22|25|sin autem in agro reppererit vir puellam quae desponsata est et adprehendens concubuerit cum illa ipse morietur solus
DEUT|22|26|puella nihil patietur nec est rea mortis quoniam sicut latro consurgit contra fratrem suum et occidit animam eius ita et puella perpessa est
DEUT|22|27|sola erat in agro clamavit et nullus adfuit qui liberaret eam
DEUT|22|28|si invenerit vir puellam virginem quae non habet sponsum et adprehendens concubuerit cum ea et res ad iudicium venerit
DEUT|22|29|dabit qui dormivit cum ea patri puellae quinquaginta siclos argenti et habebit eam uxorem quia humiliavit illam non poterit dimittere cunctis diebus vitae suae
DEUT|22|30|non accipiet homo uxorem patris sui nec revelabit operimentum eius
DEUT|23|1|non intrabit eunuchus adtritis vel amputatis testiculis et absciso veretro ecclesiam Domini
DEUT|23|2|non ingredietur mamzer hoc est de scorto natus in ecclesiam Domini usque ad decimam generationem
DEUT|23|3|Ammanites et Moabites etiam post decimam generationem non intrabunt ecclesiam Domini in aeternum
DEUT|23|4|quia noluerunt vobis occurrere cum pane et aqua in via quando egressi estis de Aegypto et quia conduxerunt contra te Balaam filium Beor de Mesopotamiam Syriae ut malediceret tibi
DEUT|23|5|et noluit Dominus Deus tuus audire Balaam vertitque maledictionem eius in benedictionem tuam eo quod diligeret te
DEUT|23|6|non facies cum eis pacem nec quaeres eis bona cunctis diebus vitae tuae in sempiternum
DEUT|23|7|non abominaberis Idumeum quia frater tuus est nec Aegyptium quia advena fuisti in terra eius
DEUT|23|8|qui nati fuerint ex eis tertia generatione intrabunt ecclesiam Domini
DEUT|23|9|quando egressus fueris adversus hostes tuos in pugnam custodies te ab omni re mala
DEUT|23|10|si fuerit inter vos homo qui nocturno pollutus sit somnio egredietur extra castra
DEUT|23|11|et non revertetur priusquam ad vesperam lavetur aqua et post solis occasum regredietur in castra
DEUT|23|12|habebis locum extra castra ad quem egrediaris ad requisita naturae
DEUT|23|13|gerens paxillum in balteo cumque sederis fodies per circuitum et egesta humo operies
DEUT|23|14|quo relevatus es Dominus enim Deus tuus ambulat in medio castrorum ut eruat te et tradat tibi inimicos tuos ut sint castra tua sancta et nihil in eis appareat foeditatis nec derelinquat te
DEUT|23|15|non trades servum domino suo qui ad te confugerit
DEUT|23|16|habitabit tecum in loco qui ei placuerit et in una urbium tuarum requiescet nec contristes eum
DEUT|23|17|non erit meretrix de filiabus Israhel neque scortator de filiis Israhel
DEUT|23|18|non offeres mercedem prostibuli nec pretium canis in domum Domini Dei tui quicquid illud est quod voverint quia abominatio est utrumque apud Dominum Deum tuum
DEUT|23|19|non fenerabis fratri tuo ad usuram pecuniam nec fruges nec quamlibet aliam rem
DEUT|23|20|sed alieno fratri autem tuo absque usura id quod indiget commodabis ut benedicat tibi Dominus Deus tuus in omni opere tuo in terra ad quam ingredieris possidendam
DEUT|23|21|cum voveris votum Domino Deo tuo non tardabis reddere quia requiret illud Dominus Deus tuus et si moratus fueris reputabit tibi in peccatum
DEUT|23|22|si nolueris polliceri absque peccato eris
DEUT|23|23|quod autem semel egressum est de labiis tuis observabis et facies sicut promisisti Domino Deo tuo et propria voluntate et ore tuo locutus es
DEUT|23|24|ingressus vineam proximi tui comede uvas quantum tibi placuerit foras autem ne efferas tecum
DEUT|23|25|si intraveris in segetem amici tui franges spicas et manu conteres falce autem non metes
DEUT|24|1|si acceperit homo uxorem et habuerit eam et non invenerit gratiam ante oculos eius propter aliquam foeditatem scribet libellum repudii et dabit in manu illius et dimittet eam de domo sua
DEUT|24|2|cumque egressa alterum maritum duxerit
DEUT|24|3|et ille quoque oderit eam dederitque ei libellum repudii et dimiserit de domo sua vel certe mortuus fuerit
DEUT|24|4|non poterit prior maritus recipere eam in uxorem quia polluta est et abominabilis facta est coram Domino ne peccare facias terram tuam quam Dominus Deus tuus tibi tradiderit possidendam
DEUT|24|5|cum acceperit homo nuper uxorem non procedet ad bellum nec ei quippiam necessitatis iniungetur publicae sed vacabit absque culpa domui suae ut uno anno laetetur cum uxore sua
DEUT|24|6|non accipies loco pignoris inferiorem et superiorem molam quia animam suam adposuit tibi
DEUT|24|7|si deprehensus fuerit homo sollicitans fratrem suum de filiis Israhel et vendito eo accipiens pretium interficietur et auferes malum de medio tui
DEUT|24|8|observa diligenter ne incurras in plagam leprae sed facies quaecumque docuerint te sacerdotes levitici generis iuxta id quod praecepi eis et imple sollicite
DEUT|24|9|mementote quae fecerit Dominus Deus vester Mariae in via cum egrederemini de Aegypto
DEUT|24|10|cum repetes a proximo tuo rem aliquam quam debet tibi non ingredieris domum eius ut pignus auferas
DEUT|24|11|sed stabis foris et ille tibi proferet quod habuerit
DEUT|24|12|sin autem pauper est non pernoctabit apud te pignus
DEUT|24|13|sed statim reddes ei ante solis occasum ut dormiens in vestimento suo benedicat tibi et habeas iustitiam coram Domino Deo tuo
DEUT|24|14|non negabis mercedem indigentis et pauperis fratris tui sive advenae qui tecum moratur in terra et intra portas tuas est
DEUT|24|15|sed eadem die reddes ei pretium laboris sui ante solis occasum quia pauper est et ex eo sustentat animam suam ne clamet contra te ad Dominum et reputetur tibi in peccatum
DEUT|24|16|non occidentur patres pro filiis nec filii pro patribus sed unusquisque pro suo peccato morietur
DEUT|24|17|non pervertes iudicium advenae et pupilli nec auferes pignoris loco viduae vestimentum
DEUT|24|18|memento quod servieris in Aegypto et eruerit te Dominus Deus tuus inde idcirco praecipio tibi ut facias hanc rem
DEUT|24|19|quando messueris segetem in agro tuo et oblitus manipulum reliqueris non reverteris ut tollas eum sed advenam et pupillum et viduam auferre patieris ut benedicat tibi Dominus Deus tuus in omni opere manuum tuarum
DEUT|24|20|si fruges colliges olivarum quicquid remanserit in arboribus non reverteris ut colligas sed relinques advenae pupillo ac viduae
DEUT|24|21|si vindemiaveris vineam tuam non colliges remanentes racemos sed cedent in usus advenae pupilli ac viduae
DEUT|24|22|memento quod et tu servieris in Aegypto et idcirco praecipiam tibi ut facias hanc rem
DEUT|25|1|si fuerit causa inter aliquos et interpellaverint iudices quem iustum esse perspexerint illi iustitiae palmam dabunt quem impium condemnabunt impietatis
DEUT|25|2|sin autem eum qui peccavit dignum viderint plagis prosternent et coram se facient verberari pro mensura peccati erit et plagarum modus
DEUT|25|3|ita dumtaxat ut quadragenarium numerum non excedant ne foede laceratus ante oculos tuos abeat frater tuus
DEUT|25|4|non ligabis os bovis terentis in area fruges tuas
DEUT|25|5|quando habitaverint fratres simul et unus ex eis absque liberis mortuus fuerit uxor defuncti non nubet alteri sed accipiet eam frater eius et suscitabit semen fratris sui
DEUT|25|6|et primogenitum ex ea filium nomine illius appellabit ut non deleatur nomen eius ex Israhel
DEUT|25|7|sin autem noluerit accipere uxorem fratris sui quae ei lege debetur perget mulier ad portam civitatis et interpellabit maiores natu dicetque non vult frater viri mei suscitare nomen fratris sui in Israhel nec me in coniugium sumere
DEUT|25|8|statimque accersiri eum facient et interrogabunt si responderit nolo eam uxorem accipere
DEUT|25|9|accedet mulier ad eum coram senioribus et tollet calciamentum de pede eius spuetque in faciem illius et dicet sic fit homini qui non aedificat domum fratris sui
DEUT|25|10|et vocabitur nomen illius in Israhel domus Disculciati
DEUT|25|11|si habuerint inter se iurgium viri et unus contra alterum rixari coeperit volensque uxor alterius eruere virum suum de manu fortioris miserit manum et adprehenderit verenda eius
DEUT|25|12|abscides manum illius nec flecteris super eam ulla misericordia
DEUT|25|13|non habebis in sacculo diversa pondera maius et minus
DEUT|25|14|nec erit in domo tua modius maior et minor
DEUT|25|15|pondus habebis iustum et verum et modius aequalis et verus erit tibi ut multo vivas tempore super terram quam Dominus Deus tuus dederit tibi
DEUT|25|16|abominatur enim Dominus eum qui facit haec et aversatur omnem iniustitiam
DEUT|25|17|memento quae fecerit tibi Amalech in via quando egrediebaris ex Aegypto
DEUT|25|18|quomodo occurrerit tibi et extremos agminis tui qui lassi residebant ceciderit quando tu eras fame et labore confectus et non timuerit Deum
DEUT|25|19|cum ergo Dominus Deus tuus dederit tibi requiem et subiecerit cunctas per circuitum nationes in terra quam tibi pollicitus est delebis nomen eius sub caelo cave ne obliviscaris
DEUT|26|1|cumque intraveris terram quam Dominus Deus tuus tibi daturus est possidendam et obtinueris eam atque habitaveris in illa
DEUT|26|2|tolles de cunctis frugibus primitias et pones in cartallo pergesque ad locum quem Dominus Deus tuus elegerit ut ibi invocetur nomen eius
DEUT|26|3|accedesque ad sacerdotem qui fuerit in diebus illis et dices ad eum profiteor hodie coram Domino Deo tuo quod ingressus sim terram pro qua iuravit patribus nostris ut daret eam nobis
DEUT|26|4|suscipiensque sacerdos cartallum de manu eius ponet ante altare Domini Dei tui
DEUT|26|5|et loqueris in conspectu Domini Dei tui Syrus persequebatur patrem meum qui descendit in Aegyptum et ibi peregrinatus est in paucissimo numero crevitque in gentem magnam et robustam et infinitae multitudinis
DEUT|26|6|adflixeruntque nos Aegyptii et persecuti sunt inponentes onera gravissima
DEUT|26|7|et clamavimus ad Dominum Deum patrum nostrorum qui exaudivit nos et respexit humilitatem nostram et laborem atque angustias
DEUT|26|8|et eduxit nos de Aegypto in manu forti et brachio extento in ingenti pavore in signis atque portentis
DEUT|26|9|et introduxit ad locum istum et tradidit nobis terram lacte et melle manantem
DEUT|26|10|et idcirco nunc offero primitias frugum terrae quam dedit Dominus mihi et dimittes eas in conspectu Domini Dei tui adorato Domino Deo tuo
DEUT|26|11|et epulaberis in omnibus bonis quae Dominus Deus tuus dederit tibi et domui tuae tu et Levites et advena qui tecum est
DEUT|26|12|quando conpleveris decimam cunctarum frugum tuarum anno decimarum tertio dabis Levitae et advenae et pupillo et viduae ut comedant intra portas tuas et saturentur
DEUT|26|13|loquerisque in conspectu Domini Dei tui abstuli quod sanctificatum est de domo mea et dedi illud Levitae et advenae pupillo et viduae sicut iussisti mihi non praeterivi mandata tua nec sum oblitus imperii
DEUT|26|14|non comedi ex eis in luctu meo nec separavi ea in qualibet inmunditia nec expendi ex his quicquam in re funebri oboedivi voci Domini Dei mei et feci omnia sicut praecepisti mihi
DEUT|26|15|respice de sanctuario tuo de excelso caelorum habitaculo et benedic populo tuo Israhel et terrae quam dedisti nobis sicut iurasti patribus nostris terrae lacte et melle mananti
DEUT|26|16|hodie Dominus Deus tuus praecepit tibi ut facias mandata haec atque iudicia et custodias et impleas ex toto corde tuo et ex tota anima tua
DEUT|26|17|Dominum elegisti hodie ut sit tibi Deus et ambules in viis eius et custodias caerimonias illius et mandata atque iudicia et oboedias eius imperio
DEUT|26|18|et Dominus elegit te hodie ut sis ei populus peculiaris sicut locutus est tibi et custodias omnia praecepta eius
DEUT|26|19|et faciat te excelsiorem cunctis gentibus quas creavit in laudem et nomen et gloriam suam ut sis populus sanctus Domini Dei tui sicut locutus est
DEUT|27|1|praecepit autem Moses et seniores Israhel populo dicentes custodite omne mandatum quod praecipio vobis hodie
DEUT|27|2|cumque transieritis Iordanem in terram quam Dominus Deus tuus dabit tibi eriges ingentes lapides et calce levigabis eos
DEUT|27|3|ut possis in eis scribere omnia verba legis huius Iordane transmisso ut introeas terram quam Dominus Deus tuus dabit tibi terram lacte et melle manantem sicut iuravit patribus tuis
DEUT|27|4|quando ergo transieritis Iordanem erige lapides quos ego hodie praecipio vobis in monte Hebal et levigabis calce
DEUT|27|5|et aedificabis ibi altare Domino Deo tuo de lapidibus quos ferrum non tetigit
DEUT|27|6|et de saxis informibus et inpolitis et offeres super eo holocausta Domino Deo tuo
DEUT|27|7|et immolabis hostias pacificas comedesque ibi et epulaberis coram Domino Deo tuo
DEUT|27|8|et scribes super lapides omnia verba legis huius plane et lucide
DEUT|27|9|dixeruntque Moses et sacerdotes levitici generis ad omnem Israhelem adtende et audi Israhel hodie factus es populus Domini Dei tui
DEUT|27|10|audies vocem eius et facies mandata atque iustitias quas ego praecipio tibi
DEUT|27|11|praecepitque Moses populo in die illo dicens
DEUT|27|12|hii stabunt ad benedicendum Domino super montem Garizim Iordane transmisso Symeon Levi Iudas Isachar Ioseph et Beniamin
DEUT|27|13|et e regione isti stabunt ad maledicendum in monte Hebal Ruben Gad et Aser Zabulon Dan et Nepthalim
DEUT|27|14|et pronuntiabunt Levitae dicentque ad omnes viros Israhel excelsa voce
DEUT|27|15|maledictus homo qui facit sculptile et conflatile abominationem Domini opus manuum artificum ponetque illud in abscondito et respondebit omnis populus et dicet amen
DEUT|27|16|maledictus qui non honorat patrem suum et matrem et dicet omnis populus amen
DEUT|27|17|maledictus qui transfert terminos proximi sui et dicet omnis populus amen
DEUT|27|18|maledictus qui errare facit caecum in itinere et dicet omnis populus amen
DEUT|27|19|maledictus qui pervertit iudicium advenae pupilli et viduae et dicet omnis populus amen
DEUT|27|20|maledictus qui dormit cum uxore patris sui et revelat operimentum lectuli eius et dicet omnis populus amen
DEUT|27|21|maledictus qui dormit cum omni iumento et dicet omnis populus amen
DEUT|27|22|maledictus qui dormit cum sorore sua filia patris sui sive matris suae et dicet omnis populus amen
DEUT|27|23|maledictus qui dormit cum socru sua et dicet omnis populus amen
DEUT|27|24|maledictus qui clam percusserit proximum suum et dicet omnis populus amen
DEUT|27|25|maledictus qui accipit munera ut percutiat animam sanguinis innocentis et dicet omnis populus amen
DEUT|27|26|maledictus qui non permanet in sermonibus legis huius nec eos opere perficit et dicet omnis populus amen
DEUT|28|1|sin autem audieris vocem Domini Dei tui ut facias atque custodias omnia mandata eius quae ego praecipio tibi hodie faciet te Dominus Deus tuus excelsiorem cunctis gentibus quae versantur in terra
DEUT|28|2|venientque super te universae benedictiones istae et adprehendent te si tamen praecepta eius audieris
DEUT|28|3|benedictus tu in civitate et benedictus in agro
DEUT|28|4|benedictus fructus ventris tui et fructus terrae tuae fructusque iumentorum tuorum greges armentorum et caulae ovium tuarum
DEUT|28|5|benedicta horrea tua et benedictae reliquiae tuae
DEUT|28|6|benedictus eris et ingrediens et egrediens
DEUT|28|7|dabit Dominus inimicos tuos qui consurgunt adversum te corruentes in conspectu tuo per unam viam venient contra te et per septem fugient a facie tua
DEUT|28|8|emittet Dominus benedictionem super cellaria tua et super omnia opera manuum tuarum benedicetque tibi in terra quam acceperis
DEUT|28|9|suscitabit te Dominus sibi in populum sanctum sicut iuravit tibi si custodieris mandata Domini Dei tui et ambulaveris in viis eius
DEUT|28|10|videbuntque omnes terrarum populi quod nomen Domini invocatum sit super te et timebunt te
DEUT|28|11|abundare te faciet Dominus omnibus bonis fructu uteri tui et fructu iumentorum tuorum fructu terrae tuae quam iuravit Dominus patribus tuis ut daret tibi
DEUT|28|12|aperiet Dominus thesaurum suum optimum caelum ut tribuat pluviam terrae tuae in tempore suo benedicet cunctis operibus manuum tuarum et fenerabis gentibus multis et ipse a nullo fenus accipies
DEUT|28|13|constituet te Dominus in caput et non in caudam et eris semper supra et non subter si audieris mandata Domini Dei tui quae ego praecipio tibi hodie et custodieris et feceris
DEUT|28|14|ac non declinaveris ab eis nec ad dextram nec ad sinistram nec secutus fueris deos alienos neque colueris eos
DEUT|28|15|quod si audire nolueris vocem Domini Dei tui ut custodias et facias omnia mandata eius et caerimonias quas ego praecipio tibi hodie venient super te omnes maledictiones istae et adprehendent te
DEUT|28|16|maledictus eris in civitate maledictus in agro
DEUT|28|17|maledictum horreum tuum et maledictae reliquiae tuae
DEUT|28|18|maledictus fructus ventris tui et fructus terrae tuae armenta boum tuorum et greges ovium tuarum
DEUT|28|19|maledictus eris ingrediens et maledictus egrediens
DEUT|28|20|mittet Dominus super te famem et esuriem et increpationem in omnia opera tua quae facies donec conterat te et perdat velociter propter adinventiones tuas pessimas in quibus reliquisti me
DEUT|28|21|adiungat Dominus tibi pestilentiam donec consumat te de terra ad quam ingredieris possidendam
DEUT|28|22|percutiat te Dominus egestate febri et frigore ardore et aestu et aere corrupto ac robigine et persequatur donec pereas
DEUT|28|23|sit caelum quod supra te est aeneum et terra quam calcas ferrea
DEUT|28|24|det Dominus imbrem terrae tuae pulverem et de caelo descendat super te cinis donec conteraris
DEUT|28|25|tradat te Dominus corruentem ante hostes tuos per unam viam egrediaris contra eos et per septem fugias et dispergaris per omnia regna terrae
DEUT|28|26|sitque cadaver tuum in escam cunctis volatilibus caeli et bestiis terrae et non sit qui abigat
DEUT|28|27|percutiat te Dominus ulcere Aegypti et parte corporis per quam stercora digeruntur scabie quoque et prurigine ita ut curari nequeas
DEUT|28|28|percutiat te Dominus amentia et caecitate ac furore mentis
DEUT|28|29|et palpes in meridie sicut palpare solet caecus in tenebris et non dirigas vias tuas omnique tempore calumniam sustineas et opprimaris violentia nec habeas qui liberet te
DEUT|28|30|uxorem accipias et alius dormiat cum ea domum aedifices et non habites in ea plantes vineam et non vindemies eam
DEUT|28|31|bos tuus immoletur coram te et non comedas ex eo asinus tuus rapiatur in conspectu tuo et non reddatur tibi oves tuae dentur inimicis tuis et non sit qui te adiuvet
DEUT|28|32|filii tui et filiae tuae tradantur alteri populo videntibus oculis tuis et deficientibus ad conspectum eorum tota die et non sit fortitudo in manu tua
DEUT|28|33|fructus terrae tuae et omnes labores tuos comedat populus quem ignoras et sis semper calumniam sustinens et oppressus cunctis diebus
DEUT|28|34|et stupens ad terrorem eorum quae videbunt oculi tui
DEUT|28|35|percutiat te Dominus ulcere pessimo in genibus et in suris sanarique non possis a planta pedis usque ad verticem tuum
DEUT|28|36|ducet Dominus te et regem tuum quem constitueris super te in gentem quam ignoras tu et patres tui et servies ibi diis alienis ligno et lapidi
DEUT|28|37|et eris perditus in proverbium ac fabulam omnibus populis ad quos te introduxerit Dominus
DEUT|28|38|sementem multam iacies in terram et modicum congregabis quia lucustae omnia devorabunt
DEUT|28|39|vineam plantabis et fodies et vinum non bibes nec colliges ex ea quippiam quoniam vastabitur vermibus
DEUT|28|40|olivas habebis in omnibus terminis tuis et non ungueris oleo quia defluent et peribunt
DEUT|28|41|filios generabis et filias et non frueris eis quoniam ducentur in captivitatem
DEUT|28|42|omnes arbores tuas et fruges terrae tuae robigo consumet
DEUT|28|43|advena qui tecum versatur in terra ascendet super te eritque sublimior tu autem descendes et eris inferior
DEUT|28|44|ipse fenerabit tibi et tu non fenerabis ei ipse erit in caput et tu eris in caudam
DEUT|28|45|et venient super te omnes maledictiones istae et persequentes adprehendent te donec intereas quia non audisti vocem Domini Dei tui nec servasti mandata eius et caerimonias quas praecepit tibi
DEUT|28|46|et erunt in te signa atque prodigia et in semine tuo usque in sempiternum
DEUT|28|47|eo quod non servieris Domino Deo tuo in gaudio cordisque laetitia propter rerum omnium abundantiam
DEUT|28|48|servies inimico tuo quem inmittet Dominus tibi in fame et siti et nuditate et omnium penuria et ponet iugum ferreum super cervicem tuam donec te conterat
DEUT|28|49|adducet Dominus super te gentem de longinquo et de extremis finibus terrae in similitudinem aquilae volantis cum impetu cuius linguam intellegere non possis
DEUT|28|50|gentem procacissimam quae non deferat seni nec misereatur parvulo
DEUT|28|51|et devoret fructum iumentorum tuorum ac fruges terrae tuae donec intereas et non relinquat tibi triticum vinum et oleum armenta boum et greges ovium donec te disperdat
DEUT|28|52|et conterat in cunctis urbibus tuis et destruantur muri tui firmi atque sublimes in quibus habebas fiduciam in omni terra tua obsideberis intra portas tuas in omni terra quam dabit tibi Dominus Deus tuus
DEUT|28|53|et comedes fructum uteri tui et carnes filiorum et filiarum tuarum quas dedit tibi Dominus Deus tuus in angustia et vastitate qua opprimet te hostis tuus
DEUT|28|54|homo delicatus in te et luxuriosus valde invidebit fratri suo et uxori quae cubat in sinu suo
DEUT|28|55|ne det eis de carnibus filiorum suorum quas comedet eo quod nihil habeat aliud in obsidione et penuria qua vastaverint te inimici tui intra omnes portas tuas
DEUT|28|56|tenera mulier et delicata quae super terram ingredi non valebat nec pedis vestigium figere propter mollitiem et teneritudinem nimiam invidebit viro suo qui cubat in sinu eius super filii et filiae carnibus
DEUT|28|57|et inluvie secundarum quae egrediuntur de medio feminum eius et super liberis qui eadem hora nati sunt comedent enim eos clam propter rerum omnium penuriam in obsidione et vastitate qua opprimet te inimicus tuus intra portas tuas
DEUT|28|58|nisi custodieris et feceris omnia verba legis huius quae scripta sunt in hoc volumine et timueris nomen eius gloriosum et terribile hoc est Dominum Deum tuum
DEUT|28|59|augebit Dominus plagas tuas et plagas seminis tui plagas magnas et perseverantes infirmitates pessimas et perpetuas
DEUT|28|60|et convertet in te omnes adflictiones Aegypti quas timuisti et adherebunt tibi
DEUT|28|61|insuper et universos languores et plagas quae non sunt scriptae in volumine legis huius inducet Dominus super te donec te conterat
DEUT|28|62|et remanebitis pauci numero qui prius eratis sicut astra caeli prae multitudine quoniam non audisti vocem Domini Dei tui
DEUT|28|63|et sicut ante laetatus est Dominus super vos bene vobis faciens vosque multiplicans sic laetabitur disperdens vos atque subvertens ut auferamini de terra ad quam ingredieris possidendam
DEUT|28|64|disperget te Dominus in omnes populos a summitate terrae usque ad terminos eius et servies ibi diis alienis quos et tu ignoras et patres tui lignis et lapidibus
DEUT|28|65|in gentibus quoque illis non quiesces neque erit requies vestigio pedis tui dabit enim tibi Dominus ibi cor pavidum et deficientes oculos et animam maerore consumptam
DEUT|28|66|et erit vita tua quasi pendens ante te timebis nocte et die et non credes vitae tuae
DEUT|28|67|mane dices quis mihi det vesperum et vespere quis mihi det mane propter cordis tui formidinem qua terreberis et propter ea quae tuis videbis oculis
DEUT|28|68|reducet te Dominus classibus in Aegyptum per viam de qua dixi tibi ut eam amplius non videres ibi venderis inimicis tuis in servos et ancillas et non erit qui emat
DEUT|29|1|haec sunt verba foederis quod praecepit Dominus Mosi ut feriret cum filiis Israhel in terra Moab praeter illud foedus quod cum eis pepigit in Horeb
DEUT|29|2|vocavitque Moses omnem Israhelem et dixit ad eos vos vidistis universa quae fecit Dominus coram vobis in terra Aegypti Pharaoni et omnibus servis eius universaeque terrae illius
DEUT|29|3|temptationes magnas quas viderunt oculi tui signa illa portentaque ingentia
DEUT|29|4|et non dedit Dominus vobis cor intellegens et oculos videntes et aures quae possint audire usque in praesentem diem
DEUT|29|5|adduxi vos quadraginta annis per desertum non sunt adtrita vestimenta vestra nec calciamenta pedum tuorum vetustate consumpta sunt
DEUT|29|6|panem non comedistis vinum et siceram non bibistis ut sciretis quia ego sum Dominus Deus vester
DEUT|29|7|et venistis ad locum hunc egressusque est Seon rex Esebon et Og rex Basan occurrens nobis ad pugnam et percussimus eos
DEUT|29|8|et tulimus terram eorum ac tradidimus possidendam Ruben et Gad et dimidiae tribui Manasse
DEUT|29|9|custodite ergo verba pacti huius et implete ea ut intellegatis universa quae facitis
DEUT|29|10|vos statis hodie cuncti coram Domino Deo vestro principes vestri ac tribus et maiores natu atque doctores omnis populus Israhel
DEUT|29|11|liberi et uxores vestrae et advena qui tecum moratur in castris exceptis lignorum caesoribus et his qui conportant aquas
DEUT|29|12|ut transeas in foedere Domini Dei tui et in iureiurando quod hodie Dominus Deus tuus percutit tecum
DEUT|29|13|ut suscitet te sibi in populum et ipse sit Deus tuus sicut locutus est tibi et sicut iuravit patribus tuis Abraham Isaac et Iacob
DEUT|29|14|nec vobis solis ego hoc foedus ferio et haec iuramenta confirmo
DEUT|29|15|sed cunctis praesentibus et absentibus
DEUT|29|16|vos enim nostis ut habitaverimus in terra Aegypti et quomodo transierimus per medium nationum quas transeuntes
DEUT|29|17|vidistis abominationes et sordes id est idola eorum lignum et lapidem argentum et aurum quae colebant
DEUT|29|18|ne forte sit inter vos vir aut mulier familia aut tribus cuius cor aversum est hodie a Domino Deo vestro ut vadat et serviat diis illarum gentium et sit inter vos radix germinans fel et amaritudinem
DEUT|29|19|cumque audierit verba iuramenti huius benedicat sibi in corde suo dicens pax erit mihi et ambulabo in pravitate cordis mei et adsumat ebria sitientem
DEUT|29|20|et Dominus non ignoscat ei sed tunc quam maxime furor eius fumet et zelus contra hominem illum et sedeant super eo omnia maledicta quae scripta sunt in hoc volumine et deleat nomen eius sub caelo
DEUT|29|21|et consumat eum in perditionem ex omnibus tribubus Israhel iuxta maledictiones quae in libro legis huius ac foederis continentur
DEUT|29|22|dicetque sequens generatio et filii qui nascentur deinceps et peregrini qui de longe venerint videntes plagas terrae illius et infirmitates quibus eam adflixerit Dominus
DEUT|29|23|sulphure et salis ardore conburens ita ut ultra non seratur nec virens quippiam germinet in exemplum subversionis Sodomae et Gomorrae Adamae et Seboim quas subvertit Dominus in ira et furore suo
DEUT|29|24|et dicent omnes gentes quare sic fecit Dominus terrae huic quae est haec ira furoris eius inmensa
DEUT|29|25|et respondebunt quia dereliquerunt pactum Domini quod pepigit cum patribus eorum quando eduxit eos de terra Aegypti
DEUT|29|26|et servierunt diis alienis et adoraverunt eos quos nesciebant et quibus non fuerant adtributi
DEUT|29|27|idcirco iratus est furor Domini contra terram istam ut induceret super eam omnia maledicta quae in hoc volumine scripta sunt
DEUT|29|28|et eiecit eos de terra sua in ira et furore et indignatione maxima proiecitque in terram alienam sicut hodie conprobatur
DEUT|29|29|abscondita Domino Deo nostro quae manifesta sunt nobis et filiis nostris usque in aeternum ut faciamus universa legis huius
DEUT|30|1|cum ergo venerint super te omnes sermones isti benedictio sive maledictio quam proposui in conspectu tuo et ductus paenitudine cordis tui in universis gentibus in quas disperserit te Dominus Deus tuus
DEUT|30|2|reversus fueris ad eum et oboedieris eius imperiis sicut ego hodie praecipio tibi cum filiis tuis in toto corde tuo et in tota anima tua
DEUT|30|3|reducet Dominus Deus tuus captivitatem tuam ac miserebitur tui et rursum congregabit te de cunctis populis in quos te ante dispersit
DEUT|30|4|si ad cardines caeli fueris dissipatus inde te retrahet Dominus Deus tuus
DEUT|30|5|et adsumet atque introducet in terram quam possederunt patres tui et obtinebis eam et benedicens tibi maioris numeri esse te faciet quam fuerunt patres tui
DEUT|30|6|circumcidet Dominus Deus tuus cor tuum et cor seminis tui ut diligas Dominum Deum tuum in toto corde tuo et in tota anima tua et possis vivere
DEUT|30|7|omnes autem maledictiones has convertet super inimicos tuos et eos qui oderunt te et persequuntur
DEUT|30|8|tu autem reverteris et audies vocem Domini Dei tui faciesque universa mandata quae ego praecipio tibi hodie
DEUT|30|9|et abundare te faciet Dominus Deus tuus in cunctis operibus manuum tuarum in subole uteri tui et in fructu iumentorum tuorum in ubertate terrae tuae et in rerum omnium largitate revertetur enim Dominus ut gaudeat super te in omnibus bonis sicut gavisus est in patribus tuis
DEUT|30|10|si tamen audieris vocem Domini Dei tui et custodieris praecepta eius et caerimonias quae in hac lege conscriptae sunt et revertaris ad Dominum Deum tuum in toto corde tuo et in tota anima tua
DEUT|30|11|mandatum hoc quod ego praecipio tibi hodie non supra te est neque procul positum
DEUT|30|12|nec in caelo situm ut possis dicere quis nostrum ad caelum valet conscendere ut deferat illud ad nos et audiamus atque opere conpleamus
DEUT|30|13|neque trans mare positum ut causeris et dicas quis e nobis transfretare poterit mare et illud ad nos usque deferre ut possimus audire et facere quod praeceptum est
DEUT|30|14|sed iuxta te est sermo valde in ore tuo et in corde tuo ut facias illum
DEUT|30|15|considera quod hodie proposuerim in conspectu tuo vitam et bonum et e contrario mortem et malum
DEUT|30|16|ut diligas Dominum Deum tuum et ambules in viis eius et custodias mandata illius et caerimonias atque iudicia et vivas ac multiplicet te benedicatque tibi in terra ad quam ingredieris possidendam
DEUT|30|17|sin autem aversum fuerit cor tuum et audire nolueris atque errore deceptus adoraveris deos alienos et servieris eis
DEUT|30|18|praedico tibi hodie quod pereas et parvo tempore moreris in terra ad quam Iordane transmisso ingredieris possidendam
DEUT|30|19|testes invoco hodie caelum et terram quod proposuerim vobis vitam et mortem bonum et malum benedictionem et maledictionem elige ergo vitam ut et tu vivas et semen tuum
DEUT|30|20|et diligas Dominum Deum tuum atque oboedias voci eius et illi adhereas ipse est enim vita tua et longitudo dierum tuorum ut habites in terra pro qua iuravit Dominus patribus tuis Abraham Isaac et Iacob ut daret eam illis
DEUT|31|1|abiit itaque Moses et locutus est omnia verba haec ad universum Israhel
DEUT|31|2|et dixit ad eos centum viginti annorum sum hodie non possum ultra egredi et ingredi praesertim cum et Dominus dixerit mihi non transibis Iordanem istum
DEUT|31|3|Dominus ergo Deus tuus transibit ante te ipse delebit omnes gentes has in conspectu tuo et possidebis eas et Iosue iste transibit ante te sicut locutus est Dominus
DEUT|31|4|facietque Dominus eis sicut fecit Seon et Og regibus Amorreorum et terrae eorum delebitque eos
DEUT|31|5|cum ergo et hos tradiderit vobis similiter facietis eis sicut praecepi vobis
DEUT|31|6|viriliter agite et confortamini nolite timere nec paveatis a conspectu eorum quia Dominus Deus tuus ipse est ductor tuus et non dimittet nec derelinquet te
DEUT|31|7|vocavitque Moses Iosue et dixit ei coram omni Israhel confortare et esto robustus tu enim introduces populum istum in terram quam daturum se patribus eorum iuravit Dominus et tu eam sorte divides
DEUT|31|8|et Dominus qui ductor vester est ipse erit tecum non dimittet nec derelinquet te noli timere nec paveas
DEUT|31|9|scripsit itaque Moses legem hanc et tradidit eam sacerdotibus filiis Levi qui portabant arcam foederis Domini et cunctis senioribus Israhelis
DEUT|31|10|praecepitque eis dicens post septem annos anno remissionis in sollemnitate tabernaculorum
DEUT|31|11|convenientibus cunctis ex Israhel ut appareant in conspectu Domini Dei tui in loco quem elegerit Dominus leges verba legis huius coram omni Israhel audientibus eis
DEUT|31|12|et in unum omni populo congregato tam viris quam mulieribus parvulis et advenis qui sunt intra portas tuas ut audientes discant et timeant Dominum Deum vestrum et custodiant impleantque omnes sermones legis huius
DEUT|31|13|filii quoque eorum qui nunc ignorant audire possint et timeant Dominum Deum suum cunctis diebus quibus versantur in terra ad quam vos Iordane transito pergitis obtinendam
DEUT|31|14|et ait Dominus ad Mosen ecce prope sunt dies mortis tuae voca Iosue et state in tabernaculo testimonii ut praecipiam ei abierunt ergo Moses et Iosue et steterunt in tabernaculo testimonii
DEUT|31|15|apparuitque Dominus ibi in columna nubis quae stetit in introitu tabernaculi
DEUT|31|16|dixitque Dominus ad Mosen ecce tu dormies cum patribus tuis et populus iste consurgens fornicabitur post deos alienos in terra ad quam ingredietur et habitabit in ea ibi derelinquet me et irritum faciet foedus quod pepigi cum eo
DEUT|31|17|et irascetur furor meus contra eum in die illo et derelinquam eum et abscondam faciem meam ab eo et erit in devorationem invenient eum omnia mala et adflictiones ita ut dicat in illo die vere quia non est Deus mecum invenerunt me haec mala
DEUT|31|18|ego autem abscondam et celabo faciem meam in die illo propter omnia mala quae fecit quia secutus est deos alienos
DEUT|31|19|nunc itaque scribite vobis canticum istud et docete filios Israhel ut memoriter teneant et ore decantent et sit mihi carmen istud pro testimonio inter filios Israhel
DEUT|31|20|introducam enim eum in terram pro qua iuravi patribus eius lacte et melle manantem cumque comederint et saturati crassique fuerint avertentur ad deos alienos et servient eis et detrahent mihi et irritum facient pactum meum
DEUT|31|21|postquam invenerint eum mala multa et adflictiones respondebit ei canticum istud pro testimonio quod nulla delebit oblivio ex ore seminis tui scio enim cogitationes eius quae facturus sit hodie antequam introducam eum in terram quam ei pollicitus sum
DEUT|31|22|scripsit ergo Moses canticum et docuit filios Israhel
DEUT|31|23|praecepitque Iosue filio Nun et ait confortare et esto robustus tu enim introduces filios Israhel in terram quam pollicitus sum et ego ero tecum
DEUT|31|24|postquam ergo scripsit Moses verba legis huius in volumine atque conplevit
DEUT|31|25|praecepit Levitis qui portabant arcam foederis Domini dicens
DEUT|31|26|tollite librum istum et ponite eum in latere arcae foederis Domini Dei vestri ut sit ibi contra te in testimonio
DEUT|31|27|ego enim scio contentionem tuam et cervicem tuam durissimam adhuc vivente me et ingrediente vobiscum semper contentiose egistis contra Dominum quanto magis cum mortuus fuero
DEUT|31|28|congregate ad me omnes maiores natu per tribus vestras atque doctores et loquar audientibus eis sermones istos et invocabo contra eos caelum et terram
DEUT|31|29|novi enim quod post mortem meam inique agetis et declinabitis cito de via quam praecepi vobis et occurrent vobis mala in extremo tempore quando feceritis malum in conspectu Domini ut inritetis eum per opera manuum vestrarum
DEUT|31|30|locutus est ergo Moses audiente universo coetu Israhel verba carminis huius et ad finem usque conplevit
DEUT|32|1|audite caeli quae loquor audiat terra verba oris mei
DEUT|32|2|concrescat in pluvia doctrina mea fluat ut ros eloquium meum quasi imber super herbam et quasi stillae super gramina
DEUT|32|3|quia nomen Domini invocabo date magnificentiam Deo nostro
DEUT|32|4|Dei perfecta sunt opera et omnes viae eius iudicia Deus fidelis et absque ulla iniquitate iustus et rectus
DEUT|32|5|peccaverunt ei non filii eius in sordibus generatio prava atque perversa
DEUT|32|6|haecine reddis Domino popule stulte et insipiens numquid non ipse est pater tuus qui possedit et fecit et creavit te
DEUT|32|7|memento dierum antiquorum cogita generationes singulas interroga patrem tuum et adnuntiabit tibi maiores tuos et dicent tibi
DEUT|32|8|quando dividebat Altissimus gentes quando separabat filios Adam constituit terminos populorum iuxta numerum filiorum Israhel
DEUT|32|9|pars autem Domini populus eius Iacob funiculus hereditatis eius
DEUT|32|10|invenit eum in terra deserta in loco horroris et vastae solitudinis circumduxit eum et docuit et custodivit quasi pupillam oculi sui
DEUT|32|11|sicut aquila provocans ad volandum pullos suos et super eos volitans expandit alas suas et adsumpsit eum atque portavit in umeris suis
DEUT|32|12|Dominus solus dux eius fuit et non erat cum eo deus alienus
DEUT|32|13|constituit eum super excelsam terram ut comederet fructus agrorum ut sugeret mel de petra oleumque de saxo durissimo
DEUT|32|14|butyrum de armento et lac de ovibus cum adipe agnorum et arietum filiorum Basan et hircos cum medulla tritici et sanguinem uvae biberet meracissimum
DEUT|32|15|incrassatus est dilectus et recalcitravit incrassatus inpinguatus dilatatus dereliquit Deum factorem suum et recessit a Deo salutari suo
DEUT|32|16|provocaverunt eum in diis alienis et in abominationibus ad iracundiam concitaverunt
DEUT|32|17|immolaverunt daemonibus et non Deo diis quos ignorabant novi recentesque venerunt quos non coluerunt patres eorum
DEUT|32|18|Deum qui te genuit dereliquisti et oblitus es Domini creatoris tui
DEUT|32|19|vidit Dominus et ad iracundiam concitatus est quia provocaverunt eum filii sui et filiae
DEUT|32|20|et ait abscondam faciem meam ab eis et considerabo novissima eorum generatio enim perversa est et infideles filii
DEUT|32|21|ipsi me provocaverunt in eo qui non erat Deus et inritaverunt in vanitatibus suis et ego provocabo eos in eo qui non est populus et in gente stulta inritabo illos
DEUT|32|22|ignis succensus est in furore meo et ardebit usque ad inferni novissima devorabitque terram cum germine suo et montium fundamenta conburet
DEUT|32|23|congregabo super eos mala et sagittas meas conplebo in eis
DEUT|32|24|consumentur fame et devorabunt eos aves morsu amarissimo dentes bestiarum inmittam in eos cum furore trahentium super terram atque serpentium
DEUT|32|25|foris vastabit eos gladius et intus pavor iuvenem simul ac virginem lactantem cum homine sene
DEUT|32|26|dixi ubinam sunt cessare faciam ex hominibus memoriam eorum
DEUT|32|27|sed propter iram inimicorum distuli ne forte superbirent hostes eorum et dicerent manus nostra excelsa et non Dominus fecit haec omnia
DEUT|32|28|gens absque consilio est et sine prudentia
DEUT|32|29|utinam saperent et intellegerent ac novissima providerent
DEUT|32|30|quomodo persequatur unus mille et duo fugent decem milia nonne ideo quia Deus suus vendidit eos et Dominus conclusit illos
DEUT|32|31|non enim est Deus noster ut deus eorum et inimici nostri sunt iudices
DEUT|32|32|de vinea Sodomorum vinea eorum et de suburbanis Gomorrae uva eorum uva fellis et botri amarissimi
DEUT|32|33|fel draconum vinum eorum et venenum aspidum insanabile
DEUT|32|34|nonne haec condita sunt apud me et signata in thesauris meis
DEUT|32|35|mea est ultio et ego retribuam in tempore ut labatur pes eorum iuxta est dies perditionis et adesse festinant tempora
DEUT|32|36|iudicabit Dominus populum suum et in servis suis miserebitur videbit quod infirmata sit manus et clausi quoque defecerint residuique consumpti sint
DEUT|32|37|et dicet ubi sunt dii eorum in quibus habebant fiduciam
DEUT|32|38|de quorum victimis comedebant adipes et bibebant vinum libaminum surgant et opitulentur vobis et in necessitate vos protegant
DEUT|32|39|videte quod ego sim solus et non sit alius deus praeter me ego occidam et ego vivere faciam percutiam et ego sanabo et non est qui de manu mea possit eruere
DEUT|32|40|levabo ad caelum manum meam et dicam vivo ego in aeternum
DEUT|32|41|si acuero ut fulgur gladium meum et arripuerit iudicium manus mea reddam ultionem hostibus meis et his qui oderunt me retribuam
DEUT|32|42|inebriabo sagittas meas sanguine et gladius meus devorabit carnes de cruore occisorum et de captivitate nudati inimicorum capitis
DEUT|32|43|laudate gentes populum eius quia sanguinem servorum suorum ulciscetur et vindictam retribuet in hostes eorum et propitius erit terrae populi sui
DEUT|32|44|venit ergo Moses et locutus est omnia verba cantici huius in auribus populi ipse et Iosue filius Nun
DEUT|32|45|conplevitque omnes sermones istos loquens ad universum Israhel
DEUT|32|46|et dixit ad eos ponite corda vestra in omnia verba quae ego testificor vobis hodie ut mandetis ea filiis vestris custodire et facere et implere universa quae scripta sunt legis huius
DEUT|32|47|quia non in cassum praecepta sunt vobis sed ut singuli in eis viverent quae facientes longo perseveretis tempore in terra ad quam Iordane transmisso ingredimini possidendam
DEUT|32|48|locutusque est Dominus ad Mosen in eadem die dicens
DEUT|32|49|ascende in montem istum Abarim id est transituum in montem Nebo qui est in terra Moab contra Hiericho et vide terram Chanaan quam ego tradam filiis Israhel obtinendam et morere in monte
DEUT|32|50|quem conscendens iungeris populis tuis sicut mortuus est Aaron frater tuus in monte Hor et adpositus populis suis
DEUT|32|51|quia praevaricati estis contra me in medio filiorum Israhel ad aquas Contradictionis in Cades deserti Sin et non sanctificastis me inter filios Israhel
DEUT|32|52|e contra videbis terram et non ingredieris in eam quam ego dabo filiis Israhel
DEUT|33|1|haec est benedictio qua benedixit Moses homo Dei filiis Israhel ante mortem suam
DEUT|33|2|et ait Dominus de Sina venit et de Seir ortus est nobis apparuit de monte Pharan et cum eo sanctorum milia in dextera eius ignea lex
DEUT|33|3|dilexit populos omnes sancti in manu illius sunt et qui adpropinquant pedibus eius accipient de doctrina illius
DEUT|33|4|legem praecepit nobis Moses hereditatem multitudinis Iacob
DEUT|33|5|erit apud rectissimum rex congregatis principibus populi cum tribubus Israhel
DEUT|33|6|vivat Ruben et non moriatur et sit parvus in numero
DEUT|33|7|haec est Iudae benedictio audi Domine vocem Iudae et ad populum suum introduc eum manus eius pugnabunt pro eo et adiutor illius contra adversarios eius erit
DEUT|33|8|Levi quoque ait perfectio tua et doctrina tua viro sancto tuo quem probasti in Temptatione et iudicasti ad aquas Contradictionis
DEUT|33|9|qui dixit patri suo et matri suae nescio vos et fratribus suis ignoro illos et nescierunt filios suos hii custodierunt eloquium tuum et pactum tuum servaverunt
DEUT|33|10|iudicia tua o Iacob et legem tuam o Israhel ponent thymiama in furore tuo et holocaustum super altare tuum
DEUT|33|11|benedic Domine fortitudini eius et opera manuum illius suscipe percute dorsa inimicorum eius et qui oderunt eum non consurgant
DEUT|33|12|et Beniamin ait amantissimus Domini habitabit confidenter in eo quasi in thalamo tota die morabitur et inter umeros illius requiescet
DEUT|33|13|Ioseph quoque ait de benedictione Domini terra eius de pomis caeli et rore atque abysso subiacente
DEUT|33|14|de pomis fructuum solis ac lunae
DEUT|33|15|de vertice antiquorum montium de pomis collium aeternorum
DEUT|33|16|et de frugibus terrae et plenitudine eius benedictio illius qui apparuit in rubo veniat super caput Ioseph et super verticem nazarei inter fratres suos
DEUT|33|17|quasi primogeniti tauri pulchritudo eius cornua rinocerotis cornua illius in ipsis ventilabit gentes usque ad terminos terrae hae sunt multitudines Ephraim et haec milia Manasse
DEUT|33|18|et Zabulon ait laetare Zabulon in exitu tuo et Isachar in tabernaculis tuis
DEUT|33|19|populos ad montem vocabunt ibi immolabunt victimas iustitiae qui inundationem maris quasi lac sugent et thesauros absconditos harenarum
DEUT|33|20|et Gad ait benedictus in latitudine Gad quasi leo requievit cepitque brachium et verticem
DEUT|33|21|et vidit principatum suum quod in parte sua doctor esset repositus qui fuit cum principibus populi et fecit iustitias Domini et iudicium suum cum Israhel
DEUT|33|22|Dan quoque ait Dan catulus leonis fluet largiter de Basan
DEUT|33|23|et Nepthalim dixit Nepthalim abundantia perfruetur et plenus erit benedictione Domini mare et meridiem possidebit
DEUT|33|24|Aser quoque ait benedictus in filiis Aser sit placens fratribus suis tinguat in oleo pedem suum
DEUT|33|25|ferrum et aes calciamentum eius sicut dies iuventutis tuae ita et senectus tua
DEUT|33|26|non est alius ut Deus rectissimi ascensor caeli auxiliator tuus magnificentia eius discurrunt nubes
DEUT|33|27|habitaculum eius sursum et subter brachia sempiterna eiciet a facie tua inimicum dicetque conterere
DEUT|33|28|habitabit Israhel confidenter et solus oculus Iacob in terra frumenti et vini caelique caligabunt rore
DEUT|33|29|beatus tu Israhel quis similis tui popule qui salvaris in Domino scutum auxilii tui et gladius gloriae tuae negabunt te inimici tui et tu eorum colla calcabis
DEUT|34|1|ascendit ergo Moses de campestribus Moab super montem Nebo in verticem Phasga contra Hiericho ostenditque ei Dominus omnem terram Galaad usque Dan
DEUT|34|2|et universum Nepthalim terramque Ephraim et Manasse et omnem terram usque ad mare Novissimum
DEUT|34|3|et australem partem et latitudinem campi Hiericho civitatis Palmarum usque Segor
DEUT|34|4|dixitque Dominus ad eum haec est terra pro qua iuravi Abraham Isaac et Iacob dicens semini tuo dabo eam vidisti eam oculis tuis et non transibis ad illam
DEUT|34|5|mortuusque est ibi Moses servus Domini in terra Moab iubente Domino
DEUT|34|6|et sepelivit eum in valle terrae Moab contra Phogor et non cognovit homo sepulchrum eius usque in praesentem diem
DEUT|34|7|Moses centum et viginti annorum erat quando mortuus est non caligavit oculus eius nec dentes illius moti sunt
DEUT|34|8|fleveruntque eum filii Israhel in campestribus Moab triginta diebus et conpleti sunt dies planctus lugentium Mosen
DEUT|34|9|Iosue vero filius Nun repletus est spiritu sapientiae quia Moses posuit super eum manus suas et oboedierunt ei filii Israhel feceruntque sicut praecepit Dominus Mosi
DEUT|34|10|et non surrexit propheta ultra in Israhel sicut Moses quem nosset Dominus facie ad faciem
DEUT|34|11|in omnibus signis atque portentis quae misit per eum ut faceret in terra Aegypti Pharaoni et omnibus servis eius universaeque terrae illius
DEUT|34|12|et cunctam manum robustam magnaque mirabilia quae fecit Moses coram universo Israhel
