1PET|1|1|Петро, апостол Ісуса Христа, захожанам Розпорошення: Понту, Галатії, Каппадокії, Азії й Віфінії, вибраним
1PET|1|2|із передбачення Бога Отця, посвяченням Духа, на покору й окроплення кров'ю Ісуса Христа: нехай примножиться вам благодать та мир!
1PET|1|3|Благословенний Бог і Отець Господа нашого Ісуса Христа, що великою Своєю милістю відродив нас до живої надії через воскресення з мертвих Ісуса Христа,
1PET|1|4|на спадщину нетлінну й непорочну та нев'янучу, заховану в небі для вас,
1PET|1|5|що ви бережені силою Божою через віру на спасіння, яке готове з'явитися останнього часу.
1PET|1|6|Тіштеся з того, засмучені трохи тепер, якщо треба, всілякими випробовуваннями,
1PET|1|7|щоб досвідчення вашої віри було дорогоцінніше за золото, яке гине, хоч і огнем випробовується, на похвалу, і честь, і славу при з'явленні Ісуса Христа.
1PET|1|8|Ви Його любите, не бачивши, і віруєте в Нього, хоч тепер не бачите, а вірувавши, радієте невимовною й славною радістю,
1PET|1|9|бо досягаєте мети віри вашої спасіння душам.
1PET|1|10|Про це спасіння розвідували та допитувалися пророки, що звіщали про благодать, призначену вам.
1PET|1|11|Вони досліджували, на котрий чи на який час показував Дух Христів, що в них був, коли Він сповіщав про Христові страждання та славу, що прийдуть по них.
1PET|1|12|Їм відкрито було, що вони не для себе самих, а для вас служили тим, що тепер звіщено вам через благовісників Духом Святим, із неба посланим, на що бажають дивитися Анголи.
1PET|1|13|Тому то, підперезавши стегна свого розуму та бувши тверезі, майте досконалу надію на благодать, що приноситься вам в з'явленні Ісуса Христа.
1PET|1|14|Як слухняні, не застосовуйтеся до попередніх пожадливостей вашого невідання,
1PET|1|15|але за Святим, що покликав вас, будьте й самі святі в усім вашім поводженні,
1PET|1|16|бо написано: Будьте святі, Я бо святий!
1PET|1|17|І коли ви Отцем звете Того, Хто кожного, не зважаючи на особу, судить за вчинок, то в страху провадьте час вашого тимчасового замешкання.
1PET|1|18|І знайте, що не тлінним сріблом або золотом відкуплені ви були від марного вашого життя, що передане вам від батьків,
1PET|1|19|але дорогоцінною кров'ю Христа, як непорочного й чистого Ягняти,
1PET|1|20|що призначений був іще перед закладинами світу, але був з'явлений вам за останнього часу.
1PET|1|21|Через Нього ви віруєте в Бога, що з мертвих Його воскресив та дав славу Йому, щоб була ваша віра й надія на Бога.
1PET|1|22|Послухом правді очистьте душі свої через Духа на нелицемірну братерську любов, і ревно від щирого серця любіть один одного,
1PET|1|23|бо народжені ви не з тлінного насіння, але з нетлінного, Словом Божим живим та тривалим.
1PET|1|24|Бо кожне тіло немов та трава, і всяка слава людини як цвіт трав'яний: засохне трава то й цвіт опаде,
1PET|1|25|а Слово Господнє повік пробуває! А це те Слово, яке звіщене вам в Євангелії.
1PET|2|1|Отож, відкладіть усяку злобу, і всякий підступ, і лицемірство, і заздрість, і всякі обмови,
1PET|2|2|і, немов новонароджені немовлята, жадайте щирого духовного молока, щоб ним вирости вам на спасіння,
1PET|2|3|якщо ви спробували, що добрий Господь.
1PET|2|4|Приступайте до Нього, до Каменя живого, дорогоцінного, що відкинули люди Його, але вибрав Бог.
1PET|2|5|І самі, немов те каміння живе, будуйтеся в дім духовий, на священство святе, щоб приносити жертви духовні, приємні для Бога через Ісуса Христа.
1PET|2|6|Бо стоїть у Писанні: Ось кладу Я на Сіоні Каменя вибраного, наріжного, дорогоцінного, і хто вірує в Нього, той не буде осоромлений!
1PET|2|7|Отож бо, для вас, хто вірує, Він коштовність, а для тих, хто не вірує камінь, що його занедбали були будівничі, той наріжним став каменем,
1PET|2|8|і камінь спотикання, і скеля спокуси, і об нього вони спотикаються, не вірячи слову, на що й призначені були.
1PET|2|9|Але ви вибраний рід, священство царське, народ святий, люд власности Божої, щоб звіщали чесноти Того, Хто покликав вас із темряви до дивного світла Свого,
1PET|2|10|колись ненарод, а тепер народ Божий, колись непомилувані, а тепер ви помилувані!
1PET|2|11|Благаю вас, любі, як приходьків та подорожніх, щоб ви здержувались від тілесних пожадливостей, що воюють проти душі.
1PET|2|12|Поводьтеся поміж поганами добре, щоб за те, за що вас обмовляють вони, немов би злочинців, побачивши добрі діла, славили Бога в день відвідання.
1PET|2|13|Отож, коріться кожному людському творінню ради Господа, чи то цареві, як найвищому,
1PET|2|14|чи то володарям, як від нього посланим для карання злочинців та для похвали доброчинців.
1PET|2|15|Бо така Божа воля, щоб доброчинці гамували неуцтво нерозумних людей,
1PET|2|16|як вільні, а не як ті, що мають волю на прикриття лихого, але як раби Божі.
1PET|2|17|Шануйте всіх, братство любіть, Бога бійтеся, царя поважайте.
1PET|2|18|Раби, коріться панам із повним страхом, не тільки добрим та тихим, але й прикрим.
1PET|2|19|Бо то вгодне, коли хто, через сумління перед Богом, терпить недолю, непоправді страждаючи.
1PET|2|20|Бо яка похвала, коли терпите ви, як вас б'ють за провини? Але коли з мукою терпите за добрі вчинки, то це вгодне Богові!
1PET|2|21|Бо на це ви покликані. Бо й Христос постраждав за нас, і залишив нам приклада, щоб пішли ми слідами Його.
1PET|2|22|Не вчинив Він гріха, і не знайшлося в устах Його підступу!
1PET|2|23|Коли був лихословлений, Він не лихословив взаємно, а коли Він страждав, не погрожував, але передав Тому, Хто судить справедливо.
1PET|2|24|Він тілом Своїм Сам підніс гріхи наші на дерево, щоб ми вмерли для гріхів та для праведности жили; Його ранами ви вздоровилися.
1PET|2|25|Ви бо були як ті вівці заблукані, та ви повернулись до Пастиря й Опікуна ваших душ.
1PET|3|1|Так само дружини, коріться своїм чоловікам, щоб і деякі, хто не кориться слову, були приєднані без слова поводженням дружин,
1PET|3|2|як побачать ваше поводження чисте в страху.
1PET|3|3|А окрасою їм нехай буде не зовнішнє, заплітання волосся та навішання золота або вбирання одеж,
1PET|3|4|але захована людина серця в нетлінні лагідного й мовчазного духа, що дорогоцінне перед Богом.
1PET|3|5|Бо так само колись прикрашали себе й святі ті жінки, що клали надію на Бога й корились своїм чоловікам.
1PET|3|6|Так Сара корилась Авраамові, і паном його називала. А ви її діти, коли добро робите та не лякаєтесь жадного страху.
1PET|3|7|Чоловіки, так само живіть разом із дружинами за розумом, як зо слабішою жіночою посудиною, і виявляйте їм честь, бо й вони є співспадкоємиці благодаті життя, щоб не спинялися ваші молитви.
1PET|3|8|Нарешті ж, будьте всі однодумні, спочутливі, братолюбні, милосердні, покірливі.
1PET|3|9|Не платіть злом за зло, або лайкою за лайку, навпаки, благословляйте, знавши, що на це вас покликано, щоб ви вспадкували благословення.
1PET|3|10|Бо хто хоче любити життя та бачити добрі дні, нехай здержить свого язика від лихого та уста свої від говорення підступу.
1PET|3|11|Ухиляйся від злого та добре чини, шукай миру й женися за ним!
1PET|3|12|Бо очі Господні до праведних, а вуха Його до їхніх прохань, а Господнє лице проти тих, хто чинить лихе!
1PET|3|13|І хто заподіє вам зле, коли будете ви оборонцями доброго?
1PET|3|14|А коли ви за правду й страждаєте, то ви блаженні! А їхнього страху не бійтеся, і не тривожтеся!
1PET|3|15|А Господа Христа святіть у ваших серцях, і завжди готовими будьте на відповідь кожному, хто в вас запитає рахунку про надію, що в вас, із лагідністю та зо страхом.
1PET|3|16|Майте добре сумління, щоб тим, за що вас обмовляють, немов би злочинців, були посоромлені лихословники вашого поводження в Христі.
1PET|3|17|Бо ліпше страждати за добрі діла, коли хоче того Божа воля, аніж за лихі.
1PET|3|18|Бо й Христос один раз постраждав був за наші гріхи, щоб привести нас до Бога, Праведний за неправедних, хоч умертвлений тілом, але Духом оживлений,
1PET|3|19|Яким Він і духам, що в в'язниці були, зійшовши, звіщав;
1PET|3|20|вони колись непокірливі були, як їх Боже довготерпіння чекало за Ноєвих днів, коли будувався ковчег, що в ньому мало, цебто вісім душ, спаслось від води.
1PET|3|21|Того образ, хрищення не тілесної нечистости позбуття, але обітниця Богові доброго сумління, спасає тепер і нас воскресенням Ісуса Христа,
1PET|3|22|що, зійшовши на небо, пробуває по Божій правиці, а Йому підкорилися Анголи, влади та сили.
1PET|4|1|Отож, коли тілом Христос постраждав за нас, то озбройтеся й ви тією самою думкою, бо хто тілом постраждав, той перестав грішити,
1PET|4|2|щоб решту часу в тілі жити вже не для пожадливостей людських, а для Божої волі.
1PET|4|3|Бо досить минулого часу, коли ви чинили волю поган, ходили в розпусті, у пожадливостях, у піяцтві, у гулянках, у піятиках, у беззаконних ідолослужбах.
1PET|4|4|Вони з того дивуються, що ви разом із ними не берете участи в розпусті, та зневажають.
1PET|4|5|Вони дадуть відповідь Тому, Хто судитиме живих та мертвих!
1PET|4|6|Бо на те й мертвим звіщувано Євангелію, щоб вони прийняли суд по-людському тілом, але жили по-Божому духом.
1PET|4|7|Кінець же всьому наблизився. Отже, будьте мудрі й пильнуйте в молитвах!
1PET|4|8|Найперше майте щиру любов один до одного, бо любов покриває багато гріхів!
1PET|4|9|Будьте гостинні один до одного без нехоті!
1PET|4|10|Служіть один одному, кожен тим даром, якого отримав, як доморядники всілякої Божої благодаті.
1PET|4|11|Коли хто говорить, говори, як Божі слова. Коли хто служить, то служи, як від сили, яку дає Бог, щоб Бог прославлявся в усьому Ісусом Христом, що Йому слава та влада на віки вічні, амінь.
1PET|4|12|Улюблені, не дивуйтесь огневі, що вам посилається на випробовування, немов би чужому випадку для вас.
1PET|4|13|Але через те, що берете ви участь у Христових стражданнях, то тіштеся, щоб і в з'явленні слави Його раділи ви й звеселялись.
1PET|4|14|Коли ж вас ганьблять за Христове Ім'я, то ви блаженні, бо на вас спочиває Дух слави й Дух Божий.
1PET|4|15|Ніхто з вас хай не страждає, як душогуб, або злодій, або злочинець, або ворохобник,
1PET|4|16|а коли як християнин, то нехай не соромиться він, але хай прославляє Бога за те.
1PET|4|17|Бо час уже суд розпочати від Божого дому; а коли він почнеться перше з нас, то який кінець тих, хто противиться Божій Євангелії?
1PET|4|18|А коли праведний ледве спасеться, то безбожний та грішний де зможе з'явитись?
1PET|4|19|Тому й ті, хто з Божої волі страждає, нехай душі свої віддадуть в доброчинстві Йому, як Створителю вірному.
1PET|5|1|Тож благаю між вами пресвітерів, співпресвітер та свідок Христових страждань, співучасник слави, що повинна з'явитись:
1PET|5|2|пасіть стадо Боже, що у вас, наглядайте не з примусу, але добровільно по-Божому, не для брудної наживи, а ревно,
1PET|5|3|не пануйте над спадком Божим, але будьте для стада за взір.
1PET|5|4|А коли Архипастир з'явиться, то одержите ви нев'янучого вінка слави.
1PET|5|5|Також молоді, коріться старшим! А всі майте покору один до одного, бо Бог противиться гордим, а смиренним дає благодать!
1PET|5|6|Тож покоріться під міцну Божу руку, щоб Він вас Свого часу повищив.
1PET|5|7|Покладіть на Нього всю вашу журбу, бо Він опікується вами!
1PET|5|8|Будьте тверезі, пильнуйте! Ваш супротивник диявол ходить, ричучи, як лев, що шукає пожерти кого.
1PET|5|9|Противтесь йому, тверді в вірі, знавши, що ті самі муки трапляються й вашому братству по світі.
1PET|5|10|А Бог усякої благодаті, що покликав вас до вічної слави Своєї в Христі, нехай Сам удосконалить вас, хто трохи потерпів, хай упевнить, зміцнить, уґрунтує.
1PET|5|11|Йому слава та влада на вічні віки, амінь.
1PET|5|12|Я коротко вам написав через Силуяна, як гадаю вірного брата. Закликаю та свідчу, що це Божа благодать правдива, що ви в ній стоїте.
1PET|5|13|Вітає вас разом вибрана Церква в Вавилоні, і Марко, мій син.
1PET|5|14|Вітайте один одного поцілунком любови. Мир вам усім у Христі! Амінь.
