ECCL|1|1|The words of the Preacher, the son of David, king in Jerusalem.
ECCL|1|2|Vanity of vanities, says the Preacher, vanity of vanities! All is vanity.
ECCL|1|3|What does man gain by all the toil at which he toils under the sun?
ECCL|1|4|A generation goes, and a generation comes, but the earth remains forever.
ECCL|1|5|The sun rises, and the sun goes down, and hastens to the place where it rises.
ECCL|1|6|The wind blows to the south and goes around to the north; around and around goes the wind, and on its circuits the wind returns.
ECCL|1|7|All streams run to the sea, but the sea is not full; to the place where the streams flow, there they flow again.
ECCL|1|8|All things are full of weariness; a man cannot utter it; the eye is not satisfied with seeing, nor the ear filled with hearing.
ECCL|1|9|What has been is what will be, and what has been done is what will be done, and there is nothing new under the sun.
ECCL|1|10|Is there a thing of which it is said, "See, this is new"? It has been already in the ages before us.
ECCL|1|11|There is no remembrance of former things, nor will there be any remembrance of later things yet to be among those who come after.
ECCL|1|12|I the Preacher have been king over Israel in Jerusalem.
ECCL|1|13|And I applied my heart to seek and to search out by wisdom all that is done under heaven. It is an unhappy business that God has given to the children of man to be busy with.
ECCL|1|14|I have seen everything that is done under the sun, and behold, all is vanity and a striving after wind.
ECCL|1|15|What is crooked cannot be made straight, and what is lacking cannot be counted.
ECCL|1|16|I said in my heart, "I have acquired great wisdom, surpassing all who were over Jerusalem before me, and my heart has had great experience of wisdom and knowledge."
ECCL|1|17|And I applied my heart to know wisdom and to know madness and folly. I perceived that this also is but a striving after wind.
ECCL|1|18|For in much wisdom is much vexation, and he who increases knowledge increases sorrow.
ECCL|2|1|I said in my heart, "Come now, I will test you with pleasure; enjoy yourself." But behold, this also was vanity.
ECCL|2|2|I said of laughter, "It is mad," and of pleasure, "What use is it?"
ECCL|2|3|I searched with my heart how to cheer my body with wine- my heart still guiding me with wisdom- and how to lay hold on folly, till I might see what was good for the children of man to do under heaven during the few days of their life.
ECCL|2|4|I made great works. I built houses and planted vineyards for myself.
ECCL|2|5|I made myself gardens and parks, and planted in them all kinds of fruit trees.
ECCL|2|6|I made myself pools from which to water the forest of growing trees.
ECCL|2|7|I bought male and female slaves, and had slaves who were born in my house. I had also great possessions of herds and flocks, more than any who had been before me in Jerusalem.
ECCL|2|8|I also gathered for myself silver and gold and the treasure of kings and provinces. I got singers, both men and women, and many concubines, the delight of the children of man.
ECCL|2|9|So I became great and surpassed all who were before me in Jerusalem. Also my wisdom remained with me.
ECCL|2|10|And whatever my eyes desired I did not keep from them. I kept my heart from no pleasure, for my heart found pleasure in all my toil, and this was my reward for all my toil.
ECCL|2|11|Then I considered all that my hands had done and the toil I had expended in doing it, and behold, all was vanity and a striving after wind, and there was nothing to be gained under the sun.
ECCL|2|12|So I turned to consider wisdom and madness and folly. For what can the man do who comes after the king? Only what has already been done.
ECCL|2|13|Then I saw that there is more gain in wisdom than in folly, as there is more gain in light than in darkness.
ECCL|2|14|The wise person has his eyes in his head, but the fool walks in darkness. And yet I perceived that the same event happens to all of them.
ECCL|2|15|Then I said in my heart, "What happens to the fool will happen to me also. Why then have I been so very wise?" And I said in my heart that this also is vanity.
ECCL|2|16|For of the wise as of the fool there is no enduring remembrance, seeing that in the days to come all will have been long forgotten. How the wise dies just like the fool!
ECCL|2|17|So I hated life, because what is done under the sun was grievous to me, for all is vanity and a striving after wind.
ECCL|2|18|I hated all my toil in which I toil under the sun, seeing that I must leave it to the man who will come after me,
ECCL|2|19|and who knows whether he will be wise or a fool? Yet he will be master of all for which I toiled and used my wisdom under the sun. This also is vanity.
ECCL|2|20|So I turned about and gave my heart up to despair over all the toil of my labors under the sun,
ECCL|2|21|because sometimes a person who has toiled with wisdom and knowledge and skill must leave everything to be enjoyed by someone who did not toil for it. This also is vanity and a great evil.
ECCL|2|22|What has a man from all the toil and striving of heart with which he toils beneath the sun?
ECCL|2|23|For all his days are full of sorrow, and his work is a vexation. Even in the night his heart does not rest. This also is vanity.
ECCL|2|24|There is nothing better for a person than that he should eat and drink and find enjoyment in his toil. This also, I saw, is from the hand of God,
ECCL|2|25|for apart from him who can eat or who can have enjoyment?
ECCL|2|26|For to the one who pleases him God has given wisdom and knowledge and joy, but to the sinner he has given the business of gathering and collecting, only to give to one who pleases God. This also is vanity and a striving after wind.
ECCL|3|1|For everything there is a season, and a time for every matter under heaven:
ECCL|3|2|a time to be born, and a time to die; a time to plant, and a time to pluck up what is planted;
ECCL|3|3|a time to kill, and a time to heal; a time to break down, and a time to build up;
ECCL|3|4|a time to weep, and a time to laugh; a time to mourn, and a time to dance;
ECCL|3|5|a time to cast away stones, and a time to gather stones together; a time to embrace, and a time to refrain from embracing;
ECCL|3|6|a time to seek, and a time to lose; a time to keep, and a time to cast away;
ECCL|3|7|a time to tear, and a time to sew; a time to keep silence, and a time to speak;
ECCL|3|8|a time to love, and a time to hate; a time for war, and a time for peace.
ECCL|3|9|What gain has the worker from his toil?
ECCL|3|10|I have seen the business that God has given to the children of man to be busy with.
ECCL|3|11|He has made everything beautiful in its time. Also, he has put eternity into man's heart, yet so that he cannot find out what God has done from the beginning to the end.
ECCL|3|12|I perceived that there is nothing better for them than to be joyful and to do good as long as they live;
ECCL|3|13|also that everyone should eat and drink and take pleasure in all his toil- this is God's gift to man.
ECCL|3|14|I perceived that whatever God does endures forever; nothing can be added to it, nor anything taken from it. God has done it, so that people fear before him.
ECCL|3|15|That which is, already has been; that which is to be, already has been; and God seeks what has been driven away.
ECCL|3|16|Moreover, I saw under the sun that in the place of justice, even there was wickedness, and in the place of righteousness, even there was wickedness.
ECCL|3|17|I said in my heart, God will judge the righteous and the wicked, for there is a time for every matter and for every work.
ECCL|3|18|I said in my heart with regard to the children of man that God is testing them that they may see that they themselves are but beasts.
ECCL|3|19|For what happens to the children of man and what happens to the beasts is the same; as one dies, so dies the other. They all have the same breath, and man has no advantage over the beasts, for all is vanity.
ECCL|3|20|All go to one place. All are from the dust, and to dust all return.
ECCL|3|21|Who knows whether the spirit of man goes upward and the spirit of the beast goes down into the earth?
ECCL|3|22|So I saw that there is nothing better than that a man should rejoice in his work, for that is his lot. Who can bring him to see what will be after him?
ECCL|4|1|Again I saw all the oppressions that are done under the sun. And behold, the tears of the oppressed, and they had no one to comfort them! On the side of their oppressors there was power, and there was no one to comfort them.
ECCL|4|2|And I thought the dead who are already dead more fortunate than the living who are still alive.
ECCL|4|3|But better than both is he who has not yet been and has not seen the evil deeds that are done under the sun.
ECCL|4|4|Then I saw that all toil and all skill in work come from a man's envy of his neighbor. This also is vanity and a striving after wind.
ECCL|4|5|The fool folds his hands and eats his own flesh.
ECCL|4|6|Better is a handful of quietness than two hands full of toil and a striving after wind.
ECCL|4|7|Again, I saw vanity under the sun:
ECCL|4|8|one person who has no other, either son or brother, yet there is no end to all his toil, and his eyes are never satisfied with riches, so that he never asks, "For whom am I toiling and depriving myself of pleasure?" This also is vanity and an unhappy business.
ECCL|4|9|Two are better than one, because they have a good reward for their toil.
ECCL|4|10|For if they fall, one will lift up his fellow. But woe to him who is alone when he falls and has not another to lift him up!
ECCL|4|11|Again, if two lie together, they keep warm, but how can one keep warm alone?
ECCL|4|12|And though a man might prevail against one who is alone, two will withstand him- a threefold cord is not quickly broken.
ECCL|4|13|Better was a poor and wise youth than an old and foolish king who no longer knew how to take advice.
ECCL|4|14|For he went from prison to the throne, though in his own kingdom he had been born poor.
ECCL|4|15|I saw all the living who move about under the sun, along with that youth who was to stand in the king's place.
ECCL|4|16|There was no end of all the people, all of whom he led. Yet those who come later will not rejoice in him. Surely this also is vanity and a striving after wind.
ECCL|5|1|Guard your steps when you go to the house of God. To draw near to listen is better than to offer the sacrifice of fools, for they do not know that they are doing evil.
ECCL|5|2|Be not rash with your mouth, nor let your heart be hasty to utter a word before God, for God is in heaven and you are on earth. Therefore let your words be few.
ECCL|5|3|For a dream comes with much business, and a fool's voice with many words.
ECCL|5|4|When you vow a vow to God, do not delay paying it, for he has no pleasure in fools. Pay what you vow.
ECCL|5|5|It is better that you should not vow than that you should vow and not pay.
ECCL|5|6|Let not your mouth lead you into sin, and do not say before the messenger that it was a mistake. Why should God be angry at your voice and destroy the work of your hands?
ECCL|5|7|For when dreams increase and words grow many, there is vanity; but God is the one you must fear.
ECCL|5|8|If you see in a province the oppression of the poor and the violation of justice and righteousness, do not be amazed at the matter, for the high official is watched by a higher, and there are yet higher ones over them.
ECCL|5|9|But this is gain for a land in every way: a king committed to cultivated fields.
ECCL|5|10|He who loves money will not be satisfied with money, nor he who loves wealth with his income; this also is vanity.
ECCL|5|11|When goods increase, they increase who eat them, and what advantage has their owner but to see them with his eyes?
ECCL|5|12|Sweet is the sleep of a laborer, whether he eats little or much, but the full stomach of the rich will not let him sleep.
ECCL|5|13|There is a grievous evil that I have seen under the sun: riches were kept by their owner to his hurt,
ECCL|5|14|and those riches were lost in a bad venture. And he is father of a son, but he has nothing in his hand.
ECCL|5|15|As he came from his mother's womb he shall go again, naked as he came, and shall take nothing for his toil that he may carry away in his hand.
ECCL|5|16|This also is a grievous evil: just as he came, so shall he go, and what gain is there to him who toils for the wind?
ECCL|5|17|Moreover, all his days he eats in darkness in much vexation and sickness and anger.
ECCL|5|18|Behold, what I have seen to be good and fitting is to eat and drink and find enjoyment in all the toil with which one toils under the sun the few days of his life that God has given him, for this is his lot.
ECCL|5|19|Everyone also to whom God has given wealth and possessions and power to enjoy them, and to accept his lot and rejoice in his toil- this is the gift of God.
ECCL|5|20|For he will not much remember the days of his life because God keeps him occupied with joy in his heart.
ECCL|6|1|There is an evil that I have seen under the sun, and it lies heavy on mankind:
ECCL|6|2|a man to whom God gives wealth, possessions, and honor, so that he lacks nothing of all that he desires, yet God does not give him power to enjoy them, but a stranger enjoys them. This is vanity; it is a grievous evil.
ECCL|6|3|If a man fathers a hundred children and lives many years, so that the days of his years are many, but his soul is not satisfied with life's good things, and he also has no burial, I say that a stillborn child is better off than he.
ECCL|6|4|For it comes in vanity and goes in darkness, and in darkness its name is covered.
ECCL|6|5|Moreover, it has not seen the sun or known anything, yet it finds rest rather than he.
ECCL|6|6|Even though he should live a thousand years twice over, yet enjoy no good- do not all go to the one place?
ECCL|6|7|All the toil of man is for his mouth, yet his appetite is not satisfied.
ECCL|6|8|For what advantage has the wise man over the fool? And what does the poor man have who knows how to conduct himself before the living?
ECCL|6|9|Better is the sight of the eyes than the wandering of the appetite: this also is vanity and a striving after wind.
ECCL|6|10|Whatever has come to be has already been named, and it is known what man is, and that he is not able to dispute with one stronger than he.
ECCL|6|11|The more words, the more vanity, and what is the advantage to man?
ECCL|6|12|For who knows what is good for man while he lives the few days of his vain life, which he passes like a shadow? For who can tell man what will be after him under the sun?
ECCL|7|1|A good name is better than precious ointment, and the day of death than the day of birth.
ECCL|7|2|It is better to go to the house of mourning than to go to the house of feasting, for this is the end of all mankind, and the living will lay it to heart.
ECCL|7|3|Sorrow is better than laughter, for by sadness of face the heart is made glad.
ECCL|7|4|The heart of the wise is in the house of mourning, but the heart of fools is in the house of mirth.
ECCL|7|5|It is better for a man to hear the rebuke of the wise than to hear the song of fools.
ECCL|7|6|For as the crackling of thorns under a pot, so is the laughter of the fools; this also is vanity.
ECCL|7|7|Surely oppression drives the wise into madness, and a bribe corrupts the heart.
ECCL|7|8|Better is the end of a thing than its beginning, and the patient in spirit is better than the proud in spirit.
ECCL|7|9|Be not quick in your spirit to become angry, for anger lodges in the bosom of fools.
ECCL|7|10|Say not, "Why were the former days better than these?" For it is not from wisdom that you ask this.
ECCL|7|11|Wisdom is good with an inheritance, an advantage to those who see the sun.
ECCL|7|12|For the protection of wisdom is like the protection of money, and the advantage of knowledge is that wisdom preserves the life of him who has it.
ECCL|7|13|Consider the work of God: who can make straight what he has made crooked?
ECCL|7|14|In the day of prosperity be joyful, and in the day of adversity consider: God has made the one as well as the other, so that man may not find out anything that will be after him.
ECCL|7|15|In my vain life I have seen everything. There is a righteous man who perishes in his righteousness, and there is a wicked man who prolongs his life in his evildoing.
ECCL|7|16|Be not overly righteous, and do not make yourself too wise. Why should you destroy yourself?
ECCL|7|17|Be not overly wicked, neither be a fool. Why should you die before your time?
ECCL|7|18|It is good that you should take hold of this, and from that withhold not your hand, for the one who fears God shall come out from both of them.
ECCL|7|19|Wisdom gives strength to the wise man more than ten rulers who are in a city.
ECCL|7|20|Surely there is not a righteous man on earth who does good and never sins.
ECCL|7|21|Do not take to heart all the things that people say, lest you hear your servant cursing you.
ECCL|7|22|Your heart knows that many times you have yourself cursed others.
ECCL|7|23|All this I have tested by wisdom. I said, "I will be wise," but it was far from me.
ECCL|7|24|That which has been is far off, and deep, very deep; who can find it out?
ECCL|7|25|I turned my heart to know and to search out and to seek wisdom and the scheme of things, and to know the wickedness of folly and the foolishness that is madness.
ECCL|7|26|And I find something more bitter than death: the woman whose heart is snares and nets, and whose hands are fetters. He who pleases God escapes her, but the sinner is taken by her.
ECCL|7|27|Behold, this is what I found, says the Preacher, while adding one thing to another to find the scheme of things-
ECCL|7|28|which my soul has sought repeatedly, but I have not found. One man among a thousand I found, but a woman among all these I have not found.
ECCL|7|29|See, this alone I found, that God made man upright, but they have sought out many schemes.
ECCL|8|1|Who is like the wise?And who knows the interpretation of a thing? A man's wisdom makes his face shine, and the hardness of his face is changed.
ECCL|8|2|I say: Keep the king's command, because of God's oath to him.
ECCL|8|3|Be not hasty to go from his presence. Do not take your stand in an evil cause, for he does whatever he pleases.
ECCL|8|4|For the word of the king is supreme, and who may say to him, "What are you doing?"
ECCL|8|5|Whoever keeps a command will know no evil thing, and the wise heart will know the proper time and the just way.
ECCL|8|6|For there is a time and a way for everything, although man's trouble lies heavy on him.
ECCL|8|7|For he does not know what is to be, for who can tell him how it will be?
ECCL|8|8|No man has power to retain the spirit, or power over the day of death. There is no discharge from war, nor will wickedness deliver those who are given to it.
ECCL|8|9|All this I observed while applying my heart to all that is done under the sun, when man had power over man to his hurt.
ECCL|8|10|Then I saw the wicked buried. They used to go in and out of the holy place and were praised in the city where they had done such things. This also is vanity.
ECCL|8|11|Because the sentence against an evil deed is not executed speedily, the heart of the children of man is fully set to do evil.
ECCL|8|12|Though a sinner does evil a hundred times and prolongs his life, yet I know that it will be well with those who fear God, because they fear before him.
ECCL|8|13|But it will not be well with the wicked, neither will he prolong his days like a shadow, because he does not fear before God.
ECCL|8|14|There is a vanity that takes place on earth, that there are righteous people to whom it happens according to the deeds of the wicked, and there are wicked people to whom it happens according to the deeds of the righteous. I said that this also is vanity.
ECCL|8|15|And I commend joy, for man has no good thing under the sun but to eat and drink and be joyful, for this will go with him in his toil through the days of his life that God has given him under the sun.
ECCL|8|16|When I applied my heart to know wisdom, and to see the business that is done on earth, how neither day nor night do one's eyes see sleep,
ECCL|8|17|then I saw all the work of God, that man cannot find out the work that is done under the sun. However much man may toil in seeking, he will not find it out. Even though a wise man claims to know, he cannot find it out.
ECCL|9|1|But all this I laid to heart, examining it all, how the righteous and the wise and their deeds are in the hand of God. Whether it is love or hate, man does not know; both are before him.
ECCL|9|2|It is the same for all, since the same event happens to the righteous and the wicked, to the good and the evil, to the clean and the unclean, to him who sacrifices and him who does not sacrifice. As is the good, so is the sinner, and he who swears is as he who shuns an oath.
ECCL|9|3|This is an evil in all that is done under the sun, that the same event happens to all. Also, the hearts of the children of man are full of evil, and madness is in their hearts while they live, and after that they go to the dead.
ECCL|9|4|But he who is joined with all the living has hope, for a living dog is better than a dead lion.
ECCL|9|5|For the living know that they will die, but the dead know nothing, and they have no more reward, for the memory of them is forgotten.
ECCL|9|6|Their love and their hate and their envy have already perished, and forever they have no more share in all that is done under the sun.
ECCL|9|7|Go, eat your bread in joy, and drink your wine with a merry heart, for God has already approved what you do.
ECCL|9|8|Let your garments be always white. Let not oil be lacking on your head.
ECCL|9|9|Enjoy life with the wife whom you love, all the days of your vain life that he has given you under the sun, because that is your portion in life and in your toil at which you toil under the sun.
ECCL|9|10|Whatever your hand finds to do, do it with your might, for there is no work or thought or knowledge or wisdom in Sheol, to which you are going.
ECCL|9|11|Again I saw that under the sun the race is not to the swift, nor the battle to the strong, nor bread to the wise, nor riches to the intelligent, nor favor to those with knowledge, but time and chance happen to them all.
ECCL|9|12|For man does not know his time. Like fish that are taken in an evil net, and like birds that are caught in a snare, so the children of man are snared at an evil time, when it suddenly falls upon them.
ECCL|9|13|I have also seen this example of wisdom under the sun, and it seemed great to me.
ECCL|9|14|There was a little city with few men in it, and a great king came against it and besieged it, building great siegeworks against it.
ECCL|9|15|But there was found in it a poor, wise man, and he by his wisdom delivered the city. Yet no one remembered that poor man.
ECCL|9|16|But I say that wisdom is better than might, though the poor man's wisdom is despised and his words are not heard.
ECCL|9|17|The words of the wise heard in quiet are better than the shouting of a ruler among fools.
ECCL|9|18|Wisdom is better than weapons of war, but one sinner destroys much good.
ECCL|10|1|Dead flies make the perfumer's ointment give off a stench; so a little folly outweighs wisdom and honor.
ECCL|10|2|A wise man's heart inclines him to the right, but a fool's heart to the left.
ECCL|10|3|Even when the fool walks on the road, he lacks sense, and he says to everyone that he is a fool.
ECCL|10|4|If the anger of the ruler rises against you, do not leave your place, for calmness will lay great offenses to rest.
ECCL|10|5|There is an evil that I have seen under the sun, as it were an error proceeding from the ruler:
ECCL|10|6|folly is set in many high places, and the rich sit in a low place.
ECCL|10|7|I have seen slaves on horses, and princes walking on the ground like slaves.
ECCL|10|8|He who digs a pit will fall into it, and a serpent will bite him who breaks through a wall.
ECCL|10|9|He who quarries stones is hurt by them, and he who splits logs is endangered by them.
ECCL|10|10|If the iron is blunt, and one does not sharpen the edge, he must use more strength, but wisdom helps one to succeed.
ECCL|10|11|If the serpent bites before it is charmed, there is no advantage to the charmer.
ECCL|10|12|The words of a wise man's mouth win him favor, but the lips of a fool consume him.
ECCL|10|13|The beginning of the words of his mouth is foolishness, and the end of his talk is evil madness.
ECCL|10|14|A fool multiplies words, though no man knows what is to be, and who can tell him what will be after him?
ECCL|10|15|The toil of a fool wearies him, for he does not know the way to the city.
ECCL|10|16|Woe to you, O land, when your king is a child, and your princes feast in the morning!
ECCL|10|17|Happy are you, O land, when your king is the son of the nobility, and your princes feast at the proper time, for strength, and not for drunkenness!
ECCL|10|18|Through sloth the roof sinks in, and through indolence the house leaks.
ECCL|10|19|Bread is made for laughter, and wine gladdens life, and money answers everything.
ECCL|10|20|Even in your thought, do not curse the king, nor in your bedroom curse the rich, for a bird of the air will carry your voice, or some winged creature tell the matter.
ECCL|11|1|Cast your bread upon the waters, for you will find it after many days.
ECCL|11|2|Give a portion to seven, or even to eight, for you know not what disaster may happen on earth.
ECCL|11|3|If the clouds are full of rain, they empty themselves on the earth, and if a tree falls to the south or to the north, in the place where the tree falls, there it will lie.
ECCL|11|4|He who observes the wind will not sow, and he who regards the clouds will not reap.
ECCL|11|5|As you do not know the way the spirit comes to the bones in the womb of a woman with child, so you do not know the work of God who makes everything.
ECCL|11|6|In the morning sow your seed, and at evening withhold not your hand, for you do not know which will prosper, this or that, or whether both alike will be good.
ECCL|11|7|Light is sweet, and it is pleasant for the eyes to see the sun.
ECCL|11|8|So if a person lives many years, let him rejoice in them all; but let him remember that the days of darkness will be many. All that comes is vanity.
ECCL|11|9|Rejoice, O young man, in your youth, and let your heart cheer you in the days of your youth. Walk in the ways of your heart and the sight of your eyes. But know that for all these things God will bring you into judgment.
ECCL|11|10|Remove vexation from your heart, and put away pain from your body, for youth and the dawn of life are vanity.
ECCL|12|1|Remember also your Creator in the days of your youth, before the evil days come and the years draw near of which you will say, "I have no pleasure in them";
ECCL|12|2|before the sun and the light and the moon and the stars are darkened and the clouds return after the rain,
ECCL|12|3|in the day when the keepers of the house tremble, and the strong men are bent, and the grinders cease because they are few, and those who look through the windows are dimmed,
ECCL|12|4|and the doors on the street are shut- when the sound of the grinding is low, and one rises up at the sound of a bird, and all the daughters of song are brought low-
ECCL|12|5|they are afraid also of what is high, and terrors are in the way; the almond tree blossoms, the grasshopper drags itself along, and desire fails, because man is going to his eternal home, and the mourners go about the streets-
ECCL|12|6|before the silver cord is snapped, or the golden bowl is broken, or the pitcher is shattered at the fountain, or the wheel broken at the cistern,
ECCL|12|7|and the dust returns to the earth as it was, and the spirit returns to God who gave it.
ECCL|12|8|Vanity of vanities, says the Preacher; all is vanity.
ECCL|12|9|Besides being wise, the Preacher also taught the people knowledge, weighing and studying and arranging many proverbs with great care.
ECCL|12|10|The Preacher sought to find words of delight, and uprightly he wrote words of truth.
ECCL|12|11|The words of the wise are like goads, and like nails firmly fixed are the collected sayings; they are given by one Shepherd.
ECCL|12|12|My son, beware of anything beyond these. Of making many books there is no end, and much study is a weariness of the flesh.
ECCL|12|13|The end of the matter; all has been heard. Fear God and keep his commandments, for this is the whole duty of man.
ECCL|12|14|For God will bring every deed into judgment, with every secret thing, whether good or evil.
