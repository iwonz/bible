EZEK|1|1|In the thirtieth year, in the fourth month on the fifth day, while I was among the exiles by the Kebar River, the heavens were opened and I saw visions of God.
EZEK|1|2|On the fifth of the month-it was the fifth year of the exile of King Jehoiachin-
EZEK|1|3|the word of the LORD came to Ezekiel the priest, the son of Buzi, by the Kebar River in the land of the Babylonians. There the hand of the LORD was upon him.
EZEK|1|4|I looked, and I saw a windstorm coming out of the north-an immense cloud with flashing lightning and surrounded by brilliant light. The center of the fire looked like glowing metal,
EZEK|1|5|and in the fire was what looked like four living creatures. In appearance their form was that of a man,
EZEK|1|6|but each of them had four faces and four wings.
EZEK|1|7|Their legs were straight; their feet were like those of a calf and gleamed like burnished bronze.
EZEK|1|8|Under their wings on their four sides they had the hands of a man. All four of them had faces and wings,
EZEK|1|9|and their wings touched one another. Each one went straight ahead; they did not turn as they moved.
EZEK|1|10|Their faces looked like this: Each of the four had the face of a man, and on the right side each had the face of a lion, and on the left the face of an ox; each also had the face of an eagle.
EZEK|1|11|Such were their faces. Their wings were spread out upward; each had two wings, one touching the wing of another creature on either side, and two wings covering its body.
EZEK|1|12|Each one went straight ahead. Wherever the spirit would go, they would go, without turning as they went.
EZEK|1|13|The appearance of the living creatures was like burning coals of fire or like torches. Fire moved back and forth among the creatures; it was bright, and lightning flashed out of it.
EZEK|1|14|The creatures sped back and forth like flashes of lightning.
EZEK|1|15|As I looked at the living creatures, I saw a wheel on the ground beside each creature with its four faces.
EZEK|1|16|This was the appearance and structure of the wheels: They sparkled like chrysolite, and all four looked alike. Each appeared to be made like a wheel intersecting a wheel.
EZEK|1|17|As they moved, they would go in any one of the four directions the creatures faced; the wheels did not turn about as the creatures went.
EZEK|1|18|Their rims were high and awesome, and all four rims were full of eyes all around.
EZEK|1|19|When the living creatures moved, the wheels beside them moved; and when the living creatures rose from the ground, the wheels also rose.
EZEK|1|20|Wherever the spirit would go, they would go, and the wheels would rise along with them, because the spirit of the living creatures was in the wheels.
EZEK|1|21|When the creatures moved, they also moved; when the creatures stood still, they also stood still; and when the creatures rose from the ground, the wheels rose along with them, because the spirit of the living creatures was in the wheels.
EZEK|1|22|Spread out above the heads of the living creatures was what looked like an expanse, sparkling like ice, and awesome.
EZEK|1|23|Under the expanse their wings were stretched out one toward the other, and each had two wings covering its body.
EZEK|1|24|When the creatures moved, I heard the sound of their wings, like the roar of rushing waters, like the voice of the Almighty, like the tumult of an army. When they stood still, they lowered their wings.
EZEK|1|25|Then there came a voice from above the expanse over their heads as they stood with lowered wings.
EZEK|1|26|Above the expanse over their heads was what looked like a throne of sapphire, and high above on the throne was a figure like that of a man.
EZEK|1|27|I saw that from what appeared to be his waist up he looked like glowing metal, as if full of fire, and that from there down he looked like fire; and brilliant light surrounded him.
EZEK|1|28|Like the appearance of a rainbow in the clouds on a rainy day, so was the radiance around him. This was the appearance of the likeness of the glory of the LORD. When I saw it, I fell facedown, and I heard the voice of one speaking.
EZEK|2|1|He said to me, "Son of man, stand up on your feet and I will speak to you."
EZEK|2|2|As he spoke, the Spirit came into me and raised me to my feet, and I heard him speaking to me.
EZEK|2|3|He said: "Son of man, I am sending you to the Israelites, to a rebellious nation that has rebelled against me; they and their fathers have been in revolt against me to this very day.
EZEK|2|4|The people to whom I am sending you are obstinate and stubborn. Say to them, 'This is what the Sovereign LORD says.'
EZEK|2|5|And whether they listen or fail to listen-for they are a rebellious house-they will know that a prophet has been among them.
EZEK|2|6|And you, son of man, do not be afraid of them or their words. Do not be afraid, though briers and thorns are all around you and you live among scorpions. Do not be afraid of what they say or terrified by them, though they are a rebellious house.
EZEK|2|7|You must speak my words to them, whether they listen or fail to listen, for they are rebellious.
EZEK|2|8|But you, son of man, listen to what I say to you. Do not rebel like that rebellious house; open your mouth and eat what I give you."
EZEK|2|9|Then I looked, and I saw a hand stretched out to me. In it was a scroll,
EZEK|2|10|which he unrolled before me. On both sides of it were written words of lament and mourning and woe.
EZEK|3|1|And he said to me, "Son of man, eat what is before you, eat this scroll; then go and speak to the house of Israel."
EZEK|3|2|So I opened my mouth, and he gave me the scroll to eat.
EZEK|3|3|Then he said to me, "Son of man, eat this scroll I am giving you and fill your stomach with it." So I ate it, and it tasted as sweet as honey in my mouth.
EZEK|3|4|He then said to me: "Son of man, go now to the house of Israel and speak my words to them.
EZEK|3|5|You are not being sent to a people of obscure speech and difficult language, but to the house of Israel-
EZEK|3|6|not to many peoples of obscure speech and difficult language, whose words you cannot understand. Surely if I had sent you to them, they would have listened to you.
EZEK|3|7|But the house of Israel is not willing to listen to you because they are not willing to listen to me, for the whole house of Israel is hardened and obstinate.
EZEK|3|8|But I will make you as unyielding and hardened as they are.
EZEK|3|9|I will make your forehead like the hardest stone, harder than flint. Do not be afraid of them or terrified by them, though they are a rebellious house."
EZEK|3|10|And he said to me, "Son of man, listen carefully and take to heart all the words I speak to you.
EZEK|3|11|Go now to your countrymen in exile and speak to them. Say to them, 'This is what the Sovereign LORD says,' whether they listen or fail to listen."
EZEK|3|12|Then the Spirit lifted me up, and I heard behind me a loud rumbling sound-May the glory of the LORD be praised in his dwelling place!-
EZEK|3|13|the sound of the wings of the living creatures brushing against each other and the sound of the wheels beside them, a loud rumbling sound.
EZEK|3|14|The Spirit then lifted me up and took me away, and I went in bitterness and in the anger of my spirit, with the strong hand of the LORD upon me.
EZEK|3|15|I came to the exiles who lived at Tel Abib near the Kebar River. And there, where they were living, I sat among them for seven days-overwhelmed.
EZEK|3|16|At the end of seven days the word of the LORD came to me:
EZEK|3|17|"Son of man, I have made you a watchman for the house of Israel; so hear the word I speak and give them warning from me.
EZEK|3|18|When I say to a wicked man, 'You will surely die,' and you do not warn him or speak out to dissuade him from his evil ways in order to save his life, that wicked man will die for his sin, and I will hold you accountable for his blood.
EZEK|3|19|But if you do warn the wicked man and he does not turn from his wickedness or from his evil ways, he will die for his sin; but you will have saved yourself.
EZEK|3|20|"Again, when a righteous man turns from his righteousness and does evil, and I put a stumbling block before him, he will die. Since you did not warn him, he will die for his sin. The righteous things he did will not be remembered, and I will hold you accountable for his blood.
EZEK|3|21|But if you do warn the righteous man not to sin and he does not sin, he will surely live because he took warning, and you will have saved yourself."
EZEK|3|22|The hand of the LORD was upon me there, and he said to me, "Get up and go out to the plain, and there I will speak to you."
EZEK|3|23|So I got up and went out to the plain. And the glory of the LORD was standing there, like the glory I had seen by the Kebar River, and I fell facedown.
EZEK|3|24|Then the Spirit came into me and raised me to my feet. He spoke to me and said: "Go, shut yourself inside your house.
EZEK|3|25|And you, son of man, they will tie with ropes; you will be bound so that you cannot go out among the people.
EZEK|3|26|I will make your tongue stick to the roof of your mouth so that you will be silent and unable to rebuke them, though they are a rebellious house.
EZEK|3|27|But when I speak to you, I will open your mouth and you shall say to them, 'This is what the Sovereign LORD says.' Whoever will listen let him listen, and whoever will refuse let him refuse; for they are a rebellious house.
EZEK|4|1|"Now, son of man, take a clay tablet, put it in front of you and draw the city of Jerusalem on it.
EZEK|4|2|Then lay siege to it: Erect siege works against it, build a ramp up to it, set up camps against it and put battering rams around it.
EZEK|4|3|Then take an iron pan, place it as an iron wall between you and the city and turn your face toward it. It will be under siege, and you shall besiege it. This will be a sign to the house of Israel.
EZEK|4|4|"Then lie on your left side and put the sin of the house of Israel upon yourself. You are to bear their sin for the number of days you lie on your side.
EZEK|4|5|I have assigned you the same number of days as the years of their sin. So for 390 days you will bear the sin of the house of Israel.
EZEK|4|6|"After you have finished this, lie down again, this time on your right side, and bear the sin of the house of Judah. I have assigned you 40 days, a day for each year.
EZEK|4|7|Turn your face toward the siege of Jerusalem and with bared arm prophesy against her.
EZEK|4|8|I will tie you up with ropes so that you cannot turn from one side to the other until you have finished the days of your siege.
EZEK|4|9|"Take wheat and barley, beans and lentils, millet and spelt; put them in a storage jar and use them to make bread for yourself. You are to eat it during the 390 days you lie on your side.
EZEK|4|10|Weigh out twenty shekels of food to eat each day and eat it at set times.
EZEK|4|11|Also measure out a sixth of a hin of water and drink it at set times.
EZEK|4|12|Eat the food as you would a barley cake; bake it in the sight of the people, using human excrement for fuel."
EZEK|4|13|The LORD said, "In this way the people of Israel will eat defiled food among the nations where I will drive them."
EZEK|4|14|Then I said, "Not so, Sovereign LORD! I have never defiled myself. From my youth until now I have never eaten anything found dead or torn by wild animals. No unclean meat has ever entered my mouth."
EZEK|4|15|"Very well," he said, "I will let you bake your bread over cow manure instead of human excrement."
EZEK|4|16|He then said to me: "Son of man, I will cut off the supply of food in Jerusalem. The people will eat rationed food in anxiety and drink rationed water in despair,
EZEK|4|17|for food and water will be scarce. They will be appalled at the sight of each other and will waste away because of their sin.
EZEK|5|1|"Now, son of man, take a sharp sword and use it as a barber's razor to shave your head and your beard. Then take a set of scales and divide up the hair.
EZEK|5|2|When the days of your siege come to an end, burn a third of the hair with fire inside the city. Take a third and strike it with the sword all around the city. And scatter a third to the wind. For I will pursue them with drawn sword.
EZEK|5|3|But take a few strands of hair and tuck them away in the folds of your garment.
EZEK|5|4|Again, take a few of these and throw them into the fire and burn them up. A fire will spread from there to the whole house of Israel.
EZEK|5|5|"This is what the Sovereign LORD says: This is Jerusalem, which I have set in the center of the nations, with countries all around her.
EZEK|5|6|Yet in her wickedness she has rebelled against my laws and decrees more than the nations and countries around her. She has rejected my laws and has not followed my decrees.
EZEK|5|7|"Therefore this is what the Sovereign LORD says: You have been more unruly than the nations around you and have not followed my decrees or kept my laws. You have not even conformed to the standards of the nations around you.
EZEK|5|8|"Therefore this is what the Sovereign LORD says: I myself am against you, Jerusalem, and I will inflict punishment on you in the sight of the nations.
EZEK|5|9|Because of all your detestable idols, I will do to you what I have never done before and will never do again.
EZEK|5|10|Therefore in your midst fathers will eat their children, and children will eat their fathers. I will inflict punishment on you and will scatter all your survivors to the winds.
EZEK|5|11|Therefore as surely as I live, declares the Sovereign LORD, because you have defiled my sanctuary with all your vile images and detestable practices, I myself will withdraw my favor; I will not look on you with pity or spare you.
EZEK|5|12|A third of your people will die of the plague or perish by famine inside you; a third will fall by the sword outside your walls; and a third I will scatter to the winds and pursue with drawn sword.
EZEK|5|13|"Then my anger will cease and my wrath against them will subside, and I will be avenged. And when I have spent my wrath upon them, they will know that I the LORD have spoken in my zeal.
EZEK|5|14|"I will make you a ruin and a reproach among the nations around you, in the sight of all who pass by.
EZEK|5|15|You will be a reproach and a taunt, a warning and an object of horror to the nations around you when I inflict punishment on you in anger and in wrath and with stinging rebuke. I the LORD have spoken.
EZEK|5|16|When I shoot at you with my deadly and destructive arrows of famine, I will shoot to destroy you. I will bring more and more famine upon you and cut off your supply of food.
EZEK|5|17|I will send famine and wild beasts against you, and they will leave you childless. Plague and bloodshed will sweep through you, and I will bring the sword against you. I the LORD have spoken."
EZEK|6|1|The word of the LORD came to me:
EZEK|6|2|"Son of man, set your face against the mountains of Israel; prophesy against them
EZEK|6|3|and say: 'O mountains of Israel, hear the word of the Sovereign LORD. This is what the Sovereign LORD says to the mountains and hills, to the ravines and valleys: I am about to bring a sword against you, and I will destroy your high places.
EZEK|6|4|Your altars will be demolished and your incense altars will be smashed; and I will slay your people in front of your idols.
EZEK|6|5|I will lay the dead bodies of the Israelites in front of their idols, and I will scatter your bones around your altars.
EZEK|6|6|Wherever you live, the towns will be laid waste and the high places demolished, so that your altars will be laid waste and devastated, your idols smashed and ruined, your incense altars broken down, and what you have made wiped out.
EZEK|6|7|Your people will fall slain among you, and you will know that I am the LORD.
EZEK|6|8|"'But I will spare some, for some of you will escape the sword when you are scattered among the lands and nations.
EZEK|6|9|Then in the nations where they have been carried captive, those who escape will remember me-how I have been grieved by their adulterous hearts, which have turned away from me, and by their eyes, which have lusted after their idols. They will loathe themselves for the evil they have done and for all their detestable practices.
EZEK|6|10|And they will know that I am the LORD; I did not threaten in vain to bring this calamity on them.
EZEK|6|11|"'This is what the Sovereign LORD says: Strike your hands together and stamp your feet and cry out "Alas!" because of all the wicked and detestable practices of the house of Israel, for they will fall by the sword, famine and plague.
EZEK|6|12|He that is far away will die of the plague, and he that is near will fall by the sword, and he that survives and is spared will die of famine. So will I spend my wrath upon them.
EZEK|6|13|And they will know that I am the LORD, when their people lie slain among their idols around their altars, on every high hill and on all the mountaintops, under every spreading tree and every leafy oak-places where they offered fragrant incense to all their idols.
EZEK|6|14|And I will stretch out my hand against them and make the land a desolate waste from the desert to Diblah -wherever they live. Then they will know that I am the LORD.'"
EZEK|7|1|The word of the LORD came to me:
EZEK|7|2|"Son of man, this is what the Sovereign LORD says to the land of Israel: The end! The end has come upon the four corners of the land.
EZEK|7|3|The end is now upon you and I will unleash my anger against you. I will judge you according to your conduct and repay you for all your detestable practices.
EZEK|7|4|I will not look on you with pity or spare you; I will surely repay you for your conduct and the detestable practices among you. Then you will know that I am the LORD.
EZEK|7|5|"This is what the Sovereign LORD says: Disaster! An unheard-of disaster is coming.
EZEK|7|6|The end has come! The end has come! It has roused itself against you. It has come!
EZEK|7|7|Doom has come upon you-you who dwell in the land. The time has come, the day is near; there is panic, not joy, upon the mountains.
EZEK|7|8|I am about to pour out my wrath on you and spend my anger against you; I will judge you according to your conduct and repay you for all your detestable practices.
EZEK|7|9|I will not look on you with pity or spare you; I will repay you in accordance with your conduct and the detestable practices among you. Then you will know that it is I the LORD who strikes the blow.
EZEK|7|10|"The day is here! It has come! Doom has burst forth, the rod has budded, arrogance has blossomed!
EZEK|7|11|Violence has grown into a rod to punish wickedness; none of the people will be left, none of that crowd-no wealth, nothing of value.
EZEK|7|12|The time has come, the day has arrived. Let not the buyer rejoice nor the seller grieve, for wrath is upon the whole crowd.
EZEK|7|13|The seller will not recover the land he has sold as long as both of them live, for the vision concerning the whole crowd will not be reversed. Because of their sins, not one of them will preserve his life.
EZEK|7|14|Though they blow the trumpet and get everything ready, no one will go into battle, for my wrath is upon the whole crowd.
EZEK|7|15|"Outside is the sword, inside are plague and famine; those in the country will die by the sword, and those in the city will be devoured by famine and plague.
EZEK|7|16|All who survive and escape will be in the mountains, moaning like doves of the valleys, each because of his sins.
EZEK|7|17|Every hand will go limp, and every knee will become as weak as water.
EZEK|7|18|They will put on sackcloth and be clothed with terror. Their faces will be covered with shame and their heads will be shaved.
EZEK|7|19|They will throw their silver into the streets, and their gold will be an unclean thing. Their silver and gold will not be able to save them in the day of the LORD 's wrath. They will not satisfy their hunger or fill their stomachs with it, for it has made them stumble into sin.
EZEK|7|20|They were proud of their beautiful jewelry and used it to make their detestable idols and vile images. Therefore I will turn these into an unclean thing for them.
EZEK|7|21|I will hand it all over as plunder to foreigners and as loot to the wicked of the earth, and they will defile it.
EZEK|7|22|I will turn my face away from them, and they will desecrate my treasured place; robbers will enter it and desecrate it.
EZEK|7|23|"Prepare chains, because the land is full of bloodshed and the city is full of violence.
EZEK|7|24|I will bring the most wicked of the nations to take possession of their houses; I will put an end to the pride of the mighty, and their sanctuaries will be desecrated.
EZEK|7|25|When terror comes, they will seek peace, but there will be none.
EZEK|7|26|Calamity upon calamity will come, and rumor upon rumor. They will try to get a vision from the prophet; the teaching of the law by the priest will be lost, as will the counsel of the elders.
EZEK|7|27|The king will mourn, the prince will be clothed with despair, and the hands of the people of the land will tremble. I will deal with them according to their conduct, and by their own standards I will judge them. Then they will know that I am the LORD."
EZEK|8|1|In the sixth year, in the sixth month on the fifth day, while I was sitting in my house and the elders of Judah were sitting before me, the hand of the Sovereign LORD came upon me there.
EZEK|8|2|I looked, and I saw a figure like that of a man. From what appeared to be his waist down he was like fire, and from there up his appearance was as bright as glowing metal.
EZEK|8|3|He stretched out what looked like a hand and took me by the hair of my head. The Spirit lifted me up between earth and heaven and in visions of God he took me to Jerusalem, to the entrance to the north gate of the inner court, where the idol that provokes to jealousy stood.
EZEK|8|4|And there before me was the glory of the God of Israel, as in the vision I had seen in the plain.
EZEK|8|5|Then he said to me, "Son of man, look toward the north." So I looked, and in the entrance north of the gate of the altar I saw this idol of jealousy.
EZEK|8|6|And he said to me, "Son of man, do you see what they are doing-the utterly detestable things the house of Israel is doing here, things that will drive me far from my sanctuary? But you will see things that are even more detestable."
EZEK|8|7|Then he brought me to the entrance to the court. I looked, and I saw a hole in the wall.
EZEK|8|8|He said to me, "Son of man, now dig into the wall." So I dug into the wall and saw a doorway there.
EZEK|8|9|And he said to me, "Go in and see the wicked and detestable things they are doing here."
EZEK|8|10|So I went in and looked, and I saw portrayed all over the walls all kinds of crawling things and detestable animals and all the idols of the house of Israel.
EZEK|8|11|In front of them stood seventy elders of the house of Israel, and Jaazaniah son of Shaphan was standing among them. Each had a censer in his hand, and a fragrant cloud of incense was rising.
EZEK|8|12|He said to me, "Son of man, have you seen what the elders of the house of Israel are doing in the darkness, each at the shrine of his own idol? They say, 'The LORD does not see us; the LORD has forsaken the land.'"
EZEK|8|13|Again, he said, "You will see them doing things that are even more detestable."
EZEK|8|14|Then he brought me to the entrance to the north gate of the house of the LORD, and I saw women sitting there, mourning for Tammuz.
EZEK|8|15|He said to me, "Do you see this, son of man? You will see things that are even more detestable than this."
EZEK|8|16|He then brought me into the inner court of the house of the LORD, and there at the entrance to the temple, between the portico and the altar, were about twenty-five men. With their backs toward the temple of the LORD and their faces toward the east, they were bowing down to the sun in the east.
EZEK|8|17|He said to me, "Have you seen this, son of man? Is it a trivial matter for the house of Judah to do the detestable things they are doing here? Must they also fill the land with violence and continually provoke me to anger? Look at them putting the branch to their nose!
EZEK|8|18|Therefore I will deal with them in anger; I will not look on them with pity or spare them. Although they shout in my ears, I will not listen to them."
EZEK|9|1|Then I heard him call out in a loud voice, "Bring the guards of the city here, each with a weapon in his hand."
EZEK|9|2|And I saw six men coming from the direction of the upper gate, which faces north, each with a deadly weapon in his hand. With them was a man clothed in linen who had a writing kit at his side. They came in and stood beside the bronze altar.
EZEK|9|3|Now the glory of the God of Israel went up from above the cherubim, where it had been, and moved to the threshold of the temple. Then the LORD called to the man clothed in linen who had the writing kit at his side
EZEK|9|4|and said to him, "Go throughout the city of Jerusalem and put a mark on the foreheads of those who grieve and lament over all the detestable things that are done in it."
EZEK|9|5|As I listened, he said to the others, "Follow him through the city and kill, without showing pity or compassion.
EZEK|9|6|Slaughter old men, young men and maidens, women and children, but do not touch anyone who has the mark. Begin at my sanctuary." So they began with the elders who were in front of the temple.
EZEK|9|7|Then he said to them, "Defile the temple and fill the courts with the slain. Go!" So they went out and began killing throughout the city.
EZEK|9|8|While they were killing and I was left alone, I fell facedown, crying out, "Ah, Sovereign LORD! Are you going to destroy the entire remnant of Israel in this outpouring of your wrath on Jerusalem?"
EZEK|9|9|He answered me, "The sin of the house of Israel and Judah is exceedingly great; the land is full of bloodshed and the city is full of injustice. They say, 'The LORD has forsaken the land; the LORD does not see.'
EZEK|9|10|So I will not look on them with pity or spare them, but I will bring down on their own heads what they have done."
EZEK|9|11|Then the man in linen with the writing kit at his side brought back word, saying, "I have done as you commanded."
EZEK|10|1|I looked, and I saw the likeness of a throne of sapphire above the expanse that was over the heads of the cherubim.
EZEK|10|2|The LORD said to the man clothed in linen, "Go in among the wheels beneath the cherubim. Fill your hands with burning coals from among the cherubim and scatter them over the city." And as I watched, he went in.
EZEK|10|3|Now the cherubim were standing on the south side of the temple when the man went in, and a cloud filled the inner court.
EZEK|10|4|Then the glory of the LORD rose from above the cherubim and moved to the threshold of the temple. The cloud filled the temple, and the court was full of the radiance of the glory of the LORD.
EZEK|10|5|The sound of the wings of the cherubim could be heard as far away as the outer court, like the voice of God Almighty when he speaks.
EZEK|10|6|When the LORD commanded the man in linen, "Take fire from among the wheels, from among the cherubim," the man went in and stood beside a wheel.
EZEK|10|7|Then one of the cherubim reached out his hand to the fire that was among them. He took up some of it and put it into the hands of the man in linen, who took it and went out.
EZEK|10|8|(Under the wings of the cherubim could be seen what looked like the hands of a man.)
EZEK|10|9|I looked, and I saw beside the cherubim four wheels, one beside each of the cherubim; the wheels sparkled like chrysolite.
EZEK|10|10|As for their appearance, the four of them looked alike; each was like a wheel intersecting a wheel.
EZEK|10|11|As they moved, they would go in any one of the four directions the cherubim faced; the wheels did not turn about as the cherubim went. The cherubim went in whatever direction the head faced, without turning as they went.
EZEK|10|12|Their entire bodies, including their backs, their hands and their wings, were completely full of eyes, as were their four wheels.
EZEK|10|13|I heard the wheels being called "the whirling wheels."
EZEK|10|14|Each of the cherubim had four faces: One face was that of a cherub, the second the face of a man, the third the face of a lion, and the fourth the face of an eagle.
EZEK|10|15|Then the cherubim rose upward. These were the living creatures I had seen by the Kebar River.
EZEK|10|16|When the cherubim moved, the wheels beside them moved; and when the cherubim spread their wings to rise from the ground, the wheels did not leave their side.
EZEK|10|17|When the cherubim stood still, they also stood still; and when the cherubim rose, they rose with them, because the spirit of the living creatures was in them.
EZEK|10|18|Then the glory of the LORD departed from over the threshold of the temple and stopped above the cherubim.
EZEK|10|19|While I watched, the cherubim spread their wings and rose from the ground, and as they went, the wheels went with them. They stopped at the entrance to the east gate of the LORD 's house, and the glory of the God of Israel was above them.
EZEK|10|20|These were the living creatures I had seen beneath the God of Israel by the Kebar River, and I realized that they were cherubim.
EZEK|10|21|Each had four faces and four wings, and under their wings was what looked like the hands of a man.
EZEK|10|22|Their faces had the same appearance as those I had seen by the Kebar River. Each one went straight ahead.
EZEK|11|1|Then the Spirit lifted me up and brought me to the gate of the house of the LORD that faces east. There at the entrance to the gate were twenty-five men, and I saw among them Jaazaniah son of Azzur and Pelatiah son of Benaiah, leaders of the people.
EZEK|11|2|The LORD said to me, "Son of man, these are the men who are plotting evil and giving wicked advice in this city.
EZEK|11|3|They say, 'Will it not soon be time to build houses? This city is a cooking pot, and we are the meat.'
EZEK|11|4|Therefore prophesy against them; prophesy, son of man."
EZEK|11|5|Then the Spirit of the LORD came upon me, and he told me to say: "This is what the LORD says: That is what you are saying, O house of Israel, but I know what is going through your mind.
EZEK|11|6|You have killed many people in this city and filled its streets with the dead.
EZEK|11|7|"Therefore this is what the Sovereign LORD says: The bodies you have thrown there are the meat and this city is the pot, but I will drive you out of it.
EZEK|11|8|You fear the sword, and the sword is what I will bring against you, declares the Sovereign LORD.
EZEK|11|9|I will drive you out of the city and hand you over to foreigners and inflict punishment on you.
EZEK|11|10|You will fall by the sword, and I will execute judgment on you at the borders of Israel. Then you will know that I am the LORD.
EZEK|11|11|This city will not be a pot for you, nor will you be the meat in it; I will execute judgment on you at the borders of Israel.
EZEK|11|12|And you will know that I am the LORD, for you have not followed my decrees or kept my laws but have conformed to the standards of the nations around you."
EZEK|11|13|Now as I was prophesying, Pelatiah son of Benaiah died. Then I fell facedown and cried out in a loud voice, "Ah, Sovereign LORD! Will you completely destroy the remnant of Israel?"
EZEK|11|14|The word of the LORD came to me:
EZEK|11|15|"Son of man, your brothers-your brothers who are your blood relatives and the whole house of Israel-are those of whom the people of Jerusalem have said, 'They are far away from the LORD; this land was given to us as our possession.'
EZEK|11|16|"Therefore say: 'This is what the Sovereign LORD says: Although I sent them far away among the nations and scattered them among the countries, yet for a little while I have been a sanctuary for them in the countries where they have gone.'
EZEK|11|17|"Therefore say: 'This is what the Sovereign LORD says: I will gather you from the nations and bring you back from the countries where you have been scattered, and I will give you back the land of Israel again.'
EZEK|11|18|"They will return to it and remove all its vile images and detestable idols.
EZEK|11|19|I will give them an undivided heart and put a new spirit in them; I will remove from them their heart of stone and give them a heart of flesh.
EZEK|11|20|Then they will follow my decrees and be careful to keep my laws. They will be my people, and I will be their God.
EZEK|11|21|But as for those whose hearts are devoted to their vile images and detestable idols, I will bring down on their own heads what they have done, declares the Sovereign LORD."
EZEK|11|22|Then the cherubim, with the wheels beside them, spread their wings, and the glory of the God of Israel was above them.
EZEK|11|23|The glory of the LORD went up from within the city and stopped above the mountain east of it.
EZEK|11|24|The Spirit lifted me up and brought me to the exiles in Babylonia in the vision given by the Spirit of God. Then the vision I had seen went up from me,
EZEK|11|25|and I told the exiles everything the LORD had shown me.
EZEK|12|1|The word of the LORD came to me:
EZEK|12|2|"Son of man, you are living among a rebellious people. They have eyes to see but do not see and ears to hear but do not hear, for they are a rebellious people.
EZEK|12|3|"Therefore, son of man, pack your belongings for exile and in the daytime, as they watch, set out and go from where you are to another place. Perhaps they will understand, though they are a rebellious house.
EZEK|12|4|During the daytime, while they watch, bring out your belongings packed for exile. Then in the evening, while they are watching, go out like those who go into exile.
EZEK|12|5|While they watch, dig through the wall and take your belongings out through it.
EZEK|12|6|Put them on your shoulder as they are watching and carry them out at dusk. Cover your face so that you cannot see the land, for I have made you a sign to the house of Israel."
EZEK|12|7|So I did as I was commanded. During the day I brought out my things packed for exile. Then in the evening I dug through the wall with my hands. I took my belongings out at dusk, carrying them on my shoulders while they watched.
EZEK|12|8|In the morning the word of the LORD came to me:
EZEK|12|9|"Son of man, did not that rebellious house of Israel ask you, 'What are you doing?'
EZEK|12|10|"Say to them, 'This is what the Sovereign LORD says: This oracle concerns the prince in Jerusalem and the whole house of Israel who are there.'
EZEK|12|11|Say to them, 'I am a sign to you.'"As I have done, so it will be done to them. They will go into exile as captives.
EZEK|12|12|"The prince among them will put his things on his shoulder at dusk and leave, and a hole will be dug in the wall for him to go through. He will cover his face so that he cannot see the land.
EZEK|12|13|I will spread my net for him, and he will be caught in my snare; I will bring him to Babylonia, the land of the Chaldeans, but he will not see it, and there he will die.
EZEK|12|14|I will scatter to the winds all those around him-his staff and all his troops-and I will pursue them with drawn sword.
EZEK|12|15|"They will know that I am the LORD, when I disperse them among the nations and scatter them through the countries.
EZEK|12|16|But I will spare a few of them from the sword, famine and plague, so that in the nations where they go they may acknowledge all their detestable practices. Then they will know that I am the LORD."
EZEK|12|17|The word of the LORD came to me:
EZEK|12|18|"Son of man, tremble as you eat your food, and shudder in fear as you drink your water.
EZEK|12|19|Say to the people of the land: 'This is what the Sovereign LORD says about those living in Jerusalem and in the land of Israel: They will eat their food in anxiety and drink their water in despair, for their land will be stripped of everything in it because of the violence of all who live there.
EZEK|12|20|The inhabited towns will be laid waste and the land will be desolate. Then you will know that I am the LORD.'"
EZEK|12|21|The word of the LORD came to me:
EZEK|12|22|"Son of man, what is this proverb you have in the land of Israel: 'The days go by and every vision comes to nothing'?
EZEK|12|23|Say to them, 'This is what the Sovereign LORD says: I am going to put an end to this proverb, and they will no longer quote it in Israel.' Say to them, 'The days are near when every vision will be fulfilled.
EZEK|12|24|For there will be no more false visions or flattering divinations among the people of Israel.
EZEK|12|25|But I the LORD will speak what I will, and it shall be fulfilled without delay. For in your days, you rebellious house, I will fulfill whatever I say, declares the Sovereign LORD.'"
EZEK|12|26|The word of the LORD came to me:
EZEK|12|27|"Son of man, the house of Israel is saying, 'The vision he sees is for many years from now, and he prophesies about the distant future.'
EZEK|12|28|"Therefore say to them, 'This is what the Sovereign LORD says: None of my words will be delayed any longer; whatever I say will be fulfilled, declares the Sovereign LORD.'"
EZEK|13|1|The word of the LORD came to me:
EZEK|13|2|"Son of man, prophesy against the prophets of Israel who are now prophesying. Say to those who prophesy out of their own imagination: 'Hear the word of the LORD!
EZEK|13|3|This is what the Sovereign LORD says: Woe to the foolish prophets who follow their own spirit and have seen nothing!
EZEK|13|4|Your prophets, O Israel, are like jackals among ruins.
EZEK|13|5|You have not gone up to the breaks in the wall to repair it for the house of Israel so that it will stand firm in the battle on the day of the LORD.
EZEK|13|6|Their visions are false and their divinations a lie. They say, "The LORD declares," when the LORD has not sent them; yet they expect their words to be fulfilled.
EZEK|13|7|Have you not seen false visions and uttered lying divinations when you say, "The LORD declares," though I have not spoken?
EZEK|13|8|"'Therefore this is what the Sovereign LORD says: Because of your false words and lying visions, I am against you, declares the Sovereign LORD.
EZEK|13|9|My hand will be against the prophets who see false visions and utter lying divinations. They will not belong to the council of my people or be listed in the records of the house of Israel, nor will they enter the land of Israel. Then you will know that I am the Sovereign LORD.
EZEK|13|10|"'Because they lead my people astray, saying, "Peace," when there is no peace, and because, when a flimsy wall is built, they cover it with whitewash,
EZEK|13|11|therefore tell those who cover it with whitewash that it is going to fall. Rain will come in torrents, and I will send hailstones hurtling down, and violent winds will burst forth.
EZEK|13|12|When the wall collapses, will people not ask you, "Where is the whitewash you covered it with?"
EZEK|13|13|"'Therefore this is what the Sovereign LORD says: In my wrath I will unleash a violent wind, and in my anger hailstones and torrents of rain will fall with destructive fury.
EZEK|13|14|I will tear down the wall you have covered with whitewash and will level it to the ground so that its foundation will be laid bare. When it falls, you will be destroyed in it; and you will know that I am the LORD.
EZEK|13|15|So I will spend my wrath against the wall and against those who covered it with whitewash. I will say to you, "The wall is gone and so are those who whitewashed it,
EZEK|13|16|those prophets of Israel who prophesied to Jerusalem and saw visions of peace for her when there was no peace, declares the Sovereign LORD."'
EZEK|13|17|"Now, son of man, set your face against the daughters of your people who prophesy out of their own imagination. Prophesy against them
EZEK|13|18|and say, 'This is what the Sovereign LORD says: Woe to the women who sew magic charms on all their wrists and make veils of various lengths for their heads in order to ensnare people. Will you ensnare the lives of my people but preserve your own?
EZEK|13|19|You have profaned me among my people for a few handfuls of barley and scraps of bread. By lying to my people, who listen to lies, you have killed those who should not have died and have spared those who should not live.
EZEK|13|20|"'Therefore this is what the Sovereign LORD says: I am against your magic charms with which you ensnare people like birds and I will tear them from your arms; I will set free the people that you ensnare like birds.
EZEK|13|21|I will tear off your veils and save my people from your hands, and they will no longer fall prey to your power. Then you will know that I am the LORD.
EZEK|13|22|Because you disheartened the righteous with your lies, when I had brought them no grief, and because you encouraged the wicked not to turn from their evil ways and so save their lives,
EZEK|13|23|therefore you will no longer see false visions or practice divination. I will save my people from your hands. And then you will know that I am the LORD.'"
EZEK|14|1|Some of the elders of Israel came to me and sat down in front of me.
EZEK|14|2|Then the word of the LORD came to me:
EZEK|14|3|"Son of man, these men have set up idols in their hearts and put wicked stumbling blocks before their faces. Should I let them inquire of me at all?
EZEK|14|4|Therefore speak to them and tell them, 'This is what the Sovereign LORD says: When any Israelite sets up idols in his heart and puts a wicked stumbling block before his face and then goes to a prophet, I the LORD will answer him myself in keeping with his great idolatry.
EZEK|14|5|I will do this to recapture the hearts of the people of Israel, who have all deserted me for their idols.'
EZEK|14|6|"Therefore say to the house of Israel, 'This is what the Sovereign LORD says: Repent! Turn from your idols and renounce all your detestable practices!
EZEK|14|7|"'When any Israelite or any alien living in Israel separates himself from me and sets up idols in his heart and puts a wicked stumbling block before his face and then goes to a prophet to inquire of me, I the LORD will answer him myself.
EZEK|14|8|I will set my face against that man and make him an example and a byword. I will cut him off from my people. Then you will know that I am the LORD.
EZEK|14|9|"'And if the prophet is enticed to utter a prophecy, I the LORD have enticed that prophet, and I will stretch out my hand against him and destroy him from among my people Israel.
EZEK|14|10|They will bear their guilt-the prophet will be as guilty as the one who consults him.
EZEK|14|11|Then the people of Israel will no longer stray from me, nor will they defile themselves anymore with all their sins. They will be my people, and I will be their God, declares the Sovereign LORD.'"
EZEK|14|12|The word of the LORD came to me:
EZEK|14|13|"Son of man, if a country sins against me by being unfaithful and I stretch out my hand against it to cut off its food supply and send famine upon it and kill its men and their animals,
EZEK|14|14|even if these three men-Noah, Daniel and Job-were in it, they could save only themselves by their righteousness, declares the Sovereign LORD.
EZEK|14|15|"Or if I send wild beasts through that country and they leave it childless and it becomes desolate so that no one can pass through it because of the beasts,
EZEK|14|16|as surely as I live, declares the Sovereign LORD, even if these three men were in it, they could not save their own sons or daughters. They alone would be saved, but the land would be desolate.
EZEK|14|17|"Or if I bring a sword against that country and say, 'Let the sword pass throughout the land,' and I kill its men and their animals,
EZEK|14|18|as surely as I live, declares the Sovereign LORD, even if these three men were in it, they could not save their own sons or daughters. They alone would be saved.
EZEK|14|19|"Or if I send a plague into that land and pour out my wrath upon it through bloodshed, killing its men and their animals,
EZEK|14|20|as surely as I live, declares the Sovereign LORD, even if Noah, Daniel and Job were in it, they could save neither son nor daughter. They would save only themselves by their righteousness.
EZEK|14|21|"For this is what the Sovereign LORD says: How much worse will it be when I send against Jerusalem my four dreadful judgments-sword and famine and wild beasts and plague-to kill its men and their animals!
EZEK|14|22|Yet there will be some survivors-sons and daughters who will be brought out of it. They will come to you, and when you see their conduct and their actions, you will be consoled regarding the disaster I have brought upon Jerusalem-every disaster I have brought upon it.
EZEK|14|23|You will be consoled when you see their conduct and their actions, for you will know that I have done nothing in it without cause, declares the Sovereign LORD."
EZEK|15|1|The word of the LORD came to me:
EZEK|15|2|"Son of man, how is the wood of a vine better than that of a branch on any of the trees in the forest?
EZEK|15|3|Is wood ever taken from it to make anything useful? Do they make pegs from it to hang things on?
EZEK|15|4|And after it is thrown on the fire as fuel and the fire burns both ends and chars the middle, is it then useful for anything?
EZEK|15|5|If it was not useful for anything when it was whole, how much less can it be made into something useful when the fire has burned it and it is charred?
EZEK|15|6|"Therefore this is what the Sovereign LORD says: As I have given the wood of the vine among the trees of the forest as fuel for the fire, so will I treat the people living in Jerusalem.
EZEK|15|7|I will set my face against them. Although they have come out of the fire, the fire will yet consume them. And when I set my face against them, you will know that I am the LORD.
EZEK|15|8|I will make the land desolate because they have been unfaithful, declares the Sovereign LORD."
EZEK|16|1|The word of the LORD came to me:
EZEK|16|2|"Son of man, confront Jerusalem with her detestable practices
EZEK|16|3|and say, 'This is what the Sovereign LORD says to Jerusalem: Your ancestry and birth were in the land of the Canaanites; your father was an Amorite and your mother a Hittite.
EZEK|16|4|On the day you were born your cord was not cut, nor were you washed with water to make you clean, nor were you rubbed with salt or wrapped in cloths.
EZEK|16|5|No one looked on you with pity or had compassion enough to do any of these things for you. Rather, you were thrown out into the open field, for on the day you were born you were despised.
EZEK|16|6|"'Then I passed by and saw you kicking about in your blood, and as you lay there in your blood I said to you, "Live!"
EZEK|16|7|I made you grow like a plant of the field. You grew up and developed and became the most beautiful of jewels. Your breasts were formed and your hair grew, you who were naked and bare.
EZEK|16|8|"'Later I passed by, and when I looked at you and saw that you were old enough for love, I spread the corner of my garment over you and covered your nakedness. I gave you my solemn oath and entered into a covenant with you, declares the Sovereign LORD, and you became mine.
EZEK|16|9|"'I bathed you with water and washed the blood from you and put ointments on you.
EZEK|16|10|I clothed you with an embroidered dress and put leather sandals on you. I dressed you in fine linen and covered you with costly garments.
EZEK|16|11|I adorned you with jewelry: I put bracelets on your arms and a necklace around your neck,
EZEK|16|12|and I put a ring on your nose, earrings on your ears and a beautiful crown on your head.
EZEK|16|13|So you were adorned with gold and silver; your clothes were of fine linen and costly fabric and embroidered cloth. Your food was fine flour, honey and olive oil. You became very beautiful and rose to be a queen.
EZEK|16|14|And your fame spread among the nations on account of your beauty, because the splendor I had given you made your beauty perfect, declares the Sovereign LORD.
EZEK|16|15|"'But you trusted in your beauty and used your fame to become a prostitute. You lavished your favors on anyone who passed by and your beauty became his.
EZEK|16|16|You took some of your garments to make gaudy high places, where you carried on your prostitution. Such things should not happen, nor should they ever occur.
EZEK|16|17|You also took the fine jewelry I gave you, the jewelry made of my gold and silver, and you made for yourself male idols and engaged in prostitution with them.
EZEK|16|18|And you took your embroidered clothes to put on them, and you offered my oil and incense before them.
EZEK|16|19|Also the food I provided for you-the fine flour, olive oil and honey I gave you to eat-you offered as fragrant incense before them. That is what happened, declares the Sovereign LORD.
EZEK|16|20|"'And you took your sons and daughters whom you bore to me and sacrificed them as food to the idols. Was your prostitution not enough?
EZEK|16|21|You slaughtered my children and sacrificed them to the idols.
EZEK|16|22|In all your detestable practices and your prostitution you did not remember the days of your youth, when you were naked and bare, kicking about in your blood.
EZEK|16|23|"'Woe! Woe to you, declares the Sovereign LORD. In addition to all your other wickedness,
EZEK|16|24|you built a mound for yourself and made a lofty shrine in every public square.
EZEK|16|25|At the head of every street you built your lofty shrines and degraded your beauty, offering your body with increasing promiscuity to anyone who passed by.
EZEK|16|26|You engaged in prostitution with the Egyptians, your lustful neighbors, and provoked me to anger with your increasing promiscuity.
EZEK|16|27|So I stretched out my hand against you and reduced your territory; I gave you over to the greed of your enemies, the daughters of the Philistines, who were shocked by your lewd conduct.
EZEK|16|28|You engaged in prostitution with the Assyrians too, because you were insatiable; and even after that, you still were not satisfied.
EZEK|16|29|Then you increased your promiscuity to include Babylonia, a land of merchants, but even with this you were not satisfied.
EZEK|16|30|"'How weak-willed you are, declares the Sovereign LORD, when you do all these things, acting like a brazen prostitute!
EZEK|16|31|When you built your mounds at the head of every street and made your lofty shrines in every public square, you were unlike a prostitute, because you scorned payment.
EZEK|16|32|"'You adulterous wife! You prefer strangers to your own husband!
EZEK|16|33|Every prostitute receives a fee, but you give gifts to all your lovers, bribing them to come to you from everywhere for your illicit favors.
EZEK|16|34|So in your prostitution you are the opposite of others; no one runs after you for your favors. You are the very opposite, for you give payment and none is given to you.
EZEK|16|35|"'Therefore, you prostitute, hear the word of the LORD!
EZEK|16|36|This is what the Sovereign LORD says: Because you poured out your wealth and exposed your nakedness in your promiscuity with your lovers, and because of all your detestable idols, and because you gave them your children's blood,
EZEK|16|37|therefore I am going to gather all your lovers, with whom you found pleasure, those you loved as well as those you hated. I will gather them against you from all around and will strip you in front of them, and they will see all your nakedness.
EZEK|16|38|I will sentence you to the punishment of women who commit adultery and who shed blood; I will bring upon you the blood vengeance of my wrath and jealous anger.
EZEK|16|39|Then I will hand you over to your lovers, and they will tear down your mounds and destroy your lofty shrines. They will strip you of your clothes and take your fine jewelry and leave you naked and bare.
EZEK|16|40|They will bring a mob against you, who will stone you and hack you to pieces with their swords.
EZEK|16|41|They will burn down your houses and inflict punishment on you in the sight of many women. I will put a stop to your prostitution, and you will no longer pay your lovers.
EZEK|16|42|Then my wrath against you will subside and my jealous anger will turn away from you; I will be calm and no longer angry.
EZEK|16|43|"'Because you did not remember the days of your youth but enraged me with all these things, I will surely bring down on your head what you have done, declares the Sovereign LORD. Did you not add lewdness to all your other detestable practices?
EZEK|16|44|"'Everyone who quotes proverbs will quote this proverb about you: "Like mother, like daughter."
EZEK|16|45|You are a true daughter of your mother, who despised her husband and her children; and you are a true sister of your sisters, who despised their husbands and their children. Your mother was a Hittite and your father an Amorite.
EZEK|16|46|Your older sister was Samaria, who lived to the north of you with her daughters; and your younger sister, who lived to the south of you with her daughters, was Sodom.
EZEK|16|47|You not only walked in their ways and copied their detestable practices, but in all your ways you soon became more depraved than they.
EZEK|16|48|As surely as I live, declares the Sovereign LORD, your sister Sodom and her daughters never did what you and your daughters have done.
EZEK|16|49|"'Now this was the sin of your sister Sodom: She and her daughters were arrogant, overfed and unconcerned; they did not help the poor and needy.
EZEK|16|50|They were haughty and did detestable things before me. Therefore I did away with them as you have seen.
EZEK|16|51|Samaria did not commit half the sins you did. You have done more detestable things than they, and have made your sisters seem righteous by all these things you have done.
EZEK|16|52|Bear your disgrace, for you have furnished some justification for your sisters. Because your sins were more vile than theirs, they appear more righteous than you. So then, be ashamed and bear your disgrace, for you have made your sisters appear righteous.
EZEK|16|53|"'However, I will restore the fortunes of Sodom and her daughters and of Samaria and her daughters, and your fortunes along with them,
EZEK|16|54|so that you may bear your disgrace and be ashamed of all you have done in giving them comfort.
EZEK|16|55|And your sisters, Sodom with her daughters and Samaria with her daughters, will return to what they were before; and you and your daughters will return to what you were before.
EZEK|16|56|You would not even mention your sister Sodom in the day of your pride,
EZEK|16|57|before your wickedness was uncovered. Even so, you are now scorned by the daughters of Edom and all her neighbors and the daughters of the Philistines-all those around you who despise you.
EZEK|16|58|You will bear the consequences of your lewdness and your detestable practices, declares the LORD.
EZEK|16|59|"'This is what the Sovereign LORD says: I will deal with you as you deserve, because you have despised my oath by breaking the covenant.
EZEK|16|60|Yet I will remember the covenant I made with you in the days of your youth, and I will establish an everlasting covenant with you.
EZEK|16|61|Then you will remember your ways and be ashamed when you receive your sisters, both those who are older than you and those who are younger. I will give them to you as daughters, but not on the basis of my covenant with you.
EZEK|16|62|So I will establish my covenant with you, and you will know that I am the LORD.
EZEK|16|63|Then, when I make atonement for you for all you have done, you will remember and be ashamed and never again open your mouth because of your humiliation, declares the Sovereign LORD.'"
EZEK|17|1|The word of the LORD came to me:
EZEK|17|2|"Son of man, set forth an allegory and tell the house of Israel a parable.
EZEK|17|3|Say to them, 'This is what the Sovereign LORD says: A great eagle with powerful wings, long feathers and full plumage of varied colors came to Lebanon. Taking hold of the top of a cedar,
EZEK|17|4|he broke off its topmost shoot and carried it away to a land of merchants, where he planted it in a city of traders.
EZEK|17|5|"'He took some of the seed of your land and put it in fertile soil. He planted it like a willow by abundant water,
EZEK|17|6|and it sprouted and became a low, spreading vine. Its branches turned toward him, but its roots remained under it. So it became a vine and produced branches and put out leafy boughs.
EZEK|17|7|"'But there was another great eagle with powerful wings and full plumage. The vine now sent out its roots toward him from the plot where it was planted and stretched out its branches to him for water.
EZEK|17|8|It had been planted in good soil by abundant water so that it would produce branches, bear fruit and become a splendid vine.'
EZEK|17|9|"Say to them, 'This is what the Sovereign LORD says: Will it thrive? Will it not be uprooted and stripped of its fruit so that it withers? All its new growth will wither. It will not take a strong arm or many people to pull it up by the roots.
EZEK|17|10|Even if it is transplanted, will it thrive? Will it not wither completely when the east wind strikes it-wither away in the plot where it grew?'"
EZEK|17|11|Then the word of the LORD came to me:
EZEK|17|12|"Say to this rebellious house, 'Do you not know what these things mean?' Say to them: 'The king of Babylon went to Jerusalem and carried off her king and her nobles, bringing them back with him to Babylon.
EZEK|17|13|Then he took a member of the royal family and made a treaty with him, putting him under oath. He also carried away the leading men of the land,
EZEK|17|14|so that the kingdom would be brought low, unable to rise again, surviving only by keeping his treaty.
EZEK|17|15|But the king rebelled against him by sending his envoys to Egypt to get horses and a large army. Will he succeed? Will he who does such things escape? Will he break the treaty and yet escape?
EZEK|17|16|"'As surely as I live, declares the Sovereign LORD, he shall die in Babylon, in the land of the king who put him on the throne, whose oath he despised and whose treaty he broke.
EZEK|17|17|Pharaoh with his mighty army and great horde will be of no help to him in war, when ramps are built and siege works erected to destroy many lives.
EZEK|17|18|He despised the oath by breaking the covenant. Because he had given his hand in pledge and yet did all these things, he shall not escape.
EZEK|17|19|"'Therefore this is what the Sovereign LORD says: As surely as I live, I will bring down on his head my oath that he despised and my covenant that he broke.
EZEK|17|20|I will spread my net for him, and he will be caught in my snare. I will bring him to Babylon and execute judgment upon him there because he was unfaithful to me.
EZEK|17|21|All his fleeing troops will fall by the sword, and the survivors will be scattered to the winds. Then you will know that I the LORD have spoken.
EZEK|17|22|"'This is what the Sovereign LORD says: I myself will take a shoot from the very top of a cedar and plant it; I will break off a tender sprig from its topmost shoots and plant it on a high and lofty mountain.
EZEK|17|23|On the mountain heights of Israel I will plant it; it will produce branches and bear fruit and become a splendid cedar. Birds of every kind will nest in it; they will find shelter in the shade of its branches.
EZEK|17|24|All the trees of the field will know that I the LORD bring down the tall tree and make the low tree grow tall. I dry up the green tree and make the dry tree flourish. "'I the LORD have spoken, and I will do it.'"
EZEK|18|1|The word of the LORD came to me:
EZEK|18|2|"What do you people mean by quoting this proverb about the land of Israel: "'The fathers eat sour grapes, and the children's teeth are set on edge'?
EZEK|18|3|"As surely as I live, declares the Sovereign LORD, you will no longer quote this proverb in Israel.
EZEK|18|4|For every living soul belongs to me, the father as well as the son-both alike belong to me. The soul who sins is the one who will die.
EZEK|18|5|"Suppose there is a righteous man who does what is just and right.
EZEK|18|6|He does not eat at the mountain shrines or look to the idols of the house of Israel. He does not defile his neighbor's wife or lie with a woman during her period.
EZEK|18|7|He does not oppress anyone, but returns what he took in pledge for a loan. He does not commit robbery but gives his food to the hungry and provides clothing for the naked.
EZEK|18|8|He does not lend at usury or take excessive interest. He withholds his hand from doing wrong and judges fairly between man and man.
EZEK|18|9|He follows my decrees and faithfully keeps my laws. That man is righteous; he will surely live, declares the Sovereign LORD.
EZEK|18|10|"Suppose he has a violent son, who sheds blood or does any of these other things
EZEK|18|11|(though the father has done none of them): "He eats at the mountain shrines. He defiles his neighbor's wife.
EZEK|18|12|He oppresses the poor and needy. He commits robbery. He does not return what he took in pledge. He looks to the idols. He does detestable things.
EZEK|18|13|He lends at usury and takes excessive interest. Will such a man live? He will not! Because he has done all these detestable things, he will surely be put to death and his blood will be on his own head.
EZEK|18|14|"But suppose this son has a son who sees all the sins his father commits, and though he sees them, he does not do such things:
EZEK|18|15|"He does not eat at the mountain shrines or look to the idols of the house of Israel. He does not defile his neighbor's wife.
EZEK|18|16|He does not oppress anyone or require a pledge for a loan. He does not commit robbery but gives his food to the hungry and provides clothing for the naked.
EZEK|18|17|He withholds his hand from sin and takes no usury or excessive interest. He keeps my laws and follows my decrees. He will not die for his father's sin; he will surely live.
EZEK|18|18|But his father will die for his own sin, because he practiced extortion, robbed his brother and did what was wrong among his people.
EZEK|18|19|"Yet you ask, 'Why does the son not share the guilt of his father?' Since the son has done what is just and right and has been careful to keep all my decrees, he will surely live.
EZEK|18|20|The soul who sins is the one who will die. The son will not share the guilt of the father, nor will the father share the guilt of the son. The righteousness of the righteous man will be credited to him, and the wickedness of the wicked will be charged against him.
EZEK|18|21|"But if a wicked man turns away from all the sins he has committed and keeps all my decrees and does what is just and right, he will surely live; he will not die.
EZEK|18|22|None of the offenses he has committed will be remembered against him. Because of the righteous things he has done, he will live.
EZEK|18|23|Do I take any pleasure in the death of the wicked? declares the Sovereign LORD. Rather, am I not pleased when they turn from their ways and live?
EZEK|18|24|"But if a righteous man turns from his righteousness and commits sin and does the same detestable things the wicked man does, will he live? None of the righteous things he has done will be remembered. Because of the unfaithfulness he is guilty of and because of the sins he has committed, he will die.
EZEK|18|25|"Yet you say, 'The way of the Lord is not just.' Hear, O house of Israel: Is my way unjust? Is it not your ways that are unjust?
EZEK|18|26|If a righteous man turns from his righteousness and commits sin, he will die for it; because of the sin he has committed he will die.
EZEK|18|27|But if a wicked man turns away from the wickedness he has committed and does what is just and right, he will save his life.
EZEK|18|28|Because he considers all the offenses he has committed and turns away from them, he will surely live; he will not die.
EZEK|18|29|Yet the house of Israel says, 'The way of the Lord is not just.' Are my ways unjust, O house of Israel? Is it not your ways that are unjust?
EZEK|18|30|"Therefore, O house of Israel, I will judge you, each one according to his ways, declares the Sovereign LORD. Repent! Turn away from all your offenses; then sin will not be your downfall.
EZEK|18|31|Rid yourselves of all the offenses you have committed, and get a new heart and a new spirit. Why will you die, O house of Israel?
EZEK|18|32|For I take no pleasure in the death of anyone, declares the Sovereign LORD. Repent and live!
EZEK|19|1|"Take up a lament concerning the princes of Israel
EZEK|19|2|and say: "'What a lioness was your mother among the lions! She lay down among the young lions and reared her cubs.
EZEK|19|3|She brought up one of her cubs, and he became a strong lion. He learned to tear the prey and he devoured men.
EZEK|19|4|The nations heard about him, and he was trapped in their pit. They led him with hooks to the land of Egypt.
EZEK|19|5|"'When she saw her hope unfulfilled, her expectation gone, she took another of her cubs and made him a strong lion.
EZEK|19|6|He prowled among the lions, for he was now a strong lion. He learned to tear the prey and he devoured men.
EZEK|19|7|He broke down their strongholds and devastated their towns. The land and all who were in it were terrified by his roaring.
EZEK|19|8|Then the nations came against him, those from regions round about. They spread their net for him, and he was trapped in their pit.
EZEK|19|9|With hooks they pulled him into a cage and brought him to the king of Babylon. They put him in prison, so his roar was heard no longer on the mountains of Israel.
EZEK|19|10|"'Your mother was like a vine in your vineyard planted by the water; it was fruitful and full of branches because of abundant water.
EZEK|19|11|Its branches were strong, fit for a ruler's scepter. It towered high above the thick foliage, conspicuous for its height and for its many branches.
EZEK|19|12|But it was uprooted in fury and thrown to the ground. The east wind made it shrivel, it was stripped of its fruit; its strong branches withered and fire consumed them.
EZEK|19|13|Now it is planted in the desert, in a dry and thirsty land.
EZEK|19|14|Fire spread from one of its main branches and consumed its fruit. No strong branch is left on it fit for a ruler's scepter.' This is a lament and is to be used as a lament."
EZEK|20|1|In the seventh year, in the fifth month on the tenth day, some of the elders of Israel came to inquire of the LORD, and they sat down in front of me.
EZEK|20|2|Then the word of the LORD came to me:
EZEK|20|3|"Son of man, speak to the elders of Israel and say to them, 'This is what the Sovereign LORD says: Have you come to inquire of me? As surely as I live, I will not let you inquire of me, declares the Sovereign LORD.'
EZEK|20|4|"Will you judge them? Will you judge them, son of man? Then confront them with the detestable practices of their fathers
EZEK|20|5|and say to them: 'This is what the Sovereign LORD says: On the day I chose Israel, I swore with uplifted hand to the descendants of the house of Jacob and revealed myself to them in Egypt. With uplifted hand I said to them, "I am the LORD your God."
EZEK|20|6|On that day I swore to them that I would bring them out of Egypt into a land I had searched out for them, a land flowing with milk and honey, the most beautiful of all lands.
EZEK|20|7|And I said to them, "Each of you, get rid of the vile images you have set your eyes on, and do not defile yourselves with the idols of Egypt. I am the LORD your God."
EZEK|20|8|"'But they rebelled against me and would not listen to me; they did not get rid of the vile images they had set their eyes on, nor did they forsake the idols of Egypt. So I said I would pour out my wrath on them and spend my anger against them in Egypt.
EZEK|20|9|But for the sake of my name I did what would keep it from being profaned in the eyes of the nations they lived among and in whose sight I had revealed myself to the Israelites by bringing them out of Egypt.
EZEK|20|10|Therefore I led them out of Egypt and brought them into the desert.
EZEK|20|11|I gave them my decrees and made known to them my laws, for the man who obeys them will live by them.
EZEK|20|12|Also I gave them my Sabbaths as a sign between us, so they would know that I the LORD made them holy.
EZEK|20|13|"'Yet the people of Israel rebelled against me in the desert. They did not follow my decrees but rejected my laws-although the man who obeys them will live by them-and they utterly desecrated my Sabbaths. So I said I would pour out my wrath on them and destroy them in the desert.
EZEK|20|14|But for the sake of my name I did what would keep it from being profaned in the eyes of the nations in whose sight I had brought them out.
EZEK|20|15|Also with uplifted hand I swore to them in the desert that I would not bring them into the land I had given them-a land flowing with milk and honey, most beautiful of all lands-
EZEK|20|16|because they rejected my laws and did not follow my decrees and desecrated my Sabbaths. For their hearts were devoted to their idols.
EZEK|20|17|Yet I looked on them with pity and did not destroy them or put an end to them in the desert.
EZEK|20|18|I said to their children in the desert, "Do not follow the statutes of your fathers or keep their laws or defile yourselves with their idols.
EZEK|20|19|I am the LORD your God; follow my decrees and be careful to keep my laws.
EZEK|20|20|Keep my Sabbaths holy, that they may be a sign between us. Then you will know that I am the LORD your God."
EZEK|20|21|"'But the children rebelled against me: They did not follow my decrees, they were not careful to keep my laws-although the man who obeys them will live by them-and they desecrated my Sabbaths. So I said I would pour out my wrath on them and spend my anger against them in the desert.
EZEK|20|22|But I withheld my hand, and for the sake of my name I did what would keep it from being profaned in the eyes of the nations in whose sight I had brought them out.
EZEK|20|23|Also with uplifted hand I swore to them in the desert that I would disperse them among the nations and scatter them through the countries,
EZEK|20|24|because they had not obeyed my laws but had rejected my decrees and desecrated my Sabbaths, and their eyes lusted after their fathers' idols.
EZEK|20|25|I also gave them over to statutes that were not good and laws they could not live by;
EZEK|20|26|I let them become defiled through their gifts-the sacrifice of every firstborn -that I might fill them with horror so they would know that I am the LORD.'
EZEK|20|27|"Therefore, son of man, speak to the people of Israel and say to them, 'This is what the Sovereign LORD says: In this also your fathers blasphemed me by forsaking me:
EZEK|20|28|When I brought them into the land I had sworn to give them and they saw any high hill or any leafy tree, there they offered their sacrifices, made offerings that provoked me to anger, presented their fragrant incense and poured out their drink offerings.
EZEK|20|29|Then I said to them: What is this high place you go to?'" (It is called Bamah to this day.)
EZEK|20|30|"Therefore say to the house of Israel: 'This is what the Sovereign LORD says: Will you defile yourselves the way your fathers did and lust after their vile images?
EZEK|20|31|When you offer your gifts-the sacrifice of your sons in the fire-you continue to defile yourselves with all your idols to this day. Am I to let you inquire of me, O house of Israel? As surely as I live, declares the Sovereign LORD, I will not let you inquire of me.
EZEK|20|32|"'You say, "We want to be like the nations, like the peoples of the world, who serve wood and stone." But what you have in mind will never happen.
EZEK|20|33|As surely as I live, declares the Sovereign LORD, I will rule over you with a mighty hand and an outstretched arm and with outpoured wrath.
EZEK|20|34|I will bring you from the nations and gather you from the countries where you have been scattered-with a mighty hand and an outstretched arm and with outpoured wrath.
EZEK|20|35|I will bring you into the desert of the nations and there, face to face, I will execute judgment upon you.
EZEK|20|36|As I judged your fathers in the desert of the land of Egypt, so I will judge you, declares the Sovereign LORD.
EZEK|20|37|I will take note of you as you pass under my rod, and I will bring you into the bond of the covenant.
EZEK|20|38|I will purge you of those who revolt and rebel against me. Although I will bring them out of the land where they are living, yet they will not enter the land of Israel. Then you will know that I am the LORD.
EZEK|20|39|"'As for you, O house of Israel, this is what the Sovereign LORD says: Go and serve your idols, every one of you! But afterward you will surely listen to me and no longer profane my holy name with your gifts and idols.
EZEK|20|40|For on my holy mountain, the high mountain of Israel, declares the Sovereign LORD, there in the land the entire house of Israel will serve me, and there I will accept them. There I will require your offerings and your choice gifts, along with all your holy sacrifices.
EZEK|20|41|I will accept you as fragrant incense when I bring you out from the nations and gather you from the countries where you have been scattered, and I will show myself holy among you in the sight of the nations.
EZEK|20|42|Then you will know that I am the LORD, when I bring you into the land of Israel, the land I had sworn with uplifted hand to give to your fathers.
EZEK|20|43|There you will remember your conduct and all the actions by which you have defiled yourselves, and you will loathe yourselves for all the evil you have done.
EZEK|20|44|You will know that I am the LORD, when I deal with you for my name's sake and not according to your evil ways and your corrupt practices, O house of Israel, declares the Sovereign LORD.'"
EZEK|20|45|The word of the LORD came to me:
EZEK|20|46|"Son of man, set your face toward the south; preach against the south and prophesy against the forest of the southland.
EZEK|20|47|Say to the southern forest: 'Hear the word of the LORD. This is what the Sovereign LORD says: I am about to set fire to you, and it will consume all your trees, both green and dry. The blazing flame will not be quenched, and every face from south to north will be scorched by it.
EZEK|20|48|Everyone will see that I the LORD have kindled it; it will not be quenched.'"
EZEK|20|49|Then I said, "Ah, Sovereign LORD! They are saying of me, 'Isn't he just telling parables?'"
EZEK|21|1|The word of the LORD came to me:
EZEK|21|2|"Son of man, set your face against Jerusalem and preach against the sanctuary. Prophesy against the land of Israel
EZEK|21|3|and say to her: 'This is what the LORD says: I am against you. I will draw my sword from its scabbard and cut off from you both the righteous and the wicked.
EZEK|21|4|Because I am going to cut off the righteous and the wicked, my sword will be unsheathed against everyone from south to north.
EZEK|21|5|Then all people will know that I the LORD have drawn my sword from its scabbard; it will not return again.'
EZEK|21|6|"Therefore groan, son of man! Groan before them with broken heart and bitter grief.
EZEK|21|7|And when they ask you, 'Why are you groaning?' you shall say, 'Because of the news that is coming. Every heart will melt and every hand go limp; every spirit will become faint and every knee become as weak as water.' It is coming! It will surely take place, declares the Sovereign LORD."
EZEK|21|8|The word of the LORD came to me:
EZEK|21|9|"Son of man, prophesy and say, 'This is what the Lord says: "'A sword, a sword, sharpened and polished-
EZEK|21|10|sharpened for the slaughter, polished to flash like lightning! "'Shall we rejoice in the scepter of my son Judah? The sword despises every such stick.
EZEK|21|11|"'The sword is appointed to be polished, to be grasped with the hand; it is sharpened and polished, made ready for the hand of the slayer.
EZEK|21|12|Cry out and wail, son of man, for it is against my people; it is against all the princes of Israel. They are thrown to the sword along with my people. Therefore beat your breast.
EZEK|21|13|"'Testing will surely come. And what if the scepter of Judah, which the sword despises, does not continue? declares the Sovereign LORD.'
EZEK|21|14|"So then, son of man, prophesy and strike your hands together. Let the sword strike twice, even three times. It is a sword for slaughter- a sword for great slaughter, closing in on them from every side.
EZEK|21|15|So that hearts may melt and the fallen be many, I have stationed the sword for slaughter at all their gates. Oh! It is made to flash like lightning, it is grasped for slaughter.
EZEK|21|16|O sword, slash to the right, then to the left, wherever your blade is turned.
EZEK|21|17|I too will strike my hands together, and my wrath will subside. I the LORD have spoken."
EZEK|21|18|The word of the LORD came to me:
EZEK|21|19|"Son of man, mark out two roads for the sword of the king of Babylon to take, both starting from the same country. Make a signpost where the road branches off to the city.
EZEK|21|20|Mark out one road for the sword to come against Rabbah of the Ammonites and another against Judah and fortified Jerusalem.
EZEK|21|21|For the king of Babylon will stop at the fork in the road, at the junction of the two roads, to seek an omen: He will cast lots with arrows, he will consult his idols, he will examine the liver.
EZEK|21|22|Into his right hand will come the lot for Jerusalem, where he is to set up battering rams, to give the command to slaughter, to sound the battle cry, to set battering rams against the gates, to build a ramp and to erect siege works.
EZEK|21|23|It will seem like a false omen to those who have sworn allegiance to him, but he will remind them of their guilt and take them captive.
EZEK|21|24|"Therefore this is what the Sovereign LORD says: 'Because you people have brought to mind your guilt by your open rebellion, revealing your sins in all that you do-because you have done this, you will be taken captive.
EZEK|21|25|"'O profane and wicked prince of Israel, whose day has come, whose time of punishment has reached its climax,
EZEK|21|26|this is what the Sovereign LORD says: Take off the turban, remove the crown. It will not be as it was: The lowly will be exalted and the exalted will be brought low.
EZEK|21|27|A ruin! A ruin! I will make it a ruin! It will not be restored until he comes to whom it rightfully belongs; to him I will give it.'
EZEK|21|28|"And you, son of man, prophesy and say, 'This is what the Sovereign LORD says about the Ammonites and their insults: "'A sword, a sword, drawn for the slaughter, polished to consume and to flash like lightning!
EZEK|21|29|Despite false visions concerning you and lying divinations about you, it will be laid on the necks of the wicked who are to be slain, whose day has come, whose time of punishment has reached its climax.
EZEK|21|30|Return the sword to its scabbard. In the place where you were created, in the land of your ancestry, I will judge you.
EZEK|21|31|I will pour out my wrath upon you and breathe out my fiery anger against you; I will hand you over to brutal men, men skilled in destruction.
EZEK|21|32|You will be fuel for the fire, your blood will be shed in your land, you will be remembered no more; for I the LORD have spoken.'"
EZEK|22|1|The word of the LORD came to me:
EZEK|22|2|"Son of man, will you judge her? Will you judge this city of bloodshed? Then confront her with all her detestable practices
EZEK|22|3|and say: 'This is what the Sovereign LORD says: O city that brings on herself doom by shedding blood in her midst and defiles herself by making idols,
EZEK|22|4|you have become guilty because of the blood you have shed and have become defiled by the idols you have made. You have brought your days to a close, and the end of your years has come. Therefore I will make you an object of scorn to the nations and a laughingstock to all the countries.
EZEK|22|5|Those who are near and those who are far away will mock you, O infamous city, full of turmoil.
EZEK|22|6|"'See how each of the princes of Israel who are in you uses his power to shed blood.
EZEK|22|7|In you they have treated father and mother with contempt; in you they have oppressed the alien and mistreated the fatherless and the widow.
EZEK|22|8|You have despised my holy things and desecrated my Sabbaths.
EZEK|22|9|In you are slanderous men bent on shedding blood; in you are those who eat at the mountain shrines and commit lewd acts.
EZEK|22|10|In you are those who dishonor their fathers' bed; in you are those who violate women during their period, when they are ceremonially unclean.
EZEK|22|11|In you one man commits a detestable offense with his neighbor's wife, another shamefully defiles his daughter-in-law, and another violates his sister, his own father's daughter.
EZEK|22|12|In you men accept bribes to shed blood; you take usury and excessive interest and make unjust gain from your neighbors by extortion. And you have forgotten me, declares the Sovereign LORD.
EZEK|22|13|"'I will surely strike my hands together at the unjust gain you have made and at the blood you have shed in your midst.
EZEK|22|14|Will your courage endure or your hands be strong in the day I deal with you? I the LORD have spoken, and I will do it.
EZEK|22|15|I will disperse you among the nations and scatter you through the countries; and I will put an end to your uncleanness.
EZEK|22|16|When you have been defiled in the eyes of the nations, you will know that I am the LORD.'"
EZEK|22|17|Then the word of the LORD came to me:
EZEK|22|18|"Son of man, the house of Israel has become dross to me; all of them are the copper, tin, iron and lead left inside a furnace. They are but the dross of silver.
EZEK|22|19|Therefore this is what the Sovereign LORD says: 'Because you have all become dross, I will gather you into Jerusalem.
EZEK|22|20|As men gather silver, copper, iron, lead and tin into a furnace to melt it with a fiery blast, so will I gather you in my anger and my wrath and put you inside the city and melt you.
EZEK|22|21|I will gather you and I will blow on you with my fiery wrath, and you will be melted inside her.
EZEK|22|22|As silver is melted in a furnace, so you will be melted inside her, and you will know that I the LORD have poured out my wrath upon you.'"
EZEK|22|23|Again the word of the LORD came to me:
EZEK|22|24|"Son of man, say to the land, 'You are a land that has had no rain or showers in the day of wrath.'
EZEK|22|25|There is a conspiracy of her princes within her like a roaring lion tearing its prey; they devour people, take treasures and precious things and make many widows within her.
EZEK|22|26|Her priests do violence to my law and profane my holy things; they do not distinguish between the holy and the common; they teach that there is no difference between the unclean and the clean; and they shut their eyes to the keeping of my Sabbaths, so that I am profaned among them.
EZEK|22|27|Her officials within her are like wolves tearing their prey; they shed blood and kill people to make unjust gain.
EZEK|22|28|Her prophets whitewash these deeds for them by false visions and lying divinations. They say, 'This is what the Sovereign LORD says'-when the LORD has not spoken.
EZEK|22|29|The people of the land practice extortion and commit robbery; they oppress the poor and needy and mistreat the alien, denying them justice.
EZEK|22|30|"I looked for a man among them who would build up the wall and stand before me in the gap on behalf of the land so I would not have to destroy it, but I found none.
EZEK|22|31|So I will pour out my wrath on them and consume them with my fiery anger, bringing down on their own heads all they have done, declares the Sovereign LORD."
EZEK|23|1|The word of the LORD came to me:
EZEK|23|2|"Son of man, there were two women, daughters of the same mother.
EZEK|23|3|They became prostitutes in Egypt, engaging in prostitution from their youth. In that land their breasts were fondled and their virgin bosoms caressed.
EZEK|23|4|The older was named Oholah, and her sister was Oholibah. They were mine and gave birth to sons and daughters. Oholah is Samaria, and Oholibah is Jerusalem.
EZEK|23|5|"Oholah engaged in prostitution while she was still mine; and she lusted after her lovers, the Assyrians-warriors
EZEK|23|6|clothed in blue, governors and commanders, all of them handsome young men, and mounted horsemen.
EZEK|23|7|She gave herself as a prostitute to all the elite of the Assyrians and defiled herself with all the idols of everyone she lusted after.
EZEK|23|8|She did not give up the prostitution she began in Egypt, when during her youth men slept with her, caressed her virgin bosom and poured out their lust upon her.
EZEK|23|9|"Therefore I handed her over to her lovers, the Assyrians, for whom she lusted.
EZEK|23|10|They stripped her naked, took away her sons and daughters and killed her with the sword. She became a byword among women, and punishment was inflicted on her.
EZEK|23|11|"Her sister Oholibah saw this, yet in her lust and prostitution she was more depraved than her sister.
EZEK|23|12|She too lusted after the Assyrians-governors and commanders, warriors in full dress, mounted horsemen, all handsome young men.
EZEK|23|13|I saw that she too defiled herself; both of them went the same way.
EZEK|23|14|"But she carried her prostitution still further. She saw men portrayed on a wall, figures of Chaldeans portrayed in red,
EZEK|23|15|with belts around their waists and flowing turbans on their heads; all of them looked like Babylonian chariot officers, natives of Chaldea.
EZEK|23|16|As soon as she saw them, she lusted after them and sent messengers to them in Chaldea.
EZEK|23|17|Then the Babylonians came to her, to the bed of love, and in their lust they defiled her. After she had been defiled by them, she turned away from them in disgust.
EZEK|23|18|When she carried on her prostitution openly and exposed her nakedness, I turned away from her in disgust, just as I had turned away from her sister.
EZEK|23|19|Yet she became more and more promiscuous as she recalled the days of her youth, when she was a prostitute in Egypt.
EZEK|23|20|There she lusted after her lovers, whose genitals were like those of donkeys and whose emission was like that of horses.
EZEK|23|21|So you longed for the lewdness of your youth, when in Egypt your bosom was caressed and your young breasts fondled.
EZEK|23|22|"Therefore, Oholibah, this is what the Sovereign LORD says: I will stir up your lovers against you, those you turned away from in disgust, and I will bring them against you from every side-
EZEK|23|23|the Babylonians and all the Chaldeans, the men of Pekod and Shoa and Koa, and all the Assyrians with them, handsome young men, all of them governors and commanders, chariot officers and men of high rank, all mounted on horses.
EZEK|23|24|They will come against you with weapons, chariots and wagons and with a throng of people; they will take up positions against you on every side with large and small shields and with helmets. I will turn you over to them for punishment, and they will punish you according to their standards.
EZEK|23|25|I will direct my jealous anger against you, and they will deal with you in fury. They will cut off your noses and your ears, and those of you who are left will fall by the sword. They will take away your sons and daughters, and those of you who are left will be consumed by fire.
EZEK|23|26|They will also strip you of your clothes and take your fine jewelry.
EZEK|23|27|So I will put a stop to the lewdness and prostitution you began in Egypt. You will not look on these things with longing or remember Egypt anymore.
EZEK|23|28|"For this is what the Sovereign LORD says: I am about to hand you over to those you hate, to those you turned away from in disgust.
EZEK|23|29|They will deal with you in hatred and take away everything you have worked for. They will leave you naked and bare, and the shame of your prostitution will be exposed. Your lewdness and promiscuity
EZEK|23|30|have brought this upon you, because you lusted after the nations and defiled yourself with their idols.
EZEK|23|31|You have gone the way of your sister; so I will put her cup into your hand.
EZEK|23|32|"This is what the Sovereign LORD says: "You will drink your sister's cup, a cup large and deep; it will bring scorn and derision, for it holds so much.
EZEK|23|33|You will be filled with drunkenness and sorrow, the cup of ruin and desolation, the cup of your sister Samaria.
EZEK|23|34|You will drink it and drain it dry; you will dash it to pieces and tear your breasts. I have spoken, declares the Sovereign LORD.
EZEK|23|35|"Therefore this is what the Sovereign LORD says: Since you have forgotten me and thrust me behind your back, you must bear the consequences of your lewdness and prostitution."
EZEK|23|36|The LORD said to me: "Son of man, will you judge Oholah and Oholibah? Then confront them with their detestable practices,
EZEK|23|37|for they have committed adultery and blood is on their hands. They committed adultery with their idols; they even sacrificed their children, whom they bore to me, as food for them.
EZEK|23|38|They have also done this to me: At that same time they defiled my sanctuary and desecrated my Sabbaths.
EZEK|23|39|On the very day they sacrificed their children to their idols, they entered my sanctuary and desecrated it. That is what they did in my house.
EZEK|23|40|"They even sent messengers for men who came from far away, and when they arrived you bathed yourself for them, painted your eyes and put on your jewelry.
EZEK|23|41|You sat on an elegant couch, with a table spread before it on which you had placed the incense and oil that belonged to me.
EZEK|23|42|"The noise of a carefree crowd was around her; Sabeans were brought from the desert along with men from the rabble, and they put bracelets on the arms of the woman and her sister and beautiful crowns on their heads.
EZEK|23|43|Then I said about the one worn out by adultery, 'Now let them use her as a prostitute, for that is all she is.'
EZEK|23|44|And they slept with her. As men sleep with a prostitute, so they slept with those lewd women, Oholah and Oholibah.
EZEK|23|45|But righteous men will sentence them to the punishment of women who commit adultery and shed blood, because they are adulterous and blood is on their hands.
EZEK|23|46|"This is what the Sovereign LORD says: Bring a mob against them and give them over to terror and plunder.
EZEK|23|47|The mob will stone them and cut them down with their swords; they will kill their sons and daughters and burn down their houses.
EZEK|23|48|"So I will put an end to lewdness in the land, that all women may take warning and not imitate you.
EZEK|23|49|You will suffer the penalty for your lewdness and bear the consequences of your sins of idolatry. Then you will know that I am the Sovereign LORD."
EZEK|24|1|In the ninth year, in the tenth month on the tenth day, the word of the LORD came to me:
EZEK|24|2|"Son of man, record this date, this very date, because the king of Babylon has laid siege to Jerusalem this very day.
EZEK|24|3|Tell this rebellious house a parable and say to them: 'This is what the Sovereign LORD says: "'Put on the cooking pot; put it on and pour water into it.
EZEK|24|4|Put into it the pieces of meat, all the choice pieces-the leg and the shoulder. Fill it with the best of these bones;
EZEK|24|5|take the pick of the flock. Pile wood beneath it for the bones; bring it to a boil and cook the bones in it.
EZEK|24|6|"'For this is what the Sovereign LORD says: "'Woe to the city of bloodshed, to the pot now encrusted, whose deposit will not go away! Empty it piece by piece without casting lots for them.
EZEK|24|7|"'For the blood she shed is in her midst: She poured it on the bare rock; she did not pour it on the ground, where the dust would cover it.
EZEK|24|8|To stir up wrath and take revenge I put her blood on the bare rock, so that it would not be covered.
EZEK|24|9|"'Therefore this is what the Sovereign LORD says: "'Woe to the city of bloodshed! I, too, will pile the wood high.
EZEK|24|10|So heap on the wood and kindle the fire. Cook the meat well, mixing in the spices; and let the bones be charred.
EZEK|24|11|Then set the empty pot on the coals till it becomes hot and its copper glows so its impurities may be melted and its deposit burned away.
EZEK|24|12|It has frustrated all efforts; its heavy deposit has not been removed, not even by fire.
EZEK|24|13|"'Now your impurity is lewdness. Because I tried to cleanse you but you would not be cleansed from your impurity, you will not be clean again until my wrath against you has subsided.
EZEK|24|14|"'I the LORD have spoken. The time has come for me to act. I will not hold back; I will not have pity, nor will I relent. You will be judged according to your conduct and your actions, declares the Sovereign LORD.'"
EZEK|24|15|The word of the LORD came to me:
EZEK|24|16|"Son of man, with one blow I am about to take away from you the delight of your eyes. Yet do not lament or weep or shed any tears.
EZEK|24|17|Groan quietly; do not mourn for the dead. Keep your turban fastened and your sandals on your feet; do not cover the lower part of your face or eat the customary food of mourners."
EZEK|24|18|So I spoke to the people in the morning, and in the evening my wife died. The next morning I did as I had been commanded.
EZEK|24|19|Then the people asked me, "Won't you tell us what these things have to do with us?"
EZEK|24|20|So I said to them, "The word of the LORD came to me:
EZEK|24|21|Say to the house of Israel, 'This is what the Sovereign LORD says: I am about to desecrate my sanctuary-the stronghold in which you take pride, the delight of your eyes, the object of your affection. The sons and daughters you left behind will fall by the sword.
EZEK|24|22|And you will do as I have done. You will not cover the lower part of your face or eat the customary food of mourners.
EZEK|24|23|You will keep your turbans on your heads and your sandals on your feet. You will not mourn or weep but will waste away because of your sins and groan among yourselves.
EZEK|24|24|Ezekiel will be a sign to you; you will do just as he has done. When this happens, you will know that I am the Sovereign LORD.'
EZEK|24|25|"And you, son of man, on the day I take away their stronghold, their joy and glory, the delight of their eyes, their heart's desire, and their sons and daughters as well-
EZEK|24|26|on that day a fugitive will come to tell you the news.
EZEK|24|27|At that time your mouth will be opened; you will speak with him and will no longer be silent. So you will be a sign to them, and they will know that I am the LORD."
EZEK|25|1|The word of the LORD came to me:
EZEK|25|2|"Son of man, set your face against the Ammonites and prophesy against them.
EZEK|25|3|Say to them, 'Hear the word of the Sovereign LORD. This is what the Sovereign LORD says: Because you said "Aha!" over my sanctuary when it was desecrated and over the land of Israel when it was laid waste and over the people of Judah when they went into exile,
EZEK|25|4|therefore I am going to give you to the people of the East as a possession. They will set up their camps and pitch their tents among you; they will eat your fruit and drink your milk.
EZEK|25|5|I will turn Rabbah into a pasture for camels and Ammon into a resting place for sheep. Then you will know that I am the LORD.
EZEK|25|6|For this is what the Sovereign LORD says: Because you have clapped your hands and stamped your feet, rejoicing with all the malice of your heart against the land of Israel,
EZEK|25|7|therefore I will stretch out my hand against you and give you as plunder to the nations. I will cut you off from the nations and exterminate you from the countries. I will destroy you, and you will know that I am the LORD.'"
EZEK|25|8|"This is what the Sovereign LORD says: 'Because Moab and Seir said, "Look, the house of Judah has become like all the other nations,"
EZEK|25|9|therefore I will expose the flank of Moab, beginning at its frontier towns-Beth Jeshimoth, Baal Meon and Kiriathaim-the glory of that land.
EZEK|25|10|I will give Moab along with the Ammonites to the people of the East as a possession, so that the Ammonites will not be remembered among the nations;
EZEK|25|11|and I will inflict punishment on Moab. Then they will know that I am the LORD.'"
EZEK|25|12|"This is what the Sovereign LORD says: 'Because Edom took revenge on the house of Judah and became very guilty by doing so,
EZEK|25|13|therefore this is what the Sovereign LORD says: I will stretch out my hand against Edom and kill its men and their animals. I will lay it waste, and from Teman to Dedan they will fall by the sword.
EZEK|25|14|I will take vengeance on Edom by the hand of my people Israel, and they will deal with Edom in accordance with my anger and my wrath; they will know my vengeance, declares the Sovereign LORD.'"
EZEK|25|15|"This is what the Sovereign LORD says: 'Because the Philistines acted in vengeance and took revenge with malice in their hearts, and with ancient hostility sought to destroy Judah,
EZEK|25|16|therefore this is what the Sovereign LORD says: I am about to stretch out my hand against the Philistines, and I will cut off the Kerethites and destroy those remaining along the coast.
EZEK|25|17|I will carry out great vengeance on them and punish them in my wrath. Then they will know that I am the LORD, when I take vengeance on them.'"
EZEK|26|1|In the eleventh year, on the first day of the month, the word of the LORD came to me:
EZEK|26|2|"Son of man, because Tyre has said of Jerusalem, 'Aha! The gate to the nations is broken, and its doors have swung open to me; now that she lies in ruins I will prosper,'
EZEK|26|3|therefore this is what the Sovereign LORD says: I am against you, O Tyre, and I will bring many nations against you, like the sea casting up its waves.
EZEK|26|4|They will destroy the walls of Tyre and pull down her towers; I will scrape away her rubble and make her a bare rock.
EZEK|26|5|Out in the sea she will become a place to spread fishnets, for I have spoken, declares the Sovereign LORD. She will become plunder for the nations,
EZEK|26|6|and her settlements on the mainland will be ravaged by the sword. Then they will know that I am the LORD.
EZEK|26|7|"For this is what the Sovereign LORD says: From the north I am going to bring against Tyre Nebuchadnezzar king of Babylon, king of kings, with horses and chariots, with horsemen and a great army.
EZEK|26|8|He will ravage your settlements on the mainland with the sword; he will set up siege works against you, build a ramp up to your walls and raise his shields against you.
EZEK|26|9|He will direct the blows of his battering rams against your walls and demolish your towers with his weapons.
EZEK|26|10|His horses will be so many that they will cover you with dust. Your walls will tremble at the noise of the war horses, wagons and chariots when he enters your gates as men enter a city whose walls have been broken through.
EZEK|26|11|The hoofs of his horses will trample all your streets; he will kill your people with the sword, and your strong pillars will fall to the ground.
EZEK|26|12|They will plunder your wealth and loot your merchandise; they will break down your walls and demolish your fine houses and throw your stones, timber and rubble into the sea.
EZEK|26|13|I will put an end to your noisy songs, and the music of your harps will be heard no more.
EZEK|26|14|I will make you a bare rock, and you will become a place to spread fishnets. You will never be rebuilt, for I the LORD have spoken, declares the Sovereign LORD.
EZEK|26|15|"This is what the Sovereign LORD says to Tyre: Will not the coastlands tremble at the sound of your fall, when the wounded groan and the slaughter takes place in you?
EZEK|26|16|Then all the princes of the coast will step down from their thrones and lay aside their robes and take off their embroidered garments. Clothed with terror, they will sit on the ground, trembling every moment, appalled at you.
EZEK|26|17|Then they will take up a lament concerning you and say to you: "'How you are destroyed, O city of renown, peopled by men of the sea! You were a power on the seas, you and your citizens; you put your terror on all who lived there.
EZEK|26|18|Now the coastlands tremble on the day of your fall; the islands in the sea are terrified at your collapse.'
EZEK|26|19|"This is what the Sovereign LORD says: When I make you a desolate city, like cities no longer inhabited, and when I bring the ocean depths over you and its vast waters cover you,
EZEK|26|20|then I will bring you down with those who go down to the pit, to the people of long ago. I will make you dwell in the earth below, as in ancient ruins, with those who go down to the pit, and you will not return or take your place in the land of the living.
EZEK|26|21|I will bring you to a horrible end and you will be no more. You will be sought, but you will never again be found, declares the Sovereign LORD."
EZEK|27|1|The word of the LORD came to me:
EZEK|27|2|"Son of man, take up a lament concerning Tyre.
EZEK|27|3|Say to Tyre, situated at the gateway to the sea, merchant of peoples on many coasts, 'This is what the Sovereign LORD says: "'You say, O Tyre, "I am perfect in beauty."
EZEK|27|4|Your domain was on the high seas; your builders brought your beauty to perfection.
EZEK|27|5|They made all your timbers of pine trees from Senir; they took a cedar from Lebanon to make a mast for you.
EZEK|27|6|Of oaks from Bashan they made your oars; of cypress wood from the coasts of Cyprus they made your deck, inlaid with ivory.
EZEK|27|7|Fine embroidered linen from Egypt was your sail and served as your banner; your awnings were of blue and purple from the coasts of Elishah.
EZEK|27|8|Men of Sidon and Arvad were your oarsmen; your skilled men, O Tyre, were aboard as your seamen.
EZEK|27|9|Veteran craftsmen of Gebal were on board as shipwrights to caulk your seams. All the ships of the sea and their sailors came alongside to trade for your wares.
EZEK|27|10|"'Men of Persia, Lydia and Put served as soldiers in your army. They hung their shields and helmets on your walls, bringing you splendor.
EZEK|27|11|Men of Arvad and Helech manned your walls on every side; men of Gammad were in your towers. They hung their shields around your walls; they brought your beauty to perfection.
EZEK|27|12|"'Tarshish did business with you because of your great wealth of goods; they exchanged silver, iron, tin and lead for your merchandise.
EZEK|27|13|"'Greece, Tubal and Meshech traded with you; they exchanged slaves and articles of bronze for your wares.
EZEK|27|14|"'Men of Beth Togarmah exchanged work horses, war horses and mules for your merchandise.
EZEK|27|15|"'The men of Rhodes traded with you, and many coastlands were your customers; they paid you with ivory tusks and ebony.
EZEK|27|16|"'Aram did business with you because of your many products; they exchanged turquoise, purple fabric, embroidered work, fine linen, coral and rubies for your merchandise.
EZEK|27|17|"'Judah and Israel traded with you; they exchanged wheat from Minnith and confections, honey, oil and balm for your wares.
EZEK|27|18|"'Damascus, because of your many products and great wealth of goods, did business with you in wine from Helbon and wool from Zahar.
EZEK|27|19|"'Danites and Greeks from Uzal bought your merchandise; they exchanged wrought iron, cassia and calamus for your wares.
EZEK|27|20|"'Dedan traded in saddle blankets with you.
EZEK|27|21|"'Arabia and all the princes of Kedar were your customers; they did business with you in lambs, rams and goats.
EZEK|27|22|"'The merchants of Sheba and Raamah traded with you; for your merchandise they exchanged the finest of all kinds of spices and precious stones, and gold.
EZEK|27|23|"'Haran, Canneh and Eden and merchants of Sheba, Asshur and Kilmad traded with you.
EZEK|27|24|In your marketplace they traded with you beautiful garments, blue fabric, embroidered work and multicolored rugs with cords twisted and tightly knotted.
EZEK|27|25|"'The ships of Tarshish serve as carriers for your wares. You are filled with heavy cargo in the heart of the sea.
EZEK|27|26|Your oarsmen take you out to the high seas. But the east wind will break you to pieces in the heart of the sea.
EZEK|27|27|Your wealth, merchandise and wares, your mariners, seamen and shipwrights, your merchants and all your soldiers, and everyone else on board will sink into the heart of the sea on the day of your shipwreck.
EZEK|27|28|The shorelands will quake when your seamen cry out.
EZEK|27|29|All who handle the oars will abandon their ships; the mariners and all the seamen will stand on the shore.
EZEK|27|30|They will raise their voice and cry bitterly over you; they will sprinkle dust on their heads and roll in ashes.
EZEK|27|31|They will shave their heads because of you and will put on sackcloth. They will weep over you with anguish of soul and with bitter mourning.
EZEK|27|32|As they wail and mourn over you, they will take up a lament concerning you: "Who was ever silenced like Tyre, surrounded by the sea?"
EZEK|27|33|When your merchandise went out on the seas, you satisfied many nations; with your great wealth and your wares you enriched the kings of the earth.
EZEK|27|34|Now you are shattered by the sea in the depths of the waters; your wares and all your company have gone down with you.
EZEK|27|35|All who live in the coastlands are appalled at you; their kings shudder with horror and their faces are distorted with fear.
EZEK|27|36|The merchants among the nations hiss at you; you have come to a horrible end and will be no more.'"
EZEK|28|1|The word of the LORD came to me:
EZEK|28|2|"Son of man, say to the ruler of Tyre, 'This is what the Sovereign LORD says: "'In the pride of your heart you say, "I am a god; I sit on the throne of a god in the heart of the seas." But you are a man and not a god, though you think you are as wise as a god.
EZEK|28|3|Are you wiser than Daniel? Is no secret hidden from you?
EZEK|28|4|By your wisdom and understanding you have gained wealth for yourself and amassed gold and silver in your treasuries.
EZEK|28|5|By your great skill in trading you have increased your wealth, and because of your wealth your heart has grown proud.
EZEK|28|6|"'Therefore this is what the Sovereign LORD says: "'Because you think you are wise, as wise as a god,
EZEK|28|7|I am going to bring foreigners against you, the most ruthless of nations; they will draw their swords against your beauty and wisdom and pierce your shining splendor.
EZEK|28|8|They will bring you down to the pit, and you will die a violent death in the heart of the seas.
EZEK|28|9|Will you then say, "I am a god," in the presence of those who kill you? You will be but a man, not a god, in the hands of those who slay you.
EZEK|28|10|You will die the death of the uncircumcised at the hands of foreigners. I have spoken, declares the Sovereign LORD.'"
EZEK|28|11|The word of the LORD came to me:
EZEK|28|12|"Son of man, take up a lament concerning the king of Tyre and say to him: 'This is what the Sovereign LORD says: "'You were the model of perfection, full of wisdom and perfect in beauty.
EZEK|28|13|You were in Eden, the garden of God; every precious stone adorned you: ruby, topaz and emerald, chrysolite, onyx and jasper, sapphire, turquoise and beryl. Your settings and mountings were made of gold; on the day you were created they were prepared.
EZEK|28|14|You were anointed as a guardian cherub, for so I ordained you. You were on the holy mount of God; you walked among the fiery stones.
EZEK|28|15|You were blameless in your ways from the day you were created till wickedness was found in you.
EZEK|28|16|Through your widespread trade you were filled with violence, and you sinned. So I drove you in disgrace from the mount of God, and I expelled you, O guardian cherub, from among the fiery stones.
EZEK|28|17|Your heart became proud on account of your beauty, and you corrupted your wisdom because of your splendor. So I threw you to the earth; I made a spectacle of you before kings.
EZEK|28|18|By your many sins and dishonest trade you have desecrated your sanctuaries. So I made a fire come out from you, and it consumed you, and I reduced you to ashes on the ground in the sight of all who were watching.
EZEK|28|19|All the nations who knew you are appalled at you; you have come to a horrible end and will be no more.'"
EZEK|28|20|The word of the LORD came to me:
EZEK|28|21|"Son of man, set your face against Sidon; prophesy against her
EZEK|28|22|and say: 'This is what the Sovereign LORD says: "'I am against you, O Sidon, and I will gain glory within you. They will know that I am the LORD, when I inflict punishment on her and show myself holy within her.
EZEK|28|23|I will send a plague upon her and make blood flow in her streets. The slain will fall within her, with the sword against her on every side. Then they will know that I am the LORD.
EZEK|28|24|"'No longer will the people of Israel have malicious neighbors who are painful briers and sharp thorns. Then they will know that I am the Sovereign LORD.
EZEK|28|25|"'This is what the Sovereign LORD says: When I gather the people of Israel from the nations where they have been scattered, I will show myself holy among them in the sight of the nations. Then they will live in their own land, which I gave to my servant Jacob.
EZEK|28|26|They will live there in safety and will build houses and plant vineyards; they will live in safety when I inflict punishment on all their neighbors who maligned them. Then they will know that I am the LORD their God.'"
EZEK|29|1|In the tenth year, in the tenth month on the twelfth day, the word of the LORD came to me:
EZEK|29|2|"Son of man, set your face against Pharaoh king of Egypt and prophesy against him and against all Egypt.
EZEK|29|3|Speak to him and say: 'This is what the Sovereign LORD says: "'I am against you, Pharaoh king of Egypt, you great monster lying among your streams. You say, "The Nile is mine; I made it for myself."
EZEK|29|4|But I will put hooks in your jaws and make the fish of your streams stick to your scales. I will pull you out from among your streams, with all the fish sticking to your scales.
EZEK|29|5|I will leave you in the desert, you and all the fish of your streams. You will fall on the open field and not be gathered or picked up. I will give you as food to the beasts of the earth and the birds of the air.
EZEK|29|6|Then all who live in Egypt will know that I am the LORD. "'You have been a staff of reed for the house of Israel.
EZEK|29|7|When they grasped you with their hands, you splintered and you tore open their shoulders; when they leaned on you, you broke and their backs were wrenched.
EZEK|29|8|"'Therefore this is what the Sovereign LORD says: I will bring a sword against you and kill your men and their animals.
EZEK|29|9|Egypt will become a desolate wasteland. Then they will know that I am the LORD. "'Because you said, "The Nile is mine; I made it,"
EZEK|29|10|therefore I am against you and against your streams, and I will make the land of Egypt a ruin and a desolate waste from Migdol to Aswan, as far as the border of Cush.
EZEK|29|11|No foot of man or animal will pass through it; no one will live there for forty years.
EZEK|29|12|I will make the land of Egypt desolate among devastated lands, and her cities will lie desolate forty years among ruined cities. And I will disperse the Egyptians among the nations and scatter them through the countries.
EZEK|29|13|"'Yet this is what the Sovereign LORD says: At the end of forty years I will gather the Egyptians from the nations where they were scattered.
EZEK|29|14|I will bring them back from captivity and return them to Upper Egypt, the land of their ancestry. There they will be a lowly kingdom.
EZEK|29|15|It will be the lowliest of kingdoms and will never again exalt itself above the other nations. I will make it so weak that it will never again rule over the nations.
EZEK|29|16|Egypt will no longer be a source of confidence for the people of Israel but will be a reminder of their sin in turning to her for help. Then they will know that I am the Sovereign LORD.'"
EZEK|29|17|In the twenty-seventh year, in the first month on the first day, the word of the LORD came to me:
EZEK|29|18|"Son of man, Nebuchadnezzar king of Babylon drove his army in a hard campaign against Tyre; every head was rubbed bare and every shoulder made raw. Yet he and his army got no reward from the campaign he led against Tyre.
EZEK|29|19|Therefore this is what the Sovereign LORD says: I am going to give Egypt to Nebuchadnezzar king of Babylon, and he will carry off its wealth. He will loot and plunder the land as pay for his army.
EZEK|29|20|I have given him Egypt as a reward for his efforts because he and his army did it for me, declares the Sovereign LORD.
EZEK|29|21|"On that day I will make a horn grow for the house of Israel, and I will open your mouth among them. Then they will know that I am the LORD."
EZEK|30|1|The word of the LORD came to me:
EZEK|30|2|"Son of man, prophesy and say: 'This is what the Sovereign LORD says: "'Wail and say, "Alas for that day!"
EZEK|30|3|For the day is near, the day of the LORD is near- a day of clouds, a time of doom for the nations.
EZEK|30|4|A sword will come against Egypt, and anguish will come upon Cush. When the slain fall in Egypt, her wealth will be carried away and her foundations torn down.
EZEK|30|5|Cush and Put, Lydia and all Arabia, Libya and the people of the covenant land will fall by the sword along with Egypt.
EZEK|30|6|"'This is what the LORD says: "'The allies of Egypt will fall and her proud strength will fail. From Migdol to Aswan they will fall by the sword within her, declares the Sovereign LORD.
EZEK|30|7|"'They will be desolate among desolate lands, and their cities will lie among ruined cities.
EZEK|30|8|Then they will know that I am the LORD, when I set fire to Egypt and all her helpers are crushed.
EZEK|30|9|"'On that day messengers will go out from me in ships to frighten Cush out of her complacency. Anguish will take hold of them on the day of Egypt's doom, for it is sure to come.
EZEK|30|10|"'This is what the Sovereign LORD says: "'I will put an end to the hordes of Egypt by the hand of Nebuchadnezzar king of Babylon.
EZEK|30|11|He and his army-the most ruthless of nations- will be brought in to destroy the land. They will draw their swords against Egypt and fill the land with the slain.
EZEK|30|12|I will dry up the streams of the Nile and sell the land to evil men; by the hand of foreigners I will lay waste the land and everything in it. I the LORD have spoken.
EZEK|30|13|"'This is what the Sovereign LORD says: "'I will destroy the idols and put an end to the images in Memphis. No longer will there be a prince in Egypt, and I will spread fear throughout the land.
EZEK|30|14|I will lay waste Upper Egypt, set fire to Zoan and inflict punishment on Thebes.
EZEK|30|15|I will pour out my wrath on Pelusium, the stronghold of Egypt, and cut off the hordes of Thebes.
EZEK|30|16|I will set fire to Egypt; Pelusium will writhe in agony. Thebes will be taken by storm; Memphis will be in constant distress.
EZEK|30|17|The young men of Heliopolis and Bubastis will fall by the sword, and the cities themselves will go into captivity.
EZEK|30|18|Dark will be the day at Tahpanhes when I break the yoke of Egypt; there her proud strength will come to an end. She will be covered with clouds, and her villages will go into captivity.
EZEK|30|19|So I will inflict punishment on Egypt, and they will know that I am the LORD.'"
EZEK|30|20|In the eleventh year, in the first month on the seventh day, the word of the LORD came to me:
EZEK|30|21|"Son of man, I have broken the arm of Pharaoh king of Egypt. It has not been bound up for healing or put in a splint so as to become strong enough to hold a sword.
EZEK|30|22|Therefore this is what the Sovereign LORD says: I am against Pharaoh king of Egypt. I will break both his arms, the good arm as well as the broken one, and make the sword fall from his hand.
EZEK|30|23|I will disperse the Egyptians among the nations and scatter them through the countries.
EZEK|30|24|I will strengthen the arms of the king of Babylon and put my sword in his hand, but I will break the arms of Pharaoh, and he will groan before him like a mortally wounded man.
EZEK|30|25|I will strengthen the arms of the king of Babylon, but the arms of Pharaoh will fall limp. Then they will know that I am the LORD, when I put my sword into the hand of the king of Babylon and he brandishes it against Egypt.
EZEK|30|26|I will disperse the Egyptians among the nations and scatter them through the countries. Then they will know that I am the LORD."
EZEK|31|1|In the eleventh year, in the third month on the first day, the word of the LORD came to me:
EZEK|31|2|"Son of man, say to Pharaoh king of Egypt and to his hordes: "'Who can be compared with you in majesty?
EZEK|31|3|Consider Assyria, once a cedar in Lebanon, with beautiful branches overshadowing the forest; it towered on high, its top above the thick foliage.
EZEK|31|4|The waters nourished it, deep springs made it grow tall; their streams flowed all around its base and sent their channels to all the trees of the field.
EZEK|31|5|So it towered higher than all the trees of the field; its boughs increased and its branches grew long, spreading because of abundant waters.
EZEK|31|6|All the birds of the air nested in its boughs, all the beasts of the field gave birth under its branches; all the great nations lived in its shade.
EZEK|31|7|It was majestic in beauty, with its spreading boughs, for its roots went down to abundant waters.
EZEK|31|8|The cedars in the garden of God could not rival it, nor could the pine trees equal its boughs, nor could the plane trees compare with its branches- no tree in the garden of God could match its beauty.
EZEK|31|9|I made it beautiful with abundant branches, the envy of all the trees of Eden in the garden of God.
EZEK|31|10|"'Therefore this is what the Sovereign LORD says: Because it towered on high, lifting its top above the thick foliage, and because it was proud of its height,
EZEK|31|11|I handed it over to the ruler of the nations, for him to deal with according to its wickedness. I cast it aside,
EZEK|31|12|and the most ruthless of foreign nations cut it down and left it. Its boughs fell on the mountains and in all the valleys; its branches lay broken in all the ravines of the land. All the nations of the earth came out from under its shade and left it.
EZEK|31|13|All the birds of the air settled on the fallen tree, and all the beasts of the field were among its branches.
EZEK|31|14|Therefore no other trees by the waters are ever to tower proudly on high, lifting their tops above the thick foliage. No other trees so well-watered are ever to reach such a height; they are all destined for death, for the earth below, among mortal men, with those who go down to the pit.
EZEK|31|15|"'This is what the Sovereign LORD says: On the day it was brought down to the grave I covered the deep springs with mourning for it; I held back its streams, and its abundant waters were restrained. Because of it I clothed Lebanon with gloom, and all the trees of the field withered away.
EZEK|31|16|I made the nations tremble at the sound of its fall when I brought it down to the grave with those who go down to the pit. Then all the trees of Eden, the choicest and best of Lebanon, all the trees that were well-watered, were consoled in the earth below.
EZEK|31|17|Those who lived in its shade, its allies among the nations, had also gone down to the grave with it, joining those killed by the sword.
EZEK|31|18|"'Which of the trees of Eden can be compared with you in splendor and majesty? Yet you, too, will be brought down with the trees of Eden to the earth below; you will lie among the uncircumcised, with those killed by the sword. "'This is Pharaoh and all his hordes, declares the Sovereign LORD.'"
EZEK|32|1|In the twelfth year, in the twelfth month on the first day, the word of the LORD came to me:
EZEK|32|2|"Son of man, take up a lament concerning Pharaoh king of Egypt and say to him: "'You are like a lion among the nations; you are like a monster in the seas thrashing about in your streams, churning the water with your feet and muddying the streams.
EZEK|32|3|"'This is what the Sovereign LORD says: "'With a great throng of people I will cast my net over you, and they will haul you up in my net.
EZEK|32|4|I will throw you on the land and hurl you on the open field. I will let all the birds of the air settle on you and all the beasts of the earth gorge themselves on you.
EZEK|32|5|I will spread your flesh on the mountains and fill the valleys with your remains.
EZEK|32|6|I will drench the land with your flowing blood all the way to the mountains, and the ravines will be filled with your flesh.
EZEK|32|7|When I snuff you out, I will cover the heavens and darken their stars; I will cover the sun with a cloud, and the moon will not give its light.
EZEK|32|8|All the shining lights in the heavens I will darken over you; I will bring darkness over your land, declares the Sovereign LORD.
EZEK|32|9|I will trouble the hearts of many peoples when I bring about your destruction among the nations, among lands you have not known.
EZEK|32|10|I will cause many peoples to be appalled at you, and their kings will shudder with horror because of you when I brandish my sword before them. On the day of your downfall each of them will tremble every moment for his life.
EZEK|32|11|"'For this is what the Sovereign LORD says: "'The sword of the king of Babylon will come against you.
EZEK|32|12|I will cause your hordes to fall by the swords of mighty men- the most ruthless of all nations. They will shatter the pride of Egypt, and all her hordes will be overthrown.
EZEK|32|13|I will destroy all her cattle from beside abundant waters no longer to be stirred by the foot of man or muddied by the hoofs of cattle.
EZEK|32|14|Then I will let her waters settle and make her streams flow like oil, declares the Sovereign LORD.
EZEK|32|15|When I make Egypt desolate and strip the land of everything in it, when I strike down all who live there, then they will know that I am the LORD.'
EZEK|32|16|"This is the lament they will chant for her. The daughters of the nations will chant it; for Egypt and all her hordes they will chant it, declares the Sovereign LORD."
EZEK|32|17|In the twelfth year, on the fifteenth day of the month, the word of the LORD came to me:
EZEK|32|18|"Son of man, wail for the hordes of Egypt and consign to the earth below both her and the daughters of mighty nations, with those who go down to the pit.
EZEK|32|19|Say to them, 'Are you more favored than others? Go down and be laid among the uncircumcised.'
EZEK|32|20|They will fall among those killed by the sword. The sword is drawn; let her be dragged off with all her hordes.
EZEK|32|21|From within the grave the mighty leaders will say of Egypt and her allies, 'They have come down and they lie with the uncircumcised, with those killed by the sword.'
EZEK|32|22|"Assyria is there with her whole army; she is surrounded by the graves of all her slain, all who have fallen by the sword.
EZEK|32|23|Their graves are in the depths of the pit and her army lies around her grave. All who had spread terror in the land of the living are slain, fallen by the sword.
EZEK|32|24|"Elam is there, with all her hordes around her grave. All of them are slain, fallen by the sword. All who had spread terror in the land of the living went down uncircumcised to the earth below. They bear their shame with those who go down to the pit.
EZEK|32|25|A bed is made for her among the slain, with all her hordes around her grave. All of them are uncircumcised, killed by the sword. Because their terror had spread in the land of the living, they bear their shame with those who go down to the pit; they are laid among the slain.
EZEK|32|26|"Meshech and Tubal are there, with all their hordes around their graves. All of them are uncircumcised, killed by the sword because they spread their terror in the land of the living.
EZEK|32|27|Do they not lie with the other uncircumcised warriors who have fallen, who went down to the grave with their weapons of war, whose swords were placed under their heads? The punishment for their sins rested on their bones, though the terror of these warriors had stalked through the land of the living.
EZEK|32|28|"You too, O Pharaoh, will be broken and will lie among the uncircumcised, with those killed by the sword.
EZEK|32|29|"Edom is there, her kings and all her princes; despite their power, they are laid with those killed by the sword. They lie with the uncircumcised, with those who go down to the pit.
EZEK|32|30|"All the princes of the north and all the Sidonians are there; they went down with the slain in disgrace despite the terror caused by their power. They lie uncircumcised with those killed by the sword and bear their shame with those who go down to the pit.
EZEK|32|31|"Pharaoh-he and all his army-will see them and he will be consoled for all his hordes that were killed by the sword, declares the Sovereign LORD.
EZEK|32|32|Although I had him spread terror in the land of the living, Pharaoh and all his hordes will be laid among the uncircumcised, with those killed by the sword, declares the Sovereign LORD."
EZEK|33|1|The word of the LORD came to me:
EZEK|33|2|"Son of man, speak to your countrymen and say to them: 'When I bring the sword against a land, and the people of the land choose one of their men and make him their watchman,
EZEK|33|3|and he sees the sword coming against the land and blows the trumpet to warn the people,
EZEK|33|4|then if anyone hears the trumpet but does not take warning and the sword comes and takes his life, his blood will be on his own head.
EZEK|33|5|Since he heard the sound of the trumpet but did not take warning, his blood will be on his own head. If he had taken warning, he would have saved himself.
EZEK|33|6|But if the watchman sees the sword coming and does not blow the trumpet to warn the people and the sword comes and takes the life of one of them, that man will be taken away because of his sin, but I will hold the watchman accountable for his blood.'
EZEK|33|7|"Son of man, I have made you a watchman for the house of Israel; so hear the word I speak and give them warning from me.
EZEK|33|8|When I say to the wicked, 'O wicked man, you will surely die,' and you do not speak out to dissuade him from his ways, that wicked man will die for his sin, and I will hold you accountable for his blood.
EZEK|33|9|But if you do warn the wicked man to turn from his ways and he does not do so, he will die for his sin, but you will have saved yourself.
EZEK|33|10|"Son of man, say to the house of Israel, 'This is what you are saying: "Our offenses and sins weigh us down, and we are wasting away because of them. How then can we live?"'
EZEK|33|11|Say to them, 'As surely as I live, declares the Sovereign LORD, I take no pleasure in the death of the wicked, but rather that they turn from their ways and live. Turn! Turn from your evil ways! Why will you die, O house of Israel?'
EZEK|33|12|"Therefore, son of man, say to your countrymen, 'The righteousness of the righteous man will not save him when he disobeys, and the wickedness of the wicked man will not cause him to fall when he turns from it. The righteous man, if he sins, will not be allowed to live because of his former righteousness.'
EZEK|33|13|If I tell the righteous man that he will surely live, but then he trusts in his righteousness and does evil, none of the righteous things he has done will be remembered; he will die for the evil he has done.
EZEK|33|14|And if I say to the wicked man, 'You will surely die,' but he then turns away from his sin and does what is just and right-
EZEK|33|15|if he gives back what he took in pledge for a loan, returns what he has stolen, follows the decrees that give life, and does no evil, he will surely live; he will not die.
EZEK|33|16|None of the sins he has committed will be remembered against him. He has done what is just and right; he will surely live.
EZEK|33|17|"Yet your countrymen say, 'The way of the Lord is not just.' But it is their way that is not just.
EZEK|33|18|If a righteous man turns from his righteousness and does evil, he will die for it.
EZEK|33|19|And if a wicked man turns away from his wickedness and does what is just and right, he will live by doing so.
EZEK|33|20|Yet, O house of Israel, you say, 'The way of the Lord is not just.' But I will judge each of you according to his own ways."
EZEK|33|21|In the twelfth year of our exile, in the tenth month on the fifth day, a man who had escaped from Jerusalem came to me and said, "The city has fallen!"
EZEK|33|22|Now the evening before the man arrived, the hand of the LORD was upon me, and he opened my mouth before the man came to me in the morning. So my mouth was opened and I was no longer silent.
EZEK|33|23|Then the word of the LORD came to me:
EZEK|33|24|"Son of man, the people living in those ruins in the land of Israel are saying, 'Abraham was only one man, yet he possessed the land. But we are many; surely the land has been given to us as our possession.'
EZEK|33|25|Therefore say to them, 'This is what the Sovereign LORD says: Since you eat meat with the blood still in it and look to your idols and shed blood, should you then possess the land?
EZEK|33|26|You rely on your sword, you do detestable things, and each of you defiles his neighbor's wife. Should you then possess the land?'
EZEK|33|27|"Say this to them: 'This is what the Sovereign LORD says: As surely as I live, those who are left in the ruins will fall by the sword, those out in the country I will give to the wild animals to be devoured, and those in strongholds and caves will die of a plague.
EZEK|33|28|I will make the land a desolate waste, and her proud strength will come to an end, and the mountains of Israel will become desolate so that no one will cross them.
EZEK|33|29|Then they will know that I am the LORD, when I have made the land a desolate waste because of all the detestable things they have done.'
EZEK|33|30|"As for you, son of man, your countrymen are talking together about you by the walls and at the doors of the houses, saying to each other, 'Come and hear the message that has come from the LORD.'
EZEK|33|31|My people come to you, as they usually do, and sit before you to listen to your words, but they do not put them into practice. With their mouths they express devotion, but their hearts are greedy for unjust gain.
EZEK|33|32|Indeed, to them you are nothing more than one who sings love songs with a beautiful voice and plays an instrument well, for they hear your words but do not put them into practice.
EZEK|33|33|"When all this comes true-and it surely will-then they will know that a prophet has been among them."
EZEK|34|1|The word of the LORD came to me:
EZEK|34|2|"Son of man, prophesy against the shepherds of Israel; prophesy and say to them: 'This is what the Sovereign LORD says: Woe to the shepherds of Israel who only take care of themselves! Should not shepherds take care of the flock?
EZEK|34|3|You eat the curds, clothe yourselves with the wool and slaughter the choice animals, but you do not take care of the flock.
EZEK|34|4|You have not strengthened the weak or healed the sick or bound up the injured. You have not brought back the strays or searched for the lost. You have ruled them harshly and brutally.
EZEK|34|5|So they were scattered because there was no shepherd, and when they were scattered they became food for all the wild animals.
EZEK|34|6|My sheep wandered over all the mountains and on every high hill. They were scattered over the whole earth, and no one searched or looked for them.
EZEK|34|7|"'Therefore, you shepherds, hear the word of the LORD:
EZEK|34|8|As surely as I live, declares the Sovereign LORD, because my flock lacks a shepherd and so has been plundered and has become food for all the wild animals, and because my shepherds did not search for my flock but cared for themselves rather than for my flock,
EZEK|34|9|therefore, O shepherds, hear the word of the LORD:
EZEK|34|10|This is what the Sovereign LORD says: I am against the shepherds and will hold them accountable for my flock. I will remove them from tending the flock so that the shepherds can no longer feed themselves. I will rescue my flock from their mouths, and it will no longer be food for them.
EZEK|34|11|"'For this is what the Sovereign LORD says: I myself will search for my sheep and look after them.
EZEK|34|12|As a shepherd looks after his scattered flock when he is with them, so will I look after my sheep. I will rescue them from all the places where they were scattered on a day of clouds and darkness.
EZEK|34|13|I will bring them out from the nations and gather them from the countries, and I will bring them into their own land. I will pasture them on the mountains of Israel, in the ravines and in all the settlements in the land.
EZEK|34|14|I will tend them in a good pasture, and the mountain heights of Israel will be their grazing land. There they will lie down in good grazing land, and there they will feed in a rich pasture on the mountains of Israel.
EZEK|34|15|I myself will tend my sheep and have them lie down, declares the Sovereign LORD.
EZEK|34|16|I will search for the lost and bring back the strays. I will bind up the injured and strengthen the weak, but the sleek and the strong I will destroy. I will shepherd the flock with justice.
EZEK|34|17|"'As for you, my flock, this is what the Sovereign LORD says: I will judge between one sheep and another, and between rams and goats.
EZEK|34|18|Is it not enough for you to feed on the good pasture? Must you also trample the rest of your pasture with your feet? Is it not enough for you to drink clear water? Must you also muddy the rest with your feet?
EZEK|34|19|Must my flock feed on what you have trampled and drink what you have muddied with your feet?
EZEK|34|20|"'Therefore this is what the Sovereign LORD says to them: See, I myself will judge between the fat sheep and the lean sheep.
EZEK|34|21|Because you shove with flank and shoulder, butting all the weak sheep with your horns until you have driven them away,
EZEK|34|22|I will save my flock, and they will no longer be plundered. I will judge between one sheep and another.
EZEK|34|23|I will place over them one shepherd, my servant David, and he will tend them; he will tend them and be their shepherd.
EZEK|34|24|I the LORD will be their God, and my servant David will be prince among them. I the LORD have spoken.
EZEK|34|25|"'I will make a covenant of peace with them and rid the land of wild beasts so that they may live in the desert and sleep in the forests in safety.
EZEK|34|26|I will bless them and the places surrounding my hill. I will send down showers in season; there will be showers of blessing.
EZEK|34|27|The trees of the field will yield their fruit and the ground will yield its crops; the people will be secure in their land. They will know that I am the LORD, when I break the bars of their yoke and rescue them from the hands of those who enslaved them.
EZEK|34|28|They will no longer be plundered by the nations, nor will wild animals devour them. They will live in safety, and no one will make them afraid.
EZEK|34|29|I will provide for them a land renowned for its crops, and they will no longer be victims of famine in the land or bear the scorn of the nations.
EZEK|34|30|Then they will know that I, the LORD their God, am with them and that they, the house of Israel, are my people, declares the Sovereign LORD.
EZEK|34|31|You my sheep, the sheep of my pasture, are people, and I am your God, declares the Sovereign LORD.'"
EZEK|35|1|The word of the LORD came to me:
EZEK|35|2|"Son of man, set your face against Mount Seir; prophesy against it
EZEK|35|3|and say: 'This is what the Sovereign LORD says: I am against you, Mount Seir, and I will stretch out my hand against you and make you a desolate waste.
EZEK|35|4|I will turn your towns into ruins and you will be desolate. Then you will know that I am the LORD.
EZEK|35|5|"'Because you harbored an ancient hostility and delivered the Israelites over to the sword at the time of their calamity, the time their punishment reached its climax,
EZEK|35|6|therefore as surely as I live, declares the Sovereign LORD, I will give you over to bloodshed and it will pursue you. Since you did not hate bloodshed, bloodshed will pursue you.
EZEK|35|7|I will make Mount Seir a desolate waste and cut off from it all who come and go.
EZEK|35|8|I will fill your mountains with the slain; those killed by the sword will fall on your hills and in your valleys and in all your ravines.
EZEK|35|9|I will make you desolate forever; your towns will not be inhabited. Then you will know that I am the LORD.
EZEK|35|10|"'Because you have said, "These two nations and countries will be ours and we will take possession of them," even though I the LORD was there,
EZEK|35|11|therefore as surely as I live, declares the Sovereign LORD, I will treat you in accordance with the anger and jealousy you showed in your hatred of them and I will make myself known among them when I judge you.
EZEK|35|12|Then you will know that I the LORD have heard all the contemptible things you have said against the mountains of Israel. You said, "They have been laid waste and have been given over to us to devour."
EZEK|35|13|You boasted against me and spoke against me without restraint, and I heard it.
EZEK|35|14|This is what the Sovereign LORD says: While the whole earth rejoices, I will make you desolate.
EZEK|35|15|Because you rejoiced when the inheritance of the house of Israel became desolate, that is how I will treat you. You will be desolate, O Mount Seir, you and all of Edom. Then they will know that I am the LORD.'"
EZEK|36|1|"Son of man, prophesy to the mountains of Israel and say, 'O mountains of Israel, hear the word of the LORD.
EZEK|36|2|This is what the Sovereign LORD says: The enemy said of you, "Aha! The ancient heights have become our possession."'
EZEK|36|3|Therefore prophesy and say, 'This is what the Sovereign LORD says: Because they ravaged and hounded you from every side so that you became the possession of the rest of the nations and the object of people's malicious talk and slander,
EZEK|36|4|therefore, O mountains of Israel, hear the word of the Sovereign LORD: This is what the Sovereign LORD says to the mountains and hills, to the ravines and valleys, to the desolate ruins and the deserted towns that have been plundered and ridiculed by the rest of the nations around you-
EZEK|36|5|this is what the Sovereign LORD says: In my burning zeal I have spoken against the rest of the nations, and against all Edom, for with glee and with malice in their hearts they made my land their own possession so that they might plunder its pastureland.'
EZEK|36|6|Therefore prophesy concerning the land of Israel and say to the mountains and hills, to the ravines and valleys: 'This is what the Sovereign LORD says: I speak in my jealous wrath because you have suffered the scorn of the nations.
EZEK|36|7|Therefore this is what the Sovereign LORD says: I swear with uplifted hand that the nations around you will also suffer scorn.
EZEK|36|8|"'But you, O mountains of Israel, will produce branches and fruit for my people Israel, for they will soon come home.
EZEK|36|9|I am concerned for you and will look on you with favor; you will be plowed and sown,
EZEK|36|10|and I will multiply the number of people upon you, even the whole house of Israel. The towns will be inhabited and the ruins rebuilt.
EZEK|36|11|I will increase the number of men and animals upon you, and they will be fruitful and become numerous. I will settle people on you as in the past and will make you prosper more than before. Then you will know that I am the LORD.
EZEK|36|12|I will cause people, my people Israel, to walk upon you. They will possess you, and you will be their inheritance; you will never again deprive them of their children.
EZEK|36|13|"'This is what the Sovereign LORD says: Because people say to you, "You devour men and deprive your nation of its children,"
EZEK|36|14|therefore you will no longer devour men or make your nation childless, declares the Sovereign LORD.
EZEK|36|15|No longer will I make you hear the taunts of the nations, and no longer will you suffer the scorn of the peoples or cause your nation to fall, declares the Sovereign LORD.'"
EZEK|36|16|Again the word of the LORD came to me:
EZEK|36|17|"Son of man, when the people of Israel were living in their own land, they defiled it by their conduct and their actions. Their conduct was like a woman's monthly uncleanness in my sight.
EZEK|36|18|So I poured out my wrath on them because they had shed blood in the land and because they had defiled it with their idols.
EZEK|36|19|I dispersed them among the nations, and they were scattered through the countries; I judged them according to their conduct and their actions.
EZEK|36|20|And wherever they went among the nations they profaned my holy name, for it was said of them, 'These are the LORD 's people, and yet they had to leave his land.'
EZEK|36|21|I had concern for my holy name, which the house of Israel profaned among the nations where they had gone.
EZEK|36|22|"Therefore say to the house of Israel, 'This is what the Sovereign LORD says: It is not for your sake, O house of Israel, that I am going to do these things, but for the sake of my holy name, which you have profaned among the nations where you have gone.
EZEK|36|23|I will show the holiness of my great name, which has been profaned among the nations, the name you have profaned among them. Then the nations will know that I am the LORD, declares the Sovereign LORD, when I show myself holy through you before their eyes.
EZEK|36|24|"'For I will take you out of the nations; I will gather you from all the countries and bring you back into your own land.
EZEK|36|25|I will sprinkle clean water on you, and you will be clean; I will cleanse you from all your impurities and from all your idols.
EZEK|36|26|I will give you a new heart and put a new spirit in you; I will remove from you your heart of stone and give you a heart of flesh.
EZEK|36|27|And I will put my Spirit in you and move you to follow my decrees and be careful to keep my laws.
EZEK|36|28|You will live in the land I gave your forefathers; you will be my people, and I will be your God.
EZEK|36|29|I will save you from all your uncleanness. I will call for the grain and make it plentiful and will not bring famine upon you.
EZEK|36|30|I will increase the fruit of the trees and the crops of the field, so that you will no longer suffer disgrace among the nations because of famine.
EZEK|36|31|Then you will remember your evil ways and wicked deeds, and you will loathe yourselves for your sins and detestable practices.
EZEK|36|32|I want you to know that I am not doing this for your sake, declares the Sovereign LORD. Be ashamed and disgraced for your conduct, O house of Israel!
EZEK|36|33|"'This is what the Sovereign LORD says: On the day I cleanse you from all your sins, I will resettle your towns, and the ruins will be rebuilt.
EZEK|36|34|The desolate land will be cultivated instead of lying desolate in the sight of all who pass through it.
EZEK|36|35|They will say, "This land that was laid waste has become like the garden of Eden; the cities that were lying in ruins, desolate and destroyed, are now fortified and inhabited."
EZEK|36|36|Then the nations around you that remain will know that I the LORD have rebuilt what was destroyed and have replanted what was desolate. I the LORD have spoken, and I will do it.'
EZEK|36|37|"This is what the Sovereign LORD says: Once again I will yield to the plea of the house of Israel and do this for them: I will make their people as numerous as sheep,
EZEK|36|38|as numerous as the flocks for offerings at Jerusalem during her appointed feasts. So will the ruined cities be filled with flocks of people. Then they will know that I am the LORD."
EZEK|37|1|The hand of the LORD was upon me, and he brought me out by the Spirit of the LORD and set me in the middle of a valley; it was full of bones.
EZEK|37|2|He led me back and forth among them, and I saw a great many bones on the floor of the valley, bones that were very dry.
EZEK|37|3|He asked me, "Son of man, can these bones live?" I said, "O Sovereign LORD, you alone know."
EZEK|37|4|Then he said to me, "Prophesy to these bones and say to them, 'Dry bones, hear the word of the LORD!
EZEK|37|5|This is what the Sovereign LORD says to these bones: I will make breath enter you, and you will come to life.
EZEK|37|6|I will attach tendons to you and make flesh come upon you and cover you with skin; I will put breath in you, and you will come to life. Then you will know that I am the LORD.'"
EZEK|37|7|So I prophesied as I was commanded. And as I was prophesying, there was a noise, a rattling sound, and the bones came together, bone to bone.
EZEK|37|8|I looked, and tendons and flesh appeared on them and skin covered them, but there was no breath in them.
EZEK|37|9|Then he said to me, "Prophesy to the breath; prophesy, son of man, and say to it, 'This is what the Sovereign LORD says: Come from the four winds, O breath, and breathe into these slain, that they may live.'"
EZEK|37|10|So I prophesied as he commanded me, and breath entered them; they came to life and stood up on their feet-a vast army.
EZEK|37|11|Then he said to me: "Son of man, these bones are the whole house of Israel. They say, 'Our bones are dried up and our hope is gone; we are cut off.'
EZEK|37|12|Therefore prophesy and say to them: 'This is what the Sovereign LORD says: O my people, I am going to open your graves and bring you up from them; I will bring you back to the land of Israel.
EZEK|37|13|Then you, my people, will know that I am the LORD, when I open your graves and bring you up from them.
EZEK|37|14|I will put my Spirit in you and you will live, and I will settle you in your own land. Then you will know that I the LORD have spoken, and I have done it, declares the LORD.'"
EZEK|37|15|The word of the LORD came to me:
EZEK|37|16|"Son of man, take a stick of wood and write on it, 'Belonging to Judah and the Israelites associated with him.' Then take another stick of wood, and write on it, 'Ephraim's stick, belonging to Joseph and all the house of Israel associated with him.'
EZEK|37|17|Join them together into one stick so that they will become one in your hand.
EZEK|37|18|"When your countrymen ask you, 'Won't you tell us what you mean by this?'
EZEK|37|19|say to them, 'This is what the Sovereign LORD says: I am going to take the stick of Joseph-which is in Ephraim's hand-and of the Israelite tribes associated with him, and join it to Judah's stick, making them a single stick of wood, and they will become one in my hand.'
EZEK|37|20|Hold before their eyes the sticks you have written on
EZEK|37|21|and say to them, 'This is what the Sovereign LORD says: I will take the Israelites out of the nations where they have gone. I will gather them from all around and bring them back into their own land.
EZEK|37|22|I will make them one nation in the land, on the mountains of Israel. There will be one king over all of them and they will never again be two nations or be divided into two kingdoms.
EZEK|37|23|They will no longer defile themselves with their idols and vile images or with any of their offenses, for I will save them from all their sinful backsliding, and I will cleanse them. They will be my people, and I will be their God.
EZEK|37|24|"'My servant David will be king over them, and they will all have one shepherd. They will follow my laws and be careful to keep my decrees.
EZEK|37|25|They will live in the land I gave to my servant Jacob, the land where your fathers lived. They and their children and their children's children will live there forever, and David my servant will be their prince forever.
EZEK|37|26|I will make a covenant of peace with them; it will be an everlasting covenant. I will establish them and increase their numbers, and I will put my sanctuary among them forever.
EZEK|37|27|My dwelling place will be with them; I will be their God, and they will be my people.
EZEK|37|28|Then the nations will know that I the LORD make Israel holy, when my sanctuary is among them forever.'"
EZEK|38|1|The word of the LORD came to me:
EZEK|38|2|"Son of man, set your face against Gog, of the land of Magog, the chief prince of Meshech and Tubal; prophesy against him
EZEK|38|3|and say: 'This is what the Sovereign LORD says: I am against you, O Gog, chief prince of Meshech and Tubal.
EZEK|38|4|I will turn you around, put hooks in your jaws and bring you out with your whole army-your horses, your horsemen fully armed, and a great horde with large and small shields, all of them brandishing their swords.
EZEK|38|5|Persia, Cush and Put will be with them, all with shields and helmets,
EZEK|38|6|also Gomer with all its troops, and Beth Togarmah from the far north with all its troops-the many nations with you.
EZEK|38|7|"'Get ready; be prepared, you and all the hordes gathered about you, and take command of them.
EZEK|38|8|After many days you will be called to arms. In future years you will invade a land that has recovered from war, whose people were gathered from many nations to the mountains of Israel, which had long been desolate. They had been brought out from the nations, and now all of them live in safety.
EZEK|38|9|You and all your troops and the many nations with you will go up, advancing like a storm; you will be like a cloud covering the land.
EZEK|38|10|"'This is what the Sovereign LORD says: On that day thoughts will come into your mind and you will devise an evil scheme.
EZEK|38|11|You will say, "I will invade a land of unwalled villages; I will attack a peaceful and unsuspecting people-all of them living without walls and without gates and bars.
EZEK|38|12|I will plunder and loot and turn my hand against the resettled ruins and the people gathered from the nations, rich in livestock and goods, living at the center of the land."
EZEK|38|13|Sheba and Dedan and the merchants of Tarshish and all her villages will say to you, "Have you come to plunder? Have you gathered your hordes to loot, to carry off silver and gold, to take away livestock and goods and to seize much plunder?"'
EZEK|38|14|"Therefore, son of man, prophesy and say to Gog: 'This is what the Sovereign LORD says: In that day, when my people Israel are living in safety, will you not take notice of it?
EZEK|38|15|You will come from your place in the far north, you and many nations with you, all of them riding on horses, a great horde, a mighty army.
EZEK|38|16|You will advance against my people Israel like a cloud that covers the land. In days to come, O Gog, I will bring you against my land, so that the nations may know me when I show myself holy through you before their eyes.
EZEK|38|17|"'This is what the Sovereign LORD says: Are you not the one I spoke of in former days by my servants the prophets of Israel? At that time they prophesied for years that I would bring you against them.
EZEK|38|18|This is what will happen in that day: When Gog attacks the land of Israel, my hot anger will be aroused, declares the Sovereign LORD.
EZEK|38|19|In my zeal and fiery wrath I declare that at that time there shall be a great earthquake in the land of Israel.
EZEK|38|20|The fish of the sea, the birds of the air, the beasts of the field, every creature that moves along the ground, and all the people on the face of the earth will tremble at my presence. The mountains will be overturned, the cliffs will crumble and every wall will fall to the ground.
EZEK|38|21|I will summon a sword against Gog on all my mountains, declares the Sovereign LORD. Every man's sword will be against his brother.
EZEK|38|22|I will execute judgment upon him with plague and bloodshed; I will pour down torrents of rain, hailstones and burning sulfur on him and on his troops and on the many nations with him.
EZEK|38|23|And so I will show my greatness and my holiness, and I will make myself known in the sight of many nations. Then they will know that I am the LORD.'
EZEK|39|1|"Son of man, prophesy against Gog and say: 'This is what the Sovereign LORD says: I am against you, O Gog, chief prince of Meshech and Tubal.
EZEK|39|2|I will turn you around and drag you along. I will bring you from the far north and send you against the mountains of Israel.
EZEK|39|3|Then I will strike your bow from your left hand and make your arrows drop from your right hand.
EZEK|39|4|On the mountains of Israel you will fall, you and all your troops and the nations with you. I will give you as food to all kinds of carrion birds and to the wild animals.
EZEK|39|5|You will fall in the open field, for I have spoken, declares the Sovereign LORD.
EZEK|39|6|I will send fire on Magog and on those who live in safety in the coastlands, and they will know that I am the LORD.
EZEK|39|7|"'I will make known my holy name among my people Israel. I will no longer let my holy name be profaned, and the nations will know that I the LORD am the Holy One in Israel.
EZEK|39|8|It is coming! It will surely take place, declares the Sovereign LORD. This is the day I have spoken of.
EZEK|39|9|"'Then those who live in the towns of Israel will go out and use the weapons for fuel and burn them up-the small and large shields, the bows and arrows, the war clubs and spears. For seven years they will use them for fuel.
EZEK|39|10|They will not need to gather wood from the fields or cut it from the forests, because they will use the weapons for fuel. And they will plunder those who plundered them and loot those who looted them, declares the Sovereign LORD.
EZEK|39|11|"'On that day I will give Gog a burial place in Israel, in the valley of those who travel east toward the Sea. It will block the way of travelers, because Gog and all his hordes will be buried there. So it will be called the Valley of Hamon Gog.
EZEK|39|12|"'For seven months the house of Israel will be burying them in order to cleanse the land.
EZEK|39|13|All the people of the land will bury them, and the day I am glorified will be a memorable day for them, declares the Sovereign LORD.
EZEK|39|14|"'Men will be regularly employed to cleanse the land. Some will go throughout the land and, in addition to them, others will bury those that remain on the ground. At the end of the seven months they will begin their search.
EZEK|39|15|As they go through the land and one of them sees a human bone, he will set up a marker beside it until the gravediggers have buried it in the Valley of Hamon Gog.
EZEK|39|16|(Also a town called Hamonah will be there.) And so they will cleanse the land.'
EZEK|39|17|"Son of man, this is what the Sovereign LORD says: Call out to every kind of bird and all the wild animals: 'Assemble and come together from all around to the sacrifice I am preparing for you, the great sacrifice on the mountains of Israel. There you will eat flesh and drink blood.
EZEK|39|18|You will eat the flesh of mighty men and drink the blood of the princes of the earth as if they were rams and lambs, goats and bulls-all of them fattened animals from Bashan.
EZEK|39|19|At the sacrifice I am preparing for you, you will eat fat till you are glutted and drink blood till you are drunk.
EZEK|39|20|At my table you will eat your fill of horses and riders, mighty men and soldiers of every kind,' declares the Sovereign LORD.
EZEK|39|21|"I will display my glory among the nations, and all the nations will see the punishment I inflict and the hand I lay upon them.
EZEK|39|22|From that day forward the house of Israel will know that I am the LORD their God.
EZEK|39|23|And the nations will know that the people of Israel went into exile for their sin, because they were unfaithful to me. So I hid my face from them and handed them over to their enemies, and they all fell by the sword.
EZEK|39|24|I dealt with them according to their uncleanness and their offenses, and I hid my face from them.
EZEK|39|25|"Therefore this is what the Sovereign LORD says: I will now bring Jacob back from captivity and will have compassion on all the people of Israel, and I will be zealous for my holy name.
EZEK|39|26|They will forget their shame and all the unfaithfulness they showed toward me when they lived in safety in their land with no one to make them afraid.
EZEK|39|27|When I have brought them back from the nations and have gathered them from the countries of their enemies, I will show myself holy through them in the sight of many nations.
EZEK|39|28|Then they will know that I am the LORD their God, for though I sent them into exile among the nations, I will gather them to their own land, not leaving any behind.
EZEK|39|29|I will no longer hide my face from them, for I will pour out my Spirit on the house of Israel, declares the Sovereign LORD."
EZEK|40|1|In the twenty-fifth year of our exile, at the beginning of the year, on the tenth of the month, in the fourteenth year after the fall of the city-on that very day the hand of the LORD was upon me and he took me there.
EZEK|40|2|In visions of God he took me to the land of Israel and set me on a very high mountain, on whose south side were some buildings that looked like a city.
EZEK|40|3|He took me there, and I saw a man whose appearance was like bronze; he was standing in the gateway with a linen cord and a measuring rod in his hand.
EZEK|40|4|The man said to me, "Son of man, look with your eyes and hear with your ears and pay attention to everything I am going to show you, for that is why you have been brought here. Tell the house of Israel everything you see."
EZEK|40|5|I saw a wall completely surrounding the temple area. The length of the measuring rod in the man's hand was six long cubits, each of which was a cubit and a handbreadth. He measured the wall; it was one measuring rod thick and one rod high.
EZEK|40|6|Then he went to the gate facing east. He climbed its steps and measured the threshold of the gate; it was one rod deep.
EZEK|40|7|The alcoves for the guards were one rod long and one rod wide, and the projecting walls between the alcoves were five cubits thick. And the threshold of the gate next to the portico facing the temple was one rod deep.
EZEK|40|8|Then he measured the portico of the gateway;
EZEK|40|9|it was eight cubits deep and its jambs were two cubits thick. The portico of the gateway faced the temple.
EZEK|40|10|Inside the east gate were three alcoves on each side; the three had the same measurements, and the faces of the projecting walls on each side had the same measurements.
EZEK|40|11|Then he measured the width of the entrance to the gateway; it was ten cubits and its length was thirteen cubits.
EZEK|40|12|In front of each alcove was a wall one cubit high, and the alcoves were six cubits square.
EZEK|40|13|Then he measured the gateway from the top of the rear wall of one alcove to the top of the opposite one; the distance was twenty-five cubits from one parapet opening to the opposite one.
EZEK|40|14|He measured along the faces of the projecting walls all around the inside of the gateway-sixty cubits. The measurement was up to the portico facing the courtyard.
EZEK|40|15|The distance from the entrance of the gateway to the far end of its portico was fifty cubits.
EZEK|40|16|The alcoves and the projecting walls inside the gateway were surmounted by narrow parapet openings all around, as was the portico; the openings all around faced inward. The faces of the projecting walls were decorated with palm trees.
EZEK|40|17|Then he brought me into the outer court. There I saw some rooms and a pavement that had been constructed all around the court; there were thirty rooms along the pavement.
EZEK|40|18|It abutted the sides of the gateways and was as wide as they were long; this was the lower pavement.
EZEK|40|19|Then he measured the distance from the inside of the lower gateway to the outside of the inner court; it was a hundred cubits on the east side as well as on the north.
EZEK|40|20|Then he measured the length and width of the gate facing north, leading into the outer court.
EZEK|40|21|Its alcoves-three on each side-its projecting walls and its portico had the same measurements as those of the first gateway. It was fifty cubits long and twenty-five cubits wide.
EZEK|40|22|Its openings, its portico and its palm tree decorations had the same measurements as those of the gate facing east. Seven steps led up to it, with its portico opposite them.
EZEK|40|23|There was a gate to the inner court facing the north gate, just as there was on the east. He measured from one gate to the opposite one; it was a hundred cubits.
EZEK|40|24|Then he led me to the south side and I saw a gate facing south. He measured its jambs and its portico, and they had the same measurements as the others.
EZEK|40|25|The gateway and its portico had narrow openings all around, like the openings of the others. It was fifty cubits long and twenty-five cubits wide.
EZEK|40|26|Seven steps led up to it, with its portico opposite them; it had palm tree decorations on the faces of the projecting walls on each side.
EZEK|40|27|The inner court also had a gate facing south, and he measured from this gate to the outer gate on the south side; it was a hundred cubits.
EZEK|40|28|Then he brought me into the inner court through the south gate, and he measured the south gate; it had the same measurements as the others.
EZEK|40|29|Its alcoves, its projecting walls and its portico had the same measurements as the others. The gateway and its portico had openings all around. It was fifty cubits long and twenty-five cubits wide.
EZEK|40|30|(The porticoes of the gateways around the inner court were twenty-five cubits wide and five cubits deep.)
EZEK|40|31|Its portico faced the outer court; palm trees decorated its jambs, and eight steps led up to it.
EZEK|40|32|Then he brought me to the inner court on the east side, and he measured the gateway; it had the same measurements as the others.
EZEK|40|33|Its alcoves, its projecting walls and its portico had the same measurements as the others. The gateway and its portico had openings all around. It was fifty cubits long and twenty-five cubits wide.
EZEK|40|34|Its portico faced the outer court; palm trees decorated the jambs on either side, and eight steps led up to it.
EZEK|40|35|Then he brought me to the north gate and measured it. It had the same measurements as the others,
EZEK|40|36|as did its alcoves, its projecting walls and its portico, and it had openings all around. It was fifty cubits long and twenty-five cubits wide.
EZEK|40|37|Its portico faced the outer court; palm trees decorated the jambs on either side, and eight steps led up to it.
EZEK|40|38|A room with a doorway was by the portico in each of the inner gateways, where the burnt offerings were washed.
EZEK|40|39|In the portico of the gateway were two tables on each side, on which the burnt offerings, sin offerings and guilt offerings were slaughtered.
EZEK|40|40|By the outside wall of the portico of the gateway, near the steps at the entrance to the north gateway were two tables, and on the other side of the steps were two tables.
EZEK|40|41|So there were four tables on one side of the gateway and four on the other-eight tables in all-on which the sacrifices were slaughtered.
EZEK|40|42|There were also four tables of dressed stone for the burnt offerings, each a cubit and a half long, a cubit and a half wide and a cubit high. On them were placed the utensils for slaughtering the burnt offerings and the other sacrifices.
EZEK|40|43|And double-pronged hooks, each a handbreadth long, were attached to the wall all around. The tables were for the flesh of the offerings.
EZEK|40|44|Outside the inner gate, within the inner court, were two rooms, one at the side of the north gate and facing south, and another at the side of the south gate and facing north.
EZEK|40|45|He said to me, "The room facing south is for the priests who have charge of the temple,
EZEK|40|46|and the room facing north is for the priests who have charge of the altar. These are the sons of Zadok, who are the only Levites who may draw near to the LORD to minister before him."
EZEK|40|47|Then he measured the court: It was square-a hundred cubits long and a hundred cubits wide. And the altar was in front of the temple.
EZEK|40|48|He brought me to the portico of the temple and measured the jambs of the portico; they were five cubits wide on either side. The width of the entrance was fourteen cubits and its projecting walls were three cubits wide on either side.
EZEK|40|49|The portico was twenty cubits wide, and twelve cubits from front to back. It was reached by a flight of stairs, and there were pillars on each side of the jambs.
EZEK|41|1|Then the man brought me to the outer sanctuary and measured the jambs; the width of the jambs was six cubits on each side.
EZEK|41|2|The entrance was ten cubits wide, and the projecting walls on each side of it were five cubits wide. He also measured the outer sanctuary; it was forty cubits long and twenty cubits wide.
EZEK|41|3|Then he went into the inner sanctuary and measured the jambs of the entrance; each was two cubits wide. The entrance was six cubits wide, and the projecting walls on each side of it were seven cubits wide.
EZEK|41|4|And he measured the length of the inner sanctuary; it was twenty cubits, and its width was twenty cubits across the end of the outer sanctuary. He said to me, "This is the Most Holy Place."
EZEK|41|5|Then he measured the wall of the temple; it was six cubits thick, and each side room around the temple was four cubits wide.
EZEK|41|6|The side rooms were on three levels, one above another, thirty on each level. There were ledges all around the wall of the temple to serve as supports for the side rooms, so that the supports were not inserted into the wall of the temple.
EZEK|41|7|The side rooms all around the temple were wider at each successive level. The structure surrounding the temple was built in ascending stages, so that the rooms widened as one went upward. A stairway went up from the lowest floor to the top floor through the middle floor.
EZEK|41|8|I saw that the temple had a raised base all around it, forming the foundation of the side rooms. It was the length of the rod, six long cubits.
EZEK|41|9|The outer wall of the side rooms was five cubits thick. The open area between the side rooms of the temple
EZEK|41|10|and the priests' rooms was twenty cubits wide all around the temple.
EZEK|41|11|There were entrances to the side rooms from the open area, one on the north and another on the south; and the base adjoining the open area was five cubits wide all around.
EZEK|41|12|The building facing the temple courtyard on the west side was seventy cubits wide. The wall of the building was five cubits thick all around, and its length was ninety cubits.
EZEK|41|13|Then he measured the temple; it was a hundred cubits long, and the temple courtyard and the building with its walls were also a hundred cubits long.
EZEK|41|14|The width of the temple courtyard on the east, including the front of the temple, was a hundred cubits.
EZEK|41|15|Then he measured the length of the building facing the courtyard at the rear of the temple, including its galleries on each side; it was a hundred cubits. The outer sanctuary, the inner sanctuary and the portico facing the court,
EZEK|41|16|as well as the thresholds and the narrow windows and galleries around the three of them-everything beyond and including the threshold was covered with wood. The floor, the wall up to the windows, and the windows were covered.
EZEK|41|17|In the space above the outside of the entrance to the inner sanctuary and on the walls at regular intervals all around the inner and outer sanctuary
EZEK|41|18|were carved cherubim and palm trees. Palm trees alternated with cherubim. Each cherub had two faces:
EZEK|41|19|the face of a man toward the palm tree on one side and the face of a lion toward the palm tree on the other. They were carved all around the whole temple.
EZEK|41|20|From the floor to the area above the entrance, cherubim and palm trees were carved on the wall of the outer sanctuary.
EZEK|41|21|The outer sanctuary had a rectangular doorframe, and the one at the front of the Most Holy Place was similar.
EZEK|41|22|There was a wooden altar three cubits high and two cubits square; its corners, its base and its sides were of wood. The man said to me, "This is the table that is before the LORD."
EZEK|41|23|Both the outer sanctuary and the Most Holy Place had double doors.
EZEK|41|24|Each door had two leaves-two hinged leaves for each door.
EZEK|41|25|And on the doors of the outer sanctuary were carved cherubim and palm trees like those carved on the walls, and there was a wooden overhang on the front of the portico.
EZEK|41|26|On the sidewalls of the portico were narrow windows with palm trees carved on each side. The side rooms of the temple also had overhangs.
EZEK|42|1|Then the man led me northward into the outer court and brought me to the rooms opposite the temple courtyard and opposite the outer wall on the north side.
EZEK|42|2|The building whose door faced north was a hundred cubits long and fifty cubits wide.
EZEK|42|3|Both in the section twenty cubits from the inner court and in the section opposite the pavement of the outer court, gallery faced gallery at the three levels.
EZEK|42|4|In front of the rooms was an inner passageway ten cubits wide and a hundred cubits long. Their doors were on the north.
EZEK|42|5|Now the upper rooms were narrower, for the galleries took more space from them than from the rooms on the lower and middle floors of the building.
EZEK|42|6|The rooms on the third floor had no pillars, as the courts had; so they were smaller in floor space than those on the lower and middle floors.
EZEK|42|7|There was an outer wall parallel to the rooms and the outer court; it extended in front of the rooms for fifty cubits.
EZEK|42|8|While the row of rooms on the side next to the outer court was fifty cubits long, the row on the side nearest the sanctuary was a hundred cubits long.
EZEK|42|9|The lower rooms had an entrance on the east side as one enters them from the outer court.
EZEK|42|10|On the south side along the length of the wall of the outer court, adjoining the temple courtyard and opposite the outer wall, were rooms
EZEK|42|11|with a passageway in front of them. These were like the rooms on the north; they had the same length and width, with similar exits and dimensions. Similar to the doorways on the north
EZEK|42|12|were the doorways of the rooms on the south. There was a doorway at the beginning of the passageway that was parallel to the corresponding wall extending eastward, by which one enters the rooms.
EZEK|42|13|Then he said to me, "The north and south rooms facing the temple courtyard are the priests' rooms, where the priests who approach the LORD will eat the most holy offerings. There they will put the most holy offerings-the grain offerings, the sin offerings and the guilt offerings-for the place is holy.
EZEK|42|14|Once the priests enter the holy precincts, they are not to go into the outer court until they leave behind the garments in which they minister, for these are holy. They are to put on other clothes before they go near the places that are for the people."
EZEK|42|15|When he had finished measuring what was inside the temple area, he led me out by the east gate and measured the area all around:
EZEK|42|16|He measured the east side with the measuring rod; it was five hundred cubits.
EZEK|42|17|He measured the north side; it was five hundred cubits by the measuring rod.
EZEK|42|18|He measured the south side; it was five hundred cubits by the measuring rod.
EZEK|42|19|Then he turned to the west side and measured; it was five hundred cubits by the measuring rod.
EZEK|42|20|So he measured the area on all four sides. It had a wall around it, five hundred cubits long and five hundred cubits wide, to separate the holy from the common.
EZEK|43|1|Then the man brought me to the gate facing east,
EZEK|43|2|and I saw the glory of the God of Israel coming from the east. His voice was like the roar of rushing waters, and the land was radiant with his glory.
EZEK|43|3|The vision I saw was like the vision I had seen when he came to destroy the city and like the visions I had seen by the Kebar River, and I fell facedown.
EZEK|43|4|The glory of the LORD entered the temple through the gate facing east.
EZEK|43|5|Then the Spirit lifted me up and brought me into the inner court, and the glory of the LORD filled the temple.
EZEK|43|6|While the man was standing beside me, I heard someone speaking to me from inside the temple.
EZEK|43|7|He said: "Son of man, this is the place of my throne and the place for the soles of my feet. This is where I will live among the Israelites forever. The house of Israel will never again defile my holy name-neither they nor their kings-by their prostitution and the lifeless idols of their kings at their high places.
EZEK|43|8|When they placed their threshold next to my threshold and their doorposts beside my doorposts, with only a wall between me and them, they defiled my holy name by their detestable practices. So I destroyed them in my anger.
EZEK|43|9|Now let them put away from me their prostitution and the lifeless idols of their kings, and I will live among them forever.
EZEK|43|10|"Son of man, describe the temple to the people of Israel, that they may be ashamed of their sins. Let them consider the plan,
EZEK|43|11|and if they are ashamed of all they have done, make known to them the design of the temple-its arrangement, its exits and entrances-its whole design and all its regulations and laws. Write these down before them so that they may be faithful to its design and follow all its regulations.
EZEK|43|12|"This is the law of the temple: All the surrounding area on top of the mountain will be most holy. Such is the law of the temple.
EZEK|43|13|"These are the measurements of the altar in long cubits, that cubit being a cubit and a handbreadth: Its gutter is a cubit deep and a cubit wide, with a rim of one span around the edge. And this is the height of the altar:
EZEK|43|14|From the gutter on the ground up to the lower ledge it is two cubits high and a cubit wide, and from the smaller ledge up to the larger ledge it is four cubits high and a cubit wide.
EZEK|43|15|The altar hearth is four cubits high, and four horns project upward from the hearth.
EZEK|43|16|The altar hearth is square, twelve cubits long and twelve cubits wide.
EZEK|43|17|The upper ledge also is square, fourteen cubits long and fourteen cubits wide, with a rim of half a cubit and a gutter of a cubit all around. The steps of the altar face east."
EZEK|43|18|Then he said to me, "Son of man, this is what the Sovereign LORD says: These will be the regulations for sacrificing burnt offerings and sprinkling blood upon the altar when it is built:
EZEK|43|19|You are to give a young bull as a sin offering to the priests, who are Levites, of the family of Zadok, who come near to minister before me, declares the Sovereign LORD.
EZEK|43|20|You are to take some of its blood and put it on the four horns of the altar and on the four corners of the upper ledge and all around the rim, and so purify the altar and make atonement for it.
EZEK|43|21|You are to take the bull for the sin offering and burn it in the designated part of the temple area outside the sanctuary.
EZEK|43|22|"On the second day you are to offer a male goat without defect for a sin offering, and the altar is to be purified as it was purified with the bull.
EZEK|43|23|When you have finished purifying it, you are to offer a young bull and a ram from the flock, both without defect.
EZEK|43|24|You are to offer them before the LORD, and the priests are to sprinkle salt on them and sacrifice them as a burnt offering to the LORD.
EZEK|43|25|"For seven days you are to provide a male goat daily for a sin offering; you are also to provide a young bull and a ram from the flock, both without defect.
EZEK|43|26|For seven days they are to make atonement for the altar and cleanse it; thus they will dedicate it.
EZEK|43|27|At the end of these days, from the eighth day on, the priests are to present your burnt offerings and fellowship offerings on the altar. Then I will accept you, declares the Sovereign LORD."
EZEK|44|1|Then the man brought me back to the outer gate of the sanctuary, the one facing east, and it was shut.
EZEK|44|2|The LORD said to me, "This gate is to remain shut. It must not be opened; no one may enter through it. It is to remain shut because the LORD, the God of Israel, has entered through it.
EZEK|44|3|The prince himself is the only one who may sit inside the gateway to eat in the presence of the LORD. He is to enter by way of the portico of the gateway and go out the same way."
EZEK|44|4|Then the man brought me by way of the north gate to the front of the temple. I looked and saw the glory of the LORD filling the temple of the LORD, and I fell facedown.
EZEK|44|5|The LORD said to me, "Son of man, look carefully, listen closely and give attention to everything I tell you concerning all the regulations regarding the temple of the LORD. Give attention to the entrance of the temple and all the exits of the sanctuary.
EZEK|44|6|Say to the rebellious house of Israel, 'This is what the Sovereign LORD says: Enough of your detestable practices, O house of Israel!
EZEK|44|7|In addition to all your other detestable practices, you brought foreigners uncircumcised in heart and flesh into my sanctuary, desecrating my temple while you offered me food, fat and blood, and you broke my covenant.
EZEK|44|8|Instead of carrying out your duty in regard to my holy things, you put others in charge of my sanctuary.
EZEK|44|9|This is what the Sovereign LORD says: No foreigner uncircumcised in heart and flesh is to enter my sanctuary, not even the foreigners who live among the Israelites.
EZEK|44|10|"'The Levites who went far from me when Israel went astray and who wandered from me after their idols must bear the consequences of their sin.
EZEK|44|11|They may serve in my sanctuary, having charge of the gates of the temple and serving in it; they may slaughter the burnt offerings and sacrifices for the people and stand before the people and serve them.
EZEK|44|12|But because they served them in the presence of their idols and made the house of Israel fall into sin, therefore I have sworn with uplifted hand that they must bear the consequences of their sin, declares the Sovereign LORD.
EZEK|44|13|They are not to come near to serve me as priests or come near any of my holy things or my most holy offerings; they must bear the shame of their detestable practices.
EZEK|44|14|Yet I will put them in charge of the duties of the temple and all the work that is to be done in it.
EZEK|44|15|"'But the priests, who are Levites and descendants of Zadok and who faithfully carried out the duties of my sanctuary when the Israelites went astray from me, are to come near to minister before me; they are to stand before me to offer sacrifices of fat and blood, declares the Sovereign LORD.
EZEK|44|16|They alone are to enter my sanctuary; they alone are to come near my table to minister before me and perform my service.
EZEK|44|17|"'When they enter the gates of the inner court, they are to wear linen clothes; they must not wear any woolen garment while ministering at the gates of the inner court or inside the temple.
EZEK|44|18|They are to wear linen turbans on their heads and linen undergarments around their waists. They must not wear anything that makes them perspire.
EZEK|44|19|When they go out into the outer court where the people are, they are to take off the clothes they have been ministering in and are to leave them in the sacred rooms, and put on other clothes, so that they do not consecrate the people by means of their garments.
EZEK|44|20|"'They must not shave their heads or let their hair grow long, but they are to keep the hair of their heads trimmed.
EZEK|44|21|No priest is to drink wine when he enters the inner court.
EZEK|44|22|They must not marry widows or divorced women; they may marry only virgins of Israelite descent or widows of priests.
EZEK|44|23|They are to teach my people the difference between the holy and the common and show them how to distinguish between the unclean and the clean.
EZEK|44|24|"'In any dispute, the priests are to serve as judges and decide it according to my ordinances. They are to keep my laws and my decrees for all my appointed feasts, and they are to keep my Sabbaths holy.
EZEK|44|25|"'A priest must not defile himself by going near a dead person; however, if the dead person was his father or mother, son or daughter, brother or unmarried sister, then he may defile himself.
EZEK|44|26|After he is cleansed, he must wait seven days.
EZEK|44|27|On the day he goes into the inner court of the sanctuary to minister in the sanctuary, he is to offer a sin offering for himself, declares the Sovereign LORD.
EZEK|44|28|"'I am to be the only inheritance the priests have. You are to give them no possession in Israel; I will be their possession.
EZEK|44|29|They will eat the grain offerings, the sin offerings and the guilt offerings; and everything in Israel devoted to the LORD will belong to them.
EZEK|44|30|The best of all the firstfruits and of all your special gifts will belong to the priests. You are to give them the first portion of your ground meal so that a blessing may rest on your household.
EZEK|44|31|The priests must not eat anything, bird or animal, found dead or torn by wild animals.
EZEK|45|1|"'When you allot the land as an inheritance, you are to present to the LORD a portion of the land as a sacred district, 25,000 cubits long and 20,000 cubits wide; the entire area will be holy.
EZEK|45|2|Of this, a section 500 cubits square is to be for the sanctuary, with 50 cubits around it for open land.
EZEK|45|3|In the sacred district, measure off a section 25,000 cubits long and 10,000 cubits wide. In it will be the sanctuary, the Most Holy Place.
EZEK|45|4|It will be the sacred portion of the land for the priests, who minister in the sanctuary and who draw near to minister before the LORD. It will be a place for their houses as well as a holy place for the sanctuary.
EZEK|45|5|An area 25,000 cubits long and 10,000 cubits wide will belong to the Levites, who serve in the temple, as their possession for towns to live in.
EZEK|45|6|"'You are to give the city as its property an area 5,000 cubits wide and 25,000 cubits long, adjoining the sacred portion; it will belong to the whole house of Israel.
EZEK|45|7|"'The prince will have the land bordering each side of the area formed by the sacred district and the property of the city. It will extend westward from the west side and eastward from the east side, running lengthwise from the western to the eastern border parallel to one of the tribal portions.
EZEK|45|8|This land will be his possession in Israel. And my princes will no longer oppress my people but will allow the house of Israel to possess the land according to their tribes.
EZEK|45|9|"'This is what the Sovereign LORD says: You have gone far enough, O princes of Israel! Give up your violence and oppression and do what is just and right. Stop dispossessing my people, declares the Sovereign LORD.
EZEK|45|10|You are to use accurate scales, an accurate ephah and an accurate bath.
EZEK|45|11|The ephah and the bath are to be the same size, the bath containing a tenth of a homer and the ephah a tenth of a homer; the homer is to be the standard measure for both.
EZEK|45|12|The shekel is to consist of twenty gerahs. Twenty shekels plus twenty-five shekels plus fifteen shekels equal one mina.
EZEK|45|13|"'This is the special gift you are to offer: a sixth of an ephah from each homer of wheat and a sixth of an ephah from each homer of barley.
EZEK|45|14|The prescribed portion of oil, measured by the bath, is a tenth of a bath from each cor (which consists of ten baths or one homer, for ten baths are equivalent to a homer).
EZEK|45|15|Also one sheep is to be taken from every flock of two hundred from the well-watered pastures of Israel. These will be used for the grain offerings, burnt offerings and fellowship offerings to make atonement for the people, declares the Sovereign LORD.
EZEK|45|16|All the people of the land will participate in this special gift for the use of the prince in Israel.
EZEK|45|17|It will be the duty of the prince to provide the burnt offerings, grain offerings and drink offerings at the festivals, the New Moons and the Sabbaths-at all the appointed feasts of the house of Israel. He will provide the sin offerings, grain offerings, burnt offerings and fellowship offerings to make atonement for the house of Israel.
EZEK|45|18|"'This is what the Sovereign LORD says: In the first month on the first day you are to take a young bull without defect and purify the sanctuary.
EZEK|45|19|The priest is to take some of the blood of the sin offering and put it on the doorposts of the temple, on the four corners of the upper ledge of the altar and on the gateposts of the inner court.
EZEK|45|20|You are to do the same on the seventh day of the month for anyone who sins unintentionally or through ignorance; so you are to make atonement for the temple.
EZEK|45|21|"'In the first month on the fourteenth day you are to observe the Passover, a feast lasting seven days, during which you shall eat bread made without yeast.
EZEK|45|22|On that day the prince is to provide a bull as a sin offering for himself and for all the people of the land.
EZEK|45|23|Every day during the seven days of the Feast he is to provide seven bulls and seven rams without defect as a burnt offering to the LORD, and a male goat for a sin offering.
EZEK|45|24|He is to provide as a grain offering an ephah for each bull and an ephah for each ram, along with a hin of oil for each ephah.
EZEK|45|25|"'During the seven days of the Feast, which begins in the seventh month on the fifteenth day, he is to make the same provision for sin offerings, burnt offerings, grain offerings and oil.
EZEK|46|1|"'This is what the Sovereign LORD says: The gate of the inner court facing east is to be shut on the six working days, but on the Sabbath day and on the day of the New Moon it is to be opened.
EZEK|46|2|The prince is to enter from the outside through the portico of the gateway and stand by the gatepost. The priests are to sacrifice his burnt offering and his fellowship offerings. He is to worship at the threshold of the gateway and then go out, but the gate will not be shut until evening.
EZEK|46|3|On the Sabbaths and New Moons the people of the land are to worship in the presence of the LORD at the entrance to that gateway.
EZEK|46|4|The burnt offering the prince brings to the LORD on the Sabbath day is to be six male lambs and a ram, all without defect.
EZEK|46|5|The grain offering given with the ram is to be an ephah, and the grain offering with the lambs is to be as much as he pleases, along with a hin of oil for each ephah.
EZEK|46|6|On the day of the New Moon he is to offer a young bull, six lambs and a ram, all without defect.
EZEK|46|7|He is to provide as a grain offering one ephah with the bull, one ephah with the ram, and with the lambs as much as he wants to give, along with a hin of oil with each ephah.
EZEK|46|8|When the prince enters, he is to go in through the portico of the gateway, and he is to come out the same way.
EZEK|46|9|"'When the people of the land come before the LORD at the appointed feasts, whoever enters by the north gate to worship is to go out the south gate; and whoever enters by the south gate is to go out the north gate. No one is to return through the gate by which he entered, but each is to go out the opposite gate.
EZEK|46|10|The prince is to be among them, going in when they go in and going out when they go out.
EZEK|46|11|"'At the festivals and the appointed feasts, the grain offering is to be an ephah with a bull, an ephah with a ram, and with the lambs as much as one pleases, along with a hin of oil for each ephah.
EZEK|46|12|When the prince provides a freewill offering to the LORD -whether a burnt offering or fellowship offerings-the gate facing east is to be opened for him. He shall offer his burnt offering or his fellowship offerings as he does on the Sabbath day. Then he shall go out, and after he has gone out, the gate will be shut.
EZEK|46|13|"'Every day you are to provide a year-old lamb without defect for a burnt offering to the LORD; morning by morning you shall provide it.
EZEK|46|14|You are also to provide with it morning by morning a grain offering, consisting of a sixth of an ephah with a third of a hin of oil to moisten the flour. The presenting of this grain offering to the LORD is a lasting ordinance.
EZEK|46|15|So the lamb and the grain offering and the oil shall be provided morning by morning for a regular burnt offering.
EZEK|46|16|"'This is what the Sovereign LORD says: If the prince makes a gift from his inheritance to one of his sons, it will also belong to his descendants; it is to be their property by inheritance.
EZEK|46|17|If, however, he makes a gift from his inheritance to one of his servants, the servant may keep it until the year of freedom; then it will revert to the prince. His inheritance belongs to his sons only; it is theirs.
EZEK|46|18|The prince must not take any of the inheritance of the people, driving them off their property. He is to give his sons their inheritance out of his own property, so that none of my people will be separated from his property.'"
EZEK|46|19|Then the man brought me through the entrance at the side of the gate to the sacred rooms facing north, which belonged to the priests, and showed me a place at the western end.
EZEK|46|20|He said to me, "This is the place where the priests will cook the guilt offering and the sin offering and bake the grain offering, to avoid bringing them into the outer court and consecrating the people."
EZEK|46|21|He then brought me to the outer court and led me around to its four corners, and I saw in each corner another court.
EZEK|46|22|In the four corners of the outer court were enclosed courts, forty cubits long and thirty cubits wide; each of the courts in the four corners was the same size.
EZEK|46|23|Around the inside of each of the four courts was a ledge of stone, with places for fire built all around under the ledge.
EZEK|46|24|He said to me, "These are the kitchens where those who minister at the temple will cook the sacrifices of the people."
EZEK|47|1|The man brought me back to the entrance of the temple, and I saw water coming out from under the threshold of the temple toward the east (for the temple faced east). The water was coming down from under the south side of the temple, south of the altar.
EZEK|47|2|He then brought me out through the north gate and led me around the outside to the outer gate facing east, and the water was flowing from the south side.
EZEK|47|3|As the man went eastward with a measuring line in his hand, he measured off a thousand cubits and then led me through water that was ankle-deep.
EZEK|47|4|He measured off another thousand cubits and led me through water that was knee-deep. He measured off another thousand and led me through water that was up to the waist.
EZEK|47|5|He measured off another thousand, but now it was a river that I could not cross, because the water had risen and was deep enough to swim in-a river that no one could cross.
EZEK|47|6|He asked me, "Son of man, do you see this?" Then he led me back to the bank of the river.
EZEK|47|7|When I arrived there, I saw a great number of trees on each side of the river.
EZEK|47|8|He said to me, "This water flows toward the eastern region and goes down into the Arabah, where it enters the Sea. When it empties into the Sea, the water there becomes fresh.
EZEK|47|9|Swarms of living creatures will live wherever the river flows. There will be large numbers of fish, because this water flows there and makes the salt water fresh; so where the river flows everything will live.
EZEK|47|10|Fishermen will stand along the shore; from En Gedi to En Eglaim there will be places for spreading nets. The fish will be of many kinds-like the fish of the Great Sea.
EZEK|47|11|But the swamps and marshes will not become fresh; they will be left for salt.
EZEK|47|12|Fruit trees of all kinds will grow on both banks of the river. Their leaves will not wither, nor will their fruit fail. Every month they will bear, because the water from the sanctuary flows to them. Their fruit will serve for food and their leaves for healing."
EZEK|47|13|This is what the Sovereign LORD says: "These are the boundaries by which you are to divide the land for an inheritance among the twelve tribes of Israel, with two portions for Joseph.
EZEK|47|14|You are to divide it equally among them. Because I swore with uplifted hand to give it to your forefathers, this land will become your inheritance.
EZEK|47|15|"This is to be the boundary of the land: "On the north side it will run from the Great Sea by the Hethlon road past Lebo Hamath to Zedad,
EZEK|47|16|Berothah and Sibraim (which lies on the border between Damascus and Hamath), as far as Hazer Hatticon, which is on the border of Hauran.
EZEK|47|17|The boundary will extend from the sea to Hazar Enan, along the northern border of Damascus, with the border of Hamath to the north. This will be the north boundary.
EZEK|47|18|"On the east side the boundary will run between Hauran and Damascus, along the Jordan between Gilead and the land of Israel, to the eastern sea and as far as Tamar. This will be the east boundary.
EZEK|47|19|"On the south side it will run from Tamar as far as the waters of Meribah Kadesh, then along the Wadi of Egypt to the Great Sea. This will be the south boundary.
EZEK|47|20|"On the west side, the Great Sea will be the boundary to a point opposite Lebo Hamath. This will be the west boundary.
EZEK|47|21|"You are to distribute this land among yourselves according to the tribes of Israel.
EZEK|47|22|You are to allot it as an inheritance for yourselves and for the aliens who have settled among you and who have children. You are to consider them as native-born Israelites; along with you they are to be allotted an inheritance among the tribes of Israel.
EZEK|47|23|In whatever tribe the alien settles, there you are to give him his inheritance," declares the Sovereign LORD.
EZEK|48|1|"These are the tribes, listed by name: At the northern frontier, Dan will have one portion; it will follow the Hethlon road to Lebo Hamath; Hazar Enan and the northern border of Damascus next to Hamath will be part of its border from the east side to the west side.
EZEK|48|2|"Asher will have one portion; it will border the territory of Dan from east to west.
EZEK|48|3|"Naphtali will have one portion; it will border the territory of Asher from east to west.
EZEK|48|4|"Manasseh will have one portion; it will border the territory of Naphtali from east to west.
EZEK|48|5|"Ephraim will have one portion; it will border the territory of Manasseh from east to west.
EZEK|48|6|"Reuben will have one portion; it will border the territory of Ephraim from east to west.
EZEK|48|7|"Judah will have one portion; it will border the territory of Reuben from east to west.
EZEK|48|8|"Bordering the territory of Judah from east to west will be the portion you are to present as a special gift. It will be 25,000 cubits wide, and its length from east to west will equal one of the tribal portions; the sanctuary will be in the center of it.
EZEK|48|9|"The special portion you are to offer to the LORD will be 25,000 cubits long and 10,000 cubits wide.
EZEK|48|10|This will be the sacred portion for the priests. It will be 25,000 cubits long on the north side, 10,000 cubits wide on the west side, 10,000 cubits wide on the east side and 25,000 cubits long on the south side. In the center of it will be the sanctuary of the LORD.
EZEK|48|11|This will be for the consecrated priests, the Zadokites, who were faithful in serving me and did not go astray as the Levites did when the Israelites went astray.
EZEK|48|12|It will be a special gift to them from the sacred portion of the land, a most holy portion, bordering the territory of the Levites.
EZEK|48|13|"Alongside the territory of the priests, the Levites will have an allotment 25,000 cubits long and 10,000 cubits wide. Its total length will be 25,000 cubits and its width 10,000 cubits.
EZEK|48|14|They must not sell or exchange any of it. This is the best of the land and must not pass into other hands, because it is holy to the LORD.
EZEK|48|15|"The remaining area, 5,000 cubits wide and 25,000 cubits long, will be for the common use of the city, for houses and for pastureland. The city will be in the center of it
EZEK|48|16|and will have these measurements: the north side 4,500 cubits, the south side 4,500 cubits, the east side 4,500 cubits, and the west side 4,500 cubits.
EZEK|48|17|The pastureland for the city will be 250 cubits on the north, 250 cubits on the south, 250 cubits on the east, and 250 cubits on the west.
EZEK|48|18|What remains of the area, bordering on the sacred portion and running the length of it, will be 10,000 cubits on the east side and 10,000 cubits on the west side. Its produce will supply food for the workers of the city.
EZEK|48|19|The workers from the city who farm it will come from all the tribes of Israel.
EZEK|48|20|The entire portion will be a square, 25,000 cubits on each side. As a special gift you will set aside the sacred portion, along with the property of the city.
EZEK|48|21|"What remains on both sides of the area formed by the sacred portion and the city property will belong to the prince. It will extend eastward from the 25,000 cubits of the sacred portion to the eastern border, and westward from the 25,000 cubits to the western border. Both these areas running the length of the tribal portions will belong to the prince, and the sacred portion with the temple sanctuary will be in the center of them.
EZEK|48|22|So the property of the Levites and the property of the city will lie in the center of the area that belongs to the prince. The area belonging to the prince will lie between the border of Judah and the border of Benjamin.
EZEK|48|23|"As for the rest of the tribes: Benjamin will have one portion; it will extend from the east side to the west side.
EZEK|48|24|"Simeon will have one portion; it will border the territory of Benjamin from east to west.
EZEK|48|25|"Issachar will have one portion; it will border the territory of Simeon from east to west.
EZEK|48|26|"Zebulun will have one portion; it will border the territory of Issachar from east to west.
EZEK|48|27|"Gad will have one portion; it will border the territory of Zebulun from east to west.
EZEK|48|28|"The southern boundary of Gad will run south from Tamar to the waters of Meribah Kadesh, then along the Wadi of Egypt to the Great Sea.
EZEK|48|29|"This is the land you are to allot as an inheritance to the tribes of Israel, and these will be their portions," declares the Sovereign LORD.
EZEK|48|30|"These will be the exits of the city: Beginning on the north side, which is 4,500 cubits long,
EZEK|48|31|the gates of the city will be named after the tribes of Israel. The three gates on the north side will be the gate of Reuben, the gate of Judah and the gate of Levi.
EZEK|48|32|"On the east side, which is 4,500 cubits long, will be three gates: the gate of Joseph, the gate of Benjamin and the gate of Dan.
EZEK|48|33|"On the south side, which measures 4,500 cubits, will be three gates: the gate of Simeon, the gate of Issachar and the gate of Zebulun.
EZEK|48|34|"On the west side, which is 4,500 cubits long, will be three gates: the gate of Gad, the gate of Asher and the gate of Naphtali.
EZEK|48|35|"The distance all around will be 18,000 cubits. "And the name of the city from that time on will be: The LORD is There."
