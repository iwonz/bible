SONG|1|1|Solomon's Song of Songs.
SONG|1|2|Let him kiss me with the kisses of his mouth- for your love is more delightful than wine.
SONG|1|3|Pleasing is the fragrance of your perfumes; your name is like perfume poured out. No wonder the maidens love you!
SONG|1|4|Take me away with you-let us hurry! Let the king bring me into his chambers. We rejoice and delight in you; we will praise your love more than wine. How right they are to adore you!
SONG|1|5|Dark am I, yet lovely, O daughters of Jerusalem, dark like the tents of Kedar, like the tent curtains of Solomon.
SONG|1|6|Do not stare at me because I am dark, because I am darkened by the sun. My mother's sons were angry with me and made me take care of the vineyards; my own vineyard I have neglected.
SONG|1|7|Tell me, you whom I love, where you graze your flock and where you rest your sheep at midday. Why should I be like a veiled woman beside the flocks of your friends?
SONG|1|8|If you do not know, most beautiful of women, follow the tracks of the sheep and graze your young goats by the tents of the shepherds.
SONG|1|9|I liken you, my darling, to a mare harnessed to one of the chariots of Pharaoh.
SONG|1|10|Your cheeks are beautiful with earrings, your neck with strings of jewels.
SONG|1|11|We will make you earrings of gold, studded with silver.
SONG|1|12|While the king was at his table, my perfume spread its fragrance.
SONG|1|13|My lover is to me a sachet of myrrh resting between my breasts.
SONG|1|14|My lover is to me a cluster of henna blossoms from the vineyards of En Gedi.
SONG|1|15|How beautiful you are, my darling! Oh, how beautiful! Your eyes are doves.
SONG|1|16|How handsome you are, my lover! Oh, how charming! And our bed is verdant.
SONG|1|17|The beams of our house are cedars; our rafters are firs.
SONG|2|1|I am a rose of Sharon, a lily of the valleys.
SONG|2|2|Like a lily among thorns is my darling among the maidens.
SONG|2|3|Like an apple tree among the trees of the forest is my lover among the young men. I delight to sit in his shade, and his fruit is sweet to my taste.
SONG|2|4|He has taken me to the banquet hall, and his banner over me is love.
SONG|2|5|Strengthen me with raisins, refresh me with apples, for I am faint with love.
SONG|2|6|His left arm is under my head, and his right arm embraces me.
SONG|2|7|Daughters of Jerusalem, I charge you by the gazelles and by the does of the field: Do not arouse or awaken love until it so desires.
SONG|2|8|Listen! My lover! Look! Here he comes, leaping across the mountains, bounding over the hills.
SONG|2|9|My lover is like a gazelle or a young stag. Look! There he stands behind our wall, gazing through the windows, peering through the lattice.
SONG|2|10|My lover spoke and said to me, "Arise, my darling, my beautiful one, and come with me.
SONG|2|11|See! The winter is past; the rains are over and gone.
SONG|2|12|Flowers appear on the earth; the season of singing has come, the cooing of doves is heard in our land.
SONG|2|13|The fig tree forms its early fruit; the blossoming vines spread their fragrance. Arise, come, my darling; my beautiful one, come with me."
SONG|2|14|My dove in the clefts of the rock, in the hiding places on the mountainside, show me your face, let me hear your voice; for your voice is sweet, and your face is lovely.
SONG|2|15|Catch for us the foxes, the little foxes that ruin the vineyards, our vineyards that are in bloom.
SONG|2|16|My lover is mine and I am his; he browses among the lilies.
SONG|2|17|Until the day breaks and the shadows flee, turn, my lover, and be like a gazelle or like a young stag on the rugged hills.
SONG|3|1|All night long on my bed I looked for the one my heart loves; I looked for him but did not find him.
SONG|3|2|I will get up now and go about the city, through its streets and squares; I will search for the one my heart loves. So I looked for him but did not find him.
SONG|3|3|The watchmen found me as they made their rounds in the city. "Have you seen the one my heart loves?"
SONG|3|4|Scarcely had I passed them when I found the one my heart loves. I held him and would not let him go till I had brought him to my mother's house, to the room of the one who conceived me.
SONG|3|5|Daughters of Jerusalem, I charge you by the gazelles and by the does of the field: Do not arouse or awaken love until it so desires.
SONG|3|6|Who is this coming up from the desert like a column of smoke, perfumed with myrrh and incense made from all the spices of the merchant?
SONG|3|7|Look! It is Solomon's carriage, escorted by sixty warriors, the noblest of Israel,
SONG|3|8|all of them wearing the sword, all experienced in battle, each with his sword at his side, prepared for the terrors of the night.
SONG|3|9|King Solomon made for himself the carriage; he made it of wood from Lebanon.
SONG|3|10|Its posts he made of silver, its base of gold. Its seat was upholstered with purple, its interior lovingly inlaid by the daughters of Jerusalem.
SONG|3|11|Come out, you daughters of Zion, and look at King Solomon wearing the crown, the crown with which his mother crowned him on the day of his wedding, the day his heart rejoiced.
SONG|4|1|How beautiful you are, my darling! Oh, how beautiful! Your eyes behind your veil are doves. Your hair is like a flock of goats descending from Mount Gilead.
SONG|4|2|Your teeth are like a flock of sheep just shorn, coming up from the washing. Each has its twin; not one of them is alone.
SONG|4|3|Your lips are like a scarlet ribbon; your mouth is lovely. Your temples behind your veil are like the halves of a pomegranate.
SONG|4|4|Your neck is like the tower of David, built with elegance; on it hang a thousand shields, all of them shields of warriors.
SONG|4|5|Your two breasts are like two fawns, like twin fawns of a gazelle that browse among the lilies.
SONG|4|6|Until the day breaks and the shadows flee, I will go to the mountain of myrrh and to the hill of incense.
SONG|4|7|All beautiful you are, my darling; there is no flaw in you.
SONG|4|8|Come with me from Lebanon, my bride, come with me from Lebanon. Descend from the crest of Amana, from the top of Senir, the summit of Hermon, from the lions' dens and the mountain haunts of the leopards.
SONG|4|9|You have stolen my heart, my sister, my bride; you have stolen my heart with one glance of your eyes, with one jewel of your necklace.
SONG|4|10|How delightful is your love, my sister, my bride! How much more pleasing is your love than wine, and the fragrance of your perfume than any spice!
SONG|4|11|Your lips drop sweetness as the honeycomb, my bride; milk and honey are under your tongue. The fragrance of your garments is like that of Lebanon.
SONG|4|12|You are a garden locked up, my sister, my bride; you are a spring enclosed, a sealed fountain.
SONG|4|13|Your plants are an orchard of pomegranates with choice fruits, with henna and nard,
SONG|4|14|nard and saffron, calamus and cinnamon, with every kind of incense tree, with myrrh and aloes and all the finest spices.
SONG|4|15|You are a garden fountain, a well of flowing water streaming down from Lebanon.
SONG|4|16|Awake, north wind, and come, south wind! Blow on my garden, that its fragrance may spread abroad. Let my lover come into his garden and taste its choice fruits.
SONG|5|1|I have come into my garden, my sister, my bride; I have gathered my myrrh with my spice. I have eaten my honeycomb and my honey; I have drunk my wine and my milk. Eat, O friends, and drink; drink your fill, O lovers.
SONG|5|2|I slept but my heart was awake. Listen! My lover is knocking: "Open to me, my sister, my darling, my dove, my flawless one. My head is drenched with dew, my hair with the dampness of the night."
SONG|5|3|I have taken off my robe- must I put it on again? I have washed my feet- must I soil them again?
SONG|5|4|My lover thrust his hand through the latch-opening; my heart began to pound for him.
SONG|5|5|I arose to open for my lover, and my hands dripped with myrrh, my fingers with flowing myrrh, on the handles of the lock.
SONG|5|6|I opened for my lover, but my lover had left; he was gone. My heart sank at his departure. I looked for him but did not find him. I called him but he did not answer.
SONG|5|7|The watchmen found me as they made their rounds in the city. They beat me, they bruised me; they took away my cloak, those watchmen of the walls!
SONG|5|8|O daughters of Jerusalem, I charge you- if you find my lover, what will you tell him? Tell him I am faint with love.
SONG|5|9|How is your beloved better than others, most beautiful of women? How is your beloved better than others, that you charge us so?
SONG|5|10|My lover is radiant and ruddy, outstanding among ten thousand.
SONG|5|11|His head is purest gold; his hair is wavy and black as a raven.
SONG|5|12|His eyes are like doves by the water streams, washed in milk, mounted like jewels.
SONG|5|13|His cheeks are like beds of spice yielding perfume. His lips are like lilies dripping with myrrh.
SONG|5|14|His arms are rods of gold set with chrysolite. His body is like polished ivory decorated with sapphires.
SONG|5|15|His legs are pillars of marble set on bases of pure gold. His appearance is like Lebanon, choice as its cedars.
SONG|5|16|His mouth is sweetness itself; he is altogether lovely. This is my lover, this my friend, O daughters of Jerusalem.
SONG|6|1|Where has your lover gone, most beautiful of women? Which way did your lover turn, that we may look for him with you?
SONG|6|2|My lover has gone down to his garden, to the beds of spices, to browse in the gardens and to gather lilies.
SONG|6|3|I am my lover's and my lover is mine; he browses among the lilies.
SONG|6|4|You are beautiful, my darling, as Tirzah, lovely as Jerusalem, majestic as troops with banners.
SONG|6|5|Turn your eyes from me; they overwhelm me. Your hair is like a flock of goats descending from Gilead.
SONG|6|6|Your teeth are like a flock of sheep coming up from the washing. Each has its twin, not one of them is alone.
SONG|6|7|Your temples behind your veil are like the halves of a pomegranate.
SONG|6|8|Sixty queens there may be, and eighty concubines, and virgins beyond number;
SONG|6|9|but my dove, my perfect one, is unique, the only daughter of her mother, the favorite of the one who bore her. The maidens saw her and called her blessed; the queens and concubines praised her.
SONG|6|10|Who is this that appears like the dawn, fair as the moon, bright as the sun, majestic as the stars in procession?
SONG|6|11|I went down to the grove of nut trees to look at the new growth in the valley, to see if the vines had budded or the pomegranates were in bloom.
SONG|6|12|Before I realized it, my desire set me among the royal chariots of my people.
SONG|6|13|Come back, come back, O Shulammite; come back, come back, that we may gaze on you! Why would you gaze on the Shulammite as on the dance of Mahanaim?
SONG|7|1|How beautiful your sandaled feet, O prince's daughter! Your graceful legs are like jewels, the work of a craftsman's hands.
SONG|7|2|Your navel is a rounded goblet that never lacks blended wine. Your waist is a mound of wheat encircled by lilies.
SONG|7|3|Your breasts are like two fawns, twins of a gazelle.
SONG|7|4|Your neck is like an ivory tower. Your eyes are the pools of Heshbon by the gate of Bath Rabbim. Your nose is like the tower of Lebanon looking toward Damascus.
SONG|7|5|Your head crowns you like Mount Carmel. Your hair is like royal tapestry; the king is held captive by its tresses.
SONG|7|6|How beautiful you are and how pleasing, O love, with your delights!
SONG|7|7|Your stature is like that of the palm, and your breasts like clusters of fruit.
SONG|7|8|I said, "I will climb the palm tree; I will take hold of its fruit." May your breasts be like the clusters of the vine, the fragrance of your breath like apples,
SONG|7|9|and your mouth like the best wine. May the wine go straight to my lover, flowing gently over lips and teeth.
SONG|7|10|I belong to my lover, and his desire is for me.
SONG|7|11|Come, my lover, let us go to the countryside, let us spend the night in the villages.
SONG|7|12|Let us go early to the vineyards to see if the vines have budded, if their blossoms have opened, and if the pomegranates are in bloom- there I will give you my love.
SONG|7|13|The mandrakes send out their fragrance, and at our door is every delicacy, both new and old, that I have stored up for you, my lover.
SONG|8|1|If only you were to me like a brother, who was nursed at my mother's breasts! Then, if I found you outside, I would kiss you, and no one would despise me.
SONG|8|2|I would lead you and bring you to my mother's house- she who has taught me. I would give you spiced wine to drink, the nectar of my pomegranates.
SONG|8|3|His left arm is under my head and his right arm embraces me.
SONG|8|4|Daughters of Jerusalem, I charge you: Do not arouse or awaken love until it so desires.
SONG|8|5|Who is this coming up from the desert leaning on her lover? Under the apple tree I roused you; there your mother conceived you, there she who was in labor gave you birth.
SONG|8|6|Place me like a seal over your heart, like a seal on your arm; for love is as strong as death, its jealousy unyielding as the grave. It burns like blazing fire, like a mighty flame.
SONG|8|7|Many waters cannot quench love; rivers cannot wash it away. If one were to give all the wealth of his house for love, it would be utterly scorned.
SONG|8|8|We have a young sister, and her breasts are not yet grown. What shall we do for our sister for the day she is spoken for?
SONG|8|9|If she is a wall, we will build towers of silver on her. If she is a door, we will enclose her with panels of cedar.
SONG|8|10|I am a wall, and my breasts are like towers. Thus I have become in his eyes like one bringing contentment.
SONG|8|11|Solomon had a vineyard in Baal Hamon; he let out his vineyard to tenants. Each was to bring for its fruit a thousand shekels of silver.
SONG|8|12|But my own vineyard is mine to give; the thousand shekels are for you, O Solomon, and two hundred are for those who tend its fruit.
SONG|8|13|You who dwell in the gardens with friends in attendance, let me hear your voice!
SONG|8|14|Come away, my lover, and be like a gazelle or like a young stag on the spice-laden mountains.
