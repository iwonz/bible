JOHN|1|1|太初有道，道與上帝同在，道就是上帝。
JOHN|1|2|這道太初與上帝同在。
JOHN|1|3|萬物都是藉著他造的，沒有一樣不是藉著他造的。凡被造的，
JOHN|1|4|在他裏面有生命 ，這生命就是人的光。
JOHN|1|5|光照在黑暗裏，黑暗卻沒有勝過光 。
JOHN|1|6|有一個人，是從上帝那裏差來的，名叫 約翰 。
JOHN|1|7|這人來是為了作見證，是為那光作見證，要使眾人藉著他而信。
JOHN|1|8|他不是那光，而是要為那光作見證。
JOHN|1|9|那光是真光，來到世上，照亮所有的人 。
JOHN|1|10|他在世界，世界是藉著他造的，世界卻不認識他。
JOHN|1|11|他來到自己的地方，自己的人並不接納他。
JOHN|1|12|凡接納他的，就是信他名的人，他就賜他們權柄作上帝的兒女。
JOHN|1|13|這些人不是從血生的，不是從情慾生的，也不是從人的意願生的，而是從上帝生的。
JOHN|1|14|道成了肉身，住在我們中間，充充滿滿地有恩典有真理，我們也見過他的榮光，正是父獨一兒子 的榮光。
JOHN|1|15|約翰 為他作見證，喊著說：「這就是我曾說：『那在我以後來的先於我，因為在我以前，他已經存在。』」
JOHN|1|16|從他的豐富裏，我們都領受了恩典，而且恩上加恩。
JOHN|1|17|律法是藉著 摩西 頒佈的；恩典和真理卻是由耶穌基督來的。
JOHN|1|18|從來沒有人見過上帝，只有在父懷裏獨一的兒子將他表明出來。
JOHN|1|19|這是 約翰 的見證： 猶太 人從 耶路撒冷 差祭司和 利未 人到 約翰 那裏去問他：「你是誰？」
JOHN|1|20|他就承認，並不隱瞞，承認說：「我不是基督。」
JOHN|1|21|他們又問他：「那麼，你是誰？是 以利亞 嗎？」他說：「我不是。」「是那位先知嗎？」他回答：「不是。」
JOHN|1|22|於是他們對他說：「你到底是誰，好讓我們回覆差我們來的人。你說，你自己是誰？」
JOHN|1|23|他說： 「我就是那在曠野呼喊的聲音： 修直主的道。」 正如 以賽亞 先知所說的。
JOHN|1|24|那些人是法利賽人差來的。
JOHN|1|25|他們就問他：「你既不是基督，不是 以利亞 ，也不是那位先知，那麼，你為甚麼施洗呢？」
JOHN|1|26|約翰 回答：「我是用水施洗，但有一位站在你們中間，是你們不認識的，
JOHN|1|27|就是那在我以後來的，我給他解鞋帶也不配。」
JOHN|1|28|這些事發生在 約旦河 東邊的 伯大尼 ， 約翰 施洗的地方。
JOHN|1|29|第二天， 約翰 看見耶穌來到他那裏，就說：「看哪，上帝的羔羊，除去世人的罪的！
JOHN|1|30|這就是我曾說『那在我以後來的先於我，因為在我以前，他已經存在』的那一位。
JOHN|1|31|我先前不認識他，如今我來用水施洗，為要使他顯明給 以色列 人。」
JOHN|1|32|約翰 又作見證說：「我曾看見聖靈彷彿鴿子從天降下，停留在他的身上。
JOHN|1|33|我先前不認識他，可是那差我來用水施洗的對我說：『你看見聖靈降下來，停留在誰的身上，誰就是用聖靈施洗的。』
JOHN|1|34|我看見了，所以作證：這一位是上帝的兒子。」
JOHN|1|35|又過了一天， 約翰 同兩個門徒站在那裏。
JOHN|1|36|他見耶穌走過，就說：「看哪，上帝的羔羊！」
JOHN|1|37|兩個門徒聽見他的話，就跟從了耶穌。
JOHN|1|38|耶穌轉過身來，看見他們跟著，就對他們說：「你們要甚麼？」他們對他說：「拉比，你在哪裏住？」（「拉比」翻出來就是老師。）
JOHN|1|39|耶穌說：「你們來看。」他們就去看他在哪裏住。這一天他們就跟他同住；那時大約是下午四點鐘。
JOHN|1|40|聽了 約翰 的話而跟從耶穌的那兩個人，其中一個是 西門．彼得 的弟弟 安得烈 。
JOHN|1|41|他先找到自己的哥哥 西門 ，對他說：「我們遇見彌賽亞了。」（「彌賽亞」翻出來就是基督。）
JOHN|1|42|於是 安得烈 領 西門 去見耶穌。耶穌看著他，說：「你是 約翰 的兒子 西門 ，你要稱為 磯法 。」（「磯法」翻出來就是 彼得 。）
JOHN|1|43|又過了一天，耶穌想要往 加利利 去。他找到 腓力 ，就對他說：「來跟從我！」
JOHN|1|44|這 腓力 是 伯賽大 人，是 安得烈 和 彼得 的同鄉。
JOHN|1|45|腓力 找到 拿但業 ，對他說：「 摩西 在律法書上所寫的，和眾先知所記的那一位，我們遇見了，就是 約瑟 的兒子 拿撒勒 人耶穌。」
JOHN|1|46|拿但業 對他說：「 拿撒勒 還能出甚麼好的嗎？」 腓力 說：「你來看。」
JOHN|1|47|耶穌看見 拿但業 向他走來，就論到他說：「看哪，這真是個 以色列 人！他心裏是沒有詭詐的。」
JOHN|1|48|拿但業 對耶穌說：「你從哪裏認識我的？」耶穌回答他說：「 腓力 還沒有呼喚你，你在無花果樹底下，我就看見你了。」
JOHN|1|49|拿但業 回答他說：「拉比！你是上帝的兒子，你是 以色列 的王。」
JOHN|1|50|耶穌回答他說：「因為我說在無花果樹底下看見你，你就信嗎？你將看見比這些更大的事呢！」
JOHN|1|51|他又說：「我實實在在地告訴你們，你們將要看見天開了，上帝的使者在人子身上，上去下來。」
JOHN|2|1|第三日，在 加利利 的 迦拿 有一個婚宴，耶穌的母親在那裏。
JOHN|2|2|耶穌和他的門徒也被請去赴宴。
JOHN|2|3|酒用完了，耶穌的母親對他說：「他們沒有酒了。」
JOHN|2|4|耶穌說：「母親 ，我與你何干呢？我的時候還沒有到。」
JOHN|2|5|他母親對用人說：「他告訴你們甚麼，你們就做吧。」
JOHN|2|6|照 猶太 人潔淨禮的規矩，有六口石缸擺在那裏，每口可以盛兩三桶 水。
JOHN|2|7|耶穌對用人說：「把缸倒滿水。」他們就倒滿了，直到缸口。
JOHN|2|8|耶穌又說：「現在舀出來，送給宴會總管。」他們就送了去。
JOHN|2|9|宴會總管嘗了那水變的酒，並不知道是哪裏來的，只有舀水的用人知道。於是宴會總管叫新郎來，
JOHN|2|10|對他說：「人家都是先擺上好酒，等客人喝夠了才擺上次的，你倒把好酒留到現在！」
JOHN|2|11|這是耶穌所行的第一個神蹟，是在 加利利 的 迦拿 行的，顯出了他的榮耀來，他的門徒就信他了。
JOHN|2|12|這事以後，耶穌與他的母親、兄弟 和門徒 都下 迦百農 去，在那裏住了不多幾天。
JOHN|2|13|猶太 人的逾越節近了，耶穌上 耶路撒冷 去。
JOHN|2|14|他看見聖殿裏有賣牛羊和鴿子的，還有兌換銀錢的人坐著，
JOHN|2|15|耶穌就拿繩子做成鞭子，把所有的，包括牛羊都趕出聖殿，倒出兌換銀錢之人的銀錢，推翻他們的桌子，
JOHN|2|16|又對賣鴿子的說：「把這些東西拿走！不要把我父的殿當作買賣的地方。」
JOHN|2|17|他的門徒就想起經上記著：「我為你的殿心裏焦急，如同火燒。」
JOHN|2|18|因此 猶太 領袖問他：「你能顯甚麼神蹟給我們看，表明你可以做這些事呢？」
JOHN|2|19|耶穌回答他們說：「你們拆毀這殿，我三日內要把它重建。」
JOHN|2|20|猶太 人問：「這殿造了四十六年，你三日內就能重建嗎？」
JOHN|2|21|但耶穌所說的殿是指他的身體。
JOHN|2|22|所以他從死人中復活以後，門徒想起他曾說過這事，就信了聖經和耶穌所說的話。
JOHN|2|23|耶穌在 耶路撒冷 過逾越節的時候，有許多人看見他所行的神蹟，就信了他的名。
JOHN|2|24|耶穌自己卻不信任他們，因為他認識所有的人，
JOHN|2|25|也用不著誰來證明人是怎樣的，因為他自己認識人的內心。
JOHN|3|1|有一個法利賽人，名叫 尼哥德慕 ，是 猶太 人的官。
JOHN|3|2|這人夜裏來見耶穌，對他說：「拉比，我們知道你是由上帝那裏來作老師的；因為你所行的神蹟，若沒有上帝同在，無人能行。」
JOHN|3|3|耶穌回答他說：「我實實在在地告訴你，人若不重生 ，就不能見上帝的國。」
JOHN|3|4|尼哥德慕 對他說：「人已經老了，如何能重生呢？豈能再進母腹生出來嗎？」
JOHN|3|5|耶穌回答：「我實實在在地告訴你，人若不是從水和聖靈生的，就不能進上帝的國。
JOHN|3|6|從肉身生的就是肉身；從靈生的就是靈。
JOHN|3|7|我說『你們必須重生』，你不要驚訝。
JOHN|3|8|風 隨著意思吹，你聽見風的聲音，卻不知道是從哪裏來，往哪裏去；凡從聖靈生的也是如此。」
JOHN|3|9|尼哥德慕 問他：「怎麼能有這些事呢？」
JOHN|3|10|耶穌回答，對他說：「你是 以色列 人的老師，還不明白這些事嗎？
JOHN|3|11|我實實在在地告訴你，我們所說的是我們知道的，我們所見證的是我們見過的，你們卻不領受我們的見證。
JOHN|3|12|我對你們說地上的事，你們尚且不信，若對你們說天上的事，如何能信呢？
JOHN|3|13|除了從天降下 的人子，沒有人升過天。
JOHN|3|14|摩西 在曠野怎樣舉蛇，人子也必須照樣被舉起來，
JOHN|3|15|要使一切信他的人都得永生。
JOHN|3|16|「上帝愛世人，甚至將他獨一的兒子 賜給他們，叫一切信他的人不致滅亡，反得永生。
JOHN|3|17|因為上帝差他的兒子到世上來，不是要定世人的罪 ，而是要使世人因他得救。
JOHN|3|18|信他的人不被定罪；不信的人已經被定罪了，因為他不信上帝獨一兒子的名。
JOHN|3|19|光來到世上，世人因自己的行為是惡的，不愛光，倒愛黑暗，這就定了他們的罪。
JOHN|3|20|凡作惡的人都恨惡光，不來接近光，恐怕他的行為被暴露。
JOHN|3|21|但實行真理的人就來接近光，為要顯明他的行為是靠上帝而行的。」
JOHN|3|22|這些事以後，耶穌和門徒到了 猶太 地區，在那裏他和他們同住，並且施洗。
JOHN|3|23|約翰 也在靠近 撒冷 的 哀嫩 施洗，因為那裏水多，眾人都去受洗。
JOHN|3|24|那時 約翰 還沒有下在監裏。
JOHN|3|25|約翰 的門徒和一個 猶太 人辯論潔淨的禮儀，
JOHN|3|26|就來見 約翰 ，對他說：「拉比，從前同你在 約旦河 的東邊，你所見證的那位，你看，他在施洗，眾人都到他那裏去了。」
JOHN|3|27|約翰 回答說：「若不是從天上賜的，人就不能得到甚麼。
JOHN|3|28|你們自己可以為我作見證，我曾說，我不是基督，只是奉差遣在他前面開路的。
JOHN|3|29|娶新娘的是新郎；新郎的朋友站在一旁聽，一聽見新郎的聲音就歡喜快樂。因此，我這喜樂得以滿足了。
JOHN|3|30|他必興旺；我必衰微。」
JOHN|3|31|「從上頭來的是在萬有之上；出於地的是屬於地，他所說的也是屬於地。從天上來的是在萬有之上。
JOHN|3|32|他把所見所聞的見證出來，只是沒有人領受他的見證。
JOHN|3|33|那領受他見證的，就印證上帝是真實的。
JOHN|3|34|上帝所差來的說上帝的話，因為上帝所賜給他的聖靈是沒有限量的。
JOHN|3|35|父愛子，已把萬有交在他手裏。
JOHN|3|36|信子的人有永生；不信子的人得不到永生，而且上帝的憤怒常在他身上。」
JOHN|4|1|耶穌 知道法利賽人聽見他收門徒和施洗比 約翰 還多， （
JOHN|4|2|其實不是耶穌親自施洗，而是他的門徒施洗，）
JOHN|4|3|他就離開 猶太 ，又回 加利利 去。
JOHN|4|4|他必須經過 撒瑪利亞 ，
JOHN|4|5|於是到了 撒瑪利亞 的一座城，名叫 敘加 ，靠近 雅各 給他兒子 約瑟 的那塊地。
JOHN|4|6|雅各井 就在那裏；耶穌因旅途疲乏，坐在井旁。那時約是正午。
JOHN|4|7|有一個 撒瑪利亞 婦人來打水。耶穌對她說：「請給我水喝。」
JOHN|4|8|因為那時門徒進城買食物去了。
JOHN|4|9|撒瑪利亞 婦人對他說：「你是 猶太 人，怎麼向我一個 撒瑪利亞 女人要水喝呢？」因為 猶太 人和 撒瑪利亞 人沒有來往。
JOHN|4|10|耶穌回答她說：「你若知道上帝的恩賜，和對你說『請給我水喝』的是誰，你早就會求他，他也早就會給了你活水。」
JOHN|4|11|婦人對耶穌說：「先生，你沒有打水的器具，井又深，哪裏去取活水呢？
JOHN|4|12|我們的祖宗 雅各 把這井留給我們，他自己和兒女以及牲畜都喝這井裏的水，難道你比他還大嗎？」
JOHN|4|13|耶穌回答，對她說：「凡喝這水的，還要再渴；
JOHN|4|14|誰喝我所賜的水，就永遠不渴。我所賜的水要在他裏面成為泉源，直湧到永生。」
JOHN|4|15|婦人對他說：「先生，請把這水賜給我，使我不渴，也不用到這裏來打水。」
JOHN|4|16|耶穌對她說：「你去，叫你的丈夫，再到這裏來。」
JOHN|4|17|婦人回答，對耶穌說：「我沒有丈夫。」耶穌說：「你說沒有丈夫是對的。
JOHN|4|18|你已經有過五個丈夫，你現在有的並不是你的丈夫。你這話是真的。」
JOHN|4|19|婦人對他說：「先生，我看你是一位先知。
JOHN|4|20|我們的祖宗在這山上敬拜上帝，你們倒說，應當敬拜的地方是在 耶路撒冷 。」
JOHN|4|21|耶穌對她說：「婦人，你要信我。時候將到，你們敬拜父，既不在這山上，也不在 耶路撒冷 。
JOHN|4|22|你們所敬拜的，你們不知道；我們所敬拜的，我們知道，因為救恩是從 猶太 人出來的。
JOHN|4|23|時候將到，現在就是了，那真正敬拜父的，要用心靈和誠實敬拜他，因為父要這樣的人敬拜他。
JOHN|4|24|上帝是靈，所以敬拜他的必須用心靈和誠實敬拜他。」
JOHN|4|25|婦人對他說：「我知道彌賽亞—就是那稱為基督的—要來；他來了，會把一切的事都告訴我們。」
JOHN|4|26|耶穌對她說：「我就是，正在跟你說話呢！」
JOHN|4|27|正在這時，門徒回來了。他們對耶穌正在和一個婦人說話感到驚訝，可是沒有人說：「你要甚麼？」或說：「你為甚麼和她說話？」
JOHN|4|28|那婦人留下水罐，往城裏去，對眾人說：
JOHN|4|29|「你們來看！有一個人把我素來所做的一切事都說了出來，難道這個人就是基督嗎？」
JOHN|4|30|他們就出城，來到耶穌那裏。
JOHN|4|31|就在這個時候，門徒求耶穌說：「拉比，請吃吧。」
JOHN|4|32|耶穌對他們說：「我有食物吃，是你們不知道的。」
JOHN|4|33|門徒就彼此說：「難道有人拿甚麼給他吃了嗎？」
JOHN|4|34|耶穌對他們說：「我的食物就是要遵行差我來那位的旨意，完成他的工作。
JOHN|4|35|你們不是說『到收割的時候還有四個月』嗎？我告訴你們，舉目向田觀看，莊稼熟了，可以收割了。
JOHN|4|36|收割的人已經得工錢 ，為永生儲存五穀，使撒種的和收割的一同快樂。
JOHN|4|37|『那人撒種，這人收割』，這話可見是真的。
JOHN|4|38|我差你們去收你們所沒有辛勞的；別人辛勞，你們享受他們辛勞的成果。」
JOHN|4|39|那城裏有好些 撒瑪利亞 人信了耶穌，因為那婦人作見證，說：「他把我素來所做的一切事都說了出來。」
JOHN|4|40|於是 撒瑪利亞 人來見耶穌，求他在他們那裏住下，他就在那裏住了兩天。
JOHN|4|41|因為耶穌的話，信的人就更多了。
JOHN|4|42|他們對那婦人說：「現在我們信，不再是因為你的話，而是我們親自聽見了，知道這人真是世界的救主。」
JOHN|4|43|過了那兩天，耶穌離開那地方，往 加利利 去。
JOHN|4|44|因為耶穌自己作過見證說：「先知在自己的家鄉是沒有人尊敬的。」
JOHN|4|45|到了 加利利 ， 加利利 人都歡迎他，因為他們也上 耶路撒冷 去過節，曾經看過他在節期間所做的一切事。
JOHN|4|46|耶穌又到了 加利利 的 迦拿 ，就是他從前變水為酒的地方。有一個大臣，他的兒子在 迦百農 病了。
JOHN|4|47|他聽見耶穌從 猶太 到了 加利利 ，就來見他，求他下去醫治他的兒子，因為他兒子快要死了。
JOHN|4|48|耶穌對他說：「若不看見神蹟奇事，你們總是不信。」
JOHN|4|49|那大臣對他說：「先生，求你趁著我的孩子還沒有死就下去吧。」
JOHN|4|50|耶穌對他說：「回去吧，你的兒子會活！」那人信耶穌所說的話，就回去了。
JOHN|4|51|正下去的時候，他的僕人迎面而來，說他的兒子活了。
JOHN|4|52|他就問甚麼時候見好的。他們對他說：「昨天下午一點鐘熱就退了。」
JOHN|4|53|他就知道這正是耶穌對他說「你的兒子會活」的時候；他自己和全家就都信了。
JOHN|4|54|這是耶穌從 猶太 回到 加利利 後所行的第二個神蹟。
JOHN|5|1|這些事以後，到了 猶太 人的一個節期，耶穌上 耶路撒冷 去。
JOHN|5|2|在 耶路撒冷 ，靠近 羊門 有一個池子， 希伯來 話叫 畢士大 ，旁邊有五個柱廊；
JOHN|5|3|裏面躺著許多病人，有失明的、瘸腿的、癱瘓的 。
JOHN|5|4|
JOHN|5|5|在那裏有一個人，病了三十八年。
JOHN|5|6|耶穌看見他躺著，知道他病了很久，就問他：「你要痊癒嗎？」
JOHN|5|7|病人回答他：「先生，水動的時候，沒有人把我放在池子裏；我正要去的時候，別人比我先下去了。」
JOHN|5|8|耶穌對他說：「起來，拿起你的褥子走吧！」
JOHN|5|9|那人立刻痊癒，就拿起自己的褥子走了。 那天是安息日，
JOHN|5|10|所以 猶太 人對那被治好了的人說：「今天是安息日，你拿褥子是不合法的。」
JOHN|5|11|他卻回答他們：「那使我痊癒的人對我說：『拿起你的褥子走吧！』」
JOHN|5|12|他們問他：「對你說『拿起褥子走』的是甚麼人？」
JOHN|5|13|那治好了的人不知道那人是誰，因為那裏人很多，耶穌已經躲開了。
JOHN|5|14|後來耶穌在聖殿裏找到他，對他說：「你已經痊癒了，不要再犯罪，免得你的遭遇更壞。」
JOHN|5|15|那人就去告訴 猶太 人，使他痊癒的是耶穌。
JOHN|5|16|所以 猶太 人迫害耶穌，因為他在安息日做了這些事。
JOHN|5|17|耶穌就回答他們：「我父做事直到如今，我也做事。」
JOHN|5|18|為了這緣故， 猶太 人越發想要殺他，因為他不但犯了安息日，而且稱上帝為他的父，把自己和上帝看為同等。
JOHN|5|19|於是耶穌回答，對他們說：「我實實在在地告訴你們，子憑著自己不能做甚麼，惟有看見父所做的，他才做；父所做的事，子也照樣做。
JOHN|5|20|父愛子，將自己所做的一切事指示給他看，還要將比這更大的事給他看，使你們驚訝。
JOHN|5|21|父怎樣叫死人復活，賜他們生命，子也照樣隨自己的意願賜人生命。
JOHN|5|22|父不審判任何人，而是把審判的事全交給子，
JOHN|5|23|為要使人都尊敬子，如同尊敬父一樣。不尊敬子的，就是不尊敬差子來的父。
JOHN|5|24|「我實實在在地告訴你們，那聽我話又信差我來那位的，就有永生，不至於被定罪，而是已經出死入生了。
JOHN|5|25|我實實在在地告訴你們，時候將到，現在就是了，死人要聽見上帝兒子的聲音，聽見的人就要活了。
JOHN|5|26|因為父怎樣自己裏面有生命，也照樣賜給他兒子自己裏面有生命，
JOHN|5|27|並且賜給他施行審判的權柄，因為他是人子。
JOHN|5|28|你們不要對這事感到驚訝，因為時候將到，凡在墳墓裏的，都要聽見他的聲音，
JOHN|5|29|並且要出來：行善的，復活得生命；作惡的，復活被定罪。
JOHN|5|30|「我憑著自己不能做甚麼。我怎麼聽見就怎麼審判，而我的審判是公平的，因為我不尋求自己的意願，只尋求差我來那位的旨意。」
JOHN|5|31|「我若為自己作見證，我的見證就不真。
JOHN|5|32|另有一位為我作見證，我也知道他為我作的見證是真的。
JOHN|5|33|你們曾差人到 約翰 那裏，他為真理作過見證。
JOHN|5|34|其實，我所受的見證不是從人來的；然而，我說這些話是為了使你們得救。
JOHN|5|35|約翰 是點亮的明燈，你們情願因他的光歡欣一時。
JOHN|5|36|但我有比 約翰 更大的見證：父交給我去完成的工作，就是我正在做的，為我作證是父差遣了我。
JOHN|5|37|那差我來的父也為我作了見證。你們從來沒有聽見他的聲音，也沒有看見他的形像。
JOHN|5|38|你們並沒有他的道存在心裏，因為你們不信他所差來的那一位。
JOHN|5|39|你們查考聖經，因你們以為其中有永生；而這經正是為我作見證的。
JOHN|5|40|然而，你們不肯到我這裏來得生命。
JOHN|5|41|「我不接受從人來的榮耀，
JOHN|5|42|但我知道，你們沒有愛上帝的心。
JOHN|5|43|我奉我父的名來了，你們並不接納我；若有別人奉自己的名來，你們倒會接納他。
JOHN|5|44|你們互相受榮耀，卻不尋求從獨一上帝來的榮耀，怎能信我呢？
JOHN|5|45|不要以為我會在父面前告你們；有一位告你們的，就是你們所仰望的 摩西 。
JOHN|5|46|如果你們信 摩西 ，也會信我，因為他寫過關於我的事。
JOHN|5|47|你們若不信他的書，怎能信我的話呢？」
JOHN|6|1|這些事以後，耶穌渡過 加利利海 ，就是 提比哩亞海 。
JOHN|6|2|有一大群人因為看見他在病人身上所行的神蹟，就跟隨他。
JOHN|6|3|耶穌上了山，和門徒一同坐在那裏。
JOHN|6|4|那時 猶太 人的逾越節近了。
JOHN|6|5|耶穌舉目看見一大群人來，就對 腓力 說：「我們到哪裏去買餅給這些人吃呢？」
JOHN|6|6|他說這話是要考驗 腓力 ，他自己原知道要怎樣做。
JOHN|6|7|腓力 回答他：「就是兩百個銀幣的餅也不夠給他們每人吃一點點。」
JOHN|6|8|有一個門徒，就是 西門．彼得 的弟弟 安得烈 ，對耶穌說：
JOHN|6|9|「這裏有一個孩子，帶著五個大麥餅和兩條魚，但是分給這麼多人還算甚麼呢？」
JOHN|6|10|耶穌說：「你們叫大家坐下。」那地方的草多，人們就坐下，男人的數目約有五千。
JOHN|6|11|耶穌拿起餅來，祝謝了，就分給坐著的人，也同樣分了魚，都照他們所要的來分。
JOHN|6|12|他們吃飽後，耶穌對門徒說：「把剩下的碎屑收拾起來，免得糟蹋了。」
JOHN|6|13|他們就把那五個大麥餅的碎屑，就是大家吃剩的，收拾起來，裝滿了十二個籃子。
JOHN|6|14|人們看見耶穌所行的神蹟，就說：「這真是那要到世上來的先知！」
JOHN|6|15|耶穌知道他們要來強迫他作王，就獨自又退到山上去了。
JOHN|6|16|到了晚上，他的門徒下到海邊，
JOHN|6|17|上了船，要過海往 迦百農 去。天已經黑了，耶穌還沒有來到他們那裏。
JOHN|6|18|忽然狂風大作，海浪翻騰。
JOHN|6|19|門徒搖櫓，約行了十里多 ，看見耶穌在海面上走，漸漸靠近了船，他們就害怕。
JOHN|6|20|耶穌對他們說：「是我，不要怕！」
JOHN|6|21|門徒就欣然接他上船，船立刻到了他們所要去的地方。
JOHN|6|22|第二天，留在海的對岸的眾人發覺那裏原來只有一條小船，而且耶穌沒有同他的門徒上船，是門徒自己去的。
JOHN|6|23|另外有幾條從 提比哩亞 來的小船，卻停靠在主祝謝後給他們吃餅的地方附近。
JOHN|6|24|這時眾人見耶穌和門徒都不在那裏，就上了船，往 迦百農 去找耶穌。
JOHN|6|25|他們在海的對岸找到他後，對他說：「拉比，你幾時到這裏來的？」
JOHN|6|26|耶穌回答他們說：「我實實在在地告訴你們，你們找我，並不是因見了神蹟，而是因吃餅吃飽了。
JOHN|6|27|不要為那會壞的食物操勞，而要為那存到永生的食物操勞。這食物是人子要賜給你們的，因為父上帝已印證了。」
JOHN|6|28|於是他們問他：「我們該做甚麼才算是做上帝的工作呢？」
JOHN|6|29|耶穌回答，對他們說：「信上帝所差來的，這就是上帝的工作。」
JOHN|6|30|於是他們對他說：「你行甚麼神蹟，好讓我們看見而信你呢？你到底要做甚麼呢？
JOHN|6|31|我們的祖宗在曠野吃過嗎哪，如經上寫著：『他從天上賜下糧食來給他們吃。』」
JOHN|6|32|於是耶穌對他們說：「我實實在在地告訴你們，那從天上來的糧不是 摩西 賜給你們的，那從天上來的真糧是我父賜給你們的。
JOHN|6|33|因為上帝的糧就是那位從天上降下來，並且賜生命給世界的。」
JOHN|6|34|於是他們對他說：「主啊，請常常把這糧賜給我們！」
JOHN|6|35|耶穌對他們說：「我就是生命的糧。到我這裏來的，絕不飢餓；信我的，永不乾渴。
JOHN|6|36|可是，我告訴過你們，你們已經看見我 ，還是不信。
JOHN|6|37|凡父所賜給我的人，必到我這裏來；到我這裏來的，我總不丟棄他。
JOHN|6|38|因為我從天上降下來，不是要按自己的意願行，而是要遵行差我來那位的旨意。
JOHN|6|39|差我來那位的旨意就是：他所賜給我的，要我一個也不失落，並且在末日使他復活。
JOHN|6|40|因為我父的旨意是要使每一個見了子而信的人得永生，並且在末日我要使他復活。」
JOHN|6|41|猶太 人因為耶穌說「我是從天上降下來的糧」，就私下議論他，
JOHN|6|42|說：「這不是 約瑟 的兒子耶穌嗎？我們豈不認得他的父母嗎？現在他怎麼說『我是從天上降下來的』呢？」
JOHN|6|43|耶穌回答，對他們說：「你們不要彼此私下議論。
JOHN|6|44|若不是差我來的父吸引人，就沒有人能到我這裏來；到我這裏來的，在末日我要使他復活。
JOHN|6|45|在先知書上寫著：『他們都要蒙上帝教導。』凡聽了父的教導而學習的，都到我這裏來。
JOHN|6|46|這不是說有人看見過父，惟獨從上帝來的，他才看見過父。
JOHN|6|47|我實實在在地告訴你們，信的人有永生。
JOHN|6|48|我就是生命的糧。
JOHN|6|49|你們的祖宗在曠野吃過嗎哪，還是死了。
JOHN|6|50|這是從天上降下來的糧，使人吃了就不死。
JOHN|6|51|我就是從天上降下來生命的糧；人若吃這糧，必永遠活著。我為世人的生命所賜下的糧就是我的肉。」
JOHN|6|52|因此， 猶太 人彼此爭論說：「這個人怎能把他的肉給我們吃呢？」
JOHN|6|53|耶穌對他們說：「我實實在在地告訴你們，你們若不吃人子的肉，不喝人子的血，在你們裏面就沒有生命。
JOHN|6|54|吃我肉、喝我血的人就有永生，並且在末日我要使他復活。
JOHN|6|55|我的肉是真正可吃的；我的血是真正可喝的。
JOHN|6|56|吃我肉、喝我血的人常在我裏面，我也常在他裏面。
JOHN|6|57|永生的父怎樣差我來，我又怎樣因父活著，照樣，吃我肉的人也要因我活著。
JOHN|6|58|這是從天上降下來的糧，不像你們的祖宗吃過嗎哪還是死了；吃這糧的人將永遠活著。」
JOHN|6|59|這些話是耶穌在 迦百農 會堂裏教導人的時候說的。
JOHN|6|60|他的門徒中有好些人聽見了，就說：「這話很難，誰聽得進呢？」
JOHN|6|61|耶穌心裏知道門徒為這話私下議論，就對他們說：「這話成了你們的絆腳石嗎？
JOHN|6|62|如果你們看見人子升到他原來所在之處，會怎麼樣呢？
JOHN|6|63|聖靈賜人生命，肉體毫無用處。我對你們所說的話就是靈，就是生命。
JOHN|6|64|可是你們中間有些人不信。」耶穌起初就知道哪些人不信他，哪一個要出賣他。
JOHN|6|65|於是耶穌說：「所以，我對你們說過，若不是蒙我父的恩賜，沒有人能到我這裏來。」
JOHN|6|66|從此，他門徒中有很多退卻了，不再和他同行。
JOHN|6|67|耶穌就對那十二使徒說：「你們也要離開嗎？」
JOHN|6|68|西門．彼得 回答他：「主啊，你有永生之道，我們還跟從誰呢？
JOHN|6|69|我們已經信了，又知道你是上帝的聖者。」
JOHN|6|70|耶穌回答他們：「我不是揀選了你們十二個嗎？但你們中間有一個是魔鬼。」
JOHN|6|71|耶穌這話是指著要出賣他的 加略 人 西門 的兒子 猶大 說的；他本是十二使徒裏的一個。
JOHN|7|1|這些事以後，耶穌周遊 加利利 ，不願在 猶太 往來，因為 猶太 人想要殺他。
JOHN|7|2|這時 猶太 人的住棚節近了。
JOHN|7|3|耶穌的兄弟們對他說：「你離開這裏上 猶太 去吧，好讓你的門徒也看見你所做的事。
JOHN|7|4|因為人要揚名，沒有在隱祕的地方行事的，如果你要做這些事，該把自己顯明給世人看。」
JOHN|7|5|原來連他的兄弟們也不信他。
JOHN|7|6|於是耶穌對他們說：「我的時機還沒有到，你們的時機卻隨時都有。
JOHN|7|7|世人不會恨你們，卻是恨我，因為我指證他們的行為是惡的。
JOHN|7|8|你們上去過節吧！我現在不上去過這節 ，因為我的時機還沒有成熟。」
JOHN|7|9|耶穌說了這些話，仍然留在 加利利 。
JOHN|7|10|但他的兄弟們上去過節以後，他也上去，不是公開去，卻似乎 是祕密地去的。
JOHN|7|11|節期間， 猶太 人尋找耶穌，說：「他在哪裏？」
JOHN|7|12|人群中有許多人對他議論紛紛，另有的說：「他是好人。」有的說：「不，他是迷惑群眾的。」
JOHN|7|13|可是沒有人公開談論他，因為他們怕 猶太 人。
JOHN|7|14|節期已過了一半，耶穌上聖殿去教導人。
JOHN|7|15|猶太 人驚訝地說：「這個人沒有學過，怎麼那樣熟悉經典呢？」
JOHN|7|16|於是耶穌回答他們，說：「我的教導不是我自己的，而是差我來那位的。
JOHN|7|17|人若立志要遵行上帝的旨意，就會知道這教導究竟是出於上帝，還是我憑著自己說的。
JOHN|7|18|憑著自己說的人是尋求自己的榮耀；但那尋求差他來那位的榮耀的人，他是真誠的，在他心裏沒有不義。
JOHN|7|19|摩西 不是傳了律法給你們嗎？你們卻沒有一個人守律法。為甚麼想要殺我呢？」
JOHN|7|20|眾人回答：「你是被鬼附了！誰想要殺你呢？」
JOHN|7|21|耶穌回答，對他們說：「我做了一件事，你們都驚訝。
JOHN|7|22|摩西 傳割禮給你們（其實割禮不是從 摩西 開始，而是從列祖開始的），你們就在安息日給人行割禮。
JOHN|7|23|人若在安息日受割禮，是為了不違背 摩西 的律法，我在安息日使一個人痊癒了，你們就向我發怒嗎？
JOHN|7|24|不要憑外表斷定是非，總要按公平斷定是非。」
JOHN|7|25|於是 耶路撒冷 人中有的說：「這個人不是他們想要殺的嗎？
JOHN|7|26|你看，他還公開講道，他們也不對他說甚麼。難道官長真的認為這是基督嗎？
JOHN|7|27|然而，我們知道這個人從哪裏來；可是基督來的時候，沒有人知道他從哪裏來。」
JOHN|7|28|那時，耶穌在聖殿裏教導人，喊著說：「你們認識我，也知道我從哪裏來；我並不是憑著自己來的。但差我來的那位是真實的，你們不認識他。
JOHN|7|29|我卻認識他，因為我從他那裏來，是他差遣了我。」
JOHN|7|30|於是他們想要捉拿耶穌，只是沒有人下手，因為他的時候還沒有到。
JOHN|7|31|但人群中有好些人信他，他們說：「基督來的時候，他所行的神蹟難道會比這人行的更多嗎？」
JOHN|7|32|法利賽人聽見群眾對耶穌這樣議論紛紛，祭司長和法利賽人就打發聖殿警衛去捉拿他。
JOHN|7|33|於是耶穌說：「我跟你們在一起的時候不會太久了，我要回到那差我來的那裏去。
JOHN|7|34|你們要找我，卻找不到；我所在的地方，你們不能去。」
JOHN|7|35|於是 猶太 人彼此問：「這人要往哪裏去，使我們找不到他呢？難道他要往散居在 希臘 的 猶太 人那裏去教導 希臘 人嗎？
JOHN|7|36|他說『你們要找我，卻找不到；我所在的地方，你們不能去』這話是甚麼意思呢？」
JOHN|7|37|節期的最後一天，就是最隆重的一天，耶穌站著，喊著說：「人若渴了，到我這裏來喝！
JOHN|7|38|信我的人，就如經上所說：『從他腹中將流出活水的江河來。』」
JOHN|7|39|耶穌這話是指信他的人要受聖靈說的；那時還沒有賜下聖靈，因為耶穌還沒有得到榮耀。
JOHN|7|40|眾人聽見這些話，有的說：「這真是那先知。」
JOHN|7|41|另有的說：「這是基督。」但也有的說：「難道基督是出自 加利利 嗎？
JOHN|7|42|經上不是說『基督是 大衛 的後裔，出自 大衛 的本鄉 伯利恆 』嗎？」
JOHN|7|43|於是眾人因耶穌而分裂了。
JOHN|7|44|其中有人要捉拿他，只是沒有人下手。
JOHN|7|45|警衛們回到祭司長和法利賽人那裏。他們對警衛說：「你們為甚麼沒有帶他來呢？」
JOHN|7|46|警衛回答：「從來沒有像他這樣說話的！」
JOHN|7|47|於是法利賽人說：「你們也受了迷惑嗎？
JOHN|7|48|難道官長或法利賽人中有信他的嗎？
JOHN|7|49|但這些不明白律法的眾人是被詛咒的！」
JOHN|7|50|其中有 尼哥德慕 ，就是從前去見過耶穌的，對他們說：
JOHN|7|51|「不先聽本人的口供，查明他所做的事，難道我們的律法還定他的罪嗎？」
JOHN|7|52|他們回答他說：「你也是出自 加利利 嗎？你去查考就知道， 加利利 是不出先知的。」 〔
JOHN|7|53|於是各人都回家去了，
JOHN|8|1|耶穌卻到 橄欖山 去。
JOHN|8|2|清早，他又回到聖殿裏。眾百姓都到他那裏去，他就坐下，教導他們。
JOHN|8|3|文士和法利賽人帶著一個犯姦淫時被捉的女人來，叫她站在當中，
JOHN|8|4|然後對耶穌說：「老師，這女人是正在犯姦淫的時候被捉到的。
JOHN|8|5|摩西 在律法書上命令我們把這樣的女人用石頭打死。那麼，你怎麼說呢？」
JOHN|8|6|他們說這話是要試探耶穌，要抓到控告他的把柄。耶穌卻彎下腰，用指頭在地上寫字。
JOHN|8|7|他們還是不住地問他，耶穌就直起腰來，對他們說：「你們中間誰沒有罪，誰就先拿石頭打她！」
JOHN|8|8|於是他又彎著腰，用指頭在地上寫字。
JOHN|8|9|他們聽見這話，從老的開始，一個一個都走開了，只剩下耶穌一人和那仍然站在中間的女人。
JOHN|8|10|耶穌就直起腰來，對她說：「婦人，那些人在哪裏呢？沒有任何人定你的罪嗎？」
JOHN|8|11|她說：「主啊，沒有。」耶穌說：「我也不定你的罪。去吧！從今以後不要再犯罪了。」〕
JOHN|8|12|耶穌又對眾人說：「我就是世界的光。跟從我的，必不在黑暗裏走，卻要得著生命的光。」
JOHN|8|13|法利賽人對他說：「你是為自己作見證，你的見證不真。」
JOHN|8|14|耶穌回答他們，對他們說：「即使我為自己作見證，我的見證還是真的，因為我知道我從哪裏來，到哪裏去。你們卻不知道我從哪裏來，到哪裏去。
JOHN|8|15|你們是以人的標準來判斷人，我不判斷任何人。
JOHN|8|16|即使我判斷人，我的判斷也是真確的，因為不是我獨自在判斷，而是差我來的父與我一同判斷。
JOHN|8|17|你們的律法也記著說：『兩個人的見證才算為真』。
JOHN|8|18|我是為自己作見證，還有差我來的父也為我作見證。」
JOHN|8|19|於是他們問他：「你的父在哪裏？」耶穌回答：「你們不認識我，也不認識我的父；若是認識我，也會認識我的父。」
JOHN|8|20|這些話是耶穌在聖殿的銀庫房裏教導人的時候說的。當時沒有人捉拿他，因為他的時候還沒有到。
JOHN|8|21|於是耶穌又對他們說：「我去了，你們會找我，而你們會死在自己的罪中；我所去的地方，你們不能去。」
JOHN|8|22|猶太 人說：「他說『我所去的地方，你們不能去』，難道他要自殺嗎？」
JOHN|8|23|耶穌對他們說：「你們是從下面來的，我是從上面來的；你們是屬這世界的，我不是屬這世界的。
JOHN|8|24|所以我對你們說，你們會死在自己的罪中，你們若不信我就是那位，就會死在自己的罪中。」
JOHN|8|25|他們就問他：「你到底是誰？」耶穌對他們說：「我從起初就告訴你們了。
JOHN|8|26|我有許多事要講論你們，判斷你們；但差我來的那位是真實的，我從他那裏所聽見的，就告訴世人。」
JOHN|8|27|他們不明白耶穌是對他們講父的事。
JOHN|8|28|所以耶穌說：「你們舉起人子以後就會知道我就是那位了，並且知道我沒有一件事是憑著自己做的。我說這些話是照著父所教導我的。
JOHN|8|29|差我來的那位與我同在；他沒有撇下我獨自一人，因為我一直行他所喜悅的事。」
JOHN|8|30|耶穌說這些話的時候，有許多人信了他。
JOHN|8|31|耶穌對信他的 猶太 人說：「你們若繼續遵守我的道，就真是我的門徒了。
JOHN|8|32|你們將認識真理，真理會使你們自由。」
JOHN|8|33|他們回答他：「我們是 亞伯拉罕 的後裔，從來沒有作過誰的奴隸，你怎麼說『會使你們自由』呢？」
JOHN|8|34|耶穌回答他們：「我實實在在地告訴你們，所有犯罪的人就是罪的奴隸。
JOHN|8|35|奴隸不能永遠住在家裏；兒子才永遠住在家裏。
JOHN|8|36|所以，上帝的兒子若使你們自由，你們就真正自由了。」
JOHN|8|37|「我知道，你們是 亞伯拉罕 的後裔，你們卻想要殺我，因為你們心裏容不下我的道。
JOHN|8|38|我所說的是在我父那裏看見的；你們所做的是在你們的父那裏聽到的。」
JOHN|8|39|他們回答耶穌：「我們的父是 亞伯拉罕 。」耶穌對他們說：「你們若是 亞伯拉罕 的兒女，就會做 亞伯拉罕 所做的事。
JOHN|8|40|我把在上帝那裏所聽見的真理告訴了你們，現在你們卻想要殺我； 亞伯拉罕 沒有做過這樣的事。
JOHN|8|41|你們是做你們父的工作。」他們就對他說：「我們不是從淫亂生的，我們只有一位父，就是上帝。」
JOHN|8|42|耶穌對他們說：「假如上帝是你們的父，你們會愛我，因為我本是出於上帝，也是從上帝而來，我不是憑著自己來，而是他差我來的。
JOHN|8|43|你們為甚麼不明白我的話呢？無非是你們聽不進我的道。
JOHN|8|44|你們是出於你們的父魔鬼，你們寧願隨著你們父的慾念而行。他從起初就是殺人的，不守真理，因他心裏沒有真理。他說謊是出於自己的本性，因他本來是說謊的，也是說謊者之父。
JOHN|8|45|但是，因為我講真理，你們就不信我。
JOHN|8|46|你們中間誰能指證我有罪呢？既然我講真理，你們為甚麼不信我呢？
JOHN|8|47|出於上帝的，必聽上帝的話；你們不聽，因為你們不是出於上帝。」
JOHN|8|48|猶太 人回答他：「我們說你是 撒瑪利亞 人，並且是被鬼附的，這話不是很對嗎？」
JOHN|8|49|耶穌回答：「我沒有被鬼附的；我尊敬我的父，你們卻不尊敬我。
JOHN|8|50|我不尋求自己的榮耀，但有一位為我尋求榮耀，判斷是非。
JOHN|8|51|我實實在在地告訴你們，人若遵守我的道，就永遠不經歷死亡。」
JOHN|8|52|於是 猶太 人對他說：「現在我們知道你是被鬼附了。 亞伯拉罕 死了，眾先知也死了，你還說：『人若遵守我的道，就永遠不經歷死亡。』
JOHN|8|53|難道你比我們的祖宗 亞伯拉罕 還大嗎？他死了，眾先知也死了，你把自己當作甚麼人呢？」
JOHN|8|54|耶穌回答：「我若榮耀自己，我的榮耀就算不了甚麼；榮耀我的是我的父，就是你們所說的你們的上帝。
JOHN|8|55|你們不認識他，我卻認識他。我若說不認識他，我就是說謊的，像你們一樣；但我認識他，也遵守他的道。
JOHN|8|56|你們的祖宗 亞伯拉罕 歡歡喜喜地仰望我的日子，他看見了，就快樂。」
JOHN|8|57|猶太 人就對他說：「你還沒有五十歲，難道見過 亞伯拉罕 嗎？」
JOHN|8|58|耶穌對他們說：「我實實在在地告訴你們，還沒有 亞伯拉罕 我就存在了。」
JOHN|8|59|於是他們拿石頭要打他，耶穌卻躲開，走出了聖殿。
JOHN|9|1|耶穌往前走的時候，看見一個生來就失明的人。
JOHN|9|2|門徒問耶穌：「拉比，這人生來失明，是誰犯了罪？是這人還是他的父母呢？」
JOHN|9|3|耶穌回答：「既不是這人犯了罪，也不是他的父母，而是要在他身上顯出上帝的作為來。
JOHN|9|4|趁著白日，我們 必須做差我 來的那位的工；黑夜來到，就沒有人能做工了。
JOHN|9|5|我在世上的時候，是世上的光。」
JOHN|9|6|耶穌說了這些話，就吐唾沫在地上，用唾沫和了泥抹在盲人的眼睛上，
JOHN|9|7|對他說：「你到 西羅亞 池子裏去洗。」（ 西羅亞 翻出來就是「奉差遣」。）於是他去，洗了，回來就看見了。
JOHN|9|8|他的鄰舍和素常見他討飯的人，就說：「這不是那從前坐著討飯的人嗎？」
JOHN|9|9|有的說：「是他」；又有的說：「不是，卻是像他。」他自己說：「是我。」
JOHN|9|10|於是他們對他說：「你的眼睛是怎麼開的呢？」
JOHN|9|11|那人回答：「有一個名叫耶穌的，他和了泥抹我的眼睛，對我說：『你到 西羅亞 池子去洗。』我去一洗，就看見了。」
JOHN|9|12|他們對他說：「那個人在哪裏？」他說：「我不知道。」
JOHN|9|13|他們把以前失明的那個人帶到法利賽人那裏。
JOHN|9|14|耶穌和泥開他眼睛的那一天是安息日。
JOHN|9|15|法利賽人又問他是怎麼得看見的。他對他們說：「他把泥抹在我的眼睛上，我一洗，就看見了。」
JOHN|9|16|於是法利賽人中有的說：「這個人不是從上帝來的，因為他不守安息日。」另有的說：「一個罪人怎能行這樣的神蹟呢？」他們之間就產生了分裂。
JOHN|9|17|於是他們又對那盲人說：「他開了你的眼睛，你說他是怎樣的人呢？」他說：「他是個先知。」
JOHN|9|18|猶太 人不信他以前是失明，後來能看見的，等到叫了他的父母來，
JOHN|9|19|問他們說：「這是你們的兒子嗎？你們說他生來是失明的，現在怎麼看見了呢？」
JOHN|9|20|他的父母就回答說：「他是我們的兒子，生來就失明，這是我們知道的。
JOHN|9|21|至於他現在怎麼能看見，我們卻不知道；是誰開了他的眼睛，我們也不知道。他已經是成人，你們問他吧，他自己會說。」
JOHN|9|22|他父母說這些話，是怕 猶太 人，因為 猶太 人已經商定，若有宣認耶穌是基督的，要把他趕出會堂。
JOHN|9|23|因此他父母說「他已經是成人，你們問他吧」。
JOHN|9|24|於是法利賽人第二次叫了那以前失明的人來，對他說：「你要將榮耀歸給上帝，我們知道這人是個罪人。」
JOHN|9|25|那人就回答：「他是不是個罪人，我不知道；有一件事我知道，我本來是失明的，現在我看見了。」
JOHN|9|26|他們就問他：「他給你做了甚麼？是怎麼開了你的眼睛？」
JOHN|9|27|他回答他們：「我已經告訴你們了，你們不聽，為甚麼又要聽呢？難道你們也要作他的門徒嗎？」
JOHN|9|28|他們就罵他：「你是他的門徒，而我們是 摩西 的門徒。
JOHN|9|29|上帝對 摩西 說話是我們知道的，可是這個人，我們不知道他從哪裏來。」
JOHN|9|30|那人回答，對他們說：「他開了我的眼睛，你們竟不知道他從哪裏來，這真是奇怪！
JOHN|9|31|我們知道上帝不聽罪人，惟有敬奉上帝、遵行他旨意的，上帝才聽他。
JOHN|9|32|從創世以來，未曾聽見有人開了生來就失明的人的眼睛。
JOHN|9|33|這人若不是從上帝來的，甚麼也不能做。」
JOHN|9|34|他們回答他說：「你完全是生在罪中的，還要來教訓我們嗎？」於是他們把他趕出去了。
JOHN|9|35|耶穌聽說他們把他趕出去，就找到他，說：「你信人子 嗎？」
JOHN|9|36|那人回答說：「主啊，人子是誰？告訴我，好讓我信他。」
JOHN|9|37|耶穌對他說：「你已經看見他，現在和你說話的就是他。」
JOHN|9|38|他說：「主啊，我信！」他就拜耶穌。
JOHN|9|39|耶穌說：「我為審判到這世上來，使不能看見的看見，能看見的反而失明。」
JOHN|9|40|同他在那裏的法利賽人聽見這些話，就對他說：「難道我們也失明了嗎？」
JOHN|9|41|耶穌對他們說：「你們若是失明的，就沒有罪了；但現在你們說『我們能看見』，你們的罪還在。」
JOHN|10|1|「我實實在在地告訴你們，那不從門進羊圈，倒從別處爬進去的，就是賊，就是強盜。
JOHN|10|2|那從門進去的才是羊的牧人。
JOHN|10|3|看門的給他開門，羊也聽他的聲音。他按著名叫自己的羊，把羊領出來。
JOHN|10|4|當他把自己的羊都放出來，就走在前面，羊也跟著他，因為牠們認得他的聲音。
JOHN|10|5|羊絕不跟陌生人，反而會逃走，因為不認得陌生人的聲音。」
JOHN|10|6|耶穌把這比方告訴他們，但他們不明白他所說的是甚麼。
JOHN|10|7|所以，耶穌又對他們說：「我實實在在地告訴你們，我就是羊的門。
JOHN|10|8|凡在我以前 來的都是賊，是強盜；羊沒有聽從他們。
JOHN|10|9|我就是門，凡從我進來的，必得安全 ，並且可進出，找到草吃。
JOHN|10|10|盜賊來，無非要偷竊，殺害，毀壞；我來了，是要羊得生命，並且得的更豐盛。
JOHN|10|11|「我是好牧人，好牧人為羊捨命。
JOHN|10|12|雇工不是牧人，羊不是他自己的，他一看見狼來，就撇下羊群逃跑；狼抓住羊，把牠們趕散。
JOHN|10|13|雇工逃走，因為他是雇工，對羊毫不關心。
JOHN|10|14|我是好牧人；我認識我的羊，我的羊也認識我，
JOHN|10|15|正如父認識我，我也認識父一樣；並且我為羊捨命。
JOHN|10|16|我另外有羊，不屬這圈裏的，我必須領牠們來，牠們也要聽我的聲音，並且要合成一群，歸一個牧人。
JOHN|10|17|為此，我父愛我，因為我把命捨去，好再取回來。
JOHN|10|18|沒有人奪去我的命，是我自己捨的；我有權捨棄，也有權再取回。這是我從我父所受的命令。」
JOHN|10|19|猶太 人為這些話又起了分裂。
JOHN|10|20|其中有好些人說：「他是被鬼附了，而且瘋了，為甚麼聽他的呢？」
JOHN|10|21|另有的說：「這不是被鬼附的人所說的話。鬼豈能開盲人的眼睛呢？」
JOHN|10|22|那時正是冬天，在 耶路撒冷 有獻殿節。
JOHN|10|23|耶穌在聖殿裏的 所羅門 廊下行走。
JOHN|10|24|猶太 人圍著他，對他說：「你讓我們猶豫不定到幾時呢？你若是基督，就明白地告訴我們。」
JOHN|10|25|耶穌回答他們：「我已經告訴你們，你們卻不信。我奉我父的名所行的事可以為我作見證。
JOHN|10|26|但是你們不信，因為你們不是我的羊。
JOHN|10|27|我的羊聽我的聲音，我認識牠們，牠們也跟從我。
JOHN|10|28|並且，我賜給他們永生；他們永不滅亡，誰也不能從我手裏把他們奪去。
JOHN|10|29|我父所賜給我的比萬有都大 ，誰也不能從我父手裏把他們奪去。
JOHN|10|30|我與父原為一。」
JOHN|10|31|猶太 人又拿起石頭來要打他。
JOHN|10|32|耶穌回應他們：「我做了許多從父那裏來的善事給你們看，你們是為哪一件拿石頭打我呢？」
JOHN|10|33|猶太 人回答他：「我們不是為了善事拿石頭打你，而是為了你說褻瀆的話；因為你是個人，卻把自己當作上帝。」
JOHN|10|34|耶穌回答他們：「你們的律法書上不是寫著『我曾說你們是諸神』嗎？
JOHN|10|35|經上的話是不能廢的；如果那些領受上帝的道的人，上帝尚且稱他們為諸神，
JOHN|10|36|那麼父所分別為聖又差到世上來的那位說『我是上帝的兒子』，你們還對他說『你說褻瀆的話』嗎？
JOHN|10|37|我若不做我父的工作，你們就不必信我；
JOHN|10|38|我若做了，你們即使不信我，也當信這些工作，好讓你們知道並且明白父在我裏面，我也在父裏面。」
JOHN|10|39|於是，他們又要捉拿他，他卻從他們手中逃脫了。
JOHN|10|40|耶穌又往 約旦河 的東邊去，到了 約翰 起初施洗的地方，就住在那裏。
JOHN|10|41|有許多人來到他那裏，說：「 約翰 沒有行過一件神蹟，但 約翰 所說有關這人的一切話都是真的。」
JOHN|10|42|在那裏，許多人信了耶穌。
JOHN|11|1|有一個患病的人，名叫 拉撒路 ，住在 伯大尼 ，就是 馬利亞 和她姐姐 馬大 的村莊。
JOHN|11|2|這 馬利亞 就是那用香膏抹主，又用頭髮擦他腳的；患病的 拉撒路 是她的弟弟。
JOHN|11|3|姊妹兩個就打發人去見耶穌，說：「主啊，你所愛的人病了。」
JOHN|11|4|耶穌聽見後卻說：「這病不至於死，而是為了上帝的榮耀，為要使上帝的兒子藉此得榮耀。」
JOHN|11|5|耶穌素來愛 馬大 和她妹妹，以及 拉撒路 。
JOHN|11|6|他聽見 拉撒路 病了，仍在原地住了兩天，
JOHN|11|7|然後對門徒說：「我們再到 猶太 去吧！」
JOHN|11|8|門徒對他說：「拉比， 猶太 人近來要拿石頭打你，你還再到那裏去嗎？」
JOHN|11|9|耶穌回答：「白天不是有十二小時嗎？人若在白天行走，就不致跌倒，因為他看見這世上的光。
JOHN|11|10|人若在黑夜行走，就會跌倒，因為他沒有光。」
JOHN|11|11|耶穌說了這些話，隨後對他們說：「我們的朋友 拉撒路 睡了，我去叫醒他。」
JOHN|11|12|門徒就說：「主啊，他若睡了，就會好的。」
JOHN|11|13|耶穌說這話是指 拉撒路 死了，他們卻以為他是指通常的睡眠。
JOHN|11|14|於是耶穌就明白地告訴他們：「 拉撒路 死了。
JOHN|11|15|為了你們的緣故，我不在那裏反而歡喜，為要使你們信。現在我們到他那裏去吧。」
JOHN|11|16|於是那稱為 低土馬 的 多馬 對其他的門徒說：「我們也去和他同死吧！」
JOHN|11|17|耶穌到了，知道 拉撒路 在墳墓裏已經四天了。
JOHN|11|18|伯大尼 離 耶路撒冷 不遠，約有六里 路。
JOHN|11|19|有好些 猶太 人來看 馬大 和 馬利亞 ，要為她們弟弟的緣故安慰她們。
JOHN|11|20|馬大 聽見耶穌來了，就出去迎接他； 馬利亞 卻仍然坐在家裏。
JOHN|11|21|馬大 對耶穌說：「主啊，你若早在這裏，我弟弟就不會死了。
JOHN|11|22|我也知道，即使現在，你無論向上帝求甚麼，上帝也必賜給你。」
JOHN|11|23|耶穌對她說：「你弟弟會復活的。」
JOHN|11|24|馬大 對他說：「我知道在末日復活的時候，他會復活。」
JOHN|11|25|耶穌對她說：「復活在我，生命也在我 。信我的人雖然死了，也必復活；
JOHN|11|26|凡活著信我的人必永遠不死。你信這話嗎？」
JOHN|11|27|馬大 對他說：「主啊，是的。我信你是基督，是上帝的兒子，就是那要臨到世界的。」
JOHN|11|28|馬大 說了這話就回去，叫她妹妹 馬利亞 ，私下說：「老師來了，他在叫你。」
JOHN|11|29|馬利亞 聽見了，急忙起來，到耶穌那裏去。
JOHN|11|30|那時，耶穌還沒有進村子，仍在 馬大 迎接他的地方。
JOHN|11|31|那些同 馬利亞 在家裏安慰她的 猶太 人，見她急忙起來，出去，就跟著她，以為她要往墳墓那裏去哭。
JOHN|11|32|馬利亞 到了耶穌那裏，看見他，就俯伏在他腳前，對他說：「主啊，你若早在這裏，我弟弟就不會死了。」
JOHN|11|33|耶穌看見她哭，並看見與她同來的 猶太 人也哭，就心裏悲嘆，又甚憂愁，
JOHN|11|34|就說：「你們把他安放在哪裏？」他們對他說：「主啊，請你來看。」
JOHN|11|35|耶穌哭了。
JOHN|11|36|猶太 人就說：「你看，他多麼愛他！」
JOHN|11|37|其中有人說：「他既然開了盲人的眼睛，難道不能叫這人不死嗎？」
JOHN|11|38|耶穌又心裏悲嘆，來到墳墓前。那墳墓是個穴，有一塊石頭擋著。
JOHN|11|39|耶穌說：「把石頭挪開！」那死者的姐姐 馬大 對他說：「主啊，他現在必定臭了，因為他已經死了四天了。」
JOHN|11|40|耶穌對她說：「我不是對你說過，你若信就必看見上帝的榮耀嗎？」
JOHN|11|41|於是他們把石頭挪開。耶穌舉目望天，說：「父啊，我感謝你，因為你已經聽了我。
JOHN|11|42|我知道你常常聽我，但我說這話是為了周圍站著的眾人，要使他們信是你差了我來的。」
JOHN|11|43|說了這些話，他大聲呼叫說：「 拉撒路 ，出來！」
JOHN|11|44|那死了的人就出來了，手腳都裹著布，臉上包著頭巾。耶穌對他們說：「解開他，讓他走！」
JOHN|11|45|於是來看 馬利亞 的 猶太 人中，有很多人見了耶穌所做的事，就信了他。
JOHN|11|46|但其中也有人去見法利賽人，把耶穌所做的事告訴他們。
JOHN|11|47|祭司長和法利賽人召開議會，說：「這人行好些神蹟，我們怎麼辦呢？
JOHN|11|48|若讓他這樣做，人人都要信他； 羅馬 人也要來毀滅我們的聖殿 和我們的民族。」
JOHN|11|49|其中有一個人，名叫 該亞法 ，那年當大祭司，對他們說：「你們甚麼都不知道，
JOHN|11|50|也不想想，一個人替百姓死，免得整個民族滅亡，這對你們是有利的。」
JOHN|11|51|他這話不是出於自己的意思，而是因他那年當大祭司，所以預言耶穌將為這民族而死。
JOHN|11|52|他不但替這民族死，還要把上帝四散的兒女都聚集起來，合成一群。
JOHN|11|53|從那日起，他們就商議要殺耶穌。
JOHN|11|54|所以，耶穌不再公開在 猶太 人中走動，卻離開那裏，往靠近曠野的鄉間去，到了一座城，名叫 以法蓮 ，就在那裏和門徒住下來。
JOHN|11|55|猶太 人的逾越節近了，有許多人從鄉下上 耶路撒冷 去，要在過節前潔淨自己。
JOHN|11|56|於是他們尋找耶穌，站在聖殿裏彼此說：「你們認為怎樣，他不會來過節吧？」
JOHN|11|57|那時，祭司長和法利賽人早已下令，若有人知道耶穌的下落，就要報告，他們好去捉拿他。
JOHN|12|1|逾越節前六天，耶穌來到 伯大尼 ，就是他使 拉撒路 從死人中復活的地方。
JOHN|12|2|有人在那裏為耶穌預備宴席； 馬大 伺候， 拉撒路 也在同耶穌坐席的人中間。
JOHN|12|3|馬利亞 拿著一斤極貴的純哪噠 香膏，抹耶穌的腳，又用自己頭髮去擦，屋裏充滿了膏的香氣。
JOHN|12|4|有一個門徒，就是那將要出賣耶穌的 加略 人 猶大 ，說：
JOHN|12|5|「為甚麼不把這香膏賣三百個銀幣去賙濟窮人呢？」
JOHN|12|6|他說這話，並不是關心窮人，而是因為他是個賊，又管錢囊，常偷取錢囊中所存的。
JOHN|12|7|耶穌說：「由她吧！她這香膏本是為我的安葬之日留著的。
JOHN|12|8|因為常有窮人和你們在一起，但是你們不常有我。」
JOHN|12|9|有一大群 猶太 人知道耶穌在那裏，就來了，不但是為耶穌的緣故，也是要看耶穌使他從死人中復活的 拉撒路 。
JOHN|12|10|於是眾祭司長商議連 拉撒路 也要殺了，
JOHN|12|11|因為有許多 猶太 人為了 拉撒路 的緣故，開始背離他們，信了耶穌。
JOHN|12|12|第二天，有一大群上來過節的人聽見耶穌要來 耶路撒冷 ，
JOHN|12|13|就拿著棕樹枝出去迎接他，喊著： 「和散那 ， 以色列 的王！ 奉主名來的是應當稱頌的！」
JOHN|12|14|耶穌找到了一匹驢駒，就騎上，如經上所記：
JOHN|12|15|「 錫安 的兒女 啊，不要懼怕！ 看哪，你的王來了； 他騎在驢駒上。」
JOHN|12|16|門徒當初不明白這些事，等到耶穌得了榮耀後才想起這些話是指他寫的，並且人們果然對他做了這些事。
JOHN|12|17|當耶穌呼喚 拉撒路 ，使他從死人中復活出墳墓的時候，同耶穌在那裏的眾人就作見證。
JOHN|12|18|眾人因聽見耶穌行了這神蹟，就去迎接他。
JOHN|12|19|法利賽人彼此說：「你們看，你們一事無成，世人都隨著他去了。」
JOHN|12|20|那時，上來過節禮拜的人中，有幾個 希臘 人。
JOHN|12|21|他們來見 加利利 的 伯賽大 人 腓力 ，請求他說：「先生，我們想見耶穌。」
JOHN|12|22|腓力 去告訴 安得烈 ，然後 安得烈 同 腓力 去告訴耶穌。
JOHN|12|23|耶穌回答他們說：「人子得榮耀的時候到了。
JOHN|12|24|我實實在在地告訴你們，一粒麥子不落在地裏死了，仍舊是一粒；若是死了，就結出許多子粒來。
JOHN|12|25|愛惜自己性命的，就喪失性命；那恨惡自己在這世上的性命的，要保全性命到永生。
JOHN|12|26|若有人服事我，就當跟從我；我在哪裏，服事我的人也要在哪裏；若有人服事我，我父必尊重他。」
JOHN|12|27|「我現在心裏憂愁，我說甚麼才好呢？說『父啊，救我脫離這時候』嗎？但我正是為這時候來的。
JOHN|12|28|父啊，願你榮耀你的名！」於是有聲音從天上來，說：「我已經榮耀了我的名，還要再榮耀。」
JOHN|12|29|站在旁邊的眾人聽見，就說：「打雷了。」另有的說：「有天使對他說話。」
JOHN|12|30|耶穌回答說：「這聲音不是為我，而是為你們來的。
JOHN|12|31|現在正是這世界受審判的時候；現在這世界的統治者要被趕出去。
JOHN|12|32|我從地上被舉起來的時候，我要吸引萬人來歸我。」
JOHN|12|33|耶穌這話是指自己將要怎樣死說的。
JOHN|12|34|眾人就回答他：「我們聽見律法書上說，基督是永存的；你怎麼說，人子必須被舉起來呢？這人子是誰呢？」
JOHN|12|35|耶穌對他們說：「光在你們中間為時不多了，應該趁著有光的時候行走，免得黑暗臨到你們；那在黑暗裏行走的，不知道往何處去。
JOHN|12|36|你們趁著有光，要信從這光，使你們成為光明之子。」 耶穌說了這些話，就離開他們隱藏了。
JOHN|12|37|他雖然在他們面前行了許多神蹟，他們還是不信他。
JOHN|12|38|這是要應驗 以賽亞 先知所說的話： 「主啊，我們所傳的有誰信呢？ 主的膀臂向誰顯露呢？」
JOHN|12|39|他們所以不能信，因為 以賽亞 又說：
JOHN|12|40|「主使他們瞎了眼， 使他們硬了心， 免得他們眼睛看見， 他們心裏明白，回轉過來， 我會醫治他們。」
JOHN|12|41|以賽亞 因看見了他的榮耀，就說了關於他的這話。
JOHN|12|42|雖然如此，官長中卻有好些信他的，只因法利賽人的緣故不敢承認，恐怕被趕出會堂。
JOHN|12|43|這是因他們愛人給的尊榮過於愛上帝給的尊榮。
JOHN|12|44|耶穌喊著說：「信我的人不是信我，而是信差我來的那位。
JOHN|12|45|看見我的，就是看見差我來的那位。
JOHN|12|46|我就是來到世上的光，使凡信我的不住在黑暗裏。
JOHN|12|47|若有人聽見我的話而不遵守，我不審判他，因為我來不是要審判世人，而是要拯救世人。
JOHN|12|48|棄絕我、不領受我話的人自有審判他的；我所講的道在末日要審判他。
JOHN|12|49|因為我沒有憑著自己講，而是差我來的父已經給我命令，叫我說甚麼，講甚麼。
JOHN|12|50|我也知道他的命令就是永生。所以，我講的正是照著父所告訴我的，我就這麼講了。」
JOHN|13|1|逾越節以前，耶穌知道自己離世歸父的時候到了。他一向愛世間屬自己的人，就愛他們到底。
JOHN|13|2|晚餐的時候，魔鬼已把出賣耶穌的意思放在 加略 人 西門 的兒子 猶大 心裏。
JOHN|13|3|耶穌知道父已把萬有交在他手裏，且知道自己是從上帝出來的，又要回到上帝那裏去，
JOHN|13|4|就離席站起來，脫了衣服，拿一條手巾束腰，
JOHN|13|5|隨後把水倒在盆裏，開始洗門徒的腳，並用束腰的手巾擦乾。
JOHN|13|6|到了 西門．彼得 跟前， 彼得 對他說：「主啊，你洗我的腳嗎？」
JOHN|13|7|耶穌回答他說：「我所做的，你現在不知道，但以後會明白。」
JOHN|13|8|彼得 對他說：「你絕對不可以洗我的腳！」耶穌回答他：「我若不洗你，你就與我無份了。」
JOHN|13|9|西門．彼得 對他說：「主啊，不僅是我的腳，連手和頭也要洗！」
JOHN|13|10|耶穌對他說：「凡洗過澡的人不需要再洗，只要把腳一洗，全身就乾淨了。你們是乾淨的，然而不都是乾淨的。」
JOHN|13|11|耶穌已知道要出賣他的是誰，因此說「你們不都是乾淨的」。
JOHN|13|12|耶穌洗完了他們的腳，就穿上衣服，又坐下，對他們說：「我為你們所做的，你們明白嗎？
JOHN|13|13|你們稱呼我老師，稱呼我主，你們說的不錯，我本來就是。
JOHN|13|14|我是你們的主，你們的老師，尚且洗你們的腳，你們也應當彼此洗腳。
JOHN|13|15|我給你們作了榜樣，為要你們照著我為你們所做的去做。
JOHN|13|16|我實實在在地告訴你們，僕人不大於主人；奉差的人也不大於差他的人。
JOHN|13|17|你們既知道這些事，若是去實行就有福了。
JOHN|13|18|我不是指著你們眾人說的，我知道我所揀選的是誰；但是要應驗經上的話：『吃我飯的人 用腳踢我。』
JOHN|13|19|事情還沒有發生，我現在先告訴你們，讓你們到事情發生的時候好信我就是那位。
JOHN|13|20|我實實在在地告訴你們，接納我所差遣的就是接納我；接納我的就是接納差遣我的那位。」
JOHN|13|21|耶穌說了這些話，心裏憂愁，於是明確地說：「我實實在在地告訴你們，你們中間有一個人要出賣我。」
JOHN|13|22|門徒彼此相看，猜不出他說的是誰。
JOHN|13|23|門徒中有一個人，是耶穌所愛的，側身挨近耶穌的胸懷。
JOHN|13|24|西門．彼得 就對這個人示意，要問耶穌是指著誰說的。
JOHN|13|25|於是那人緊靠著耶穌的胸膛，問他：「主啊，是誰呢？」
JOHN|13|26|耶穌回答：「我蘸一點餅給誰，就是誰。」耶穌就蘸了一點餅，遞給 加略 人 西門 的兒子 猶大 。
JOHN|13|27|他接 了那餅以後，撒但就進入他的心。於是耶穌對他說：「你要做的，快做吧！」
JOHN|13|28|同席的人沒有一個知道耶穌為甚麼對他說這話。
JOHN|13|29|有人因 猶大 管錢囊，以為耶穌是對他說「你去買我們過節所需要的東西」，或是叫他拿些甚麼給窮人。
JOHN|13|30|猶大 受 了那點餅以後立刻出去。那時候是夜間了。
JOHN|13|31|猶大 出去後，耶穌說：「如今人子得了榮耀，上帝在人子身上也得了榮耀。
JOHN|13|32|如果上帝因人子得了榮耀 ，上帝也要因自己榮耀人子，並且要立刻榮耀他。
JOHN|13|33|孩子們！我與你們同在的時候不多了；你們會找我，但我所去的地方，你們不能去。這話我曾對 猶太 人說過，現在也照樣對你們說。
JOHN|13|34|我賜給你們一條新命令，乃是叫你們彼此相愛；我怎樣愛你們，你們也要怎樣彼此相愛。
JOHN|13|35|你們若彼此相愛，眾人因此就認出你們是我的門徒了。」
JOHN|13|36|西門．彼得 問耶穌：「主啊，你去哪裏？」耶穌回答：「我所去的地方，你現在不能跟我去，以後卻要跟我去。」
JOHN|13|37|彼得 對他說：「主啊，為甚麼我現在不能跟你去？我願意為你捨命。」
JOHN|13|38|耶穌回答：「你願意為我捨命嗎？我實實在在地告訴你，雞叫以前，你要三次不認我。」
JOHN|14|1|「你們心裏不要憂愁；你們信上帝，也當信我。
JOHN|14|2|在我父的家裏有許多住處；若是沒有，我就早已告訴你們了。我去原是為你們預備地去方。
JOHN|14|3|我若去為你們預備了地方，就必再來接你們到我那裏去，我在哪裏，叫你們也在哪裏。
JOHN|14|4|我往哪裏去，你們知道那條路。」
JOHN|14|5|多馬 對他說：「主啊，我們不知道你去哪裏，怎麼能知道那條路呢？」
JOHN|14|6|耶穌對他說：「我就是道路、真理、生命；若不藉著我，沒有人能到父那裏去。
JOHN|14|7|既然你們認識了我，也會認識我的父。從今以後，你們就認識他，並且已經看見他了。」
JOHN|14|8|腓力 對他說：「主啊，將父顯給我們看，我們就知足了。」
JOHN|14|9|耶穌對他說：「 腓力 ，我與你們在一起這麼久了，你還不認識我嗎？看見我的就是看見了父，你怎麼還說『將父顯給我們看』呢？
JOHN|14|10|我在父裏面，父在我裏面，你不信嗎？我對你們所說的話不是憑著自己說的，而是住在我裏面的父在做他的工作。
JOHN|14|11|你們要信我，我在父裏面，父在我裏面；即使不信，也要因我所做的工作信我。
JOHN|14|12|我實實在在地告訴你們，我所做的工作，信我的人也要做，並且要做得比這些更大，因為我到父那裏去。
JOHN|14|13|你們奉我的名無論求甚麼，我必成全，為了使父因兒子得榮耀。
JOHN|14|14|你們若奉我的名向我求甚麼，我必成全。」
JOHN|14|15|「你們若愛我，就會遵守我的命令。
JOHN|14|16|我要求父，父就賜給你們另外一位保惠師 ，使他永遠與你們同在。
JOHN|14|17|他就是真理的靈，是世人不能接受的。因為他們既看不見他，也不認識他；你們卻認識他，因他常與你們同在，也要在你們裏面。
JOHN|14|18|我不會撇下你們為孤兒，我必到你們這裏來。
JOHN|14|19|再過不久，世人不再看見我，你們卻會看見我，因為我活著，你們也要活著。
JOHN|14|20|到那日，你們就會知道我在父裏面，你們在我裏面，我也在你們裏面。
JOHN|14|21|有了我的命令而又遵守的人，就是愛我的；愛我的人，我父要愛他，我也要愛他，並且要親自向他顯現。」
JOHN|14|22|猶大 （不是 加略 人 猶大 ）問耶穌：「主啊，為甚麼親自向我們顯現，而不向世人顯現呢？」
JOHN|14|23|耶穌回答他說：「凡愛我的人就會遵守我的道，我父也會愛他，並且我們要到他那裏去，與他同住。
JOHN|14|24|不愛我的人就不遵守我的道。你們所聽見的道不是我的，而是差我來之父的。
JOHN|14|25|「我還與你們在一起的時候，已對你們說了這些事。
JOHN|14|26|但保惠師，就是父因我的名所要差來的聖靈，他要把一切的事教導你們，並且要使你們想起我對你們所說的一切話。
JOHN|14|27|我留下平安給你們，我把我的平安賜給你們。我所賜給你們的，不像世人所賜的。你們心裏不要憂愁，也不要膽怯。
JOHN|14|28|你們聽見我對你們說過，我去了還要回到你們這裏來。你們若愛我，就會因我到父那裏去而喜樂，因為父比我大。
JOHN|14|29|現在事情還沒有發生，我預先告訴你們，使你們在事情發生的時候會信。
JOHN|14|30|我不再和你們多說了，因為這世界的統治者將到，他在我身上一無所能。
JOHN|14|31|我這麼做是照著父命令我的，為了讓世人知道我愛父。起來，我們走吧！」
JOHN|15|1|「我就是真葡萄樹，我父是栽培的人。
JOHN|15|2|凡屬我不結果子的枝子，他就剪掉；凡結果子的，他就修剪乾淨，使枝子結果子更多。
JOHN|15|3|現在你們因我講給你們的道已經潔淨了。
JOHN|15|4|你們要常在我裏面，我也常在你們裏面。枝子若不常在葡萄樹上，自己就不能結果子；你們若不常在我裏面，也是這樣。
JOHN|15|5|我就是葡萄樹，你們是枝子。常在我裏面的，我也常在他裏面，這人就多結果子，因為離了我，你們就不能做甚麼。
JOHN|15|6|人若不常在我裏面，就像枝子被丟在外面，枯乾了，人撿起來，扔進火裏燒了。
JOHN|15|7|你們若常在我裏面，我的話也常在你們裏面，凡你們想要的，祈求，就給你們成全。
JOHN|15|8|你們多結果子，我父就因此得榮耀，你們也就是 我的門徒了。
JOHN|15|9|我愛你們，正如父愛我一樣；你們要常在我的愛裏。
JOHN|15|10|你們若遵守我的命令，就會常在我的愛裏，正如我遵守了我父的命令，常在他的愛裏。
JOHN|15|11|「我已對你們說了這些事，是要讓我的喜樂存在你們心裏，並讓你們的喜樂得以滿足。
JOHN|15|12|你們要彼此相愛，像我愛你們一樣，這是我的命令。
JOHN|15|13|人為朋友捨命，人的愛心沒有比這個更大的了。
JOHN|15|14|你們若遵行我所命令的，就是我的朋友。
JOHN|15|15|以後我不再稱你們為僕人，因為僕人不知道主人所做的事；但我稱你們為朋友，因為我從我父所聽見的一切都已經讓你們知道了。
JOHN|15|16|不是你們揀選了我，而是我揀選了你們，並且派你們去結果子，讓你們的果子得以長存，好使你們奉我的名，無論向父求甚麼，他會賜給你們。
JOHN|15|17|我這樣命令你們，是要你們彼此相愛。」
JOHN|15|18|「世人若恨你們，你們要知道，他們在恨你們以前已經恨我了。
JOHN|15|19|你們若屬世界，世界會愛屬自己的；只因你們不屬世界，而是我從世界中揀選了你們，所以世界就恨你們。
JOHN|15|20|你們要記得我對你們說過的話：『僕人不大於主人。』他們若迫害了我，也會迫害你們，他們若遵守了我的話，也會遵守你們的話。
JOHN|15|21|但他們要因我的名向你們做這一切的事，因為他們不認識差我來的那位。
JOHN|15|22|我若沒有來教導他們，他們就沒有罪；但如今他們的罪無可推諉了。
JOHN|15|23|恨我的也恨我的父。
JOHN|15|24|我若沒有在他們中間做過別人未曾做的事，他們就沒有罪；但如今連我與我的父，他們也看見了，也恨惡了。
JOHN|15|25|這是要應驗他們律法上所寫的話：『他們無故地恨我。』
JOHN|15|26|「但我要從父那裏差保惠師來，就是從父出來的那真理的靈，他來的時候要為我作見證。
JOHN|15|27|你們也要作見證，因為你們從起初就與我同在。」
JOHN|16|1|「我對你們說了這些事，是要使你們不至於跌倒。
JOHN|16|2|人要把你們趕出會堂，而且時候將到，凡殺你們的還以為是在事奉上帝。
JOHN|16|3|他們這樣做，是因為沒有認識父，也沒有認識我。
JOHN|16|4|我對你們說了這些事，是要在他們做這些事的時候，你們會想起我對你們說過的話。」 「我起先沒有對你們說這些事，因為我一直與你們同在。
JOHN|16|5|現在我要到差我來的父那裏去，你們中間卻沒有人問我『你去哪裏？』
JOHN|16|6|只因我對你們說了這些事，你們就滿心憂愁。
JOHN|16|7|然而，我把真情告訴你們，我去對你們是有益的。我若不去，保惠師就不會到你們這裏來；我若去，就差他到你們這裏來。
JOHN|16|8|他來的時候，要為罪、為義，為審判，指證世人；
JOHN|16|9|為罪，是因他們不信我；
JOHN|16|10|為義，是因我到父那裏去，你們將不再見到我；
JOHN|16|11|為審判，是因這世界的統治者已受了審判。
JOHN|16|12|「我還有好些事要告訴你們，但你們現在擔當不了 。
JOHN|16|13|但真理的靈來的時候，他要引導你們進入一切真理。因為他不是憑著自己說的，而是把他所聽見的都說出來，並且要把將要來的事向你們傳達。
JOHN|16|14|他要榮耀我，因為他要把從我領受的向你們傳達。
JOHN|16|15|凡父所有的都是我的，所以我說，他要把從我領受的向你們傳達。」
JOHN|16|16|「不久，你們將不再見到我；再過不久，你們還要見到我。」
JOHN|16|17|有幾個門徒彼此說：「他對我們說『不久，你們將不再見到我；再過不久，你們還要見到我』；又說『因我到父那裏去』。這是甚麼意思呢？」
JOHN|16|18|於是門徒說：「他說 『不久』到底是甚麼意思呢？我們不明白他說甚麼。」
JOHN|16|19|耶穌看出他們要問他，就對他們說：「我說『不久，你們將不再見到我；再過不久，你們還要見到我』，你們為這話彼此詢問嗎？
JOHN|16|20|我實實在在地告訴你們，你們將要痛哭，哀號，世人反要歡喜。你們將要憂愁，然而你們的憂愁要變成喜樂。
JOHN|16|21|婦人生產的時候會憂愁，因為她的時候到了；但孩子一生出來，就不再記得那痛苦了，因為歡喜有一個人生在世上了。
JOHN|16|22|你們現在也是憂愁，但我要再見到你們，你們的心就會有喜樂了；這喜樂沒有人能奪去。
JOHN|16|23|到那日，你們甚麼也不會問我了。我實實在在地告訴你們，你們奉我的名無論向父求甚麼，他會賜給你們 。
JOHN|16|24|直到現在，你們沒有奉我的名求甚麼，如今你們求就必得著，使你們的喜樂得以滿足。」
JOHN|16|25|「這些事，我是用比方對你們說的；時候將到，我不再用比方對你們說，而是要把父的事明白地告訴你們。
JOHN|16|26|到那日，你們要奉我的名祈求；我並不對你們說，我要為你們向父祈求。
JOHN|16|27|父自己愛你們，因為你們已經愛我，又信我是從上帝 而來的。
JOHN|16|28|我從父而來，到了世界 ，又離開世界，到父那裏去。」
JOHN|16|29|門徒說：「你看，如今你是明說，不用比方了。
JOHN|16|30|現在我們曉得你凡事都知道，也不需要有人問你；從此我們信你是從上帝而來的。」
JOHN|16|31|耶穌回答他們：「現在你們信了嗎？
JOHN|16|32|看哪，時候將到，其實已經到了，你們要分散，各歸自己的地方，留下我獨自一人；然而我不是獨自一人，因為有父與我同在。
JOHN|16|33|我對你們說了這些事，是要使你們在我裏面有平安。在世上你們有苦難，但你們要有勇氣 ，我已經勝過世界。」
JOHN|17|1|耶穌說了這些話，就舉目望天，說：「父啊，時候到了，願你榮耀你的兒子，使兒子也榮耀你；
JOHN|17|2|因為你曾賜給他權柄掌管凡血肉之軀的，使他把永生賜給你所賜給他的人。
JOHN|17|3|認識你—獨一的真神，並且認識你所差來的耶穌基督，這就是永生。
JOHN|17|4|我在地上已經榮耀你，你交給我做的工作，我已完成了。
JOHN|17|5|父啊，現在求你使我在你面前得榮耀，就是在未有世界以前，我同你享有的榮耀。
JOHN|17|6|「你從世上賜給我的人，我已把你的名顯明給他們。他們本是你的，你把他們賜給我，他們也遵守了你的道。
JOHN|17|7|現在他們知道，你所賜給我的一切都是從你那裏來的；
JOHN|17|8|因為你所賜給我的話，我已經賜給他們，他們也領受了，又確實知道，我是從你出來的，並且信你差了我來。
JOHN|17|9|我為他們祈求，不為世人祈求，卻為你所賜給我的人祈求，因他們本是你的。
JOHN|17|10|凡是我的都是你的，你的也是我的，並且我因他們得了榮耀。
JOHN|17|11|我到你那裏去；我不再留在世上，他們卻在世上。聖父啊，求你因你的名，就是你所賜給我的名，保守他們，使他們像我們一樣合而為一。
JOHN|17|12|我與他們同在的時候，我奉你的名，就是你所賜給我的名，保守了他們，我也護衛了他們；其中除了那滅亡之子，沒有一個滅亡的，好使經上的話得以應驗。
JOHN|17|13|現在我到你那裏去，我在世上說這些話，是要他們心裏充滿了我的喜樂。
JOHN|17|14|我已把你的道賜給他們；世界恨他們，因為他們不屬世界，正如我不屬世界一樣。
JOHN|17|15|我不求你把他們從世上接走，只求你保全他們，使他們脫離那惡者。
JOHN|17|16|他們不屬世界，正如我不屬世界一樣。
JOHN|17|17|求你用真理使他們成聖；你的道就是真理。
JOHN|17|18|你怎樣差我到世上，我也照樣差他們到世上。
JOHN|17|19|我為他們的緣故使自己分別為聖，為要使他們也因真理成聖。
JOHN|17|20|「我不但為這些人祈求，也為那些藉著他們的話信我的人祈求，
JOHN|17|21|使他們都合而為一。正如父你在我裏面，我在你裏面，使他們也在我們裏面，好讓世人信是你差我來的。
JOHN|17|22|你所賜給我的榮耀，我已賜給他們，使他們合而為一，像我們合而為一。
JOHN|17|23|我在他們裏面，你在我裏面，使他們完完全全合而為一，讓世人知道是你差我來的，也知道你愛他們，如同愛我一樣。
JOHN|17|24|父啊，我在哪裏，願你所賜給我的人也同我在哪裏，使他們看見你所賜給我的榮耀，因為創世以前，你已經愛我了。
JOHN|17|25|公義的父啊，世人未曾認識你，我卻認識你，這些人也知道是你差我來的。
JOHN|17|26|我已讓他們認識你的名，還要讓他們認識，好讓你愛我的愛在他們裏面，我也在他們裏面。」
JOHN|18|1|耶穌說了這些話，就同門徒出去，過了 汲淪溪 。在那裏有一個園子，他和門徒進去了。
JOHN|18|2|出賣耶穌的 猶大 也知道那地方，因為耶穌和門徒屢次在那裏聚集。
JOHN|18|3|猶大 領了一隊兵，以及祭司長和法利賽人的聖殿警衛，拿著燈籠、火把和兵器來到園裏。
JOHN|18|4|耶穌知道將要臨到自己的一切事，就出來對他們說：「你們找誰？」
JOHN|18|5|他們回答他：「 拿撒勒 人耶穌。」耶穌對他們說：「我就是。」出賣他的 猶大 也同他們站在一起。
JOHN|18|6|耶穌一對他們說「我就是」，他們就退後，倒在地上。
JOHN|18|7|他又問他們：「你們找誰？」他們說：「 拿撒勒 人耶穌。」
JOHN|18|8|耶穌回答：「我已經告訴你們，我就是。你們若找的是我，就讓這些人走吧。」
JOHN|18|9|這要應驗耶穌說過的話：「你所賜給我的人，我一個也不失落。」
JOHN|18|10|西門．彼得 帶著一把刀，就拔出來，把大祭司的僕人砍了一刀，削掉了他的右耳，那僕人名叫 馬勒古 。
JOHN|18|11|於是耶穌對 彼得 說：「收刀入鞘吧！我父給我的杯，我豈可不喝呢？」
JOHN|18|12|那隊兵、千夫長和 猶太 人的警衛拿住耶穌，把他捆綁了，
JOHN|18|13|先帶到 亞那 面前，因為他是那年的大祭司 該亞法 的岳父。
JOHN|18|14|這 該亞法 就是從前向 猶太 人忠告說「一個人替百姓死是有利的」那個人。
JOHN|18|15|西門．彼得 跟著耶穌，另一個門徒也跟著；那門徒是大祭司所認識的，他就同耶穌進了大祭司的院子。
JOHN|18|16|彼得 卻站在門外。大祭司所認識的那個門徒出來，對看門的使女說了一聲，就領 彼得 進去。
JOHN|18|17|那看門的使女對 彼得 說：「你不也是這人的門徒嗎？」他說：「我不是。」
JOHN|18|18|僕人和警衛因為天冷生了炭火，站在那裏取暖； 彼得 也同他們站著取暖。
JOHN|18|19|於是，大祭司盤問耶穌有關他的門徒和他教導的事。
JOHN|18|20|耶穌回答他：「我一向都是公開地對世人講話，我常在會堂和聖殿裏，就是 猶太 人聚集的地方教導人，我私下並沒有講甚麼。
JOHN|18|21|你為甚麼問我呢？去問那些聽過我講話的人，我所說的，他們都知道。」
JOHN|18|22|耶穌說了這些話，旁邊站著的一個警衛打了他一耳光，說：「你這樣回答大祭司嗎？」
JOHN|18|23|耶穌回答他：「假如我說的不對，你指證不對的地方；假如我說的對，你為甚麼打我呢？」
JOHN|18|24|於是 亞那 把耶穌綁著押解到大祭司 該亞法 那裏。
JOHN|18|25|西門．彼得 正站著取暖，有人對他說：「你不也是他的門徒嗎？」 彼得 不承認，說：「我不是。」
JOHN|18|26|大祭司的一個僕人，是被 彼得 削掉耳朵那人的親屬，說：「我不是看見你同他在園子裏嗎？」
JOHN|18|27|彼得 又不承認，立刻雞就叫了。
JOHN|18|28|他們把耶穌從 該亞法 那裏押解到總督府。那時是清早。他們自己卻不進總督府，恐怕染了污穢，不能吃逾越節的宴席。
JOHN|18|29|於是 彼拉多 出來，到他們那裏，說：「你們告這人是為甚麼事呢？」
JOHN|18|30|他們回答他說：「這人若不作惡，我們就不會把他交給你了。」
JOHN|18|31|彼拉多 對他們說：「你們自己帶他去，按著你們的律法問他吧！」 猶太 人說：「我們沒有殺人的權柄。」
JOHN|18|32|這是要應驗耶穌所說，指自己將要怎樣死的話。
JOHN|18|33|於是 彼拉多 又進了總督府，叫耶穌來，對他說：「你是 猶太 人的王嗎？」
JOHN|18|34|耶穌回答：「這話是你說的，還是別人論到我時對你說的呢？」
JOHN|18|35|彼拉多 回答：「難道我是 猶太 人嗎？你的同胞和祭司長把你交給我。你做了甚麼事呢？」
JOHN|18|36|耶穌回答：「我的國不屬於這世界；我的國若屬於這世界，我的部下就會為我戰鬥，使我不至於被交給 猶太 人。只是我的國不屬於這世界。」
JOHN|18|37|於是 彼拉多 對他說：「那麼，你是王了？」耶穌回答：「是你說我是王。我為此而生，也為此來到世界，為了給真理作見證。凡屬真理的人都聽我的話。」
JOHN|18|38|彼拉多 對他說：「真理是甚麼呢？」 說了這話， 彼拉多 又出來到 猶太 人那裏，對他們說：「我查不出他有甚麼罪狀。
JOHN|18|39|但你們有個規矩，在逾越節要我給你們釋放一個人，你們要我給你們釋放這 猶太 人的王嗎？」
JOHN|18|40|他們又再喊著說：「不要這人！要 巴拉巴 ！」這 巴拉巴 是個強盜。
JOHN|19|1|於是， 彼拉多 命令把耶穌帶去鞭打了。
JOHN|19|2|士兵用荊棘編了冠冕，戴在他頭上，給他穿上紫袍，
JOHN|19|3|又走到他面前，說：「萬歲， 猶太 人的王！」他們就打他耳光。
JOHN|19|4|彼拉多 又出來對眾人說：「看，我帶他出來見你們，讓你們知道我查不出他有甚麼罪狀。」
JOHN|19|5|耶穌出來，戴著荊棘冠冕，穿著紫袍。 彼拉多 對他們說：「看哪，這個人！」
JOHN|19|6|祭司長和聖殿警衛看見他，就喊著說：「釘十字架！釘十字架！」 彼拉多 對他們說：「你們自己把他帶去釘十字架吧！我查不出他有甚麼罪狀。」
JOHN|19|7|猶太 人回答他：「我們有律法，按照律法，他是該死的，因為他自以為是上帝的兒子。」
JOHN|19|8|彼拉多 聽見這話，越發害怕，
JOHN|19|9|又進了總督府，對耶穌說：「你是哪裏來的？」耶穌卻不回答。
JOHN|19|10|於是 彼拉多 對他說：「你不對我說話嗎？難道你不知道我有權柄釋放你，也有權柄把你釘十字架嗎？」
JOHN|19|11|耶穌回答他：「若不是從上頭賜給你的，你就毫無權柄辦我，所以，把我交給你的那人罪更重了。」
JOHN|19|12|從此， 彼拉多 想要釋放耶穌，無奈 猶太 人喊著說：「你若釋放這個人，你就不是凱撒的忠臣 。凡自立為王的就是背叛凱撒。」
JOHN|19|13|彼拉多 聽見這些話，就帶耶穌出來，到了一個地方，叫「鋪華石處」， 希伯來 話叫 厄巴大 ，就在那裏坐堂。
JOHN|19|14|那日是逾越節的預備日，約在正午。 彼拉多 對 猶太 人說：「看哪，你們的王！」
JOHN|19|15|他們就喊著：「除掉他！除掉他！把他釘十字架！」 彼拉多 對他們說：「要我把你們的王釘十字架嗎？」祭司長回答：「除了凱撒，我們沒有王。」
JOHN|19|16|於是 彼拉多 把耶穌交給他們去釘十字架。 他們就把耶穌帶了去。
JOHN|19|17|耶穌背著自己的十字架出來，到了一個地方，名叫「髑髏地」， 希伯來 話叫 各各他 。
JOHN|19|18|他們就在那裏把他釘在十字架上，還有兩個人和他一同被釘，一邊一個，耶穌在中間。
JOHN|19|19|彼拉多 又寫了一個牌子，釘在十字架上，寫的是：「 猶太 人的王， 拿撒勒 人耶穌。」
JOHN|19|20|有許多 猶太 人念這牌子，因為耶穌被釘十字架的地方靠近城，而且牌子是用 希伯來 、 羅馬 、 希臘 三種文字寫的。
JOHN|19|21|猶太 人的祭司長就對 彼拉多 說：「不要寫『 猶太 人的王』，要寫『那人說：我是 猶太 人的王』。」
JOHN|19|22|彼拉多 回答：「我寫了就寫了。」
JOHN|19|23|士兵把耶穌釘在十字架上以後，把他的衣服拿來分為四份，每人一份。他們又拿他的內衣，這件內衣沒有縫，是上下一片織成的。
JOHN|19|24|他們就彼此說：「我們不要撕開，我們抽籤，看是誰的。」這要應驗經上的話說： 「他們分了我的外衣， 為我的內衣抽籤。」 士兵果然做了這些事。
JOHN|19|25|站在耶穌十字架旁邊的，有他的母親、姨母、 革羅罷 的妻子 馬利亞 ，和 抹大拉 的 馬利亞 。
JOHN|19|26|耶穌見母親和他所愛的那門徒站在旁邊，就對母親說：「母親 ，看，你的兒子！」
JOHN|19|27|又對那門徒說：「看，你的母親！」從那刻起，那門徒就接她到自己家裏去了。
JOHN|19|28|這事以後，耶穌知道各樣的事已經成了，為使經上的話應驗，就說：「我渴了。」
JOHN|19|29|有一個盛滿了醋的罐子放在那裏，他們就拿海綿蘸滿了醋，綁在牛膝草上，送到他嘴邊。
JOHN|19|30|耶穌嘗了那醋，說：「成了！」就低下頭，斷了氣 。
JOHN|19|31|因為這日是預備日，又因為那安息日是個大日子， 猶太 人就來求 彼拉多 叫人打斷他們的腿，把他們搬走，免得屍首在安息日留在十字架上。
JOHN|19|32|於是士兵來，把第一個人的腿，和與耶穌同釘的另一個人的腿，都打斷了。
JOHN|19|33|當他們來到耶穌那裏，見他已經死了，就沒有打斷他的腿。
JOHN|19|34|然而有一個士兵拿槍扎他的肋旁，立刻有血和水流出來。
JOHN|19|35|看見這事的人作了見證—他的見證是真的，他知道自己所說的是真的—好讓你們也信。
JOHN|19|36|這些事發生，為要應驗經上的話：「他的骨頭一根也不可折斷。」
JOHN|19|37|另有經文也說：「他們要仰望自己所扎的人。」
JOHN|19|38|這些事以後， 亞利馬太 的 約瑟 來求 彼拉多 ，要把耶穌的身體領去。他是耶穌的門徒，只因怕 猶太 人，就暗地裏作門徒。 彼拉多 准許了，他就把耶穌的身體領走。
JOHN|19|39|尼哥德慕 也來了，就是先前夜裏去見耶穌的那位，他帶著約一百斤的沒藥和沉香。
JOHN|19|40|他們照 猶太 人喪葬的規矩，用細麻布加上香料，把耶穌的身體裹好了。
JOHN|19|41|在耶穌釘十字架的地方有一個園子，園子裏有一座新墓穴，是從來沒有葬過人的。
JOHN|19|42|因為那天是 猶太 人的預備日，而那墳墓又在附近，他們就把耶穌安放在那裏。
JOHN|20|1|七日的第一日清早，天還黑的時候， 抹大拉 的 馬利亞 來到墳墓，看見石頭已從墳墓挪開了，
JOHN|20|2|就跑來見 西門．彼得 和耶穌所愛的那個門徒，對他們說：「有人從墳墓裏把主移走了，我們不知道他們把他放在哪裏。」
JOHN|20|3|彼得 和那門徒就出來，往墳墓去。
JOHN|20|4|兩個人同跑，那門徒比 彼得 跑得快，先到了墳墓，
JOHN|20|5|低頭往裏看，看見細麻布還放在那裏，只是沒有進去。
JOHN|20|6|西門．彼得 隨後也到了，進了墳墓，看見細麻布放在那裏，
JOHN|20|7|又看見耶穌的裹頭巾沒有和細麻布放在一起，是另在一處捲著。
JOHN|20|8|然後先到墳墓的那門徒也進去，他看見就信了。
JOHN|20|9|他們還不明白聖經所說耶穌必須從死人中復活的意思。
JOHN|20|10|於是兩個門徒回自己的住處去了。
JOHN|20|11|馬利亞 卻站在墳墓外面哭。她哭的時候，低頭往墳墓裏看，
JOHN|20|12|看見兩個天使穿著白衣，在安放耶穌身體的地方坐著，一個在頭，一個在腳。
JOHN|20|13|天使對她說：「婦人，你為甚麼哭？」她對他們說：「因為有人把我主移走了，我不知道他們把他放在哪裏。」
JOHN|20|14|說了這些話，她轉過身來，看見耶穌站在那裏，卻不知道他是耶穌。
JOHN|20|15|耶穌問她：「婦人，你為甚麼哭？你找誰？」 馬利亞 以為他是看園子的，就對他說：「先生，若是你把他移了去，請告訴我，你把他放在哪裏，我去把他移回來。」
JOHN|20|16|耶穌對她說：「 馬利亞 。」 馬利亞 轉過身來，用 希伯來 話對他說：「拉波尼！」（「拉波尼」就是老師的意思。）
JOHN|20|17|耶穌對她說：「不要拉住我，因為我還沒有升上去見我的父。你到我弟兄那裏去告訴他們，我要升上去見我的父，也是你們的父，見我的上帝，也是你們的上帝。」
JOHN|20|18|抹大拉 的 馬利亞 就向門徒報信：「我已經看見了主。」她又把主對她說的話告訴他們。
JOHN|20|19|那日（就是七日的第一日）晚上，門徒因怕 猶太 人，所在的地方門都關了。耶穌來，站在當中，對他們說：「願你們平安！」
JOHN|20|20|說了這話，他把手和肋旁給他們看。門徒一看見主就喜樂了。
JOHN|20|21|於是耶穌又對他們說：「願你們平安！父怎樣差遣了我，我也照樣差遣你們。」
JOHN|20|22|說了這話，他向他們吹一口氣，說：「領受聖靈吧！
JOHN|20|23|你們赦免誰的罪，誰的罪就得赦免；你們不赦免誰的罪，誰的罪就不得赦免。」
JOHN|20|24|那十二使徒中，有個叫 低土馬 的 多馬 ，耶穌來的時候，他沒有和他們在一起。
JOHN|20|25|其他的門徒就對他說：「我們已經看見主了。」 多馬 卻對他們說：「除非我看見他手上的釘痕，用我的指頭探入那釘痕，用我的手探入他的肋旁，我絕不信。」
JOHN|20|26|過了八日，門徒又在屋裏， 多馬 也和他們在一起。門都關了，耶穌來，站在當中，說：「願你們平安！」
JOHN|20|27|然後他對 多馬 說：「把你的指頭伸到這裏來，看看我的手；把你的手伸過來，探入我的肋旁。不要疑惑，總要信！」
JOHN|20|28|多馬 回答，對他說：「我的主！我的上帝！」
JOHN|20|29|耶穌對他說：「你因為看見了我才信嗎？那沒有看見卻信的有福了。」
JOHN|20|30|耶穌在他門徒面前另外行了許多神蹟，沒有記錄在這書上。
JOHN|20|31|但記載這些事是要使你們信 耶穌是基督，是上帝的兒子，並且使你們信他，好因著他的名得生命。
JOHN|21|1|這些事以後，耶穌在 提比哩亞 海邊又向門徒顯現。他怎樣顯現記在下面。
JOHN|21|2|西門．彼得 、叫 低土馬 的 多馬 、 加利利 的 迦拿 人 拿但業 、 西庇太 的兩個兒子，和另外兩個門徒，都在一起。
JOHN|21|3|西門．彼得 對他們說：「我打魚去。」他們對他說：「我們也和你一起去。」他們就出去，上了船；那一夜並沒有打著甚麼。
JOHN|21|4|天剛亮的時候，耶穌站在岸上，門徒卻不知道他是耶穌。
JOHN|21|5|耶穌就對他們說：「孩子們！你們有吃的沒有？」他們回答他：「沒有。」
JOHN|21|6|耶穌對他們說：「你們把網撒在船的右邊，就會得到。」於是他們撒下網去，竟拉不上來了，因為魚很多。
JOHN|21|7|耶穌所愛的那門徒對 彼得 說：「是主！」那時 西門．彼得 赤著身子，一聽見是主，就束上外衣，跳進海裏。
JOHN|21|8|其餘的門徒因離岸不遠，約有二百肘，就坐著小船把那網魚拉過來。
JOHN|21|9|他們上了岸，看見那裏有炭火，上面有魚和餅。
JOHN|21|10|耶穌對他們說：「把剛才打的魚拿幾條來。」
JOHN|21|11|西門．彼得 就上船，把網拉到岸上，網裏滿了大魚，共一百五十三條；雖然魚這樣多，網卻沒有破。
JOHN|21|12|耶穌對他們說：「你們來吃早飯。」門徒中沒有一個敢問他：「你是誰？」因為他們知道他是主。
JOHN|21|13|耶穌走過來，拿餅給他們，也照樣拿魚給他們。
JOHN|21|14|耶穌從死人中復活後向門徒顯現，這是第三次。
JOHN|21|15|他們吃完了早飯，耶穌對 西門．彼得 說：「 約翰 的兒子 西門 ，你愛我比這些更深嗎？」 彼得 對他說：「主啊，是的，你知道我愛你。」耶穌對他說：「你餵養我的小羊。」
JOHN|21|16|耶穌第二次又對他說：「 約翰 的兒子 西門 ，你愛我嗎？」 彼得 對他說：「主啊，是的，你知道我愛你。」耶穌說：「你牧養我的羊。」
JOHN|21|17|耶穌第三次對他說：「 約翰 的兒子 西門 ，你愛我嗎？」 彼得 因為耶穌第三次對他說「你愛我嗎」，就憂愁，對耶穌說：「主啊，你無所不知，你知道我愛你。」耶穌說：「你餵養我的羊。
JOHN|21|18|我實實在在地告訴你，你年輕的時候，自己束上帶子，隨意往來；但年老的時候，你要伸出手來，別人要把你束上，帶你到不願意去的地方。」
JOHN|21|19|耶穌說這話，是指 彼得 會怎樣死來榮耀上帝。說了這話，耶穌對他說：「你跟從我吧！」
JOHN|21|20|彼得 轉過身來，看見耶穌所愛的那門徒跟著，就是在晚餐時靠著耶穌胸膛說「主啊，出賣你的是誰」的那門徒。
JOHN|21|21|彼得 看見他，就問耶穌：「主啊，這個人怎樣呢？」
JOHN|21|22|耶穌對他說：「假如我要他等到我來的時候還在，跟你有甚麼關係呢？你跟從我吧！」
JOHN|21|23|於是這話在弟兄中間流傳，說那門徒不死。其實，耶穌不是說他不死，而是對 彼得 說：「假如我要他等到我來的時候還在，跟你有甚麼關係呢？ 」
JOHN|21|24|這門徒就是為這些事作見證、並且記載這些事的，我們知道他的見證是真的。
JOHN|21|25|耶穌所行的事還有許多，若是一一都寫出來，我想，就是全世界也容不下所要寫的書。
