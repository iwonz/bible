HEB|1|1|古时候，上帝藉着众先知多次多方向列祖说话，
HEB|1|2|末世，藉着他儿子向我们说话，又立他为承受万有的，也藉着他创造宇宙。
HEB|1|3|他是上帝荣耀的光辉，是上帝本体的真像，常用他大能的命令托住万有。他洗净了人的罪，就坐在高天至大者的右边。
HEB|1|4|他所承受的名比天使的名更尊贵，所以他远比天使崇高。
HEB|1|5|上帝曾对哪一个天使说过： “你是我的儿子； 我今日生了你”？ 又说过： “我要作他的父； 他要作我的子”呢？
HEB|1|6|再者，上帝引领他长子 进入世界的时候，说： “上帝的使者都要拜他。”
HEB|1|7|关于使者，他说： “上帝以风为使者， 以火焰为仆役。”
HEB|1|8|关于子，他却说： “上帝啊，你的宝座是永永远远的； 你国度的权杖是正直的权杖。
HEB|1|9|你喜爱公义，恨恶罪恶； 所以上帝，就是你的上帝，用喜乐油膏你， 胜过膏你的同伴。”
HEB|1|10|他又说： “主啊，你起初立了地的根基， 天也是你手所造的。
HEB|1|11|天地都会消灭，你却长存； 天地都会像衣服渐渐旧了；
HEB|1|12|你要将天地卷起来，像卷一件外衣， 天地像衣服都会改变。 你却永不改变； 你的年数没有穷尽。”
HEB|1|13|上帝曾对哪一个天使说： “你坐在我的右边， 等我使你的仇敌作你的脚凳”？
HEB|1|14|众天使不都是事奉的灵，奉差遣为那将要承受救恩的人服务的吗？
HEB|2|1|所以，我们必须越发注意所听见的道，免得我们随流失去。
HEB|2|2|既然那藉着天使所传的话是确定的，凡违背不听从的，都受了该受的报应；
HEB|2|3|我们若忽略这么大的救恩，怎能逃避呢？这拯救起先是主亲自讲的，后来是听见的人给我们证实了。
HEB|2|4|上帝又按自己的旨意，更用神迹奇事、百般的异能，和圣灵所给的恩赐，与他们一同作见证。
HEB|2|5|我们所说将来的世界，上帝没有交给天使管辖。
HEB|2|6|但有人在某处证明说： “人算什么，你竟顾念他； 世人算什么，你竟眷顾他。
HEB|2|7|你使他暂时比天使微小 ， 赐他荣耀尊贵为冠冕， 你派他管理你手所造的，
HEB|2|8|使万物都服在他的脚下。” 既然使万物都服他 ，就没有剩下一样不服他的了。只是如今我们还不见万物都服他；
HEB|2|9|惟独见那成为暂时比天使微小的耶稣，因为受了死的痛苦，得了尊贵荣耀为冠冕，好使他因着上帝的恩，为人人经历了死亡。
HEB|2|10|原来那为万物所属、为万物所本的，为要领许多儿子进入荣耀，使救他们的元帅因受苦难而得以完全，本是合宜的。
HEB|2|11|因那使人成圣的，和那些得以成圣的，都是出于一。为这缘故，他称他们为弟兄也不以为耻，
HEB|2|12|说： “我要将你的名传给我的弟兄， 在会众中我要颂扬你。”
HEB|2|13|他又说： “我要依赖他。” 他又说： “看哪！我与上帝所给我的儿女都在这里。”
HEB|2|14|既然儿女同有血肉之躯，他也照样亲自成了血肉之躯，为能藉着死败坏那掌管死权的，就是魔鬼，
HEB|2|15|并要释放那些一生因怕死而作奴隶的人。
HEB|2|16|诚然，他并没有帮助天使，而是帮助了 亚伯拉罕 的后裔。
HEB|2|17|所以，他凡事应当与他的弟兄相同，为要在上帝的事上成为慈悲忠信的大祭司，为百姓的罪献上赎罪祭。
HEB|2|18|既然他自己被试探而受苦，他能帮助被试探的人。
HEB|3|1|同蒙天召的圣洁弟兄啊，要思想我们所宣认为使者、为大祭司的耶稣；
HEB|3|2|他向指派他的尽忠，如同 摩西 向上帝的全 家尽忠一样。
HEB|3|3|他比 摩西 配得更多的荣耀，好像建造房屋的人比房屋更尊荣；
HEB|3|4|因为房屋都必有人建造，但建造万物的是上帝。
HEB|3|5|摩西 作为仆人，向上帝的全家尽忠，为将来要谈论的事作证；
HEB|3|6|但是基督作为儿子，治理上帝的家。我们若坚持因盼望而有的胆量和夸耀，我们就是他的家了。
HEB|3|7|所以，正如圣灵所说： “今日，你们若听他的话，
HEB|3|8|就不可硬着心，像在背叛之时， 就如在旷野受试探之日。
HEB|3|9|在那里，你们的祖宗试探我， 并且观看我的作为，
HEB|3|10|有四十年之久。 所以，我厌烦那世代， 说：他们的心常常迷糊， 竟不知道我的道路！
HEB|3|11|我在怒中起誓： 他们断不可进入我的安息！”
HEB|3|12|弟兄们，你们要谨慎，免得你们中间有人存着邪恶不信的心，离弃了永生的上帝。
HEB|3|13|总要趁着还有今日，天天彼此相劝，免得你们中间有人被罪迷惑，心肠刚硬了。
HEB|3|14|只要我们将起初确实的信心坚持到底，就在基督里有份了。
HEB|3|15|经上说： “今日，你们若听他的话， 就不可硬着心，像在背叛之时。”
HEB|3|16|听见他而又背叛他的是谁呢？岂不是跟着 摩西 从 埃及 出来的众人吗？
HEB|3|17|上帝向谁发怒四十年之久呢？岂不是那些犯罪而陈尸在旷野的人吗？
HEB|3|18|他向谁起誓，不容他们进入他的安息呢？岂不是向那些不信从的人吗？
HEB|3|19|这样看来，他们不能进入安息是因为不信的缘故了。
HEB|4|1|所以，既然进入他安息的应许依旧存在，我们就该存畏惧的心，免得我们 中间有人似乎没有得到安息。
HEB|4|2|因为的确有福音传给我们像传给他们一样；只是所听见的道对他们无益，因为他们没有以信心与所听见的道配合。
HEB|4|3|但我们已经信的人进入安息，正如上帝所说： “我在怒中起誓： 他们断不可进入我的安息！” 其实造物之工，从创世以来已经完成了。
HEB|4|4|论到第七日，有一处说：“到第七日，上帝就歇了他一切工作。”
HEB|4|5|又有一处说：“他们断不可进入我的安息！”
HEB|4|6|既有这安息保留着让一些人进入，那些先前听见福音的人，因不信从而不得进去，
HEB|4|7|所以上帝多年后藉着 大卫 的书，又定了一天—“今日”，如以上所引的说： “今日，你们若听他的话， 就不可硬着心。”
HEB|4|8|若是 约书亚 已使他们享了安息，后来上帝就不会再提别的日子了。
HEB|4|9|这样看来，另有一安息日的安息为上帝的子民保留着。
HEB|4|10|因为那些进入安息的，也是歇了自己的工作，正如上帝歇了他的工作一样。
HEB|4|11|所以，我们务必竭力进入那安息，免得有人学了不顺从而跌倒了。
HEB|4|12|上帝的道是活泼的，是有功效的，比一切两刃的剑更锋利，甚至魂与灵、骨节与骨髓，都能刺入、剖开，连心中的思念和主意都能辨明。
HEB|4|13|被造的，没有一样在他面前不是显露的；万物在他眼前都是赤露敞开的，我们必须向他交账。
HEB|4|14|既然我们有一位伟大、进入高天的大祭司，就是耶稣—上帝的儿子，我们应当持定所宣认的道。
HEB|4|15|因为我们的大祭司并非不能体恤我们的软弱；他也在各方面受过试探，与我们一样，只是他没有犯罪。
HEB|4|16|所以，我们只管坦然无惧地来到施恩的宝座前，为要得怜悯，蒙恩惠，作及时的帮助。
HEB|5|1|凡从人间挑选的大祭司都是奉派替人办理属上帝的事，要为罪献上礼物和祭物 。
HEB|5|2|他能体谅无知和迷失的人，因为他自己也是被软弱所困，
HEB|5|3|因此他理当为百姓和自己的罪献祭。
HEB|5|4|没有人可擅自取得大祭司的尊荣，惟有蒙上帝所选召的才可以，像 亚伦 一样。
HEB|5|5|同样，基督也没有自取作大祭司的荣耀，而是在乎向他说话的那一位，他说： “你是我的儿子， 我今日生了你。”
HEB|5|6|就如又有一处说： “你是照着 麦基洗德 的体系 永远为祭司。”
HEB|5|7|基督在他肉身的日子，曾大声哀哭，流泪祷告，恳求那能救他免死的上帝，就因他的虔诚蒙了应允。
HEB|5|8|他虽然为儿子，还是因所受的苦难学了顺从。
HEB|5|9|既然他得以完全，就为凡顺从他的人成了永远得救的根源，
HEB|5|10|并蒙上帝照着 麦基洗德 的体系宣称他为大祭司。
HEB|5|11|论到这事，我们有好些话要说，可是很难解释，因为你们听不进去。
HEB|5|12|按时间说，你们早该作教师了，谁知还需要有人再将上帝圣言基础的要道教导你们；你们成了那需要吃奶、不能吃干粮的人。
HEB|5|13|凡只能吃奶的，就不熟练仁义的道理，因为他是婴孩。
HEB|5|14|惟独长大成人的才能吃干粮，他们的心窍因练习而灵活，能分辨善恶了。
HEB|6|1|所以，我们应当离开基督道理的基础，竭力进到成熟的地步；不必再立根基，就如懊悔致死的行为、信靠上帝、
HEB|6|2|各样洗礼、按手礼、死人复活，以及永远的审判等的教导。
HEB|6|3|上帝若准许，我们就这样做。
HEB|6|4|论到那些已经蒙了光照、尝过天恩的滋味、又于圣灵有份、并尝过上帝的话的美味，和来世权能的人，若再离弃真道，就不可能使他们重新懊悔了；因为他们亲自把上帝的儿子重钉十字架，公然羞辱他。
HEB|6|5|
HEB|6|6|
HEB|6|7|就如一块田地吸收过屡次下的雨水，生长蔬菜，合乎耕种的人用，就从上帝得福。
HEB|6|8|这块田地若长荆棘和蒺藜，必被废弃，近于诅咒，结局就是焚烧。
HEB|6|9|亲爱的，虽然这样说，我们仍深信你们有更好的情况，更接近救恩。
HEB|6|10|因为上帝并非不公义，竟忘记你们的工作和你们为他的名所显的爱心，就是你们过去和现在伺候圣徒的爱心。
HEB|6|11|我们盼望你们各人都显出同样的热忱，一直到底，好达成所确信的指望。
HEB|6|12|这样你们才不会懒惰，却成为效法那些藉着信和忍耐承受应许的人。
HEB|6|13|当初上帝应许 亚伯拉罕 的时候，因为没有比自己更大的可以指着起誓，就指着自己起誓，
HEB|6|14|说：“我必多多赐福给你；我必使你大大增多。”
HEB|6|15|这样， 亚伯拉罕 因恒心等待而得了所应许的。
HEB|6|16|人都是指着比自己大的起誓，并且以起誓作保证，了结各样的争论。
HEB|6|17|照样，上帝愿意为那承受应许的人更有力地显明他的旨意不可更改，他以起誓作保证。
HEB|6|18|藉这两件不可更改的事—在这些事上，上帝绝不会说谎—我们这些逃往避难所的人能得到强有力的鼓励，去抓住那摆在我们前头的指望。
HEB|6|19|我们有这指望，如同灵魂的锚，又坚固又牢靠，进入幔子后面的至圣所。
HEB|6|20|为我们作先锋的耶稣，既照着 麦基洗德 的体系成了永远的大祭司，已经进入了。
HEB|7|1|这 麦基洗德 就是 撒冷 王，是至高上帝的祭司。他在 亚伯拉罕 打败诸王回来的时候迎接他，并给他祝福。
HEB|7|2|亚伯拉罕 也将自己所得来的一切，取十分之一给他。他头一个名字翻译出来是“公义的王”，他又名“ 撒冷 王”，是和平王的意思。
HEB|7|3|他无父、无母、无族谱、无生之始、无命之终，是与上帝的儿子相似，他永远作祭司。
HEB|7|4|你们想一想，这个人多么伟大啊！连先祖 亚伯拉罕 都拿战利品的十分之一给他。
HEB|7|5|那得祭司职分的 利未 子孙，奉命照例向百姓取十分之一，这百姓是自己的弟兄，虽是从 亚伯拉罕 亲身生的，还是照例取十分之一。
HEB|7|6|惟独 麦基洗德 那不与他们同族谱的，从 亚伯拉罕 收取了十分之一，并且给蒙应许的 亚伯拉罕 祝福。
HEB|7|7|向来位分大的给位分小的祝福，这是无可争议的。
HEB|7|8|在这事上，一方面，收取十分之一的都是必死的人；另一方面，收取十分之一的却是那位被证实是活着的。
HEB|7|9|我们可以说，那接受十分之一的 利未 也是藉着 亚伯拉罕 纳了十分之一，
HEB|7|10|因为 麦基洗德 迎接 亚伯拉罕 的时候， 利未 还在他先祖的身体里面。
HEB|7|11|那么，如果百姓藉着 利未 人的祭司职任能达到完全—因为百姓是在这职分下领受律法的—为什么还需要按照 麦基洗德 的体系另外兴起一位祭司，而不按照 亚伦 的体系呢？
HEB|7|12|既然祭司的职分已更改，律法也需要更改。
HEB|7|13|因为这些话所指的人本属别的支派，那支派里从来没有一人在祭坛前事奉的。
HEB|7|14|很明显地，我们的主是从 犹大 出来的；但关于这支派， 摩西 并没有提到祭司。
HEB|7|15|倘若有另一位像 麦基洗德 的祭司兴起来，我的话就更显而易见了。
HEB|7|16|他成为祭司，并不是照属肉身的条例，而是照无穷 生命的大能。
HEB|7|17|因为有给他作见证的说： “你是照着 麦基洗德 的体系 永远为祭司。”
HEB|7|18|一方面，先前的诫命因软弱无能而废掉了，
HEB|7|19|（律法本来就不能成就什么）；另一方面，一个更好的指望被引进来，靠这指望，我们就可以亲近上帝。
HEB|7|20|再者，耶稣成为祭司，并不是没有上帝的誓言；其他的祭司被指派时并没有这种誓言，
HEB|7|21|只有耶稣是起誓立的，因为那位立他的对他说： “主起了誓， 绝不改变。 你是永远为祭司。”
HEB|7|22|既是起誓立的，耶稣也作了更美之约的中保。
HEB|7|23|一方面，那些成为祭司的数目本来多，是因为受死亡限制不能长久留住。
HEB|7|24|另一方面，这位既是永远留住的，他具有不可更换的祭司职任。
HEB|7|25|所以，凡靠着他进到上帝面前的人，他都能拯救到底，因为他长远活着为他们祈求。
HEB|7|26|这样一位圣洁、无邪恶、无玷污、远离罪人、高过诸天的大祭司，对我们是最合适的；
HEB|7|27|他不像那些大祭司，每日必须先为自己的罪，后为百姓的罪献祭，因为他只一次将自己献上就把这事成全了。
HEB|7|28|律法所立的大祭司本是有弱点的人，但在律法以后，上帝以起誓的话立了儿子为大祭司，成为完全，直到永远。
HEB|8|1|我们所讲的事，其中第一要紧的就是：我们有这样一位大祭司，他已经坐在天上至大者宝座的右边，
HEB|8|2|在圣所，就是在真帐幕里作仆役；这帐幕是主所支搭的，不是人所支搭的。
HEB|8|3|凡大祭司都是为献礼物和祭物设立的，所以这位大祭司也必须有所献上。
HEB|8|4|他若在地上，就不用作祭司，因为已经有照律法献礼物的祭司了。
HEB|8|5|他们所供奉的本是天上之事的样式和影像，正如 摩西 将要造帐幕的时候，上帝警戒他，说：“要谨慎，一切都要照着在山上指示你的样式去做。”
HEB|8|6|如今耶稣已经得了更优越的事奉，正如他作更美之约的中保；这约原是凭更美之应许立的。
HEB|8|7|第一个约若没有瑕疵，就无须寻求第二个约了。
HEB|8|8|所以上帝指责他们说： “主说，看哪，日子将到， 我要与 以色列 家 和 犹大 家另立新的约；
HEB|8|9|不像我拉着他们祖宗的手 领他们出 埃及 地的时候， 与他们所立的约； 因为他们不恒心守我的约， 所以我也不理他们；这是主说的。
HEB|8|10|主又说： 那些日子以后， 我与 以色列 家所立的约是这样： 我要将我的律法放在他们的心思里， 写在他们的心上； 我要作他们的上帝， 他们要作我的子民。
HEB|8|11|他们各人不用教导自己的乡亲和自己的弟兄，说：你要认识主； 因为从最小的到最大的， 他们都要认识我。
HEB|8|12|我要宽恕他们的不义， 绝不再记得他们的罪恶。”
HEB|8|13|既然上帝提到“新的约”，那么第一个约就成为旧的了；而那渐旧渐衰的必然很快消逝了。
HEB|9|1|原来连第一个约都有敬拜的礼仪和属世界的圣幕。
HEB|9|2|因为那预备好了的帐幕，第一层叫圣所，里面有灯台、供桌和供饼。
HEB|9|3|第二层幔子后又有一层帐幕，叫至圣所，
HEB|9|4|有金香坛和四周包金的约柜，柜里有盛吗哪的金罐、 亚伦 那根发过芽的杖和两块约版；
HEB|9|5|柜上面有荣耀的基路伯罩着施恩座。有关这一切我现在不能一一细说。
HEB|9|6|这些物件既如此预备齐了，众祭司就不断地进第一层帐幕行拜上帝的礼。
HEB|9|7|至于第二层帐幕，惟有大祭司一年一次独自进去，没有一次不带着血，为自己献上，也为百姓无意所犯的过错献上。
HEB|9|8|圣灵藉此指明，第一层帐幕仍存在的时候，进入至圣所的路还没有显示。
HEB|9|9|那第一层帐幕是现今时代的一个预表，表示所献的礼物和祭物都不能使敬拜的人在良心上得以完全。
HEB|9|10|这些事只不过是有关饮食和各种洁净的规矩，是属肉体的条例，它的功效是直到新次序的时期来到为止。
HEB|9|11|但现在基督已经来到，作了已实现的美事的大祭司，经过那更大更全备的帐幕，不是人手所造，也不是属于这世界的；
HEB|9|12|他不用山羊和牛犊的血，而是用自己的血，只一次进入至圣所就获得了永远的赎罪。
HEB|9|13|若山羊和公牛的血，以及母牛犊的灰，洒在不洁的人身上，尚且使人成圣，身体洁净，
HEB|9|14|何况基督的血，他藉着永远的灵把自己无瑕疵地献给上帝，更能洗净我们 的良心，除去致死的行为，好事奉那位永生的上帝。
HEB|9|15|为此，基督作了新约的中保；因为他的死，赎了人在第一个约之时所犯的罪过，使蒙召的人能得着所应许永远的产业。
HEB|9|16|凡有遗嘱，必须证实立遗嘱的人已经死了。
HEB|9|17|因为人死了，遗嘱才有效力；立遗嘱的人尚在，遗嘱就不能生效。
HEB|9|18|所以，第一个约也是用血立的。
HEB|9|19|因为 摩西 当日照着律法将各样诫命传给众百姓，就拿朱红色绒和牛膝草，把牛犊、山羊 的血和水洒在书上，又洒在众百姓身上，
HEB|9|20|说：“这血就是上帝与你们立约的凭据。”
HEB|9|21|他又照样把血洒在帐幕和敬拜用的各样器皿上。
HEB|9|22|按着律法，几乎每样东西都是用血洁净的；没有流血，就没有赦罪。
HEB|9|23|这样，照着天上样式做的物件必须用这些礼仪去洁净，但那天上的一切，自然当用更美的祭物去洁净。
HEB|9|24|因为基督并没有进了人手所造的圣所—这不过是真圣所的影像—而是进到天上，如今为我们出现在上帝面前。
HEB|9|25|他也无须多次将自己献上，像大祭司每年带着牛羊的血进入至圣所。
HEB|9|26|如果这样，他从创世以来就必须多次受苦了。但如今，他在今世的末期显现，仅一次把自己献为祭，好除掉罪。
HEB|9|27|按着命定，人人都有一死，死后且有审判。
HEB|9|28|同样，基督既然一次献上，担当了许多人的罪，将来要第二次显现，与罪无关，而是为了拯救热切等候他的人。
HEB|10|1|既然律法只不过是未来美好事物的影子，不是本体的真像，就不能藉着每年常献一样的祭物，使那些进前来的人完全。
HEB|10|2|若不然，献祭的事岂不早已停止了吗？因为敬拜的人仅只一次洁净，良心就不再觉得有罪了。
HEB|10|3|但是这些祭物使人每年都想起罪来，
HEB|10|4|因为公牛和山羊的血不能除罪。
HEB|10|5|所以，基督到世上来的时候，就说： “祭物和礼物不是你所要的， 但你曾给我预备了身体。
HEB|10|6|燔祭和赎罪祭 是你不喜欢的。
HEB|10|7|那时我说： 看哪！我来了，我的事在经卷上已经记载了； 上帝啊！我来为要照你的旨意行。”
HEB|10|8|以上说：“祭物和礼物，以及燔祭和赎罪祭，不是你所要的，也不是你喜欢的。”这都是按着律法献的。
HEB|10|9|他接着说：“看哪！我来了，为要照你的旨意行。”可见他除去在先的，为要立定在后的。
HEB|10|10|我们凭着这旨意，藉着耶稣基督，仅只一次献上他的身体就得以成圣。
HEB|10|11|所有的祭司天天站着事奉上帝，屡次献上一样的祭物，这祭物永不能除罪。
HEB|10|12|但基督献了一次永远有效的赎罪祭，就坐在上帝的右边，
HEB|10|13|从此等候他的仇敌成为他的脚凳。
HEB|10|14|因为他仅只一次献祭，就使那些得以成圣的人永远完全。
HEB|10|15|圣灵也对我们作证，因为他说过：
HEB|10|16|“主说：那些日子以后， 我与他们所立的约是这样的： 我要将我的律法放在他们的心上， 又要写在他们的心思里。”
HEB|10|17|并说： “他们的罪恶和他们的过犯， 我绝不再记得。”
HEB|10|18|这些罪过既已蒙赦免，就不用再为罪献祭了。
HEB|10|19|所以，弟兄们，既然我们靠着耶稣的血得以坦然进入至圣所，
HEB|10|20|是藉着他给我们开了一条又新又活的路，从幔子经过，这幔子就是他的身体。
HEB|10|21|既然我们有一位伟大祭司治理上帝的家，
HEB|10|22|那么，我们该用诚心和充足的信心，同已蒙洁净、无亏的良心，和清水洗净了的身体来亲近上帝。
HEB|10|23|我们要坚守所宣认的指望，毫不动摇，因为应许我们的那位是信实的。
HEB|10|24|我们要彼此相顾，激发爱心，勉励行善；
HEB|10|25|不可停止聚会，好像那些停止惯了的人，倒要彼此劝勉，既然知道那日子临近，就更当如此。
HEB|10|26|如果我们领受真理的知识以后仍故意犯罪，就不再有赎罪的祭物，
HEB|10|27|惟有战战兢兢等候审判和那将吞灭众敌人的烈火了。
HEB|10|28|任何人干犯 摩西 的律法，凭两个或三个证人，尚且必须处死，不得宽赦，
HEB|10|29|更何况践踏上帝儿子的人，他们将那使他成圣之约的血当作不洁净，又亵慢施恩的圣灵的人，你们想，他不该受更严厉的惩罚吗？
HEB|10|30|因为我们知道谁说： “伸冤在我， 我必报应。” 又说： “主要审判他的百姓。”
HEB|10|31|落在永生上帝的手里真是可怕呀！
HEB|10|32|你们要追念往日；你们蒙了光照以后，忍受了许多痛苦的挣扎：
HEB|10|33|一面在众人面前公然被毁谤，遭患难；一面陪伴那些受这样苦难的人。
HEB|10|34|你们同情那些遭监禁的人，也欣然忍受你们的家业被人抢去，因为你们知道自己有更美好更长存的家业。
HEB|10|35|所以，不可丢弃你们无惧的心，存这样的心必得大赏赐。
HEB|10|36|你们必须忍耐，使你们行完了上帝的旨意，可以获得所应许的。
HEB|10|37|因为 “还有一点点时候， 那要来的就来，必不迟延。
HEB|10|38|只是我的义人必因信得生； 他若退缩，我心就不喜欢他。”
HEB|10|39|我们却不是退缩以致沉沦的那等人，而是有信心以致得生命的人。
HEB|11|1|信就是对所盼望之事有把握，对未见之事有确据。
HEB|11|2|古人因着这信获得了赞许。
HEB|11|3|因着信，我们知道这宇宙是藉上帝的话造成的。这样，看得见的是从看不见的造出来的。
HEB|11|4|因着信， 亚伯 献祭给上帝比 该隐 所献的更美，因此获得了赞许为义人，上帝亲自悦纳了他的礼物。他虽然死了，却因这信仍旧在说话。
HEB|11|5|因着信， 以诺 被接去，得以不见死，人也找不着他，因为上帝已经把他接去了；只是他被接去以前，已讨得上帝的喜悦而蒙赞许。
HEB|11|6|没有信，就不能讨上帝的喜悦，因为到上帝面前来的人必须信有上帝，并且信他会赏赐寻求他的人。
HEB|11|7|因着信， 挪亚 既蒙上帝指示他未见的事，动了敬畏的心，造了方舟，使他全家得救。藉此他定了那世代的罪，自己也承受了那从信而来的义。
HEB|11|8|因着信， 亚伯拉罕 蒙召的时候就遵命出去，往将来要承受为基业的地方去；他出去的时候还不知往哪里去。
HEB|11|9|因着信，他就在所应许之地作客，好像在异乡，居住在帐棚里，与蒙同一个应许的 以撒 和 雅各 一样。
HEB|11|10|因为他等候着那座有根基的城，就是上帝所设计和建造的。
HEB|11|11|因着信， 撒拉 自己已过了生育的年龄还能怀孕，因为她认为应许她的那位是可信的 ；
HEB|11|12|所以，从一个仿佛已死的人竟生出子孙，如同天上的星那样众多，海边的沙那样无数。
HEB|11|13|这些人都是存着信心死的，并没有得着所应许的，却从远处观望，且欢喜迎接。他们承认自己在地上是客旅，是寄居的。
HEB|11|14|说这样话的人是表明自己要寻找一个家乡。
HEB|11|15|他们若想念所离开的家乡，还有回去的机会。
HEB|11|16|其实他们所羡慕的是一个更美的，就是在天上的家乡。所以，上帝并不因他们称他为上帝 而觉得羞耻，因为他已经为他们预备了一座城。
HEB|11|17|因着信， 亚伯拉罕 被考验的时候把 以撒 献上，这就是那领受了应许的人甘心把自己独生的儿子献上。
HEB|11|18|论到这儿子，上帝曾说：“从 以撒 生的才要称为你的后裔。”
HEB|11|19|他认为上帝甚至能使人从死人中复活，意味着他得回了他的儿子。
HEB|11|20|因着信， 以撒 指着将来的事给 雅各 、 以扫 祝福。
HEB|11|21|因着信， 雅各 临死的时候给 约瑟 的两个儿子个别祝福，扶着拐杖敬拜上帝。
HEB|11|22|因着信， 约瑟 临终的时候提到 以色列 人将来要出 埃及 ，并为自己的骸骨留下遗言。
HEB|11|23|因着信， 摩西 生下来，他的父母见他是个俊美的孩子，把他藏了三个月，并不怕王的命令。
HEB|11|24|因着信， 摩西 长大了不肯称为法老女儿之子。
HEB|11|25|他宁可和上帝的百姓一同受苦，也不愿在罪中享受片刻的欢乐。
HEB|11|26|他把为弥赛亚受凌辱看得比 埃及 的财物更宝贵，因为他想望所要得的赏赐。
HEB|11|27|因着信，他离开 埃及 ，不怕王的愤怒，因为他恒心忍耐，如同看见那不能看见的上帝。
HEB|11|28|因着信，他设立逾越节，在门上洒血，免得那毁灭者加害 以色列 人的长子。
HEB|11|29|因着信，他们过 红海 如行干地； 埃及 人试着要过去就被淹没了。
HEB|11|30|因着信， 以色列 人围绕 耶利哥城 七日，城墙就倒塌了。
HEB|11|31|因着信，妓女 喇合 曾友善地接待探子，就没有跟那些不顺从的人一同灭亡。
HEB|11|32|我还要说什么呢？若要一一细说 基甸 、 巴拉 、 参孙 、 耶弗他 、 大卫 、 撒母耳 和众先知的事，时间就不够了。
HEB|11|33|他们藉着信，制伏了敌国，行了公义，得了应许，堵住了狮子的口，
HEB|11|34|灭了烈火的威力，在锋利的刀剑下逃生，从软弱变为刚强，争战中显出勇猛，打退外邦的全军。
HEB|11|35|有些妇人得回从死人中复活的亲人。又有人忍受严刑，拒绝被释放，为要得着更美好的复活。
HEB|11|36|又有人忍受戏弄、鞭打、捆锁、监禁、各等的磨炼；
HEB|11|37|他们被石头打死，被锯锯死， 被刀杀，披着绵羊山羊的皮各处奔跑，受贫穷、患难、虐待。
HEB|11|38|这世界配不上他们，他们在旷野、山岭、山洞、地穴，飘流无定。
HEB|11|39|这些人都是因信获得了赞许，却仍未得着所应许的，
HEB|11|40|因为上帝给我们预备了更美好的事，若没有我们，他们就不能达到完全。
HEB|12|1|所以，既然我们有这许多见证人如同云彩围绕着我们，就该卸下各样重担和紧紧缠累的罪，以坚忍的心奔那摆在我们前头的路程，
HEB|12|2|仰望我们信心的创始成终者耶稣，他因那摆在前面的喜乐，轻看羞辱，忍受了十字架的苦难，如今已坐在上帝宝座的右边。
HEB|12|3|你们要仔细想想这位忍受了罪人如此顶撞的耶稣，你们就不致心灰意懒了。
HEB|12|4|你们与罪恶争斗，还没有抵抗到流血的地步。
HEB|12|5|你们又忘了上帝劝你们如同劝儿女的那些话，说： “我儿啊，不可轻看主的管教， 被他责备的时候不可灰心；
HEB|12|6|因为主所爱的，他必管教， 又鞭打他所接纳的每一个孩子。”
HEB|12|7|为了受管教，你们要忍受。上帝待你们如同待儿女。哪有儿女不被父亲管教的呢？
HEB|12|8|管教原是众儿女共同所领受的；你们若不受管教，就是私生子，不是儿女了。
HEB|12|9|再者，我们曾有肉身之父管教我们，我们尚且敬重他，何况灵性之父，我们岂不更当顺服他而得生命吗？
HEB|12|10|肉身之父都是短时间随己意管教我们，惟有灵性之父管教我们是要我们得益处，使我们在他的圣洁上有份。
HEB|12|11|凡管教的事，当时不觉得快乐，反觉得痛苦；后来却为那经过锻鍊的人结出平安的果子，就是义的果子。
HEB|12|12|所以，你们要把下垂的手举起来，发酸的腿挺直；
HEB|12|13|要为自己的脚把道路修直了，使瘸了的腿不再脱臼，反而得到痊愈。
HEB|12|14|你们要追求与众人和睦，并要追求圣洁；人非圣洁不能见主。
HEB|12|15|要谨慎，免得有人失去了上帝的恩典；免得有毒根生出来扰乱你们，因而使许多人沾染污秽，
HEB|12|16|免得有人淫乱，或不敬虔如 以扫 ，他因一点点食物把自己长子的名分卖了。
HEB|12|17|后来你们知道，他想要承受父亲的祝福，竟被拒绝，虽然流着泪苦求，却得不着门路使他父亲回心转意。
HEB|12|18|你们不是来到那可触摸的山，那里有火焰、密云、黑暗、暴风、
HEB|12|19|角声，和说话的声音；当时那些听见这声音的，都求不要再向他们说话，
HEB|12|20|因为他们担当不起所命令他们的话，说：“靠近这山的，即使是走兽，也要用石头打死。”
HEB|12|21|所见的景象极其可怕，以致 摩西 说：“我恐惧战兢。”
HEB|12|22|但是你们是来到 锡安山 ，永生上帝的城，就是天上的 耶路撒冷 ，那里有千千万万的天使，
HEB|12|23|有名字记录在天上众长子的盛会，有审判众人的上帝和成为完全的义人的灵魂，
HEB|12|24|并新约的中保耶稣，以及所洒的血；这血所说的信息比 亚伯 的血所说的更美。
HEB|12|25|你们总要谨慎，不可拒绝那向你们说话的，因为那些拒绝了在地上警戒他们的，尚且不能逃罪，何况我们违背那从天上警戒我们的呢？
HEB|12|26|当时他的声音震动了地，但如今他应许说：“再一次我不单要震动地，还要震动天。”
HEB|12|27|这“再一次”的话是指明被震动的要像受造之物一样被挪去，使那不被震动的能常存。
HEB|12|28|所以，既然我们得了不能被震动的国度，就要感恩，照着上帝所喜悦的，用虔诚、敬畏的心事奉上帝，
HEB|12|29|因为我们的上帝是吞灭的火。
HEB|13|1|你们务要常存弟兄相爱的心。
HEB|13|2|不可忘记用爱心接待旅客，因为曾经有人这样做，在无意中接待了天使。
HEB|13|3|要记念受监禁的人，好像与他们同受监禁；要记念受虐待的人，好像你们也亲身受虐待一样。
HEB|13|4|婚姻，人人都当尊重，共眠的床也不可污秽，因为淫乱和通奸的人，上帝必审判。
HEB|13|5|不可贪爱钱财，要以自己所有的为满足，因为上帝曾说：“我绝不撇下你，也绝不丢弃你。”
HEB|13|6|所以，我们可以勇敢地说： “主是我的帮助， 我必不惧怕。 人能把我怎么样呢？”
HEB|13|7|从前引导你们、传上帝的道给你们的人，你们要记念他们，效法他们的信心，回顾他们为人的结局。
HEB|13|8|耶稣基督昨日、今日，一直到永远，是一样的。
HEB|13|9|你们不要被种种怪异的教训勾引了去，因为人的心靠恩典得坚固才是好的，并不是靠饮食。那在饮食上用心的，从来没有得到益处。
HEB|13|10|我们有一祭坛，上面的祭物是那些在会幕中供职的人无权可吃的。
HEB|13|11|因为牲畜的血被大祭司带入至圣所作赎罪祭，牲畜的体却在营外烧掉。
HEB|13|12|所以，耶稣也在城门外受苦，为要用自己的血使百姓成圣。
HEB|13|13|这样，我们也当走出营外，到他那里去，忍受他所受的凌辱。
HEB|13|14|在这里，我们本没有永存的城，而是在寻求那将要来的城。
HEB|13|15|我们应当藉着耶稣，常常以颂赞为祭献给上帝，这是那宣认他名的人嘴唇所结的果子。
HEB|13|16|只是不可忘记行善和分享，因为这样的祭物是上帝所喜悦的。
HEB|13|17|你们要服从那些引导你们的，并且要顺服，因为他们为你们的灵魂时刻警醒，像在上帝面前交账的人，让他们在交账的时候有喜乐，而不是叹息，叹息就对你们无益了。
HEB|13|18|请你们为我们祷告；因为我们自觉良心无亏，愿意凡事按正道而行。
HEB|13|19|我更求你们为我祷告，使我快些回到你们那里去。
HEB|13|20|但愿赐平安 的上帝，就是那凭永约之血，把群羊的大牧人—我们主耶稣从死人中领出来的上帝，
HEB|13|21|在各样善事上装备你们，使你们遵行他的旨意；又藉着耶稣基督在我们 里面行他所喜悦的事。愿荣耀归给他，直到永永远远 。阿们！
HEB|13|22|弟兄们，我简略地写信给你们，希望你们听我劝勉的话。
HEB|13|23|你们该知道，我们的弟兄 提摩太 已经重获自由了；他若很快就来，我必同他去见你们。
HEB|13|24|请你们向带领你们的诸位和众圣徒问安。从 意大利 来的人也向你们问安。
HEB|13|25|愿恩惠与你们众人同在。
