AMOS|1|1|Verba Amos, qui fuit in pastori bus de Thecua; quae vidit super Israel in diebus Oziae regis Iudae et in diebus Ieroboam filii Ioas regis Israel, duobus annis ante terraemotum.
AMOS|1|2|Et dixit: Dominus de Sion rugitet de Ierusalem dat vocem suam;et lugent pascua pastorum,et exsiccatur vertex Carmeli ".
AMOS|1|3|Haec dicit Dominus: Super tribus sceleribus Damasciet super quattuor verbum non revocabo:eo quod trituraverint in plaustris ferreis Galaad,
AMOS|1|4|mittam ignem in domum Hazael,et devorabit aedes Benadad;
AMOS|1|5|conteram vectem Damasciet disperdam habitatorem de Biceatavenet tenentem sceptrum de Betheden;et transferetur populus Syriae Cir ",dicit Dominus.
AMOS|1|6|Haec dicit Dominus: Super tribus sceleribus Gazaeet super quattuor verbum non revocabo:eo quod transtulerint captivitatem perfectam,ut traderent eam in Edom,
AMOS|1|7|mittam ignem in murum Gazae,et devorabit aedes eius;
AMOS|1|8|disperdam habitatorem de Azotoet tenentem sceptrum de Ascalone;convertam manum meam super Accaron,et peribunt reliqui Philisthinorum ",dicit Dominus Deus.
AMOS|1|9|Haec dicit Dominus: Super tribus sceleribus Tyriet super quattuor verbum non revocabo:eo quod tradiderint captivitatem perfectam in Edomet non sint recordati foederis fratrum,
AMOS|1|10|mittam ignem in murum Tyri,et devorabit aedes eius ".
AMOS|1|11|Haec dicit Dominus: Super tribus sceleribus Edomet super quattuor verbum non revocabo:eo quod persecutus sit in gladio fratrem suumet violaverit misericordiam eiuset tenuerit ultra furorem suumet indignationem suam servaverit usque in finem,
AMOS|1|12|mittam ignem in Theman,et devorabit aedes Bosrae ".
AMOS|1|13|Haec dicit Dominus: Super tribus sceleribus filiorum Ammonet super quattuor verbum non revocabo:eo quod dissecuerint praegnantes Galaadad dilatandum terminum suum,
AMOS|1|14|succendam ignem in muro Rabba,et devorabit aedes eius in ululatu in die belliet in turbine in die procellae;
AMOS|1|15|et ibit rex eorum in captivitatem,ipse et principes eius simul ",dicit Dominus.
AMOS|2|1|Haec dicit Dominus: Super tribus sceleribus Moabet super quattuor verbum non revocabo:eo quod incenderit ossa regis Edomusque ad cinerem,
AMOS|2|2|mittam ignem in Moab,et devorabit aedes Carioth,et morietur in tumultu Moab,in clamore et voce tubae;
AMOS|2|3|disperdam iudicem de medio eiuset omnes principes eius interficiam cum eo ",dicit Dominus.
AMOS|2|4|Haec dicit Dominus: Super tribus sceleribus Iudaeet super quattuor verbum non revocabo:eo quod abiecerint legem Dominiet mandata eius non custodierintC deceperunt enim eos idola sua,post quae abierant patres eorum C
AMOS|2|5|mittam ignem in Iudam,et devorabit aedes Ierusalem ".
AMOS|2|6|Haec dicit Dominus: Super tribus sceleribus Israelet super quattuor verbum non revocabo:eo quod vendiderint pro argento iustumet pauperem pro calceamentis;
AMOS|2|7|qui contriverint super pulverem terrae capita pauperumet viam humilium declinaverint,et filius ac pater eius iverint ad puellam,ut violarent nomen sanctum meum;
AMOS|2|8|et super vestimentis pignoratis accubuerintiuxta omne altareet vinum damnatorum biberintin domo Dei sui.
AMOS|2|9|Ego autem exterminaveramAmorraeum a facie eorum,cuius altitudo sicut altitudo cedrorum,et fortitudo quasi quercuum;exterminaveram fructum eius desuperet radices eius subter.
AMOS|2|10|Ego ascendere vos fecide terra Aegyptiet duxi vos in desertoquadraginta annis,ut possideretis terram Amorraei;
AMOS|2|11|et suscitavi de filiis vestris prophetas et de iuvenibus vestris nazaraeos.Numquid non ita est, filii Israel?,dicit Dominus.
AMOS|2|12|Et propinastis nazaraeis vinumet prophetis mandastis dicentes:Ne prophetetis".
AMOS|2|13|Ecce ego comprimam vos ad solum,sicut comprimit plaustrumonustum feno;
AMOS|2|14|deerit fuga a veloce,et fortis non firmabit virtutem suam,et robustus non salvabit animam suam;
AMOS|2|15|tenens arcum non stabit,et velox pedibus suis non salvabitur;ascensor equi non salvabit animam suam,
AMOS|2|16|et fortissimus corde inter robustosnudus fugiet in illa die ",dicit Dominus.
AMOS|3|1|Audite verbum hoc, quod locutus est Dominus super vos, filii Israel, super omnem cognationem, quam eduxi de terra Aegypti, dicens:
AMOS|3|2|" Tantummodo vos cognoviex omnibus cognationibus terrae;idcirco visitabo super vosomnes iniquitates vestras.
AMOS|3|3|Numquid ambulabunt duo pariter, nisi convenerint?
AMOS|3|4|Numquid rugiet leo in saltu,nisi habuerit praedam?Numquid dabit catulus leonis vocem de cubili suo,nisi aliquid apprehenderit?
AMOS|3|5|Numquid cadet avis super terramabsque laqueo?Numquid laxatur laqueus de terra, antequam quid ceperit?
AMOS|3|6|Si clanget tuba in civitate,populus non expavescet?Si erit malum in civitate,nonne Dominus fecit?
AMOS|3|7|Nihil enim faciet Dominus Deus,nisi revelaverit secretum suumad servos suos prophetas.
AMOS|3|8|Leo rugit,quis non timebit?Dominus Deus locutus est,quis non prophetabit?
AMOS|3|9|Auditum facite in aedibus Assyriaeet in aedibus terrae Aegyptiet dicite: "Congregamini super montes Samariae";et videte insanias multas in medio eiuset oppressos in sinu eius.
AMOS|3|10|Et nescierunt facere rectum,dicit Dominus,thesaurizantes violentiam et rapinasin aedibus suis ".
AMOS|3|11|Propterea haec dicit Dominus Deus: Inimicus circumdabit terram,et detrahetur ex te fortitudo tua,et diripientur aedes tuae ".
AMOS|3|12|Haec dicit Dominus: Quomodo si eruat pastor de ore leonisduo crura aut extremum auriculae, sic eruentur filii Israel,qui habitant in Samaria,in margine lectuliet in Damasci grabato.
AMOS|3|13|Audite et contestamini in domo Iacob,dicit Dominus, Deus exercituum:
AMOS|3|14|In die cum visitavero praevaricationes Israel,super eum visitabo et super altaria Bethel,et amputabuntur cornua altariset cadent in terram;
AMOS|3|15|et percutiam domum hiemalemcum domo aestiva,et peribunt domus eburneae,et dissipabuntur aedes magnae ",dicit Dominus.
AMOS|4|1|Audite verbum hoc,vaccae Basan,quae estis in monte Samariae,quae opprimitis egenoset vexatis pauperes,quae dicitis dominis vestris: Affer, ut bibamus ".
AMOS|4|2|Iuravit Dominus Deusin sanctitate sua: Ecce dies venient super vos,et levabunt vos in contiset posteros vestros in hamis piscatoriis;
AMOS|4|3|et per aperturas exibitis altera contra alteramet proiciemini in Armon ",dicit Dominus.
AMOS|4|4|" Venite in Bethel et impie agite,ad Galgalam et multiplicate praevaricationem;et offerte mane victimas vestras,tribus diebus decimas vestras,
AMOS|4|5|et sacrificate de fermentato laudemet vocate voluntarias oblationes et annuntiate;sic enim diligitis, filii Israel ",dicit Dominus Deus.
AMOS|4|6|" Unde et ego dedi vobisvacuitatem dentium in cunctis urbibus vestriset indigentiam panis in omnibus locis vestris;et non estis reversi ad me ",dicit Dominus.
AMOS|4|7|" Ego quoque prohibui a vobis imbrem,cum adhuc tres menses superessent usque ad messem;et plui super unam civitatemet super alteram civitatem non plui: pars una compluta est,et pars, super quam non plui, aruit.
AMOS|4|8|Tunc fugiebant duae, tres civitatesad unam civitatem, ut biberent aquam,et non satiabantur;sed non redistis ad me ",dicit Dominus.
AMOS|4|9|" Percussi vos in vento urente et in aurugine;multitudinem hortorum vestrorum et vinearum vestrarum,ficeta vestra et oliveta vestracomedit eruca;sed non redistis ad me ",dicit Dominus.
AMOS|4|10|" Misi in vos pestemsicut pestem Aegypti,percussi in gladio iuvenes vestros,captis equis vestris;et ascendere feci putredinemcastrorum vestrorum in nares vestras;sed non redistis ad me ",dicit Dominus.
AMOS|4|11|" Subverti vos,sicut subvertit Deus Sodomam et Gomorram,et facti estis quasi torrisraptus ab incendio;sed non redistis ad me ",dicit Dominus.
AMOS|4|12|Quapropter haec faciam tibi, Israel,et quia haec faciam tibi,praeparare in occursum Dei tui, Israel;
AMOS|4|13|quia ecce formans montes et creans ventumet annuntians homini cogitationem eius,faciens auroram et tenebraset gradiens super excelsa terrae;Dominus, Deus exercituum, nomen eius.
AMOS|5|1|Audite verbum istud,quod ego levo super vos,planctum, domus Israel:
AMOS|5|2|Cecidit, non adiciet ut resurgatvirgo Israel;proiecta est in terram suam,non est qui suscitet eam.
AMOS|5|3|Quia haec dicit Dominus Deus: Urbs, de qua egrediebantur mille,relinquentur in ea centum;et de qua egrediebantur centum,relinquentur in ea decempro domo Israel ".
AMOS|5|4|Quia haec dicit Dominus domui Israel: Quaerite me et vivetis;
AMOS|5|5|et nolite quaerere Bethelet in Galgalam nolite intrareet in Bersabee nolite transire,quia Galgala captiva ducetur,et Bethel erit iniquitas ".
AMOS|5|6|Quaerite Dominum et vivite;ne forte invadat sicut ignisdomum Ioseph,et devoret, et non sitqui exstinguat Bethel.
AMOS|5|7|Qui convertunt in absinthium iudiciumet iustitiam in terram deiciunt.
AMOS|5|8|Qui facit stellas Pliadis et Orionemet convertit in mane tenebraset diem in noctem obscurat;qui vocat aquas mariset effundit eas super faciem terrae;Dominus nomen eius.
AMOS|5|9|Qui micare facit vastitatem super robustumet vastitatem super arcem affert.
AMOS|5|10|Odio habuerunt corripientem in portaet loquentem perfecte abominati sunt.
AMOS|5|11|Idcirco, pro eo quod conculcastis pauperemet portionem frumenti abstulistis ab eo,domos quadro lapide aedificastiset non habitabitis in eis,vineas plantastis amantissimaset non bibetis vinum earum.
AMOS|5|12|Quia cognovi multa scelera vestraet fortia peccata vestra,opprimentes iustum, accipientes munuset pauperes deprimentes in porta.
AMOS|5|13|Ideo prudens in tempore illo tacet,quia tempus malum est.
AMOS|5|14|Quaerite bonum et non malum,ut vivatis,ita ut sit Dominus, Deus exercituum,vobiscum, sicut dixistis.
AMOS|5|15|Odite malum et diligite bonumet constituite in porta iudicium,si forte misereatur Dominus, Deus exercituum,reliquiis Ioseph.
AMOS|5|16|Propterea haec dicit Dominus,Deus exercituum, dominator: In omnibus plateis planctus,et in cunctis viis dicetur: "Vae, vae!";et vocabunt agricolam ad luctumet ad planctum eos, qui sciunt lamentationem.
AMOS|5|17|Et in omnibus vineis erit luctus,quia pertransibo in medio tui ",dicit Dominus.
AMOS|5|18|Vae desiderantibus diem Domini!Ad quid vobis dies Domini?Tenebrae et non lux.
AMOS|5|19|Quomodo si fugiat vir a facie leonis,et occurrat ei ursus;et ingrediatur domumet innitatur manu sua super parietem,et mordeat eum coluber.
AMOS|5|20|Numquid non tenebrae dies Domini et non lux?Et caligo sine splendore in ea?
AMOS|5|21|" Odi, proieci festivitates vestraset non delector coetibus vestris.
AMOS|5|22|Quod si obtuleritis mihi holocautomata,oblationes vestras non suscipiamet sacrificia pinguium vestrorum non respiciam.
AMOS|5|23|Aufer a me tumultum carminum tuorum,et canticum lyrarum tuarum non audiam.
AMOS|5|24|Et affluat quasi aqua iudicium,et iustitia quasi torrens perennis.
AMOS|5|25|Numquid hostias et oblationes obtulistis mihi in desertoquadraginta annis, domus Israel?
AMOS|5|26|Et portastis Saccut regem vestrum,et Caivan, imagines vestras,sidus deorum vestrorum, quae fecistis vobis.
AMOS|5|27|Et migrare vos faciam trans Damascum ",dicit Dominus; Deus exercituum nomen eius.
AMOS|6|1|Vae, qui tranquilli sunt in Sionet confidunt in monte Samariae;designati primitiae populorum,ad quos venit domus Israel!
AMOS|6|2|Transite in Chalanne et videte;et ite inde in Emath magnamet descendite in Geth Palaestinorum.Numquid meliores regnis istis vos,aut latior terminus eorum termino vestro est?
AMOS|6|3|Qui removetis diem malumet appropinquare facitis solium violentiae.
AMOS|6|4|Qui dormiunt in lectis eburneis,recumbentes in stratis suis,comedentes agnos de gregeet vitulos de medio armenti;
AMOS|6|5|canentes ad vocem psalterii,sicut David excogitant sibi vasa cantici;
AMOS|6|6|bibentes vinum in phialis,optimis unguentis delibuti,et non sunt contristati super ruina Ioseph.
AMOS|6|7|Quapropter nunc migrabunt in capite transmigrantium,et auferetur factio lascivientium.
AMOS|6|8|Iuravit Dominus Deus in anima sua,dicit Dominus, Deus exercituum: Detestor ego superbiam Iacobet domos eius odiet tradam civitatem et plenitudinem eius ".
AMOS|6|9|Quod si reliqui fuerintdecem viri in domo una,et ipsi morientur;
AMOS|6|10|et tollet eum propinquus suuset comburet eum, ut efferat ossa de domo,et dicet ei, qui in penetralibus domus est: Numquid adhuc est penes te? ".Et respondebit: "Non est";et dicet ei: "Tace!";non est qui recordetur nominis Domini.
AMOS|6|11|Quia ecce Dominus mandatet percutiet domum maiorem ruiniset domum minorem scissionibus.
AMOS|6|12|Numquid currunt in petris equi,aut aratur mare in bobus,quoniam convertistis in venenum iudiciumet fructum iustitiae in absinthium?
AMOS|6|13|Qui laetantur pro Lodabar,qui dicunt: " Numquid non in fortitudine nostracepimus nobis Carnaim? ".
AMOS|6|14|" Ecce enim suscitabo super vos, domus Israel,dicit Dominus, Deus exercituum, gentem;et oppriment vos ab introitu Emathusque ad torrentem Arabae ".
AMOS|7|1|Haec ostendit mihi Dominus Deus: et ecce, ipse formabat lo custas in principio, cum germinarent serotinae fruges; et ecce fruges serotinae post fruges demessas regis.
AMOS|7|2|Et factum est, cum consummasset comedere herbam terrae, dixi: "Domine Deus, propitius esto, obsecro; quomodo stabit Iacob, quia parvulus est? ".
AMOS|7|3|Misertus est Dominus super hoc. " Non erit ", dixit Dominus Deus.
AMOS|7|4|Haec ostendit mihi Dominus Deus: et ecce, vocabat ad iudicium per ignem Dominus Deus, et devoravit abyssum magnam et comedit simul partem.
AMOS|7|5|Et dixi: " Domine Deus, quiesce, obsecro; quomodo stabit Iacob, quia parvulus est? ".
AMOS|7|6|Misertus est Dominus super hoc. " Sed et istud non erit ", dicit Dominus Deus.
AMOS|7|7|Haec ostendit mihi Dominus Deus: ecce vir stans super murum litum, et in manu eius trulla caementarii.
AMOS|7|8|Et dixit Dominus ad me: " Quid tu vides, Amos? ". Et dixi: " Trullam caementarii ". Et dixit Dominus: "Ecce ego ponam trullam in medio populi mei Israel; non adiciam ultra ignoscere ei.
AMOS|7|9|Et demolientur excelsa Isaac, et sanctuaria Israel desolabuntur, et consurgam super domum Ieroboam in gladio ".
AMOS|7|10|Et misit Amasias sacerdos Bethel ad Ieroboam regem Israel dicens: " Conspiravit contra te Amos in medio domus Israel; non poterit terra sustinere universos sermones eius.
AMOS|7|11|Haec enim dicit Amos: "In gladio morietur Ieroboam, et Israel captivus migrabit de terra sua" ".
AMOS|7|12|Et dixit Amasias ad Amos: " Qui vides, gradere. Fuge in terram Iudae et comede ibi panem et prophetabis ibi;
AMOS|7|13|et in Bethel non adicies ultra ut prophetes, quia sanctuarium regis est, et domus regni est ".
AMOS|7|14|Responditque Amos et dixit ad Amasiam: Non sum prophetaet non sum filius prophetae;sed armentarius ego sum, vellicans sycomoros.
AMOS|7|15|Et tulit me Dominus,cum sequerer gregem,et dixit Dominus ad me:Vade, propheta ad populum meum Israel".
AMOS|7|16|Et nunc audi verbum Domini. Tu dicis: "Non prophetabis super Israel et non stillabis verba super domum Isaac".
AMOS|7|17|Propter hoc haec dicit Dominus: "Uxor tua in civitate fornicabitur, et filii tui et filiae tuae in gladio cadent, et humus tua funiculo metietur; et tu in terra polluta morieris, et Israel captivus migrabit de terra sua".
AMOS|8|1|Haec ostendit mihi Dominus Deus:et ecce canistrum pomorum.
AMOS|8|2|Et dixit: " Quid tu vides, Amos? ".Et dixi: " Canistrum pomorum ".Et dixit Dominus ad me: Venit finis super populum meum Israel;non adiciam ultra ignoscere ei.
AMOS|8|3|Et lugent cantatrices palatii in die illa,dicit Dominus Deus;multa erunt cadavera,in omni loco proicientur: silentium.
AMOS|8|4|Audite hoc, qui conteritis pauperemet deficere facitis egenos terrae,
AMOS|8|5|dicentes: "Quando transibit neomenia,et venumdabimus merces?Et sabbatum, et aperiemus frumentum,ut imminuamus mensuram et augeamus siclumet supponamus stateras dolosas,
AMOS|8|6|ut possideamus in argento egenoset pauperem pro calceamentiset quisquilias frumenti vendamus?"".
AMOS|8|7|Iuravit Dominus in superbia Iacob: Non obliviscar in perpetuum omnia opera eorum.
AMOS|8|8|Numquid super isto non commovebitur terra,et lugebit omnis habitator eius,et ascendet quasi fluvius universa,fervebit et decrescet quasi flumen Aegypti?
AMOS|8|9|Et erit: in die illa,dicit Dominus Deus,occidere faciam solem in meridieet tenebrescere faciam terram in die luminis
AMOS|8|10|et convertam festivitates vestras in luctumet omnia cantica vestra in planctum;et inducam super omnes lumbos saccumet super omne caput calvitium;et ponam eam quasi luctum unigenitiet novissima eius quasi diem amarum.
AMOS|8|11|Ecce dies veniunt,dicit Dominus,et mittam famem in terram;non famem panis neque sitim aquae,sed audiendi verbum Domini ".
AMOS|8|12|Et fugient a mari usque ad mare;et ab aquilone usque ad orientem circuibunt,quaerentes verbum Domini,et non invenient.
AMOS|8|13|In die illa deficient virgines pulchraeet adulescentes in siti.
AMOS|8|14|Qui iurant in delicto Samariaeet dicunt: " Vivit Deus tuus, Dan! "et " Vivit via, Bersabee! ",et cadent et non resurgent ultra.
AMOS|9|1|Vidi Dominumstantem super altare,et dixit: "Percute capitellum,et commoveantur superliminaria;frange eos in capite omnes,et novissimum eorum in gladio interficiam;non fugiet ex eis fugitivus,et non salvabitur superstes eis.
AMOS|9|2|Si descenderint usque ad infernum,inde manus mea educet eos;et si ascenderint usque in caelum,inde detraham eos.
AMOS|9|3|Et si absconditi fuerint in vertice Carmeli,inde quaeram et auferam eos;et si celaverint se ab oculis meisin profundo maris,ibi mandabo serpenti, et mordebit eos;
AMOS|9|4|et si abierint in captivitatemcoram inimicis suis,ibi mandabo gladio, et occidet eos,et ponam oculos meos super eosin malum et non in bonum ".
AMOS|9|5|Et Dominus, Deus exercituum,qui tangit terram, et tabescet.Et lugebunt omnes habitantes in ea;et ascendet sicut fluvius ea omniset decrescet sicut flumen Aegypti.
AMOS|9|6|Qui aedificat in caelo ascensus suoset cameram suam super terram fundat,qui vocat aquas mariset effundit eas super faciem terrae;Dominus nomen eius.
AMOS|9|7|" Numquid non ut filii Aethiopumvos estis mihi, filii Israel?,ait Dominus.Numquid non Israel ascendere fecide terra Aegyptiet Philisthim de Caphtoret Syros de Cir?
AMOS|9|8|Ecce oculi Domini Deisuper regnum peccans,et conteram illuda facie terrae;verumtamen conterens non conteramdomum Iacob,dicit Dominus.
AMOS|9|9|Ecce enim mandabo egoet concutiam in omnibus gentibus domum Israel,sicut concutitur triticum in cribro,et non cadet lapillus super terram.
AMOS|9|10|In gladio morientur omnes peccatores populi mei,qui dicunt: "Non appropinquabit et non venietsuper nos malum".
AMOS|9|11|In die illa suscitabotabernaculum David, quod cecidit,et reaedificabo rupturas eius;et ea, quae corruerant, instauraboet reaedificabo illud sicut diebus antiquis,
AMOS|9|12|ut possideantreliquias Edomet omnes nationes,super quas invocatum est nomen meum,dicit Dominus, qui faciet haec.
AMOS|9|13|Ecce dies veniunt,dicit Dominus,et comprehendet arator messorem,et calcator uvae mittentem semen; et stillabunt montes mustum,et omnes colles liquefient.
AMOS|9|14|Et convertam captivitatem populi mei Israel;et aedificabunt civitates vastatas et inhabitabuntet plantabunt vineas et bibent vinum earumet facient hortos et comedent fructus eorum.
AMOS|9|15|Et plantabo eos super humum suam,et non evellentur ultrade terra sua, quam dedi eis ",dicit Dominus Deus tuus.
