JOSH|1|1|По смерти Моисея, раба Господня, Господь сказал Иисусу, сыну Навину, служителю Моисееву:
JOSH|1|2|Моисей, раб Мой, умер; итак встань, перейди через Иордан сей, ты и весь народ сей, в землю, которую Я даю им, сынам Израилевым.
JOSH|1|3|Всякое место, на которое ступят стопы ног ваших, Я даю вам, как Я сказал Моисею:
JOSH|1|4|от пустыни и Ливана сего до реки великой, реки Евфрата, всю землю Хеттеев; и до великого моря к западу солнца будут пределы ваши.
JOSH|1|5|Никто не устоит пред тобою во все дни жизни твоей; и как Я был с Моисеем, так буду и с тобою: не отступлю от тебя и не оставлю тебя.
JOSH|1|6|Будь тверд и мужествен; ибо ты народу сему передашь во владение землю, которую Я клялся отцам их дать им;
JOSH|1|7|только будь тверд и очень мужествен, и тщательно храни и исполняй весь закон, который завещал тебе Моисей, раб Мой; не уклоняйся от него ни направо ни налево, дабы поступать благоразумно во всех предприятиях твоих.
JOSH|1|8|Да не отходит сия книга закона от уст твоих; но поучайся в ней день и ночь, дабы в точности исполнять все, что в ней написано: тогда ты будешь успешен в путях твоих и будешь поступать благоразумно.
JOSH|1|9|Вот Я повелеваю тебе: будь тверд и мужествен, не страшись и не ужасайся; ибо с тобою Господь Бог твой везде, куда ни пойдешь.
JOSH|1|10|И дал Иисус повеление надзирателям народа и сказал:
JOSH|1|11|пройдите по стану и дайте повеление народу и скажите: заготовляйте себе пищу для пути, потому что, спустя три дня, вы пойдете за Иордан сей, дабы придти взять землю, которую Господь Бог [отцов] ваших дает вам в наследие.
JOSH|1|12|А колену Рувимову, Гадову и половине колена Манассиина Иисус сказал:
JOSH|1|13|вспомните, что заповедал вам Моисей, раб Господень, говоря: Господь Бог ваш успокоил вас и дал вам землю сию;
JOSH|1|14|жены ваши, дети ваши и скот ваш пусть останутся в земле, которую дал вам Моисей за Иорданом; а вы все, могущие сражаться, вооружившись идите пред братьями вашими и помогайте им,
JOSH|1|15|доколе Господь не успокоит братьев ваших, как и вас; доколе и они не получат в наследие землю, которую Господь Бог ваш дает им; тогда возвратитесь в наследие ваше и владейте землею, которую Моисей, раб Господень, дал вам за Иорданом к востоку солнца.
JOSH|1|16|Они в ответ Иисусу сказали: все, что ни повелишь нам, сделаем, и куда ни пошлешь нас, пойдем;
JOSH|1|17|как слушали мы Моисея, так будем слушать и тебя: только Господь, Бог твой, да будет с тобою, как Он был с Моисеем;
JOSH|1|18|всякий, кто воспротивится повелению твоему и не послушает слов твоих во всем, что ты ни повелишь ему, будет предан смерти. Только будь тверд и мужествен!
JOSH|2|1|И послал Иисус, сын Навин, из Ситтима двух соглядатаев тайно и сказал: пойдите, осмотрите землю и Иерихон. [Два юноши] пошли и пришли в дом блудницы, которой имя Раав, и остались ночевать там.
JOSH|2|2|И сказано было царю Иерихонскому: вот, какие–то люди из сынов Израилевых пришли сюда в эту ночь, чтобы высмотреть землю.
JOSH|2|3|Царь Иерихонский послал сказать Рааве: выдай людей, пришедших к тебе, которые вошли в твой дом, ибо они пришли высмотреть всю землю.
JOSH|2|4|Но женщина взяла двух человек тех и скрыла их и сказала: точно приходили ко мне люди, но я не знала, откуда они;
JOSH|2|5|когда же в сумерки надлежало затворять ворота, тогда они ушли; не знаю, куда они пошли; гонитесь скорее за ними, вы догоните их.
JOSH|2|6|А сама отвела их на кровлю и скрыла их в снопах льна, разложенных у нее на кровле.
JOSH|2|7|[Посланные] гнались за ними по дороге к Иордану до самой переправы; ворота же [тотчас] затворили, после того как вышли погнавшиеся за ними.
JOSH|2|8|Прежде нежели они легли спать, она взошла к ним на кровлю
JOSH|2|9|и сказала им: я знаю, что Господь отдал землю сию вам, ибо вы навели на нас ужас, и все жители земли сей пришли от вас в робость;
JOSH|2|10|ибо мы слышали, как Господь иссушил пред вами воду Чермного моря, когда вы шли из Египта, и как поступили вы с двумя царями Аморрейскими за Иорданом, с Сигоном и Огом, которых вы истребили;
JOSH|2|11|когда мы услышали об этом, ослабело сердце наше, и ни в ком [из нас] не стало духа против вас; ибо Господь Бог ваш есть Бог на небе вверху и на земле внизу;
JOSH|2|12|итак поклянитесь мне Господом что, как я сделала вам милость, так и вы сделаете милость дому отца моего, и дайте мне верный знак,
JOSH|2|13|что вы сохраните в живых отца моего и матерь мою, и братьев моих и сестер моих, и всех, кто есть у них, и избавите души наши от смерти.
JOSH|2|14|Эти люди сказали ей: душа наша вместо вас [да будет предана] смерти, если вы не откроете сего дела нашего; когда же Господь предаст нам землю, мы окажем тебе милость и истину.
JOSH|2|15|И спустила она их по веревке чрез окно, ибо дом ее был в городской стене, и она жила в стене;
JOSH|2|16|и сказала им: идите на гору, чтобы не встретили вас преследующие, и скрывайтесь там три дня, доколе не возвратятся погнавшиеся [за вами]; а после пойдете в путь ваш.
JOSH|2|17|И сказали ей те люди: мы свободны будем от твоей клятвы, которою ты нас закляла, [если не сделаешь так]:
JOSH|2|18|вот, когда мы придем в эту землю, ты привяжи червленую веревку к окну, чрез которое ты нас спустила, а отца твоего и матерь твою и братьев твоих, все семейство отца твоего собери к себе в дом твой;
JOSH|2|19|и если кто–нибудь выйдет из дверей твоего дома вон, того кровь на голове его, а мы свободны [будем от сей клятвы твоей]; а кто будет с тобою в [твоем] доме, того кровь на голове нашей, если чья рука коснется его;
JOSH|2|20|если же ты откроешь сие наше дело, то мы также свободны будем от клятвы твоей, которою ты нас закляла.
JOSH|2|21|Она сказала: да будет по словам вашим! И отпустила их, и они пошли, а она привязала к окну червленую веревку.
JOSH|2|22|Они пошли и пришли на гору, и пробыли там три дня, доколе не возвратились гнавшиеся [за ними]. Гнавшиеся искали их по всей дороге и не нашли.
JOSH|2|23|Таким образом два сии человека пошли назад, сошли с горы, перешли [Иордан] и пришли к Иисусу, сыну Навину, и пересказали ему все, что с ними случилось.
JOSH|2|24|И сказали Иисусу: Господь предал всю землю сию в руки наши, и все жители земли в страхе от нас.
JOSH|3|1|И встал Иисус рано поутру, и двинулись они от Ситтима и пришли к Иордану, он и все сыны Израилевы, и ночевали там, еще не переходя [его].
JOSH|3|2|Чрез три дня пошли надзиратели по стану
JOSH|3|3|и дали народу повеление, говоря: когда увидите ковчег завета Господа Бога вашего и священников [и] левитов, несущих его, то и вы двиньтесь с места своего и идите за ним;
JOSH|3|4|впрочем расстояние между вами и им должно быть до двух тысяч локтей мерою; не подходите к нему близко, чтобы знать вам путь, по которому идти; ибо вы не ходили сим путем ни вчера, ни третьего дня.
JOSH|3|5|И сказал Иисус народу: освятитесь, ибо завтра сотворит Господь среди вас чудеса.
JOSH|3|6|Священникам же сказал Иисус: возьмите ковчег завета, и идите пред народом. [Священники] взяли ковчег завета, и пошли пред народом.
JOSH|3|7|Тогда Господь сказал Иисусу: в сей день Я начну прославлять тебя пред очами всех [сынов] Израиля, дабы они узнали, что как Я был с Моисеем, так буду и с тобою;
JOSH|3|8|а ты дай повеление священникам, несущим ковчег завета, и скажи: как только войдете в воды Иордана, остановитесь в Иордане.
JOSH|3|9|Иисус сказал сынам Израилевым: подойдите сюда и выслушайте слова Господа, Бога вашего.
JOSH|3|10|И сказал Иисус: из сего узнаете, что среди вас есть Бог живый, Который прогонит от вас Хананеев и Хеттеев, и Евеев, и Ферезеев, и Гергесеев, и Аморреев, и Иевусеев:
JOSH|3|11|вот, ковчег завета Господа всей земли пойдет пред вами чрез Иордан;
JOSH|3|12|и возьмите себе двенадцать человек из колен Израилевых, по одному человеку из колена;
JOSH|3|13|и как только стопы ног священников, несущих ковчег Господа, Владыки всей земли, ступят в воду Иордана, вода Иорданская иссякнет, текущая же сверху вода остановится стеною.
JOSH|3|14|Итак, когда народ двинулся от своих шатров, чтобы переходить Иордан, и священники понесли ковчег завета пред народом,
JOSH|3|15|то, лишь только несущие ковчег вошли в Иордан, и ноги священников, несших ковчег, погрузились в воду Иордана – Иордан же выступает из всех берегов своих во все дни жатвы пшеницы, –
JOSH|3|16|вода, текущая сверху, остановилась и стала стеною на весьма большое расстояние, до города Адама, который подле Цартана; а текущая в море равнины, в море Соленое, ушла и иссякла.
JOSH|3|17|И народ переходил против Иерихона; священники же, несшие ковчег завета Господня, стояли на суше среди Иордана твердою ногою. Все [сыны] Израилевы переходили по суше, доколе весь народ не перешел чрез Иордан.
JOSH|4|1|Когда весь народ перешел чрез Иордан, Господь сказал Иисусу:
JOSH|4|2|возьмите себе из народа двенадцать человек, по одному человеку из колена,
JOSH|4|3|и дайте им повеление и скажите: возьмите себе отсюда, из средины Иордана, где стояли ноги священников неподвижно, двенадцать камней, и перенесите их с собою, и положите их на ночлеге, где будете ночевать в эту ночь.
JOSH|4|4|Иисус призвал двенадцать человек, которых назначил из Сынов израилевых, по одному человеку из колена,
JOSH|4|5|и сказал им Иисус: пойдите пред ковчегом Господа Бога вашего в средину Иордана и [возьмите оттуда] и положите на плечо свое каждый по одному камню, по числу колен сынов Израилевых,
JOSH|4|6|чтобы они были у вас знамением; когда спросят вас в последующее время сыны ваши и скажут: "к чему у вас эти камни?",
JOSH|4|7|вы скажете им: "[в память того], что вода Иордана разделилась пред ковчегом завета Господа; когда он переходил чрез Иордан, тогда вода Иордана разделилась"; таким образом камни сии будут для сынов Израилевых памятником на век.
JOSH|4|8|И сделали сыны Израилевы так, как приказал Иисус: взяли двенадцать камней из Иордана, как говорил Господь Иисусу, по числу колен сынов Израилевых, и перенесли их с собою на ночлег, и положили их там.
JOSH|4|9|И [другие] двенадцать камней поставил Иисус среди Иордана на месте, где стояли ноги священников, несших ковчег завета. Они там и до сего дня.
JOSH|4|10|Священники, несшие ковчег, стояли среди Иордана, доколе не окончено было все, что Господь повелел Иисусу сказать народу, так, как завещал Моисей Иисусу; а народ между тем поспешно переходил.
JOSH|4|11|Когда весь народ перешел Иордан, тогда перешел и ковчег [завета] Господня, и священники пред народом;
JOSH|4|12|и сыны Рувима и сыны Гада и половина колена Манассиина перешли вооруженные впереди сынов Израилевых, как говорил им Моисей.
JOSH|4|13|Около сорока тысяч вооруженных на брань перешло пред Господом на равнины Иерихонские, чтобы сразиться.
JOSH|4|14|В тот день прославил Господь Иисуса пред очами всего Израиля и стали бояться его, как боялись Моисея, во все дни жизни его.
JOSH|4|15|И сказал Господь Иисусу, говоря:
JOSH|4|16|прикажи священникам, несущим ковчег откровения, выйти из Иордана.
JOSH|4|17|Иисус приказал священникам и сказал: выйдите из Иордана.
JOSH|4|18|И когда священники, несшие ковчег завета Господня, вышли из Иордана, то, лишь только стопы ног их ступили на сушу, вода Иордана устремилась по своему месту и пошла, как вчера и третьего дня, выше всех берегов своих.
JOSH|4|19|И вышел народ из Иордана в десятый день первого месяца и поставил стан в Галгале, на восточной стороне Иерихона.
JOSH|4|20|И двенадцать камней, которые взяли они из Иордана, Иисус поставил в Галгале
JOSH|4|21|и сказал сынам Израилевым: когда спросят в последующее время сыны ваши отцов своих: "что значат эти камни?",
JOSH|4|22|скажите сынам вашим: "Израиль перешел чрез Иордан сей по суше",
JOSH|4|23|ибо Господь Бог ваш иссушил воды Иордана для вас, доколе вы не перешли его, так же, как Господь Бог ваш сделал с Чермным морем, которое иссушил пред нами, доколе мы не перешли его,
JOSH|4|24|дабы все народы земли познали, что рука Господня сильна, и дабы вы боялись Господа Бога вашего во все дни.
JOSH|5|1|Когда все цари Аморрейские, которые жили по эту сторону Иордана к морю, и все цари Ханаанские, которые при море, услышали, что Господь иссушил воды Иордана пред сынами Израилевыми, доколе переходили они, тогда ослабело сердце их, и не стало уже в них духа против сынов Израилевых.
JOSH|5|2|В то время сказал Господь Иисусу: сделай себе острые ножи и обрежь сынов Израилевых во второй раз.
JOSH|5|3|И сделал себе Иисус острые ножи и обрезал сынов Израилевых на [месте, названном]: Холм обрезания.
JOSH|5|4|Вот причина, почему обрезал Иисус [сынов Израилевых], весь народ, вышедший из Египта, мужеского пола, все способные к войне умерли в пустыне на пути, по исшествии из Египта;
JOSH|5|5|весь же вышедший народ был обрезан, но весь народ, родившийся в пустыне на пути, после того как вышел из Египта, не был обрезан;
JOSH|5|6|ибо сыны Израилевы сорок года ходили в пустыне, доколе не перемер весь народ, способный к войне, вышедший из Египта, которые не слушали гласа Господня, и которым Господь клялся, что они не увидят земли, которую Господь с клятвою обещал отцам их, дать нам землю, где течет молоко и мед,
JOSH|5|7|а вместо их воздвиг сынов их. Сих обрезал Иисус, ибо они были необрезаны; потому что их, на пути, не обрезывали.
JOSH|5|8|Когда весь народ был обрезан, оставался он на своем месте в стане, доколе не выздоровел.
JOSH|5|9|И сказал Господь Иисусу: ныне Я снял с вас посрамление Египетское. Почему и называется то место "Галгал", даже до сего дня.
JOSH|5|10|И стояли сыны Израилевы станом в Галгале и совершили Пасху в четырнадцатый день месяца вечером на равнинах Иерихонских;
JOSH|5|11|и на другой день Пасхи стали есть из произведений земли сей, опресноки и сушеные зерна в самый тот день;
JOSH|5|12|а манна перестала падать на другой день после того, как они стали есть произведения земли, и не было более манны у сынов Израилевых, но они ели в тот год произведения земли Ханаанской.
JOSH|5|13|Иисус, находясь близ Иерихона, взглянул, и видит, и вот стоит пред ним человек, и в руке его обнаженный меч. Иисус подошел к нему и сказал ему: наш ли ты, или из неприятелей наших?
JOSH|5|14|Он сказал: нет; я вождь воинства Господня, теперь пришел [сюда]. Иисус пал лицем своим на землю, и поклонился и сказал ему: что господин мой скажет рабу своему?
JOSH|5|15|Вождь воинства Господня сказал Иисусу: сними обувь твою с ног твоих, ибо место, на котором ты стоишь, свято. Иисус так и сделал.
JOSH|6|1|Иерихон заперся и был заперт от [страха] сынов Израилевых: никто не выходил [из него] и никто не входил.
JOSH|6|2|Тогда сказал Господь Иисусу: вот, Я предаю в руки твои Иерихон и царя его, [и находящихся в нем] людей сильных;
JOSH|6|3|пойдите вокруг города все способные к войне и обходите город однажды [в день]; и это делай шесть дней;
JOSH|6|4|и семь священников пусть несут семь труб юбилейных пред ковчегом; а в седьмой день обойдите вокруг города семь раз, и священники пусть трубят трубами;
JOSH|6|5|когда затрубит юбилейный рог, когда услышите звук трубы, тогда весь народ пусть воскликнет громким голосом, и стена города обрушится до своего основания, и [весь] народ пойдет [в город, устремившись] каждый с своей стороны.
JOSH|6|6|И призвал Иисус, сын Навин, священников [Израилевых] и сказал им: несите ковчег завета; а семь священников пусть несут семь труб юбилейных пред ковчегом Господним.
JOSH|6|7|И сказал народу: пойдите и обойдите вокруг города; вооруженные же пусть идут пред ковчегом Господним.
JOSH|6|8|Как скоро Иисус сказал народу, семь священников, несших семь труб юбилейных пред Господом, пошли и затрубили трубами, и ковчег завета Господня шел за ними;
JOSH|6|9|вооруженные же шли впереди священников, которые трубили трубами; а идущие позади следовали за ковчегом, во время шествия трубя трубами.
JOSH|6|10|Народу же Иисус дал повеление и сказал: не восклицайте и не давайте слышать голоса вашего, и чтобы слово не выходило из уст ваших до [того] дня, доколе я не скажу вам: "воскликните!" и тогда воскликните.
JOSH|6|11|Таким образом ковчег [завета] Господня пошел вокруг города и обошел однажды; и пришли в стан и ночевали в стане.
JOSH|6|12|[На другой день] Иисус встал рано поутру, и священники понесли ковчег [завета] Господня;
JOSH|6|13|и семь священников, несших семь труб юбилейных пред ковчегом Господним, шли и трубили трубами; вооруженные же шли впереди их, а идущие позади следовали за ковчегом [завета] Господня и идучи трубили трубами.
JOSH|6|14|Таким образом и на другой день обошли вокруг города однажды и возвратились в стан. И делали это шесть дней.
JOSH|6|15|В седьмой день встали рано, при появлении зари, и обошли таким же образом вокруг города семь раз; только в этот день обошли вокруг города семь раз.
JOSH|6|16|Когда в седьмой раз священники трубили трубами, Иисус сказал народу: воскликните, ибо Господь предал вам город!
JOSH|6|17|город будет под заклятием, и все, что в нем, Господу; только Раав блудница пусть останется в живых, она и всякий, кто у нее в доме; потому что она укрыла посланных, которых мы посылали;
JOSH|6|18|но вы берегитесь заклятого, чтоб и самим не подвергнуться заклятию, если возьмете что–нибудь из заклятого, и чтобы на стан [сынов] Израилевых не навести заклятия и не сделать ему беды;
JOSH|6|19|и все серебро и золото, и сосуды медные и железные да будут святынею Господу и войдут в сокровищницу Господню.
JOSH|6|20|Народ воскликнул, и затрубили трубами. Как скоро услышал народ голос трубы, воскликнул народ громким голосом, и обрушилась стена [города] до своего основания, и народ пошел в город, каждый с своей стороны, и взяли город.
JOSH|6|21|И предали заклятию все, что в городе, и мужей и жен, и молодых и старых, и волов, и овец, и ослов, [все истребили] мечом.
JOSH|6|22|А двум юношам, высматривавшим землю, Иисус сказал: пойдите в дом оной блудницы и выведите оттуда ее и всех, которые у нее, так как вы поклялись ей.
JOSH|6|23|И пошли юноши, высматривавшие [город, в дом женщины] и вывели Раав и отца ее и мать ее, и братьев ее, и всех, которые у нее [были], и всех родственников ее вывели, и поставили их вне стана Израильского.
JOSH|6|24|А город и все, что в нем, сожгли огнем; только серебро и золото и сосуды медные и железные отдали, в сокровищницу дома Господня.
JOSH|6|25|Раав же блудницу и дом отца ее и всех, которые у нее [были], Иисус оставил в живых, и она живет среди Израиля до сего дня, потому что она укрыла посланных, которых посылал Иисус для высмотрения Иерихона.
JOSH|6|26|В то время Иисус поклялся и сказал: проклят пред Господом тот, кто восставит и построит город сей Иерихон; на первенце своем он положит основание его и на младшем своем поставит врата его.
JOSH|6|27|И Господь был с Иисусом, и слава его носилась по всей земле.
JOSH|7|1|Но сыны Израилевы сделали преступление [и взяли] из заклятого. Ахан, сын Хармия, сына Завдия, сына Зары, из колена Иудина, взял из заклятого, и гнев Господень возгорелся на сынов Израиля.
JOSH|7|2|Иисус из Иерихона послал людей в Гай, что близ Беф–Авена, с восточной стороны Вефиля, и сказал им: пойдите, осмотрите землю. Они пошли и осмотрели Гай.
JOSH|7|3|И возвратившись к Иисусу, сказали ему: не весь народ пусть идет, а пусть пойдет около двух тысяч или около трех тысяч человек, и поразят Гай; всего народа не утруждай туда, ибо их мало [там].
JOSH|7|4|Итак пошло туда из народа около трех тысяч человек, но они обратились в бегство от жителей Гайских;
JOSH|7|5|жители Гайские убили из них до тридцати шести человек, и преследовали их от ворот до Севарим и разбили их на спуске с горы; отчего сердце народа растаяло и стало, как вода.
JOSH|7|6|Иисус разодрал одежды свои и пал лицем своим на землю пред ковчегом Господним [и лежал] до самого вечера, он и старейшины Израилевы, и посыпали прахом головы свои.
JOSH|7|7|И сказал Иисус: о, Господи Владыка! для чего Ты перевел народ сей чрез Иордан, дабы предать нас в руки Аморреев и погубить нас? о, если бы мы остались и жили за Иорданом!
JOSH|7|8|О, Господи! что сказать мне после того, как Израиль обратил тыл врагам своим?
JOSH|7|9|Хананеи и все жители земли услышат и окружат нас и истребят имя наше с земли. И что сделаешь [тогда] имени Твоему великому?
JOSH|7|10|Господь сказал Иисусу: встань, для чего ты пал на лице твое?
JOSH|7|11|Израиль согрешил, и преступили они завет Мой, который Я завещал им; и взяли из заклятого, и украли, и утаили, и положили между своими вещами;
JOSH|7|12|за то сыны Израилевы не могли устоять пред врагами своими и обратили тыл врагам своим, ибо они подпали заклятию; не буду более с вами, если не истребите из среды вашей заклятого.
JOSH|7|13|Встань, освяти народ и скажи: освятитесь к утру, ибо так говорит Господь Бог Израилев: "заклятое среди тебя, Израиль; посему ты не можешь устоять пред врагами твоим, доколе не отдалишь от себя заклятого";
JOSH|7|14|завтра подходите [все] по коленам вашим; колено же, которое укажет Господь, пусть подходит по племенам; племя, которое укажет Господь, пусть подходит по семействам; семейство, которое укажет Господь, пусть подходит по одному человеку;
JOSH|7|15|и обличенного в [похищении] заклятого пусть сожгут огнем, его и все, что у него, за то, что он преступил завет Господень и сделал беззаконие среди Израиля.
JOSH|7|16|Иисус, встав рано поутру, велел подходить Израилю по коленам его, и указано колено Иудино;
JOSH|7|17|потом велел подходить племенам Иуды, и указано племя Зары; велел подходить племени Зарину по семействам, и указано [семейство] Завдиево;
JOSH|7|18|велел подходить семейству его по одному человеку, и указан Ахан, сын Хармия, сына Завдия, сына Зары, из колена Иудина.
JOSH|7|19|Тогда Иисус сказал Ахану: сын мой! воздай славу Господу, Богу Израилеву и сделай пред Ним исповедание и объяви мне, что ты сделал; не скрой от меня.
JOSH|7|20|В ответ Иисусу Ахан сказал: точно, я согрешил пред Господом Богом Израилевым и сделал то и то:
JOSH|7|21|между добычею увидел я одну прекрасную Сеннаарскую одежду и двести сиклей серебра и слиток золота весом в пятьдесят сиклей; это мне полюбилось и я взял это; и вот, оно спрятано в земле среди шатра моего, и серебро под ним.
JOSH|7|22|Иисус послал людей, и они побежали в шатер; и вот, [все] это спрятано было в шатре его, и серебро под ним.
JOSH|7|23|Они взяли это из шатра и принесли к Иисусу и ко всем сынам Израилевым и положили пред Господом.
JOSH|7|24|Иисус и все Израильтяне с ним взяли Ахана, сына Зарина, и серебро, и одежду, и слиток золота, и сыновей его и дочерей его, и волов его и ослов его, и овец его и шатер его, и все, что у него [было], и вывели их на долину Ахор.
JOSH|7|25|И сказал Иисус: за то, что ты навел на нас беду, Господь на тебя наводит беду в день сей. И побили его все Израильтяне камнями, и сожгли их огнем, и наметали на них камни.
JOSH|7|26|И набросали на него большую груду камней, [которая уцелела] и до сего дня. После сего утихла ярость гнева Господня. Посему то место называется долиною Ахор даже до сего дня.
JOSH|8|1|Господь сказал Иисусу: не бойся и не ужасайся; возьми с собою весь народ, способный к войне, и встав пойди к Гаю; вот, Я предаю в руки твои царя Гайского и народ его, город его и землю его;
JOSH|8|2|сделай с Гаем и царем его то же, что сделал ты с Иерихоном и царем его, только добычу его и скот его разделите себе; сделай засаду позади города.
JOSH|8|3|Иисус и весь народ, способный к войне, встал, чтобы идти к Гаю, и выбрал Иисус тридцать тысяч человек храбрых и послал их ночью,
JOSH|8|4|и дал им приказание и сказал: смотрите, вы будете составлять засаду у города позади города; не отходите далеко от города и будьте все готовы;
JOSH|8|5|а я и весь народ, который со мною, подойдем к городу; и когда [жители Гая] выступят против нас, как и прежде, то мы побежим от них;
JOSH|8|6|они пойдут за нами, так что мы отвлечем их от города; ибо они скажут: "бегут от нас, как и прежде"; когда мы побежим от них,
JOSH|8|7|тогда вы встаньте из засады и завладейте городом, и Господь Бог ваш предаст его в руки ваши;
JOSH|8|8|когда возьмете город, зажгите город огнем, по слову Господню сделайте; смотрите, я повелеваю вам.
JOSH|8|9|Таким образом послал их Иисус, и они пошли в засаду и засели между Вефилем и между Гаем, с западной стороны Гая; а Иисус в ту ночь ночевал среди народа.
JOSH|8|10|Встав рано поутру, Иисус осмотрел народ, и пошел он и старейшины Израилевы впереди народа к Гаю;
JOSH|8|11|и весь народ, способный к войне, который был с ним, пошел, приблизился и подошел к городу,
JOSH|8|12|и поставил стан с северной стороны Гая, а между ним и Гаем была долина. Потом взял он около пяти тысяч человек и посадил их в засаде между Вефилем и Гаем, с западной стороны города.
JOSH|8|13|И народ расположил весь стан, который был с северной стороны города, так, что задняя часть была с западной стороны города. И пришел Иисус в ту ночь на средину долины.
JOSH|8|14|Когда увидел это царь Гайский, тотчас с жителями города, встав рано, выступил против Израиля на сражение, он и весь народ его, на назначенное место пред равниною; а он не знал, что для него есть засада позади города.
JOSH|8|15|Иисус и весь Израиль, будто пораженные ими, побежали к пустыне;
JOSH|8|16|а они кликнули весь народ, который был в городе, чтобы преследовать их, и, преследуя Иисуса, отдалились от города;
JOSH|8|17|в Гае и Вефиле не осталось ни одного человека, который не погнался бы за Израилем; и город свой они оставили отворенным, преследуя Израиля.
JOSH|8|18|Тогда Господь сказал Иисусу: простри копье, которое в руке твоей, к Гаю, ибо Я предам его в руки твои. Иисус простер копье, которое было в его руке, к городу.
JOSH|8|19|Сидевшие в засаде тотчас встали с места своего и побежали, как скоро он простер руку свою, вошли в город и взяли его и тотчас зажгли город огнем.
JOSH|8|20|Жители Гая, оглянувшись назад, увидели, что дым от города восходил к небу. И не было для них места, куда бы бежать – ни туда, ни сюда; ибо народ, бежавший к пустыне, обратился на преследователей.
JOSH|8|21|Иисус и весь Израиль, увидев, что сидевшие в засаде взяли город, и дым от города восходил [к небу], возвратились и стали поражать жителей Гая;
JOSH|8|22|а те из города вышли навстречу им, так что они находились в средине между Израильтянами, [из которых] одни были с той стороны, а другие с другой; так поражали их, что не оставили ни одного из них, уцелевшего или убежавшего;
JOSH|8|23|а царя Гайского взяли живого и привели его к Иисусу.
JOSH|8|24|Когда Израильтяне перебили всех жителей Гая на поле, в пустыне, куда они преследовали их, и когда все они до последнего пали от острия меча, тогда все Израильтяне обратились к Гаю и поразили его острием меча.
JOSH|8|25|Падших в тот день мужей и жен, всех жителей Гая, было двенадцать тысяч.
JOSH|8|26|Иисус не опускал руки своей, которую простер с копьем, доколе не предал заклятию всех жителей Гая;
JOSH|8|27|только скот и добычу города сего [сыны] Израиля разделили между собою, по слову Господа, которое [Господь] сказал Иисусу.
JOSH|8|28|И сожег Иисус Гай и обратил его в вечные развалины, в пустыню, до сего дня;
JOSH|8|29|а царя Гайского повесил на дереве, до вечера; по захождении же солнца приказал Иисус, и сняли труп его с дерева, и бросили его у ворот городских, и набросали над ним большую груду камней, [которая уцелела] даже до сего дня.
JOSH|8|30|Тогда Иисус устроил жертвенник Господу Богу Израилеву на горе Гевал,
JOSH|8|31|как заповедал Моисей, раб Господень, сынам Израилевым, о чем написано в книге закона Моисеева, – жертвенник из камней цельных, на которые не поднимали железа; и принесли на нем всесожжение Господу и совершили жертвы мирные.
JOSH|8|32|И написал [Иисус] там на камнях список с закона Моисеева, который он написал пред сынами Израилевыми.
JOSH|8|33|Весь Израиль, старейшины его и надзиратели [его] и судьи его, стали с той и другой стороны ковчега против священников [и] левитов, носящих ковчег завета Господня, как пришельцы, так и природные жители, одна половина их у горы Гаризим, а другая половина у горы Гевал, как прежде повелел Моисей, раб Господень, благословлять народ Израилев.
JOSH|8|34|И потом прочитал [Иисус] все слова закона, благословение и проклятие, как написано в книге закона;
JOSH|8|35|из всего, что Моисей заповедал [Иисусу], не было [ни одного] слова, которого Иисус не прочитал бы пред всем собранием Израиля, и женами, и детьми, и пришельцами, находившимися среди них.
JOSH|9|1|Услышав сие, все цари, которые за Иорданом, на горе и на равнине и по всему берегу великого моря, близ Ливана, Хеттеи, Аморреи, Хананеи, Ферезеи, Евеи и Иевусеи,
JOSH|9|2|собрались вместе, дабы единодушно сразиться с Иисусом и Израилем.
JOSH|9|3|Но жители Гаваона, услышав, что Иисус сделал с Иерихоном и Гаем,
JOSH|9|4|употребили хитрость: пошли, запаслись хлебом на дорогу и положили ветхие мешки на ослов своих и ветхие, изорванные и заплатанные мехи вина;
JOSH|9|5|и обувь на ногах их была ветхая с заплатами, и одежда на них ветхая; и весь дорожный хлеб их был сухой и заплесневелый.
JOSH|9|6|Они пришли к Иисусу в стан [Израильский] в Галгал и сказали ему и всем Израильтянам: из весьма дальней земли пришли мы; итак заключите с нами союз.
JOSH|9|7|Израильтяне же сказали Евеям: может быть, вы живете близ нас? как нам заключить с вами союз?
JOSH|9|8|Они сказали Иисусу: мы рабы твои. Иисус же сказал им: кто вы и откуда пришли?
JOSH|9|9|Они сказали ему: из весьма дальней земли пришли рабы твои во имя Господа Бога твоего; ибо мы слышали славу Его и все, что сделал Он в Египте,
JOSH|9|10|и все, что Он сделал двум царям Аморрейским, которые по ту сторону Иордана, Сигону, царю Есевонскому, и Огу, царю Васанскому, который [жил] в Астарофе.
JOSH|9|11|[Слыша сие], старейшины наши и все жители нашей земли сказали нам: возьмите в руки ваши хлеба на дорогу и пойдите навстречу им и скажите им: "мы рабы ваши; итак заключите с нами союз".
JOSH|9|12|Этот хлеб наш из домов наших мы взяли теплый в тот день, когда пошли к вам, а теперь вот, он сделался сухой и заплесневелый;
JOSH|9|13|и эти мехи с вином, которые мы налили новые, вот, изорвались; и эта одежда наша и обувь наша обветшала от весьма дальней дороги.
JOSH|9|14|Израильтяне взяли их хлеба, а Господа не вопросили.
JOSH|9|15|И заключил Иисус с ними мир и постановил с ними условие в том, что он сохранит им жизнь; и поклялись им начальники общества.
JOSH|9|16|А чрез три дня, как заключили они с ними союз, услышали, что они соседи их и живут близ них;
JOSH|9|17|ибо сыны Израилевы, отправившись в путь, пришли в города их на третий день; города же их [были]: Гаваон, Кефира, Беероф и Кириаф–Иарим.
JOSH|9|18|сыны Израилевы не побили их, потому что начальники общества клялись им Господом Богом Израилевым. За это все общество [Израилево] возроптало на начальников.
JOSH|9|19|Все начальники сказали всему обществу: мы клялись им Господом Богом Израилевым и потому не можем коснуться их;
JOSH|9|20|а вот что сделаем с ними: оставим их в живых, чтобы не постиг нас гнев за клятву, которою мы клялись им.
JOSH|9|21|И сказали им начальники: пусть они живут, но будут рубить дрова и черпать воду для всего общества. [И сделало все общество] так, как сказали им начальники.
JOSH|9|22|Иисус призвал их и сказал: для чего вы обманули нас, сказав: "мы весьма далеко от вас", тогда как вы живете близ нас?
JOSH|9|23|за это прокляты вы! без конца вы будете рабами, будете рубить дрова и черпать воду для дома Бога моего!
JOSH|9|24|Они в ответ Иисусу сказали: дошло до сведения рабов твоих, что Господь Бог твой повелел Моисею, рабу Своему, дать вам всю землю и погубить всех жителей сей земли пред лицем вашим; посему мы весьма боялись, чтобы вы не лишили нас жизни, и сделали это дело;
JOSH|9|25|теперь вот мы в руке твоей: как лучше и справедливее тебе покажется поступить с нами, так и поступи.
JOSH|9|26|И поступил с ними так: избавил их от руки сынов Израилевых, и они не умертвили их;
JOSH|9|27|и определил в тот день Иисус, чтобы они рубили дрова и черпали воду для общества и для жертвенника Господня; – посему жители Гаваона сделались дровосеками и водоносами для жертвенника Божия, – даже до сего дня, на месте, какое ни избрал бы [Господь].
JOSH|10|1|Когда Адониседек, царь Иерусалимский, услышал, что Иисус взял Гай и предал его заклятию, и что так же поступил с Гаем и царем его, как поступил с Иерихоном и царем его, и что жители Гаваона заключили мир с Израилем и остались среди их,
JOSH|10|2|тогда он весьма испугался, потому что Гаваон [был] город большой, как один из царских городов, и больше Гая, и все жители его люди храбрые.
JOSH|10|3|Посему Адониседек, царь Иерусалимский, послал к Гогаму, царю Хевронскому, и к Фираму, царю Иармуфскому, и к Яфию, царю Лахисскому, и к Девиру, царю Еглонскому, чтобы сказать:
JOSH|10|4|придите ко мне и помогите мне поразить Гаваон за то, что он заключил мир с Иисусом и сынами Израилевыми.
JOSH|10|5|Они собрались, и пошли пять царей Аморрейских: царь Иерусалимский, царь Хевронский, царь Иармуфский, царь Лахисский, царь Еглонский, они и все ополчение их, и расположились станом подле Гаваона, чтобы воевать против него.
JOSH|10|6|Жители Гаваона послали к Иисусу в стан [Израильский], в Галгал, сказать: не отними руки твоей от рабов твоих; приди к нам скорее, спаси нас и подай нам помощь; ибо собрались против нас все цари Аморрейские, живущие на горах.
JOSH|10|7|Иисус пошел из Галгала сам, и с ним весь народ, способный к войне, и все мужи храбрые.
JOSH|10|8|И сказал Господь Иисусу: не бойся их, ибо Я предал их в руки твои: никто из них не устоит пред лицем твоим.
JOSH|10|9|И пришел на них Иисус внезапно, [потому что] всю ночь шел он из Галгала.
JOSH|10|10|Господь привел их в смятение при виде Израильтян, и они поразили их в Гаваоне сильным поражением, и преследовали их по дороге к возвышенности Вефорона, и поражали их до Азека и до Македа.
JOSH|10|11|Когда же они бежали от Израильтян по скату горы Вефоронской, Господь бросал на них с небес большие камни до самого Азека, и они умирали; больше было тех, которые умерли от камней града, нежели тех, которых умертвили сыны Израилевы мечом.
JOSH|10|12|Иисус воззвал к Господу в тот день, в который предал Господь Аморрея в руки Израилю, когда побил их в Гаваоне, и они побиты были пред лицем сынов Израилевых, и сказал пред Израильтянами: стой, солнце, над Гаваоном, и луна, над долиною Аиалонскою!
JOSH|10|13|И остановилось солнце, и луна стояла, доколе народ мстил врагам своим. Не это ли написано в книге Праведного: "стояло солнце среди неба и не спешило к западу почти целый день"?
JOSH|10|14|И не было такого дня ни прежде ни после того, в который Господь [так] слушал бы гласа человеческого. Ибо Господь сражался за Израиля.
JOSH|10|15|Потом возвратился Иисус и весь Израиль с ним в стан, в Галгал.
JOSH|10|16|А те пять царей убежали и скрылись в пещере в Македе.
JOSH|10|17|Когда донесено было Иисусу и сказано: "нашлись пять царей, они скрываются в пещере в Македе",
JOSH|10|18|Иисус сказал: "привалите большие камни к отверстию пещеры и приставьте к ней людей стеречь их;
JOSH|10|19|а вы не останавливайтесь, но преследуйте врагов ваших и истребляйте заднюю часть войска их и не давайте им уйти в города их, ибо Господь Бог ваш предал их в руки ваши".
JOSH|10|20|После того, как Иисус и сыны Израилевы совершенно поразили их весьма великим поражением, и оставшиеся из них убежали в города укрепленные,
JOSH|10|21|весь народ возвратился в стан к Иисусу в Макед с миром, и никто на сынов Израилевых не пошевелил языком своим.
JOSH|10|22|Тогда Иисус сказал: откройте отверстие пещеры и выведите ко мне из пещеры пятерых царей тех.
JOSH|10|23|Так и сделали: вывели к нему из пещеры пятерых царей тех: царя Иерусалимского, царя Хевронского, царя Иармуфского, царя Лахисского и царя Еглонского.
JOSH|10|24|Когда вывели царей сих к Иисусу, Иисус призвал всех Израильтян и сказал вождям воинов, ходившим с ним: подойдите, наступите ногами вашими на выи царей сих. Они подошли и наступили ногами своими на выи их.
JOSH|10|25|Иисус сказал им: не бойтесь и не ужасайтесь, будьте тверды и мужественны; ибо так поступит Господь со всеми врагами вашими, с которыми будете воевать.
JOSH|10|26|Потом поразил их Иисус и убил их и повесил их на пяти деревах; и висели они на деревах до вечера.
JOSH|10|27|При захождении солнца приказал Иисус, и сняли их с дерев, и бросили их в пещеру, в которой они скрывались, и привалили большие камни к отверстию пещеры, [которые там] даже до сего дня.
JOSH|10|28|В тот же день взял Иисус Макед, и поразил [его] мечом и царя его, и предал заклятию их и все дышащее, что находилось в нем: никого не оставил, кто бы уцелел; и поступил с царем Македским так же, как поступил с царем Иерихонским.
JOSH|10|29|И пошел Иисус и все Израильтяне с ним из Македа к Ливне и воевал против Ливны;
JOSH|10|30|и предал Господь и ее в руки Израиля, и царя ее, и истребил ее Иисус мечом и все дышащее, что [находилось] в ней: никого не оставил в ней, кто бы уцелел, и поступил с царем ее так же, как поступил с царем Иерихонским.
JOSH|10|31|Из Ливны пошел Иисус и все Израильтяне с ним к Лахису и расположился подле него станом и воевал против него;
JOSH|10|32|и предал Господь Лахис в руки Израиля, и взял он его на другой день, и поразил его мечом и все дышащее, что было в нем, так, как поступил с Ливною.
JOSH|10|33|Тогда пришел на помощь Лахису Горам, царь Газерский; но Иисус поразил его и народ его [мечом] так, что никого у него не оставил, кто бы уцелел.
JOSH|10|34|И пошел Иисус и все Израильтяне с ним из Лахиса к Еглону и расположились подле него станом и воевали против него;
JOSH|10|35|И взяли его в тот же день и поразили его мечом, и все дышащее, что находилось в нем в тот день, предал он заклятию, как поступил с Лахисом.
JOSH|10|36|И пошел Иисус и все Израильтяне с ним из Еглона к Хеврону и воевали против него;
JOSH|10|37|и взяли его и поразили его мечом, и царя его, и все города его, и все дышащее, что находилось в нем; никого не оставил, кто уцелел бы, как поступил он и с Еглоном: предал заклятию его и все дышащее, что находилось в нем.
JOSH|10|38|Потом обратился Иисус и весь Израиль с ним к Давиру и воевал против него;
JOSH|10|39|и взял его и царя его и все города его, и поразили их мечом, и предали заклятию все дышащее, что находилось в нем: никого не осталось, кто уцелел бы; как поступил с Хевроном и царем его, так поступил с Давиром и царем его, и как поступил с Ливною и царем ее.
JOSH|10|40|И поразил Иисус всю землю нагорную и полуденную, и низменные места и землю, лежащую у гор, и всех царей их: никого не оставил, кто уцелел бы, и все дышащее предал заклятию, как повелел Господь Бог Израилев;
JOSH|10|41|поразил их Иисус от Кадес–Варни до Газы, и всю землю Гошен даже до Гаваона;
JOSH|10|42|и всех царей сих и земли их Иисус взял одним разом, ибо Господь Бог Израилев сражался за Израиля.
JOSH|10|43|Потом Иисус и все Израильтяне с ним возвратились в стан, в Галгал.
JOSH|11|1|Услышав [сие], Иавин, царь Асорский, послал к Иоваву, царю Мадонскому, и к царю Шимронскому, и к царю Ахсафскому,
JOSH|11|2|и к царям, которые [жили] к северу на горе и на равнине с южной стороны Хиннарофа, и на низменных местах, и в Нафоф–Доре к западу,
JOSH|11|3|к Хананеям, [которые жили] к востоку и к морю, к Аморреям и Хеттеям, к Ферезеям и к Иевусеям, [жившим] на горе, и к Евеям, [жившим] подле Ермона в земле Массифе.
JOSH|11|4|И выступили они и все ополчение их с ними, многочисленный народ, который множеством равнялся песку на берегу морском; и коней и колесниц [было] весьма много.
JOSH|11|5|И собрались все цари сии, и пришли и расположились станом вместе при водах Меромских, чтобы сразиться с Израилем.
JOSH|11|6|Но Господь сказал Иисусу: не бойся их, ибо завтра, около сего времени, Я предам всех [их] на избиение [сынам] Израиля; коням же их перережь жилы и колесницы их сожги огнем.
JOSH|11|7|Иисус и с ним весь народ, способный к войне, внезапно вышли на них к водам Меромским и напали на них.
JOSH|11|8|И предал их Господь в руки Израильтян, и поразили они их, и преследовали их до Сидона великого и до Мисрефоф–Маима, и до долины Мицфы к востоку, и перебили их, так что никого из них не осталось, кто уцелел бы.
JOSH|11|9|И поступил Иисус с ними так, как сказал ему Господь: коням их перерезал жилы и колесницы их сожег огнем.
JOSH|11|10|В то же время возвратившись Иисус взял Асор и царя его убил мечом (Асор же прежде был главою всех царств сих);
JOSH|11|11|и побили все дышащее, что было в нем, мечом, предав заклятию: не осталось ни одной души; а Асор сожег он огнем.
JOSH|11|12|И все города царей сих и всех царей их взял Иисус и побил мечом, предав их заклятию, как повелел Моисей, раб Господень;
JOSH|11|13|впрочем всех городов, лежавших на возвышенности, не жгли Израильтяне, кроме одного Асора, [который] сжег Иисус.
JOSH|11|14|А всю добычу городов сих и скот разграбили сыны Израилевы себе; людей же всех перебили мечом, так что истребили [всех] их: не оставили ни одной души.
JOSH|11|15|Как повелел Господь Моисею, рабу Своему, так Моисей заповедал Иисусу, а Иисус так и сделал: не отступил ни от одного слова во всем, что повелел Господь Моисею.
JOSH|11|16|Таким образом Иисус взял всю эту нагорную землю, всю землю полуденную, всю землю Гошен и низменные места, и равнину и гору Израилеву, и низменные места,
JOSH|11|17|от горы Халак, простирающейся к Сеиру, до Ваал–Гада в долине Ливанской, подле горы Ермона, и всех царей их взял, поразил их и убил.
JOSH|11|18|Долгое время вел Иисус войну со всеми сими царями.
JOSH|11|19|Не было города, который заключил бы мир с сынами Израилевыми, кроме Евеев, жителей Гаваона: все взяли они войною;
JOSH|11|20|ибо от Господа было то, что они ожесточили сердце свое и войною встречали Израиля – для того, чтобы преданы были заклятию и чтобы не было им помилования, но чтобы истреблены были так, как повелел Господь Моисею.
JOSH|11|21|В то же время пришел Иисус и поразил Енакимов на горе, в Хевроне, в Давире, в Анаве, на всей горе Иудиной и на всей горе Израилевой; с городами их предал их Иисус заклятию;
JOSH|11|22|не осталось [ни одного] из Енакимов в земле сынов Израилевых, остались только в Газе, в Гефе и в Азоте.
JOSH|11|23|Таким образом взял Иисус всю землю, как говорил Господь Моисею, и отдал ее Иисусу в удел Израильтянам, по разделению между коленами их. И успокоилась земля от войны.
JOSH|12|1|Вот цари той земли, которых поразили сыны Израилевы и которых землю взяли в наследие по ту сторону Иордана к востоку солнца, от потока Арнона до горы Ермона, и всю равнину к востоку:
JOSH|12|2|Сигон, царь Аморрейский, живший в Есевоне, владевший от Ароера, что при береге потока Арнона, и от средины потока, половиною Галаада, до потока Иавока, предела Аммонитян,
JOSH|12|3|и равниною до самого моря Хиннерефского к востоку и до моря равнины, моря Соленого, к востоку по дороге к Беф–Иешимофу, а к югу местами, лежащими при подошве Фасги;
JOSH|12|4|сопредельный [ему] Ог, царь Васанский, последний из Рефаимов, живший в Астарофе и в Едреи,
JOSH|12|5|владевший горою Ермоном и Салхою и всем Васаном, до предела Гессурского и Маахского, и половиною Галаада, до предела Сигона, царя Есевонского.
JOSH|12|6|Моисей, раб Господень, и сыны Израилевы убили их; и дал ее Моисей, раб Господень, в наследие [колену] Рувимову и Гадову и половине колена Манассиина.
JOSH|12|7|И вот цари [Аморрейской] земли, которых поразил Иисус и сыны Израилевы по эту сторону Иордана к западу, от Ваал–Гада на долине Ливанской до Халака, горы, простирающейся к Сеиру, которую отдал Иисус коленам Израилевым в наследие, по разделению их,
JOSH|12|8|на горе, на низменных местах, на равнине, на местах, лежащих при горах, и в пустыне и на юге, Хеттеев, Аморреев, Хананеев, Ферезеев, Евеев и Иевусеев:
JOSH|12|9|один царь Иерихона, один царь Гая, что близ Вефиля,
JOSH|12|10|один царь Иерусалима, один царь Хеврона,
JOSH|12|11|один царь Иармуфа, один царь Лахиса,
JOSH|12|12|один царь Еглона, один царь Газера,
JOSH|12|13|один царь Давира, один царь Гадера,
JOSH|12|14|один царь Хормы, один царь Арада,
JOSH|12|15|один царь Ливны, один царь Одоллама,
JOSH|12|16|один царь Македа, один царь Вефиля,
JOSH|12|17|один царь Таппуаха, один царь Хефера.
JOSH|12|18|Один царь Афека, один царь Шарона,
JOSH|12|19|один царь Мадона, один царь Асора,
JOSH|12|20|один царь Шимрон–Мерона, один царь Ахсафа,
JOSH|12|21|один царь Фаанаха, один царь Мегиддона,
JOSH|12|22|один царь Кедеса, один царь Иокнеама при Кармиле,
JOSH|12|23|один царь Дора при Нафаф–Доре, один царь Гоима в Галгале,
JOSH|12|24|один царь Фирцы. Всех царей тридцать один.
JOSH|13|1|Когда Иисус состарился, вошел в лета [преклонные], тогда Господь сказал ему: ты состарился, вошел в лета [преклонные], а земли брать в наследие остается еще очень много.
JOSH|13|2|Остается сия земля: все округи Филистимские и вся [земля] Гессурская.
JOSH|13|3|От Сихора, что пред Египтом, до пределов Екрона к северу, считаются Ханаанскими пять владельцев Филистимских: Газский, Азотский, Аскалонский, Гефский, Екронский и Аввейский;
JOSH|13|4|к югу же вся земля Ханаанская от Меары Сидонской до Афека, до пределов Аморрейских,
JOSH|13|5|также земля Гевла и весь Ливан к востоку солнца от Ваал–Гада, [что] подле горы Ермона, до входа в Емаф.
JOSH|13|6|Всех горных жителей от Ливана до Мисрефоф–Маима, всех Сидонян Я изгоню от лица сынов Израилевых. Раздели же ее в удел Израилю, как Я повелел тебе;
JOSH|13|7|раздели землю сию в удел девяти коленам и половине колена Манассиина.
JOSH|13|8|А [колено] Рувимово и Гадово с другою половиною колена Манассиина получили удел свой от Моисея за Иорданом к востоку, как дал им Моисей, раб Господень,
JOSH|13|9|от Ароера, который на берегу потока Арнона, и город, который среди потока, и всю равнину Медеву до Дивона;
JOSH|13|10|также все города Сигона, царя Аморрейского, который царствовал в Есевоне, до пределов Аммонитских,
JOSH|13|11|также Галаад и область Гессурскую и Маахскую, и всю гору Ермон и весь Васан до Салхи,
JOSH|13|12|все царство Ога Васанского, который царствовал в Астарофе и в Едреи. Он оставался один из Рефаимов, которых Моисей поразил и прогнал.
JOSH|13|13|Но сыны Израилевы не выгнали жителей Гессура и Маахи, и живет Гессур и Мааха среди Израиля до сего дня.
JOSH|13|14|Только колену Левиину не дал он удела: жертвы Господа Бога Израилева суть удел его, как сказал ему Господь.
JOSH|13|15|колену сынов Рувимовых по племенам их дал [удел] Моисей:
JOSH|13|16|пределом их был Ароер, который на берегу потока Арнона, и город, который среди потока, и вся равнина при Медеве,
JOSH|13|17|Есевон и все города его, которые на равнине, и Дивон, Вамоф–Ваали Беф–Ваал–Меон,
JOSH|13|18|Иааца, Кедемоф и Мефааф,
JOSH|13|19|Кириафаим, Сивма и Цереф–Шахар на горе Емек,
JOSH|13|20|Беф–Фегор и места при подошве Фасги и Беф–Иешимоф,
JOSH|13|21|и все города на равнине, и все царство Сигона, царя Аморрейского, который царствовал в Есевоне, которого убил Моисей, равно как и вождей Мадиамских: Евия, и Рекема, и Цура, и Хура, и Реву, князей Сигоновых, живших в земле [той];
JOSH|13|22|также Валаама, сына Веорова, прорицателя, убили сыны Израилевы мечом в числе убитых ими.
JOSH|13|23|Пределом сынов Рувимовых был Иордан. Вот удел сынов Рувимовых по племенам их, города и села их.
JOSH|13|24|Моисей дал также [удел] колену Гадову, сынам Гадовым, по племенам их:
JOSH|13|25|пределом их был Иазер и все города Галаадские, и половина земли сынов Аммоновых до Ароера, что пред Раввою,
JOSH|13|26|и [земли] от Есевона до Рамаф–Мицфы и Ветонима и от Маханаима до пределов Давира,
JOSH|13|27|и на долине Беф–Гарам и Беф–Нимра и Сокхоф и Цафон, остаток царства Сигона, царя Есевонского; пределом его был Иордан до моря Хиннерефского за Иорданом к востоку.
JOSH|13|28|Вот удел сынов Гадовых по племенам их, города и села их.
JOSH|13|29|Моисей дал [удел] и половине колена Манассиина, который [принадлежал] половине колена сынов Манассииных, по племенам их;
JOSH|13|30|предел их был: от Маханаима весь Васан, все царство Ога, царя Васанского, и все селения Иаировы, что в Васане, шестьдесят городов;
JOSH|13|31|а половина Галаада и Астароф и Едрея, царственные города Ога Васанского, [даны] сынам Махира, сына Манассиина, половине сынов Махировых, по племенам их.
JOSH|13|32|Вот что Моисей дал в удел на равнинах Моавитских за Иорданом против Иерихона к востоку.
JOSH|13|33|Но колену Левиину Моисей не дал удела: Господь Бог Израилев Сам есть удел их, как Он говорил им.
JOSH|14|1|Вот что получили в удел сыны Израилевы в земле Ханаанской, что разделили им в удел Елеазар священник и Иисус, сын Навин, и начальники поколений в коленах сынов Израилевых;
JOSH|14|2|по жребию делили они, как повелел Господь чрез Моисея, девяти коленам и половине колена [Манассиина],
JOSH|14|3|ибо двум коленам и половине колена [Манассиина] Моисей дал удел за Иорданом, левитам же не дал удела между ними;
JOSH|14|4|ибо от сынов Иосифовых произошли два колена: Манассиино и Ефремово; посему они и не дали левитам части в земле, [а только] города для жительства с предместиями их для скота их и для [других] выгод их.
JOSH|14|5|Как повелел Господь Моисею, так [и] сделали сыны Израилевы, когда делили на уделы землю.
JOSH|14|6|Сыны Иудины пришли в Галгал к Иисусу. И сказал ему Халев, сын Иефоннии, Кенезеянин: ты знаешь, что говорил Господь Моисею, человеку Божию, о мне и о тебе в Кадес–Варне;
JOSH|14|7|я был сорока лет, когда Моисей, раб Господень, посылал меня из Кадес–Варни осмотреть землю, и я принес ему в ответ, что было у меня на сердце:
JOSH|14|8|братья мои, которые ходили со мною, привели в робость сердце народа, а я в точности следовал Господу Богу моему;
JOSH|14|9|и клялся Моисей в тот день и сказал: "земля, по которой ходила нога твоя, будет уделом тебе и детям твоим на век, ибо ты в точности последовал Господу Богу моему";
JOSH|14|10|итак, вот, Господь сохранил меня в живых, как Он говорил; уже сорок пять лет [прошло] от того времени, когда Господь сказал Моисею слово сие, и Израиль ходил по пустыне; теперь, вот, мне восемьдесят пять лет;
JOSH|14|11|но и ныне я столько же крепок, как и тогда, когда посылал меня Моисей: сколько тогда было у меня силы, столько и теперь есть для того, чтобы воевать и выходить и входить;
JOSH|14|12|итак дай мне сию гору, о которой говорил Господь в тот день; ибо ты слышал в тот день, что там [живут] сыны Енаковы, и города [у них] большие и укрепленные; может быть, Господь [будет] со мною, и я изгоню их, как говорил Господь.
JOSH|14|13|Иисус благословил его, и дал в удел Халеву, сыну Иефонниину, Хеврон.
JOSH|14|14|Таким образом Хеврон остался уделом Халева, сына Иефонниина, Кенезеянина, до сего дня, за то, что он в точности последовал [повелению] Господа Бога Израилева.
JOSH|14|15|Имя Хеврону прежде было Кириаф–Арбы, как назывался между сынами Енака один человек великий. И земля успокоилась от войны.
JOSH|15|1|Жребий колену сынов Иудиных, по племенам их, выпал такой: в смежности с Идумеею была пустыня Син, к югу, при конце Фемана;
JOSH|15|2|южным пределом их был край моря Соленого от простирающегося к югу залива;
JOSH|15|3|на юге идет он к возвышенности Акраввимской, проходит Цин и, восходя с южной стороны к Кадес–Варне, проходит Хецрон и, восходя до Аддара, поворачивает к Каркае,
JOSH|15|4|потом проходит Ацмон, идет к потоку Египетскому, так что конец сего предела есть море. Сей будет южный ваш предел.
JOSH|15|5|Пределом же к востоку море Соленое, до устья Иордана; а предел с северной стороны [начинается] от залива моря, от устья Иордана;
JOSH|15|6|отсюда предел восходит к Беф–Хогле и проходит с северной стороны к Беф–Араве, и идет предел вверх до камня Богана, сына Рувимова;
JOSH|15|7|потом восходит предел к Давиру от долины Ахор и на севере поворачивает к Галгалу, который против возвышенности Адуммима, лежащего с южной стороны потока; отсюда предел проходит к водам Ен–Шемеша и оканчивается у Ен–Рогела;
JOSH|15|8|отсюда предел идет вверх к долине сына Енномова с южной стороны Иевуса, который [есть] Иерусалим, и восходит предел на вершину горы, которая к западу против долины Енномовой, которая на краю долины Рефаимов к северу;
JOSH|15|9|от вершины горы предел поворачивает к источнику вод Нефтоах и идет к городам горы Ефрона, и поворачивает предел к Ваалу, который [есть] Кириаф–Иарим;
JOSH|15|10|потом поворачивает предел от Ваала к морю к горе Сеиру, и идет северною стороною горы Иеарим, которая [есть] Кесалон, и, нисходя к Вефсамису, проходит чрез Фимну;
JOSH|15|11|отсюда предел идет северною стороною Екрона, и поворачивает предел к Шикарону, проходит чрез гору Ваал и доходит до Иавнеила, и оканчивается предел у моря. Западный предел составляет великое море.
JOSH|15|12|Вот предел сынов Иудиных с племенами их со всех сторон.
JOSH|15|13|И Халеву, сыну Иефонниину, [Иисус] дал часть среди сынов Иудиных, как повелел Господь Иисусу; Кириаф–Арбы, отца Енакова, иначе Хеврон.
JOSH|15|14|И выгнал оттуда Халев трех сынов Енаковых: Шешая, Ахимана и Фалмая, детей Енаковых.
JOSH|15|15|Отсюда пошел против жителей Давира (имя Давиру прежде [было] Кириаф–Сефер).
JOSH|15|16|И сказал Халев: кто поразит Кириаф–Сефер и возьмет его, тому отдам Ахсу, дочь мою, в жену.
JOSH|15|17|И взял его Гофониил, сын Кеназа, брата Халевова, и отдал он в жену ему Ахсу, дочь свою.
JOSH|15|18|Когда надлежало ей идти, ее научили просить у отца ее поле, и она сошла с осла. Халев сказал ей: что тебе?
JOSH|15|19|Она сказала: дай мне благословение; ты дал мне землю полуденную, дай мне и источники вод. И дал он ей источники верхние и источники нижние.
JOSH|15|20|Вот удел колена сынов Иудиных, по племенам их:
JOSH|15|21|города с края колена сынов Иудиных в смежности с Идумеею на юге были: Кавцеил, Едер и Иагур,
JOSH|15|22|Кина, Димона, Адада,
JOSH|15|23|Кедес, Асор и Ифнан,
JOSH|15|24|Зиф, Телем и Валоф,
JOSH|15|25|Гацор–Хадафа, Кириаф, Хецрон, иначе Гацор,
JOSH|15|26|Амам, Шема и Молада,
JOSH|15|27|Хацар–Гадда, Хешмон и Веф–Палет,
JOSH|15|28|Хацар–Шуал, Вирсавия и Визиофея,
JOSH|15|29|Ваала, Иим и Ацем,
JOSH|15|30|Елфолад, Кесил и Хорма,
JOSH|15|31|Циклаг, Мадмана и Сансана,
JOSH|15|32|Леваоф, Шелихим, Аин и Риммон: всех двадцать девять городов с их селами.
JOSH|15|33|На низменных местах: Ештаол, Цора и Ашна,
JOSH|15|34|Заноах, Ен–Ганним, Таппуах и Гаенам,
JOSH|15|35|Иармуф, Одоллам, Сохо и Азека,
JOSH|15|36|Шаараим, Адифаим, Гедера или Гедерофаим: четырнадцать городов с их селами.
JOSH|15|37|Ценан, Хадаша, Мигдал–Гад,
JOSH|15|38|Дилеан, Мицфе и Иокфеил,
JOSH|15|39|Лахис, Воцкаф и Еглон,
JOSH|15|40|Хаббон, Лахмас и Хифлис,
JOSH|15|41|Гедероф, Беф–Дагон, Наема и Макед: шестнадцать городов с их селами.
JOSH|15|42|Ливна, Ефер и Ашан,
JOSH|15|43|Иффах, Ашна и Нецив,
JOSH|15|44|Кеила, Ахзив и Мареша: девять городов с их селами.
JOSH|15|45|Екрон с зависящими от него [городами] и селами его,
JOSH|15|46|и от Екрона к морю все, что находится около Азота, с селами их,
JOSH|15|47|Азот, зависящие от него города и села его, Газа, зависящие от нее города и села ее, до самого потока Египетского и великого моря, которое [есть] предел.
JOSH|15|48|На горах: Шамир, Иаттир и Сохо,
JOSH|15|49|Данна, Кириаф–Санна, иначе Давир,
JOSH|15|50|Анаф, Ештемо и Аним,
JOSH|15|51|Гошен, Холон и Гило: одиннадцать городов с их селами.
JOSH|15|52|Арав, Дума и Ешан,
JOSH|15|53|Ианум, Беф–Таппуах и Афека,
JOSH|15|54|Хумта, Кириаф–Арбы, иначе Хеврон, и Цигор: девять городов с их селами.
JOSH|15|55|Маон, Кармил, Зиф и Юта,
JOSH|15|56|Изреель, Иокдам и Заноах,
JOSH|15|57|Каин, Гива и Фимна: десять городов с их селами.
JOSH|15|58|Халхул, Беф–Цур и Гедор,
JOSH|15|59|Маараф, Беф–Аноф и Елтекон: шесть городов с их селами.
JOSH|15|60|Кириаф–Ваал, иначе Кириаф–Иарим, и Аравва: два города с их селами.
JOSH|15|61|В пустыне: Беф–Арава, Миддин и Секаха,
JOSH|15|62|Нившан, Ир–Мелах и Ен–Геди: шесть городов с их селами.
JOSH|15|63|Но Иевусеев, жителей Иерусалима, не могли изгнать сыны Иудины, и потому Иевусеи живут с сынами Иуды в Иерусалиме даже до сего дня.
JOSH|16|1|Потом выпал жребий сынам Иосифа: от Иордана подле Иерихона, у вод Иерихонских на восток, пустыня, простирающаяся от Иерихона к горе Вефильской;
JOSH|16|2|от Вефиля идет [предел] к Лузу и переходит к пределу Архи до Атарофа,
JOSH|16|3|и спускается к морю, к пределу Иафлета, до предела нижнего Беф–Орона и до Газера, и оканчивается у моря.
JOSH|16|4|Это получили в удел сыны Иосифа: Манассия и Ефрем.
JOSH|16|5|Предел сынов Ефремовых по племенам их был сей: от востока пределом удела их был Атароф–Адар до Беф–Орона верхнего;
JOSH|16|6|потом идет предел к морю северною стороною Михмефафа и поворачивает к восточной стороне Фаанаф–Силома и проходит его с восточной стороны Ианоха;
JOSH|16|7|от Ианоха, нисходя к Атарофу и Наарафу, примыкает к Иерихону и доходит до Иордана;
JOSH|16|8|от Таппуаха идет предел к морю, к потоку Кане, и оканчивается морем. Вот удел колена сынов Ефремовых, по племенам их.
JOSH|16|9|И города отделены сынам Ефремовым в уделе сынов Манассииных, все города с селами их.
JOSH|16|10|Но [Ефремляне] не изгнали Хананеев, живших в Газере; посему Хананеи жили среди Ефремлян до сего дня, платя им дань.
JOSH|17|1|И выпал жребий колену Манассии, так как он был первенец Иосифа. Махиру, первенцу Манассии, отцу Галаада, который [был] храбр на войне, достался Галаад и Васан.
JOSH|17|2|Достались [уделы] и прочим сынам Манассии, по племенам их, и сынам Авиезера, и сынам Хелека, и сынам Асриила, и сынам Шехема, и сынам Хефера, и сынам Шемиды. Вот дети Манассии, сына Иосифова, мужеского пола, по племенам их.
JOSH|17|3|У Салпаада же, сына Хеферова, сына Галаадова, сына Махирова, сына Манассиина, не было сыновей, а [только] дочери. Вот имена дочерей его: Махла, Ноа, Хогла, Милка и Фирца.
JOSH|17|4|Они пришли к священнику Елеазару и к Иисусу, сыну Навину, и к начальникам, и сказали: Господь повелел Моисею дать нам удел между братьями нашими. И дан им удел, по повелению Господню, между братьями отца их.
JOSH|17|5|И выпало Манассии десять участков, кроме земли Галаадской и Васанской, которая за Иорданом;
JOSH|17|6|ибо дочери Манассии получили удел среди сыновей его, а земля Галаадская досталась прочим сыновьям Манассии.
JOSH|17|7|Предел Манассии идет от Асира к Михмефафу, который против Сихема; отсюда предел идет направо к жителям Ен–Таппуаха.
JOSH|17|8|Земля Таппуах досталась Манассии, а [город] Таппуах у предела Манассиина – сынам Ефремовым.
JOSH|17|9|Отсюда предел нисходит к потоку Кане, с южной стороны потока. Города сии [принадлежат] Ефрему, [хотя находятся] среди городов Манассии. Предел Манассии – на северной стороне потока и оканчивается морем.
JOSH|17|10|Что к югу, то Ефремово, а что к северу, то Манассиино; море же было пределом их; к Асиру примыкали они с северной стороны и к Иссахару с восточной.
JOSH|17|11|У Иссахара и Асира [принадлежат] Манассии Беф–Сан и зависящие от него места, Ивлеам и зависящие от него места, жители Дора и зависящие от него места, жители Ен–Дора и зависящие от него места, жители Фаанаха и зависящие от него места, жители Мегиддона и зависящие от него места, и третья часть Нафефа.
JOSH|17|12|Сыны Манассиины не могли выгнать [жителей] городов сих, и Хананеи остались жить в земле сей.
JOSH|17|13|Когда же сыны Израилевы пришли в силу, тогда Хананеев сделали они данниками, но изгнать не изгнали их.
JOSH|17|14|Сыны Иосифа говорили Иисусу и сказали: почему ты дал мне в удел один жребий и один участок, тогда как я многолюден, потому что так благословил меня Господь?
JOSH|17|15|Иисус сказал им: если ты многолюден, то пойди в леса и там, в земле Ферезеев и Рефаимов, расчисти себе [место], если гора Ефремова для тебя тесна.
JOSH|17|16|Сыны Иосифа сказали: не останется за нами гора, потому что железные колесницы у всех Хананеев, живущих на долине, как у тех, которые в Беф–Сане и в зависящих от него местах, так и у тех, которые на долине Изреельской.
JOSH|17|17|Но Иисус сказал дому Иосифову, Ефрему и Манассии: ты многолюден и сила у тебя велика; не один жребий будет у тебя:
JOSH|17|18|и гора будет твоею, и лес сей; ты расчистишь его, и он будет твой до самого конца его; ибо ты изгонишь Хананеев, хотя у них колесницы железные, и хотя они сильны.
JOSH|18|1|Все общество сынов Израилевых собралось в Силом, и поставили там скинию собрания, ибо земля была покорена ими.
JOSH|18|2|Из сынов же Израилевых оставалось семь колен, которые еще не получили удела своего.
JOSH|18|3|И сказал Иисус сынам Израилевым: долго ли вы будете нерадеть о том, чтобы пойти [и] взять в наследие землю, которую дал вам Господь Бог отцов ваших?
JOSH|18|4|дайте от себя по три человека из колена; я пошлю их, и они встав пройдут по земле и опишут ее, как надобно разделить им на уделы, и придут ко мне;
JOSH|18|5|пусть разделят ее на семь уделов; Иуда пусть остается в пределе своем на юге, а дом Иосифов пусть остается в пределе своем на севере;
JOSH|18|6|а вы распишите землю на семь уделов и представьте мне сюда: я брошу вам жребий здесь пред лицем Господа Бога нашего;
JOSH|18|7|а левитам нет части между вами, ибо священство Господне есть удел их; Гад же, Рувим и половина колена Манассиина получили удел свой за Иорданом к востоку, который дал им Моисей, раб Господень.
JOSH|18|8|Эти люди встали и пошли. Иисус же пошедшим описывать землю дал такое приказание: пойдите, обойдите землю, опишите ее и возвратитесь ко мне; а я здесь брошу вам жребий пред лицем Господним, в Силоме.
JOSH|18|9|Они пошли, прошли по земле, и описали ее, по городам ее, на семь уделов, в книге, и пришли к Иисусу в стан, в Силом.
JOSH|18|10|Иисус бросил им жребий в Силоме пред Господом, и разделил там Иисус землю сынам Израилевым по участкам их.
JOSH|18|11|[Первый] жребий вышел колену сынов Вениаминовых, по племенам их. Предел их по жребию шел между сынами Иуды и между сынами Иосифа;
JOSH|18|12|предел их на северной стороне начинается у Иордана, и проходит предел сей подле Иерихона с севера, и восходит на гору к западу, и оканчивается в пустыне Бефавен;
JOSH|18|13|оттуда предел идет к Лузу, к южной стороне Луза, иначе Вефиля, и нисходит предел к Атароф–Адару, к горе, которая на южной стороне Беф–Орона нижнего;
JOSH|18|14|потом предел поворачивает и склоняется к морской стороне на юг от горы, которая на юге пред Беф–Ороном, и оканчивается у Кириаф–Ваала, иначе Кириаф–Иарима, города сынов Иудиных. Это западная сторона.
JOSH|18|15|Южною же стороною от Кириаф–Иарима идет предел к морю и доходит до источника вод Нефтоаха;
JOSH|18|16|потом предел нисходит к концу горы, которая пред долиною сына Енномова, на долине Рефаимов, к северу, и нисходит долиною Еннома к южной стороне Иевуса, и идет к Ен–Рогелу;
JOSH|18|17|потом поворачивает от севера и идет к Ен–Шемешу, и идет к Гелилофу, который против возвышенности Адуммима, и нисходит к камню Богана, сына Рувимова;
JOSH|18|18|потом проходит близ равнины к северу и нисходит на равнину;
JOSH|18|19|отсюда проходит предел подле Беф–Хоглы к северу, и оканчивается предел у северного залива моря Соленого, у южного конца Иордана. Вот предел южный. С восточной же стороны пределом служит Иордан.
JOSH|18|20|Вот удел сынов Вениаминовых, с пределами его со всех сторон, по племенам их.
JOSH|18|21|Города колену сынов Вениаминовых, по племенам их, принадлежали сии: Иерихон, Беф–Хогла и Емек–Кециц,
JOSH|18|22|Беф–Арава, Цемараим и Вефиль,
JOSH|18|23|Аввим, Фара и Офра,
JOSH|18|24|Кефар–Аммонай, Афни и Гева: двенадцать городов с их селами.
JOSH|18|25|Гаваон, Рама и Бероф,
JOSH|18|26|Мицфе, Кефира и Моца,
JOSH|18|27|Рекем, Ирфеил и Фарала,
JOSH|18|28|Цела, Елеф и Иевус, иначе Иерусалим, Гивеаф и Кириаф: четырнадцать городов с их селами. Вот удел сынов Вениаминовых, по племенам их.
JOSH|19|1|Второй жребий вышел Симеону, колену сынов Симеоновых, по племенам их; и был удел их среди удела сынов Иудиных.
JOSH|19|2|В уделе их были: Вирсавия или Шева, Молада,
JOSH|19|3|Хацар–Шуал, Вала и Ацем,
JOSH|19|4|Елтолад, Вефул и Хорма,
JOSH|19|5|Циклаг, Беф–Маркавоф и Хацар–Суса,
JOSH|19|6|Беф–Леваоф и Шарухен: тринадцать городов с их селами.
JOSH|19|7|Аин, Риммон, Ефер и Ашан: четыре города с селами их,
JOSH|19|8|и все села, которые находились вокруг городов сих даже до Ваалаф–Беера, или южной Рамы. Вот удел колена сынов Симеоновых, по племенам их.
JOSH|19|9|От участка сынов Иудиных [выделен] удел [колену] сынов Симеоновых. Так как участок сынов Иудиных был слишком велик для них, то сыны Симеоновы и получили удел среди их удела.
JOSH|19|10|Третий жребий выпал сынам Завулоновым по племенам их, и простирался предел удела их до Сарида;
JOSH|19|11|предел их восходит к морю и Марале и примыкает к Дабешефу и примыкает к потоку, который пред Иокнеамом;
JOSH|19|12|от Сарида идет назад к восточной стороне, к востоку солнца, до предела Кислоф–Фавора; отсюда идет к Даврафу и восходит к Иафие;
JOSH|19|13|отсюда проходит к востоку в Геф–Хефер, в Итту–Кацин, и идет к Риммону, Мифоару и Нее;
JOSH|19|14|и поворачивает предел от севера к Ханнафону и оканчивается долиною Ифтах–Ел;
JOSH|19|15|далее: Каттаф, Нагалал, Шимрон, Идеала и Вифлеем: двенадцать городов с их селами.
JOSH|19|16|Вот удел сынов Завулоновых, по их племенам; вот города и села их.
JOSH|19|17|Четвертый жребий вышел Иссахару, сынам Иссахара, по племенам их;
JOSH|19|18|пределом их был: Изреель, Кесуллоф и Сунем,
JOSH|19|19|Хафараим, Шион и Анахараф,
JOSH|19|20|Раввиф, Кишион и Авец,
JOSH|19|21|Ремеф, Ен–Ганним, Ен–Хадда и Беф–Пацец;
JOSH|19|22|и примыкает предел к Фавору и Шагациме и Вефсамису, и оканчивается предел их у Иордана: шестнадцать городов с селами их.
JOSH|19|23|Вот удел колена сынов Иссахаровых по племенам их; вот города и села их.
JOSH|19|24|Пятый жребий вышел колену сынов Асировых, по племенам их;
JOSH|19|25|пределом их были: Хелкаф, Хали, Ветен и Ахсаф,
JOSH|19|26|Аламелех, Амад и Мишал; и примыкает [предел] к Кармилу с западной стороны и к Шихор–Ливнафу;
JOSH|19|27|потом идет назад к востоку солнца в Беф–Дагон, и примыкает к Завулону и к долине Ифтах–Ел с севера, в Беф–Емек и Неиел, и идет у Кавула, с левой стороны;
JOSH|19|28|далее: Еврон, Рехов, Хаммон и Кана, до Сидона великого;
JOSH|19|29|потом предел возвращается к Раме до укрепленного города Тира, и поворачивает предел к Хоссе, и оканчивается у моря, в местечке Ахзиве;
JOSH|19|30|далее: Умма, Афек и Рехов: двадцать два города с селами их.
JOSH|19|31|Вот удел колена сынов Асировых, по племенам их; вот города и села их.
JOSH|19|32|Шестой жребий вышел сынам Неффалима, сынам Неффалима по племенам их;
JOSH|19|33|предел их шел от Хелефа [и] от дубравы, [что] в Цананниме, к Адами–Некеву и Иавнеилу, до Лаккума, и оканчивался у Иордана;
JOSH|19|34|отсюда возвращается предел на запад к Азноф–Фавору и идет оттуда к Хуккоку, и примыкает к Завулону с юга, и к Асиру примыкает с запада, и к Иуде у Иордана, от востока солнца.
JOSH|19|35|Города укрепленные: Циддим, Цер, Хамаф, Раккаф и Хиннереф,
JOSH|19|36|Адама, Рама и Асор,
JOSH|19|37|Кедес, Едрея и Ен–Гацор,
JOSH|19|38|Иреон, Мигдал–Ел, Хорем, Беф–Анаф и Вефсамис: девятнадцать городов с их селами.
JOSH|19|39|Вот удел колена сынов Неффалимовых по племенам их; вот города и села их.
JOSH|19|40|Колену сынов Дановых, по племенам их, вышел жребий седьмой;
JOSH|19|41|пределом удела их были: Цора, Ештаол и Ир–Шемеш,
JOSH|19|42|Шаалаввин, Аиалон и Ифла,
JOSH|19|43|Елон, Фимнафа и Екрон,
JOSH|19|44|Елтеке, Гиввефон и Ваалаф,
JOSH|19|45|Игуд, Бене–Верак и Гаф–Риммон,
JOSH|19|46|Ме–Иаркон и Ракон с пределом близ Иоппии. И вышел предел сынов Дановых мал для них.
JOSH|19|47|И сыны Дановы пошли войною на Ласем и взяли его, и поразили его мечом, и получили его в наследие, и поселились в нем, и назвали Ласем Даном по имени Дана, отца своего.
JOSH|19|48|Вот удел колена сынов Дановых, по племенам их; вот города и села их.
JOSH|19|49|Когда окончили разделение земли, по пределам ее, тогда сыны Израилевы дали среди себя удел Иисусу, сыну Навину:
JOSH|19|50|по повелению Господню дали ему город Фамнаф–Сараи, которого он просил, на горе Ефремовой; и построил он город и жил в нем.
JOSH|19|51|Вот уделы, которые Елеазар священник, Иисус, сын Навин, и начальники поколений разделили коленам сынов Израилевых, по жребию, в Силоме, пред лицем Господним, у входа скинии собрания. И кончили разделение земли.
JOSH|20|1|И сказал Господь Иисусу, говоря:
JOSH|20|2|скажи сынам Израилевым: сделайте у себя города убежища, о которых Я говорил вам чрез Моисея,
JOSH|20|3|чтобы мог убегать туда убийца, убивший человека по ошибке, без умысла; пусть [города сии] будут у вас убежищем от мстящего за кровь.
JOSH|20|4|И кто убежит в один из городов сих, пусть станет у ворот города и расскажет вслух старейшин города сего дело свое; и они примут его к себе в город и дадут ему место, чтоб он жил у них;
JOSH|20|5|и когда погонится за ним мстящий за кровь, то они не должны выдавать в руки его убийцу, потому что он без умысла убил ближнего своего, не имел к нему ненависти ни вчера, ни третьего дня;
JOSH|20|6|пусть он живет в этом городе, доколе не предстанет пред общество на суд, доколе не умрет великий священник, который будет в те дни. А потом пусть возвратится убийца и пойдет в город свой и в дом свой, в город, из которого он убежал.
JOSH|20|7|И отделили Кедес в Галилее на горе Неффалимовой, Сихем на горе Ефремовой, и Кириаф–Арбы, иначе Хеврон, на горе Иудиной;
JOSH|20|8|за Иорданом, против Иерихона к востоку, отделили: Бецер в пустыне, на равнине, от колена Рувимова, и Рамоф в Галааде от колена Гадова, и Голан в Васане от колена Манассиина;
JOSH|20|9|сии города назначены для всех сынов Израилевых и для пришельцев, живущих у них, дабы убегал туда всякий, убивший человека по ошибке, дабы не умер он от руки мстящего за кровь, доколе не предстанет пред общество [на суд].
JOSH|21|1|Начальники поколений левитских пришли к Елеазару священнику и к Иисусу, сыну Навину, и к начальникам поколений сынов Израилевых,
JOSH|21|2|и говорили им в Силоме, в земле Ханаанской, и сказали: Господь повелел чрез Моисея дать нам города для жительства и предместья их для скота нашего.
JOSH|21|3|И дали сыны Израилевы левитам из уделов своих, по повелению Господню, сии города с предместьями их.
JOSH|21|4|Вышел жребий племенам Каафовым; и досталось по жребию сынам Аарона священника, левитам, от колена Иудина, и от колена Симеонова, и от колена Вениаминова, тринадцать городов;
JOSH|21|5|а прочим сынам Каафа от племен колен Ефремова, и от колена Данова, и от половины колена Манассиина, по жребию, [досталось] десять городов;
JOSH|21|6|сынам Гирсоновым – от племен колена Иссахарова, и от колена Асирова, и от колена Неффалимова, и от половины колена Манассиина в Васане, по жребию, [досталось] тринадцать городов;
JOSH|21|7|сынам Мерариным, по их племенам, от колена Рувимова, от колена Гадова и от колена Завулонова – двенадцать городов.
JOSH|21|8|И отдали сыны Израилевы левитам сии города с предместьями их, как повелел Господь чрез Моисея, по жребию.
JOSH|21|9|От колена сынов Иудиных, и от колена сынов Симеоновых, дали города, которые [здесь] названы по имени:
JOSH|21|10|сынам Аарона, из племен Каафовых, из сынов Левия, так как жребий их был первый,
JOSH|21|11|дали Кириаф–Арбы, отца Енакова, иначе Хеврон, на горе Иудиной, и предместья его вокруг его;
JOSH|21|12|а поле сего города и села его отдали в собственность Халеву, сыну Иефонниину.
JOSH|21|13|Итак сынам Аарона священника дали город убежища для убийцы – Хеврон и предместья его, Ливну и предместья ее,
JOSH|21|14|Иаттир и предместья его, Ештемо и предместья его,
JOSH|21|15|Холон и предместья его, Давир и предместья его,
JOSH|21|16|Аин и предместья его, Ютту и предместья ее, Беф–Шемеш и предместья его: девять городов от двух колен сих;
JOSH|21|17|а от колена Вениаминова: Гаваон и предместья его, Геву и предместья ее,
JOSH|21|18|Анафоф и предместья его, Алмон и предместья его: четыре города.
JOSH|21|19|Всех городов сынам Аароновым, священникам, [досталось] тринадцать городов с предместьями их.
JOSH|21|20|И племенам сынов Каафовых, левитов, прочим из сынов Каафовых, по жребию их, достались города от колена Ефремова;
JOSH|21|21|дали им город убежища для убийцы – Сихем и предместья его, на горе Ефремовой, Гезер и предместья его,
JOSH|21|22|Кивцаим и предместья его, Беф–Орон и предместья его: четыре города;
JOSH|21|23|от колена Данова: Елфеке и предместья его, Гиввефон и предместья его,
JOSH|21|24|Аиалон и предместья его, Гаф–Риммон и предместья его: четыре города;
JOSH|21|25|от половины колена Манассиина: Фаанах и предместья его, Гаф–Риммон и предместья его: два города.
JOSH|21|26|Всех городов с предместьями их прочим племенам сынов Каафовых [досталось] десять.
JOSH|21|27|А сынам Гирсоновым, из племен левитских [дали]: от половины колена Манассиина город убежища для убийцы – Голан в Васане и предместья его, и Беештеру и предместья ее: два города;
JOSH|21|28|от колена Иссахарова: Кишион и предместья его, Давраф и предместья его,
JOSH|21|29|Иармуф и предместья его, Ен–Ганним и предместья его: четыре города;
JOSH|21|30|от колена Асирова: Мишал и предместья его, Авдон и предместья его,
JOSH|21|31|Хелкаф и предместья его, Рехов и предместья его: четыре города;
JOSH|21|32|от колена Неффалимова город убежища для убийцы – Кедес в Галилее и предместья его, Хамоф–Дор и предместья его, Карфан и предместья его: три города.
JOSH|21|33|Всех городов сынам Гирсоновым, по племенам их, [досталось] тринадцать городов с предместьями их.
JOSH|21|34|Племенам сынов Мерариных, остальным левитам, [дали]: от колена Завулонова Иокнеам и предместья его, Карфу и предместья ее,
JOSH|21|35|Димну и предместья ее, Нагалал и предместья его: четыре города;
JOSH|21|36|от колена Рувимова Бецер и предместья его, Иааца и предместья ее,
JOSH|21|37|Кедемоф и предместья его, Мефааф и предместья его: четыре города;
JOSH|21|38|от колена Гадова: города убежища для убийцы – Рамоф в Галааде и предместья его, Маханаим и предместья его,
JOSH|21|39|Есевон и предместья его, Иазер и предместья его: всех городов четыре.
JOSH|21|40|Всех городов сынам Мерариным по племенам их, остальным племенам левитским, по жребию досталось двенадцать городов.
JOSH|21|41|Всех городов левитских среди владения сынов Израилевых [было] сорок восемь городов с предместьями их.
JOSH|21|42|При городах сих были при каждом городе предместья вокруг него: так было при всех городах сих.
JOSH|21|43|Таким образом отдал Господь Израилю всю землю, которую дать клялся отцам их, и они получили ее в наследие и поселились на ней.
JOSH|21|44|И дал им Господь покой со всех сторон, как клялся отцам их, и никто из всех врагов их не устоял против них; всех врагов их предал Господь в руки их.
JOSH|21|45|Не осталось неисполнившимся ни одно слово из всех добрых слов, которые Господь говорил дому Израилеву; все сбылось.
JOSH|22|1|Тогда Иисус призвал [колено] Рувимово, Гадово и половину колена Манассиина и сказал им:
JOSH|22|2|вы исполнили все, что повелел вам Моисей, раб Господень, и слушались слов моих во всем, что я приказывал вам;
JOSH|22|3|вы не оставляли братьев своих в продолжение многих дней до сего дня и исполнили, что надлежало исполнить по повелению Господа, Бога вашего:
JOSH|22|4|ныне Господь, Бог ваш, успокоил братьев ваших, как говорил им; итак возвратитесь и пойдите в шатры ваши, в землю вашего владения, которую дал вам Моисей, раб Господень, за Иорданом;
JOSH|22|5|только старайтесь тщательно исполнять заповеди и закон, который завещал вам Моисей, раб Господень: любить Господа Бога вашего, ходить всеми путями Его, хранить заповеди Его, прилепляться к Нему и служить Ему всем сердцем вашим и всею душею вашею.
JOSH|22|6|Потом Иисус благословил их и отпустил их, и они разошлись по шатрам своим.
JOSH|22|7|Одной половине колена Манассиина дал Моисей удел в Васане, а другой половине его дал Иисус [удел] с братьями его по эту сторону Иордана к западу. И когда отпускал их Иисус в шатры их и благословил их,
JOSH|22|8|то сказал им: с великим богатством возвращаетесь вы в шатры ваши, с великим множеством скота, с серебром, с золотом, с медью и с железом, и с великим множеством одежд; разделите же добычу, [взятую] у врагов ваших, с братьями своими.
JOSH|22|9|И возвратились, и пошли сыны Рувимовы и сыны Гадовы и половина колена Манассиина от сынов Израилевых из Силома, который в земле Ханаанской, чтоб идти в землю Галаад, в землю своего владения, которую получили во владение по повелению Господню, [данному] чрез Моисея.
JOSH|22|10|Придя в окрестности Иордана, что в земле Ханаанской, сыны Рувимовы и сыны Гадовы и половина колена Манассиина соорудили там подле Иордана жертвенник, жертвенник большой по виду.
JOSH|22|11|И услышали сыны Израилевы, что говорят: вот, сыны Рувимовы и сыны Гадовы и половина колена Манассиина соорудили жертвенник на земле Ханаанской, в окрестностях Иордана, напротив сынов Израилевых.
JOSH|22|12|Когда услышали [сие] сыны Израилевы, то собралось все общество сынов Израилевых в Силом, чтоб идти против них войною.
JOSH|22|13|Впрочем сыны Израилевы [прежде] послали к сынам Рувимовым и к сынам Гадовым и к половине колена Манассиина в землю Галаадскую Финееса, сына Елеазара, священника,
JOSH|22|14|и с ним десять начальников, по начальнику поколения от всех колен Израилевых; каждый из них был начальником поколения в тысячах Израилевых.
JOSH|22|15|И пришли они к сынам Рувимовым и к сынам Гадовым и к половине колена Манассиина в землю Галаад и говорили им и сказали:
JOSH|22|16|так говорит все общество Господне: что это за преступление сделали вы пред Богом Израилевым, отступив ныне от Господа, соорудив себе жертвенник и восстав ныне против Господа?
JOSH|22|17|Разве мало для нас беззакония Фегорова, от которого мы не очистились до сего дня и [за которое] поражено было общество Господне?
JOSH|22|18|А вы отступаете сегодня от Господа! Сегодня вы восстаете против Господа, а завтра прогневается [Господь] на все общество Израилево;
JOSH|22|19|если же земля вашего владения кажется вам нечистою, то перейдите в землю владения Господня, в которой находится скиния Господня, возьмите удел среди нас, но не восставайте против Господа и против нас не восставайте, сооружая себе жертвенник, кроме жертвенника Господа, Бога нашего;
JOSH|22|20|не [один] ли Ахан, сын Зары, сделал преступление, [взяв] из заклятого, а гнев был на все общество Израилево? не один он умер за свое беззаконие.
JOSH|22|21|Сыны Рувимовы и сыны Гадовы и половина колена Манассиина в ответ [на сие] говорили начальникам тысяч Израилевых:
JOSH|22|22|Бог богов Господь, Бог богов Господь, Он знает, и Израиль да знает! Если мы восстаем и отступаем от Господа, то да не пощадит нас [Господь] в сей день!
JOSH|22|23|Если мы соорудили жертвенник для того, чтоб отступить от Господа, и для того, чтобы приносить на нем всесожжение и приношение хлебное и чтобы совершать на нем жертвы мирные, то да взыщет Сам Господь!
JOSH|22|24|Но мы сделали сие по опасению того, чтобы в последующее время не сказали ваши сыны нашим сынам: "что вам до Господа Бога Израилева!
JOSH|22|25|Господь поставил пределом между нами и вами, сыны Рувимовы и сыны Гадовы, Иордан: нет вам части в Господе". Таким образом ваши сыны не допустили бы наших сынов чтить Господа.
JOSH|22|26|Поэтому мы сказали: соорудим себе жертвенник не для всесожжения и не для жертв,
JOSH|22|27|но чтобы он между нами и вами, между последующими родами нашими, был свидетелем, что мы можем служить Господу всесожжениями нашими и жертвами нашими и благодарениями нашими, и чтобы в последующее время не сказали ваши сыны сынам нашим: "нет вам части в Господе".
JOSH|22|28|Мы говорили: если скажут так нам и родам нашим в последующее время, то мы скажем: видите подобие жертвенника Господа, которое сделали отцы наши не для всесожжения и не для жертвы, но чтобы это было свидетелем между нами и вами.
JOSH|22|29|Да не будет этого, чтобы восстать нам против Господа и отступить ныне от Господа, и соорудить жертвенник для всесожжения и для приношения хлебного и для жертв, кроме жертвенника Господа Бога нашего, который пред скиниею Его.
JOSH|22|30|Финеес священник, начальники общества и головы тысяч Израилевых, которые были с ним, услышав слова, которые говорили сыны Рувимовы и сыны Гадовы и сыны Манассиины, одобрили их.
JOSH|22|31|И сказал Финеес, сын Елеазара, священник, сынам Рувимовым и сынам Гадовым и сынам Манассииным: сегодня мы узнали, что Господь среди нас, что вы не сделали пред Господом преступления сего; теперь вы избавили сынов Израиля от руки Господней.
JOSH|22|32|И возвратился Финеес, сын Елеазара, священник, и начальники от сынов Рувимовых и от сынов Гадовых в землю Ханаанскую к сынам Израилевым и принесли им ответ.
JOSH|22|33|И сыны Израилевы одобрили это, и благословили сыны Израилевы Бога и отложили идти против них войною, чтобы разорить землю, на которой жили сыны Рувимовы и сыны Гадовы.
JOSH|22|34|И назвали сыны Рувимовы и сыны Гадовы жертвенник: [Ед], потому что, [сказали они,] он свидетель между нами, что Господь есть Бог наш.
JOSH|23|1|Спустя много времени после того, как Господь успокоил Израиля от всех врагов его со всех сторон, Иисус состарился, вошел в [преклонные] лета.
JOSH|23|2|И призвал Иисус всех [сынов] Израилевых, старейшин их, начальников их, судей их и надзирателей их, и сказал им: я состарился, вошел в [преклонные] лета.
JOSH|23|3|Вы видели все, что сделал Господь Бог ваш пред лицем вашим со всеми сими народами, ибо Господь Бог ваш Сам сражался за вас.
JOSH|23|4|Вот, я разделил вам по жребию оставшиеся народы сии в удел коленам вашим, все народы, которые я истребил, от Иордана до великого моря, на запад солнца.
JOSH|23|5|Господь Бог ваш Сам прогонит их от вас, и истребит их пред вами, дабы вы получили в наследие землю их, как говорил вам Господь Бог ваш.
JOSH|23|6|Посему во всей точности старайтесь хранить и исполнять все написанное в книге закона Моисеева, не уклоняясь от него ни направо, ни налево.
JOSH|23|7|Не сообщайтесь с сими народами, которые остались между вами, не воспоминайте имени богов их, не клянитесь [ими] и не служите им и не поклоняйтесь им,
JOSH|23|8|но прилепитесь к Господу Богу вашему, как вы делали до сего дня.
JOSH|23|9|Господь прогнал от вас народы великие и сильные, и пред вами никто не устоял до сего дня;
JOSH|23|10|один из вас прогоняет тысячу, ибо Господь Бог ваш Сам сражается за вас, как говорил вам.
JOSH|23|11|Посему всячески старайтесь любить Господа Бога вашего.
JOSH|23|12|Если же вы отвратитесь и пристанете к оставшимся из народов сих, которые остались между вами, и вступите в родство с ними и будете ходить к ним и они к вам,
JOSH|23|13|то знайте, что Господь Бог ваш не будет уже прогонять от вас народы сии, но они будут для вас петлею и сетью, бичом для ребр ваших и терном для глаз ваших, доколе не будете истреблены с сей доброй земли, которую дал вам Господь Бог ваш.
JOSH|23|14|Вот, я ныне отхожу в путь всей земли. А вы знаете всем сердцем вашим и всею душею вашею, что не осталось тщетным ни одно слово из всех добрых слов, которые говорил о вас Господь Бог ваш; все сбылось для вас, ни одно слово не осталось неисполнившимся.
JOSH|23|15|Но как сбылось над вами всякое доброе слово, которое говорил вам Господь Бог ваш, так Господь исполнит над вами всякое злое слово, доколе не истребит вас с этой доброй земли, которую дал вам Господь Бог ваш.
JOSH|23|16|Если вы преступите завет Господа Бога вашего, который Он поставил с вами, и пойдете и будете служить другим богам и поклоняться им, то возгорится на вас гнев Господень, и скоро сгибнете с этой доброй земли, которую дал вам [Господь].
JOSH|24|1|И собрал Иисус все колена Израилевы в Сихем и призвал старейшин Израиля и начальников его, и судей его и надзирателей его, и предстали пред [Господа] Бога.
JOSH|24|2|И сказал Иисус всему народу: так говорит Господь Бог Израилев: "за рекою жили отцы ваши издревле, Фарра, отец Авраама и отец Нахора, и служили иным богам.
JOSH|24|3|Но Я взял отца вашего Авраама из–за реки и водил его по всей земле Ханаанской, и размножил семя его и дал ему Исаака.
JOSH|24|4|Исааку дал Иакова и Исава. Исаву дал Я гору Сеир в наследие; Иаков же и сыны его перешли в Египет
JOSH|24|5|И послал Я Моисея и Аарона и поразил Египет язвами, которые делал Я среди его, и потом вывел вас.
JOSH|24|6|Я вывел отцов ваших из Египта, и вы пришли к [Чермному] морю. Тогда Египтяне гнались за отцами вашими с колесницами и всадниками до Чермного моря;
JOSH|24|7|но они возопили к Господу, и Он положил тьму между вами и Египтянами и навел на них море, которое их и покрыло. Глаза ваши видели, что Я сделал в Египте. [Потом] много времени пробыли вы в пустыне.
JOSH|24|8|И привел Я вас к земле Аморреев, живших за Иорданом; они сразились с вами, но Я предал их в руки ваши, и вы получили в наследие землю их, и Я истребил их пред вами.
JOSH|24|9|Восстал Валак, сын Сепфоров, царь Моавитский, и пошел войною на Израиля, и послал и призвал Валаама, сына Веорова, чтоб он проклял вас;
JOSH|24|10|но Я не хотел послушать Валаама, – и он благословил вас, и Я избавил вас из рук его.
JOSH|24|11|Вы перешли Иордан и пришли к Иерихону. И стали воевать с вами жители Иерихона, Аморреи, и Ферезеи, и Хананеи, и Хеттеи, и Гергесеи, и Евеи, и Иевусеи, но Я предал их в руки ваши.
JOSH|24|12|Я послал пред вами шершней, которые прогнали их от вас, двух царей Аморрейских; не мечом твоим и не луком твоим [сделано это].
JOSH|24|13|И дал Я вам землю, над которою ты не трудился, и города, которых вы не строили, и вы живете в них; из виноградных и масличных садов, которых вы не насаждали, вы едите [плоды]".
JOSH|24|14|Итак бойтесь Господа и служите Ему в чистоте и искренности; отвергните богов, которым служили отцы ваши за рекою и в Египте, а служите Господу.
JOSH|24|15|Если же не угодно вам служить Господу, то изберите себе ныне, кому служить, богам ли, которым служили отцы ваши, бывшие за рекою, или богам Аморреев, в земле которых живете; а я и дом мой будем служить Господу.
JOSH|24|16|И отвечал народ и сказал: нет, не будет того, чтобы мы оставили Господа и стали служить другим богам!
JOSH|24|17|Ибо Господь – Бог наш, Он вывел нас и отцов наших из земли Египетской, из дома рабства, и делал пред глазами нашими великие знамения и хранил нас на всем пути, по которому мы шли, и среди всех народов, чрез которые мы проходили.
JOSH|24|18|Господь прогнал от нас все народы и Аморреев, живших в сей земле. Посему и мы будем служить Господу, ибо Он – Бог наш.
JOSH|24|19|Иисус сказал народу: не возможете служить Господу, ибо Он Бог святый, Бог ревнитель, не потерпит беззакония вашего и грехов ваших.
JOSH|24|20|Если вы оставите Господа и будете служить чужим богам, то Он наведет на вас зло и истребит вас, после того как благотворил вам.
JOSH|24|21|И сказал народ Иисусу: нет, мы Господу будем служить.
JOSH|24|22|Иисус сказал народу: вы свидетели о себе, что вы избрали себе Господа – служить Ему? Они отвечали: свидетели.
JOSH|24|23|Итак отвергните чужих богов, которые у вас, и обратите сердце свое к Господу Богу Израилеву.
JOSH|24|24|Народ сказал Иисусу: Господу Богу нашему будем служить и гласа Его будем слушать.
JOSH|24|25|И заключил Иисус с народом завет в тот день и дал ему постановления и закон в Сихеме.
JOSH|24|26|И вписал Иисус слова сии в книгу закона Божия, и взял большой камень и положил его там под дубом, который подле святилища Господня.
JOSH|24|27|И сказал Иисус всему народу: вот, камень сей будет нам свидетелем, ибо он слышал все слова Господа, которые Он говорил с нами; он да будет свидетелем против вас, чтобы вы не солгали пред Богом вашим.
JOSH|24|28|И отпустил Иисус народ, каждого в свой удел.
JOSH|24|29|После сего умер Иисус, сын Навин, раб Господень, будучи ста десяти лет.
JOSH|24|30|И похоронили его в пределе его удела в Фамнаф–Сараи, что на горе Ефремовой, на север от горы Гааша.
JOSH|24|31|И служил Израиль Господу во все дни Иисуса и во все дни старейшин, которых жизнь продлилась после Иисуса и которые видели все дела Господа, какие Он сделал Израилю.
JOSH|24|32|И кости Иосифа, которые вынесли сыны Израилевы из Египта, схоронили в Сихеме, в участке поля, которое купил Иаков у сынов Еммора, отца Сихемова, за сто монет и которое досталось в удел сынам Иосифовым.
JOSH|24|33|[После сего] умер и Елеазар, сын Аарона, и похоронили его на холме Финееса, сына его, который дан ему на горе Ефремовой.
JOSH|24|34|[В тот день сыны Израилевы, взяв ковчег Божий, носили с собою, и Финеес был священником вместо Елеазара, отца своего, доколе не умер и не был погребен в [городе] своем Гаваофе.
JOSH|24|35|И сыны Израилевы пошли каждый в свое место и в свой город.
JOSH|24|36|И стали сыны Израилевы служить Астарте и Астарофу и богам окрестных народов; и предал их Господь в руки Еглона, царя Моавитского, и он владел ими восемнадцать лет.
