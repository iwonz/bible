TITUS|1|1|Павел, раб Божий, Апостол же Иисуса Христа, по вере избранных Божиих и познанию истины, [относящейся] к благочестию,
TITUS|1|2|в надежде вечной жизни, которую обещал неизменный в слове Бог прежде вековых времен,
TITUS|1|3|а в свое время явил Свое слово в проповеди, вверенной мне по повелению Спасителя нашего, Бога, –
TITUS|1|4|Титу, истинному сыну по общей вере: благодать, милость и мир от Бога Отца и Господа Иисуса Христа, Спасителя нашего.
TITUS|1|5|Для того я оставил тебя в Крите, чтобы ты довершил недоконченное и поставил по всем городам пресвитеров, как я тебе приказывал:
TITUS|1|6|если кто непорочен, муж одной жены, детей имеет верных, не укоряемых в распутстве или непокорности.
TITUS|1|7|Ибо епископ должен быть непорочен, как Божий домостроитель, не дерзок, не гневлив, не пьяница, не бийца, не корыстолюбец,
TITUS|1|8|но страннолюбив, любящий добро, целомудрен, справедлив, благочестив, воздержан,
TITUS|1|9|держащийся истинного слова, согласного с учением, чтобы он был силен и наставлять в здравом учении и противящихся обличать.
TITUS|1|10|Ибо есть много и непокорных, пустословов и обманщиков, особенно из обрезанных,
TITUS|1|11|каковым должно заграждать уста: они развращают целые домы, уча, чему не должно, из постыдной корысти.
TITUS|1|12|Из них же самих один стихотворец сказал: "Критяне всегда лжецы, злые звери, утробы ленивые".
TITUS|1|13|Свидетельство это справедливо. По сей причине обличай их строго, дабы они были здравы в вере,
TITUS|1|14|не внимая Иудейским басням и постановлениям людей, отвращающихся от истины.
TITUS|1|15|Для чистых все чисто; а для оскверненных и неверных нет ничего чистого, но осквернены и ум их и совесть.
TITUS|1|16|Они говорят, что знают Бога, а делами отрекаются, будучи гнусны и непокорны и не способны ни к какому доброму делу.
TITUS|2|1|Ты же говори то, что сообразно с здравым учением:
TITUS|2|2|чтобы старцы были бдительны, степенны, целомудренны, здравы в вере, в любви, в терпении;
TITUS|2|3|чтобы старицы также одевались прилично святым, не были клеветницы, не порабощались пьянству, учили добру;
TITUS|2|4|чтобы вразумляли молодых любить мужей, любить детей,
TITUS|2|5|быть целомудренными, чистыми, попечительными о доме, добрыми, покорными своим мужьям, да не порицается слово Божие.
TITUS|2|6|Юношей также увещевай быть целомудренными.
TITUS|2|7|Во всем показывай в себе образец добрых дел, в учительстве чистоту, степенность, неповрежденность,
TITUS|2|8|слово здравое, неукоризненное, чтобы противник был посрамлен, не имея ничего сказать о нас худого.
TITUS|2|9|Рабов [увещевай] повиноваться своим господам, угождать им во всем, не прекословить,
TITUS|2|10|не красть, но оказывать всю добрую верность, дабы они во всем были украшением учению Спасителя нашего, Бога.
TITUS|2|11|Ибо явилась благодать Божия, спасительная для всех человеков,
TITUS|2|12|научающая нас, чтобы мы, отвергнув нечестие и мирские похоти, целомудренно, праведно и благочестиво жили в нынешнем веке,
TITUS|2|13|ожидая блаженного упования и явления славы великого Бога и Спасителя нашего Иисуса Христа,
TITUS|2|14|Который дал Себя за нас, чтобы избавить нас от всякого беззакония и очистить Себе народ особенный, ревностный к добрым делам.
TITUS|2|15|Сие говори, увещевай и обличай со всякою властью, чтобы никто не пренебрегал тебя.
TITUS|3|1|Напоминай им повиноваться и покоряться начальству и властям, быть готовыми на всякое доброе дело,
TITUS|3|2|никого не злословить, быть не сварливыми, но тихими, и оказывать всякую кротость ко всем человекам.
TITUS|3|3|Ибо и мы были некогда несмысленны, непокорны, заблуждшие, были рабы похотей и различных удовольствий, жили в злобе и зависти, были гнусны, ненавидели друг друга.
TITUS|3|4|Когда же явилась благодать и человеколюбие Спасителя нашего, Бога,
TITUS|3|5|Он спас нас не по делам праведности, которые бы мы сотворили, а по Своей милости, банею возрождения и обновления Святым Духом,
TITUS|3|6|Которого излил на нас обильно через Иисуса Христа, Спасителя нашего,
TITUS|3|7|чтобы, оправдавшись Его благодатью, мы по упованию соделались наследниками вечной жизни.
TITUS|3|8|Слово это верно; и я желаю, чтобы ты подтверждал о сем, дабы уверовавшие в Бога старались быть прилежными к добрым делам: это хорошо и полезно человекам.
TITUS|3|9|Глупых же состязаний и родословий, и споров и распрей о законе удаляйся, ибо они бесполезны и суетны.
TITUS|3|10|Еретика, после первого и второго вразумления, отвращайся,
TITUS|3|11|зная, что таковой развратился и грешит, будучи самоосужден.
TITUS|3|12|Когда пришлю к тебе Артему или Тихика, поспеши придти ко мне в Никополь, ибо я положил там провести зиму.
TITUS|3|13|Зину законника и Аполлоса позаботься отправить так, чтобы у них ни в чем не было недостатка.
TITUS|3|14|Пусть и наши учатся упражняться в добрых делах, [в] [удовлетворении] необходимым нуждам, дабы не были бесплодны.
TITUS|3|15|Приветствуют тебя все находящиеся со мною. Приветствуй любящих нас в вере. Благодать со всеми вами. Аминь.
