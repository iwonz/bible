JOSH|1|1|Now after the death of Moses the servant of the LORD it came to pass, that the LORD spake unto Joshua the son of Nun, Moses' minister, saying,
JOSH|1|2|Moses my servant is dead; now therefore arise, go over this Jordan, thou, and all this people, unto the land which I do give to them, even to the children of Israel.
JOSH|1|3|Every place that the sole of your foot shall tread upon, that have I given unto you, as I said unto Moses.
JOSH|1|4|From the wilderness and this Lebanon even unto the great river, the river Euphrates, all the land of the Hittites, and unto the great sea toward the going down of the sun, shall be your coast.
JOSH|1|5|There shall not any man be able to stand before thee all the days of thy life: as I was with Moses, so I will be with thee: I will not fail thee, nor forsake thee.
JOSH|1|6|Be strong and of a good courage: for unto this people shalt thou divide for an inheritance the land, which I sware unto their fathers to give them.
JOSH|1|7|Only be thou strong and very courageous, that thou mayest observe to do according to all the law, which Moses my servant commanded thee: turn not from it to the right hand or to the left, that thou mayest prosper whithersoever thou goest.
JOSH|1|8|This book of the law shall not depart out of thy mouth; but thou shalt meditate therein day and night, that thou mayest observe to do according to all that is written therein: for then thou shalt make thy way prosperous, and then thou shalt have good success.
JOSH|1|9|Have not I commanded thee? Be strong and of a good courage; be not afraid, neither be thou dismayed: for the LORD thy God is with thee whithersoever thou goest.
JOSH|1|10|Then Joshua commanded the officers of the people, saying,
JOSH|1|11|Pass through the host, and command the people, saying, Prepare you victuals; for within three days ye shall pass over this Jordan, to go in to possess the land, which the LORD your God giveth you to possess it.
JOSH|1|12|And to the Reubenites, and to the Gadites, and to half the tribe of Manasseh, spake Joshua, saying,
JOSH|1|13|Remember the word which Moses the servant of the LORD commanded you, saying, The LORD your God hath given you rest, and hath given you this land.
JOSH|1|14|Your wives, your little ones, and your cattle, shall remain in the land which Moses gave you on this side Jordan; but ye shall pass before your brethren armed, all the mighty men of valor, and help them;
JOSH|1|15|Until the LORD have given your brethren rest, as he hath given you, and they also have possessed the land which the LORD your God giveth them: then ye shall return unto the land of your possession, and enjoy it, which Moses the LORD's servant gave you on this side Jordan toward the sunrising.
JOSH|1|16|And they answered Joshua, saying, All that thou commandest us we will do, and whithersoever thou sendest us, we will go.
JOSH|1|17|According as we hearkened unto Moses in all things, so will we hearken unto thee: only the LORD thy God be with thee, as he was with Moses.
JOSH|1|18|Whosoever he be that doth rebel against thy commandment, and will not hearken unto thy words in all that thou commandest him, he shall be put to death: only be strong and of a good courage.
JOSH|2|1|And Joshua the son of Nun sent out of Shittim two men to spy secretly, saying, Go view the land, even Jericho. And they went, and came into an harlot's house, named Rahab, and lodged there.
JOSH|2|2|And it was told the king of Jericho, saying, Behold, there came men in hither to night of the children of Israel to search out the country.
JOSH|2|3|And the king of Jericho sent unto Rahab, saying, Bring forth the men that are come to thee, which are entered into thine house: for they be come to search out all the country.
JOSH|2|4|And the woman took the two men, and hid them, and said thus, There came men unto me, but I wist not whence they were:
JOSH|2|5|And it came to pass about the time of shutting of the gate, when it was dark, that the men went out: whither the men went I wot not: pursue after them quickly; for ye shall overtake them.
JOSH|2|6|But she had brought them up to the roof of the house, and hid them with the stalks of flax, which she had laid in order upon the roof.
JOSH|2|7|And the men pursued after them the way to Jordan unto the fords: and as soon as they which pursued after them were gone out, they shut the gate.
JOSH|2|8|And before they were laid down, she came up unto them upon the roof;
JOSH|2|9|And she said unto the men, I know that the LORD hath given you the land, and that your terror is fallen upon us, and that all the inhabitants of the land faint because of you.
JOSH|2|10|For we have heard how the LORD dried up the water of the Red sea for you, when ye came out of Egypt; and what ye did unto the two kings of the Amorites, that were on the other side Jordan, Sihon and Og, whom ye utterly destroyed.
JOSH|2|11|And as soon as we had heard these things, our hearts did melt, neither did there remain any more courage in any man, because of you: for the LORD your God, he is God in heaven above, and in earth beneath.
JOSH|2|12|Now therefore, I pray you, swear unto me by the LORD, since I have showed you kindness, that ye will also show kindness unto my father's house, and give me a true token:
JOSH|2|13|And that ye will save alive my father, and my mother, and my brethren, and my sisters, and all that they have, and deliver our lives from death.
JOSH|2|14|And the men answered her, Our life for yours, if ye utter not this our business. And it shall be, when the LORD hath given us the land, that we will deal kindly and truly with thee.
JOSH|2|15|Then she let them down by a cord through the window: for her house was upon the town wall, and she dwelt upon the wall.
JOSH|2|16|And she said unto them, Get you to the mountain, lest the pursuers meet you; and hide yourselves there three days, until the pursuers be returned: and afterward may ye go your way.
JOSH|2|17|And the men said unto her, We will be blameless of this thine oath which thou hast made us swear.
JOSH|2|18|Behold, when we come into the land, thou shalt bind this line of scarlet thread in the window which thou didst let us down by: and thou shalt bring thy father, and thy mother, and thy brethren, and all thy father's household, home unto thee.
JOSH|2|19|And it shall be, that whosoever shall go out of the doors of thy house into the street, his blood shall be upon his head, and we will be guiltless: and whosoever shall be with thee in the house, his blood shall be on our head, if any hand be upon him.
JOSH|2|20|And if thou utter this our business, then we will be quit of thine oath which thou hast made us to swear.
JOSH|2|21|And she said, According unto your words, so be it. And she sent them away, and they departed: and she bound the scarlet line in the window.
JOSH|2|22|And they went, and came unto the mountain, and abode there three days, until the pursuers were returned: and the pursuers sought them throughout all the way, but found them not.
JOSH|2|23|So the two men returned, and descended from the mountain, and passed over, and came to Joshua the son of Nun, and told him all things that befell them:
JOSH|2|24|And they said unto Joshua, Truly the LORD hath delivered into our hands all the land; for even all the inhabitants of the country do faint because of us.
JOSH|3|1|And Joshua rose early in the morning; and they removed from Shittim, and came to Jordan, he and all the children of Israel, and lodged there before they passed over.
JOSH|3|2|And it came to pass after three days, that the officers went through the host;
JOSH|3|3|And they commanded the people, saying, When ye see the ark of the covenant of the LORD your God, and the priests the Levites bearing it, then ye shall remove from your place, and go after it.
JOSH|3|4|Yet there shall be a space between you and it, about two thousand cubits by measure: come not near unto it, that ye may know the way by which ye must go: for ye have not passed this way heretofore.
JOSH|3|5|And Joshua said unto the people, Sanctify yourselves: for to morrow the LORD will do wonders among you.
JOSH|3|6|And Joshua spake unto the priests, saying, Take up the ark of the covenant, and pass over before the people. And they took up the ark of the covenant, and went before the people.
JOSH|3|7|And the LORD said unto Joshua, This day will I begin to magnify thee in the sight of all Israel, that they may know that, as I was with Moses, so I will be with thee.
JOSH|3|8|And thou shalt command the priests that bear the ark of the covenant, saying, When ye are come to the brink of the water of Jordan, ye shall stand still in Jordan.
JOSH|3|9|And Joshua said unto the children of Israel, Come hither, and hear the words of the LORD your God.
JOSH|3|10|And Joshua said, Hereby ye shall know that the living God is among you, and that he will without fail drive out from before you the Canaanites, and the Hittites, and the Hivites, and the Perizzites, and the Girgashites, and the Amorites, and the Jebusites.
JOSH|3|11|Behold, the ark of the covenant of the LORD of all the earth passeth over before you into Jordan.
JOSH|3|12|Now therefore take you twelve men out of the tribes of Israel, out of every tribe a man.
JOSH|3|13|And it shall come to pass, as soon as the soles of the feet of the priests that bear the ark of the LORD, the LORD of all the earth, shall rest in the waters of Jordan, that the waters of Jordan shall be cut off from the waters that come down from above; and they shall stand upon an heap.
JOSH|3|14|And it came to pass, when the people removed from their tents, to pass over Jordan, and the priests bearing the ark of the covenant before the people;
JOSH|3|15|And as they that bare the ark were come unto Jordan, and the feet of the priests that bare the ark were dipped in the brim of the water, (for Jordan overfloweth all his banks all the time of harvest,)
JOSH|3|16|That the waters which came down from above stood and rose up upon an heap very far from the city Adam, that is beside Zaretan: and those that came down toward the sea of the plain, even the salt sea, failed, and were cut off: and the people passed over right against Jericho.
JOSH|3|17|And the priests that bare the ark of the covenant of the LORD stood firm on dry ground in the midst of Jordan, and all the Israelites passed over on dry ground, until all the people were passed clean over Jordan.
JOSH|4|1|And it came to pass, when all the people were clean passed over Jordan, that the LORD spake unto Joshua, saying,
JOSH|4|2|Take you twelve men out of the people, out of every tribe a man,
JOSH|4|3|And command ye them, saying, Take you hence out of the midst of Jordan, out of the place where the priests' feet stood firm, twelve stones, and ye shall carry them over with you, and leave them in the lodging place, where ye shall lodge this night.
JOSH|4|4|Then Joshua called the twelve men, whom he had prepared of the children of Israel, out of every tribe a man:
JOSH|4|5|And Joshua said unto them, Pass over before the ark of the LORD your God into the midst of Jordan, and take you up every man of you a stone upon his shoulder, according unto the number of the tribes of the children of Israel:
JOSH|4|6|That this may be a sign among you, that when your children ask their fathers in time to come, saying, What mean ye by these stones?
JOSH|4|7|Then ye shall answer them, That the waters of Jordan were cut off before the ark of the covenant of the LORD; when it passed over Jordan, the waters of Jordan were cut off: and these stones shall be for a memorial unto the children of Israel for ever.
JOSH|4|8|And the children of Israel did so as Joshua commanded, and took up twelve stones out of the midst of Jordan, as the LORD spake unto Joshua, according to the number of the tribes of the children of Israel, and carried them over with them unto the place where they lodged, and laid them down there.
JOSH|4|9|And Joshua set up twelve stones in the midst of Jordan, in the place where the feet of the priests which bare the ark of the covenant stood: and they are there unto this day.
JOSH|4|10|For the priests which bare the ark stood in the midst of Jordan, until everything was finished that the LORD commanded Joshua to speak unto the people, according to all that Moses commanded Joshua: and the people hasted and passed over.
JOSH|4|11|And it came to pass, when all the people were clean passed over, that the ark of the LORD passed over, and the priests, in the presence of the people.
JOSH|4|12|And the children of Reuben, and the children of Gad, and half the tribe of Manasseh, passed over armed before the children of Israel, as Moses spake unto them:
JOSH|4|13|About forty thousand prepared for war passed over before the LORD unto battle, to the plains of Jericho.
JOSH|4|14|On that day the LORD magnified Joshua in the sight of all Israel; and they feared him, as they feared Moses, all the days of his life.
JOSH|4|15|And the LORD spake unto Joshua, saying,
JOSH|4|16|Command the priests that bear the ark of the testimony, that they come up out of Jordan.
JOSH|4|17|Joshua therefore commanded the priests, saying, Come ye up out of Jordan.
JOSH|4|18|And it came to pass, when the priests that bare the ark of the covenant of the LORD were come up out of the midst of Jordan, and the soles of the priests' feet were lifted up unto the dry land, that the waters of Jordan returned unto their place, and flowed over all his banks, as they did before.
JOSH|4|19|And the people came up out of Jordan on the tenth day of the first month, and encamped in Gilgal, in the east border of Jericho.
JOSH|4|20|And those twelve stones, which they took out of Jordan, did Joshua pitch in Gilgal.
JOSH|4|21|And he spake unto the children of Israel, saying, When your children shall ask their fathers in time to come, saying, What mean these stones?
JOSH|4|22|Then ye shall let your children know, saying, Israel came over this Jordan on dry land.
JOSH|4|23|For the LORD your God dried up the waters of Jordan from before you, until ye were passed over, as the LORD your God did to the Red sea, which he dried up from before us, until we were gone over:
JOSH|4|24|That all the people of the earth might know the hand of the LORD, that it is mighty: that ye might fear the LORD your God for ever.
JOSH|5|1|And it came to pass, when all the kings of the Amorites, which were on the side of Jordan westward, and all the kings of the Canaanites, which were by the sea, heard that the LORD had dried up the waters of Jordan from before the children of Israel, until we were passed over, that their heart melted, neither was there spirit in them any more, because of the children of Israel.
JOSH|5|2|At that time the LORD said unto Joshua, Make thee sharp knives, and circumcise again the children of Israel the second time.
JOSH|5|3|And Joshua made him sharp knives, and circumcised the children of Israel at the hill of the foreskins.
JOSH|5|4|And this is the cause why Joshua did circumcise: All the people that came out of Egypt, that were males, even all the men of war, died in the wilderness by the way, after they came out of Egypt.
JOSH|5|5|Now all the people that came out were circumcised: but all the people that were born in the wilderness by the way as they came forth out of Egypt, them they had not circumcised.
JOSH|5|6|For the children of Israel walked forty years in the wilderness, till all the people that were men of war, which came out of Egypt, were consumed, because they obeyed not the voice of the LORD: unto whom the LORD sware that he would not show them the land, which the LORD sware unto their fathers that he would give us, a land that floweth with milk and honey.
JOSH|5|7|And their children, whom he raised up in their stead, them Joshua circumcised: for they were uncircumcised, because they had not circumcised them by the way.
JOSH|5|8|And it came to pass, when they had done circumcising all the people, that they abode in their places in the camp, till they were whole.
JOSH|5|9|And the LORD said unto Joshua, This day have I rolled away the reproach of Egypt from off you. Wherefore the name of the place is called Gilgal unto this day.
JOSH|5|10|And the children of Israel encamped in Gilgal, and kept the passover on the fourteenth day of the month at even in the plains of Jericho.
JOSH|5|11|And they did eat of the old corn of the land on the morrow after the passover, unleavened cakes, and parched corn in the selfsame day.
JOSH|5|12|And the manna ceased on the morrow after they had eaten of the old corn of the land; neither had the children of Israel manna any more; but they did eat of the fruit of the land of Canaan that year.
JOSH|5|13|And it came to pass, when Joshua was by Jericho, that he lifted up his eyes and looked, and, behold, there stood a man over against him with his sword drawn in his hand: and Joshua went unto him, and said unto him, Art thou for us, or for our adversaries?
JOSH|5|14|And he said, Nay; but as captain of the host of the LORD am I now come. And Joshua fell on his face to the earth, and did worship, and said unto him, What saith my Lord unto his servant?
JOSH|5|15|And the captain of the LORD's host said unto Joshua, Loose thy shoe from off thy foot; for the place whereon thou standest is holy. And Joshua did so.
JOSH|6|1|Now Jericho was straitly shut up because of the children of Israel: none went out, and none came in.
JOSH|6|2|And the LORD said unto Joshua, See, I have given into thine hand Jericho, and the king thereof, and the mighty men of valor.
JOSH|6|3|And ye shall compass the city, all ye men of war, and go round about the city once. Thus shalt thou do six days.
JOSH|6|4|And seven priests shall bear before the ark seven trumpets of rams' horns: and the seventh day ye shall compass the city seven times, and the priests shall blow with the trumpets.
JOSH|6|5|And it shall come to pass, that when they make a long blast with the ram's horn, and when ye hear the sound of the trumpet, all the people shall shout with a great shout; and the wall of the city shall fall down flat, and the people shall ascend up every man straight before him.
JOSH|6|6|And Joshua the son of Nun called the priests, and said unto them, Take up the ark of the covenant, and let seven priests bear seven trumpets of rams' horns before the ark of the LORD.
JOSH|6|7|And he said unto the people, Pass on, and compass the city, and let him that is armed pass on before the ark of the LORD.
JOSH|6|8|And it came to pass, when Joshua had spoken unto the people, that the seven priests bearing the seven trumpets of rams' horns passed on before the LORD, and blew with the trumpets: and the ark of the covenant of the LORD followed them.
JOSH|6|9|And the armed men went before the priests that blew with the trumpets, and the rearward came after the ark, the priests going on, and blowing with the trumpets.
JOSH|6|10|And Joshua had commanded the people, saying, Ye shall not shout, nor make any noise with your voice, neither shall any word proceed out of your mouth, until the day I bid you shout; then shall ye shout.
JOSH|6|11|So the ark of the LORD compassed the city, going about it once: and they came into the camp, and lodged in the camp.
JOSH|6|12|And Joshua rose early in the morning, and the priests took up the ark of the LORD.
JOSH|6|13|And seven priests bearing seven trumpets of rams' horns before the ark of the LORD went on continually, and blew with the trumpets: and the armed men went before them; but the rearward came after the ark of the LORD, the priests going on, and blowing with the trumpets.
JOSH|6|14|And the second day they compassed the city once, and returned into the camp: so they did six days.
JOSH|6|15|And it came to pass on the seventh day, that they rose early about the dawning of the day, and compassed the city after the same manner seven times: only on that day they compassed the city seven times.
JOSH|6|16|And it came to pass at the seventh time, when the priests blew with the trumpets, Joshua said unto the people, Shout; for the LORD hath given you the city.
JOSH|6|17|And the city shall be accursed, even it, and all that are therein, to the LORD: only Rahab the harlot shall live, she and all that are with her in the house, because she hid the messengers that we sent.
JOSH|6|18|And ye, in any wise keep yourselves from the accursed thing, lest ye make yourselves accursed, when ye take of the accursed thing, and make the camp of Israel a curse, and trouble it.
JOSH|6|19|But all the silver, and gold, and vessels of brass and iron, are consecrated unto the LORD: they shall come into the treasury of the LORD.
JOSH|6|20|So the people shouted when the priests blew with the trumpets: and it came to pass, when the people heard the sound of the trumpet, and the people shouted with a great shout, that the wall fell down flat, so that the people went up into the city, every man straight before him, and they took the city.
JOSH|6|21|And they utterly destroyed all that was in the city, both man and woman, young and old, and ox, and sheep, and ass, with the edge of the sword.
JOSH|6|22|But Joshua had said unto the two men that had spied out the country, Go into the harlot's house, and bring out thence the woman, and all that she hath, as ye sware unto her.
JOSH|6|23|And the young men that were spies went in, and brought out Rahab, and her father, and her mother, and her brethren, and all that she had; and they brought out all her kindred, and left them without the camp of Israel.
JOSH|6|24|And they burnt the city with fire, and all that was therein: only the silver, and the gold, and the vessels of brass and of iron, they put into the treasury of the house of the LORD.
JOSH|6|25|And Joshua saved Rahab the harlot alive, and her father's household, and all that she had; and she dwelleth in Israel even unto this day; because she hid the messengers, which Joshua sent to spy out Jericho.
JOSH|6|26|And Joshua adjured them at that time, saying, Cursed be the man before the LORD, that riseth up and buildeth this city Jericho: he shall lay the foundation thereof in his firstborn, and in his youngest son shall he set up the gates of it.
JOSH|6|27|So the LORD was with Joshua; and his fame was noised throughout all the country.
JOSH|7|1|But the children of Israel committed a trespass in the accursed thing: for Achan, the son of Carmi, the son of Zabdi, the son of Zerah, of the tribe of Judah, took of the accursed thing: and the anger of the LORD was kindled against the children of Israel.
JOSH|7|2|And Joshua sent men from Jericho to Ai, which is beside Bethaven, on the east of Bethel, and spake unto them, saying, Go up and view the country. And the men went up and viewed Ai.
JOSH|7|3|And they returned to Joshua, and said unto him, Let not all the people go up; but let about two or three thousand men go up and smite Ai; and make not all the people to labor thither; for they are but few.
JOSH|7|4|So there went up thither of the people about three thousand men: and they fled before the men of Ai.
JOSH|7|5|And the men of Ai smote of them about thirty and six men: for they chased them from before the gate even unto Shebarim, and smote them in the going down: wherefore the hearts of the people melted, and became as water.
JOSH|7|6|And Joshua rent his clothes, and fell to the earth upon his face before the ark of the LORD until the eventide, he and the elders of Israel, and put dust upon their heads.
JOSH|7|7|And Joshua said, Alas, O LORD God, wherefore hast thou at all brought this people over Jordan, to deliver us into the hand of the Amorites, to destroy us? would to God we had been content, and dwelt on the other side Jordan!
JOSH|7|8|O LORD, what shall I say, when Israel turneth their backs before their enemies!
JOSH|7|9|For the Canaanites and all the inhabitants of the land shall hear of it, and shall environ us round, and cut off our name from the earth: and what wilt thou do unto thy great name?
JOSH|7|10|And the LORD said unto Joshua, Get thee up; wherefore liest thou thus upon thy face?
JOSH|7|11|Israel hath sinned, and they have also transgressed my covenant which I commanded them: for they have even taken of the accursed thing, and have also stolen, and dissembled also, and they have put it even among their own stuff.
JOSH|7|12|Therefore the children of Israel could not stand before their enemies, but turned their backs before their enemies, because they were accursed: neither will I be with you any more, except ye destroy the accursed from among you.
JOSH|7|13|Up, sanctify the people, and say, Sanctify yourselves against to morrow: for thus saith the LORD God of Israel, There is an accursed thing in the midst of thee, O Israel: thou canst not stand before thine enemies, until ye take away the accursed thing from among you.
JOSH|7|14|In the morning therefore ye shall be brought according to your tribes: and it shall be, that the tribe which the LORD taketh shall come according to the families thereof; and the family which the LORD shall take shall come by households; and the household which the LORD shall take shall come man by man.
JOSH|7|15|And it shall be, that he that is taken with the accursed thing shall be burnt with fire, he and all that he hath: because he hath transgressed the covenant of the LORD, and because he hath wrought folly in Israel.
JOSH|7|16|So Joshua rose up early in the morning, and brought Israel by their tribes; and the tribe of Judah was taken:
JOSH|7|17|And he brought the family of Judah; and he took the family of the Zarhites: and he brought the family of the Zarhites man by man; and Zabdi was taken:
JOSH|7|18|And he brought his household man by man; and Achan, the son of Carmi, the son of Zabdi, the son of Zerah, of the tribe of Judah, was taken.
JOSH|7|19|And Joshua said unto Achan, My son, give, I pray thee, glory to the LORD God of Israel, and make confession unto him; and tell me now what thou hast done; hide it not from me.
JOSH|7|20|And Achan answered Joshua, and said, Indeed I have sinned against the LORD God of Israel, and thus and thus have I done:
JOSH|7|21|When I saw among the spoils a goodly Babylonish garment, and two hundred shekels of silver, and a wedge of gold of fifty shekels weight, then I coveted them, and took them; and, behold, they are hid in the earth in the midst of my tent, and the silver under it.
JOSH|7|22|So Joshua sent messengers, and they ran unto the tent; and, behold, it was hid in his tent, and the silver under it.
JOSH|7|23|And they took them out of the midst of the tent, and brought them unto Joshua, and unto all the children of Israel, and laid them out before the LORD.
JOSH|7|24|And Joshua, and all Israel with him, took Achan the son of Zerah, and the silver, and the garment, and the wedge of gold, and his sons, and his daughters, and his oxen, and his asses, and his sheep, and his tent, and all that he had: and they brought them unto the valley of Achor.
JOSH|7|25|And Joshua said, Why hast thou troubled us? the LORD shall trouble thee this day. And all Israel stoned him with stones, and burned them with fire, after they had stoned them with stones.
JOSH|7|26|And they raised over him a great heap of stones unto this day. So the LORD turned from the fierceness of his anger. Wherefore the name of that place was called, The valley of Achor, unto this day.
JOSH|8|1|And the LORD said unto Joshua, Fear not, neither be thou dismayed: take all the people of war with thee, and arise, go up to Ai: see, I have given into thy hand the king of Ai, and his people, and his city, and his land:
JOSH|8|2|And thou shalt do to Ai and her king as thou didst unto Jericho and her king: only the spoil thereof, and the cattle thereof, shall ye take for a prey unto yourselves: lay thee an ambush for the city behind it.
JOSH|8|3|So Joshua arose, and all the people of war, to go up against Ai: and Joshua chose out thirty thousand mighty men of valor, and sent them away by night.
JOSH|8|4|And he commanded them, saying, Behold, ye shall lie in wait against the city, even behind the city: go not very far from the city, but be ye all ready:
JOSH|8|5|And I, and all the people that are with me, will approach unto the city: and it shall come to pass, when they come out against us, as at the first, that we will flee before them,
JOSH|8|6|(For they will come out after us) till we have drawn them from the city; for they will say, They flee before us, as at the first: therefore we will flee before them.
JOSH|8|7|Then ye shall rise up from the ambush, and seize upon the city: for the LORD your God will deliver it into your hand.
JOSH|8|8|And it shall be, when ye have taken the city, that ye shall set the city on fire: according to the commandment of the LORD shall ye do. See, I have commanded you.
JOSH|8|9|Joshua therefore sent them forth: and they went to lie in ambush, and abode between Bethel and Ai, on the west side of Ai: but Joshua lodged that night among the people.
JOSH|8|10|And Joshua rose up early in the morning, and numbered the people, and went up, he and the elders of Israel, before the people to Ai.
JOSH|8|11|And all the people, even the people of war that were with him, went up, and drew nigh, and came before the city, and pitched on the north side of Ai: now there was a valley between them and Ai.
JOSH|8|12|And he took about five thousand men, and set them to lie in ambush between Bethel and Ai, on the west side of the city.
JOSH|8|13|And when they had set the people, even all the host that was on the north of the city, and their liers in wait on the west of the city, Joshua went that night into the midst of the valley.
JOSH|8|14|And it came to pass, when the king of Ai saw it, that they hasted and rose up early, and the men of the city went out against Israel to battle, he and all his people, at a time appointed, before the plain; but he wist not that there were liers in ambush against him behind the city.
JOSH|8|15|And Joshua and all Israel made as if they were beaten before them, and fled by the way of the wilderness.
JOSH|8|16|And all the people that were in Ai were called together to pursue after them: and they pursued after Joshua, and were drawn away from the city.
JOSH|8|17|And there was not a man left in Ai or Bethel, that went not out after Israel: and they left the city open, and pursued after Israel.
JOSH|8|18|And the LORD said unto Joshua, Stretch out the spear that is in thy hand toward Ai; for I will give it into thine hand. And Joshua stretched out the spear that he had in his hand toward the city.
JOSH|8|19|And the ambush arose quickly out of their place, and they ran as soon as he had stretched out his hand: and they entered into the city, and took it, and hasted and set the city on fire.
JOSH|8|20|And when the men of Ai looked behind them, they saw, and, behold, the smoke of the city ascended up to heaven, and they had no power to flee this way or that way: and the people that fled to the wilderness turned back upon the pursuers.
JOSH|8|21|And when Joshua and all Israel saw that the ambush had taken the city, and that the smoke of the city ascended, then they turned again, and slew the men of Ai.
JOSH|8|22|And the other issued out of the city against them; so they were in the midst of Israel, some on this side, and some on that side: and they smote them, so that they let none of them remain or escape.
JOSH|8|23|And the king of Ai they took alive, and brought him to Joshua.
JOSH|8|24|And it came to pass, when Israel had made an end of slaying all the inhabitants of Ai in the field, in the wilderness wherein they chased them, and when they were all fallen on the edge of the sword, until they were consumed, that all the Israelites returned unto Ai, and smote it with the edge of the sword.
JOSH|8|25|And so it was, that all that fell that day, both of men and women, were twelve thousand, even all the men of Ai.
JOSH|8|26|For Joshua drew not his hand back, wherewith he stretched out the spear, until he had utterly destroyed all the inhabitants of Ai.
JOSH|8|27|Only the cattle and the spoil of that city Israel took for a prey unto themselves, according unto the word of the LORD which he commanded Joshua.
JOSH|8|28|And Joshua burnt Ai, and made it an heap for ever, even a desolation unto this day.
JOSH|8|29|And the king of Ai he hanged on a tree until eventide: and as soon as the sun was down, Joshua commanded that they should take his carcass down from the tree, and cast it at the entering of the gate of the city, and raise thereon a great heap of stones, that remaineth unto this day.
JOSH|8|30|Then Joshua built an altar unto the LORD God of Israel in mount Ebal,
JOSH|8|31|As Moses the servant of the LORD commanded the children of Israel, as it is written in the book of the law of Moses, an altar of whole stones, over which no man hath lift up any iron: and they offered thereon burnt offerings unto the LORD, and sacrificed peace offerings.
JOSH|8|32|And he wrote there upon the stones a copy of the law of Moses, which he wrote in the presence of the children of Israel.
JOSH|8|33|And all Israel, and their elders, and officers, and their judges, stood on this side the ark and on that side before the priests the Levites, which bare the ark of the covenant of the LORD, as well the stranger, as he that was born among them; half of them over against mount Gerizim, and half of them over against mount Ebal; as Moses the servant of the LORD had commanded before, that they should bless the people of Israel.
JOSH|8|34|And afterward he read all the words of the law, the blessings and cursings, according to all that is written in the book of the law.
JOSH|8|35|There was not a word of all that Moses commanded, which Joshua read not before all the congregation of Israel, with the women, and the little ones, and the strangers that were conversant among them.
JOSH|9|1|And it came to pass, when all the kings which were on this side Jordan, in the hills, and in the valleys, and in all the coasts of the great sea over against Lebanon, the Hittite, and the Amorite, the Canaanite, the Perizzite, the Hivite, and the Jebusite, heard thereof;
JOSH|9|2|That they gathered themselves together, to fight with Joshua and with Israel, with one accord.
JOSH|9|3|And when the inhabitants of Gibeon heard what Joshua had done unto Jericho and to Ai,
JOSH|9|4|They did work wilily, and went and made as if they had been ambassadors, and took old sacks upon their asses, and wine bottles, old, and rent, and bound up;
JOSH|9|5|And old shoes and clouted upon their feet, and old garments upon them; and all the bread of their provision was dry and mouldy.
JOSH|9|6|And they went to Joshua unto the camp at Gilgal, and said unto him, and to the men of Israel, We be come from a far country: now therefore make ye a league with us.
JOSH|9|7|And the men of Israel said unto the Hivites, Peradventure ye dwell among us; and how shall we make a league with you?
JOSH|9|8|And they said unto Joshua, We are thy servants. And Joshua said unto them, Who are ye? and from whence come ye?
JOSH|9|9|And they said unto him, From a very far country thy servants are come because of the name of the LORD thy God: for we have heard the fame of him, and all that he did in Egypt,
JOSH|9|10|And all that he did to the two kings of the Amorites, that were beyond Jordan, to Sihon king of Heshbon, and to Og king of Bashan, which was at Ashtaroth.
JOSH|9|11|Wherefore our elders and all the inhabitants of our country spake to us, saying, Take victuals with you for the journey, and go to meet them, and say unto them, We are your servants: therefore now make ye a league with us.
JOSH|9|12|This our bread we took hot for our provision out of our houses on the day we came forth to go unto you; but now, behold, it is dry, and it is mouldy:
JOSH|9|13|And these bottles of wine, which we filled, were new; and, behold, they be rent: and these our garments and our shoes are become old by reason of the very long journey.
JOSH|9|14|And the men took of their victuals, and asked not counsel at the mouth of the LORD.
JOSH|9|15|And Joshua made peace with them, and made a league with them, to let them live: and the princes of the congregation sware unto them.
JOSH|9|16|And it came to pass at the end of three days after they had made a league with them, that they heard that they were their neighbors, and that they dwelt among them.
JOSH|9|17|And the children of Israel journeyed, and came unto their cities on the third day. Now their cities were Gibeon, and Chephirah, and Beeroth, and Kirjathjearim.
JOSH|9|18|And the children of Israel smote them not, because the princes of the congregation had sworn unto them by the LORD God of Israel. And all the congregation murmured against the princes.
JOSH|9|19|But all the princes said unto all the congregation, We have sworn unto them by the LORD God of Israel: now therefore we may not touch them.
JOSH|9|20|This we will do to them; we will even let them live, lest wrath be upon us, because of the oath which we sware unto them.
JOSH|9|21|And the princes said unto them, Let them live; but let them be hewers of wood and drawers of water unto all the congregation; as the princes had promised them.
JOSH|9|22|And Joshua called for them, and he spake unto them, saying, Wherefore have ye beguiled us, saying, We are very far from you; when ye dwell among us?
JOSH|9|23|Now therefore ye are cursed, and there shall none of you be freed from being bondmen, and hewers of wood and drawers of water for the house of my God.
JOSH|9|24|And they answered Joshua, and said, Because it was certainly told thy servants, how that the LORD thy God commanded his servant Moses to give you all the land, and to destroy all the inhabitants of the land from before you, therefore we were sore afraid of our lives because of you, and have done this thing.
JOSH|9|25|And now, behold, we are in thine hand: as it seemeth good and right unto thee to do unto us, do.
JOSH|9|26|And so did he unto them, and delivered them out of the hand of the children of Israel, that they slew them not.
JOSH|9|27|And Joshua made them that day hewers of wood and drawers of water for the congregation, and for the altar of the LORD, even unto this day, in the place which he should choose.
JOSH|10|1|Now it came to pass, when Adonizedec king of Jerusalem had heard how Joshua had taken Ai, and had utterly destroyed it; as he had done to Jericho and her king, so he had done to Ai and her king; and how the inhabitants of Gibeon had made peace with Israel, and were among them;
JOSH|10|2|That they feared greatly, because Gibeon was a great city, as one of the royal cities, and because it was greater than Ai, and all the men thereof were mighty.
JOSH|10|3|Wherefore Adonizedec king of Jerusalem, sent unto Hoham king of Hebron, and unto Piram king of Jarmuth, and unto Japhia king of Lachish, and unto Debir king of Eglon, saying,
JOSH|10|4|Come up unto me, and help me, that we may smite Gibeon: for it hath made peace with Joshua and with the children of Israel.
JOSH|10|5|Therefore the five kings of the Amorites, the king of Jerusalem, the king of Hebron, the king of Jarmuth, the king of Lachish, the king of Eglon, gathered themselves together, and went up, they and all their hosts, and encamped before Gibeon, and made war against it.
JOSH|10|6|And the men of Gibeon sent unto Joshua to the camp to Gilgal, saying, Slack not thy hand from thy servants; come up to us quickly, and save us, and help us: for all the kings of the Amorites that dwell in the mountains are gathered together against us.
JOSH|10|7|So Joshua ascended from Gilgal, he, and all the people of war with him, and all the mighty men of valor.
JOSH|10|8|And the LORD said unto Joshua, Fear them not: for I have delivered them into thine hand; there shall not a man of them stand before thee.
JOSH|10|9|Joshua therefore came unto them suddenly, and went up from Gilgal all night.
JOSH|10|10|And the LORD discomfited them before Israel, and slew them with a great slaughter at Gibeon, and chased them along the way that goeth up to Bethhoron, and smote them to Azekah, and unto Makkedah.
JOSH|10|11|And it came to pass, as they fled from before Israel, and were in the going down to Bethhoron, that the LORD cast down great stones from heaven upon them unto Azekah, and they died: they were more which died with hailstones than they whom the children of Israel slew with the sword.
JOSH|10|12|Then spake Joshua to the LORD in the day when the LORD delivered up the Amorites before the children of Israel, and he said in the sight of Israel, Sun, stand thou still upon Gibeon; and thou, Moon, in the valley of Ajalon.
JOSH|10|13|And the sun stood still, and the moon stayed, until the people had avenged themselves upon their enemies. Is not this written in the book of Jasher? So the sun stood still in the midst of heaven, and hasted not to go down about a whole day.
JOSH|10|14|And there was no day like that before it or after it, that the LORD hearkened unto the voice of a man: for the LORD fought for Israel.
JOSH|10|15|And Joshua returned, and all Israel with him, unto the camp to Gilgal.
JOSH|10|16|But these five kings fled, and hid themselves in a cave at Makkedah.
JOSH|10|17|And it was told Joshua, saying, The five kings are found hid in a cave at Makkedah.
JOSH|10|18|And Joshua said, Roll great stones upon the mouth of the cave, and set men by it for to keep them:
JOSH|10|19|And stay ye not, but pursue after your enemies, and smite the hindmost of them; suffer them not to enter into their cities: for the LORD your God hath delivered them into your hand.
JOSH|10|20|And it came to pass, when Joshua and the children of Israel had made an end of slaying them with a very great slaughter, till they were consumed, that the rest which remained of them entered into fenced cities.
JOSH|10|21|And all the people returned to the camp to Joshua at Makkedah in peace: none moved his tongue against any of the children of Israel.
JOSH|10|22|Then said Joshua, Open the mouth of the cave, and bring out those five kings unto me out of the cave.
JOSH|10|23|And they did so, and brought forth those five kings unto him out of the cave, the king of Jerusalem, the king of Hebron, the king of Jarmuth, the king of Lachish, and the king of Eglon.
JOSH|10|24|And it came to pass, when they brought out those kings unto Joshua, that Joshua called for all the men of Israel, and said unto the captains of the men of war which went with him, Come near, put your feet upon the necks of these kings. And they came near, and put their feet upon the necks of them.
JOSH|10|25|And Joshua said unto them, Fear not, nor be dismayed, be strong and of good courage: for thus shall the LORD do to all your enemies against whom ye fight.
JOSH|10|26|And afterward Joshua smote them, and slew them, and hanged them on five trees: and they were hanging upon the trees until the evening.
JOSH|10|27|And it came to pass at the time of the going down of the sun, that Joshua commanded, and they took them down off the trees, and cast them into the cave wherein they had been hid, and laid great stones in the cave's mouth, which remain until this very day.
JOSH|10|28|And that day Joshua took Makkedah, and smote it with the edge of the sword, and the king thereof he utterly destroyed, them, and all the souls that were therein; he let none remain: and he did to the king of Makkedah as he did unto the king of Jericho.
JOSH|10|29|Then Joshua passed from Makkedah, and all Israel with him, unto Libnah, and fought against Libnah:
JOSH|10|30|And the LORD delivered it also, and the king thereof, into the hand of Israel; and he smote it with the edge of the sword, and all the souls that were therein; he let none remain in it; but did unto the king thereof as he did unto the king of Jericho.
JOSH|10|31|And Joshua passed from Libnah, and all Israel with him, unto Lachish, and encamped against it, and fought against it:
JOSH|10|32|And the LORD delivered Lachish into the hand of Israel, which took it on the second day, and smote it with the edge of the sword, and all the souls that were therein, according to all that he had done to Libnah.
JOSH|10|33|Then Horam king of Gezer came up to help Lachish; and Joshua smote him and his people, until he had left him none remaining.
JOSH|10|34|And from Lachish Joshua passed unto Eglon, and all Israel with him; and they encamped against it, and fought against it:
JOSH|10|35|And they took it on that day, and smote it with the edge of the sword, and all the souls that were therein he utterly destroyed that day, according to all that he had done to Lachish.
JOSH|10|36|And Joshua went up from Eglon, and all Israel with him, unto Hebron; and they fought against it:
JOSH|10|37|And they took it, and smote it with the edge of the sword, and the king thereof, and all the cities thereof, and all the souls that were therein; he left none remaining, according to all that he had done to Eglon; but destroyed it utterly, and all the souls that were therein.
JOSH|10|38|And Joshua returned, and all Israel with him, to Debir; and fought against it:
JOSH|10|39|And he took it, and the king thereof, and all the cities thereof; and they smote them with the edge of the sword, and utterly destroyed all the souls that were therein; he left none remaining: as he had done to Hebron, so he did to Debir, and to the king thereof; as he had done also to Libnah, and to her king.
JOSH|10|40|So Joshua smote all the country of the hills, and of the south, and of the vale, and of the springs, and all their kings: he left none remaining, but utterly destroyed all that breathed, as the LORD God of Israel commanded.
JOSH|10|41|And Joshua smote them from Kadeshbarnea even unto Gaza, and all the country of Goshen, even unto Gibeon.
JOSH|10|42|And all these kings and their land did Joshua take at one time, because the LORD God of Israel fought for Israel.
JOSH|10|43|And Joshua returned, and all Israel with him, unto the camp to Gilgal.
JOSH|11|1|And it came to pass, when Jabin king of Hazor had heard those things, that he sent to Jobab king of Madon, and to the king of Shimron, and to the king of Achshaph,
JOSH|11|2|And to the kings that were on the north of the mountains, and of the plains south of Chinneroth, and in the valley, and in the borders of Dor on the west,
JOSH|11|3|And to the Canaanite on the east and on the west, and to the Amorite, and the Hittite, and the Perizzite, and the Jebusite in the mountains, and to the Hivite under Hermon in the land of Mizpeh.
JOSH|11|4|And they went out, they and all their hosts with them, much people, even as the sand that is upon the sea shore in multitude, with horses and chariots very many.
JOSH|11|5|And when all these kings were met together, they came and pitched together at the waters of Merom, to fight against Israel.
JOSH|11|6|And the LORD said unto Joshua, Be not afraid because of them: for to morrow about this time will I deliver them up all slain before Israel: thou shalt hough their horses, and burn their chariots with fire.
JOSH|11|7|So Joshua came, and all the people of war with him, against them by the waters of Merom suddenly; and they fell upon them.
JOSH|11|8|And the LORD delivered them into the hand of Israel, who smote them, and chased them unto great Zidon, and unto Misrephothmaim, and unto the valley of Mizpeh eastward; and they smote them, until they left them none remaining.
JOSH|11|9|And Joshua did unto them as the LORD bade him: he houghed their horses, and burnt their chariots with fire.
JOSH|11|10|And Joshua at that time turned back, and took Hazor, and smote the king thereof with the sword: for Hazor beforetime was the head of all those kingdoms.
JOSH|11|11|And they smote all the souls that were therein with the edge of the sword, utterly destroying them: there was not any left to breathe: and he burnt Hazor with fire.
JOSH|11|12|And all the cities of those kings, and all the kings of them, did Joshua take, and smote them with the edge of the sword, and he utterly destroyed them, as Moses the servant of the LORD commanded.
JOSH|11|13|But as for the cities that stood still in their strength, Israel burned none of them, save Hazor only; that did Joshua burn.
JOSH|11|14|And all the spoil of these cities, and the cattle, the children of Israel took for a prey unto themselves; but every man they smote with the edge of the sword, until they had destroyed them, neither left they any to breathe.
JOSH|11|15|As the LORD commanded Moses his servant, so did Moses command Joshua, and so did Joshua; he left nothing undone of all that the LORD commanded Moses.
JOSH|11|16|So Joshua took all that land, the hills, and all the south country, and all the land of Goshen, and the valley, and the plain, and the mountain of Israel, and the valley of the same;
JOSH|11|17|Even from the mount Halak, that goeth up to Seir, even unto Baalgad in the valley of Lebanon under mount Hermon: and all their kings he took, and smote them, and slew them.
JOSH|11|18|Joshua made war a long time with all those kings.
JOSH|11|19|There was not a city that made peace with the children of Israel, save the Hivites the inhabitants of Gibeon: all other they took in battle.
JOSH|11|20|For it was of the LORD to harden their hearts, that they should come against Israel in battle, that he might destroy them utterly, and that they might have no favor, but that he might destroy them, as the LORD commanded Moses.
JOSH|11|21|And at that time came Joshua, and cut off the Anakims from the mountains, from Hebron, from Debir, from Anab, and from all the mountains of Judah, and from all the mountains of Israel: Joshua destroyed them utterly with their cities.
JOSH|11|22|There was none of the Anakims left in the land of the children of Israel: only in Gaza, in Gath, and in Ashdod, there remained.
JOSH|11|23|So Joshua took the whole land, according to all that the LORD said unto Moses; and Joshua gave it for an inheritance unto Israel according to their divisions by their tribes. And the land rested from war.
JOSH|12|1|Now these are the kings of the land, which the children of Israel smote, and possessed their land on the other side Jordan toward the rising of the sun, from the river Arnon unto mount Hermon, and all the plain on the east:
JOSH|12|2|Sihon king of the Amorites, who dwelt in Heshbon, and ruled from Aroer, which is upon the bank of the river Arnon, and from the middle of the river, and from half Gilead, even unto the river Jabbok, which is the border of the children of Ammon;
JOSH|12|3|And from the plain to the sea of Chinneroth on the east, and unto the sea of the plain, even the salt sea on the east, the way to Bethjeshimoth; and from the south, under Ashdothpisgah:
JOSH|12|4|And the coast of Og king of Bashan, which was of the remnant of the giants, that dwelt at Ashtaroth and at Edrei,
JOSH|12|5|And reigned in mount Hermon, and in Salcah, and in all Bashan, unto the border of the Geshurites and the Maachathites, and half Gilead, the border of Sihon king of Heshbon.
JOSH|12|6|Them did Moses the servant of the LORD and the children of Israel smite: and Moses the servant of the LORD gave it for a possession unto the Reubenites, and the Gadites, and the half tribe of Manasseh.
JOSH|12|7|And these are the kings of the country which Joshua and the children of Israel smote on this side Jordan on the west, from Baalgad in the valley of Lebanon even unto the mount Halak, that goeth up to Seir; which Joshua gave unto the tribes of Israel for a possession according to their divisions;
JOSH|12|8|In the mountains, and in the valleys, and in the plains, and in the springs, and in the wilderness, and in the south country; the Hittites, the Amorites, and the Canaanites, the Perizzites, the Hivites, and the Jebusites:
JOSH|12|9|The king of Jericho, one; the king of Ai, which is beside Bethel, one;
JOSH|12|10|The king of Jerusalem, one; the king of Hebron, one;
JOSH|12|11|The king of Jarmuth, one; the king of Lachish, one;
JOSH|12|12|The king of Eglon, one; the king of Gezer, one;
JOSH|12|13|The king of Debir, one; the king of Geder, one;
JOSH|12|14|The king of Hormah, one; the king of Arad, one;
JOSH|12|15|The king of Libnah, one; the king of Adullam, one;
JOSH|12|16|The king of Makkedah, one; the king of Bethel, one;
JOSH|12|17|The king of Tappuah, one; the king of Hepher, one;
JOSH|12|18|The king of Aphek, one; the king of Lasharon, one;
JOSH|12|19|The king of Madon, one; the king of Hazor, one;
JOSH|12|20|The king of Shimronmeron, one; the king of Achshaph, one;
JOSH|12|21|The king of Taanach, one; the king of Megiddo, one;
JOSH|12|22|The king of Kedesh, one; the king of Jokneam of Carmel, one;
JOSH|12|23|The king of Dor in the coast of Dor, one; the king of the nations of Gilgal, one;
JOSH|12|24|The king of Tirzah, one: all the kings thirty and one.
JOSH|13|1|Now Joshua was old and stricken in years; and the LORD said unto him, Thou art old and stricken in years, and there remaineth yet very much land to be possessed.
JOSH|13|2|This is the land that yet remaineth: all the borders of the Philistines, and all Geshuri,
JOSH|13|3|From Sihor, which is before Egypt, even unto the borders of Ekron northward, which is counted to the Canaanite: five lords of the Philistines; the Gazathites, and the Ashdothites, the Eshkalonites, the Gittites, and the Ekronites; also the Avites:
JOSH|13|4|From the south, all the land of the Canaanites, and Mearah that is beside the Sidonians unto Aphek, to the borders of the Amorites:
JOSH|13|5|And the land of the Giblites, and all Lebanon, toward the sunrising, from Baalgad under mount Hermon unto the entering into Hamath.
JOSH|13|6|All the inhabitants of the hill country from Lebanon unto Misrephothmaim, and all the Sidonians, them will I drive out from before the children of Israel: only divide thou it by lot unto the Israelites for an inheritance, as I have commanded thee.
JOSH|13|7|Now therefore divide this land for an inheritance unto the nine tribes, and the half tribe of Manasseh,
JOSH|13|8|With whom the Reubenites and the Gadites have received their inheritance, which Moses gave them, beyond Jordan eastward, even as Moses the servant of the LORD gave them;
JOSH|13|9|From Aroer, that is upon the bank of the river Arnon, and the city that is in the midst of the river, and all the plain of Medeba unto Dibon;
JOSH|13|10|And all the cities of Sihon king of the Amorites, which reigned in Heshbon, unto the border of the children of Ammon;
JOSH|13|11|And Gilead, and the border of the Geshurites and Maachathites, and all mount Hermon, and all Bashan unto Salcah;
JOSH|13|12|All the kingdom of Og in Bashan, which reigned in Ashtaroth and in Edrei, who remained of the remnant of the giants: for these did Moses smite, and cast them out.
JOSH|13|13|Nevertheless the children of Israel expelled not the Geshurites, nor the Maachathites: but the Geshurites and the Maachathites dwell among the Israelites until this day.
JOSH|13|14|Only unto the tribes of Levi he gave none inheritance; the sacrifices of the LORD God of Israel made by fire are their inheritance, as he said unto them.
JOSH|13|15|And Moses gave unto the tribe of the children of Reuben inheritance according to their families.
JOSH|13|16|And their coast was from Aroer, that is on the bank of the river Arnon, and the city that is in the midst of the river, and all the plain by Medeba;
JOSH|13|17|Heshbon, and all her cities that are in the plain; Dibon, and Bamothbaal, and Bethbaalmeon,
JOSH|13|18|And Jahaza, and Kedemoth, and Mephaath,
JOSH|13|19|And Kirjathaim, and Sibmah, and Zarethshahar in the mount of the valley,
JOSH|13|20|And Bethpeor, and Ashdothpisgah, and Bethjeshimoth,
JOSH|13|21|And all the cities of the plain, and all the kingdom of Sihon king of the Amorites, which reigned in Heshbon, whom Moses smote with the princes of Midian, Evi, and Rekem, and Zur, and Hur, and Reba, which were dukes of Sihon, dwelling in the country.
JOSH|13|22|Balaam also the son of Beor, the soothsayer, did the children of Israel slay with the sword among them that were slain by them.
JOSH|13|23|And the border of the children of Reuben was Jordan, and the border thereof. This was the inheritance of the children of Reuben after their families, the cities and the villages thereof.
JOSH|13|24|And Moses gave inheritance unto the tribe of Gad, even unto the children of Gad according to their families.
JOSH|13|25|And their coast was Jazer, and all the cities of Gilead, and half the land of the children of Ammon, unto Aroer that is before Rabbah;
JOSH|13|26|And from Heshbon unto Ramathmizpeh, and Betonim; and from Mahanaim unto the border of Debir;
JOSH|13|27|And in the valley, Betharam, and Bethnimrah, and Succoth, and Zaphon, the rest of the kingdom of Sihon king of Heshbon, Jordan and his border, even unto the edge of the sea of Chinnereth on the other side Jordan eastward.
JOSH|13|28|This is the inheritance of the children of Gad after their families, the cities, and their villages.
JOSH|13|29|And Moses gave inheritance unto the half tribe of Manasseh: and this was the possession of the half tribe of the children of Manasseh by their families.
JOSH|13|30|And their coast was from Mahanaim, all Bashan, all the kingdom of Og king of Bashan, and all the towns of Jair, which are in Bashan, threescore cities:
JOSH|13|31|And half Gilead, and Ashtaroth, and Edrei, cities of the kingdom of Og in Bashan, were pertaining unto the children of Machir the son of Manasseh, even to the one half of the children of Machir by their families.
JOSH|13|32|These are the countries which Moses did distribute for inheritance in the plains of Moab, on the other side Jordan, by Jericho, eastward.
JOSH|13|33|But unto the tribe of Levi Moses gave not any inheritance: the LORD God of Israel was their inheritance, as he said unto them.
JOSH|14|1|And these are the countries which the children of Israel inherited in the land of Canaan, which Eleazar the priest, and Joshua the son of Nun, and the heads of the fathers of the tribes of the children of Israel, distributed for inheritance to them.
JOSH|14|2|By lot was their inheritance, as the LORD commanded by the hand of Moses, for the nine tribes, and for the half tribe.
JOSH|14|3|For Moses had given the inheritance of two tribes and an half tribe on the other side Jordan: but unto the Levites he gave none inheritance among them.
JOSH|14|4|For the children of Joseph were two tribes, Manasseh and Ephraim: therefore they gave no part unto the Levites in the land, save cities to dwell in, with their suburbs for their cattle and for their substance.
JOSH|14|5|As the LORD commanded Moses, so the children of Israel did, and they divided the land.
JOSH|14|6|Then the children of Judah came unto Joshua in Gilgal: and Caleb the son of Jephunneh the Kenezite said unto him, Thou knowest the thing that the LORD said unto Moses the man of God concerning me and thee in Kadeshbarnea.
JOSH|14|7|Forty years old was I when Moses the servant of the LORD sent me from Kadeshbarnea to espy out the land; and I brought him word again as it was in mine heart.
JOSH|14|8|Nevertheless my brethren that went up with me made the heart of the people melt: but I wholly followed the LORD my God.
JOSH|14|9|And Moses sware on that day, saying, Surely the land whereon thy feet have trodden shall be thine inheritance, and thy children's for ever, because thou hast wholly followed the LORD my God.
JOSH|14|10|And now, behold, the LORD hath kept me alive, as he said, these forty and five years, even since the LORD spake this word unto Moses, while the children of Israel wandered in the wilderness: and now, lo, I am this day fourscore and five years old.
JOSH|14|11|As yet I am as strong this day as I was in the day that Moses sent me: as my strength was then, even so is my strength now, for war, both to go out, and to come in.
JOSH|14|12|Now therefore give me this mountain, whereof the LORD spake in that day; for thou heardest in that day how the Anakims were there, and that the cities were great and fenced: if so be the LORD will be with me, then I shall be able to drive them out, as the LORD said.
JOSH|14|13|And Joshua blessed him, and gave unto Caleb the son of Jephunneh Hebron for an inheritance.
JOSH|14|14|Hebron therefore became the inheritance of Caleb the son of Jephunneh the Kenezite unto this day, because that he wholly followed the LORD God of Israel.
JOSH|14|15|And the name of Hebron before was Kirjatharba; which Arba was a great man among the Anakims. And the land had rest from war.
JOSH|15|1|This then was the lot of the tribe of the children of Judah by their families; even to the border of Edom the wilderness of Zin southward was the uttermost part of the south coast.
JOSH|15|2|And their south border was from the shore of the salt sea, from the bay that looketh southward:
JOSH|15|3|And it went out to the south side to Maalehacrabbim, and passed along to Zin, and ascended up on the south side unto Kadeshbarnea, and passed along to Hezron, and went up to Adar, and fetched a compass to Karkaa:
JOSH|15|4|From thence it passed toward Azmon, and went out unto the river of Egypt; and the goings out of that coast were at the sea: this shall be your south coast.
JOSH|15|5|And the east border was the salt sea, even unto the end of Jordan. And their border in the north quarter was from the bay of the sea at the uttermost part of Jordan:
JOSH|15|6|And the border went up to Bethhogla, and passed along by the north of Betharabah; and the border went up to the stone of Bohan the son of Reuben:
JOSH|15|7|And the border went up toward Debir from the valley of Achor, and so northward, looking toward Gilgal, that is before the going up to Adummim, which is on the south side of the river: and the border passed toward the waters of Enshemesh, and the goings out thereof were at Enrogel:
JOSH|15|8|And the border went up by the valley of the son of Hinnom unto the south side of the Jebusite; the same is Jerusalem: and the border went up to the top of the mountain that lieth before the valley of Hinnom westward, which is at the end of the valley of the giants northward:
JOSH|15|9|And the border was drawn from the top of the hill unto the fountain of the water of Nephtoah, and went out to the cities of mount Ephron; and the border was drawn to Baalah, which is Kirjathjearim:
JOSH|15|10|And the border compassed from Baalah westward unto mount Seir, and passed along unto the side of mount Jearim, which is Chesalon, on the north side, and went down to Bethshemesh, and passed on to Timnah:
JOSH|15|11|And the border went out unto the side of Ekron northward: and the border was drawn to Shicron, and passed along to mount Baalah, and went out unto Jabneel; and the goings out of the border were at the sea.
JOSH|15|12|And the west border was to the great sea, and the coast thereof. This is the coast of the children of Judah round about according to their families.
JOSH|15|13|And unto Caleb the son of Jephunneh he gave a part among the children of Judah, according to the commandment of the LORD to Joshua, even the city of Arba the father of Anak, which city is Hebron.
JOSH|15|14|And Caleb drove thence the three sons of Anak, Sheshai, and Ahiman, and Talmai, the children of Anak.
JOSH|15|15|And he went up thence to the inhabitants of Debir: and the name of Debir before was Kirjathsepher.
JOSH|15|16|And Caleb said, He that smiteth Kirjathsepher, and taketh it, to him will I give Achsah my daughter to wife.
JOSH|15|17|And Othniel the son of Kenaz, the brother of Caleb, took it: and he gave him Achsah his daughter to wife.
JOSH|15|18|And it came to pass, as she came unto him, that she moved him to ask of her father a field: and she lighted off her ass; and Caleb said unto her, What wouldest thou?
JOSH|15|19|Who answered, Give me a blessing; for thou hast given me a south land; give me also springs of water. And he gave her the upper springs, and the nether springs.
JOSH|15|20|This is the inheritance of the tribe of the children of Judah according to their families.
JOSH|15|21|And the uttermost cities of the tribe of the children of Judah toward the coast of Edom southward were Kabzeel, and Eder, and Jagur,
JOSH|15|22|And Kinah, and Dimonah, and Adadah,
JOSH|15|23|And Kedesh, and Hazor, and Ithnan,
JOSH|15|24|Ziph, and Telem, and Bealoth,
JOSH|15|25|And Hazor, Hadattah, and Kerioth, and Hezron, which is Hazor,
JOSH|15|26|Amam, and Shema, and Moladah,
JOSH|15|27|And Hazargaddah, and Heshmon, and Bethpalet,
JOSH|15|28|And Hazarshual, and Beersheba, and Bizjothjah,
JOSH|15|29|Baalah, and Iim, and Azem,
JOSH|15|30|And Eltolad, and Chesil, and Hormah,
JOSH|15|31|And Ziklag, and Madmannah, and Sansannah,
JOSH|15|32|And Lebaoth, and Shilhim, and Ain, and Rimmon: all the cities are twenty and nine, with their villages:
JOSH|15|33|And in the valley, Eshtaol, and Zoreah, and Ashnah,
JOSH|15|34|And Zanoah, and Engannim, Tappuah, and Enam,
JOSH|15|35|Jarmuth, and Adullam, Socoh, and Azekah,
JOSH|15|36|And Sharaim, and Adithaim, and Gederah, and Gederothaim; fourteen cities with their villages:
JOSH|15|37|Zenan, and Hadashah, and Migdalgad,
JOSH|15|38|And Dilean, and Mizpeh, and Joktheel,
JOSH|15|39|Lachish, and Bozkath, and Eglon,
JOSH|15|40|And Cabbon, and Lahmam, and Kithlish,
JOSH|15|41|And Gederoth, Bethdagon, and Naamah, and Makkedah; sixteen cities with their villages:
JOSH|15|42|Libnah, and Ether, and Ashan,
JOSH|15|43|And Jiphtah, and Ashnah, and Nezib,
JOSH|15|44|And Keilah, and Achzib, and Mareshah; nine cities with their villages:
JOSH|15|45|Ekron, with her towns and her villages:
JOSH|15|46|From Ekron even unto the sea, all that lay near Ashdod, with their villages:
JOSH|15|47|Ashdod with her towns and her villages, Gaza with her towns and her villages, unto the river of Egypt, and the great sea, and the border thereof:
JOSH|15|48|And in the mountains, Shamir, and Jattir, and Socoh,
JOSH|15|49|And Dannah, and Kirjathsannah, which is Debir,
JOSH|15|50|And Anab, and Eshtemoh, and Anim,
JOSH|15|51|And Goshen, and Holon, and Giloh; eleven cities with their villages:
JOSH|15|52|Arab, and Dumah, and Eshean,
JOSH|15|53|And Janum, and Bethtappuah, and Aphekah,
JOSH|15|54|And Humtah, and Kirjatharba, which is Hebron, and Zior; nine cities with their villages:
JOSH|15|55|Maon, Carmel, and Ziph, and Juttah,
JOSH|15|56|And Jezreel, and Jokdeam, and Zanoah,
JOSH|15|57|Cain, Gibeah, and Timnah; ten cities with their villages:
JOSH|15|58|Halhul, Bethzur, and Gedor,
JOSH|15|59|And Maarath, and Bethanoth, and Eltekon; six cities with their villages:
JOSH|15|60|Kirjathbaal, which is Kirjathjearim, and Rabbah; two cities with their villages:
JOSH|15|61|In the wilderness, Betharabah, Middin, and Secacah,
JOSH|15|62|And Nibshan, and the city of Salt, and Engedi; six cities with their villages.
JOSH|15|63|As for the Jebusites the inhabitants of Jerusalem, the children of Judah could not drive them out; but the Jebusites dwell with the children of Judah at Jerusalem unto this day.
JOSH|16|1|And the lot of the children of Joseph fell from Jordan by Jericho, unto the water of Jericho on the east, to the wilderness that goeth up from Jericho throughout mount Bethel,
JOSH|16|2|And goeth out from Bethel to Luz, and passeth along unto the borders of Archi to Ataroth,
JOSH|16|3|And goeth down westward to the coast of Japhleti, unto the coast of Bethhoron the nether, and to Gezer; and the goings out thereof are at the sea.
JOSH|16|4|So the children of Joseph, Manasseh and Ephraim, took their inheritance.
JOSH|16|5|And the border of the children of Ephraim according to their families was thus: even the border of their inheritance on the east side was Atarothaddar, unto Bethhoron the upper;
JOSH|16|6|And the border went out toward the sea to Michmethah on the north side; and the border went about eastward unto Taanathshiloh, and passed by it on the east to Janohah;
JOSH|16|7|And it went down from Janohah to Ataroth, and to Naarath, and came to Jericho, and went out at Jordan.
JOSH|16|8|The border went out from Tappuah westward unto the river Kanah; and the goings out thereof were at the sea. This is the inheritance of the tribe of the children of Ephraim by their families.
JOSH|16|9|And the separate cities for the children of Ephraim were among the inheritance of the children of Manasseh, all the cities with their villages.
JOSH|16|10|And they drave not out the Canaanites that dwelt in Gezer: but the Canaanites dwell among the Ephraimites unto this day, and serve under tribute.
JOSH|17|1|There was also a lot for the tribe of Manasseh; for he was the firstborn of Joseph; to wit, for Machir the firstborn of Manasseh, the father of Gilead: because he was a man of war, therefore he had Gilead and Bashan.
JOSH|17|2|There was also a lot for the rest of the children of Manasseh by their families; for the children of Abiezer, and for the children of Helek, and for the children of Asriel, and for the children of Shechem, and for the children of Hepher, and for the children of Shemida: these were the male children of Manasseh the son of Joseph by their families.
JOSH|17|3|But Zelophehad, the son of Hepher, the son of Gilead, the son of Machir, the son of Manasseh, had no sons, but daughters: and these are the names of his daughters, Mahlah, and Noah, Hoglah, Milcah, and Tirzah.
JOSH|17|4|And they came near before Eleazar the priest, and before Joshua the son of Nun, and before the princes, saying, The LORD commanded Moses to give us an inheritance among our brethren. Therefore according to the commandment of the LORD he gave them an inheritance among the brethren of their father.
JOSH|17|5|And there fell ten portions to Manasseh, beside the land of Gilead and Bashan, which were on the other side Jordan;
JOSH|17|6|Because the daughters of Manasseh had an inheritance among his sons: and the rest of Manasseh's sons had the land of Gilead.
JOSH|17|7|And the coast of Manasseh was from Asher to Michmethah, that lieth before Shechem; and the border went along on the right hand unto the inhabitants of Entappuah.
JOSH|17|8|Now Manasseh had the land of Tappuah: but Tappuah on the border of Manasseh belonged to the children of Ephraim;
JOSH|17|9|And the coast descended unto the river Kanah, southward of the river: these cities of Ephraim are among the cities of Manasseh: the coast of Manasseh also was on the north side of the river, and the outgoings of it were at the sea:
JOSH|17|10|Southward it was Ephraim's, and northward it was Manasseh's, and the sea is his border; and they met together in Asher on the north, and in Issachar on the east.
JOSH|17|11|And Manasseh had in Issachar and in Asher Bethshean and her towns, and Ibleam and her towns, and the inhabitants of Dor and her towns, and the inhabitants of Endor and her towns, and the inhabitants of Taanach and her towns, and the inhabitants of Megiddo and her towns, even three countries.
JOSH|17|12|Yet the children of Manasseh could not drive out the inhabitants of those cities; but the Canaanites would dwell in that land.
JOSH|17|13|Yet it came to pass, when the children of Israel were waxen strong, that they put the Canaanites to tribute, but did not utterly drive them out.
JOSH|17|14|And the children of Joseph spake unto Joshua, saying, Why hast thou given me but one lot and one portion to inherit, seeing I am a great people, forasmuch as the LORD hath blessed me hitherto?
JOSH|17|15|And Joshua answered them, If thou be a great people, then get thee up to the wood country, and cut down for thyself there in the land of the Perizzites and of the giants, if mount Ephraim be too narrow for thee.
JOSH|17|16|And the children of Joseph said, The hill is not enough for us: and all the Canaanites that dwell in the land of the valley have chariots of iron, both they who are of Bethshean and her towns, and they who are of the valley of Jezreel.
JOSH|17|17|And Joshua spake unto the house of Joseph, even to Ephraim and to Manasseh, saying, Thou art a great people, and hast great power: thou shalt not have one lot only:
JOSH|17|18|But the mountain shall be thine; for it is a wood, and thou shalt cut it down: and the outgoings of it shall be thine: for thou shalt drive out the Canaanites, though they have iron chariots, and though they be strong.
JOSH|18|1|And the whole congregation of the children of Israel assembled together at Shiloh, and set up the tabernacle of the congregation there. And the land was subdued before them.
JOSH|18|2|And there remained among the children of Israel seven tribes, which had not yet received their inheritance.
JOSH|18|3|And Joshua said unto the children of Israel, How long are ye slack to go to possess the land, which the LORD God of your fathers hath given you?
JOSH|18|4|Give out from among you three men for each tribe: and I will send them, and they shall rise, and go through the land, and describe it according to the inheritance of them; and they shall come again to me.
JOSH|18|5|And they shall divide it into seven parts: Judah shall abide in their coast on the south, and the house of Joseph shall abide in their coasts on the north.
JOSH|18|6|Ye shall therefore describe the land into seven parts, and bring the description hither to me, that I may cast lots for you here before the LORD our God.
JOSH|18|7|But the Levites have no part among you; for the priesthood of the LORD is their inheritance: and Gad, and Reuben, and half the tribe of Manasseh, have received their inheritance beyond Jordan on the east, which Moses the servant of the LORD gave them.
JOSH|18|8|And the men arose, and went away: and Joshua charged them that went to describe the land, saying, Go and walk through the land, and describe it, and come again to me, that I may here cast lots for you before the LORD in Shiloh.
JOSH|18|9|And the men went and passed through the land, and described it by cities into seven parts in a book, and came again to Joshua to the host at Shiloh.
JOSH|18|10|And Joshua cast lots for them in Shiloh before the LORD: and there Joshua divided the land unto the children of Israel according to their divisions.
JOSH|18|11|And the lot of the tribe of the children of Benjamin came up according to their families: and the coast of their lot came forth between the children of Judah and the children of Joseph.
JOSH|18|12|And their border on the north side was from Jordan; and the border went up to the side of Jericho on the north side, and went up through the mountains westward; and the goings out thereof were at the wilderness of Bethaven.
JOSH|18|13|And the border went over from thence toward Luz, to the side of Luz, which is Bethel, southward; and the border descended to Atarothadar, near the hill that lieth on the south side of the nether Bethhoron.
JOSH|18|14|And the border was drawn thence, and compassed the corner of the sea southward, from the hill that lieth before Bethhoron southward; and the goings out thereof were at Kirjathbaal, which is Kirjathjearim, a city of the children of Judah: this was the west quarter.
JOSH|18|15|And the south quarter was from the end of Kirjathjearim, and the border went out on the west, and went out to the well of waters of Nephtoah:
JOSH|18|16|And the border came down to the end of the mountain that lieth before the valley of the son of Hinnom, and which is in the valley of the giants on the north, and descended to the valley of Hinnom, to the side of Jebusi on the south, and descended to Enrogel,
JOSH|18|17|And was drawn from the north, and went forth to Enshemesh, and went forth toward Geliloth, which is over against the going up of Adummim, and descended to the stone of Bohan the son of Reuben,
JOSH|18|18|And passed along toward the side over against Arabah northward, and went down unto Arabah:
JOSH|18|19|And the border passed along to the side of Bethhoglah northward: and the outgoings of the border were at the north bay of the salt sea at the south end of Jordan: this was the south coast.
JOSH|18|20|And Jordan was the border of it on the east side. This was the inheritance of the children of Benjamin, by the coasts thereof round about, according to their families.
JOSH|18|21|Now the cities of the tribe of the children of Benjamin according to their families were Jericho, and Bethhoglah, and the valley of Keziz,
JOSH|18|22|And Betharabah, and Zemaraim, and Bethel,
JOSH|18|23|And Avim, and Pharah, and Ophrah,
JOSH|18|24|And Chepharhaammonai, and Ophni, and Gaba; twelve cities with their villages:
JOSH|18|25|Gibeon, and Ramah, and Beeroth,
JOSH|18|26|And Mizpeh, and Chephirah, and Mozah,
JOSH|18|27|And Rekem, and Irpeel, and Taralah,
JOSH|18|28|And Zelah, Eleph, and Jebusi, which is Jerusalem, Gibeath, and Kirjath; fourteen cities with their villages. This is the inheritance of the children of Benjamin according to their families.
JOSH|19|1|And the second lot came forth to Simeon, even for the tribe of the children of Simeon according to their families: and their inheritance was within the inheritance of the children of Judah.
JOSH|19|2|And they had in their inheritance Beersheba, and Sheba, and Moladah,
JOSH|19|3|And Hazarshual, and Balah, and Azem,
JOSH|19|4|And Eltolad, and Bethul, and Hormah,
JOSH|19|5|And Ziklag, and Bethmarcaboth, and Hazarsusah,
JOSH|19|6|And Bethlebaoth, and Sharuhen; thirteen cities and their villages:
JOSH|19|7|Ain, Remmon, and Ether, and Ashan; four cities and their villages:
JOSH|19|8|And all the villages that were round about these cities to Baalathbeer, Ramath of the south. This is the inheritance of the tribe of the children of Simeon according to their families.
JOSH|19|9|Out of the portion of the children of Judah was the inheritance of the children of Simeon: for the part of the children of Judah was too much for them: therefore the children of Simeon had their inheritance within the inheritance of them.
JOSH|19|10|And the third lot came up for the children of Zebulun according to their families: and the border of their inheritance was unto Sarid:
JOSH|19|11|And their border went up toward the sea, and Maralah, and reached to Dabbasheth, and reached to the river that is before Jokneam;
JOSH|19|12|And turned from Sarid eastward toward the sunrising unto the border of Chislothtabor, and then goeth out to Daberath, and goeth up to Japhia,
JOSH|19|13|And from thence passeth on along on the east to Gittahhepher, to Ittahkazin, and goeth out to Remmonmethoar to Neah;
JOSH|19|14|And the border compasseth it on the north side to Hannathon: and the outgoings thereof are in the valley of Jiphthahel:
JOSH|19|15|And Kattath, and Nahallal, and Shimron, and Idalah, and Bethlehem: twelve cities with their villages.
JOSH|19|16|This is the inheritance of the children of Zebulun according to their families, these cities with their villages.
JOSH|19|17|And the fourth lot came out to Issachar, for the children of Issachar according to their families.
JOSH|19|18|And their border was toward Jezreel, and Chesulloth, and Shunem,
JOSH|19|19|And Haphraim, and Shihon, and Anaharath,
JOSH|19|20|And Rabbith, and Kishion, and Abez,
JOSH|19|21|And Remeth, and Engannim, and Enhaddah, and Bethpazzez;
JOSH|19|22|And the coast reacheth to Tabor, and Shahazimah, and Bethshemesh; and the outgoings of their border were at Jordan: sixteen cities with their villages.
JOSH|19|23|This is the inheritance of the tribe of the children of Issachar according to their families, the cities and their villages.
JOSH|19|24|And the fifth lot came out for the tribe of the children of Asher according to their families.
JOSH|19|25|And their border was Helkath, and Hali, and Beten, and Achshaph,
JOSH|19|26|And Alammelech, and Amad, and Misheal; and reacheth to Carmel westward, and to Shihorlibnath;
JOSH|19|27|And turneth toward the sunrising to Bethdagon, and reacheth to Zebulun, and to the valley of Jiphthahel toward the north side of Bethemek, and Neiel, and goeth out to Cabul on the left hand,
JOSH|19|28|And Hebron, and Rehob, and Hammon, and Kanah, even unto great Zidon;
JOSH|19|29|And then the coast turneth to Ramah, and to the strong city Tyre; and the coast turneth to Hosah; and the outgoings thereof are at the sea from the coast to Achzib:
JOSH|19|30|Ummah also, and Aphek, and Rehob: twenty and two cities with their villages.
JOSH|19|31|This is the inheritance of the tribe of the children of Asher according to their families, these cities with their villages.
JOSH|19|32|The sixth lot came out to the children of Naphtali, even for the children of Naphtali according to their families.
JOSH|19|33|And their coast was from Heleph, from Allon to Zaanannim, and Adami, Nekeb, and Jabneel, unto Lakum; and the outgoings thereof were at Jordan:
JOSH|19|34|And then the coast turneth westward to Aznothtabor, and goeth out from thence to Hukkok, and reacheth to Zebulun on the south side, and reacheth to Asher on the west side, and to Judah upon Jordan toward the sunrising.
JOSH|19|35|And the fenced cities are Ziddim, Zer, and Hammath, Rakkath, and Chinnereth,
JOSH|19|36|And Adamah, and Ramah, and Hazor,
JOSH|19|37|And Kedesh, and Edrei, and Enhazor,
JOSH|19|38|And Iron, and Migdalel, Horem, and Bethanath, and Bethshemesh; nineteen cities with their villages.
JOSH|19|39|This is the inheritance of the tribe of the children of Naphtali according to their families, the cities and their villages.
JOSH|19|40|And the seventh lot came out for the tribe of the children of Dan according to their families.
JOSH|19|41|And the coast of their inheritance was Zorah, and Eshtaol, and Irshemesh,
JOSH|19|42|And Shaalabbin, and Ajalon, and Jethlah,
JOSH|19|43|And Elon, and Thimnathah, and Ekron,
JOSH|19|44|And Eltekeh, and Gibbethon, and Baalath,
JOSH|19|45|And Jehud, and Beneberak, and Gathrimmon,
JOSH|19|46|And Mejarkon, and Rakkon, with the border before Japho.
JOSH|19|47|And the coast of the children of Dan went out too little for them: therefore the children of Dan went up to fight against Leshem, and took it, and smote it with the edge of the sword, and possessed it, and dwelt therein, and called Leshem, Dan, after the name of Dan their father.
JOSH|19|48|This is the inheritance of the tribe of the children of Dan according to their families, these cities with their villages.
JOSH|19|49|When they had made an end of dividing the land for inheritance by their coasts, the children of Israel gave an inheritance to Joshua the son of Nun among them:
JOSH|19|50|According to the word of the LORD they gave him the city which he asked, even Timnathserah in mount Ephraim: and he built the city, and dwelt therein.
JOSH|19|51|These are the inheritances, which Eleazar the priest, and Joshua the son of Nun, and the heads of the fathers of the tribes of the children of Israel, divided for an inheritance by lot in Shiloh before the LORD, at the door of the tabernacle of the congregation. So they made an end of dividing the country.
JOSH|20|1|The LORD also spake unto Joshua, saying,
JOSH|20|2|Speak to the children of Israel, saying, Appoint out for you cities of refuge, whereof I spake unto you by the hand of Moses:
JOSH|20|3|That the slayer that killeth any person unawares and unwittingly may flee thither: and they shall be your refuge from the avenger of blood.
JOSH|20|4|And when he that doth flee unto one of those cities shall stand at the entering of the gate of the city, and shall declare his cause in the ears of the elders of that city, they shall take him into the city unto them, and give him a place, that he may dwell among them.
JOSH|20|5|And if the avenger of blood pursue after him, then they shall not deliver the slayer up into his hand; because he smote his neighbor unwittingly, and hated him not beforetime.
JOSH|20|6|And he shall dwell in that city, until he stand before the congregation for judgment, and until the death of the high priest that shall be in those days: then shall the slayer return, and come unto his own city, and unto his own house, unto the city from whence he fled.
JOSH|20|7|And they appointed Kedesh in Galilee in mount Naphtali, and Shechem in mount Ephraim, and Kirjatharba, which is Hebron, in the mountain of Judah.
JOSH|20|8|And on the other side Jordan by Jericho eastward, they assigned Bezer in the wilderness upon the plain out of the tribe of Reuben, and Ramoth in Gilead out of the tribe of Gad, and Golan in Bashan out of the tribe of Manasseh.
JOSH|20|9|These were the cities appointed for all the children of Israel, and for the stranger that sojourneth among them, that whosoever killeth any person at unawares might flee thither, and not die by the hand of the avenger of blood, until he stood before the congregation.
JOSH|21|1|Then came near the heads of the fathers of the Levites unto Eleazar the priest, and unto Joshua the son of Nun, and unto the heads of the fathers of the tribes of the children of Israel;
JOSH|21|2|And they spake unto them at Shiloh in the land of Canaan, saying, The LORD commanded by the hand of Moses to give us cities to dwell in, with the suburbs thereof for our cattle.
JOSH|21|3|And the children of Israel gave unto the Levites out of their inheritance, at the commandment of the LORD, these cities and their suburbs.
JOSH|21|4|And the lot came out for the families of the Kohathites: and the children of Aaron the priest, which were of the Levites, had by lot out of the tribe of Judah, and out of the tribe of Simeon, and out of the tribe of Benjamin, thirteen cities.
JOSH|21|5|And the rest of the children of Kohath had by lot out of the families of the tribe of Ephraim, and out of the tribe of Dan, and out of the half tribe of Manasseh, ten cities.
JOSH|21|6|And the children of Gershon had by lot out of the families of the tribe of Issachar, and out of the tribe of Asher, and out of the tribe of Naphtali, and out of the half tribe of Manasseh in Bashan, thirteen cities.
JOSH|21|7|The children of Merari by their families had out of the tribe of Reuben, and out of the tribe of Gad, and out of the tribe of Zebulun, twelve cities.
JOSH|21|8|And the children of Israel gave by lot unto the Levites these cities with their suburbs, as the LORD commanded by the hand of Moses.
JOSH|21|9|And they gave out of the tribe of the children of Judah, and out of the tribe of the children of Simeon, these cities which are here mentioned by name.
JOSH|21|10|Which the children of Aaron, being of the families of the Kohathites, who were of the children of Levi, had: for theirs was the first lot.
JOSH|21|11|And they gave them the city of Arba the father of Anak, which city is Hebron, in the hill country of Judah, with the suburbs thereof round about it.
JOSH|21|12|But the fields of the city, and the villages thereof, gave they to Caleb the son of Jephunneh for his possession.
JOSH|21|13|Thus they gave to the children of Aaron the priest Hebron with her suburbs, to be a city of refuge for the slayer; and Libnah with her suburbs,
JOSH|21|14|And Jattir with her suburbs, and Eshtemoa with her suburbs,
JOSH|21|15|And Holon with her suburbs, and Debir with her suburbs,
JOSH|21|16|And Ain with her suburbs, and Juttah with her suburbs, and Bethshemesh with her suburbs; nine cities out of those two tribes.
JOSH|21|17|And out of the tribe of Benjamin, Gibeon with her suburbs, Geba with her suburbs,
JOSH|21|18|Anathoth with her suburbs, and Almon with her suburbs; four cities.
JOSH|21|19|All the cities of the children of Aaron, the priests, were thirteen cities with their suburbs.
JOSH|21|20|And the families of the children of Kohath, the Levites which remained of the children of Kohath, even they had the cities of their lot out of the tribe of Ephraim.
JOSH|21|21|For they gave them Shechem with her suburbs in mount Ephraim, to be a city of refuge for the slayer; and Gezer with her suburbs,
JOSH|21|22|And Kibzaim with her suburbs, and Bethhoron with her suburbs; four cities.
JOSH|21|23|And out of the tribe of Dan, Eltekeh with her suburbs, Gibbethon with her suburbs,
JOSH|21|24|Aijalon with her suburbs, Gathrimmon with her suburbs; four cities.
JOSH|21|25|And out of the half tribe of Manasseh, Tanach with her suburbs, and Gathrimmon with her suburbs; two cities.
JOSH|21|26|All the cities were ten with their suburbs for the families of the children of Kohath that remained.
JOSH|21|27|And unto the children of Gershon, of the families of the Levites, out of the other half tribe of Manasseh they gave Golan in Bashan with her suburbs, to be a city of refuge for the slayer; and Beeshterah with her suburbs; two cities.
JOSH|21|28|And out of the tribe of Issachar, Kishon with her suburbs, Dabareh with her suburbs,
JOSH|21|29|Jarmuth with her suburbs, Engannim with her suburbs; four cities.
JOSH|21|30|And out of the tribe of Asher, Mishal with her suburbs, Abdon with her suburbs,
JOSH|21|31|Helkath with her suburbs, and Rehob with her suburbs; four cities.
JOSH|21|32|And out of the tribe of Naphtali, Kedesh in Galilee with her suburbs, to be a city of refuge for the slayer; and Hammothdor with her suburbs, and Kartan with her suburbs; three cities.
JOSH|21|33|All the cities of the Gershonites according to their families were thirteen cities with their suburbs.
JOSH|21|34|And unto the families of the children of Merari, the rest of the Levites, out of the tribe of Zebulun, Jokneam with her suburbs, and Kartah with her suburbs,
JOSH|21|35|Dimnah with her suburbs, Nahalal with her suburbs; four cities.
JOSH|21|36|And out of the tribe of Reuben, Bezer with her suburbs, and Jahazah with her suburbs,
JOSH|21|37|Kedemoth with her suburbs, and Mephaath with her suburbs; four cities.
JOSH|21|38|And out of the tribe of Gad, Ramoth in Gilead with her suburbs, to be a city of refuge for the slayer; and Mahanaim with her suburbs,
JOSH|21|39|Heshbon with her suburbs, Jazer with her suburbs; four cities in all.
JOSH|21|40|So all the cities for the children of Merari by their families, which were remaining of the families of the Levites, were by their lot twelve cities.
JOSH|21|41|All the cities of the Levites within the possession of the children of Israel were forty and eight cities with their suburbs.
JOSH|21|42|These cities were every one with their suburbs round about them: thus were all these cities.
JOSH|21|43|And the LORD gave unto Israel all the land which he sware to give unto their fathers; and they possessed it, and dwelt therein.
JOSH|21|44|And the LORD gave them rest round about, according to all that he sware unto their fathers: and there stood not a man of all their enemies before them; the LORD delivered all their enemies into their hand.
JOSH|21|45|There failed not ought of any good thing which the LORD had spoken unto the house of Israel; all came to pass.
JOSH|22|1|Then Joshua called the Reubenites, and the Gadites, and the half tribe of Manasseh,
JOSH|22|2|And said unto them, Ye have kept all that Moses the servant of the LORD commanded you, and have obeyed my voice in all that I commanded you:
JOSH|22|3|Ye have not left your brethren these many days unto this day, but have kept the charge of the commandment of the LORD your God.
JOSH|22|4|And now the LORD your God hath given rest unto your brethren, as he promised them: therefore now return ye, and get you unto your tents, and unto the land of your possession, which Moses the servant of the LORD gave you on the other side Jordan.
JOSH|22|5|But take diligent heed to do the commandment and the law, which Moses the servant of the LORD charged you, to love the LORD your God, and to walk in all his ways, and to keep his commandments, and to cleave unto him, and to serve him with all your heart and with all your soul.
JOSH|22|6|So Joshua blessed them, and sent them away: and they went unto their tents.
JOSH|22|7|Now to the one half of the tribe of Manasseh Moses had given possession in Bashan: but unto the other half thereof gave Joshua among their brethren on this side Jordan westward. And when Joshua sent them away also unto their tents, then he blessed them,
JOSH|22|8|And he spake unto them, saying, Return with much riches unto your tents, and with very much cattle, with silver, and with gold, and with brass, and with iron, and with very much raiment: divide the spoil of your enemies with your brethren.
JOSH|22|9|And the children of Reuben and the children of Gad and the half tribe of Manasseh returned, and departed from the children of Israel out of Shiloh, which is in the land of Canaan, to go unto the country of Gilead, to the land of their possession, whereof they were possessed, according to the word of the LORD by the hand of Moses.
JOSH|22|10|And when they came unto the borders of Jordan, that are in the land of Canaan, the children of Reuben and the children of Gad and the half tribe of Manasseh built there an altar by Jordan, a great altar to see to.
JOSH|22|11|And the children of Israel heard say, Behold, the children of Reuben and the children of Gad and the half tribe of Manasseh have built an altar over against the land of Canaan, in the borders of Jordan, at the passage of the children of Israel.
JOSH|22|12|And when the children of Israel heard of it, the whole congregation of the children of Israel gathered themselves together at Shiloh, to go up to war against them.
JOSH|22|13|And the children of Israel sent unto the children of Reuben, and to the children of Gad, and to the half tribe of Manasseh, into the land of Gilead, Phinehas the son of Eleazar the priest,
JOSH|22|14|And with him ten princes, of each chief house a prince throughout all the tribes of Israel; and each one was an head of the house of their fathers among the thousands of Israel.
JOSH|22|15|And they came unto the children of Reuben, and to the children of Gad, and to the half tribe of Manasseh, unto the land of Gilead, and they spake with them, saying,
JOSH|22|16|Thus saith the whole congregation of the LORD, What trespass is this that ye have committed against the God of Israel, to turn away this day from following the LORD, in that ye have builded you an altar, that ye might rebel this day against the LORD?
JOSH|22|17|Is the iniquity of Peor too little for us, from which we are not cleansed until this day, although there was a plague in the congregation of the LORD,
JOSH|22|18|But that ye must turn away this day from following the LORD? and it will be, seeing ye rebel to day against the LORD, that to morrow he will be wroth with the whole congregation of Israel.
JOSH|22|19|Notwithstanding, if the land of your possession be unclean, then pass ye over unto the land of the possession of the LORD, wherein the LORD's tabernacle dwelleth, and take possession among us: but rebel not against the LORD, nor rebel against us, in building you an altar beside the altar of the LORD our God.
JOSH|22|20|Did not Achan the son of Zerah commit a trespass in the accursed thing, and wrath fell on all the congregation of Israel? and that man perished not alone in his iniquity.
JOSH|22|21|Then the children of Reuben and the children of Gad and the half tribe of Manasseh answered, and said unto the heads of the thousands of Israel,
JOSH|22|22|The LORD God of gods, the LORD God of gods, he knoweth, and Israel he shall know; if it be in rebellion, or if in transgression against the LORD, (save us not this day,)
JOSH|22|23|That we have built us an altar to turn from following the LORD, or if to offer thereon burnt offering or meat offering, or if to offer peace offerings thereon, let the LORD himself require it;
JOSH|22|24|And if we have not rather done it for fear of this thing, saying, In time to come your children might speak unto our children, saying, What have ye to do with the LORD God of Israel?
JOSH|22|25|For the LORD hath made Jordan a border between us and you, ye children of Reuben and children of Gad; ye have no part in the LORD: so shall your children make our children cease from fearing the LORD.
JOSH|22|26|Therefore we said, Let us now prepare to build us an altar, not for burnt offering, nor for sacrifice:
JOSH|22|27|But that it may be a witness between us, and you, and our generations after us, that we might do the service of the LORD before him with our burnt offerings, and with our sacrifices, and with our peace offerings; that your children may not say to our children in time to come, Ye have no part in the LORD.
JOSH|22|28|Therefore said we, that it shall be, when they should so say to us or to our generations in time to come, that we may say again, Behold the pattern of the altar of the LORD, which our fathers made, not for burnt offerings, nor for sacrifices; but it is a witness between us and you.
JOSH|22|29|God forbid that we should rebel against the LORD, and turn this day from following the LORD, to build an altar for burnt offerings, for meat offerings, or for sacrifices, beside the altar of the LORD our God that is before his tabernacle.
JOSH|22|30|And when Phinehas the priest, and the princes of the congregation and heads of the thousands of Israel which were with him, heard the words that the children of Reuben and the children of Gad and the children of Manasseh spake, it pleased them.
JOSH|22|31|And Phinehas the son of Eleazar the priest said unto the children of Reuben, and to the children of Gad, and to the children of Manasseh, This day we perceive that the LORD is among us, because ye have not committed this trespass against the LORD: now ye have delivered the children of Israel out of the hand of the LORD.
JOSH|22|32|And Phinehas the son of Eleazar the priest, and the princes, returned from the children of Reuben, and from the children of Gad, out of the land of Gilead, unto the land of Canaan, to the children of Israel, and brought them word again.
JOSH|22|33|And the thing pleased the children of Israel; and the children of Israel blessed God, and did not intend to go up against them in battle, to destroy the land wherein the children of Reuben and Gad dwelt.
JOSH|22|34|And the children of Reuben and the children of Gad called the altar Ed: for it shall be a witness between us that the LORD is God.
JOSH|23|1|And it came to pass a long time after that the LORD had given rest unto Israel from all their enemies round about, that Joshua waxed old and stricken in age.
JOSH|23|2|And Joshua called for all Israel, and for their elders, and for their heads, and for their judges, and for their officers, and said unto them, I am old and stricken in age:
JOSH|23|3|And ye have seen all that the LORD your God hath done unto all these nations because of you; for the LORD your God is he that hath fought for you.
JOSH|23|4|Behold, I have divided unto you by lot these nations that remain, to be an inheritance for your tribes, from Jordan, with all the nations that I have cut off, even unto the great sea westward.
JOSH|23|5|And the LORD your God, he shall expel them from before you, and drive them from out of your sight; and ye shall possess their land, as the LORD your God hath promised unto you.
JOSH|23|6|Be ye therefore very courageous to keep and to do all that is written in the book of the law of Moses, that ye turn not aside therefrom to the right hand or to the left;
JOSH|23|7|That ye come not among these nations, these that remain among you; neither make mention of the name of their gods, nor cause to swear by them, neither serve them, nor bow yourselves unto them:
JOSH|23|8|But cleave unto the LORD your God, as ye have done unto this day.
JOSH|23|9|For the LORD hath driven out from before you great nations and strong: but as for you, no man hath been able to stand before you unto this day.
JOSH|23|10|One man of you shall chase a thousand: for the LORD your God, he it is that fighteth for you, as he hath promised you.
JOSH|23|11|Take good heed therefore unto yourselves, that ye love the LORD your God.
JOSH|23|12|Else if ye do in any wise go back, and cleave unto the remnant of these nations, even these that remain among you, and shall make marriages with them, and go in unto them, and they to you:
JOSH|23|13|Know for a certainty that the LORD your God will no more drive out any of these nations from before you; but they shall be snares and traps unto you, and scourges in your sides, and thorns in your eyes, until ye perish from off this good land which the LORD your God hath given you.
JOSH|23|14|And, behold, this day I am going the way of all the earth: and ye know in all your hearts and in all your souls, that not one thing hath failed of all the good things which the LORD your God spake concerning you; all are come to pass unto you, and not one thing hath failed thereof.
JOSH|23|15|Therefore it shall come to pass, that as all good things are come upon you, which the LORD your God promised you; so shall the LORD bring upon you all evil things, until he have destroyed you from off this good land which the LORD your God hath given you.
JOSH|23|16|When ye have transgressed the covenant of the LORD your God, which he commanded you, and have gone and served other gods, and bowed yourselves to them; then shall the anger of the LORD be kindled against you, and ye shall perish quickly from off the good land which he hath given unto you.
JOSH|24|1|And Joshua gathered all the tribes of Israel to Shechem, and called for the elders of Israel, and for their heads, and for their judges, and for their officers; and they presented themselves before God.
JOSH|24|2|And Joshua said unto all the people, Thus saith the LORD God of Israel, Your fathers dwelt on the other side of the flood in old time, even Terah, the father of Abraham, and the father of Nachor: and they served other gods.
JOSH|24|3|And I took your father Abraham from the other side of the flood, and led him throughout all the land of Canaan, and multiplied his seed, and gave him Isaac.
JOSH|24|4|And I gave unto Isaac Jacob and Esau: and I gave unto Esau mount Seir, to possess it; but Jacob and his children went down into Egypt.
JOSH|24|5|I sent Moses also and Aaron, and I plagued Egypt, according to that which I did among them: and afterward I brought you out.
JOSH|24|6|And I brought your fathers out of Egypt: and ye came unto the sea; and the Egyptians pursued after your fathers with chariots and horsemen unto the Red sea.
JOSH|24|7|And when they cried unto the LORD, he put darkness between you and the Egyptians, and brought the sea upon them, and covered them; and your eyes have seen what I have done in Egypt: and ye dwelt in the wilderness a long season.
JOSH|24|8|And I brought you into the land of the Amorites, which dwelt on the other side Jordan; and they fought with you: and I gave them into your hand, that ye might possess their land; and I destroyed them from before you.
JOSH|24|9|Then Balak the son of Zippor, king of Moab, arose and warred against Israel, and sent and called Balaam the son of Beor to curse you:
JOSH|24|10|But I would not hearken unto Balaam; therefore he blessed you still: so I delivered you out of his hand.
JOSH|24|11|And you went over Jordan, and came unto Jericho: and the men of Jericho fought against you, the Amorites, and the Perizzites, and the Canaanites, and the Hittites, and the Girgashites, the Hivites, and the Jebusites; and I delivered them into your hand.
JOSH|24|12|And I sent the hornet before you, which drave them out from before you, even the two kings of the Amorites; but not with thy sword, nor with thy bow.
JOSH|24|13|And I have given you a land for which ye did not labor, and cities which ye built not, and ye dwell in them; of the vineyards and oliveyards which ye planted not do ye eat.
JOSH|24|14|Now therefore fear the LORD, and serve him in sincerity and in truth: and put away the gods which your fathers served on the other side of the flood, and in Egypt; and serve ye the LORD.
JOSH|24|15|And if it seem evil unto you to serve the LORD, choose you this day whom ye will serve; whether the gods which your fathers served that were on the other side of the flood, or the gods of the Amorites, in whose land ye dwell: but as for me and my house, we will serve the LORD.
JOSH|24|16|And the people answered and said, God forbid that we should forsake the LORD, to serve other gods;
JOSH|24|17|For the LORD our God, he it is that brought us up and our fathers out of the land of Egypt, from the house of bondage, and which did those great signs in our sight, and preserved us in all the way wherein we went, and among all the people through whom we passed:
JOSH|24|18|And the LORD drave out from before us all the people, even the Amorites which dwelt in the land: therefore will we also serve the LORD; for he is our God.
JOSH|24|19|And Joshua said unto the people, Ye cannot serve the LORD: for he is an holy God; he is a jealous God; he will not forgive your transgressions nor your sins.
JOSH|24|20|If ye forsake the LORD, and serve strange gods, then he will turn and do you hurt, and consume you, after that he hath done you good.
JOSH|24|21|And the people said unto Joshua, Nay; but we will serve the LORD.
JOSH|24|22|And Joshua said unto the people, Ye are witnesses against yourselves that ye have chosen you the LORD, to serve him. And they said, We are witnesses.
JOSH|24|23|Now therefore put away, said he, the strange gods which are among you, and incline your heart unto the LORD God of Israel.
JOSH|24|24|And the people said unto Joshua, The LORD our God will we serve, and his voice will we obey.
JOSH|24|25|So Joshua made a covenant with the people that day, and set them a statute and an ordinance in Shechem.
JOSH|24|26|And Joshua wrote these words in the book of the law of God, and took a great stone, and set it up there under an oak, that was by the sanctuary of the LORD.
JOSH|24|27|And Joshua said unto all the people, Behold, this stone shall be a witness unto us; for it hath heard all the words of the LORD which he spake unto us: it shall be therefore a witness unto you, lest ye deny your God.
JOSH|24|28|So Joshua let the people depart, every man unto his inheritance.
JOSH|24|29|And it came to pass after these things, that Joshua the son of Nun, the servant of the LORD, died, being an hundred and ten years old.
JOSH|24|30|And they buried him in the border of his inheritance in Timnathserah, which is in mount Ephraim, on the north side of the hill of Gaash.
JOSH|24|31|And Israel served the LORD all the days of Joshua, and all the days of the elders that overlived Joshua, and which had known all the works of the LORD, that he had done for Israel.
JOSH|24|32|And the bones of Joseph, which the children of Israel brought up out of Egypt, buried they in Shechem, in a parcel of ground which Jacob bought of the sons of Hamor the father of Shechem for an hundred pieces of silver: and it became the inheritance of the children of Joseph.
JOSH|24|33|And Eleazar the son of Aaron died; and they buried him in a hill that pertained to Phinehas his son, which was given him in mount Ephraim.
