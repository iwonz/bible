JAS|1|1|James, a servant of God and of the Lord Jesus Christ, To the twelve tribes in the Dispersion: Greetings.
JAS|1|2|Count it all joy, my brothers, when you meet trials of various kinds,
JAS|1|3|for you know that the testing of your faith produces steadfastness.
JAS|1|4|And let steadfastness have its full effect, that you may be perfect and complete, lacking in nothing.
JAS|1|5|If any of you lacks wisdom, let him ask God, who gives generously to all without reproach, and it will be given him.
JAS|1|6|But let him ask in faith, with no doubting, for the one who doubts is like a wave of the sea that is driven and tossed by the wind.
JAS|1|7|For that person must not suppose that he will receive anything from the Lord;
JAS|1|8|he is a double-minded man, unstable in all his ways.
JAS|1|9|Let the lowly brother boast in his exaltation,
JAS|1|10|and the rich in his humiliation, because like a flower of the grass he will pass away.
JAS|1|11|For the sun rises with its scorching heat and withers the grass; its flower falls, and its beauty perishes. So also will the rich man fade away in the midst of his pursuits.
JAS|1|12|Blessed is the man who remains steadfast under trial, for when he has stood the test he will receive the crown of life, which God has promised to those who love him.
JAS|1|13|Let no one say when he is tempted, "I am being tempted by God," for God cannot be tempted with evil, and he himself tempts no one.
JAS|1|14|But each person is tempted when he is lured and enticed by his own desire.
JAS|1|15|Then desire when it has conceived gives birth to sin, and sin when it is fully grown brings forth death.
JAS|1|16|Do not be deceived, my beloved brothers.
JAS|1|17|Every good gift and every perfect gift is from above, coming down from the Father of lights with whom there is no variation or shadow due to change.
JAS|1|18|Of his own will he brought us forth by the word of truth, that we should be a kind of firstfruits of his creation.
JAS|1|19|Know this, my beloved brothers: let every person be quick to hear, slow to speak, slow to anger;
JAS|1|20|for the anger of man does not produce the righteousness that God requires.
JAS|1|21|Therefore put away all filthiness and rampant wickedness and receive with meekness the implanted word, which is able to save your souls.
JAS|1|22|But be doers of the word, and not hearers only, deceiving yourselves.
JAS|1|23|For if anyone is a hearer of the word and not a doer, he is like a man who looks intently at his natural face in a mirror.
JAS|1|24|For he looks at himself and goes away and at once forgets what he was like.
JAS|1|25|But the one who looks into the perfect law, the law of liberty, and perseveres, being no hearer who forgets but a doer who acts, he will be blessed in his doing.
JAS|1|26|If anyone thinks he is religious and does not bridle his tongue but deceives his heart, this person's religion is worthless.
JAS|1|27|Religion that is pure and undefiled before God and the Father is this: to visit orphans and widows in their affliction, and to keep oneself unstained from the world.
JAS|2|1|My brothers, show no partiality as you hold the faith in our Lord Jesus Christ, the Lord of glory.
JAS|2|2|For if a man wearing a gold ring and fine clothing comes into your assembly, and a poor man in shabby clothing also comes in,
JAS|2|3|and if you pay attention to the one who wears the fine clothing and say, "You sit here in a good place," while you say to the poor man, "You stand over there," or, "Sit down at my feet,"
JAS|2|4|have you not then made distinctions among yourselves and become judges with evil thoughts?
JAS|2|5|Listen, my beloved brothers, has not God chosen those who are poor in the world to be rich in faith and heirs of the kingdom, which he has promised to those who love him?
JAS|2|6|But you have dishonored the poor man. Are not the rich the ones who oppress you, and the ones who drag you into court?
JAS|2|7|Are they not the ones who blaspheme the honorable name by which you were called?
JAS|2|8|If you really fulfill the royal law according to the Scripture, "You shall love your neighbor as yourself," you are doing well.
JAS|2|9|But if you show partiality, you are committing sin and are convicted by the law as transgressors.
JAS|2|10|For whoever keeps the whole law but fails in one point has become accountable for all of it.
JAS|2|11|For he who said, "Do not commit adultery," also said, "Do not murder." If you do not commit adultery but do murder, you have become a transgressor of the law.
JAS|2|12|So speak and so act as those who are to be judged under the law of liberty.
JAS|2|13|For judgment is without mercy to one who has shown no mercy. Mercy triumphs over judgment.
JAS|2|14|What good is it, my brothers, if someone says he has faith but does not have works? Can that faith save him?
JAS|2|15|If a brother or sister is poorly clothed and lacking in daily food,
JAS|2|16|and one of you says to them, "Go in peace, be warmed and filled," without giving them the things needed for the body, what good is that?
JAS|2|17|So also faith by itself, if it does not have works, is dead.
JAS|2|18|But someone will say, "You have faith and I have works." Show me your faith apart from your works, and I will show you my faith by my works.
JAS|2|19|You believe that God is one; you do well. Even the demons believe- and shudder!
JAS|2|20|Do you want to be shown, you foolish person, that faith apart from works is useless?
JAS|2|21|Was not Abraham our father justified by works when he offered up his son Isaac on the altar?
JAS|2|22|You see that faith was active along with his works, and faith was completed by his works;
JAS|2|23|and the Scripture was fulfilled that says, "Abraham believed God, and it was counted to him as righteousness"- and he was called a friend of God.
JAS|2|24|You see that a person is justified by works and not by faith alone.
JAS|2|25|And in the same way was not also Rahab the prostitute justified by works when she received the messengers and sent them out by another way?
JAS|2|26|For as the body apart from the spirit is dead, so also faith apart from works is dead.
JAS|3|1|Not many of you should become teachers, my brothers, for you know that we who teach will be judged with greater strictness.
JAS|3|2|For we all stumble in many ways, and if anyone does not stumble in what he says, he is a perfect man, able also to bridle his whole body.
JAS|3|3|If we put bits into the mouths of horses so that they obey us, we guide their whole bodies as well.
JAS|3|4|Look at the ships also: though they are so large and are driven by strong winds, they are guided by a very small rudder wherever the will of the pilot directs.
JAS|3|5|So also the tongue is a small member, yet it boasts of great things. How great a forest is set ablaze by such a small fire!
JAS|3|6|And the tongue is a fire, a world of unrighteousness. The tongue is set among our members, staining the whole body, setting on fire the entire course of life, and set on fire by hell.
JAS|3|7|For every kind of beast and bird, of reptile and sea creature, can be tamed and has been tamed by mankind,
JAS|3|8|but no human being can tame the tongue. It is a restless evil, full of deadly poison.
JAS|3|9|With it we bless our Lord and Father, and with it we curse people who are made in the likeness of God.
JAS|3|10|From the same mouth come blessing and cursing. My brothers, these things ought not to be so.
JAS|3|11|Does a spring pour forth from the same opening both fresh and salt water?
JAS|3|12|Can a fig tree, my brothers, bear olives, or a grapevine produce figs? Neither can a salt pond yield fresh water.
JAS|3|13|Who is wise and understanding among you? By his good conduct let him show his works in the meekness of wisdom.
JAS|3|14|But if you have bitter jealousy and selfish ambition in your hearts, do not boast and be false to the truth.
JAS|3|15|This is not the wisdom that comes down from above, but is earthly, unspiritual, demonic.
JAS|3|16|For where jealousy and selfish ambition exist, there will be disorder and every vile practice.
JAS|3|17|But the wisdom from above is first pure, then peaceable, gentle, open to reason, full of mercy and good fruits, impartial and sincere.
JAS|3|18|And a harvest of righteousness is sown in peace by those who make peace.
JAS|4|1|What causes quarrels and what causes fights among you? Is it not this, that your passions are at war within you?
JAS|4|2|You desire and do not have, so you murder. You covet and cannot obtain, so you fight and quarrel. You do not have, because you do not ask.
JAS|4|3|You ask and do not receive, because you ask wrongly, to spend it on your passions.
JAS|4|4|You adulterous people! Do you not know that friendship with the world is enmity with God? Therefore whoever wishes to be a friend of the world makes himself an enemy of God.
JAS|4|5|Or do you suppose it is to no purpose that the Scripture says, "He yearns jealously over the spirit that he has made to dwell in us"?
JAS|4|6|But he gives more grace. Therefore it says, "God opposes the proud, but gives grace to the humble."
JAS|4|7|Submit yourselves therefore to God. Resist the devil, and he will flee from you.
JAS|4|8|Draw near to God, and he will draw near to you. Cleanse your hands, you sinners, and purify your hearts, you double-minded.
JAS|4|9|Be wretched and mourn and weep. Let your laughter be turned to mourning and your joy to gloom.
JAS|4|10|Humble yourselves before the Lord, and he will exalt you.
JAS|4|11|Do not speak evil against one another, brothers. The one who speaks against a brother or judges his brother, speaks evil against the law and judges the law. But if you judge the law, you are not a doer of the law but a judge.
JAS|4|12|There is only one lawgiver and judge, he who is able to save and to destroy. But who are you to judge your neighbor?
JAS|4|13|Come now, you who say, "Today or tomorrow we will go into such and such a town and spend a year there and trade and make a profit"-
JAS|4|14|yet you do not know what tomorrow will bring. What is your life? For you are a mist that appears for a little time and then vanishes.
JAS|4|15|Instead you ought to say, "If the Lord wills, we will live and do this or that."
JAS|4|16|As it is, you boast in your arrogance. All such boasting is evil.
JAS|4|17|So whoever knows the right thing to do and fails to do it, for him it is sin.
JAS|5|1|Come now, you rich, weep and howl for the miseries that are coming upon you.
JAS|5|2|Your riches have rotted and your garments are moth-eaten.
JAS|5|3|Your gold and silver have corroded, and their corrosion will be evidence against you and will eat your flesh like fire. You have laid up treasure in the last days.
JAS|5|4|Behold, the wages of the laborers who mowed your fields, which you kept back by fraud, are crying out against you, and the cries of the harvesters have reached the ears of the Lord of hosts.
JAS|5|5|You have lived on the earth in luxury and in self-indulgence. You have fattened your hearts in a day of slaughter.
JAS|5|6|You have condemned; you have murdered the righteous person. He does not resist you.
JAS|5|7|Be patient, therefore, brothers, until the coming of the Lord. See how the farmer waits for the precious fruit of the earth, being patient about it, until it receives the early and the late rains.
JAS|5|8|You also, be patient. Establish your hearts, for the coming of the Lord is at hand.
JAS|5|9|Do not grumble against one another, brothers, so that you may not be judged; behold, the Judge is standing at the door.
JAS|5|10|As an example of suffering and patience, brothers, take the prophets who spoke in the name of the Lord.
JAS|5|11|Behold, we consider those blessed who remained steadfast. You have heard of the steadfastness of Job, and you have seen the purpose of the Lord, how the Lord is compassionate and merciful.
JAS|5|12|But above all, my brothers, do not swear, either by heaven or by earth or by any other oath, but let your "yes" be yes and your "no" be no, so that you may not fall under condemnation.
JAS|5|13|Is anyone among you suffering? Let him pray. Is anyone cheerful? Let him sing praise.
JAS|5|14|Is anyone among you sick? Let him call for the elders of the church, and let them pray over him, anointing him with oil in the name of the Lord.
JAS|5|15|And the prayer of faith will save the one who is sick, and the Lord will raise him up. And if he has committed sins, he will be forgiven.
JAS|5|16|Therefore, confess your sins to one another and pray for one another, that you may be healed. The prayer of a righteous person has great power as it is working.
JAS|5|17|Elijah was a man with a nature like ours, and he prayed fervently that it might not rain, and for three years and six months it did not rain on the earth.
JAS|5|18|Then he prayed again, and heaven gave rain, and the earth bore its fruit.
JAS|5|19|My brothers, if anyone among you wanders from the truth and someone brings him back,
JAS|5|20|let him know that whoever brings back a sinner from his wandering will save his soul from death and will cover a multitude of sins.
