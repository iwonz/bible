1SAM|1|1|Был один человек из Рамафаим–Цофима, с горы Ефремовой, имя ему Елкана, сын Иерохама, сына Илия, сына Тоху, сына Цуфа, – Ефрафянин;
1SAM|1|2|у него были две жены: имя одной Анна, а имя другой Феннана; у Феннаны были дети, у Анны же не было детей.
1SAM|1|3|И ходил этот человек из города своего в положенные дни поклоняться и приносить жертву Господу Саваофу в Силом; там [были Илий и] два сына его, Офни и Финеес, священниками Господа.
1SAM|1|4|В тот день, когда Елкана приносил жертву, давал Феннане, жене своей, и всем сыновьям ее и дочерям ее части;
1SAM|1|5|Анне же давал часть особую, ибо любил Анну, хотя Господь заключил чрево ее.
1SAM|1|6|Соперница ее сильно огорчала ее, побуждая ее к ропоту на то, что Господь заключил чрево ее.
1SAM|1|7|Так бывало каждый год, когда ходила она в дом Господень; та огорчала ее, а эта плакала и не ела.
1SAM|1|8|И сказал ей Елкана, муж ее: Анна! что ты плачешь и почему не ешь, и отчего скорбит сердце твое? не лучше ли я для тебя десяти сыновей?
1SAM|1|9|И встала Анна после того, как они ели и пили в Силоме. Илий же священник сидел тогда на седалище у входа в храм Господень.
1SAM|1|10|И была она в скорби души, и молилась Господу, и горько плакала,
1SAM|1|11|и дала обет, говоря: Господи Саваоф! если Ты призришь на скорбь рабы Твоей и вспомнишь обо мне, и не забудешь рабы Твоей и дашь рабе Твоей дитя мужеского пола, то я отдам его Господу на все дни жизни его, и бритва не коснется головы его.
1SAM|1|12|Между тем как она долго молилась пред Господом, Илий смотрел на уста ее;
1SAM|1|13|и как Анна говорила в сердце своем, а уста ее только двигались, и не было слышно голоса ее, то Илий счел ее пьяною.
1SAM|1|14|И сказал ей Илий: доколе ты будешь пьяною? вытрезвись от вина твоего.
1SAM|1|15|И отвечала Анна, и сказала: нет, господин мой; я – жена, скорбящая духом, вина и сикера я не пила, но изливаю душу мою пред Господом;
1SAM|1|16|не считай рабы твоей негодною женщиною, ибо от великой печали моей и от скорби моей я говорила доселе.
1SAM|1|17|И отвечал Илий и сказал: иди с миром, и Бог Израилев исполнит прошение твое, чего ты просила у Него.
1SAM|1|18|Она же сказала: да найдет раба твоя милость в очах твоих! И пошла она в путь свой, и ела, и лице ее не было уже [печально], как прежде.
1SAM|1|19|И встали они поутру, и поклонились пред Господом, и возвратились, и пришли в дом свой в Раму. И познал Елкана Анну, жену свою, и вспомнил о ней Господь.
1SAM|1|20|Чрез несколько времени зачала Анна и родила сына и дала ему имя: Самуил, ибо, [говорила она], от Господа я испросила его.
1SAM|1|21|И пошел муж ее Елкана и все семейство его совершить годичную жертву Господу и обеты свои.
1SAM|1|22|Анна же не пошла, сказав мужу своему: когда младенец отнят будет от груди и подрастет, тогда я отведу его, и он явится пред Господом и останется там навсегда.
1SAM|1|23|И сказал ей Елкана, муж ее: делай, что тебе угодно; оставайся, доколе не вскормишь его грудью; только да утвердит Господь слово, [вышедшее из уст твоих]. И осталась жена [его], и кормила грудью сына своего, доколе не вскормила.
1SAM|1|24|Когда же вскормила его, пошла с ним в Силом, [взяв] три тельца и одну ефу муки и мех вина, и пришла в дом Господа в Силом; отрок же был еще дитя.
1SAM|1|25|и закололи тельца; и привела отрока к Илию
1SAM|1|26|и сказала: о, господин мой! да живет душа твоя, господин мой! я – та самая женщина, которая здесь при тебе стояла и молилась Господу;
1SAM|1|27|о сем дитяти молилась я, и исполнил мне Господь прошение мое, чего я просила у Него;
1SAM|1|28|и я отдаю его Господу на все дни жизни его, служить Господу. И поклонилась там Господу.
1SAM|2|1|И молилась Анна и говорила: возрадовалось сердце мое в Господе; вознесся рог мой в Боге моем; широко разверзлись уста мои на врагов моих, ибо я радуюсь о спасении Твоем.
1SAM|2|2|Нет [столь] святаго, как Господь; ибо нет другого, кроме Тебя; и нет твердыни, как Бог наш.
1SAM|2|3|Не умножайте речей надменных; дерзкие слова да не исходят из уст ваших; ибо Господь есть Бог ведения, и дела у Него взвешены.
1SAM|2|4|Лук сильных преломляется, а немощные препоясываются силою;
1SAM|2|5|сытые работают из хлеба, а голодные отдыхают; даже бесплодная рождает семь раз, а многочадная изнемогает.
1SAM|2|6|Господь умерщвляет и оживляет, низводит в преисподнюю и возводит;
1SAM|2|7|Господь делает нищим и обогащает, унижает и возвышает.
1SAM|2|8|Из праха подъемлет Он бедного, из брения возвышает нищего, посаждая с вельможами, и престол славы дает им в наследие; ибо у Господа основания земли, и Он утвердил на них вселенную.
1SAM|2|9|Стопы святых Своих Он блюдет, а беззаконные во тьме исчезают; ибо не силою крепок человек.
1SAM|2|10|Господь сотрет препирающихся с Ним; с небес возгремит на них. [Господь] будет судить концы земли, и даст крепость царю Своему и вознесет рог помазанника Своего.
1SAM|2|11|и пошел Елкана в Раму в дом свой, а отрок остался служить Господу при Илии священнике.
1SAM|2|12|Сыновья же Илия были люди негодные; они не знали Господа
1SAM|2|13|и долга священников в отношении к народу. Когда кто приносил жертву, отрок священнический, во время варения мяса, приходил с вилкой в руке своей
1SAM|2|14|и опускал ее в котел, или в кастрюлю, или на сковороду, или в горшок, и что вынет вилка, то брал себе священник. Так поступали они со всеми Израильтянами, приходившими туда в Силом.
1SAM|2|15|Даже прежде, нежели сожигали тук, приходил отрок священнический и говорил приносившему жертву: дай мяса на жаркое священнику; он не возьмет у тебя вареного мяса, а дай сырое.
1SAM|2|16|И [если] кто говорил ему: пусть сожгут прежде тук, как должно, и [потом] возьми себе, сколько пожелает душа твоя, то он говорил: нет, теперь же дай, а если нет, то силою возьму.
1SAM|2|17|И грех этих молодых людей был весьма велик пред Господом, ибо они отвращали от жертвоприношений Господу.
1SAM|2|18|Отрок же Самуил служил пред Господом, надевая льняной ефод.
1SAM|2|19|Верхнюю одежду малую делала ему мать его и приносила ему ежегодно, когда приходила с мужем своим для принесения положенной жертвы.
1SAM|2|20|И благословил Илий Елкану и жену его и сказал: да даст тебе Господь детей от жены сей вместо данного, которого ты отдал Господу! И пошли они в место свое.
1SAM|2|21|И посетил Господь Анну, и зачала она и родила еще трех сыновей и двух дочерей; а отрок Самуил возрастал у Господа.
1SAM|2|22|Илий же был весьма стар и слышал все, как поступают сыновья его со всеми Израильтянами, и что они спят с женщинами, собиравшимися у входа в скинию собрания.
1SAM|2|23|И сказал им: для чего вы делаете такие дела? ибо я слышу худые речи о вас от всего народа.
1SAM|2|24|Нет, дети мои, нехороша молва, которую я слышу: вы развращаете народ Господень;
1SAM|2|25|если согрешит человек против человека, то помолятся о нем Богу; если же человек согрешит против Господа, то кто будет ходатаем о нем? Но они не слушали голоса отца своего, ибо Господь решил уже предать их смерти.
1SAM|2|26|Отрок же Самуил более и более приходил в возраст и в благоволение у Господа и у людей.
1SAM|2|27|И пришел человек Божий к Илию и сказал ему: так говорит Господь: не открылся ли Я дому отца твоего, когда еще были они в Египте, в доме фараона?
1SAM|2|28|И не избрал ли его из всех колен Израилевых Себе во священника, чтоб он восходил к жертвеннику Моему, чтобы воскурял фимиам, чтобы носил ефод предо Мною? И не дал ли Я дому отца твоего от всех огнем сожигаемых жертв сынов Израилевых?
1SAM|2|29|Для чего же вы попираете ногами жертвы Мои и хлебные приношения Мои, которые заповедал Я для жилища [Моего], и для чего ты предпочитаешь Мне сыновей своих, утучняя себя начатками всех приношений народа Моего – Израиля?
1SAM|2|30|Посему так говорит Господь Бог Израилев: Я сказал [тогда]: "дом твой и дом отца твоего будут ходить пред лицем Моим вовек". Но теперь говорит Господь: да не будет так, ибо Я прославлю прославляющих Меня, а бесславящие Меня будут посрамлены.
1SAM|2|31|Вот, наступают дни, в [которые] Я подсеку мышцу твою и мышцу дома отца твоего, так что не будет старца в доме твоем;
1SAM|2|32|и ты будешь видеть бедствие жилища Моего, при всем том, что [Господь] благотворит Израилю и не будет в доме твоем старца во все дни,
1SAM|2|33|Я не отрешу у тебя [всех] от жертвенника Моего, чтобы томить глаза твои и мучить душу твою; но все потомство дома твоего будет умирать в средних летах.
1SAM|2|34|И вот тебе знамение, которое последует с двумя сыновьями твоими, Офни и Финеесом: оба они умрут в один день.
1SAM|2|35|И поставлю Себе священника верного; он будет поступать по сердцу Моему и по душе Моей; и дом его сделаю твердым, и он будет ходить пред помазанником Моим во все дни;
1SAM|2|36|и всякий, оставшийся из дома твоего, придет кланяться ему из–за геры серебра и куска хлеба и скажет: "причисли меня к какой–либо левитской должности, чтоб иметь пропитание".
1SAM|3|1|Отрок Самуил служил Господу при Илии; слово Господне было редко в те дни, видения [были] не часты.
1SAM|3|2|И было в то время, когда Илий лежал на своем месте, – глаза же его начали смежаться, и он не мог видеть, –
1SAM|3|3|и светильник Божий еще не погас, и Самуил лежал в храме Господнем, где ковчег Божий;
1SAM|3|4|воззвал Господь к Самуилу: И отвечал он: вот я!
1SAM|3|5|И побежал к Илию и сказал: вот я! ты звал меня. Но тот сказал: я не звал тебя; пойди назад, ложись. И он пошел и лег.
1SAM|3|6|Но Господь в другой раз воззвал к Самуилу: Он встал, и пришел к Илию вторично, и сказал: вот я! ты звал меня. Но тот сказал: я не звал тебя, сын мой; пойди назад, ложись.
1SAM|3|7|Самуил еще не знал тогда [голоса] Господа, и еще не открывалось ему слово Господне.
1SAM|3|8|И воззвал Господь к Самуилу еще в третий раз. Он встал и пришел к Илию и сказал: вот я! ты звал меня. Тогда понял Илий, что Господь зовет отрока.
1SAM|3|9|И сказал Илий Самуилу: пойди назад и ложись, и когда [Зовущий] позовет тебя, ты скажи: говори, Господи, ибо слышит раб Твой. И пошел Самуил и лег на месте своем.
1SAM|3|10|И пришел Господь, и стал, и воззвал, как в тот и другой раз: Самуил, Самуил! И сказал Самуил: говори, [Господи], ибо слышит раб Твой.
1SAM|3|11|И сказал Господь Самуилу: вот, Я сделаю дело в Израиле, о котором кто услышит, у того зазвенит в обоих ушах;
1SAM|3|12|в тот день Я исполню над Илием все то, что Я говорил о доме его; Я начну и окончу;
1SAM|3|13|Я объявил ему, что Я накажу дом его на веки за ту вину, что он знал, как сыновья его нечествуют, и не обуздывал их;
1SAM|3|14|и посему клянусь дому Илия, что вина дома Илиева не загладится ни жертвами, ни приношениями хлебными вовек.
1SAM|3|15|И спал Самуил до утра, и отворил двери дома Господня; и боялся Самуил объявить видение сие Илию.
1SAM|3|16|Но Илий позвал Самуила и сказал: сын мой Самуил! Тот сказал: вот я!
1SAM|3|17|И сказал [Илий]: что сказано тебе? не скрой от меня; то и то сделает с тобою Бог, и еще больше сделает, если ты утаишь от меня что–либо из всего того, что сказано тебе.
1SAM|3|18|И объявил ему Самуил все и не скрыл от него [ничего]. Тогда сказал [Илий]: Он – Господь; что Ему угодно, то да сотворит.
1SAM|3|19|И возрос Самуил, и Господь был с ним; и не осталось ни одного из слов его неисполнившимся.
1SAM|3|20|И узнал весь Израиль от Дана до Вирсавии, что Самуил удостоен быть пророком Господним.
1SAM|3|21|И продолжал Господь являться в Силоме после того, как открыл Себя Самуилу в Силоме чрез слово Господне.
1SAM|4|1|И было слово Самуила ко всему Израилю. И выступили Израильтяне против Филистимлян на войну и расположились станом при Авен–Езере, а Филистимляне расположились при Афеке.
1SAM|4|2|И выстроились Филистимляне против Израильтян, и произошла битва, и были поражены Израильтяне Филистимлянами, которые побили на поле сражения около четырех тысяч человек.
1SAM|4|3|И пришел народ в стан; и сказали старейшины Израилевы: за что поразил нас Господь сегодня пред Филистимлянами? возьмем себе из Силома ковчег завета Господня, и он пойдет среди нас и спасет нас от руки врагов наших.
1SAM|4|4|И послал народ в Силом, и принесли оттуда ковчег завета Господа Саваофа, седящего на херувимах; а при ковчеге завета Божия были и два сына Илиевы, Офни и Финеес.
1SAM|4|5|И когда прибыл ковчег завета Господня в стан, весь Израиль поднял такой сильный крик, что земля стонала.
1SAM|4|6|И услышали Филистимляне шум восклицаний и сказали: отчего такие громкие восклицания в стане Евреев? И узнали, что ковчег Господень прибыл в стан.
1SAM|4|7|И устрашились Филистимляне, ибо сказали: Бог тот пришел к ним в стан. И сказали: горе нам! ибо не бывало подобного ни вчера, ни третьего дня;
1SAM|4|8|горе нам! кто избавит нас от руки этого сильного Бога? Это – тот Бог, Который поразил Египтян всякими казнями в пустыне;
1SAM|4|9|укрепитесь и будьте мужественны, Филистимляне, чтобы вам не быть в порабощении у Евреев, как они у вас в порабощении; будьте мужественны и сразитесь с ними.
1SAM|4|10|И сразились Филистимляне, и поражены были Израильтяне, и каждый побежал в шатер свой, и было поражение весьма великое, и пало из Израильтян тридцать тысяч пеших.
1SAM|4|11|И ковчег Божий был взят, и два сына Илиевы, Офни и Финеес, умерли.
1SAM|4|12|И побежал один Вениамитянин с места сражения и пришел в Силом в тот же день; одежда на нем была разодрана и прах на голове его.
1SAM|4|13|Когда пришел он, Илий сидел на седалище при дороге у ворот и смотрел, ибо сердце его трепетало за ковчег Божий. И когда человек тот пришел и объявил в городе, то громко восстенал весь город.
1SAM|4|14|И услышал Илий звуки вопля и сказал: отчего такой шум? И тотчас подошел человек тот и объявил Илию.
1SAM|4|15|Илий был тогда девяноста восьми лет; и глаза его померкли, и он не мог видеть.
1SAM|4|16|И сказал тот человек Илию: я пришел из стана, сегодня же бежал я с места сражения. И сказал [Илий]: что произошло, сын мой?
1SAM|4|17|И отвечал вестник и сказал: побежал Израиль пред Филистимлянами, и поражение великое произошло в народе, и оба сына твои, Офни и Финеес, умерли, и ковчег Божий взят.
1SAM|4|18|Когда упомянул он о ковчеге Божием, [Илий] упал с седалища навзничь у ворот, сломал себе хребет и умер; ибо он [был] стар и тяжел. Был же он судьею Израиля сорок лет.
1SAM|4|19|Невестка его, жена Финеесова, была беременна уже пред родами. И когда услышала она известие о взятии ковчега Божия и о смерти свекра своего и мужа своего, то упала на колени и родила, ибо приступили к ней боли ее.
1SAM|4|20|И когда умирала она, стоявшие при ней женщины говорили ей: не бойся, ты родила сына. Но она не отвечала и не обращала внимания.
1SAM|4|21|И назвала младенца: Ихавод, сказав: "отошла слава от Израиля" – со взятием ковчега Божия и [со смертью] свекра ее и мужа ее.
1SAM|4|22|Она сказала: отошла слава от Израиля, ибо взят ковчег Божий.
1SAM|5|1|Филистимляне же взяли ковчег Божий и принесли его из Авен–Езера в Азот.
1SAM|5|2|И взяли Филистимляне ковчег Божий, и внесли его в храм Дагона, и поставили его подле Дагона.
1SAM|5|3|И встали Азотяне рано на другой день, и вот, Дагон лежит лицем своим к земле пред ковчегом Господним. И взяли они Дагона и опять поставили его на свое место.
1SAM|5|4|И встали они поутру на следующий день, и вот, Дагон лежит ниц на земле пред ковчегом Господним; голова Дагонова и обе руки его [лежали] отсеченные, каждая особо, на пороге, осталось только туловище Дагона.
1SAM|5|5|Посему жрецы Дагоновы и все приходящие в капище Дагона в Азот не ступают на порог Дагонов до сего дня.
1SAM|5|6|И отяготела рука Господня над Азотянами, и Он поражал их и наказал их мучительными наростами, в Азоте и в окрестностях его.
1SAM|5|7|И увидели это Азотяне и сказали: да не останется ковчег Бога Израилева у нас, ибо тяжка рука Его и для нас и для Дагона, бога нашего.
1SAM|5|8|И послали, и собрали к себе всех владетелей Филистимских, и сказали: что нам делать с ковчегом Бога Израилева? И сказали: пусть ковчег Бога Израилева перейдет в Геф. И отправили ковчег Бога Израилева в Геф.
1SAM|5|9|После того, как отправили его, была рука Господа на городе – ужас весьма великий, и поразил Господь жителей города от малого до большого, и показались на них наросты.
1SAM|5|10|И отослали они ковчег Божий в Аскалон; и когда пришел ковчег Божий в Аскалон, возопили Аскалонитяне, говоря: принесли к нам ковчег Бога Израилева, чтоб умертвить нас и народ наш.
1SAM|5|11|И послали, и собрали всех владетелей Филистимских, и сказали: отошлите ковчег Бога Израилева; пусть он возвратится в свое место, чтобы не умертвил он нас и народа нашего. Ибо смертельный ужас был во всем городе; весьма отяготела рука Божия на них.
1SAM|5|12|И те, которые не умерли, поражены были наростами, так что вопль города восходил до небес.
1SAM|6|1|И пробыл ковчег Господень в области Филистимской семь месяцев.
1SAM|6|2|И призвали Филистимляне жрецов и прорицателей, и сказали: что нам делать с ковчегом Господним? научите нас, как нам отпустить его в свое место.
1SAM|6|3|Те сказали: если вы хотите отпустить ковчег Бога Израилева, то не отпускайте его ни с чем, но принесите Ему жертву повинности; тогда исцелитесь и узнаете, за что не отступает от вас рука Его.
1SAM|6|4|И сказали они: какую жертву повинности должны мы принести Ему? Те сказали: по числу владетелей Филистимских пять наростов золотых и пять мышей золотых; ибо казнь одна на всех вас и на владетелях ваших;
1SAM|6|5|итак сделайте изваяния наростов ваших и изваяния мышей ваших, опустошающих землю, и воздайте славу Богу Израилеву; может быть, Он облегчит руку Свою над вами и над богами вашими и над землею вашею;
1SAM|6|6|и для чего вам ожесточать сердце ваше, как ожесточили сердце свое Египтяне и фараон? вот, когда Господь показал силу Свою над ними, то они отпустили их, и те пошли;
1SAM|6|7|итак возьмите, сделайте одну колесницу новую и возьмите двух первородивших коров, на которых не было ярма, и впрягите коров в колесницу, а телят их отведите от них домой;
1SAM|6|8|и возьмите ковчег Господень, и поставьте его на колесницу, а золотые вещи, которые принесете Ему в жертву повинности, положите в ящик сбоку его; и отпустите его, и пусть пойдет;
1SAM|6|9|и смотрите, если он пойдет к пределам своим, к Вефсамису, то он великое сие зло сделал нам; если же нет, то мы будем знать, что не его рука поразила нас, а сделалось это с нами случайно.
1SAM|6|10|И сделали они так: и взяли двух первородивших коров и впрягли их в колесницу, а телят их удержали дома;
1SAM|6|11|и поставили ковчег Господа на колесницу и ящик с золотыми мышами и изваяниями наростов.
1SAM|6|12|И пошли коровы прямо на дорогу к Вефсамису; одною дорогою шли, шли и мычали, но не уклонялись ни направо, ни налево; владетели же Филистимские следовали за ними до пределов Вефсамиса.
1SAM|6|13|[Жители] Вефсамиса жали тогда пшеницу в долине, и взглянув увидели ковчег Господень, и обрадовались, что увидели его.
1SAM|6|14|Колесница же пришла на поле Иисуса Вефсамитянина и остановилась там; и был тут большой камень, и раскололи колесницу на дрова, а коров принесли во всесожжение Господу.
1SAM|6|15|Левиты сняли ковчег Господа и ящик, бывший при нем, в котором [были] золотые вещи, и поставили на большом том камне; жители же Вефсамиса принесли в тот день всесожжения и закололи жертвы Господу.
1SAM|6|16|И пять владетелей Филистимских видели [это] и возвратились в тот день в Аккарон.
1SAM|6|17|Золотые эти наросты, которые принесли Филистимляне в жертву повинности Господу, были: один за Азот, один за Газу, один за Аскалон, один за Геф, один за Аккарон;
1SAM|6|18|а золотые мыши [были] по числу всех городов Филистимских – пяти владетелей, от городов укрепленных и до открытых сел, до большого камня, на котором поставили ковчег Господа и [который находится] до сего дня на поле Иисуса Вефсамитянина.
1SAM|6|19|И поразил Он жителей Вефсамиса за то, что они заглядывали в ковчег Господа, и убил из народа пятьдесят тысяч семьдесят человек; и заплакал народ, ибо поразил Господь народ поражением великим.
1SAM|6|20|И сказали жители Вефсамиса: кто может стоять пред Господом, сим святым Богом? и к кому Он пойдет от нас?
1SAM|6|21|И послали послов к жителям Кириаф–Иарима сказать: Филистимляне возвратили ковчег Господа; придите, возьмите его к себе.
1SAM|7|1|И пришли жители Кириаф–Иарима, и взяли ковчег Господа, и принесли его в дом Аминадава, на холм, а Елеазара, сына его, посвятили, чтобы он хранил ковчег Господа.
1SAM|7|2|С того дня, как остался ковчег в Кириаф–Иариме, прошло много времени, лет двадцать. И обратился весь дом Израилев к Господу.
1SAM|7|3|И сказал Самуил всему дому Израилеву, говоря: если вы всем сердцем своим обращаетесь к Господу, то удалите из среды себя богов иноземных и Астарт и расположите сердце ваше к Господу, и служите Ему одному, и Он избавит вас от руки Филистимлян.
1SAM|7|4|И удалили сыны Израилевы Ваалов и Астарт и стали служить одному Господу.
1SAM|7|5|И сказал Самуил: соберите всех Израильтян в Массифу и я помолюсь о вас Господу.
1SAM|7|6|И собрались в Массифу, и черпали воду, и проливали пред Господом, и постились в тот день, говоря: согрешили мы пред Господом. И судил Самуил сынов Израилевых в Массифе.
1SAM|7|7|Когда же услышали Филистимляне, что собрались сыны Израилевы в Массифу, тогда пошли владетели Филистимские на Израиля. Израильтяне, услышав [о том], убоялись Филистимлян.
1SAM|7|8|И сказали сыны Израилевы Самуилу: не переставай взывать о нас к Господу Богу нашему, чтоб он спас нас от руки Филистимлян.
1SAM|7|9|И взял Самуил одного ягненка от сосцов, и принес его во всесожжение Господу, и воззвал Самуил к Господу о Израиле, и услышал его Господь.
1SAM|7|10|И когда Самуил возносил всесожжение, Филистимляне пришли воевать с Израилем. Но Господь возгремел в тот день сильным громом над Филистимлянами и навел на них ужас, и они были поражены пред Израилем.
1SAM|7|11|И выступили Израильтяне из Массифы, и преследовали Филистимлян, и поражали их до места под Вефхором.
1SAM|7|12|И взял Самуил один камень, и поставил между Массифою и между Сеном, и назвал его Авен–Езер, сказав: до сего места помог нам Господь.
1SAM|7|13|Так усмирены были Филистимляне, и не стали более ходить в пределы Израилевы; и была рука Господня на Филистимлянах во все дни Самуила.
1SAM|7|14|И возвращены были Израилю города, которые взяли Филистимляне у Израиля, от Аккарона и до Гефа, и пределы их освободил Израиль из рук Филистимлян, и был мир между Израилем и Аморреями.
1SAM|7|15|И был Самуил судьею Израиля во все дни жизни своей:
1SAM|7|16|из года в год он ходил и обходил Вефиль, и Галгал и Массифу и судил Израиля во всех сих местах;
1SAM|7|17|потом возвращался в Раму; ибо [там] был дом его, и там судил он Израиля, и построил там жертвенник Господу.
1SAM|8|1|Когда же состарился Самуил, то поставил сыновей своих судьями над Израилем.
1SAM|8|2|Имя старшему сыну его Иоиль, а имя второму [сыну] его Авия; они [были] судьями в Вирсавии.
1SAM|8|3|Но сыновья его не ходили путями его, а уклонились в корысть и брали подарки, и судили превратно.
1SAM|8|4|И собрались все старейшины Израиля, и пришли к Самуилу в Раму,
1SAM|8|5|и сказали ему: вот, ты состарился, а сыновья твои не ходят путями твоими; итак поставь над нами царя, чтобы он судил нас, как у прочих народов.
1SAM|8|6|И не понравилось слово сие Самуилу, когда они сказали: дай нам царя, чтобы он судил нас. И молился Самуил Господу.
1SAM|8|7|И сказал Господь Самуилу: послушай голоса народа во всем, что они говорят тебе; ибо не тебя они отвергли, но отвергли Меня, чтоб Я не царствовал над ними;
1SAM|8|8|как они поступали с того дня, в который Я вывел их из Египта, и до сего дня, оставляли Меня и служили иным богам, так поступают они с тобою;
1SAM|8|9|итак послушай голоса их; только представь им и объяви им права царя, который будет царствовать над ними.
1SAM|8|10|И пересказал Самуил все слова Господа народу, просящему у него царя,
1SAM|8|11|и сказал: вот какие будут права царя, который будет царствовать над вами: сыновей ваших он возьмет и приставит их к колесницам своим и [сделает] всадниками своими, и будут они бегать пред колесницами его;
1SAM|8|12|и поставит [их] у себя тысяченачальниками и пятидесятниками, и чтобы они возделывали поля его, и жали хлеб его, и делали ему воинское оружие и колесничный прибор его;
1SAM|8|13|и дочерей ваших возьмет, чтоб они составляли масти, варили кушанье и пекли хлебы;
1SAM|8|14|и поля ваши и виноградные и масличные сады ваши лучшие возьмет, и отдаст слугам своим;
1SAM|8|15|и от посевов ваших и из виноградных садов ваших возьмет десятую часть и отдаст евнухам своим и слугам своим;
1SAM|8|16|и рабов ваших и рабынь ваших, и юношей ваших лучших, и ослов ваших возьмет и употребит на свои дела;
1SAM|8|17|от мелкого скота вашего возьмет десятую часть, и сами вы будете ему рабами;
1SAM|8|18|и восстенаете тогда от царя вашего, которого вы избрали себе; и не будет Господь отвечать вам тогда.
1SAM|8|19|Но народ не согласился послушаться голоса Самуила, и сказал: нет, пусть царь будет над нами,
1SAM|8|20|и мы будем как прочие народы: будет судить нас царь наш, и ходить пред нами, и вести войны наши.
1SAM|8|21|И выслушал Самуил все слова народа, и пересказал их вслух Господа.
1SAM|8|22|И сказал Господь Самуилу: послушай голоса их и поставь им царя. И сказал Самуил Израильтянам: пойдите каждый в свой город.
1SAM|9|1|Был некто из сынов Вениамина, имя его Кис, сын Авиила, сына Церона, сына Бехорафа, сына Афия, сына некоего Вениамитянина, человек знатный.
1SAM|9|2|У него был сын, имя его Саул, молодой и красивый; и не было никого из Израильтян красивее его; он от плеч своих был выше всего народа.
1SAM|9|3|И пропали ослицы у Киса, отца Саулова, и сказал Кис Саулу, сыну своему: возьми с собою одного из слуг и встань, пойди, поищи ослиц.
1SAM|9|4|И прошел он гору Ефремову и прошел землю Шалишу, но не нашли; и прошли землю Шаалим, и [там их] нет; и прошел он землю Вениаминову, и не нашли.
1SAM|9|5|Когда они пришли в землю Цуф, Саул сказал слуге своему, который был с ним: пойдем назад, чтобы отец мой, оставив ослиц, не стал беспокоиться о нас.
1SAM|9|6|Но слуга сказал ему: вот в этом городе есть человек Божий, человек уважаемый; все, что он ни скажет, сбывается; сходим теперь туда; может быть, он укажет нам путь наш, по которому нам идти.
1SAM|9|7|И сказал Саул слуге своему: вот мы пойдем, а что мы принесем тому человеку? ибо хлеба не стало в сумах наших, и подарка нет, чтобы поднести человеку Божию; что у нас?
1SAM|9|8|И опять отвечал слуга Саулу и сказал: вот в руке моей четверть сикля серебра; я отдам человеку Божию, и он укажет нам путь наш.
1SAM|9|9|Прежде у Израиля, когда кто–нибудь шел вопрошать Бога, говорили так: "пойдем к прозорливцу"; ибо тот, кого [называют] ныне пророком, прежде назывался прозорливцем.
1SAM|9|10|И сказал Саул слуге своему: хорошо ты говоришь; пойдем. И пошли в город, где человек Божий.
1SAM|9|11|Когда они поднимались вверх в город, то встретили девиц, вышедших черпать воду, и сказали им: есть ли здесь прозорливец?
1SAM|9|12|Те отвечали им и сказали: есть; вот, он впереди тебя; только поспешай, ибо он сегодня пришел в город, потому что сегодня у народа жертвоприношение на высоте;
1SAM|9|13|когда придете в город, застанете его, пока он еще не пошел на ту высоту, на обед; ибо народ не начнет есть, доколе он не придет; потому что он благословит жертву, и после того станут есть званые; итак ступайте, теперь еще застанете его.
1SAM|9|14|И пошли они в город. Когда же вошли в средину города, то вот и Самуил выходит навстречу им, чтоб идти на высоту.
1SAM|9|15|А Господь открыл Самуилу за день до прихода Саулова и сказал:
1SAM|9|16|завтра в это время Я пришлю к тебе человека из земли Вениаминовой, и ты помажь его в правителя народу Моему – Израилю, и он спасет народ Мой от руки Филистимлян; ибо Я призрел на народ Мой, так как вопль его достиг до Меня.
1SAM|9|17|Когда Самуил увидел Саула, то Господь сказал ему: вот человек, о котором Я говорил тебе; он будет управлять народом Моим.
1SAM|9|18|И подошел Саул к Самуилу в воротах и спросил его: скажи мне, где дом прозорливца?
1SAM|9|19|И отвечал Самуил Саулу, и сказал: я прозорливец, иди впереди меня на высоту; и вы будете обедать со мною сегодня, и отпущу тебя утром, и все, что у тебя на сердце, скажу тебе;
1SAM|9|20|а об ослицах, которые у тебя пропали уже три дня, не заботься; они нашлись. И кому все вожделенное в Израиле? Не тебе ли и всему дому отца твоего?
1SAM|9|21|И отвечал Саул и сказал: не сын ли я Вениамина, одного из меньших колен Израилевых? И племя мое не малейшее ли между всеми племенами колена Вениаминова? К чему же ты говоришь мне это?
1SAM|9|22|И взял Самуил Саула и слугу его, и ввел их в комнату, и дал им первое место между званными, которых было около тридцати человек.
1SAM|9|23|И сказал Самуил повару: подай ту часть, которую я дал тебе и о которой я сказал тебе: "отложи ее у себя".
1SAM|9|24|И взял повар плечо и что было при нем и положил пред Саулом. И сказал [Самуил]: вот это оставлено, положи пред собою [и] ешь, ибо к сему времени сбережено [это] для тебя, когда я созывал народ. И обедал Саул с Самуилом в тот день.
1SAM|9|25|И сошли они с высоты в город, и Самуил разговаривал с Саулом на кровле.
1SAM|9|26|Утром встали они так: когда взошла заря, Самуил воззвал к Саулу на кровлю и сказал: встань, я провожу тебя. И встал Саул, и вышли оба они из дома, он и Самуил.
1SAM|9|27|Когда подходили они к концу города, Самуил сказал Саулу: скажи слуге, чтобы он пошел впереди нас, – и он пошел вперед; – а ты остановись теперь, и я открою тебе, что сказал Бог.
1SAM|10|1|И взял Самуил сосуд с елеем и вылил на голову его, и поцеловал его и сказал: вот, Господь помазывает тебя в правителя наследия Своего:
1SAM|10|2|когда ты теперь пойдешь от меня, то встретишь двух человек близ гроба Рахили, на пределах Вениаминовых, в Целцахе, и они скажут тебе: "нашлись ослицы, которых ты ходил искать, и вот отец твой, забыв об ослицах, беспокоится о вас, говоря: что с сыном моим?"
1SAM|10|3|И пойдешь оттуда далее и придешь к дубраве Фаворской, и встретят тебя там три человека, идущих к Богу в Вефиль: один несет трех козлят, другой несет три хлеба, а третий несет мех с вином;
1SAM|10|4|и будут приветствовать они тебя и дадут тебе два хлеба, и ты возьмешь из рук их.
1SAM|10|5|После того ты придешь на холм Божий, где охранный отряд Филистимский; и когда войдешь там в город, встретишь сонм пророков, сходящих с высоты, и пред ними псалтирь и тимпан, и свирель и гусли, и они пророчествуют;
1SAM|10|6|и найдет на тебя Дух Господень, и ты будешь пророчествовать с ними и сделаешься иным человеком.
1SAM|10|7|Когда эти знамения сбудутся с тобою, тогда делай, что может рука твоя, ибо с тобою Бог.
1SAM|10|8|И ты пойди прежде меня в Галгал, куда и я приду к тебе для принесения всесожжений и мирных жертв; семь дней жди, доколе я не приду к тебе, и тогда укажу тебе, что тебе делать.
1SAM|10|9|Как скоро Саул обратился, чтоб идти от Самуила, Бог дал ему иное сердце, и сбылись все те знамения в тот же день.
1SAM|10|10|Когда пришли они к холму, вот встречается им сонм пророков, и сошел на него Дух Божий, и он пророчествовал среди них.
1SAM|10|11|Все знавшие его вчера и третьего дня, увидев, что он с пророками пророчествует, говорили в народе друг другу: что это сталось с сыном Кисовым? неужели и Саул во пророках?
1SAM|10|12|И отвечал один из бывших там и сказал: а у тех кто отец? Посему вошло в пословицу: "неужели и Саул во пророках?"
1SAM|10|13|И перестал он пророчествовать, и пошел на высоту.
1SAM|10|14|И сказал дядя Саулов ему и слуге его: куда вы ходили? Он сказал: искать ослиц, но, видя, что [их] нет, зашли к Самуилу.
1SAM|10|15|И сказал дядя Саулов: расскажи мне, что сказал вам Самуил.
1SAM|10|16|И сказал Саул дяде своему: он объявил нам, что ослицы нашлись. А того, что сказал ему Самуил о царстве, не открыл ему.
1SAM|10|17|И созвал Самуил народ к Господу в Массифу
1SAM|10|18|и сказал сынам Израилевым: так говорит Господь Бог Израилев: Я вывел Израиля из Египта и избавил вас от руки Египтян и от руки всех царств, угнетавших вас.
1SAM|10|19|А вы теперь отвергли Бога вашего, Который спасает вас от всех бедствий ваших и скорбей ваших, и сказали Ему: "царя поставь над нами". Итак предстаньте теперь пред Господом по коленам вашим и по племенам вашим.
1SAM|10|20|И велел Самуил подходить всем коленам Израилевым, и указано колено Вениаминово.
1SAM|10|21|И велел подходить колену Вениаминову по племенам его, и указано племя Матриево; и приводят племя Матриево по мужам, и назван Саул, сын Кисов; и искали его, и не находили.
1SAM|10|22|И вопросили еще Господа: придет ли еще он сюда? И сказал Господь: вот он скрывается в обозе.
1SAM|10|23|И побежали и взяли его оттуда, и он стал среди народа и был от плеч своих выше всего народа.
1SAM|10|24|И сказал Самуил всему народу: видите ли, кого избрал Господь? подобного ему нет во всем народе. Тогда весь народ воскликнул и сказал: да живет царь!
1SAM|10|25|И изложил Самуил народу права царства, и написал в книгу, и положил пред Господом. И отпустил весь народ, каждого в дом свой.
1SAM|10|26|Также и Саул пошел в дом свой, в Гиву; и пошли с ним храбрые, которых сердца коснулся Бог.
1SAM|10|27|А негодные люди говорили: ему ли спасать нас? И презрели его и не поднесли ему даров; но он как бы не замечал того.
1SAM|11|1|И пришел Наас Аммонитянин и осадил Иавис Галаадский. И сказали все жители Иависа Наасу: заключи с нами союз, и мы будем служить тебе.
1SAM|11|2|И сказал им Наас Аммонитянин: я заключу с вами союз, но с тем, чтобы выколоть у каждого из вас правый глаз и тем положить бесчестие на всего Израиля.
1SAM|11|3|И сказали ему старейшины Иависа: дай нам сроку семь дней, чтобы послать нам послов во все пределы Израильские, и если никто не поможет нам, то мы выйдем к тебе.
1SAM|11|4|И пришли послы в Гиву Саулову и пересказали слова сии вслух народа; и весь народ поднял вопль и заплакал.
1SAM|11|5|И вот, пришел Саул позади волов с поля и сказал: что [сделалось] с народом, что он плачет? И пересказали ему слова жителей Иависа.
1SAM|11|6|И сошел Дух Божий на Саула, когда он услышал слова сии, и сильно воспламенился гнев его;
1SAM|11|7|и взял он пару волов, и рассек их на части, и послал во все пределы Израильские чрез тех послов, объявляя, что так будет поступлено с волами того, кто не пойдет вслед Саула и Самуила. И напал страх Господень на народ, и выступили [все], как один человек.
1SAM|11|8|[Саул] осмотрел их в Везеке, и нашлось сынов Израилевых триста тысяч и мужей Иудиных тридцать тысяч.
1SAM|11|9|И сказали пришедшим послам: так скажите жителям Иависа Галаадского: завтра будет к вам помощь, когда обогреет солнце. И пришли послы и объявили жителям Иависа, и они обрадовались.
1SAM|11|10|И сказали жители Иависа [Наасу]: завтра выйдем к вам, и поступайте с нами, как вам угодно.
1SAM|11|11|В следующий день Саул разделил народ на три отряда, и они проникли в средину стана во время утренней стражи и поразили Аммонитян до дневного зноя; оставшиеся рассеялись, так что не осталось из них двоих вместе.
1SAM|11|12|Тогда сказал народ Самуилу: кто говорил: "Саулу ли царствовать над нами"? дайте этих людей, и мы умертвим их.
1SAM|11|13|Но Саул сказал: в сей день никого не должно умерщвлять, ибо сегодня Господь совершил спасение в Израиле.
1SAM|11|14|И сказал Самуил народу: пойдем в Галгал, и обновим там царство.
1SAM|11|15|И пошел весь народ в Галгал, и поставили там Саула царем пред Господом в Галгале, и принесли там мирные жертвы пред Господом. И весьма веселились там Саул и все Израильтяне.
1SAM|12|1|И сказал Самуил всему Израилю: вот, я послушался голоса вашего во всем, что вы говорили мне, и поставил над вами царя,
1SAM|12|2|и вот, царь ходит пред вами; а я состарился и поседел; и сыновья мои с вами; я же ходил пред вами от юности моей и до сего дня;
1SAM|12|3|вот я; свидетельствуйте на меня пред Господом и пред помазанником Его, у кого взял я вола, у кого взял осла, кого обидел и кого притеснил, у кого взял дар и закрыл в [деле] его глаза мои, – и я возвращу вам.
1SAM|12|4|И отвечали: ты не обижал нас и не притеснял нас и ничего ни у кого не взял.
1SAM|12|5|И сказал он им: свидетель на вас Господь, и свидетель помазанник Его в сей день, что вы не нашли ничего за мною. И сказали: свидетель.
1SAM|12|6|Тогда Самуил сказал народу: [свидетель] Господь, Который поставил Моисея и Аарона и Который вывел отцов ваших из земли Египетской.
1SAM|12|7|Теперь же предстаньте, и я буду судиться с вами пред Господом о всех благодеяниях, которые оказал Он вам и отцам вашим.
1SAM|12|8|Когда пришел Иаков в Египет, и отцы ваши возопили к Господу, то Господь послал Моисея и Аарона, и они вывели отцов ваших из Египта и поселили их на месте сем.
1SAM|12|9|Но они забыли Господа Бога своего, и Он предал их в руки Сисары, военачальника Асорского, и в руки Филистимлян и в руки царя Моавитского, [которые] воевали против них.
1SAM|12|10|Но когда они возопили к Господу и сказали: "согрешили мы, ибо оставили Господа и стали служить Ваалам и Астартам, теперь избавь нас от руки врагов наших, и мы будем служить Тебе",
1SAM|12|11|тогда Господь послал Иероваала, и Варака, и Иеффая, и Самуила, и избавил вас от руки врагов ваших, окружавших вас, и вы жили безопасно.
1SAM|12|12|Но увидев, что Наас, царь Аммонитский, идет против вас, вы сказали мне: "нет, царь пусть царствует над нами", тогда как Господь Бог ваш – Царь ваш.
1SAM|12|13|Итак, вот царь, которого вы избрали, которого вы требовали: вот, Господь поставил над вами царя.
1SAM|12|14|Если будете бояться Господа и служить Ему и слушать гласа Его, и не станете противиться повелениям Господа, и будете и вы и царь ваш, который царствует над вами, [ходить] вслед Господа, Бога вашего.
1SAM|12|15|а если не будете слушать гласа Господа и станете противиться повелениям Господа, то рука Господа будет против вас, [как была] против отцов ваших.
1SAM|12|16|Теперь станьте и посмотрите на дело великое, которое Господь совершит пред глазами вашими:
1SAM|12|17|не жатва ли пшеницы ныне? Но я воззову к Господу, и пошлет Он гром и дождь, и вы узнаете и увидите, как велик грех, который вы сделали пред очами Господа, прося себе царя.
1SAM|12|18|И воззвал Самуил к Господу, и Господь послал гром и дождь в тот день; и пришел весь народ в большой страх от Господа и Самуила.
1SAM|12|19|И сказал весь народ Самуилу: помолись о рабах твоих пред Господом Богом твоим, чтобы не умереть нам; ибо ко всем грехам нашим мы прибавили еще грех, когда просили себе царя.
1SAM|12|20|И отвечал Самуил народу: не бойтесь, грех этот вами сделан, но вы не отступайте только от Господа и служите Господу всем сердцем вашим
1SAM|12|21|и не обращайтесь вслед ничтожных [богов], которые не принесут пользы и не избавят; ибо они – ничто;
1SAM|12|22|Господь же не оставит народа Своего ради великого имени Своего, ибо Господу угодно было избрать вас народом Своим;
1SAM|12|23|и я также не допущу себе греха пред Господом, чтобы перестать молиться за вас, и буду наставлять вас на путь добрый и прямой;
1SAM|12|24|только бойтесь Господа и служите Ему истинно, от всего сердца вашего, ибо вы видели, какие великие дела Он сделал с вами;
1SAM|12|25|если же вы будете делать зло, то и вы и царь ваш погибнете.
1SAM|13|1|Год был по воцарении Саула, и другой год царствовал он над Израилем, как выбрал Саул себе три тысячи из Израильтян:
1SAM|13|2|две тысячи были с Саулом в Михмасе и на горе Вефильской, тысяча же была с Ионафаном в Гиве Вениаминовой; а прочий народ отпустил он по домам своим.
1SAM|13|3|И разбил Ионафан охранный отряд Филистимский, который был в Гиве; и услышали об этом Филистимляне, а Саул протрубил трубою по всей стране, возглашая: да услышат Евреи!
1SAM|13|4|Когда весь Израиль услышал, что разбил Саул охранный отряд Филистимский и что Израиль сделался ненавистным для Филистимлян, то народ собрался к Саулу в Галгал.
1SAM|13|5|И собрались Филистимляне на войну против Израиля: тридцать тысяч колесниц и шесть тысяч конницы, и народа множество, как песок на берегу моря; и пришли и расположились станом в Михмасе, с восточной стороны Беф–Авена.
1SAM|13|6|Израильтяне, видя, что они в опасности, потому что народ был стеснен, укрывались в пещерах и в ущельях, и между скалами, и в башнях, и во рвах;
1SAM|13|7|а [некоторые] из Евреев переправились за Иордан в страну Гадову и Галаадскую; Саул же находился еще в Галгале, и весь народ, бывший с ним, находился в страхе.
1SAM|13|8|И ждал он семь дней, до срока, [назначенного] Самуилом, а Самуил не приходил в Галгал; и стал народ разбегаться от него.
1SAM|13|9|И сказал Саул: приведите ко мне, что [назначено] для жертвы всесожжения и для жертв мирных. И вознес всесожжение.
1SAM|13|10|Но едва кончил он возношение всесожжения, вот, приходит Самуил; и вышел Саул к нему навстречу, чтобы приветствовать его.
1SAM|13|11|Но Самуил сказал: что ты сделал? Саул отвечал: я видел, что народ разбегается от меня, а ты не приходил к назначенному времени; Филистимляне же собрались в Михмасе;
1SAM|13|12|тогда подумал я: "теперь придут на меня Филистимляне в Галгал, а я еще не вопросил Господа", и потому решился принести всесожжение.
1SAM|13|13|И сказал Самуил Саулу: худо поступил ты, что не исполнил повеления Господа Бога твоего, которое дано было тебе, ибо ныне упрочил бы Господь царствование твое над Израилем навсегда;
1SAM|13|14|но теперь не устоять царствованию твоему; Господь найдет Себе мужа по сердцу Своему, и повелит ему Господь быть вождем народа Своего, так как ты не исполнил того, что было повелено тебе Господом.
1SAM|13|15|И встал Самуил и пошел из Галгала в Гиву Вениаминову; а Саул пересчитал людей, бывших с ним, до шестисот человек.
1SAM|13|16|Саул с сыном своим Ионафаном и людьми, находившимися при них, засели в Гиве Вениаминовой; Филистимляне же стояли станом в Михмасе.
1SAM|13|17|И вышли из стана Филистимского три отряда для опустошения земли: один направился по дороге к Офре, в округ Суаль,
1SAM|13|18|другой отряд направился по дороге Вефоронской, а третий направился по дороге к границе долины Цевоим, к пустыне.
1SAM|13|19|Кузнецов не было во всей земле Израильской; ибо Филистимляне опасались, чтобы Евреи не сделали меча или копья.
1SAM|13|20|И должны были ходить все Израильтяне к Филистимлянам оттачивать свои сошники, и свои заступы, и свои топоры, и свои кирки,
1SAM|13|21|когда сделается щербина на острие у сошников, и у заступов, и у вил, и у топоров, или нужно рожон поправить.
1SAM|13|22|Поэтому во время войны не было ни меча, ни копья у всего народа, бывшего с Саулом и Ионафаном, а [только] нашлись они у Саула и Ионафана, сына его.
1SAM|13|23|И вышел передовой отряд Филистимский к переправе Михмасской.
1SAM|14|1|В один день сказал Ионафан, сын Саулов, слуге оруженосцу своему: ступай, перейдем к отряду Филистимскому, что на той стороне. А отцу своему не сказал [об этом].
1SAM|14|2|Саул же находился в окраине Гивы, под гранатовым деревом, что в Мигроне. С ним было около шестисот человек народа
1SAM|14|3|и Ахия, сын Ахитува, брата Иохаведа, сына Финееса, сына Илия, священник Господа в Силоме, носивший ефод. Народ же не знал, что Ионафан пошел.
1SAM|14|4|Между переходами, по которым Ионафан искал пробраться к отряду Филистимскому, была острая скала с одной стороны и острая скала с другой: имя одной Боцец, а имя другой Сене;
1SAM|14|5|одна скала выдавалась с севера к Михмасу, другая с юга к Гиве.
1SAM|14|6|И сказал Ионафан слуге оруженосцу своему: ступай, перейдем к отряду этих необрезанных; может быть, Господь поможет нам, ибо для Господа нетрудно спасти чрез многих, или немногих.
1SAM|14|7|И отвечал оруженосец: делай все, что на сердце у тебя; иди, вот я с тобою, куда тебе угодно.
1SAM|14|8|И сказал Ионафан: вот, мы перейдем к этим людям и станем на виду у них;
1SAM|14|9|если они так скажут нам: "остановитесь, пока мы подойдем к вам", то мы остановимся на своих местах и не взойдем к ним;
1SAM|14|10|а если так скажут: "поднимитесь к нам", то мы взойдем, ибо Господь предал их в руки наши; и это будет знаком для нас.
1SAM|14|11|Когда оба они стали на виду у отряда Филистимского, то Филистимляне сказали: вот, Евреи выходят из ущелий, в которых попрятались они.
1SAM|14|12|И закричали люди, составлявшие отряд, к Ионафану и оруженосцу его, говоря: взойдите к нам, и мы вам скажем нечто. Тогда Ионафан сказал оруженосцу своему: следуй за мною, ибо Господь предал их в руки Израиля.
1SAM|14|13|И начал всходить Ионафан, [цепляясь] руками и ногами, и оруженосец его за ним. И падали [Филистимляне] пред Ионафаном, а оруженосец добивал их за ним.
1SAM|14|14|И пало от этого первого поражения, нанесенного Ионафаном и оруженосцем его, около двадцати человек, на половине поля, обрабатываемого парою волов в день.
1SAM|14|15|И произошел ужас в стане на поле и во всем народе; передовые отряды и опустошавшие землю пришли в трепет; дрогнула вся земля, и был ужас великий от Господа.
1SAM|14|16|И увидели стражи Саула в Гиве Вениаминовой, что толпа рассеивается и бежит туда и сюда.
1SAM|14|17|И сказал Саул к народу, бывшему с ним; пересмотрите и узнайте, кто из наших вышел. И пересмотрели, и вот нет Ионафана и оруженосца его.
1SAM|14|18|И сказал Саул Ахии: "принеси кивот Божий", ибо кивот Божий в то время был с сынами Израильскими.
1SAM|14|19|Саул еще говорил к священнику, как смятение в стане Филистимском более и более [распространялось и] увеличивалось. Тогда сказал Саул священнику: сложи руки твои.
1SAM|14|20|И воскликнул Саул и весь народ, бывший с ним, и пришли к месту сражения, и вот, там меч каждого [обращен] был против ближнего своего; смятение [было] очень великое.
1SAM|14|21|Тогда и Евреи, которые вчера и третьего дня были у Филистимлян и которые повсюду ходили с ними в стане, пристали к Израильтянам, находившимся с Саулом и Ионафаном;
1SAM|14|22|и все Израильтяне, скрывавшиеся в горе Ефремовой, услышав, что Филистимляне побежали, также пристали к своим в сражении.
1SAM|14|23|И спас Господь в тот день Израиля; битва же простерлась даже до Беф–Авена.
1SAM|14|24|Люди Израильские были истомлены в тот день; а Саул заклял народ, сказав: проклят, кто вкусит хлеба до вечера, доколе я не отомщу врагам моим. И никто из народа не вкусил пищи.
1SAM|14|25|И пошел весь народ в лес, и был там на поляне мед.
1SAM|14|26|И вошел народ в лес, говоря: вот, течет мед. Но никто не протянул руки своей ко рту своему, ибо народ боялся заклятия.
1SAM|14|27|Ионафан же не слышал, когда отец его заклинал народ, и, протянув конец палки, которая была в руке его, обмокнул ее в сот медовый и обратил рукою к устам своим, и просветлели глаза его.
1SAM|14|28|И сказал ему один из народа, говоря: отец твой заклял народ, сказав: "проклят, кто сегодня вкусит пищи"; от этого народ истомился.
1SAM|14|29|И сказал Ионафан: смутил отец мой землю; смотрите, у меня просветлели глаза, когда я вкусил немного этого меду;
1SAM|14|30|если бы поел сегодня народ из добычи, какую нашел у врагов своих, то не большее ли было бы поражение Филистимлян?
1SAM|14|31|И поражали Филистимлян в тот день от Михмаса до Аиалона, и народ очень истомился.
1SAM|14|32|И кинулся народ на добычу, и брали овец, волов и телят, и заколали на земле, и ел народ с кровью.
1SAM|14|33|И возвестили Саулу, говоря: вот, народ грешит пред Господом, ест с кровью. И сказал Саул: вы согрешили; привалите ко мне теперь большой камень.
1SAM|14|34|Потом сказал Саул: пройдите между народом и скажите ему: пусть каждый приводит ко мне своего вола и каждый свою овцу, и заколайте здесь и ешьте, и не грешите пред Господом, не ешьте с кровью. И приводили все из народа, каждый своею рукою, вола своего ночью, и заколали там.
1SAM|14|35|И устроил Саул жертвенник Господу: то был первый жертвенник, поставленный им Господу.
1SAM|14|36|И сказал Саул: пойдем [в погоню] за Филистимлянами ночью и оберем их до рассвета и не оставим у них ни одного человека. И сказали: делай все, что хорошо в глазах твоих. Священник же сказал: приступим здесь к Богу.
1SAM|14|37|И вопросил Саул Бога: идти ли мне [в погоню] за Филистимлянами? предашь ли их в руки Израиля? Но Он не отвечал ему в тот день.
1SAM|14|38|Тогда сказал Саул: пусть подойдут сюда все начальники народа и разведают и узнают, на ком грех ныне?
1SAM|14|39|ибо, – жив Господь, спасший Израиля, – если окажется и на Ионафане, сыне моем, то и он умрет непременно. Но никто не отвечал ему из всего народа.
1SAM|14|40|И сказал [Саул] всем Израильтянам: станьте вы по одну сторону, а я и сын мой Ионафан станем по другую сторону. И отвечал народ Саулу: делай, что хорошо в глазах твоих.
1SAM|14|41|И сказал Саул: Господи, Боже Израилев! дай знамение. И уличены были Ионафан и Саул, а народ вышел [правым].
1SAM|14|42|Тогда сказал Саул: бросьте жребий между мною и между Ионафаном, сыном моим. и пал жребий на Ионафана.
1SAM|14|43|И сказал Саул Ионафану: расскажи мне, что сделал ты? И рассказал ему Ионафан и сказал: я отведал концом палки, которая в руке моей, немного меду; и вот, я должен умереть.
1SAM|14|44|И сказал Саул: пусть то и то сделает мне Бог, и еще больше сделает; ты, Ионафан, должен сегодня умереть!
1SAM|14|45|Но народ сказал Саулу: Ионафану ли умереть, который доставил столь великое спасение Израилю? Да не будет этого! Жив Господь, и волос не упадет с головы его на землю, ибо с Богом он действовал ныне. И освободил народ Ионафана, и не умер он.
1SAM|14|46|И возвратился Саул от преследования Филистимлян; Филистимляне же пошли в свое место.
1SAM|14|47|И утвердил Саул свое царствование над Израилем, и воевал со всеми окрестными врагами своими, с Моавом и с Аммонитянами, и с Едомом и с царями Совы и с Филистимлянами, и везде, против кого ни обращался, имел успех.
1SAM|14|48|И устроил войско, и поразил Амалика, и освободил Израиля от руки грабителей его.
1SAM|14|49|Сыновья у Саула были: Ионафан, Иессуи и Мелхисуа; а имена двух дочерей его: имя старшей – Мерова, а имя младшей – Мелхола.
1SAM|14|50|Имя же жены Сауловой – Ахиноамь, дочь Ахимааца; а имя начальника войска его – Авенир, сын Нира, дяди Саулова.
1SAM|14|51|Кис, отец Саулов, и Нир, отец Авенира, были сыновьями Авиила.
1SAM|14|52|И была упорная война против Филистимлян во все время Саулово. И когда Саул видел какого–либо человека сильного и воинственного, брал его к себе.
1SAM|15|1|И сказал Самуил Саулу: Господь послал меня помазать тебя царем над народом Его, над Израилем; теперь послушай гласа Господа.
1SAM|15|2|Так говорит Господь Саваоф: вспомнил Я о том, что сделал Амалик Израилю, как он противостал ему на пути, когда он шел из Египта;
1SAM|15|3|теперь иди и порази Амалика, и истреби все, что у него; и не давай пощады ему, но предай смерти от мужа до жены, от отрока до грудного младенца, от вола до овцы, от верблюда до осла.
1SAM|15|4|И собрал Саул народ и насчитал их в Телаиме двести тысяч Израильтян пеших и десять тысяч из колена Иудина.
1SAM|15|5|И дошел Саул до города Амаликова, и сделал засаду в долине.
1SAM|15|6|И сказал Саул Кинеянам: пойдите, отделитесь, выйдите из среды Амалика, чтобы мне не погубить вас с ним, ибо вы оказали благосклонность всем Израильтянам, когда они шли из Египта. И отделились Кинеяне из среды Амалика.
1SAM|15|7|И поразил Саул Амалика от Хавилы до окрестностей Сура, что пред Египтом;
1SAM|15|8|и Агага, царя Амаликова, захватил живого, а народ весь истребил мечом.
1SAM|15|9|Но Саул и народ пощадили Агага и лучших из овец и волов и откормленных ягнят, и все хорошее, и не хотели истребить, а все вещи маловажные и худые истребили.
1SAM|15|10|И было слово Господа к Самуилу такое:
1SAM|15|11|жалею, что поставил Я Саула царем, ибо он отвратился от Меня и слова Моего не исполнил. И опечалился Самуил и взывал к Господу целую ночь.
1SAM|15|12|И встал Самуил рано утром [и пошел] навстречу Саулу. И известили Самуила, что Саул ходил на Кармил и там поставил себе памятник, и сошел в Галгал.
1SAM|15|13|Когда пришел Самуил к Саулу, то Саул сказал ему: благословен ты у Господа; я исполнил слово Господа.
1SAM|15|14|И сказал Самуил: а что это за блеяние овец в ушах моих и мычание волов, которое я слышу?
1SAM|15|15|И сказал Саул: привели их от Амалика, так как народ пощадил лучших из овец и волов для жертвоприношения Господу Богу твоему; прочее же мы истребили.
1SAM|15|16|И сказал Самуил Саулу: подожди, я скажу тебе, что сказал мне Господь ночью. И сказал ему Саул: говори.
1SAM|15|17|И сказал Самуил: не малым ли ты был в глазах твоих, когда сделался главою колен Израилевых, и Господь помазал тебя царем над Израилем?
1SAM|15|18|И послал тебя Господь в путь, сказав: "иди и предай заклятию нечестивых Амаликитян и воюй против них, доколе не уничтожишь их".
1SAM|15|19|Зачем же ты не послушал гласа Господа и бросился на добычу, и сделал зло пред очами Господа?
1SAM|15|20|И сказал Саул Самуилу: я послушал гласа Господа и пошел в путь, куда послал меня Господь, и привел Агага, царя Амаликитского, а Амалика истребил;
1SAM|15|21|народ же из добычи, из овец и волов, взял лучшее из заклятого, для жертвоприношения Господу Богу твоему, в Галгале.
1SAM|15|22|И отвечал Самуил: неужели всесожжения и жертвы столько же приятны Господу, как послушание гласу Господа? Послушание лучше жертвы и повиновение лучше тука овнов;
1SAM|15|23|ибо непокорность есть [такой же] грех, что волшебство, и противление [то же, что] идолопоклонство; за то, что ты отверг слово Господа, и Он отверг тебя, чтобы ты не был царем.
1SAM|15|24|И сказал Саул Самуилу: согрешил я, ибо преступил повеление Господа и слово твое; но я боялся народа и послушал голоса их;
1SAM|15|25|теперь же сними с меня грех мой и воротись со мною, чтобы я поклонился Господу.
1SAM|15|26|И отвечал Самуил Саулу: не ворочусь я с тобою, ибо ты отверг слово Господа, и Господь отверг тебя, чтобы ты не был царем над Израилем.
1SAM|15|27|И обратился Самуил, чтобы уйти. Но [Саул] ухватился за край одежды его и разодрал ее.
1SAM|15|28|Тогда сказал Самуил: ныне отторг Господь царство Израильское от тебя и отдал его ближнему твоему, лучшему тебя;
1SAM|15|29|и не скажет неправды и не раскается Верный Израилев; ибо не человек Он, чтобы раскаяться Ему.
1SAM|15|30|И сказал [Саул]: я согрешил, но почти меня ныне пред старейшинами народа моего и пред Израилем и воротись со мною, и я поклонюсь Господу Богу твоему.
1SAM|15|31|И возвратился Самуил за Саулом, и поклонился Саул Господу.
1SAM|15|32|Потом сказал Самуил: приведите ко мне Агага, царя Амаликитского. И подошел к нему Агаг дрожащий, и сказал Агаг: конечно горечь смерти миновалась?
1SAM|15|33|Но Самуил сказал: как меч твой жен лишал детей, так мать твоя между женами пусть лишена будет [сына]. И разрубил Самуил Агага пред Господом в Галгале.
1SAM|15|34|И отошел Самуил в Раму, а Саул пошел в дом свой, в Гиву Саулову.
1SAM|15|35|И более не видался Самуил с Саулом до дня смерти своей; но печалился Самуил о Сауле, потому что Господь раскаялся, что воцарил Саула над Израилем.
1SAM|16|1|И сказал Господь Самуилу: доколе будешь ты печалиться о Сауле, которого Я отверг, чтоб он не был царем над Израилем? Наполни рог твой елеем и пойди; Я пошлю тебя к Иессею Вифлеемлянину, ибо между сыновьями его Я усмотрел Себе царя.
1SAM|16|2|И сказал Самуил: как я пойду? Саул услышит и убьет меня. Господь сказал: возьми в руку твою телицу из стада и скажи: "я пришел для жертвоприношения Господу";
1SAM|16|3|и пригласи Иессея к жертве; Я укажу тебе, что делать тебе, и ты помажешь Мне того, о котором Я скажу тебе.
1SAM|16|4|И сделал Самуил так, как сказал ему Господь. Когда пришел он в Вифлеем, то старейшины города с трепетом вышли навстречу ему и сказали: мирен ли приход твой?
1SAM|16|5|И отвечал он: мирен, для жертвоприношения Господу пришел я; освятитесь и идите со мною к жертвоприношению. И освятил Иессея и сыновей его и пригласил их к жертве.
1SAM|16|6|И когда они пришли, он, увидев Елиава, сказал: верно, сей пред Господом помазанник Его!
1SAM|16|7|Но Господь сказал Самуилу: не смотри на вид его и на высоту роста его; Я отринул его; Я [смотрю не так], как смотрит человек; ибо человек смотрит на лице, а Господь смотрит на сердце.
1SAM|16|8|И позвал Иессей Аминадава и подвел его к Самуилу, и сказал Самуил: и этого не избрал Господь.
1SAM|16|9|И подвел Иессей Самму, и сказал [Самуил]: и этого не избрал Господь.
1SAM|16|10|Так подводил Иессей к Самуилу семерых сыновей своих, но Самуил сказал Иессею: [никого] из этих не избрал Господь.
1SAM|16|11|И сказал Самуил Иессею: все ли дети здесь? И отвечал Иессей: есть еще меньший; он пасет овец. И сказал Самуил Иессею: пошли и возьми его, ибо мы не сядем обедать, доколе не придет он сюда.
1SAM|16|12|И послал [Иессей] и привели его. Он был белокур, с красивыми глазами и приятным лицем. И сказал Господь: встань, помажь его, ибо это он.
1SAM|16|13|И взял Самуил рог с елеем и помазал его среди братьев его, и почивал Дух Господень на Давиде с того дня и после; Самуил же встал и отошел в Раму.
1SAM|16|14|А от Саула отступил Дух Господень, и возмущал его злой дух от Господа.
1SAM|16|15|И сказали слуги Сауловы ему: вот, злой дух от Бога возмущает тебя;
1SAM|16|16|пусть господин наш прикажет слугам своим, [которые] пред тобою, поискать человека, искусного в игре на гуслях, и когда придет на тебя злой дух от Бога, то он, играя рукою своею, будет успокоивать тебя.
1SAM|16|17|И отвечал Саул слугам своим: найдите мне человека, хорошо играющего, и представьте его ко мне.
1SAM|16|18|Тогда один из слуг его сказал: вот, я видел у Иессея Вифлеемлянина сына, умеющего играть, человека храброго и воинственного, и разумного в речах и видного собою, и Господь с ним.
1SAM|16|19|И послал Саул вестников к Иессею и сказал: пошли ко мне Давида, сына твоего, который при стаде.
1SAM|16|20|И взял Иессей осла с хлебом и мех с вином и одного козленка, и послал с Давидом, сыном своим, к Саулу.
1SAM|16|21|И пришел Давид к Саулу и служил пред ним, и очень понравился ему и сделался его оруженосцем.
1SAM|16|22|И послал Саул сказать Иессею: пусть Давид служит при мне, ибо он снискал благоволение в глазах моих.
1SAM|16|23|И когда дух от Бога бывал на Сауле, то Давид, взяв гусли, играл, – и отраднее и лучше становилось Саулу, и дух злой отступал от него.
1SAM|17|1|Филистимляне собрали войска свои для войны и собрались в Сокхофе, что в Иудее, и расположились станом между Сокхофом и Азеком в Ефес–Даммиме.
1SAM|17|2|А Саул и Израильтяне собрались и расположились станом в долине дуба и приготовились к войне против Филистимлян.
1SAM|17|3|И стали Филистимляне на горе с одной стороны, и Израильтяне на горе с другой стороны, а между ними была долина.
1SAM|17|4|И выступил из стана Филистимского единоборец, по имени Голиаф, из Гефа; ростом он – шести локтей и пяди.
1SAM|17|5|Медный шлем на голове его; и одет он был в чешуйчатую броню, и вес брони его – пять тысяч сиклей меди;
1SAM|17|6|медные наколенники на ногах его, и медный щит за плечами его;
1SAM|17|7|и древко копья его, как навой у ткачей; а самое копье его в шестьсот сиклей железа, и пред ним шел оруженосец.
1SAM|17|8|И стал [он] и кричал к полкам Израильским, говоря им: зачем вышли вы воевать? Не Филистимлянин ли я, а вы рабы Сауловы? Выберите у себя человека, и пусть сойдет ко мне;
1SAM|17|9|если он может сразиться со мною и убьет меня, то мы будем вашими рабами; если же я одолею его и убью его, то вы будете нашими рабами и будете служить нам.
1SAM|17|10|И сказал Филистимлянин: сегодня я посрамлю полки Израильские; дайте мне человека, и мы сразимся вдвоем.
1SAM|17|11|И услышали Саул и все Израильтяне эти слова Филистимлянина, и очень испугались и ужаснулись.
1SAM|17|12|Давид же был сын Ефрафянина из Вифлеема Иудина, по имени Иессея, у которого было восемь сыновей. Этот человек во дни Саула достиг старости и был старший между мужами.
1SAM|17|13|Три старших сына Иессеевы пошли с Саулом на войну; имена трех сыновей его, пошедших на войну: старший – Елиав, второй за ним – Аминадав, и третий – Самма;
1SAM|17|14|Давид же был меньший. Трое старших пошли с Саулом,
1SAM|17|15|а Давид возвратился от Саула, чтобы пасти овец отца своего в Вифлееме.
1SAM|17|16|И выступал Филистимлянин тот утром и вечером и выставлял себя сорок дней.
1SAM|17|17|И сказал Иессей Давиду, сыну своему: возьми для братьев своих ефу сушеных зерен и десять этих хлебов и отнеси поскорее в стан к твоим братьям;
1SAM|17|18|а эти десять сыров отнеси тысяченачальнику и наведайся о здоровье братьев и узнай о нуждах их.
1SAM|17|19|Саул и они и все Израильтяне [находились] в долине дуба и готовились к сражению с Филистимлянами.
1SAM|17|20|И встал Давид рано утром, и поручил овец сторожу, и, взяв ношу, пошел, как приказал ему Иессей, и пришел к обозу, когда войско выведено было в строй и с криком готовилось к сражению.
1SAM|17|21|И расположили Израильтяне и Филистимляне строй против строя.
1SAM|17|22|Давид оставил свою ношу обозному сторожу и побежал в ряды и, придя, спросил братьев своих о здоровье.
1SAM|17|23|И вот, когда он разговаривал с ними, единоборец, по имени Голиаф, Филистимлянин из Гефа, выступает из рядов Филистимских и говорит те слова, и Давид услышал [их].
1SAM|17|24|И все Израильтяне, увидев этого человека, убегали от него и весьма боялись.
1SAM|17|25|И говорили Израильтяне: видите этого выступающего человека? Он выступает, чтобы поносить Израиля. Если бы кто убил его, одарил бы того царь великим богатством, и дочь свою выдал бы за него, и дом отца его сделал бы свободным в Израиле.
1SAM|17|26|И сказал Давид людям, стоящим с ним: что сделают тому, кто убьет этого Филистимлянина и снимет поношение с Израиля? ибо кто этот необрезанный Филистимлянин, что так поносит воинство Бога живаго?
1SAM|17|27|И сказал ему народ те же слова, говоря: вот что сделано будет тому человеку, который убьет его.
1SAM|17|28|И услышал Елиав, старший брат Давида, что говорил он с людьми, и рассердился Елиав на Давида и сказал: зачем ты сюда пришел и на кого оставил немногих овец тех в пустыне? Я знаю высокомерие твое и дурное сердце твое, ты пришел посмотреть на сражение.
1SAM|17|29|И сказал Давид: что же я сделал? не слова ли это?
1SAM|17|30|И отворотился от него к другому и говорил те же слова, и отвечал ему народ по–прежнему.
1SAM|17|31|И услышали слова, которые говорил Давид, и пересказали Саулу, и тот призвал его.
1SAM|17|32|И сказал Давид Саулу: пусть никто не падает духом из–за него; раб твой пойдет и сразится с этим Филистимлянином.
1SAM|17|33|И сказал Саул Давиду: не можешь ты идти против этого Филистимлянина, чтобы сразиться с ним, ибо ты еще юноша, а он воин от юности своей.
1SAM|17|34|И сказал Давид Саулу: раб твой пас овец у отца своего, и когда, бывало, приходил лев или медведь и уносил овцу из стада,
1SAM|17|35|то я гнался за ним и нападал на него и отнимал из пасти его; а если он бросался на меня, то я брал его за космы и поражал его и умерщвлял его;
1SAM|17|36|и льва и медведя убивал раб твой, и с этим Филистимлянином необрезанным будет то же, что с ними, потому что так поносит воинство Бога живаго.
1SAM|17|37|И сказал Давид: Господь, Который избавлял меня от льва и медведя, избавит меня и от руки этого Филистимлянина. И сказал Саул Давиду: иди, и да будет Господь с тобою.
1SAM|17|38|И одел Саул Давида в свои одежды, и возложил на голову его медный шлем, и надел на него броню.
1SAM|17|39|И опоясался Давид мечом его сверх одежды и начал ходить, ибо не привык [к такому вооружению]; потом сказал Давид Саулу: я не могу ходить в этом, я не привык. И снял Давид все это с себя.
1SAM|17|40|И взял посох свой в руку свою, и выбрал себе пять гладких камней из ручья, и положил их в пастушескую сумку, которая была с ним; и с сумкою и с пращею в руке своей выступил против Филистимлянина.
1SAM|17|41|Выступил и Филистимлянин, идя и приближаясь к Давиду, и оруженосец шел впереди его.
1SAM|17|42|И взглянул Филистимлянин и, увидев Давида, с презрением посмотрел на него, ибо он был молод, белокур и красив лицем.
1SAM|17|43|И сказал Филистимлянин Давиду: что ты идешь на меня с палкою? разве я собака? И проклял Филистимлянин Давида своими богами.
1SAM|17|44|И сказал Филистимлянин Давиду: подойди ко мне, и я отдам тело твое птицам небесным и зверям полевым.
1SAM|17|45|А Давид отвечал Филистимлянину: ты идешь против меня с мечом и копьем и щитом, а я иду против тебя во имя Господа Саваофа, Бога воинств Израильских, которые ты поносил;
1SAM|17|46|ныне предаст тебя Господь в руку мою, и я убью тебя, и сниму с тебя голову твою, и отдам трупы войска Филистимского птицам небесным и зверям земным, и узнает вся земля, что есть Бог в Израиле;
1SAM|17|47|и узнает весь этот сонм, что не мечом и копьем спасает Господь, ибо это война Господа, и Он предаст вас в руки наши.
1SAM|17|48|Когда Филистимлянин поднялся и стал подходить и приближаться навстречу Давиду, Давид поспешно побежал к строю навстречу Филистимлянину.
1SAM|17|49|И опустил Давид руку свою в сумку и взял оттуда камень, и бросил из пращи и поразил Филистимлянина в лоб, так что камень вонзился в лоб его, и он упал лицем на землю.
1SAM|17|50|Так одолел Давид Филистимлянина пращею и камнем, и поразил Филистимлянина и убил его; меча же не было в руках Давида.
1SAM|17|51|Тогда Давид подбежал и, наступив на Филистимлянина, взял меч его и вынул его из ножен, ударил его и отсек им голову его; Филистимляне, увидев, что силач их умер, побежали.
1SAM|17|52|И поднялись мужи Израильские и Иудейские, и воскликнули и гнали Филистимлян до входа в долину и до ворот Аккарона. И падали поражаемые Филистимляне по дороге Шааримской до Гефа и до Аккарона.
1SAM|17|53|И возвратились сыны Израилевы из погони за Филистимлянами и разграбили стан их.
1SAM|17|54|И взял Давид голову Филистимлянина и отнес ее в Иерусалим, а оружие его положил в шатре своем.
1SAM|17|55|Когда Саул увидел Давида, выходившего против Филистимлянина, то сказал Авениру, начальнику войска: Авенир, чей сын этот юноша? Авенир сказал: да живет душа твоя, царь; я не знаю.
1SAM|17|56|И сказал царь: так спроси, чей сын этот юноша?
1SAM|17|57|Когда же Давид возвращался после поражения Филистимлянина, то Авенир взял его и привел к Саулу, и голова Филистимлянина была в руке его.
1SAM|17|58|И спросил его Саул: чей ты сын, юноша? И отвечал Давид: сын раба твоего Иессея из Вифлеема.
1SAM|18|1|Когда кончил [Давид] разговор с Саулом, душа Ионафана прилепилась к душе его, и полюбил его Ионафан, как свою душу.
1SAM|18|2|И взял его Саул в тот день и не позволил ему возвратиться в дом отца его.
1SAM|18|3|Ионафан же заключил с Давидом союз, ибо полюбил его, как свою душу.
1SAM|18|4|И снял Ионафан верхнюю одежду свою, которая была на нем, и отдал ее Давиду, также и прочие одежды свои, и меч свой, и лук свой, и пояс свой.
1SAM|18|5|И Давид действовал благоразумно везде, куда ни посылал его Саул, и сделал его Саул начальником над военными людьми; и это понравилось всему народу и слугам Сауловым.
1SAM|18|6|Когда они шли, при возвращении Давида с победы над Филистимлянином, то женщины из всех городов Израильских выходили навстречу Саулу царю с пением и плясками, с торжественными тимпанами и с кимвалами.
1SAM|18|7|И восклицали игравшие женщины, говоря: Саул победил тысячи, а Давид – десятки тысяч!
1SAM|18|8|И Саул сильно огорчился, и неприятно было ему это слово, и он сказал: Давиду дали десятки тысяч, а мне тысячи; ему недостает только царства.
1SAM|18|9|И с того дня и потом подозрительно смотрел Саул на Давида.
1SAM|18|10|И было на другой день: напал злой дух от Бога на Саула, и он бесновался в доме своем, а Давид играл рукою своею на струнах, как и в другие дни; в руке у Саула было копье.
1SAM|18|11|И бросил Саул копье, подумав: пригвожду Давида к стене; но Давид два раза уклонился от него.
1SAM|18|12|И стал бояться Саул Давида, потому что Господь был с ним, а от Саула отступил.
1SAM|18|13|И удалил его Саул от себя и поставил его у себя тысяченачальником, и он выходил и входил пред народом.
1SAM|18|14|И Давид во всех делах своих поступал благоразумно, и Господь [был] с ним.
1SAM|18|15|И Саул видел, что он очень благоразумен, и боялся его.
1SAM|18|16|А весь Израиль и Иуда любили Давида, ибо он выходил и входил пред ними.
1SAM|18|17|И сказал Саул Давиду: вот старшая дочь моя, Мерова; я дам ее тебе в жену, только будь у меня храбрым и веди войны Господни. Ибо Саул думал: пусть не моя рука будет на нем, но рука Филистимлян будет на нем.
1SAM|18|18|Но Давид сказал Саулу: кто я, и что жизнь моя и род отца моего в Израиле, чтобы мне быть зятем царя?
1SAM|18|19|А когда наступило время отдать Мерову, дочь Саула, Давиду, то она выдана была в замужество за Адриэла из Мехолы.
1SAM|18|20|Но Давида полюбила [другая] дочь Саула, Мелхола; и когда возвестили [об этом] Саулу, то это было приятно ему.
1SAM|18|21|Саул думал: отдам ее за него, и она будет ему сетью, и рука Филистимлян будет на нем. И сказал Саул Давиду: чрез другую ты породнишься ныне со мною.
1SAM|18|22|И приказал Саул слугам своим: скажите Давиду тайно: вот, царь благоволит к тебе, и все слуги его любят тебя; итак будь зятем царя.
1SAM|18|23|И передали слуги Сауловы в уши Давиду все слова эти. И сказал Давид: разве легко кажется вам быть зятем царя? я – человек бедный и незначительный.
1SAM|18|24|И донесли Саулу слуги его и сказали: вот что говорит Давид.
1SAM|18|25|И сказал Саул: так скажите Давиду: царь не хочет вена, кроме ста краеобрезаний Филистимских, в отмщение врагам царя. Ибо Саул имел в мыслях погубить Давида руками Филистимлян.
1SAM|18|26|И пересказали слуги его Давиду эти слова, и понравилось Давиду сделаться зятем царя.
1SAM|18|27|Еще не прошли назначенные дни, как Давид встал и пошел сам и люди его с ним, и убил двести человек Филистимлян, и принес Давид краеобрезания их, и представил их в полном количестве царю, чтобы сделаться зятем царя. И выдал Саул за него Мелхолу, дочь свою, в замужество.
1SAM|18|28|И увидел Саул и узнал, что Господь с Давидом, и что Мелхола, дочь Саула, любила [Давида].
1SAM|18|29|И стал Саул еще больше бояться Давида и сделался врагом его на всю жизнь.
1SAM|18|30|И когда вожди Филистимские вышли [на войну], Давид, с самого выхода их, действовал благоразумнее всех слуг Сауловых, и весьма прославилось имя его.
1SAM|19|1|И говорил Саул Ионафану, сыну своему, и всем слугам своим, чтобы умертвить Давида; но Ионафан, сын Саула, очень любил Давида.
1SAM|19|2|И известил Ионафан Давида, говоря: отец мой Саул ищет умертвить тебя; итак берегись завтра; скройся и будь в потаенном месте;
1SAM|19|3|а я выйду и стану подле отца моего на поле, где ты будешь, и поговорю о тебе отцу моему, и что увижу, расскажу тебе.
1SAM|19|4|И говорил Ионафан доброе о Давиде Саулу, отцу своему, и сказал ему: да не грешит царь против раба своего Давида, ибо он ничем не согрешил против тебя, и дела его весьма полезны для тебя;
1SAM|19|5|он подвергал опасности душу свою, чтобы поразить Филистимлянина, и Господь соделал великое спасение всему Израилю; ты видел [это] и радовался; для чего же ты хочешь согрешить [против] невинной крови и умертвить Давида без причины?
1SAM|19|6|И послушал Саул голоса Ионафана и поклялся Саул: жив Господь, [Давид] не умрет.
1SAM|19|7|И позвал Ионафан Давида, и пересказал ему Ионафан все слова сии, и привел Ионафан Давида к Саулу, и он был при нем, как вчера и третьего дня.
1SAM|19|8|Опять началась война, и вышел Давид, и воевал с Филистимлянами, и нанес им великое поражение, и они побежали от него.
1SAM|19|9|И злой дух от Бога напал на Саула, и он сидел в доме своем, и копье его было в руке его, а Давид играл рукою своею на струнах.
1SAM|19|10|И хотел Саул пригвоздить Давида копьем к стене, но Давид отскочил от Саула, и копье вонзилось в стену; Давид же убежал и спасся в ту ночь.
1SAM|19|11|И послал Саул слуг в дом к Давиду, чтобы стеречь его и убить его до утра. И сказала Давиду Мелхола, жена его: если ты не спасешь души твоей в эту ночь, то завтра будешь убит.
1SAM|19|12|И спустила Мелхола Давида из окна, и он пошел, и убежал и спасся.
1SAM|19|13|Мелхола же взяла статую и положила на постель, а в изголовье ее положила козью кожу, и покрыла одеждою.
1SAM|19|14|И послал Саул слуг, чтобы взять Давида; но [Мелхола] сказала: он болен.
1SAM|19|15|И послал Саул слуг, чтобы осмотреть Давида, говоря: принесите его ко мне на постели, чтоб убить его.
1SAM|19|16|И пришли слуги, и вот, на постели статуя, а в изголовье ее козья кожа.
1SAM|19|17|Тогда Саул сказал Мелхоле: для чего ты так обманула меня и отпустила врага моего, чтоб он убежал? И сказала Мелхола Саулу: он сказал мне: отпусти меня, иначе я убью тебя.
1SAM|19|18|И убежал Давид и спасся, и пришел к Самуилу в Раму и рассказал ему все, что делал с ним Саул. И пошел он с Самуилом, и остановились они в Навафе.
1SAM|19|19|И донесли Саулу, говоря: вот, Давид в Навафе, в Раме.
1SAM|19|20|И послал Саул слуг взять Давида, и [когда] увидели они сонм пророков пророчествующих и Самуила, начальствующего над ними, то Дух Божий сошел на слуг Саула, и они стали пророчествовать.
1SAM|19|21|Донесли [об этом] Саулу, и он послал других слуг, но и эти стали пророчествовать. Потом послал Саул третьих слуг, и эти стали пророчествовать.
1SAM|19|22|Саул сам пошел в Раму, и дошел до большого источника, что в Сефе, и спросил, говоря: где Самуил и Давид? И сказали: вот, в Навафе, в Раме.
1SAM|19|23|И пошел он туда в Наваф в Раме, и на него сошел Дух Божий, и он шел и пророчествовал, доколе не пришел в Наваф в Раме.
1SAM|19|24|И снял и он одежды свои, и пророчествовал пред Самуилом, и весь день тот и всю ту ночь лежал неодетый; поэтому говорят: "неужели и Саул во пророках?"
1SAM|20|1|Давид убежал из Навафа в Раме и пришел и сказал Ионафану: что сделал я, в чем неправда моя, чем согрешил я пред отцом твоим, что он ищет души моей?
1SAM|20|2|И сказал ему [Ионафан]: нет, ты не умрешь; вот, отец мой не делает ни большого, ни малого дела, не открыв ушам моим; для чего же бы отцу моему скрывать от меня это дело? этого не будет.
1SAM|20|3|Давид клялся и говорил: отец твой хорошо знает, что я нашел благоволение в очах твоих, и потому говорит сам в себе: "пусть не знает о том Ионафан, чтобы не огорчился"; но жив Господь и жива душа твоя! один только шаг между мною и смертью.
1SAM|20|4|И сказал Ионафан Давиду: чего желает душа твоя, я сделаю для тебя.
1SAM|20|5|И сказал Давид Ионафану: вот, завтра новомесячие, и я должен сидеть с царем за столом; но отпусти меня, и я скроюсь в поле до вечера третьего дня.
1SAM|20|6|Если отец твой спросит обо мне, ты скажи: "Давид выпросился у меня сходить в свой город Вифлеем; потому что там годичное жертвоприношение всего родства его".
1SAM|20|7|Если на это он скажет: "хорошо", то мир рабу твоему; а если он разгневается, то знай, что злое дело решено у него.
1SAM|20|8|Ты же сделай милость рабу твоему, – ибо ты принял раба твоего в завет Господень с тобою, – и если есть какая вина на мне, то умертви ты меня; зачем тебе вести меня к отцу твоему?
1SAM|20|9|И сказал Ионафан: никак не будет этого с тобою; ибо, если я узнаю наверное, что у отца моего решено злое дело совершить над тобою, то неужели не извещу тебя об этом?
1SAM|20|10|И сказал Давид Ионафану: кто известит меня, если отец твой ответит тебе сурово?
1SAM|20|11|И сказал Ионафан Давиду: иди, выйдем в поле. И вышли оба в поле.
1SAM|20|12|И сказал Ионафан Давиду: жив Господь Бог Израилев! я завтра около этого времени, или послезавтра, выпытаю у отца моего; и если он благосклонен к Давиду, и я тогда же не пошлю к тебе и не открою пред ушами твоими,
1SAM|20|13|пусть то и то сделает Господь с Ионафаном и еще больше сделает. Если же отец мой замышляет сделать тебе зло, и это открою в уши твои, и отпущу тебя, и тогда иди с миром: и да будет Господь с тобою, как был с отцом моим!
1SAM|20|14|Но и ты, если я буду еще жив, окажи мне милость Господню.
1SAM|20|15|А если я умру, то не отними милости твоей от дома моего во веки, даже и тогда, когда Господь истребит с лица земли всех врагов Давида.
1SAM|20|16|Так заключил Ионафан завет с домом Давида [и сказал]: да взыщет Господь с врагов Давида!
1SAM|20|17|И снова Ионафан клялся Давиду своею любовью к нему, ибо любил его, как свою душу.
1SAM|20|18|И сказал ему Ионафан: завтра новомесячие, и о тебе спросят, ибо место твое будет не занято;
1SAM|20|19|поэтому на третий день ты спустись и поспеши на то место, где скрывался ты прежде, и сядь у камня Азель;
1SAM|20|20|а я в ту сторону пущу три стрелы, как будто стреляя в цель;
1SAM|20|21|потом пошлю отрока, [говоря]: "пойди, найди стрелы"; и если я скажу отроку: "вот, стрелы сзади тебя, возьми их", то приди ко мне, ибо мир тебе, и, жив Господь, ничего [тебе не будет];
1SAM|20|22|если же так скажу отроку: "вот, стрелы впереди тебя", то ты уходи, ибо отпускает тебя Господь;
1SAM|20|23|а тому, что мы говорили, я и ты, [свидетель] Господь между мною и тобою во веки.
1SAM|20|24|И скрылся Давид на поле. И наступило новомесячие, и сел царь обедать.
1SAM|20|25|Царь сел на своем месте, по обычаю, на седалище у стены, и Ионафан встал, и Авенир сел подле Саула; место же Давида осталось праздным.
1SAM|20|26|И не сказал Саул в тот день ничего, ибо подумал, что это случайность, что [Давид] нечист, не очистился.
1SAM|20|27|Наступил и второй день новомесячия, а место Давида оставалось праздным. Тогда сказал Саул сыну своему Ионафану: почему сын Иессеев не пришел к обеду ни вчера, ни сегодня?
1SAM|20|28|И отвечал Ионафан Саулу: Давид выпросился у меня в Вифлеем;
1SAM|20|29|он говорил: "отпусти меня, ибо у нас в городе родственное жертвоприношение, и мой брат пригласил меня; итак, если я нашел благоволение в очах твоих, схожу я и повидаюсь со своими братьями"; поэтому он и не пришел к обеду царя.
1SAM|20|30|Тогда сильно разгневался Саул на Ионафана и сказал ему: сын негодный и непокорный! разве я не знаю, что ты подружился с сыном Иессеевым на срам себе и на срам матери твоей?
1SAM|20|31|ибо во все дни, доколе сын Иессеев будет жить на земле, не устоишь ни ты, ни царство твое; теперь же пошли и приведи его ко мне, ибо он обречен на смерть.
1SAM|20|32|И отвечал Ионафан Саулу, отцу своему, и сказал ему: за что умерщвлять его? что он сделал?
1SAM|20|33|Тогда Саул бросил копье в него, чтобы поразить его. И Ионафан понял, что отец его решился убить Давида.
1SAM|20|34|И встал Ионафан из–за стола в великом гневе и не обедал во второй день новомесячия, потому что скорбел о Давиде и потому что обидел его отец его.
1SAM|20|35|На другой день утром вышел Ионафан в поле, во время, которое назначил Давиду, и малый отрок с ним.
1SAM|20|36|И сказал он отроку: беги, ищи стрелы, которые я пускаю. Отрок побежал, а он пускал стрелы так, что они летели дальше [отрока].
1SAM|20|37|И побежал отрок туда, куда Ионафан пускал стрелы, и закричал Ионафан вслед отроку и сказал: смотри, стрела впереди тебя.
1SAM|20|38|И опять кричал Ионафан вслед отроку: скорей беги, не останавливайся. И собрал отрок Ионафанов стрелы и пришел к своему господину.
1SAM|20|39|Отрок же не знал ничего; только Ионафан и Давид знали, в чем дело.
1SAM|20|40|И отдал Ионафан оружие свое отроку, бывшему при нем, и сказал ему: ступай, отнеси в город.
1SAM|20|41|Отрок пошел, а Давид поднялся с южной стороны и пал лицем своим на землю и трижды поклонился; и целовали они друг друга, и плакали оба вместе, но Давид плакал более.
1SAM|20|42|И сказал Ионафан Давиду: иди с миром; а в чем клялись мы оба именем Господа, говоря: "Господь да будет между мною и между тобою и между семенем моим и семенем твоим", то да будет на веки. И встал [Давид] и пошел, а Ионафан возвратился в город.
1SAM|21|1|И пришел Давид в Номву к Ахимелеху священнику, и смутился Ахимелех при встрече с Давидом и сказал ему: почему ты один, и никого нет с тобою?
1SAM|21|2|И сказал Давид Ахимелеху священнику: царь поручил мне дело и сказал мне: "пусть никто не знает, за чем я послал тебя и что поручил тебе"; поэтому людей я оставил на известном месте;
1SAM|21|3|итак, что есть у тебя под рукою, дай мне, хлебов пять, или что найдется.
1SAM|21|4|И отвечал священник Давиду, говоря: нет у меня под рукою простого хлеба, а есть хлеб священный; если только люди [твои] воздержались от женщин!
1SAM|21|5|И отвечал Давид священнику и сказал ему: женщин при нас не было ни вчера, ни третьего дня, со времени, как я вышел, и сосуды отроков чисты, а если дорога нечиста, то [хлеб] останется чистым в сосудах.
1SAM|21|6|И дал ему священник священного хлеба; ибо не было у него хлеба, кроме хлебов предложения, которые взяты были от лица Господа, чтобы по снятии их положить теплые хлебы.
1SAM|21|7|Там находился в тот день пред Господом один из слуг Сауловых, по имени Доик, Идумеянин, начальник пастухов Сауловых.
1SAM|21|8|И сказал Давид Ахимелеху: нет ли здесь у тебя под рукою копья или меча? ибо я не взял с собою ни меча, ни другого оружия, так как поручение царя было спешное.
1SAM|21|9|И сказал священник: вот меч Голиафа Филистимлянина, которого ты поразил в долине дуба, завернутый в одежду, позади ефода; если хочешь, возьми его; другого кроме этого нет здесь. И сказал Давид: нет ему подобного, дай мне его.
1SAM|21|10|И встал Давид, и убежал в тот же день от Саула, и пришел к Анхусу, царю Гефскому.
1SAM|21|11|И сказали Анхусу слуги его: не это ли Давид, царь той страны? не ему ли пели в хороводах и говорили: "Саул поразил тысячи, а Давид – десятки тысяч"?
1SAM|21|12|Давид положил слова эти в сердце своем и сильно боялся Анхуса, царя Гефского.
1SAM|21|13|И изменил лице свое пред ними, и притворился безумным в их глазах, и чертил на дверях, и пускал слюну по бороде своей.
1SAM|21|14|И сказал Анхус рабам своим: видите, он человек сумасшедший; для чего вы привели его ко мне?
1SAM|21|15|разве мало у меня сумасшедших, что вы привели его, чтобы он юродствовал предо мною?
1SAM|21|16|неужели он войдет в дом мой?
1SAM|22|1|И вышел Давид оттуда и убежал в пещеру Одолламскую, и услышали братья его и весь дом отца его и пришли к нему туда.
1SAM|22|2|И собрались к нему все притесненные и все должники и все огорченные душею, и сделался он начальником над ними; и было с ним около четырехсот человек.
1SAM|22|3|Оттуда пошел Давид в Массифу Моавитскую и сказал царю Моавитскому: пусть отец мой и мать моя побудут у вас, доколе я не узнаю, что сделает со мною Бог.
1SAM|22|4|И привел их к царю Моавитскому, и жили они у него все время, доколе Давид был в оном убежище.
1SAM|22|5|Но пророк Гад сказал Давиду: не оставайся в этом убежище, но ступай, иди в землю Иудину. И пошел Давид и пришел в лес Херет.
1SAM|22|6|И услышал Саул, что Давид появился и люди, бывшие с ним. Саул сидел тогда в Гиве под дубом на горе, с копьем в руке, и все слуги его окружали его.
1SAM|22|7|И сказал Саул слугам своим, окружавшим его: послушайте, сыны Вениаминовы, неужели всем вам даст сын Иессея поля и виноградники и всех вас поставит тысяченачальниками и сотниками,
1SAM|22|8|что вы все сговорились против меня, и никто не открыл мне, когда сын мой вступил в дружбу с сыном Иессея, и никто из вас не пожалел о мне и не открыл мне, что сын мой возбудил против меня раба моего строить мне ковы, как это ныне видно?
1SAM|22|9|И отвечал Доик Идумеянин, стоявший со слугами Сауловыми, и сказал: я видел, как сын Иессея приходил в Номву к Ахимелеху, сыну Ахитува,
1SAM|22|10|и тот вопросил о нем Господа, и дал ему продовольствие, и меч Голиафа Филистимлянина отдал ему.
1SAM|22|11|И послал царь призвать Ахимелеха, сына Ахитувова, священника, и весь дом отца его, священников, что в Номве; и пришли они все к царю.
1SAM|22|12|И сказал Саул: послушай, сын Ахитува. И тот отвечал: вот я, господин мой.
1SAM|22|13|И сказал ему Саул: для чего вы сговорились против меня, ты и сын Иессея, что ты дал ему хлебы и меч и вопросил о нем Бога, чтоб он восстал против меня и строил мне ковы, как это ныне видно?
1SAM|22|14|И отвечал Ахимелех царю и сказал: кто из всех рабов твоих верен как Давид? он и зять царя, и исполнитель повелений твоих, и почтен в доме твоем.
1SAM|22|15|Теперь ли я стал вопрошать для него Бога? Нет, не обвиняй в этом, царь, раба твоего и весь дом отца моего, ибо во всем этом деле не знает раб твой ни малого, ни великого.
1SAM|22|16|И сказал царь: ты должен умереть, Ахимелех, ты и весь дом отца твоего.
1SAM|22|17|И сказал царь телохранителям, стоявшим при нем: ступайте, умертвите священников Господних, ибо и их рука с Давидом, и они знали, что он убежал, и не открыли мне. Но слуги царя не хотели поднять рук своих на убиение священников Господних.
1SAM|22|18|И сказал царь Доику: ступай ты и умертви священников. И пошел Доик Идумеянин, и напал на священников, и умертвил в тот день восемьдесят пять мужей, носивших льняной ефод;
1SAM|22|19|и Номву, город священников, поразил мечом; и мужчин и женщин, и юношей и младенцев, и волов и ослов и овец поразил мечом.
1SAM|22|20|Спасся один только сын Ахимелеха, сына Ахитува, по имени Авиафар, и убежал к Давиду.
1SAM|22|21|И рассказал Авиафар Давиду, что Саул умертвил священников Господних.
1SAM|22|22|И сказал Давид Авиафару: я знал в тот день, когда там был Доик Идумеянин, что он непременно донесет Саулу; я виновен во всех душах дома отца твоего;
1SAM|22|23|останься у меня, не бойся, ибо кто будет искать моей души, будет искать и твоей души; ты будешь у меня под охранением.
1SAM|23|1|И известили Давида, говоря: вот, Филистимляне напали на Кеиль и расхищают гумна.
1SAM|23|2|И вопросил Давид Господа, говоря: идти ли мне, и поражу ли я этих Филистимлян? И отвечал Господь Давиду: иди, ты поразишь Филистимлян и спасешь Кеиль.
1SAM|23|3|Но бывшие с Давидом сказали ему: вот, мы боимся здесь в Иудее, как же нам идти в Кеиль против ополчений Филистимских?
1SAM|23|4|Тогда снова вопросил Давид Господа, и отвечал ему Господь и сказал: встань и иди в Кеиль, ибо Я предам Филистимлян в руки твои.
1SAM|23|5|И пошел Давид с людьми своими в Кеиль, и воевал с Филистимлянами, и угнал скот их, и нанес им великое поражение, и спас Давид жителей Кеиля.
1SAM|23|6|Когда Авиафар, сын Ахимелеха, прибежал к Давиду в Кеиль, то принес с собою и ефод.
1SAM|23|7|И донесли Саулу, что Давид пришел в Кеиль, и Саул сказал: Бог предал его в руки мои, ибо он запер себя, войдя в город с воротами и запорами.
1SAM|23|8|И созвал Саул весь народ на войну, чтоб идти к Кеилю, осадить Давида и людей его.
1SAM|23|9|Когда узнал Давид, что Саул задумал против него злое, сказал священнику Авиафару: принеси ефод.
1SAM|23|10|И сказал Давид: Господи Боже Израилев! раб Твой услышал, что Саул хочет придти в Кеиль, разорить город ради меня.
1SAM|23|11|Предадут ли меня жители Кеиля в руки его? И придет ли сюда Саул, как слышал раб Твой? Господи Боже Израилев! открой рабу Твоему. И сказал Господь: придет.
1SAM|23|12|И сказал Давид: предадут ли жители Кеиля меня и людей моих в руки Саула? И сказал Господь: предадут.
1SAM|23|13|Тогда поднялся Давид и люди его, около шестисот человек, и вышли из Кеиля и ходили, где могли. Саулу же было донесено, что Давид убежал из Кеиля, и тогда он отменил поход.
1SAM|23|14|Давид же пребывал в пустыне в неприступных местах и потом на горе в пустыне Зиф. Саул искал его всякий день; но Бог не предал [Давида] в руки его.
1SAM|23|15|И видел Давид, что Саул вышел искать души его; Давид же был в пустыне Зиф в лесу.
1SAM|23|16|И встал Ионафан, сын Саула, и пришел к Давиду в лес, и укрепил его упованием на Бога,
1SAM|23|17|и сказал ему: не бойся, ибо не найдет тебя рука отца моего Саула, и ты будешь царствовать над Израилем, а я буду вторым по тебе; и Саул, отец мой, знает это.
1SAM|23|18|И заключили они между собою завет пред лицем Господа; и Давид остался в лесу, а Ионафан пошел в дом свой.
1SAM|23|19|И пришли Зифеи к Саулу в Гиву, говоря: вот, Давид скрывается у нас в неприступных местах, в лесу, на холме Гахила, что направо от Иесимона;
1SAM|23|20|итак по желанию души твоей, царь, иди; а наше дело будет предать его в руки царя.
1SAM|23|21|И сказал им Саул: благословенны вы у Господа за то, что пожалели о мне;
1SAM|23|22|идите, удостоверьтесь еще, разведайте [и] высмотрите место его, где будет нога его, [и] кто видел его там, ибо мне говорят, что он очень хитер;
1SAM|23|23|и высмотрите, и разведайте о всех убежищах, в которых он скрывается, и возвратитесь ко мне с верным известием, и я пойду с вами; и если он в этой земле, я буду искать его во всех тысячах Иудиных.
1SAM|23|24|И встали они и пошли в Зиф прежде Саула. Давид же и люди его были в пустыне Маон, на равнине, направо от Иесимона.
1SAM|23|25|И пошел Саул с людьми своими искать [его]. Но Давида известили об этом, и он перешел к скале и оставался в пустыне Маон. И услышал Саул, и погнался за Давидом в пустыню Маон.
1SAM|23|26|И шел Саул по одной стороне горы, а Давид с людьми своими был на другой стороне горы. И когда Давид спешил уйти от Саула, а Саул с людьми своими шел в обход Давиду и людям его, чтобы захватить их;
1SAM|23|27|тогда пришел к Саулу вестник, говоря: поспешай и приходи, ибо Филистимляне напали на землю.
1SAM|23|28|И возвратился Саул от преследования Давида и пошел навстречу Филистимлянам; посему и назвали это место: Села–Гаммахлекоф.
1SAM|24|1|И вышел Давид оттуда и жил в безопасных местах Ен–Гадди.
1SAM|24|2|Когда Саул возвратился от Филистимлян, его известили, говоря: вот, Давид в пустыне Ен–Гадди.
1SAM|24|3|И взял Саул три тысячи отборных мужей из всего Израиля и пошел искать Давида и людей его по горам, где живут серны.
1SAM|24|4|И пришел к загону овечьему, при дороге; там была пещера, и зашел туда Саул для нужды; Давид же и люди его сидели в глубине пещеры.
1SAM|24|5|И говорили Давиду люди его: вот день, о котором говорил тебе Господь: "вот, Я предам врага твоего в руки твои, и сделаешь с ним, что тебе угодно". Давид встал и тихонько отрезал край от верхней одежды Саула.
1SAM|24|6|Но после сего больно стало сердцу Давида, что он отрезал край от одежды Саула.
1SAM|24|7|И сказал он людям своим: да не попустит мне Господь сделать это господину моему, помазаннику Господню, чтобы наложить руку мою на него, ибо он помазанник Господень.
1SAM|24|8|И удержал Давид людей своих сими словами и не дал им восстать на Саула. А Саул встал и вышел из пещеры на дорогу.
1SAM|24|9|Потом встал и Давид, и вышел из пещеры, и закричал вслед Саула, говоря: господин мой, царь! Саул оглянулся назад, и Давид пал лицем на землю и поклонился [ему].
1SAM|24|10|И сказал Давид Саулу: зачем ты слушаешь речи людей, которые говорят: "вот, Давид умышляет зло на тебя"?
1SAM|24|11|Вот, сегодня видят глаза твои, что Господь предавал тебя ныне в руки мои в пещере; и мне говорили, чтоб убить тебя; но я пощадил тебя и сказал: "не подниму руки моей на господина моего, ибо он помазанник Господа".
1SAM|24|12|Отец мой! посмотри на край одежды твоей в руке моей; я отрезал край одежды твоей, а тебя не убил: узнай и убедись, что нет в руке моей зла, ни коварства, и я не согрешил против тебя; а ты ищешь души моей, чтоб отнять ее.
1SAM|24|13|Да рассудит Господь между мною и тобою, и да отмстит тебе Господь за меня; но рука моя не будет на тебе,
1SAM|24|14|как говорит древняя притча: "от беззаконных исходит беззаконие". А рука моя не будет на тебе.
1SAM|24|15|Против кого вышел царь Израильский? За кем ты гоняешься? За мертвым псом, за одною блохою.
1SAM|24|16|Господь да будет судьею и рассудит между мною и тобою. Он рассмотрит, разберет дело мое, и спасет меня от руки твоей.
1SAM|24|17|Когда кончил Давид говорить слова сии к Саулу, Саул сказал: твой ли это голос, сын мой Давид? И возвысил Саул голос свой, и плакал,
1SAM|24|18|и сказал Давиду: ты правее меня, ибо ты воздал мне добром, а я воздавал тебе злом;
1SAM|24|19|ты показал это сегодня, поступив со мною милостиво, когда Господь предавал меня в руки твои, ты не убил меня.
1SAM|24|20|Кто, найдя врага своего, отпустил бы его в добрый путь? Господь воздаст тебе добром за то, что сделал ты мне сегодня.
1SAM|24|21|И теперь я знаю, что ты непременно будешь царствовать, и царство Израилево будет твердо в руке твоей.
1SAM|24|22|Итак поклянись мне Господом, что ты не искоренишь потомства моего после меня и не уничтожишь имени моего в доме отца моего.
1SAM|24|23|И поклялся Давид Саулу. И пошел Саул в дом свой, Давид же и люди его взошли в место укрепленное.
1SAM|25|1|И умер Самуил; и собрались все Израильтяне, и плакали по нем, и погребли его в доме его, в Раме. Давид встал и сошел к пустыне Фаран.
1SAM|25|2|Был некто в Маоне, а имение его на Кармиле, человек очень богатый; у него было три тысячи овец и тысяча коз; и был он при стрижке овец своих на Кармиле.
1SAM|25|3|Имя человека того – Навал, а имя жены его – Авигея; эта женщина [была] весьма умная и красивая лицем, а он – человек жестокий и злой нравом; он был из рода Халева.
1SAM|25|4|И услышал Давид в пустыне, что Навал стрижет овец своих.
1SAM|25|5|И послал Давид десять отроков, и сказал Давид отрокам: взойдите на Кармил и пойдите к Навалу, и приветствуйте его от моего имени,
1SAM|25|6|и скажите так: "мир тебе, мир дому твоему, мир всему твоему;
1SAM|25|7|ныне я услышал, что у тебя стригут [овец]. Вот, пастухи твои были с нами, и мы не обижали их, и ничего у них не пропало во все время их пребывания на Кармиле;
1SAM|25|8|спроси слуг твоих, и они скажут тебе; итак да найдут отроки благоволение в глазах твоих, ибо в добрый день пришли мы; дай же рабам твоим и сыну твоему Давиду, что найдет рука твоя".
1SAM|25|9|И пошли люди Давидовы, и сказали Навалу от имени Давида все эти слова, и умолкли.
1SAM|25|10|И Навал, отвечал слугам Давидовым, и сказал: кто такой Давид, и кто такой сын Иессеев? ныне стало много рабов, бегающих от господ своих;
1SAM|25|11|неужели мне взять хлебы мои и воду мою, и мясо, приготовленное мною для стригущих овец у меня, и отдать людям, о которых не знаю, откуда они?
1SAM|25|12|И пошли назад люди Давида своим путем и возвратились, и пришли и пересказали ему все слова сии.
1SAM|25|13|Тогда Давид сказал людям своим: опояшьтесь каждый мечом своим. И все опоясались мечами своими, опоясался и сам Давид своим мечом, и пошли за Давидом около четырехсот человек, а двести остались при обозе.
1SAM|25|14|Авигею же, жену Навала, известил один из слуг, сказав: вот, Давид присылал из пустыни послов приветствовать нашего господина, но он обошелся с ними грубо;
1SAM|25|15|а эти люди очень добры к нам, не обижали нас, и ничего не пропало у нас во все время, когда мы ходили с ними, быв в поле;
1SAM|25|16|они были для нас оградою и днем и ночью во все время, когда мы пасли стада вблизи их;
1SAM|25|17|итак подумай и посмотри, что делать; ибо неминуемо угрожает беда господину нашему и всему дому его, а он – человек злой, нельзя говорить с ним.
1SAM|25|18|Тогда Авигея поспешно взяла двести хлебов, и два меха с вином, и пять овец приготовленных, и пять мер сушеных зерен, и сто связок изюму, и двести связок смокв, и навьючила на ослов,
1SAM|25|19|и сказала слугам своим: ступайте впереди меня, вот, я пойду за вами. А мужу своему Навалу ничего не сказала.
1SAM|25|20|Когда же она, сидя на осле, спускалась по извилинам горы, вот, навстречу ей идет Давид и люди его, и она встретилась с ними.
1SAM|25|21|И Давид сказал: да, напрасно я охранял в пустыне все имущество этого человека, и ничего не пропало из принадлежащего ему; он платит мне злом за добро;
1SAM|25|22|пусть то и то сделает Бог с врагами Давида, и еще больше сделает, если до рассвета утреннего из всего, что принадлежит Навалу, я оставлю мочащегося к стене.
1SAM|25|23|Когда Авигея увидела Давида, то поспешила сойти с осла и пала пред Давидом на лице свое и поклонилась до земли;
1SAM|25|24|и пала к ногам его и сказала: на мне грех, господин мой; позволь рабе твоей говорить в уши твои и послушай слов рабы твоей.
1SAM|25|25|Пусть господин мой не обращает внимания на этого злого человека, на Навала; ибо каково имя его, таков и он. Навал – имя его, и безумие его с ним. А я, раба твоя, не видела слуг господина моего, которых ты присылал.
1SAM|25|26|И ныне, господин мой, жив Господь и жива душа твоя, Господь не попустит тебе идти на пролитие крови и удержит руку твою от мщения, и ныне да будут, как Навал, враги твои и злоумышляющие против господина моего.
1SAM|25|27|Вот эти дары, которые принесла раба твоя господину моему, чтобы дать их отрокам, служащим господину моему.
1SAM|25|28|Прости вину рабы твоей; Господь непременно устроит господину моему дом твердый, ибо войны Господа ведет господин мой, и зло не найдется в тебе во всю жизнь твою.
1SAM|25|29|Если восстанет человек преследовать тебя и искать души твоей, то душа господина моего будет завязана в узле жизни у Господа Бога твоего, а душу врагов твоих бросит Он как бы пращею.
1SAM|25|30|И когда сделает Господь господину моему все, что говорил о тебе доброго, и поставит тебя вождем над Израилем,
1SAM|25|31|то не будет это сердцу господина моего огорчением и беспокойством, что не пролил напрасно крови и сберег себя от мщения. И Господь облагодетельствует господина моего, и вспомнишь рабу твою.
1SAM|25|32|И сказал Давид Авигее: благословен Господь Бог Израилев, Который послал тебя ныне навстречу мне,
1SAM|25|33|и благословен разум твой, и благословенна ты за то, что ты теперь не допустила меня идти на пролитие крови и отмстить за себя.
1SAM|25|34|Но, – жив Господь Бог Израилев, удержавший меня от нанесения зла тебе, – если бы ты не поспешила и не пришла навстречу мне, то до рассвета утреннего я не оставил бы Навалу мочащегося к стене.
1SAM|25|35|И принял Давид из рук ее то, что она принесла ему, и сказал ей: иди с миром в дом твой; вот, я послушался голоса твоего и почтил лице твое.
1SAM|25|36|И пришла Авигея к Навалу, и вот, у него пир в доме его, как пир царский, и сердце Навала было весело; он же был очень пьян; и не сказала ему ни слова, ни большого, ни малого, до утра.
1SAM|25|37|Утром же, когда Навал отрезвился, жена его рассказала ему об этом, и замерло в нем сердце его, и стал он, как камень.
1SAM|25|38|Дней через десять поразил Господь Навала, и он умер.
1SAM|25|39|И услышал Давид, что Навал умер, и сказал: благословен Господь, воздавший за посрамление, нанесенное мне Навалом, и сохранивший раба Своего от зла; Господь обратил злобу Навала на его же голову. И послал Давид сказать Авигее, что он берет ее себе в жену.
1SAM|25|40|И пришли слуги Давидовы к Авигее на Кармил и сказали ей так: Давид послал нас к тебе, чтобы взять тебя ему в жену.
1SAM|25|41|Она встала и поклонилась лицем до земли и сказала: вот, раба твоя [готова] быть служанкою, чтобы омывать ноги слуг господина моего.
1SAM|25|42|И собралась Авигея поспешно и села на осла, и пять служанок сопровождали ее; и пошла она за послами Давида и сделалась его женою.
1SAM|25|43|И Ахиноаму из Изрееля взял Давид, и обе они были его женами.
1SAM|25|44|Саул же отдал дочь свою Мелхолу, жену Давидову, Фалтию, сыну Лаиша, что из Галлима.
1SAM|26|1|Пришли Зифеи к Саулу в Гиву и сказали: вот, Давид скрывается у нас на холме Гахила, что направо от Иесимона.
1SAM|26|2|И встал Саул и спустился в пустыню Зиф, и с ним три тысячи отборных мужей Израильских, чтоб искать Давида в пустыне Зиф.
1SAM|26|3|И расположился Саул на холме Гахила, что направо от Иесимона, при дороге; Давид же находился в пустыне и видел, что Саул шел за ним в пустыню;
1SAM|26|4|и послал Давид соглядатаев и узнал, что Саул действительно пришел.
1SAM|26|5|И встал Давид, и пошел к месту, на котором Саул расположился станом, и увидел Давид место, где спал Саул и Авенир, сын Ниров, военачальник его. Саул же спал в шатре, а народ расположился вокруг него.
1SAM|26|6|И обратился Давид и сказал Ахимелеху Хеттеянину и Авессе, сыну Саруину, брату Иоава, говоря: кто пойдет со мною к Саулу в стан? И отвечал Авесса: я пойду с тобою.
1SAM|26|7|И пришел Давид с Авессою к людям [Сауловым] ночью; и вот, Саул лежит, спит в шатре, и копье его воткнуто в землю у изголовья его; Авенир же и народ лежат вокруг него.
1SAM|26|8|Авесса сказал Давиду: предал Бог ныне врага твоего в руки твои; итак позволь, я пригвожду его копьем к земле одним ударом и не повторю [удара].
1SAM|26|9|Но Давид сказал Авессе: не убивай его; ибо кто, подняв руку на помазанника Господня, останется ненаказанным?
1SAM|26|10|И сказал Давид: жив Господь! пусть поразит его Господь, или придет день его, и он умрет, или пойдет на войну и погибнет; меня же да не попустит Господь поднять руку мою на помазанника Господня;
1SAM|26|11|а возьми его копье, которое у изголовья его, и сосуд с водою, и пойдем к себе.
1SAM|26|12|И взял Давид копье и сосуд с водою у изголовья Саула, и пошли они к себе; и никто не видел, и никто не знал, и никто не проснулся, но все спали, ибо сон от Господа напал на них.
1SAM|26|13|И перешел Давид на другую сторону и стал на вершине горы вдали; большое расстояние [было] между ними.
1SAM|26|14|И воззвал Давид к народу и Авениру, сыну Нирову, говоря: отвечай, Авенир. И отвечал Авенир и сказал: кто ты, что кричишь и [беспокоишь] царя?
1SAM|26|15|И сказал Давид Авениру: не муж ли ты, и кто равен тебе в Израиле? Для чего же ты не бережешь господина твоего, царя? ибо приходил некто из народа, чтобы погубить царя, господина твоего.
1SAM|26|16|Нехорошо ты это делаешь; жив Господь! вы достойны смерти за то, что не бережете господина вашего, помазанника Господня. Посмотри, где копье царя и сосуд с водою, что [были] у изголовья его?
1SAM|26|17|И узнал Саул голос Давида и сказал: твой ли это голос, сын мой Давид? И сказал Давид: мой голос, господин мой, царь.
1SAM|26|18|И сказал [еще]: за что господин мой преследует раба своего? что я сделал? какое зло в руке моей?
1SAM|26|19|И ныне пусть выслушает господин мой, царь, слова раба своего: если Господь возбудил тебя против меня, то да будет это от тебя благовонною жертвою; если же – сыны человеческие, то прокляты они пред Господом, ибо они изгнали меня ныне, чтобы не принадлежать мне к наследию Господа, говоря: "ступай, служи богам чужим".
1SAM|26|20|Да не прольется же кровь моя на землю пред лицем Господа; ибо царь Израилев вышел искать одну блоху, как гоняются за куропаткою по горам.
1SAM|26|21|И сказал Саул: согрешил я; возвратись, сын мой Давид, ибо я не буду больше делать тебе зла, потому что душа моя была дорога ныне в глазах твоих; безумно поступал я и очень много погрешал.
1SAM|26|22|И отвечал Давид и сказал: вот копье царя; пусть один из отроков придет и возьмет его;
1SAM|26|23|и да воздаст Господь каждому по правде его и по истине его, так как Господь предавал тебя в руки [мои], но я не захотел поднять руки моей на помазанника Господня;
1SAM|26|24|и пусть, как драгоценна была жизнь твоя ныне в глазах моих, так ценится моя жизнь в очах Господа, и да избавит меня от всякой беды!
1SAM|26|25|И сказал Саул Давиду: благословен ты, сын мой Давид; и дело сделаешь, и превозмочь превозможешь. И пошел Давид своим путем, а Саул возвратился в свое место.
1SAM|27|1|И сказал Давид в сердце своем: когда–нибудь попаду я в руки Саула, и нет для меня ничего лучшего, как убежать в землю Филистимскую; и отстанет от меня Саул [и не будет] искать меня более по всем пределам Израильским, и я спасусь от руки его.
1SAM|27|2|И встал Давид, и отправился сам и шестьсот мужей, бывших с ним, к Анхусу, сыну Маоха, царю Гефскому.
1SAM|27|3|И жил Давид у Анхуса в Гефе, сам и люди его, каждый с семейством своим, Давид и обе жены его – Ахиноама Изреелитянка и Авигея, [бывшая] жена Навала, Кармилитянка.
1SAM|27|4|И донесли Саулу, что Давид убежал в Геф, и не стал он более искать его.
1SAM|27|5|И сказал Давид Анхусу: если я приобрел благоволение в глазах твоих, то пусть дано будет мне место в одном из малых городов, и я буду жить там; для чего рабу твоему жить в царском городе вместе с тобою?
1SAM|27|6|Тогда дал ему Анхус Секелаг, посему Секелаг и остался за царями Иудейскими доныне.
1SAM|27|7|Всего времени, какое прожил Давид в стране Филистимской, было год и четыре месяца.
1SAM|27|8|И выходил Давид с людьми своими и нападал на Гессурян и Гирзеян и Амаликитян, которые издавна населяли эту страну до Сура и даже до земли Египетской.
1SAM|27|9|И опустошал Давид ту страну, и не оставлял в живых ни мужчины, ни женщины, и забирал овец, и волов, и ослов, и верблюдов, и одежду; и возвращался, и приходил к Анхусу.
1SAM|27|10|И сказал Анхус Давиду: на кого нападали ныне? Давид сказал: на полуденную страну Иудеи и на полуденную страну Иерахмеела и на полуденную страну Кенеи.
1SAM|27|11|И не оставлял Давид в живых ни мужчины, ни женщины, и не приводил в Геф, говоря: они могут донести на нас и сказать: "так поступил Давид, и таков образ действий его во все время пребывания в стране Филистимской".
1SAM|27|12|И доверился Анхус Давиду, говоря: он опротивел народу своему Израилю и будет слугою моим вовек.
1SAM|28|1|В то время Филистимляне собрали войска свои для войны, чтобы воевать с Израилем. И сказал Анхус Давиду: да будет тебе известно, что ты пойдешь со мною в ополчение, ты и люди твои.
1SAM|28|2|И сказал Давид Анхусу: ныне ты узнаешь, что сделает раб твой. И сказал Анхус Давиду: за то я сделаю тебя хранителем головы моей на все время.
1SAM|28|3|И умер Самуил, и оплакивали его все Израильтяне и погребли его в Раме, в городе его. Саул же изгнал волшебников и гадателей из страны.
1SAM|28|4|И собрались Филистимляне и пошли и стали станом в Сонаме; собрал и Саул весь народ Израильский, и стали станом на Гелвуе.
1SAM|28|5|И увидел Саул стан Филистимский и испугался, и крепко дрогнуло сердце его.
1SAM|28|6|И вопросил Саул Господа; но Господь не отвечал ему ни во сне, ни чрез урим, ни чрез пророков.
1SAM|28|7|Тогда Саул сказал слугам своим: сыщите мне женщину волшебницу, и я пойду к ней и спрошу ее. И отвечали ему слуги его: здесь в Аэндоре есть женщина волшебница.
1SAM|28|8|И снял с себя Саул одежды свои и надел другие, и пошел сам и два человека с ним, и пришли они к женщине ночью. И сказал ей [Саул]: прошу тебя, поворожи мне и выведи мне, о ком я скажу тебе.
1SAM|28|9|Но женщина отвечала ему: ты знаешь, что сделал Саул, как выгнал он из страны волшебников и гадателей; для чего же ты расставляешь сеть душе моей на погибель мне?
1SAM|28|10|И поклялся ей Саул Господом, говоря: жив Господь! не будет тебе беды за это дело.
1SAM|28|11|Тогда женщина спросила: кого же вывесть тебе? И отвечал он: Самуила выведи мне.
1SAM|28|12|И увидела женщина Самуила и громко вскрикнула; и обратилась женщина к Саулу, говоря: зачем ты обманул меня? ты – Саул.
1SAM|28|13|И сказал ей царь: не бойся; что ты видишь? И отвечала женщина: вижу как бы бога, выходящего из земли.
1SAM|28|14|Какой он видом? – спросил у нее [Саул]. Она сказала: выходит из земли муж престарелый, одетый в длинную одежду. Тогда узнал Саул, что это Самуил, и пал лицем на землю и поклонился.
1SAM|28|15|И сказал Самуил Саулу: для чего ты тревожишь меня, чтобы я вышел? И отвечал Саул: тяжело мне очень; Филистимляне воюют против меня, а Бог отступил от меня и более не отвечает мне ни чрез пророков, ни во сне; потому я вызвал тебя, чтобы ты научил меня, что мне делать.
1SAM|28|16|И сказал Самуил: для чего же ты спрашиваешь меня, когда Господь отступил от тебя и сделался врагом твоим?
1SAM|28|17|Господь сделает то, что говорил чрез меня; отнимет Господь царство из рук твоих и отдаст его ближнему твоему, Давиду.
1SAM|28|18|Так как ты не послушал гласа Господня и не выполнил ярости гнева Его на Амалика, то Господь и делает это над тобою ныне.
1SAM|28|19|И предаст Господь Израиля вместе с тобою в руки Филистимлян: завтра ты и сыны твои [будете] со мною, и стан Израильский предаст Господь в руки Филистимлян.
1SAM|28|20|Тогда Саул вдруг пал всем телом своим на землю, ибо сильно испугался слов Самуила; притом и силы не стало в нем, ибо он не ел хлеба весь тот день и всю ночь.
1SAM|28|21|И подошла женщина та к Саулу, и увидела, что он очень испугался, и сказала: вот, раба твоя послушалась голоса твоего и подвергала жизнь свою опасности и исполнила приказание, которое ты дал мне;
1SAM|28|22|теперь прошу, послушайся и ты голоса рабы твоей: я предложу тебе кусок хлеба, поешь, и будет в тебе крепость, когда пойдешь в путь.
1SAM|28|23|Но он отказался и сказал: не буду есть. И стали уговаривать его слуги его, а также и женщина; и он послушался голоса их, и встал с земли и сел на ложе.
1SAM|28|24|У женщины же был в доме откормленный теленок, и она поспешила заколоть его и, взяв муки, замесила и испекла опресноки,
1SAM|28|25|и предложила Саулу и слугам его, и они поели, и встали, и ушли в ту же ночь.
1SAM|29|1|И собрали Филистимляне все ополчения свои в Афеке, а Израильтяне расположились станом у источника, что в Изрееле.
1SAM|29|2|Князья Филистимские шли с сотнями и тысячами, Давид же и люди его шли позади с Анхусом.
1SAM|29|3|И говорили князья Филистимские: это что за Евреи? Анхус отвечал князьям Филистимским: разве не знаете, что это Давид, раб Саула, царя Израильского? он при мне уже более года, и я не нашел в нем ничего худого со времени его прихода до сего дня.
1SAM|29|4|И вознегодовали на него князья Филистимские, и сказали ему князья Филистимские: отпусти ты этого человека, пусть он сидит в своем месте, которое ты ему назначил, чтоб он не шел с нами на войну и не сделался противником нашим на войне. Чем он может умилостивить господина своего, как не головами сих мужей?
1SAM|29|5|Не тот ли это Давид, которому пели в хороводах, говоря: "Саул поразил тысячи, а Давид – десятки тысяч"?
1SAM|29|6|И призвал Анхус Давида и сказал ему: жив Господь! ты честен, и глазам моим приятно было бы, чтобы ты выходил и входил со мною в ополчении; ибо я не заметил в тебе худого со времени прихода твоего ко мне до сего дня; но в глазах князей ты не хорош.
1SAM|29|7|Итак, возвратись теперь, и иди с миром и не раздражай князей Филистимских.
1SAM|29|8|Но Давид сказал Анхусу: что я сделал, и что ты нашел в рабе твоем с того времени, как я пред лицем твоим, и до сего дня, почему бы мне не идти и не воевать с врагами господина моего, царя?
1SAM|29|9|И отвечал Анхус Давиду: будь уверен, что в моих глазах ты хорош, как Ангел Божий; но князья Филистимские сказали: "пусть он не идет с нами на войну".
1SAM|29|10|Итак встань утром, ты и рабы господина твоего, которые пришли с тобою; и встаньте поутру, и когда светло будет, идите.
1SAM|29|11|И встал Давид, сам и люди его, чтобы идти утром и возвратиться в землю Филистимскую. А Филистимляне пошли [на войну] в Изреель.
1SAM|30|1|В третий день после того, как Давид и люди его пошли в Секелаг, Амаликитяне напали с юга на Секелаг и взяли Секелаг и сожгли его огнем,
1SAM|30|2|а женщин [и всех], бывших в нем, от малого до большого, не умертвили, но увели в плен, и ушли своим путем.
1SAM|30|3|И пришел Давид и люди его к городу, и вот, он сожжен огнем, а жены их и сыновья их и дочери их взяты в плен.
1SAM|30|4|И поднял Давид и народ, бывший с ним, вопль, и плакали, доколе не стало в них силы плакать.
1SAM|30|5|Взяты были в плен и обе жены Давида: Ахиноама Изреелитянка и Авигея, [бывшая] жена Навала, Кармилитянка.
1SAM|30|6|Давид сильно был смущен, так как народ хотел побить его камнями; ибо скорбел душею весь народ, каждый о сыновьях своих и дочерях своих.
1SAM|30|7|Но Давид укрепился [надеждою] на Господа Бога своего, и сказал Давид Авиафару священнику, сыну Ахимелехову: принеси мне ефод. И принес Авиафар ефод к Давиду.
1SAM|30|8|И вопросил Давид Господа, говоря: преследовать ли мне это полчище, и догоню ли их? И сказано ему: преследуй, догонишь и отнимешь.
1SAM|30|9|И пошел Давид сам и шестьсот мужей, бывших с ним; и пришли к потоку Восор и усталые остановились там.
1SAM|30|10|И преследовал Давид сам и четыреста человек; двести же человек остановились, потому что были не в силах перейти поток Восорский.
1SAM|30|11|И нашли Египтянина в поле, и привели его к Давиду, и дали ему хлеба, и он ел, и напоили его водою;
1SAM|30|12|и дали ему часть связки смокв и две связки изюму, и он ел и укрепился, ибо он не ел хлеба и не пил воды три дня и три ночи.
1SAM|30|13|И сказал ему Давид: чей ты и откуда ты? И сказал он: я – отрок Египтянина, раб одного Амаликитянина, и бросил меня господин мой, ибо уже три дня, как я заболел;
1SAM|30|14|мы вторгались в полуденную часть Керети и в область Иудину и в полуденную часть Халева, а Секелаг сожгли огнем.
1SAM|30|15|И сказал ему Давид: доведешь ли меня до этого полчища? И сказал он: поклянись мне Богом, что ты не умертвишь меня и не предашь меня в руки господина моего, и я доведу тебя до этого полчища.
1SAM|30|16|и он повел его; и вот, [Амаликитяне], рассыпавшись по всей той стране, едят и пьют и празднуют по причине великой добычи, которую они взяли из земли Филистимской и из земли Иудейской.
1SAM|30|17|и поражал их Давид от сумерек до вечера другого дня, и никто из них не спасся, кроме четырехсот юношей, которые сели на верблюдов и убежали.
1SAM|30|18|И отнял Давид все, что взяли Амаликитяне, и обеих жен своих отнял Давид.
1SAM|30|19|И не пропало у них ничего, ни малого, ни большого, ни из сыновей, ни из дочерей, ни из добычи, ни из всего, что [Амаликитяне] взяли у них; все возвратил Давид,
1SAM|30|20|и взял Давид весь мелкий и крупный скот, и гнали его пред своим скотом и говорили: это – добыча Давида.
1SAM|30|21|И пришел Давид к тем двум стам человек, которые не были в силах идти за ним, и [которых] он оставил у потока Восор, и вышли они навстречу Давиду и навстречу людям, бывшим с ним. И подошел Давид к этим людям и приветствовал их.
1SAM|30|22|Тогда злые и негодные из людей, ходивших с Давидом, стали говорить: за то, что они не ходили с нами, не дадим им из добычи, которую мы отняли; пусть каждый возьмет только свою жену и детей и идет.
1SAM|30|23|Но Давид сказал: не делайте так, братья мои, после того, как Господь дал нам это и сохранил нас и предал в руки наши полчище, приходившее против нас.
1SAM|30|24|И кто послушает вас в этом деле? Какова часть ходившим на войну, такова часть должна быть и оставшимся при обозе: на всех должно разделить.
1SAM|30|25|Так было с этого времени и после; и поставил он это в закон и в правило для Израиля до сего дня.
1SAM|30|26|И пришел Давид в Секелаг и послал из добычи к старейшинам Иудиным, друзьям своим, говоря: "вот вам подарок из добычи, [взятой] у врагов Господних", –
1SAM|30|27|тем, которые в Вефиле, и в Рамофе южном, и в Иаттире.
1SAM|30|28|и в Ароере, и в Шифмофе, и в Естемоа,
1SAM|30|29|и в Рахале, и в городах Иерахмеельских, и в городах Кенейских,
1SAM|30|30|и в Хорме, и в Хорашане, и в Атахе,
1SAM|30|31|и в Хевроне, и во всех местах, где ходил Давид сам и люди его.
1SAM|31|1|Филистимляне же воевали с Израильтянами, и побежали мужи Израильские от Филистимлян и пали пораженные на горе Гелвуе.
1SAM|31|2|И догнали Филистимляне Саула и сыновей его, и убили Филистимляне Ионафана, и Аминадава, и Малхисуа, сыновей Саула.
1SAM|31|3|И битва против Саула сделалась жестокая, и стрелки из луков поражали его, и он очень изранен был стрелками.
1SAM|31|4|И сказал Саул оруженосцу своему: обнажи твой меч и заколи меня им, чтобы не пришли эти необрезанные и не убили меня и не издевались надо мною. Но оруженосец не хотел, ибо очень боялся. Тогда Саул взял меч свой и пал на него.
1SAM|31|5|Оруженосец его, увидев, что Саул умер, и сам пал на свой меч и умер с ним.
1SAM|31|6|Так умер в тот день Саул и три сына его, и оруженосец его, а также и все люди его вместе.
1SAM|31|7|Израильтяне, жившие на стороне долины и за Иорданом, видя, что люди Израилевы побежали и что умер Саул и сыновья его, оставили города свои и бежали, а Филистимляне пришли и засели в них.
1SAM|31|8|На другой день Филистимляне пришли грабить убитых, и нашли Саула и трех сыновей его, павших на горе Гелвуйской.
1SAM|31|9|И отсекли ему голову, и сняли с него оружие и послали по всей земле Филистимской, чтобы возвестить о сем в капищах идолов своих и народу;
1SAM|31|10|и положили оружие его в капище Астарты, а тело его повесили на стене Беф–Сана.
1SAM|31|11|И услышали жители Иависа Галаадского о том, как поступили Филистимляне с Саулом,
1SAM|31|12|и поднялись все люди сильные, и шли всю ночь, и взяли тело Саула и тела сыновей его со стены Беф–Сана, и пришли в Иавис, и сожгли их там;
1SAM|31|13|и взяли кости их, и погребли под дубом в Иависе, и постились семь дней.
