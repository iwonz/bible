HEB|1|1|God, who at sundry times and in divers manners spake in time past unto the fathers by the prophets,
HEB|1|2|Hath in these last days spoken unto us by his Son, whom he hath appointed heir of all things, by whom also he made the worlds;
HEB|1|3|Who being the brightness of his glory, and the express image of his person, and upholding all things by the word of his power, when he had by himself purged our sins, sat down on the right hand of the Majesty on high:
HEB|1|4|Being made so much better than the angels, as he hath by inheritance obtained a more excellent name than they.
HEB|1|5|For unto which of the angels said he at any time, Thou art my Son, this day have I begotten thee? And again, I will be to him a Father, and he shall be to me a Son?
HEB|1|6|And again, when he bringeth in the firstbegotten into the world, he saith, And let all the angels of God worship him.
HEB|1|7|And of the angels he saith, Who maketh his angels spirits, and his ministers a flame of fire.
HEB|1|8|But unto the Son he saith, Thy throne, O God, is for ever and ever: a sceptre of righteousness is the sceptre of thy kingdom.
HEB|1|9|Thou hast loved righteousness, and hated iniquity; therefore God, even thy God, hath anointed thee with the oil of gladness above thy fellows.
HEB|1|10|And, Thou, Lord, in the beginning hast laid the foundation of the earth; and the heavens are the works of thine hands:
HEB|1|11|They shall perish; but thou remainest; and they all shall wax old as doth a garment;
HEB|1|12|And as a vesture shalt thou fold them up, and they shall be changed: but thou art the same, and thy years shall not fail.
HEB|1|13|But to which of the angels said he at any time, Sit on my right hand, until I make thine enemies thy footstool?
HEB|1|14|Are they not all ministering spirits, sent forth to minister for them who shall be heirs of salvation?
HEB|2|1|Therefore we ought to give the more earnest heed to the things which we have heard, lest at any time we should let them slip.
HEB|2|2|For if the word spoken by angels was stedfast, and every transgression and disobedience received a just recompence of reward;
HEB|2|3|How shall we escape, if we neglect so great salvation; which at the first began to be spoken by the Lord, and was confirmed unto us by them that heard him;
HEB|2|4|God also bearing them witness, both with signs and wonders, and with divers miracles, and gifts of the Holy Ghost, according to his own will?
HEB|2|5|For unto the angels hath he not put in subjection the world to come, whereof we speak.
HEB|2|6|But one in a certain place testified, saying, What is man, that thou art mindful of him? or the son of man that thou visitest him?
HEB|2|7|Thou madest him a little lower than the angels; thou crownedst him with glory and honour, and didst set him over the works of thy hands:
HEB|2|8|Thou hast put all things in subjection under his feet. For in that he put all in subjection under him, he left nothing that is not put under him. But now we see not yet all things put under him.
HEB|2|9|But we see Jesus, who was made a little lower than the angels for the suffering of death, crowned with glory and honour; that he by the grace of God should taste death for every man.
HEB|2|10|For it became him, for whom are all things, and by whom are all things, in bringing many sons unto glory, to make the captain of their salvation perfect through sufferings.
HEB|2|11|For both he that sanctifieth and they who are sanctified are all of one: for which cause he is not ashamed to call them brethren,
HEB|2|12|Saying, I will declare thy name unto my brethren, in the midst of the church will I sing praise unto thee.
HEB|2|13|And again, I will put my trust in him. And again, Behold I and the children which God hath given me.
HEB|2|14|Forasmuch then as the children are partakers of flesh and blood, he also himself likewise took part of the same; that through death he might destroy him that had the power of death, that is, the devil;
HEB|2|15|And deliver them who through fear of death were all their lifetime subject to bondage.
HEB|2|16|For verily he took not on him the nature of angels; but he took on him the seed of Abraham.
HEB|2|17|Wherefore in all things it behoved him to be made like unto his brethren, that he might be a merciful and faithful high priest in things pertaining to God, to make reconciliation for the sins of the people.
HEB|2|18|For in that he himself hath suffered being tempted, he is able to succour them that are tempted.
HEB|3|1|Wherefore, holy brethren, partakers of the heavenly calling, consider the Apostle and High Priest of our profession, Christ Jesus;
HEB|3|2|Who was faithful to him that appointed him, as also Moses was faithful in all his house.
HEB|3|3|For this man was counted worthy of more glory than Moses, inasmuch as he who hath builded the house hath more honour than the house.
HEB|3|4|For every house is builded by some man; but he that built all things is God.
HEB|3|5|And Moses verily was faithful in all his house, as a servant, for a testimony of those things which were to be spoken after;
HEB|3|6|But Christ as a son over his own house; whose house are we, if we hold fast the confidence and the rejoicing of the hope firm unto the end.
HEB|3|7|Wherefore (as the Holy Ghost saith, To day if ye will hear his voice,
HEB|3|8|Harden not your hearts, as in the provocation, in the day of temptation in the wilderness:
HEB|3|9|When your fathers tempted me, proved me, and saw my works forty years.
HEB|3|10|Wherefore I was grieved with that generation, and said, They do alway err in their heart; and they have not known my ways.
HEB|3|11|So I sware in my wrath, They shall not enter into my rest.)
HEB|3|12|Take heed, brethren, lest there be in any of you an evil heart of unbelief, in departing from the living God.
HEB|3|13|But exhort one another daily, while it is called To day; lest any of you be hardened through the deceitfulness of sin.
HEB|3|14|For we are made partakers of Christ, if we hold the beginning of our confidence stedfast unto the end;
HEB|3|15|While it is said, To day if ye will hear his voice, harden not your hearts, as in the provocation.
HEB|3|16|For some, when they had heard, did provoke: howbeit not all that came out of Egypt by Moses.
HEB|3|17|But with whom was he grieved forty years? was it not with them that had sinned, whose carcases fell in the wilderness?
HEB|3|18|And to whom sware he that they should not enter into his rest, but to them that believed not?
HEB|3|19|So we see that they could not enter in because of unbelief.
HEB|4|1|Let us therefore fear, lest, a promise being left us of entering into his rest, any of you should seem to come short of it.
HEB|4|2|For unto us was the gospel preached, as well as unto them: but the word preached did not profit them, not being mixed with faith in them that heard it.
HEB|4|3|For we which have believed do enter into rest, as he said, As I have sworn in my wrath, if they shall enter into my rest: although the works were finished from the foundation of the world.
HEB|4|4|For he spake in a certain place of the seventh day on this wise, And God did rest the seventh day from all his works.
HEB|4|5|And in this place again, If they shall enter into my rest.
HEB|4|6|Seeing therefore it remaineth that some must enter therein, and they to whom it was first preached entered not in because of unbelief:
HEB|4|7|Again, he limiteth a certain day, saying in David, To day, after so long a time; as it is said, To day if ye will hear his voice, harden not your hearts.
HEB|4|8|For if Joshua had given them rest, then would he not afterward have spoken of another day.
HEB|4|9|There remaineth therefore a rest to the people of God.
HEB|4|10|For he that is entered into his rest, he also hath ceased from his own works, as God did from his.
HEB|4|11|Let us labour therefore to enter into that rest, lest any man fall after the same example of unbelief.
HEB|4|12|For the word of God is quick, and powerful, and sharper than any twoedged sword, piercing even to the dividing asunder of soul and spirit, and of the joints and marrow, and is a discerner of the thoughts and intents of the heart.
HEB|4|13|Neither is there any creature that is not manifest in his sight: but all things are naked and opened unto the eyes of him with whom we have to do.
HEB|4|14|Seeing then that we have a great high priest, that is passed into the heavens, Jesus the Son of God, let us hold fast our profession.
HEB|4|15|For we have not an high priest which cannot be touched with the feeling of our infirmities; but was in all points tempted like as we are, yet without sin.
HEB|4|16|Let us therefore come boldly unto the throne of grace, that we may obtain mercy, and find grace to help in time of need.
HEB|5|1|For every high priest taken from among men is ordained for men in things pertaining to God, that he may offer both gifts and sacrifices for sins:
HEB|5|2|Who can have compassion on the ignorant, and on them that are out of the way; for that he himself also is compassed with infirmity.
HEB|5|3|And by reason hereof he ought, as for the people, so also for himself, to offer for sins.
HEB|5|4|And no man taketh this honour unto himself, but he that is called of God, as was Aaron.
HEB|5|5|So also Christ glorified not himself to be made an high priest; but he that said unto him, Thou art my Son, to day have I begotten thee.
HEB|5|6|As he saith also in another place, Thou art a priest for ever after the order of Melchisedec.
HEB|5|7|Who in the days of his flesh, when he had offered up prayers and supplications with strong crying and tears unto him that was able to save him from death, and was heard in that he feared;
HEB|5|8|Though he were a Son, yet learned he obedience by the things which he suffered;
HEB|5|9|And being made perfect, he became the author of eternal salvation unto all them that obey him;
HEB|5|10|Called of God an high priest after the order of Melchisedec.
HEB|5|11|Of whom we have many things to say, and hard to be uttered, seeing ye are dull of hearing.
HEB|5|12|For when for the time ye ought to be teachers, ye have need that one teach you again which be the first principles of the oracles of God; and are become such as have need of milk, and not of strong meat.
HEB|5|13|For every one that useth milk is unskilful in the word of righteousness: for he is a babe.
HEB|5|14|But strong meat belongeth to them that are of full age, even those who by reason of use have their senses exercised to discern both good and evil.
HEB|6|1|Therefore leaving the principles of the doctrine of Christ, let us go on unto perfection; not laying again the foundation of repentance from dead works, and of faith toward God,
HEB|6|2|Of the doctrine of baptisms, and of laying on of hands, and of resurrection of the dead, and of eternal judgment.
HEB|6|3|And this will we do, if God permit.
HEB|6|4|For it is impossible for those who were once enlightened, and have tasted of the heavenly gift, and were made partakers of the Holy Ghost,
HEB|6|5|And have tasted the good word of God, and the powers of the world to come,
HEB|6|6|If they shall fall away, to renew them again unto repentance; seeing they crucify to themselves the Son of God afresh, and put him to an open shame.
HEB|6|7|For the earth which drinketh in the rain that cometh oft upon it, and bringeth forth herbs meet for them by whom it is dressed, receiveth blessing from God:
HEB|6|8|But that which beareth thorns and briers is rejected, and is nigh unto cursing; whose end is to be burned.
HEB|6|9|But, beloved, we are persuaded better things of you, and things that accompany salvation, though we thus speak.
HEB|6|10|For God is not unrighteous to forget your work and labour of love, which ye have shewed toward his name, in that ye have ministered to the saints, and do minister.
HEB|6|11|And we desire that every one of you do shew the same diligence to the full assurance of hope unto the end:
HEB|6|12|That ye be not slothful, but followers of them who through faith and patience inherit the promises.
HEB|6|13|For when God made promise to Abraham, because he could swear by no greater, he sware by himself,
HEB|6|14|Saying, Surely blessing I will bless thee, and multiplying I will multiply thee.
HEB|6|15|And so, after he had patiently endured, he obtained the promise.
HEB|6|16|For men verily swear by the greater: and an oath for confirmation is to them an end of all strife.
HEB|6|17|Wherein God, willing more abundantly to shew unto the heirs of promise the immutability of his counsel, confirmed it by an oath:
HEB|6|18|That by two immutable things, in which it was impossible for God to lie, we might have a strong consolation, who have fled for refuge to lay hold upon the hope set before us:
HEB|6|19|Which hope we have as an anchor of the soul, both sure and stedfast, and which entereth into that within the veil;
HEB|6|20|Whither the forerunner is for us entered, even Jesus, made an high priest for ever after the order of Melchisedec.
HEB|7|1|For this Melchisedec, king of Salem, priest of the most high God, who met Abraham returning from the slaughter of the kings, and blessed him;
HEB|7|2|To whom also Abraham gave a tenth part of all; first being by interpretation King of righteousness, and after that also King of Salem, which is, King of peace;
HEB|7|3|Without father, without mother, without descent, having neither beginning of days, nor end of life; but made like unto the Son of God; abideth a priest continually.
HEB|7|4|Now consider how great this man was, unto whom even the patriarch Abraham gave the tenth of the spoils.
HEB|7|5|And verily they that are of the sons of Levi, who receive the office of the priesthood, have a commandment to take tithes of the people according to the law, that is, of their brethren, though they come out of the loins of Abraham:
HEB|7|6|But he whose descent is not counted from them received tithes of Abraham, and blessed him that had the promises.
HEB|7|7|And without all contradiction the less is blessed of the better.
HEB|7|8|And here men that die receive tithes; but there he receiveth them, of whom it is witnessed that he liveth.
HEB|7|9|And as I may so say, Levi also, who receiveth tithes, payed tithes in Abraham.
HEB|7|10|For he was yet in the loins of his father, when Melchisedec met him.
HEB|7|11|If therefore perfection were by the Levitical priesthood, (for under it the people received the law,) what further need was there that another priest should rise after the order of Melchisedec, and not be called after the order of Aaron?
HEB|7|12|For the priesthood being changed, there is made of necessity a change also of the law.
HEB|7|13|For he of whom these things are spoken pertaineth to another tribe, of which no man gave attendance at the altar.
HEB|7|14|For it is evident that our Lord sprang out of Juda; of which tribe Moses spake nothing concerning priesthood.
HEB|7|15|And it is yet far more evident: for that after the similitude of Melchisedec there ariseth another priest,
HEB|7|16|Who is made, not after the law of a carnal commandment, but after the power of an endless life.
HEB|7|17|For he testifieth, Thou art a priest for ever after the order of Melchisedec.
HEB|7|18|For there is verily a disannulling of the commandment going before for the weakness and unprofitableness thereof.
HEB|7|19|For the law made nothing perfect, but the bringing in of a better hope did; by the which we draw nigh unto God.
HEB|7|20|And inasmuch as not without an oath he was made priest:
HEB|7|21|(For those priests were made without an oath; but this with an oath by him that said unto him, The Lord sware and will not repent, Thou art a priest for ever after the order of Melchisedec:)
HEB|7|22|By so much was Jesus made a surety of a better testament.
HEB|7|23|And they truly were many priests, because they were not suffered to continue by reason of death:
HEB|7|24|But this man, because he continueth ever, hath an unchangeable priesthood.
HEB|7|25|Wherefore he is able also to save them to the uttermost that come unto God by him, seeing he ever liveth to make intercession for them.
HEB|7|26|For such an high priest became us, who is holy, harmless, undefiled, separate from sinners, and made higher than the heavens;
HEB|7|27|Who needeth not daily, as those high priests, to offer up sacrifice, first for his own sins, and then for the people's: for this he did once, when he offered up himself.
HEB|7|28|For the law maketh men high priests which have infirmity; but the word of the oath, which was since the law, maketh the Son, who is consecrated for evermore.
HEB|8|1|Now of the things which we have spoken this is the sum: We have such an high priest, who is set on the right hand of the throne of the Majesty in the heavens;
HEB|8|2|A minister of the sanctuary, and of the true tabernacle, which the Lord pitched, and not man.
HEB|8|3|For every high priest is ordained to offer gifts and sacrifices: wherefore it is of necessity that this man have somewhat also to offer.
HEB|8|4|For if he were on earth, he should not be a priest, seeing that there are priests that offer gifts according to the law:
HEB|8|5|Who serve unto the example and shadow of heavenly things, as Moses was admonished of God when he was about to make the tabernacle: for, See, saith he, that thou make all things according to the pattern shewed to thee in the mount.
HEB|8|6|But now hath he obtained a more excellent ministry, by how much also he is the mediator of a better covenant, which was established upon better promises.
HEB|8|7|For if that first covenant had been faultless, then should no place have been sought for the second.
HEB|8|8|For finding fault with them, he saith, Behold, the days come, saith the Lord, when I will make a new covenant with the house of Israel and with the house of Judah:
HEB|8|9|Not according to the covenant that I made with their fathers in the day when I took them by the hand to lead them out of the land of Egypt; because they continued not in my covenant, and I regarded them not, saith the Lord.
HEB|8|10|For this is the covenant that I will make with the house of Israel after those days, saith the Lord; I will put my laws into their mind, and write them in their hearts: and I will be to them a God, and they shall be to me a people:
HEB|8|11|And they shall not teach every man his neighbour, and every man his brother, saying, Know the Lord: for all shall know me, from the least to the greatest.
HEB|8|12|For I will be merciful to their unrighteousness, and their sins and their iniquities will I remember no more.
HEB|8|13|In that he saith, A new covenant, he hath made the first old. Now that which decayeth and waxeth old is ready to vanish away.
HEB|9|1|Then verily the first covenant had also ordinances of divine service, and a worldly sanctuary.
HEB|9|2|For there was a tabernacle made; the first, wherein was the candlestick, and the table, and the shewbread; which is called the sanctuary.
HEB|9|3|And after the second veil, the tabernacle which is called the Holiest of all;
HEB|9|4|Which had the golden censer, and the ark of the covenant overlaid round about with gold, wherein was the golden pot that had manna, and Aaron's rod that budded, and the tables of the covenant;
HEB|9|5|And over it the cherubims of glory shadowing the mercyseat; of which we cannot now speak particularly.
HEB|9|6|Now when these things were thus ordained, the priests went always into the first tabernacle, accomplishing the service of God.
HEB|9|7|But into the second went the high priest alone once every year, not without blood, which he offered for himself, and for the errors of the people:
HEB|9|8|The Holy Ghost this signifying, that the way into the holiest of all was not yet made manifest, while as the first tabernacle was yet standing:
HEB|9|9|Which was a figure for the time then present, in which were offered both gifts and sacrifices, that could not make him that did the service perfect, as pertaining to the conscience;
HEB|9|10|Which stood only in meats and drinks, and divers washings, and carnal ordinances, imposed on them until the time of reformation.
HEB|9|11|But Christ being come an high priest of good things to come, by a greater and more perfect tabernacle, not made with hands, that is to say, not of this building;
HEB|9|12|Neither by the blood of goats and calves, but by his own blood he entered in once into the holy place, having obtained eternal redemption for us.
HEB|9|13|For if the blood of bulls and of goats, and the ashes of an heifer sprinkling the unclean, sanctifieth to the purifying of the flesh:
HEB|9|14|How much more shall the blood of Christ, who through the eternal Spirit offered himself without spot to God, purge your conscience from dead works to serve the living God?
HEB|9|15|And for this cause he is the mediator of the new testament, that by means of death, for the redemption of the transgressions that were under the first testament, they which are called might receive the promise of eternal inheritance.
HEB|9|16|For where a testament is, there must also of necessity be the death of the testator.
HEB|9|17|For a testament is of force after men are dead: otherwise it is of no strength at all while the testator liveth.
HEB|9|18|Whereupon neither the first testament was dedicated without blood.
HEB|9|19|For when Moses had spoken every precept to all the people according to the law, he took the blood of calves and of goats, with water, and scarlet wool, and hyssop, and sprinkled both the book, and all the people,
HEB|9|20|Saying, This is the blood of the testament which God hath enjoined unto you.
HEB|9|21|Moreover he sprinkled with blood both the tabernacle, and all the vessels of the ministry.
HEB|9|22|And almost all things are by the law purged with blood; and without shedding of blood is no remission.
HEB|9|23|It was therefore necessary that the patterns of things in the heavens should be purified with these; but the heavenly things themselves with better sacrifices than these.
HEB|9|24|For Christ is not entered into the holy places made with hands, which are the figures of the true; but into heaven itself, now to appear in the presence of God for us:
HEB|9|25|Nor yet that he should offer himself often, as the high priest entereth into the holy place every year with blood of others;
HEB|9|26|For then must he often have suffered since the foundation of the world: but now once in the end of the world hath he appeared to put away sin by the sacrifice of himself.
HEB|9|27|And as it is appointed unto men once to die, but after this the judgment:
HEB|9|28|So Christ was once offered to bear the sins of many; and unto them that look for him shall he appear the second time without sin unto salvation.
HEB|10|1|For the law having a shadow of good things to come, and not the very image of the things, can never with those sacrifices which they offered year by year continually make the comers thereunto perfect.
HEB|10|2|For then would they not have ceased to be offered? because that the worshippers once purged should have had no more conscience of sins.
HEB|10|3|But in those sacrifices there is a remembrance again made of sins every year.
HEB|10|4|For it is not possible that the blood of bulls and of goats should take away sins.
HEB|10|5|Wherefore when he cometh into the world, he saith, Sacrifice and offering thou wouldest not, but a body hast thou prepared me:
HEB|10|6|In burnt offerings and sacrifices for sin thou hast had no pleasure.
HEB|10|7|Then said I, Lo, I come (in the volume of the book it is written of me,) to do thy will, O God.
HEB|10|8|Above when he said, Sacrifice and offering and burnt offerings and offering for sin thou wouldest not, neither hadst pleasure therein; which are offered by the law;
HEB|10|9|Then said he, Lo, I come to do thy will, O God. He taketh away the first, that he may establish the second.
HEB|10|10|By the which will we are sanctified through the offering of the body of Jesus Christ once for all.
HEB|10|11|And every priest standeth daily ministering and offering oftentimes the same sacrifices, which can never take away sins:
HEB|10|12|But this man, after he had offered one sacrifice for sins for ever, sat down on the right hand of God;
HEB|10|13|From henceforth expecting till his enemies be made his footstool.
HEB|10|14|For by one offering he hath perfected for ever them that are sanctified.
HEB|10|15|Whereof the Holy Ghost also is a witness to us: for after that he had said before,
HEB|10|16|This is the covenant that I will make with them after those days, saith the Lord, I will put my laws into their hearts, and in their minds will I write them;
HEB|10|17|And their sins and iniquities will I remember no more.
HEB|10|18|Now where remission of these is, there is no more offering for sin.
HEB|10|19|Having therefore, brethren, boldness to enter into the holiest by the blood of Jesus,
HEB|10|20|By a new and living way, which he hath consecrated for us, through the veil, that is to say, his flesh;
HEB|10|21|And having an high priest over the house of God;
HEB|10|22|Let us draw near with a true heart in full assurance of faith, having our hearts sprinkled from an evil conscience, and our bodies washed with pure water.
HEB|10|23|Let us hold fast the profession of our faith without wavering; (for he is faithful that promised;)
HEB|10|24|And let us consider one another to provoke unto love and to good works:
HEB|10|25|Not forsaking the assembling of ourselves together, as the manner of some is; but exhorting one another: and so much the more, as ye see the day approaching.
HEB|10|26|For if we sin wilfully after that we have received the knowledge of the truth, there remaineth no more sacrifice for sins,
HEB|10|27|But a certain fearful looking for of judgment and fiery indignation, which shall devour the adversaries.
HEB|10|28|He that despised Moses' law died without mercy under two or three witnesses:
HEB|10|29|Of how much sorer punishment, suppose ye, shall he be thought worthy, who hath trodden under foot the Son of God, and hath counted the blood of the covenant, wherewith he was sanctified, an unholy thing, and hath done despite unto the Spirit of grace?
HEB|10|30|For we know him that hath said, Vengeance belongeth unto me, I will recompense, saith the Lord. And again, The Lord shall judge his people.
HEB|10|31|It is a fearful thing to fall into the hands of the living God.
HEB|10|32|But call to remembrance the former days, in which, after ye were illuminated, ye endured a great fight of afflictions;
HEB|10|33|Partly, whilst ye were made a gazingstock both by reproaches and afflictions; and partly, whilst ye became companions of them that were so used.
HEB|10|34|For ye had compassion of me in my bonds, and took joyfully the spoiling of your goods, knowing in yourselves that ye have in heaven a better and an enduring substance.
HEB|10|35|Cast not away therefore your confidence, which hath great recompence of reward.
HEB|10|36|For ye have need of patience, that, after ye have done the will of God, ye might receive the promise.
HEB|10|37|For yet a little while, and he that shall come will come, and will not tarry.
HEB|10|38|Now the just shall live by faith: but if any man draw back, my soul shall have no pleasure in him.
HEB|10|39|But we are not of them who draw back unto perdition; but of them that believe to the saving of the soul.
HEB|11|1|Now faith is the substance of things hoped for, the evidence of things not seen.
HEB|11|2|For by it the elders obtained a good report.
HEB|11|3|Through faith we understand that the worlds were framed by the word of God, so that things which are seen were not made of things which do appear.
HEB|11|4|By faith Abel offered unto God a more excellent sacrifice than Cain, by which he obtained witness that he was righteous, God testifying of his gifts: and by it he being dead yet speaketh.
HEB|11|5|By faith Enoch was translated that he should not see death; and was not found, because God had translated him: for before his translation he had this testimony, that he pleased God.
HEB|11|6|But without faith it is impossible to please him: for he that cometh to God must believe that he is, and that he is a rewarder of them that diligently seek him.
HEB|11|7|By faith Noah, being warned of God of things not seen as yet, moved with fear, prepared an ark to the saving of his house; by the which he condemned the world, and became heir of the righteousness which is by faith.
HEB|11|8|By faith Abraham, when he was called to go out into a place which he should after receive for an inheritance, obeyed; and he went out, not knowing whither he went.
HEB|11|9|By faith he sojourned in the land of promise, as in a strange country, dwelling in tabernacles with Isaac and Jacob, the heirs with him of the same promise:
HEB|11|10|For he looked for a city which hath foundations, whose builder and maker is God.
HEB|11|11|Through faith also Sara herself received strength to conceive seed, and was delivered of a child when she was past age, because she judged him faithful who had promised.
HEB|11|12|Therefore sprang there even of one, and him as good as dead, so many as the stars of the sky in multitude, and as the sand which is by the sea shore innumerable.
HEB|11|13|These all died in faith, not having received the promises, but having seen them afar off, and were persuaded of them, and embraced them, and confessed that they were strangers and pilgrims on the earth.
HEB|11|14|For they that say such things declare plainly that they seek a country.
HEB|11|15|And truly, if they had been mindful of that country from whence they came out, they might have had opportunity to have returned.
HEB|11|16|But now they desire a better country, that is, an heavenly: wherefore God is not ashamed to be called their God: for he hath prepared for them a city.
HEB|11|17|By faith Abraham, when he was tried, offered up Isaac: and he that had received the promises offered up his only begotten son,
HEB|11|18|Of whom it was said, That in Isaac shall thy seed be called:
HEB|11|19|Accounting that God was able to raise him up, even from the dead; from whence also he received him in a figure.
HEB|11|20|By faith Isaac blessed Jacob and Esau concerning things to come.
HEB|11|21|By faith Jacob, when he was a dying, blessed both the sons of Joseph; and worshipped, leaning upon the top of his staff.
HEB|11|22|By faith Joseph, when he died, made mention of the departing of the children of Israel; and gave commandment concerning his bones.
HEB|11|23|By faith Moses, when he was born, was hid three months of his parents, because they saw he was a proper child; and they were not afraid of the king's commandment.
HEB|11|24|By faith Moses, when he was come to years, refused to be called the son of Pharaoh's daughter;
HEB|11|25|Choosing rather to suffer affliction with the people of God, than to enjoy the pleasures of sin for a season;
HEB|11|26|Esteeming the reproach of Christ greater riches than the treasures in Egypt: for he had respect unto the recompence of the reward.
HEB|11|27|By faith he forsook Egypt, not fearing the wrath of the king: for he endured, as seeing him who is invisible.
HEB|11|28|Through faith he kept the passover, and the sprinkling of blood, lest he that destroyed the firstborn should touch them.
HEB|11|29|By faith they passed through the Red sea as by dry land: which the Egyptians assaying to do were drowned.
HEB|11|30|By faith the walls of Jericho fell down, after they were compassed about seven days.
HEB|11|31|By faith the harlot Rahab perished not with them that believed not, when she had received the spies with peace.
HEB|11|32|And what shall I more say? for the time would fail me to tell of Gedeon, and of Barak, and of Samson, and of Jephthae; of David also, and Samuel, and of the prophets:
HEB|11|33|Who through faith subdued kingdoms, wrought righteousness, obtained promises, stopped the mouths of lions.
HEB|11|34|Quenched the violence of fire, escaped the edge of the sword, out of weakness were made strong, waxed valiant in fight, turned to flight the armies of the aliens.
HEB|11|35|Women received their dead raised to life again: and others were tortured, not accepting deliverance; that they might obtain a better resurrection:
HEB|11|36|And others had trial of cruel mockings and scourgings, yea, moreover of bonds and imprisonment:
HEB|11|37|They were stoned, they were sawn asunder, were tempted, were slain with the sword: they wandered about in sheepskins and goatskins; being destitute, afflicted, tormented;
HEB|11|38|(Of whom the world was not worthy:) they wandered in deserts, and in mountains, and in dens and caves of the earth.
HEB|11|39|And these all, having obtained a good report through faith, received not the promise:
HEB|11|40|God having provided some better thing for us, that they without us should not be made perfect.
HEB|12|1|Wherefore seeing we also are compassed about with so great a cloud of witnesses, let us lay aside every weight, and the sin which doth so easily beset us, and let us run with patience the race that is set before us,
HEB|12|2|Looking unto Jesus the author and finisher of our faith; who for the joy that was set before him endured the cross, despising the shame, and is set down at the right hand of the throne of God.
HEB|12|3|For consider him that endured such contradiction of sinners against himself, lest ye be wearied and faint in your minds.
HEB|12|4|Ye have not yet resisted unto blood, striving against sin.
HEB|12|5|And ye have forgotten the exhortation which speaketh unto you as unto children, My son, despise not thou the chastening of the Lord, nor faint when thou art rebuked of him:
HEB|12|6|For whom the Lord loveth he chasteneth, and scourgeth every son whom he receiveth.
HEB|12|7|If ye endure chastening, God dealeth with you as with sons; for what son is he whom the father chasteneth not?
HEB|12|8|But if ye be without chastisement, whereof all are partakers, then are ye bastards, and not sons.
HEB|12|9|Furthermore we have had fathers of our flesh which corrected us, and we gave them reverence: shall we not much rather be in subjection unto the Father of spirits, and live?
HEB|12|10|For they verily for a few days chastened us after their own pleasure; but he for our profit, that we might be partakers of his holiness.
HEB|12|11|Now no chastening for the present seemeth to be joyous, but grievous: nevertheless afterward it yieldeth the peaceable fruit of righteousness unto them which are exercised thereby.
HEB|12|12|Wherefore lift up the hands which hang down, and the feeble knees;
HEB|12|13|And make straight paths for your feet, lest that which is lame be turned out of the way; but let it rather be healed.
HEB|12|14|Follow peace with all men, and holiness, without which no man shall see the Lord:
HEB|12|15|Looking diligently lest any man fail of the grace of God; lest any root of bitterness springing up trouble you, and thereby many be defiled;
HEB|12|16|Lest there be any fornicator, or profane person, as Esau, who for one morsel of meat sold his birthright.
HEB|12|17|For ye know how that afterward, when he would have inherited the blessing, he was rejected: for he found no place of repentance, though he sought it carefully with tears.
HEB|12|18|For ye are not come unto the mount that might be touched, and that burned with fire, nor unto blackness, and darkness, and tempest,
HEB|12|19|And the sound of a trumpet, and the voice of words; which voice they that heard intreated that the word should not be spoken to them any more:
HEB|12|20|(For they could not endure that which was commanded, And if so much as a beast touch the mountain, it shall be stoned, or thrust through with a dart:
HEB|12|21|And so terrible was the sight, that Moses said, I exceedingly fear and quake:)
HEB|12|22|But ye are come unto mount Sion, and unto the city of the living God, the heavenly Jerusalem, and to an innumerable company of angels,
HEB|12|23|To the general assembly and church of the firstborn, which are written in heaven, and to God the Judge of all, and to the spirits of just men made perfect,
HEB|12|24|And to Jesus the mediator of the new covenant, and to the blood of sprinkling, that speaketh better things that that of Abel.
HEB|12|25|See that ye refuse not him that speaketh. For if they escaped not who refused him that spake on earth, much more shall not we escape, if we turn away from him that speaketh from heaven:
HEB|12|26|Whose voice then shook the earth: but now he hath promised, saying, Yet once more I shake not the earth only, but also heaven.
HEB|12|27|And this word, Yet once more, signifieth the removing of those things that are shaken, as of things that are made, that those things which cannot be shaken may remain.
HEB|12|28|Wherefore we receiving a kingdom which cannot be moved, let us have grace, whereby we may serve God acceptably with reverence and godly fear:
HEB|12|29|For our God is a consuming fire.
HEB|13|1|Let brotherly love continue.
HEB|13|2|Be not forgetful to entertain strangers: for thereby some have entertained angels unawares.
HEB|13|3|Remember them that are in bonds, as bound with them; and them which suffer adversity, as being yourselves also in the body.
HEB|13|4|Marriage is honourable in all, and the bed undefiled: but whoremongers and adulterers God will judge.
HEB|13|5|Let your conversation be without covetousness; and be content with such things as ye have: for he hath said, I will never leave thee, nor forsake thee.
HEB|13|6|So that we may boldly say, The Lord is my helper, and I will not fear what man shall do unto me.
HEB|13|7|Remember them which have the rule over you, who have spoken unto you the word of God: whose faith follow, considering the end of their conversation.
HEB|13|8|Jesus Christ the same yesterday, and to day, and for ever.
HEB|13|9|Be not carried about with divers and strange doctrines. For it is a good thing that the heart be established with grace; not with meats, which have not profited them that have been occupied therein.
HEB|13|10|We have an altar, whereof they have no right to eat which serve the tabernacle.
HEB|13|11|For the bodies of those beasts, whose blood is brought into the sanctuary by the high priest for sin, are burned without the camp.
HEB|13|12|Wherefore Jesus also, that he might sanctify the people with his own blood, suffered without the gate.
HEB|13|13|Let us go forth therefore unto him without the camp, bearing his reproach.
HEB|13|14|For here have we no continuing city, but we seek one to come.
HEB|13|15|By him therefore let us offer the sacrifice of praise to God continually, that is, the fruit of our lips giving thanks to his name.
HEB|13|16|But to do good and to communicate forget not: for with such sacrifices God is well pleased.
HEB|13|17|Obey them that have the rule over you, and submit yourselves: for they watch for your souls, as they that must give account, that they may do it with joy, and not with grief: for that is unprofitable for you.
HEB|13|18|Pray for us: for we trust we have a good conscience, in all things willing to live honestly.
HEB|13|19|But I beseech you the rather to do this, that I may be restored to you the sooner.
HEB|13|20|Now the God of peace, that brought again from the dead our Lord Jesus, that great shepherd of the sheep, through the blood of the everlasting covenant,
HEB|13|21|Make you perfect in every good work to do his will, working in you that which is wellpleasing in his sight, through Jesus Christ; to whom be glory for ever and ever. Amen.
HEB|13|22|And I beseech you, brethren, suffer the word of exhortation: for I have written a letter unto you in few words.
HEB|13|23|Know ye that our brother Timothy is set at liberty; with whom, if he come shortly, I will see you.
HEB|13|24|Salute all them that have the rule over you, and all the saints. They of Italy salute you.
HEB|13|25|Grace be with you all. Amen.
