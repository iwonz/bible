NAH|1|1|Oraculum Nineve. Liber visio nis Nahum Elcesaei.
NAH|1|2|Deus aemulator et ulciscens Dominus,ulciscens Dominus et habens furorem,ulciscens Dominus in hostes suoset servans iram inimicis suis.
NAH|1|3|Dominus patiens et magnus fortitudine,nullumque impunitum derelinquet Dominus.In tempestate et turbine via eius,et nubes pulvis pedum eius.
NAH|1|4|Increpans mare et exsiccans illudet omnia flumina ad desertum deducens.Elanguit Basan et Carmelus,et flos Libani elanguit.
NAH|1|5|Montes commoti sunt ab eo,et colles conturbati;et contremuit terra a facie eiuset orbis et omnes habitantes in eo.
NAH|1|6|Ante faciem indignationis eius quis stabit,et quis resistet in aestu furoris eius? Indignatio eius effusa est ut ignis,et petrae dissolutae sunt ab eo.
NAH|1|7|Bonus Dominus,refugium in die tribulationiset sciens sperantes in se
NAH|1|8|et in diluvio transeunte;consummationem faciet adversariorum suorum,et inimicos eius persequentur tenebrae.
NAH|1|9|Quid cogitatis contra Dominum?Consummationem ipse faciet;non consurget duplex tribulatio.
NAH|1|10|Sicut spinae condensae se invicem complectenteset sicut potatores inebriaticonsumentur quasi stipula omnino arida.
NAH|1|11|Ex te exivit cogitans contra Dominum malitiam,mente pertractans praevaricationem.
NAH|1|12|Haec dicit Dominus: Et si incolumes fuerint et numerosi,sic quoque attondentur et pertransibunt;afflixi te et non affligam te ultra.
NAH|1|13|Et nunc conteram virgam eius de dorso tuoet vincula tua disrumpam ".
NAH|1|14|Et praecipiet super te Dominus: Non seminabitur ex nomine tuo amplius.De domo dei tui disperdam sculptile et conflatile;ponam sepulcrum tuum,quia inhonoratus es ".
NAH|2|1|Ecce super montes pedes evan gelizantiset annuntiantis pacem.Celebra, Iuda, festivitates tuaset redde vota tua,quia non adiciet ultra ut pertranseat in te Belial:totus interiit.
NAH|2|2|Ascendit, qui dispergat, contra te. Custodi munitionem,contemplare viam, conforta lumbos, robora virtutem valde ".
NAH|2|3|Quia restituet Dominus magnificentiam Iacobsicut magnificentiam Israel,quia praedones praedati sunt eoset propagines eorum corruperunt.
NAH|2|4|Clipeus fortium eius ruber,viri exercitus in coccineis;ignitae laminae ferreae curruum,quando praeparat bellum,et equites agitantur.
NAH|2|5|In viis furibundae currunt quadrigae,invicem colliduntur in plateis;aspectus eorum quasi lampades,quasi fulgura discurrentia.
NAH|2|6|Recordatur fortium suorum,ruunt in itineribus suis;currunt ad murum,et praeparatur umbraculum.
NAH|2|7|Portae fluviorum apertae sunt,palatium tremit.
NAH|2|8|Et speciosa denudatur, tollitur,et ancillae eius gemunt ut columbae et percutiunt corda sua.
NAH|2|9|Et Nineve quasi piscina aquarum,cuius aquae fugiunt. State, state! ";sed non est qui revertatur.
NAH|2|10|" Diripite argentum, diripite aurum! ".Et non est finis divitiarum;thesaurus ex omnibus vasis desiderabilibus.
NAH|2|11|Dissipata et vastata et dilacerata,et cor tabescens,et dissolutio geniculorum;et tremor in cunctis renibus,et facies omnium eorum candentes.
NAH|2|12|Ubi est habitaculum leonum,et spelunca catulorum leonum,ad quam ivit leo, ut duceret illuc catulum leonis,et non erat qui exterreret?
NAH|2|13|Leo cepit sufficienter catulis suiset necavit leaenis suis;et implevit praeda speluncas suaset cubile suum rapina.
NAH|2|14|" Ecce ego ad te,dicit Dominus exercituum,et succendam usque ad fumum quadrigas tuas;et leunculos tuos comedet gladius,et exterminabo de terra praedam tuam,et non audietur ultra vox nuntiorum tuorum ".
NAH|3|1|Vae, civitas sanguinum,universa mendaciipraeda plena!Non recedet a te rapina.
NAH|3|2|Vox flagellorum et vox strepitus rotarum,equi frementes et quadrigae ferventes,equites irruentes
NAH|3|3|et gladii micantes et hastae fulguranteset multitudo interfectorum et acervi mortuorum;nec est finis cadaverum,et corruunt super corpora.
NAH|3|4|Hoc propter multitudinem fornicationum meretricisspeciosae et gratae et habentis maleficia,quae vendidit gentes fornicationibus suiset nationes maleficiis suis.
NAH|3|5|" Ecce ego ad te,dicit Dominus exercituum;et levabo vestimentum tuum in faciem tuamet ostendam gentibus nuditatem tuamet regnis ignominiam tuam.
NAH|3|6|Et proiciam super te abominationeset contumeliis te afficiam;et ponam te in exemplum.
NAH|3|7|Et erit: omnis, qui viderit te,resiliet a te et dicet:Vastata est Nineve!Quis dolebit super eam?Unde quaeram consolatorem tibi?".
NAH|3|8|Numquid melior es quam Noamon,quae habitabat in fluminibus?Aquae in circuitu eius:cuius vallum mare,aquae muri eius.
NAH|3|9|Chus fuit fortitudo eiuset Aegyptus, cuius non est finis;Phut et Libyes fuerunt in auxilio eius.
NAH|3|10|Sed et ipsa in transmigrationem ducta est,ivit in captivitatem.Parvuli eius elisi suntin capite omnium viarum;et super inclitos eius miserunt sortem,et omnes optimates eius constricti sunt in compedibus.
NAH|3|11|Et tu ergo inebriaberis,eris despecta;et tu quaeresrefugium ab inimico.
NAH|3|12|Omnes munitiones tuae sicut ficuscum ficis praecocibus:si concussae fuerint,cadent in os comedentis.
NAH|3|13|Ecce populus tuus,mulieres in medio tui;inimicis tuis late patebuntportae terrae tuae;devorabit ignis vectes tuos.
NAH|3|14|Aquam propter obsidionem hauri tibi,firma munitiones tuas;intra in lutum et calca argillam,tene typum laterum.
NAH|3|15|Ibi comedet te ignis,peribis gladio,devorabit te ut bruchus.Augere ut bruchus,multiplicare ut locusta.
NAH|3|16|Plures fecisti negotiatores tuosquam stellae sint caeli;bruchus exuit pellemet avolavit.
NAH|3|17|Custodes tui quasi locustae,et scribae tui quasi agmen locustarum,quae considunt in saepibusin die frigoris;sol ortus est,et avolaverunt,non est cognitus locus earum,ubi fuerint.
NAH|3|18|Dormiunt pastores tui, rex Assyriae,requiescunt principes tui;dispersus est populus tuus in montibus,et non est qui congreget.
NAH|3|19|Non est remedium fracturae tuae,insanabilis est plaga tua;omnes, qui audierint auditionem tuam,plaudent manibus super te,quia super quem non transiitmalitia tua semper? ".
