2JOHN|1|1|The elder,
2JOHN|1|2|To the chosen lady and her children, whom I love in the truth--and not I only, but also all who know the truth--because of the truth, which lives in us and will be with us forever:
2JOHN|1|3|Grace, mercy and peace from God the Father and from Jesus Christ, the Father's Son, will be with us in truth and love.
2JOHN|1|4|It has given me great joy to find some of your children walking in the truth, just as the Father commanded us.
2JOHN|1|5|And now, dear lady, I am not writing you a new command but one we have had from the beginning. I ask that we love one another.
2JOHN|1|6|And this is love: that we walk in obedience to his commands. As you have heard from the beginning, his command is that you walk in love.
2JOHN|1|7|Many deceivers, who do not acknowledge Jesus Christ as coming in the flesh, have gone out into the world. Any such person is the deceiver and the antichrist.
2JOHN|1|8|Watch out that you do not lose what you have worked for, but that you may be rewarded fully.
2JOHN|1|9|Anyone who runs ahead and does not continue in the teaching of Christ does not have God; whoever continues in the teaching has both the Father and the Son.
2JOHN|1|10|If anyone comes to you and does not bring this teaching, do not take him into your house or welcome him.
2JOHN|1|11|Anyone who welcomes him shares in his wicked work.
2JOHN|1|12|I have much to write to you, but I do not want to use paper and ink. Instead, I hope to visit you and talk with you face to face, so that our joy may be complete.
2JOHN|1|13|The children of your chosen sister send their greetings.
