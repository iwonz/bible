MATT|1|1|Книга родоводу Ісуса Христа, Сина Давидового, Сина Авраамового:
MATT|1|2|Авраам породив Ісака, а Ісак породив Якова, а Яків породив Юду й братів його.
MATT|1|3|Юда ж породив Фареса та Зару від Тамари. Фарес же породив Есрома, а Есром породив Арама.
MATT|1|4|А Арам породив Амінадава, Амінадав же породив Наассона, а Наассон породив Салмона.
MATT|1|5|Салмон же породив Вооза від Рахави, а Вооз породив Йовіда від Рути, Йовід же породив Єссея.
MATT|1|6|А Єссей породив царя Давида, Давид же породив Соломона від Урієвої.
MATT|1|7|Соломон же породив Ровоама, а Ровоам породив Авію, а Авія породив Асафа.
MATT|1|8|Асаф же породив Йосафата, а Йосафат породив Йорама, Йорам же породив Озію.
MATT|1|9|Озія ж породив Йоатама, а Йоатам породив Ахаза, Ахаз же породив Єзекію.
MATT|1|10|А Єзекія породив Манасію, Манасія ж породив Амоса, а Амос породив Йосію.
MATT|1|11|Йосія ж породив Йоякима, Йояким породив Єхонію й братів його за вавилонського переселення.
MATT|1|12|А по вавилонськім переселенні Єхонія породив Салатіїля, а Салатіїль породив Зоровавеля.
MATT|1|13|Зоровавель же породив Авіюда, а Авіюд породив Еліякима, а Еліяким породив Азора.
MATT|1|14|Азор же породив Садока, а Садок породив Ахіма, а Ахім породив Еліюда.
MATT|1|15|Еліюд же породив Елеазара, а Елеазар породив Маттана, а Маттан породив Якова.
MATT|1|16|А Яків породив Йосипа, мужа Марії, що з неї родився Ісус, званий Христос.
MATT|1|17|А всіх поколінь від Авраама аж до Давида чотирнадцять поколінь, і від Давида аж до вавилонського переселення чотирнадцять поколінь, і від вавилонського переселення до Христа поколінь чотирнадцять.
MATT|1|18|Народження ж Ісуса Христа сталося так. Коли Його матір Марію заручено з Йосипом, то перш, ніж зійшлися вони, виявилося, що вона має в утробі від Духа Святого.
MATT|1|19|А Йосип, муж її, бувши праведний, і не бажавши ославити її, хотів тайкома відпустити її.
MATT|1|20|Коли ж він те подумав, ось з'явивсь йому Ангол Господній у сні, промовляючи: Йосипе, сину Давидів, не бійся прийняти Марію, дружину свою, бо зачате в ній то від Духа Святого.
MATT|1|21|І вона вродить Сина, ти ж даси Йому йменна Ісус, бо спасе Він людей Своїх від їхніх гріхів.
MATT|1|22|А все оце сталось, щоб збулося сказане пророком від Господа, який провіщає:
MATT|1|23|Ось діва в утробі зачне, і Сина породить, і назвуть Йому Ймення Еммануїл, що в перекладі є: З нами Бог.
MATT|1|24|Як прокинувся ж Йосип зо сну, то зробив, як звелів йому Ангол Господній, і прийняв він дружину свою.
MATT|1|25|І не знав він її, аж Сина свого первородженого вона породила, а він дав Йому ймення Ісус.
MATT|2|1|Коли ж народився Ісус у Віфлеємі Юдейськім, за днів царя Ірода, то ось мудреці прибули до Єрусалиму зо сходу,
MATT|2|2|і питали: Де народжений Цар Юдейський? Бо на сході ми бачили зорю Його, і прибули поклонитись Йому.
MATT|2|3|І, як зачув це цар Ірод, занепокоївся, і з ним увесь Єрусалим.
MATT|2|4|І, зібравши всіх первосвящеників і книжників людських, він випитував у них, де має Христос народитись?
MATT|2|5|Вони ж відказали йому: У Віфлеємі Юдейськім, бо в пророка написано так:
MATT|2|6|І ти, Віфлеєме, земле Юдина, не менший нічим між осадами Юдиними, бо з тебе з'явиться Вождь, що буде Він пасти народ Мій ізраїльський.
MATT|2|7|Тоді Ірод покликав таємно отих мудреців, і докладно випитував їх про час, коли з'явилась зоря.
MATT|2|8|І він відіслав їх до Віфлеєму, говорячи: Ідіть, і пильно розвідайтеся про Дитятко; а як знайдете, сповістіть мене, щоб і я міг піти й поклонитись Йому.
MATT|2|9|Вони ж царя вислухали й відійшли. І ось зоря, що на сході вони її бачили, ішла перед ними, аж прийшла й стала зверху, де Дитятко було.
MATT|2|10|А бачивши зорю, вони надзвичайно зраділи.
MATT|2|11|І, ввійшовши до дому, знайшли там Дитятко з Марією, Його матір'ю. І вони впали ницьма, і вклонились Йому. І, відчинивши скарбниці свої, піднесли Йому свої дари: золото, ладан та смирну.
MATT|2|12|А вві сні остережені, щоб не вертатись до Ірода, відійшли вони іншим шляхом до своєї землі.
MATT|2|13|Як вони ж відійшли, ось Ангол Господній з'явивсь у сні Йосипові та й сказав: Уставай, візьми Дитятко та матір Його, і втікай до Єгипту, і там зоставайся, аж поки скажу тобі, бо Дитятка шукатиме Ірод, щоб Його погубити.
MATT|2|14|І він устав, узяв Дитятко та матір Його вночі, та й пішов до Єгипту.
MATT|2|15|І він там зоставався аж до смерти Іродової, щоб збулося сказане від Господа пророком, який провіщає: Із Єгипту покликав Я Сина Свого.
MATT|2|16|Спостеріг тоді Ірод, що ті мудреці насміялися з нього, та й розгнівався дуже, і послав повбивати в Віфлеємі й по всій тій околиці всіх дітей від двох років і менше, за часом, що його в мудреців він був випитав.
MATT|2|17|Тоді справдилось те, що сказав Єремія пророк, промовляючи:
MATT|2|18|Чути голос у Рамі, плач і ридання та голосіння велике: Рахиль плаче за дітьми своїми, і не дається розважити себе, бо нема їх...
MATT|2|19|Коли ж Ірод умер, ось Ангол Господній з'явився в Єгипті вві сні Йосипові, та й промовив:
MATT|2|20|Уставай, візьми Дитятко та матір Його, та йди в землю Ізраїлеву, бо вимерли ті, хто шукав був душу Дитини.
MATT|2|21|І він устав, узяв Дитятко та матір Його, і прийшов у землю Ізраїлеву.
MATT|2|22|Та прочувши, що царює в Юдеї Архелай, замість Ірода, батька свого, побоявся піти туди він. А вві сні остережений, відійшов до країв галілейських.
MATT|2|23|А прибувши, оселився у місті, на ім'я Назарет, щоб збулося пророками сказане, що Він Назарянин буде званий.
MATT|3|1|Тими ж днями приходить Іван Христитель, і проповідує в пустині юдейській,
MATT|3|2|та й каже: Покайтесь, бо наблизилось Царство Небесне!
MATT|3|3|Бо він той, що про нього сказав був Ісая пророк, промовляючи: Голос того, хто кличе: В пустині готуйте дорогу для Господа, рівняйте стежки Йому!
MATT|3|4|Сам же Іван мав одежу собі з верблюжого волосу, і пояс ремінний на стегнах своїх; а пожива для нього була сарана та мед польовий.
MATT|3|5|Тоді до нього виходив Єрусалим, і вся Юдея, і вся йорданська околиця,
MATT|3|6|і в річці Йордані христились від нього, і визнавали гріхи свої.
MATT|3|7|Як побачив же він багатьох фарисеїв та саддукеїв, що приходять на хрищення, то промовив до них: Роде зміїний, хто вас надоумив утікати від гніву майбутнього?
MATT|3|8|Отож, учиніть гідний плід покаяння!
MATT|3|9|І не думайте говорити в собі: Ми маємо отця Авраама. Кажу бо я вам, що Бог може піднести дітей Авраамові з цього каміння!
MATT|3|10|Бо вже до коріння дерев і сокира прикладена: кожне ж дерево, що доброго плоду не родить, буде зрубане та й в огонь буде вкинене.
MATT|3|11|Я хрищу вас водою на покаяння, але Той, Хто йде по мені, потужніший від мене: я недостойний понести взуття Йому! Він христитиме вас Святим Духом й огнем.
MATT|3|12|У руці Своїй має Він віячку, і перечистить Свій тік: пшеницю Свою Він збере до засіків, а полову попалить ув огні невгасимім.
MATT|3|13|Тоді прибуває Ісус із Галілеї понад Йордан до Івана, щоб христитись від нього.
MATT|3|14|Але перешкоджав він Йому й говорив: Я повинен христитись від Тебе, і чи Тобі йти до мене?
MATT|3|15|А Ісус відповів і сказав йому: Допусти це тепер, бо так годиться нам виповнити усю правду. Тоді допустив він Його.
MATT|3|16|І охристившись Ісус, зараз вийшов із води. І ось небо розкрилось, і побачив Іван Духа Божого, що спускався, як голуб, і сходив на Нього.
MATT|3|17|І ось голос почувся із неба: Це Син Мій Улюблений, що Його Я вподобав!
MATT|4|1|Потому Ісус був поведений Духом у пустиню, щоб диявол Його спокушав.
MATT|4|2|І постив Він сорок день і сорок ночей, а вкінці зголоднів.
MATT|4|3|І ось приступив до Нього спокусник, і сказав: Коли Ти Син Божий, скажи, щоб каміння це стало хлібами!
MATT|4|4|А Він відповів і промовив: Написано: Не хлібом самим буде жити людина, але кожним словом, що походить із уст Божих.
MATT|4|5|Тоді забирає диявол Його в святе місто, і ставить Його на наріжника храму,
MATT|4|6|та й каже Йому: Коли Ти Син Божий, то кинься додолу, бож написано: Він накаже про Тебе Своїм Анголам, і вони на руках понесуть Тебе, щоб об камінь коли не спіткнув Ти Своєї ноги.
MATT|4|7|Ісус відказав йому: Ще написано: Не спокушуй Господа Бога свого!
MATT|4|8|Знов диявол бере Його на височезную гору, і показує Йому всі царства на світі та їхнюю славу,
MATT|4|9|та й каже до Нього: Це все Тобі дам, якщо впадеш і мені Ти поклонишся!
MATT|4|10|Тоді каже до нього Ісус: Відійди, сатано! Бож написано: Господеві Богові своєму вклоняйся, і служи Одному Йому!
MATT|4|11|Тоді позоставив диявол Його. І ось Анголи приступили, і служили Йому.
MATT|4|12|Як довідавсь Ісус, що Івана ув'язнено, перейшов у Галілею.
MATT|4|13|І, покинувши Він Назарета, прийшов й оселився в Капернаумі приморськім, на границі країн Завулонової й Нефталимової,
MATT|4|14|щоб справдилось те, що сказав був Ісая пророк, промовляючи:
MATT|4|15|Завулонова земле, і Нефталимова земле, за Йорданом при морській дорозі, Галілеє поганська!
MATT|4|16|Народ, що в темноті сидів, світло велике побачив, а тим, хто сидів у країні смертельної тіні, засяяло світло.
MATT|4|17|Із того часу Ісус розпочав проповідувати й промовляти: Покайтеся, бо наблизилось Царство Небесне!
MATT|4|18|Як проходив же Він поблизу Галілейського моря, то побачив двох братів: Симона, що зветься Петром, та Андрія, його брата, що невода в море закидали, бо рибалки були.
MATT|4|19|І Він каже до них: Ідіть за Мною, Я зроблю вас ловцями людей!
MATT|4|20|І вони зараз покинули сіті, та й пішли вслід за Ним.
MATT|4|21|І, далі пішовши звідти, Він побачив двох інших братів, Зеведеєвого сина Якова та Івана, його брата, із Зеведеєм, їхнім батьком, що лагодили свого невода в човні, і покликав Він їх.
MATT|4|22|Вони зараз залишили човна та батька свого, та й пішли вслід за Ним.
MATT|4|23|І ходив Він по всій Галілеї, по їхніх синагогах навчаючи, та Євангелію Царства проповідуючи, і вздоровлюючи всяку недугу, і всяку неміч між людьми.
MATT|4|24|А чутка про Нього пішла по всій Сирії. І водили до Нього недужих усіх, хто терпів на різні хвороби та муки, і біснуватих, і сновид, і розслаблених, і Він їх уздоровляв.
MATT|4|25|І багато людей ішло за Ним і з Галілеї, і з Десятимістя, і з Єрусалиму, і з Юдеї, і з Зайордання.
MATT|5|1|І, побачивши натовп, Він вийшов на гору. А як сів, підійшли Його учні до Нього.
MATT|5|2|І, відкривши уста Свої, Він навчати їх став, промовляючи:
MATT|5|3|Блаженні вбогі духом, бо їхнєє Царство Небесне.
MATT|5|4|Блаженні засмучені, бо вони будуть утішені.
MATT|5|5|Блаженні лагідні, бо землю вспадкують вони.
MATT|5|6|Блаженні голодні та спрагнені правди, бо вони нагодовані будуть.
MATT|5|7|Блаженні милостиві, бо помилувані вони будуть.
MATT|5|8|Блаженні чисті серцем, бо вони будуть бачити Бога.
MATT|5|9|Блаженні миротворці, бо вони синами Божими стануть.
MATT|5|10|Блаженні вигнані за правду, бо їхнє Царство Небесне.
MATT|5|11|Блаженні ви, як ганьбити та гнати вас будуть, і будуть облудно на вас наговорювати всяке слово лихе ради Мене.
MATT|5|12|Радійте та веселіться, нагорода бо ваша велика на небесах! Бо так гнали й пророків, що були перед вами.
MATT|5|13|Ви сіль землі. Коли сіль ізвітріє, то чим насолити її? Не придасться вона вже нінащо, хіба щоб надвір була висипана та потоптана людьми.
MATT|5|14|Ви світло для світу. Не може сховатися місто, що стоїть на верховині гори.
MATT|5|15|І не запалюють світильника, щоб поставити його під посудину, але на свічник, і світить воно всім у домі.
MATT|5|16|Отак ваше світло нехай світить перед людьми, щоб вони бачили ваші добрі діла, та прославляли Отця вашого, що на небі.
MATT|5|17|Не подумайте, ніби Я руйнувати Закон чи Пророків прийшов, Я не руйнувати прийшов, але виконати.
MATT|5|18|Поправді ж кажу вам: доки небо й земля не минеться, ані йота єдина, ані жаден значок із Закону не минеться, аж поки не збудеться все.
MATT|5|19|Хто ж порушить одну з найменших цих заповідей, та й людей так навчить, той буде найменшим у Царстві Небеснім; а хто виконає та й навчить, той стане великим у Царстві Небеснім.
MATT|5|20|Кажу бо Я вам: коли праведність ваша не буде рясніша, як книжників та фарисеїв, то не ввійдете в Царство Небесне!
MATT|5|21|Ви чули, що було стародавнім наказане: Не вбивай, а хто вб'є, підпадає він судові.
MATT|5|22|А Я вам кажу, що кожен, хто гнівається на брата свого, підпадає вже судові. А хто скаже на брата свого: рака, підпадає верховному судові, а хто скаже дурний, підпадає геєнні огненній.
MATT|5|23|Тому, коли принесеш ти до жертівника свого дара, та тут ізгадаєш, що брат твій щось має на тебе,
MATT|5|24|залиши отут дара свого перед жертівником, і піди, примирись перше з братом своїм, і тоді повертайся, і принось свого дара.
MATT|5|25|Зо своїм супротивником швидко мирися, доки з ним на дорозі ще ти, щоб тебе супротивник судді не віддав, а суддя щоб прислужникові тебе не передав, і щоб тебе до в'язниці не вкинули.
MATT|5|26|Поправді кажу тобі: Не вийдеш ізвідти, поки не віддаси ти й останнього шеляга!
MATT|5|27|Ви чули, що сказано: Не чини перелюбу.
MATT|5|28|А Я вам кажу, що кожен, хто на жінку подивиться із пожадливістю, той уже вчинив із нею перелюб у серці своїм.
MATT|5|29|Коли праве око твоє спокушає тебе, його вибери, і кинь від себе: бо краще тобі, щоб загинув один із твоїх членів, аніж до геєнни все тіло твоє було вкинене.
MATT|5|30|І як правиця твоя спокушає тебе, відітни її й кинь від себе: бо краще тобі, щоб загинув один із твоїх членів, аніж до геєнни все тіло твоє було вкинене.
MATT|5|31|Також сказано: Хто дружину свою відпускає, нехай дасть їй листа розводового.
MATT|5|32|А Я вам кажу, що кожен, хто пускає дружину свою, крім провини розпусти, той доводить її до перелюбу. І хто з відпущеною побереться, той чинить перелюб.
MATT|5|33|Ще ви чули, що було стародавнім наказане: Не клянись неправдиво, але виконуй клятви свої перед Господом.
MATT|5|34|А Я вам кажу не клястися зовсім: ані небом, бо воно престол Божий;
MATT|5|35|ні землею, бо підніжок для ніг Його це; ані Єрусалимом, бо він місто Царя Великого;
MATT|5|36|не клянись головою своєю, бо навіть однієї волосинки ти не можеш учинити білою чи чорною.
MATT|5|37|Ваше ж слово хай буде: так-так, ні-ні. А що більше над це, то те від лукавого.
MATT|5|38|Ви чули, що сказано: Око за око, і зуб за зуба.
MATT|5|39|А Я вам кажу не противитись злому. І коли вдарить тебе хто у праву щоку твою, підстав йому й другу.
MATT|5|40|А хто хоче тебе позивати й забрати сорочку твою, віддай і плаща йому.
MATT|5|41|А хто силувати тебе буде відбути подорожнє на милю одну, іди з ним навіть дві.
MATT|5|42|Хто просить у тебе то дай, а хто хоче позичити в тебе не відвертайсь від нього.
MATT|5|43|Ви чули, що сказано: Люби свого ближнього, і ненавидь свого ворога.
MATT|5|44|А Я вам кажу: Любіть ворогів своїх, благословляйте тих, хто вас проклинає, творіть добро тим, хто ненавидить вас, і моліться за тих, хто вас переслідує,
MATT|5|45|щоб вам бути синами Отця вашого, що на небі, що наказує сходити сонцю Своєму над злими й над добрими, і дощ посилає на праведних і на неправедних.
MATT|5|46|Коли бо ви любите тих, хто вас любить, то яку нагороду ви маєте? Хіба не те саме й митники роблять?
MATT|5|47|І коли ви вітаєте тільки братів своїх, то що ж особливого робите? Чи й погани не чинять отак?
MATT|5|48|Отож, будьте досконалі, як досконалий Отець ваш Небесний!
MATT|6|1|Стережіться виставляти свою милостиню перед людьми, щоб бачили вас; а як ні, то не матимете нагороди від Отця вашого, що на небі.
MATT|6|2|Отож, коли чиниш ти милостиню, не сурми перед себе, як то роблять оті лицеміри по синагогах та вулицях, щоб хвалили їх люди. Поправді кажу вам: вони мають уже нагороду свою!
MATT|6|3|А як ти чиниш милостиню, хай не знатиме ліва рука твоя, що робить правиця твоя,
MATT|6|4|щоб таємна була твоя милостиня, а Отець твій, що бачить таємне, віддасть тобі явно.
MATT|6|5|А як молитеся, то не будьте, як ті лицеміри, що люблять ставати й молитися по синагогах та на перехрестях, щоб їх бачили люди. Поправді кажу вам: вони мають уже нагороду свою!
MATT|6|6|А ти, коли молишся, увійди до своєї комірчини, зачини свої двері, і помолися Отцеві своєму, що в таїні; а Отець твій, що бачить таємне, віддасть тобі явно.
MATT|6|7|А як молитеся, не проказуйте зайвого, як ті погани, бо думають, ніби вони будуть вислухані за своє велемовство.
MATT|6|8|Отож, не вподобляйтеся їм, бо знає Отець ваш, чого потребуєте, ще раніше за ваше прохання!
MATT|6|9|Ви ж моліться отак: Отче наш, що єси на небесах! Нехай святиться Ім'я Твоє,
MATT|6|10|нехай прийде Царство Твоє, нехай буде воля Твоя, як на небі, так і на землі.
MATT|6|11|Хліба нашого насущного дай нам сьогодні.
MATT|6|12|І прости нам довги наші, як і ми прощаємо винуватцям нашим.
MATT|6|13|І не введи нас у випробовування, але визволи нас від лукавого. Бо Твоє є царство, і сила, і слава навіки. Амінь.
MATT|6|14|Бо як людям ви простите прогріхи їхні, то простить і вам ваш Небесний Отець.
MATT|6|15|А коли ви не будете людям прощати, то й Отець ваш не простить вам прогріхів ваших.
MATT|6|16|А як постите, то не будьте сумні, як оті лицеміри: вони бо зміняють обличчя свої, щоб бачили люди, що постять вони. Поправді кажу вам: вони мають уже нагороду свою!
MATT|6|17|А ти, коли постиш, намасти свою голову, і лице своє вмий,
MATT|6|18|щоб ти посту свого не виявив людям, а Отцеві своєму, що в таїні; і Отець твій, що бачить таємне, віддасть тобі явно.
MATT|6|19|Не складайте скарбів собі на землі, де нищить їх міль та іржа, і де злодії підкопуються й викрадають.
MATT|6|20|Складайте ж собі скарби на небі, де ні міль, ні іржа їх не нищить, і де злодії до них не підкопуються та не крадуть.
MATT|6|21|Бо де скарб твій, там буде й серце твоє!
MATT|6|22|Око то світильник для тіла. Тож як око твоє буде здорове, то й усе тіло твоє буде світле.
MATT|6|23|А коли б твоє око лихе було, то й усе тіло твоє буде темне. Отож, коли світло, що в тобі, є темрява, то яка ж то велика та темрява!
MATT|6|24|Ніхто двом панам служити не може, бо або одного зненавидить, а другого буде любити, або буде триматись одного, а другого знехтує. Не можете Богові служити й мамоні.
MATT|6|25|Через те вам кажу: Не журіться про життя своє що будете їсти та що будете пити, ні про тіло своє, у що зодягнетеся. Чи ж не більше від їжі життя, а від одягу тіло?
MATT|6|26|Погляньте на птахів небесних, що не сіють, не жнуть, не збирають у клуні, та проте ваш Небесний Отець їх годує. Чи ж ви не багато вартніші за них?
MATT|6|27|Хто ж із вас, коли журиться, зможе додати до зросту свого бодай ліктя одного?
MATT|6|28|І про одяг чого ви клопочетесь? Погляньте на польові лілеї, як зростають вони, не працюють, ані не прядуть.
MATT|6|29|А Я вам кажу, що й сам Соломон у всій славі своїй не вдягався отак, як одна з них.
MATT|6|30|І коли польову ту траву, що сьогодні ось є, а взавтра до печі вкидається, Бог отак зодягає, скільки ж краще зодягне Він вас, маловірні!
MATT|6|31|Отож, не журіться, кажучи: Що ми будемо їсти, чи: Що будемо пити, або: У що ми зодягнемось?
MATT|6|32|Бож усього того погани шукають; але знає Отець ваш Небесний, що всього того вам потрібно.
MATT|6|33|Шукайте ж найперш Царства Божого й правди Його, а все це вам додасться.
MATT|6|34|Отож, не журіться про завтрашній день, бо завтра за себе само поклопочеться. Кожний день має досить своєї турботи!
MATT|7|1|Не судіть, щоб і вас не судили;
MATT|7|2|бо яким судом судити будете, таким же осудять і вас, і якою мірою будете міряти, такою відміряють вам.
MATT|7|3|І чого в оці брата свого ти заскалку бачиш, колоди ж у власному оці не чуєш?
MATT|7|4|Або як ти скажеш до брата свого: Давай вийму я заскалку з ока твого, коли он колода у власному оці?
MATT|7|5|Лицеміре, вийми перше колоду із власного ока, а потім побачиш, як вийняти заскалку з ока брата твого.
MATT|7|6|Не давайте святого псам, і не розсипайте перел своїх перед свиньми, щоб вони не потоптали їх ногами своїми, і, обернувшись, щоб не розшматували й вас...
MATT|7|7|Просіть і буде вам дано, шукайте і знайдете, стукайте і відчинять вам;
MATT|7|8|бо кожен, хто просить одержує, хто шукає знаходить, а хто стукає відчинять йому.
MATT|7|9|Чи ж то серед вас є людина, що подасть своєму синові каменя, коли хліба проситиме він?
MATT|7|10|Або коли риби проситиме, то подасть йому гадину?
MATT|7|11|Тож як ви, бувши злі, потрапите добрі дари своїм дітям давати, скільки ж більше Отець ваш Небесний подасть добра тим, хто проситиме в Нього!
MATT|7|12|Тож усе, чого тільки бажаєте, щоб чинили вам люди, те саме чиніть їм і ви. Бо в цьому Закон і Пророки.
MATT|7|13|Увіходьте тісними ворітьми, бо просторі ворота й широка дорога, що веде до погибелі, і нею багато-хто ходять.
MATT|7|14|Бо тісні ті ворота, і вузька та дорога, що веде до життя, і мало таких, що знаходять її!
MATT|7|15|Стережіться фальшивих пророків, що приходять до вас ув одежі овечій, а всередині хижі вовки.
MATT|7|16|По їхніх плодах ви пізнаєте їх. Бо хіба ж виноград на тернині збирають, або фіґи із будяків?
MATT|7|17|Так ото родить добрі плоди кожне дерево добре, а дерево зле плоди родить лихі.
MATT|7|18|Не може родить добре дерево плоду лихого, ані дерево зле плодів добрих родити.
MATT|7|19|Усяке ж дерево, що доброго плоду не родить, зрубується та в огонь укидається.
MATT|7|20|Ото ж бо, по їхніх плодах ви пізнаєте їх!
MATT|7|21|Не кожен, хто каже до Мене: Господи, Господи! увійде в Царство Небесне, але той, хто виконує волю Мого Отця, що на небі.
MATT|7|22|Багато-хто скажуть Мені того дня: Господи, Господи, хіба ми не Ім'ям Твоїм пророкували, хіба не Ім'ям Твоїм демонів ми виганяли, або не Ім'ям Твоїм чуда великі творили?
MATT|7|23|І їм оголошу Я тоді: Я ніколи не знав вас... Відійдіть від Мене, хто чинить беззаконня!
MATT|7|24|Отож, кожен, хто слухає цих Моїх слів і виконує їх, подібний до чоловіка розумного, що свій дім збудував на камені.
MATT|7|25|І линула злива, і розлилися річки, і буря знялася, і на дім отой кинулась, та не впав, бо на камені був він заснований.
MATT|7|26|А кожен, хто слухає цих Моїх слів, та їх не виконує, подібний до чоловіка того необачного, що свій дім збудував на піску.
MATT|7|27|І линула злива, і розлилися річки, і буря знялася й на дім отой кинулась, і він упав. І велика була та руїна його!
MATT|7|28|І ото, як Ісус закінчив ці слова, то народ дивувався з науки Його.
MATT|7|29|Бо навчав Він їх, як можновладний, а не як ті книжники їхні.
MATT|8|1|А коли Він зійшов із гори, услід за Ним ішов натовп великий.
MATT|8|2|І ось підійшов прокажений, уклонився Йому та й сказав: Коли, Господи, хочеш, Ти можеш очистити мене!
MATT|8|3|А Ісус простяг руку, і доторкнувся до нього, говорячи: Хочу, будь чистий! І тієї хвилини очистився той від своєї прокази.
MATT|8|4|І говорить до нього Ісус: Гляди, не розповідай нікому. Але йди, покажися священикові, та дар принеси, якого Мойсей заповів, їм на свідоцтво.
MATT|8|5|А коли Він до Капернауму ввійшов, то до Нього наблизився сотник, та й благати зачав Його,
MATT|8|6|кажучи: Господи, мій слуга лежить удома розслаблений, і тяжко страждає.
MATT|8|7|Він говорить йому: Я прийду й уздоровлю його.
MATT|8|8|А сотник Йому відповів: Недостойний я, Господи, щоб зайшов Ти під стріху мою... Та промов тільки слово, і видужає мій слуга!
MATT|8|9|Бо й я людина підвладна, і вояків під собою я маю; і одному кажу: піди то йде він, а тому: прийди і приходить, або рабові своєму: зроби те і він зробить.
MATT|8|10|Почувши таке, Ісус здивувався, і промовив до тих, хто йшов услід за Ним: Поправді кажу вам: навіть серед Ізраїля Я не знайшов був такої великої віри!
MATT|8|11|Кажу ж вам, що багато-хто прийдуть від сходу та заходу, і засядуть у Царстві Небеснім із Авраамом, Ісаком та Яковом.
MATT|8|12|Сини ж Царства повкидані будуть до темряви зовнішньої буде там плач і скрегіт зубів!...
MATT|8|13|І сказав Ісус сотникові: Іди, і як повірив ти, нехай так тобі й станеться! І тієї ж години одужав слуга його.
MATT|8|14|Як прийшов же Ісус до Петрового дому, то побачив тещу його, що лежала в гарячці.
MATT|8|15|І Він доторкнувся руки її, і гарячка покинула ту... І встала вона, та й Йому прислуговувала!
MATT|8|16|А коли настав вечір, привели багатьох біснуватих до Нього, і Він словом Своїм вигнав духів, а недужих усіх уздоровив,
MATT|8|17|щоб справдилося, що сказав був Ісая пророк, промовляючи: Він узяв наші немочі, і недуги поніс.
MATT|8|18|А як угледів Ісус навколо Себе багато народу, наказав переплинути на той бік.
MATT|8|19|І приступив один книжник та й до Нього сказав: Учителю, я піду за Тобою, хоч би куди ти пішов!
MATT|8|20|Промовляє до нього Ісус: Мають нори лисиці, а гнізда небесні пташки, Син же Людський не має де й голови прихилити...
MATT|8|21|А інший із учнів промовив до Нього: Дозволь мені, Господи, перше піти та батька свого поховати.
MATT|8|22|А Ісус йому каже: Іди за Мною, і зостав мертвим ховати мерців своїх!
MATT|8|23|І коли Він до човна вступив, за Ним увійшли Його учні.
MATT|8|24|І ось буря велика зірвалась на морі, аж човен зачав заливатися хвилями. А Він спав...
MATT|8|25|І кинулись учні, і збудили Його та й благали: Рятуй, Господи, гинемо!
MATT|8|26|А Він відповів їм: Чого полохливі ви, маловірні? Тоді встав, заказав бурі й морю, і тиша велика настала...
MATT|8|27|А народ дивувався й казав: Хто ж це такий, що вітри та море слухняні Йому?
MATT|8|28|І, як прибув Він на той бік, до землі Гадаринської, перестріли Його два біснуваті, що вийшли з могильних печер, дуже люті, так що ніхто не міг переходити тією дорогою.
MATT|8|29|І ось, вони стали кричати, говорячи: Що Тобі, Сину Божий, до нас? Прийшов Ти сюди передчасно нас мучити?
MATT|8|30|А оподаль від них пасся гурт великий свиней.
MATT|8|31|І просилися демони, кажучи: Коли виженеш нас, то пошли нас у той гурт свиней.
MATT|8|32|А Він відповів їм: Ідіть. І вийшли вони, і пішли в гурт свиней. І ось кинувся з кручі до моря ввесь гурт, і потопився в воді.
MATT|8|33|Пастухи ж повтікали; а коли прибули вони в місто, то про все розповіли, і про біснуватих.
MATT|8|34|І ось, усе місто вийшло назустріч Ісусові. Як Його ж угледіли, то стали благати, щоб пішов Собі з їхнього краю!..
MATT|9|1|І, сівши до човна, Він переплинув, і до міста Свого прибув.
MATT|9|2|І ото, принесли до Нього розслабленого, що на ложі лежав. І, як побачив Ісус їхню віру, сказав розслабленому: Будь бадьорий, сину! Прощаються тобі гріхи твої!
MATT|9|3|І ось, дехто із книжників стали казати про себе: Він богозневажає.
MATT|9|4|Ісус же думки їхні знав і сказав: Чого думаєте ви лукаве в серцях своїх?
MATT|9|5|Що легше, сказати: Прощаються тобі гріхи, чи сказати: Уставай та й ходи?
MATT|9|6|Але щоб ви знали, що прощати гріхи на землі має владу Син Людський, тож каже Він розслабленому: Уставай, візьми ложе своє, та й іди у свій дім!
MATT|9|7|Той устав і пішов у свій дім.
MATT|9|8|А натовп, побачивши це, налякався, і славив Бога, що людям Він дав таку владу!...
MATT|9|9|А коли Ісус звідти проходив, побачив чоловіка, на ймення Матвія, що сидів на митниці, та й каже йому: Іди за Мною! Той устав, і пішов услід за Ним.
MATT|9|10|І сталось, як Ісус сидів при столі у домі, ось зійшлося багато митників і грішників, і вони посідали з Ним та з Його учнями.
MATT|9|11|Як побачили ж те фарисеї, то сказали до учнів Його: Чому то Вчитель ваш їсть із митниками та із грішниками?
MATT|9|12|А Він це почув та й сказав: Лікаря не потребують здорові, а слабі!
MATT|9|13|Ідіть же, і навчіться, що то є: Милости хочу, а не жертви. Бо Я не прийшов кликати праведних, але грішників до покаяння.
MATT|9|14|Тоді приступили до Нього Іванові учні та й кажуть: Чому постимо ми й фарисеї, а учні Твої не постять?
MATT|9|15|Ісус же промовив до них: Хіба можуть гості весільні сумувати, поки з ними ще є молодий? Але прийдуть ті дні, коли заберуть молодого від них, тоді й постити будуть вони.
MATT|9|16|До одежі ж старої ніхто не вставляє латки з сукна сирового, бо збіжиться воно, і дірка стане ще гірша.
MATT|9|17|І не вливають вина молодого в старі бурдюки, а то бурдюки розірвуться, і вино розіллється, і бурдюки пропадуть; а вливають вино молоде до нових бурдюків, і одне й друге збережено буде.
MATT|9|18|Коли Він говорив це до них, підійшов ось один із старших, уклонився Йому та й говорить: Дочка моя хвилі цієї померла. Та прийди, поклади Свою руку на неї, і вона оживе.
MATT|9|19|І підвівся Ісус, і пішов услід за ним, також учні Його.
MATT|9|20|І ото одна жінка, що дванадцять літ хворою на кровотечу була, приступила ззаду, і доторкнулась до краю одежі Його.
MATT|9|21|Бо вона говорила про себе: Коли хоч доторкнуся одежі Його, то одужаю.
MATT|9|22|Ісус, обернувшись, побачив її та й сказав: Будь бадьорою, дочко, твоя віра спасла тебе! І одужала жінка з тієї години.
MATT|9|23|А Ісус, як прибув до господи старшого, і вздрів дударів та юрбу голосільників,
MATT|9|24|то сказав: Відійдіть, бо не вмерло дівча, але спить. І насміхалися з Нього.
MATT|9|25|А коли народ випроваджено, Він увійшов, узяв за руку її, і дівчина встала!
MATT|9|26|І вістка про це розійшлася по всій тій країні.
MATT|9|27|Коли ж Ісус звідти вертався, ішли за Ним два сліпці, що кричали й казали: Змилуйсь над нами, Сину Давидів!
MATT|9|28|І коли Він додому прийшов, приступили до Нього сліпці. А Ісус до них каже: Чи ж вірите ви, що Я можу вчинити оце? Говорять до Нього вони: Так, Господи.
MATT|9|29|Тоді Він доторкнувся до їхніх очей і сказав: Нехай станеться вам згідно з вашою вірою!
MATT|9|30|І очі відкрилися їм. А Ісус наказав їм суворо, говорячи: Глядіть, щоб ніхто не довідавсь про це!
MATT|9|31|А вони відійшли, та й розголосили про Нього по всій тій країні.
MATT|9|32|Коли ж ті виходили, то ось привели до Нього чоловіка німого, що був біснуватий.
MATT|9|33|І як демон був вигнаний, німий заговорив. І дивувався народ і казав: Ніколи таке не траплялося серед Ізраїля!
MATT|9|34|Фарисеї ж казали: Виганяє Він демонів силою князя демонів.
MATT|9|35|І обходив Ісус всі міста та оселі, навчаючи в їхніх синагогах, та Євангелію Царства проповідуючи, і вздоровлюючи всяку недугу та неміч усяку.
MATT|9|36|А як бачив людей, змилосерджувався Він над ними, бо були вони змучені та розпорошені, як ті вівці, що не мають пастуха.
MATT|9|37|Тоді Він казав Своїм учням: Жниво справді велике, та робітників мало;
MATT|9|38|тож благайте Господаря жнива, щоб на жниво Своє Він робітників вислав.
MATT|10|1|І закликав Він дванадцятьох Своїх учнів, і владу їм дав над нечистими духами, щоб їх виганяли вони, і щоб уздоровляли всіляку недугу та неміч всіляку.
MATT|10|2|А ймення апостолів дванадцятьох отакі: перший Симон, що Петром прозивається, і Андрій, брат його; Яків, син Зеведеїв, та Іван, брат його;
MATT|10|3|Пилип і Варфоломій, Хома й митник Матвій; Яків, син Алфеїв, і Тадей;
MATT|10|4|Симон Кананіт, та Юда Іскаріотський, що й видав Його.
MATT|10|5|Цих Дванадцятьох Ісус вислав, і їм наказав, промовляючи: На путь до поган не ходіть, і до самарянського міста не входьте,
MATT|10|6|але йдіть радніш до овечок загинулих дому Ізраїлевого.
MATT|10|7|А ходячи, проповідуйте та говоріть, що наблизилось Царство Небесне.
MATT|10|8|Уздоровляйте недужих, воскрешайте померлих, очищайте прокажених, виганяйте демонів. Ви дармо дістали, дармо й давайте.
MATT|10|9|Не беріть ані золота, ані срібла, ані мідяків до своїх поясів,
MATT|10|10|ані торби в дорогу, ані двох одеж, ні сандаль, ані палиці. Бо вартий робітник своєї поживи.
MATT|10|11|А як зайдете в місто якесь чи в село, то розвідайте, хто там достойний, і там перебудьте, аж поки не вийдете.
MATT|10|12|А входячи в дім, вітайте його, промовляючи: Мир дому цьому!
MATT|10|13|І коли буде достойний той дім, нехай зійде на нього ваш мир; а як недостойний він буде, то мир ваш нехай до вас вернеться.
MATT|10|14|А як хто вас не прийме, і ваших слів не послухає, то, виходячи з дому чи з міста того, обтрусіть порох із ніг своїх.
MATT|10|15|Поправді кажу вам: легше буде країні содомській й гоморській дня судного, аніж місту тому!
MATT|10|16|Оце посилаю Я вас, як овець між вовки. Будьте ж мудрі, як змії, і невинні, як голубки.
MATT|10|17|Стережіться ж людей, бо вони на суди видаватимуть вас, та по синагогах своїх бичувати вас будуть.
MATT|10|18|І до правителів та до царів поведуть вас за Мене, на свідчення їм і поганам.
MATT|10|19|А коли видаватимуть вас, не журіться, як або що говорити: тієї години буде вам дане, що маєте ви говорити,
MATT|10|20|бо не ви промовлятимете, але Дух Отця вашого в вас промовлятиме.
MATT|10|21|І видасть на смерть брата брат, а батько дитину. І діти повстануть супроти батьків, і їх повбивають.
MATT|10|22|І за Ім'я Моє будуть усі вас ненавидіти. А хто витерпить аж до кінця, той буде спасений.
MATT|10|23|А коли будуть вас переслідувати в однім місті, утікайте до іншого. Поправді кажу вам, не встигнете ви обійти міст Ізраїлевих, як прийде Син Людський.
MATT|10|24|Учень не більший за вчителя, а раб понад пана свого.
MATT|10|25|Доволі для учня, коли буде він, як учитель його, а раб як господар його. Коли Вельзевулом назвали господаря дому, скільки ж більше назвуть так домашніх його!
MATT|10|26|Але не лякайтеся їх. Немає нічого захованого, що воно не відкриється, ані потаємного, що не виявиться.
MATT|10|27|Що кажу Я вам потемки, говоріть те при світлі, що ж на вухо ви чуєте проповідуйте те на дахах.
MATT|10|28|І не лякайтеся тих, хто тіло вбиває, а душі вбити не може; але бійтеся більше того, хто може й душу, і тіло вам занапастити в геєнні.
MATT|10|29|Чи не два горобці продаються за гріш? А на землю із них ні один не впаде без волі Отця вашого.
MATT|10|30|А вам і волосся все на голові пораховано.
MATT|10|31|Отож, не лякайтесь, бо вартніші ви за багатьох горобців.
MATT|10|32|Отже, кожного, хто Мене визнає перед людьми, того перед Небесним Отцем Моїм визнаю й Я.
MATT|10|33|Хто ж Мене відцурається перед людьми, того й Я відцураюся перед Небесним Отцем Моїм.
MATT|10|34|Не думайте, що Я прийшов, щоб мир на землю принести, Я не мир принести прийшов, а меча.
MATT|10|35|Я ж прийшов порізнити чоловіка з батьком його, дочку з її матір'ю, і невістку з свекрухою її.
MATT|10|36|І: вороги чоловікові домашні його!
MATT|10|37|Хто більш, як Мене, любить батька чи матір, той Мене недостойний. І хто більш, як Мене, любить сина чи дочку, той Мене недостойний.
MATT|10|38|І хто не візьме свого хреста, і не піде за Мною слідом, той Мене недостойний.
MATT|10|39|Хто душу свою зберігає, той погубить її, хто ж за Мене погубить душу свою, той знайде її.
MATT|10|40|Хто вас приймає приймає Мене, хто ж приймає Мене, приймає Того, Хто послав Мене.
MATT|10|41|Хто приймає пророка, як пророка, той дістане нагороду пророчу, хто ж приймає праведника, як праведника, той дістане нагороду праведничу.
MATT|10|42|І хто напоїть, як учня, кого з малих цих бодай кухлем водиці холодної, поправді кажу вам, той не згубить нагороди своєї.
MATT|11|1|І сталось, коли Ісус перестав навчати дванадцятьох Своїх учнів, Він звідти пішов, щоб учити, і по їхніх містах проповідувати.
MATT|11|2|Прочувши ж Іван у в'язниці про дії Христові, послав через учнів своїх,
MATT|11|3|щоб Його запитати: Чи Ти Той, Хто має прийти, чи чекати нам Іншого?
MATT|11|4|Ісус же промовив у відповідь їм: Ідіть, і перекажіть Іванові, що ви чуєте й бачите:
MATT|11|5|Сліпі прозрівають, і криві ходять, стають чистими прокажені, і чують глухі, і померлі встають, а вбогим звіщається Добра Новина...
MATT|11|6|І блаженний, хто через Мене спокуси не матиме!
MATT|11|7|Як вони ж відійшли, Ісус про Івана почав говорити народові: На що ви ходили в пустиню дивитися? Чи на очерет, що вітер гойдає його?
MATT|11|8|Та на що ви дивитись ходили? Може на чоловіка, у м'які шати одягненого? Аджеж ті, хто носить м'яке, по палатах царських.
MATT|11|9|По що ж ви ходили? Може бачити пророка? Так, кажу вам, навіть більш, як пророка.
MATT|11|10|Бо це ж той, що про нього написано: Ось перед обличчя Твоє посилаю Свого посланця, який перед Тобою дорогу Твою приготує!
MATT|11|11|Поправді кажу вам: Між народженими від жінок не було більшого над Івана Христителя! Та найменший у Царстві Небеснім той більший від нього!
MATT|11|12|Від днів же Івана Христителя й досі Царство Небесне здобувається силою, і ті, хто вживає зусилля, хапають його.
MATT|11|13|Усі бо Пророки й Закон до Івана провіщували.
MATT|11|14|Коли ж хочете знати, то Ілля він, що має прийти.
MATT|11|15|Хто має вуха, нехай слухає!
MATT|11|16|До кого ж цей рід прирівняю? До хлоп'ят він подібний, що на ринку сидять та вигукують іншим,
MATT|11|17|і кажуть: Ми вам грали, а ви не танцювали, ми співали вам жалібно, та не плакали ви...
MATT|11|18|Бо прийшов був Іван, що не їв і не пив, вони ж кажуть: Він демона має.
MATT|11|19|Прийшов же Син Людський, що їсть і п'є, вони ж кажуть: Чоловік ось, ласун і п'яниця, Він приятель митників і грішників. І виправдалася мудрість своїми ділами.
MATT|11|20|Ісус тоді став докоряти містам, де відбулося найбільш Його чуд, що вони не покаялись:
MATT|11|21|Горе тобі, Хоразіне, горе тобі, Віфсаїдо! Бо коли б то в Тирі й Сидоні були відбулися ті чуда, що сталися в вас, то давно б вони каялися в волосяниці та в попелі.
MATT|11|22|Але кажу вам: Легше буде дня судного Тиру й Сидону, ніж вам!
MATT|11|23|А ти, Капернауме, що до неба піднісся, аж до аду ти зійдеш. Бо коли б у Содомі були відбулися ті чуда, що в тобі вони стались, то лишився б він був по сьогоднішній день.
MATT|11|24|Але кажу вам, що содомській землі буде легше дня судного, аніж тобі!...
MATT|11|25|Того часу, навчаючи, промовив Ісус: Прославляю Тебе, Отче, Господи неба й землі, що втаїв Ти оце від премудрих і розумних, та його немовлятам відкрив.
MATT|11|26|Так, Отче, бо Тобі так було до вподоби!
MATT|11|27|Передав Мені все Мій Отець. І Сина не знає ніхто, крім Отця, і Отця не знає ніхто, окрім Сина, та кому Син захоче відкрити.
MATT|11|28|Прийдіть до Мене, усі струджені та обтяжені, і Я вас заспокою!
MATT|11|29|Візьміть на себе ярмо Моє, і навчіться від Мене, бо Я тихий і серцем покірливий, і знайдете спокій душам своїм.
MATT|11|30|Бож ярмо Моє любе, а тягар Мій легкий!
MATT|12|1|Того часу Ісус переходив ланами в суботу. А учні Його зголодніли були, і стали зривати колосся та їсти.
MATT|12|2|Побачили ж це фарисеї, та й кажуть Йому: Он учні Твої роблять те, чого не годиться робити в суботу...
MATT|12|3|А Він відповів їм: Чи ж ви не читали, що зробив був Давид, коли сам зголоднів і ті, хто був із ним?
MATT|12|4|Як він увійшов до Божого дому, і спожив хліби показні, яких їсти не можна було ні йому, ані тим, хто був із ним, а тільки самим священикам?
MATT|12|5|Або ви не читали в Законі що в суботу священики порушують суботу у храмі, і невинні вони?
MATT|12|6|А Я вам кажу, що тут Більший, як храм!
MATT|12|7|Коли б знали ви, що то є: Милости хочу, а не жертви, то ви не судили б невинних...
MATT|12|8|Бо Син Людський Господь і суботі!
MATT|12|9|І, вийшовши звідти, прибув Він до їхньої синагоги.
MATT|12|10|І ото, був там чоловік, що мав суху руку. І, щоб обвинити Ісуса, запитали Його: Чи вздоровляти годиться в суботу?
MATT|12|11|А Він їм сказав: Чи знайдеться між вами людина, яка, одну мавши вівцю, не піде по неї, і не врятує її, як вона впаде в яму в суботу?
MATT|12|12|А скільки ж людина вартніша за тую овечку! Тому можна чинити добро й у суботу!
MATT|12|13|І каже тоді чоловікові: Простягни свою руку! Той простяг, і стала здорова вона, як і друга...
MATT|12|14|Фарисеї ж пішли, і зібрали нараду на Нього, як би Його погубити?...
MATT|12|15|А Ісус, розізнавши, пішов Собі звідти. І багато пішло вслід за Ним, і Він їх уздоровив усіх.
MATT|12|16|А Він наказав їм суворо Його не виявляти,
MATT|12|17|щоб справдилось те, що сказав був Ісая пророк, промовляючи:
MATT|12|18|Ото Мій Отрок, що Я вибрав Його, Мій Улюблений, що Його полюбила душа Моя! Вкладу Свого Духа в Нього, і Він суд проголосить поганам.
MATT|12|19|Він не буде змагатися, ані кричати, і на вулицях чути не буде ніхто Його голосу.
MATT|12|20|Він очеретини надломленої не доломить, і ґнота догасаючого не погасить, поки не допровадить присуду до перемоги...
MATT|12|21|І погани надіятись будуть на Ймення Його!
MATT|12|22|Тоді привели до Нього німого сліпця, що був біснуватий, і Він уздоровив його, так що німий став говорити та бачити.
MATT|12|23|І дивувались усі люди й казали: Чи ж не Син це Давидів?
MATT|12|24|Фарисеї ж, почувши, сказали: Він демонів не виганяє інакше, тільки як Вельзевулом, князем демонів.
MATT|12|25|А Він знав думки їхні, і промовив до них: Кожне царство, поділене супроти себе, запустіє. І кожне місто чи дім, поділені супроти себе, не втримаються.
MATT|12|26|І коли сатана сатану виганяє, то ділиться супроти себе; як же втримається царство його?
MATT|12|27|І коли Вельзевулом виганяю Я демонів, то ким виганяють сини ваші? Тому вони стануть вам суддями.
MATT|12|28|А коли ж Духом Божим вигоню Я демонів, то настало для вас Царство Боже.
MATT|12|29|Або як то хто може вдертися в дім дужого, та пограбувати добро його, якщо перше не зв'яже дужого? І аж тоді він господу його пограбує.
MATT|12|30|Хто не зо Мною, той супроти Мене; і хто не збирає зо Мною, той розкидає.
MATT|12|31|Тому то кажу вам: усякий гріх, навіть богозневага, проститься людям, але богозневага на Духа не проститься!
MATT|12|32|І як скаже хто слово на Людського Сина, то йому проститься те; а коли скаже проти Духа Святого, не проститься того йому ані в цім віці, ані в майбутнім!
MATT|12|33|Або виростіть дерево добре, то й плід його добрий, або виростіть дерево зле, то й плід його злий. Пізнається бо дерево з плоду!
MATT|12|34|Роде зміїний! Як ви можете мовити добре, бувши злі? Бо чим серце наповнене, те говорять уста.
MATT|12|35|Добра людина з доброго скарбу добре виносить, а лукава людина зо скарбу лихого виносить лихе.
MATT|12|36|Кажу ж вам, що за кожне слово пусте, яке скажуть люди, дадуть вони відповідь судного дня!
MATT|12|37|Бо зо слів своїх будеш виправданий, і зо слів своїх будеш засуджений.
MATT|12|38|Тоді дехто із книжників та фарисеїв озвались до Нього й сказали: Учителю, хочемо побачити ознаку від Тебе.
MATT|12|39|А Ісус відповів їм: Рід лукавий і перелюбний шукає ознаки, та ознаки йому не дадуть, окрім ознаки пророка Йони.
MATT|12|40|Як Йона перебув у середині китовій три дні і три ночі, так перебуде три дні та три ночі й Син Людський у серці землі.
MATT|12|41|Ніневітяни стануть на суд із цим родом, і осудять його, вони бо покаялися через Йонину проповідь. А тут ото Більший, ніж Йона!
MATT|12|42|Цариця з півдня на суд стане з родом оцим, і засудить його, бо вона з кінця світу прийшла Соломонову мудрість послухати. А тут ото Більший, аніж Соломон!
MATT|12|43|А коли дух нечистий виходить із людини, то блукає місцями безвідними, відпочинку шукаючи, та не знаходить.
MATT|12|44|Тоді він говорить: Вернуся до дому свого, звідки вийшов. А як вернеться він, то хату знаходить порожню, заметену й прибрану.
MATT|12|45|Тоді він іде, та й приводить сімох духів інших, лютіших за себе, і входять вони та й живуть тут. І буде останнє людині тій гірше за перше... Так буде й лукавому родові цьому!
MATT|12|46|Коли Він іще промовляв до народу, аж ось мати й брати Його осторонь стали, бажаючи з Ним говорити.
MATT|12|47|І сказав хтось Йому: Ото мати Твоя й Твої браття стоять онде осторонь, і говорити з Тобою бажають.
MATT|12|48|А Він відповів тому, хто Йому говорив, і сказав: Хто мати Моя? І хто браття Мої?
MATT|12|49|І, показавши рукою Своєю на учнів Своїх, Він промовив: Ото Моя мати та браття Мої!
MATT|12|50|Бо хто волю Мого Отця, що на небі, чинитиме, той Мені брат, і сестра, і мати!
MATT|13|1|Того ж дня Ісус вийшов із дому, та й сів біля моря.
MATT|13|2|І безліч народу зібралась до Нього, так що Він увійшов був до човна та й сів, а ввесь натовп стояв понад берегом.
MATT|13|3|І багато навчав Він їх притчами, кажучи: Ось вийшов сіяч, щоб посіяти.
MATT|13|4|І як сіяв він зерна, упали одні край дороги, і пташки налетіли, та їх повидзьобували.
MATT|13|5|Другі ж упали на ґрунт кам'янистий, де не мали багато землі, і негайно посходили, бо земля неглибока була;
MATT|13|6|а як сонце зійшло, то зів'яли, і коріння не мавши, посохли.
MATT|13|7|А інші попадали в терен, і вигнався терен, і їх поглушив.
MATT|13|8|Інші ж упали на добрую землю і зродили: одне в сто раз, друге в шістдесят, а те втридцятеро.
MATT|13|9|Хто має вуха, щоб слухати, нехай слухає!
MATT|13|10|І учні Його приступили й сказали до Нього: Чому притчами Ти промовляєш до них?
MATT|13|11|А Він відповів і промовив: Тому, що вам дано пізнати таємниці Царства Небесного, їм же не дано.
MATT|13|12|Бо хто має, то дасться йому та додасться, хто ж не має, забереться від нього й те, що він має.
MATT|13|13|Я тому говорю до них притчами, що вони, дивлячися, не бачать, і слухаючи, не чують, і не розуміють.
MATT|13|14|І над ними збувається пророцтво Ісаї, яке промовляє: Почуєте слухом, і не зрозумієте, дивитися будете оком, і не побачите...
MATT|13|15|Затовстіло бо серце людей цих, тяжко чують вухами вони, і зажмурили очі свої, щоб коли не побачити очима й не почути вухами, і не зрозуміти їм серцем, і не навернутись, щоб Я їх уздоровив!
MATT|13|16|Очі ж ваші блаженні, що бачать, і вуха ваші, що чують.
MATT|13|17|Бо поправді кажу вам, що багато пророків і праведних бажали побачити, що бачите ви, та не бачили, і почути, що чуєте ви, і не чули.
MATT|13|18|Послухайте ж притчу про сіяча.
MATT|13|19|До кожного, хто слухає слово про Царство, але не розуміє, приходить лукавий, і краде посіяне в серці його; це те, що посіяне понад дорогою.
MATT|13|20|А посіяне на кам'янистому ґрунті, це той, хто слухає слово, і з радістю зараз приймає його;
MATT|13|21|але кореня в ньому нема, тому він непостійний; коли ж утиск або переслідування настають за слово, то він зараз спокушується.
MATT|13|22|А між терен посіяне, це той, хто слухає слово, але клопоти віку цього та омана багатства заглушують слово, і воно зостається без плоду.
MATT|13|23|А посіяне в добрій землі, це той, хто слухає слово й його розуміє, і плід він приносить, і дає один у сто раз, другий у шістдесят, а той утридцятеро.
MATT|13|24|Іншу притчу подав Він їм, кажучи: Царство Небесне подібне до чоловіка, що посіяв був добре насіння на полі своїм.
MATT|13|25|А коли люди спали, прийшов ворог його, і куколю між пшеницю насіяв, та й пішов.
MATT|13|26|А як виросло збіжжя та кинуло колос, тоді показався і кукіль.
MATT|13|27|І прийшли господареві раби, та й кажуть йому: Пане, чи ж не добре насіння ти сіяв на полі своїм? Звідки ж узявся кукіль?
MATT|13|28|А він їм відказав: Чоловік супротивник накоїв оце. А раби відказали йому: Отож, чи не хочеш, щоб пішли ми і його повиполювали?
MATT|13|29|Але він відказав: Ні, щоб, виполюючи той кукіль, ви не вирвали разом із ним і пшеницю.
MATT|13|30|Залишіть, хай разом обоє ростуть аж до жнив; а в жнива накажу я женцям: Зберіть перше кукіль і його пов'яжіть у снопки, щоб їх попалити; пшеницю ж спровадьте до клуні моєї.
MATT|13|31|Іншу притчу подав Він їм, кажучи: Царство Небесне подібне до зерна гірчичного, що взяв чоловік і посіяв на полі своїм.
MATT|13|32|Воно найдрібніше з увсього насіння, але, коли виросте, більше воно за зілля, і стає деревом, так що птаство небесне злітається, і кублиться в віттях його.
MATT|13|33|Іншу притчу Він їм розповів: Царство Небесне подібне до розчини, що її бере жінка, і кладе на три мірі муки, аж поки все вкисне.
MATT|13|34|Це все в притчах Ісус говорив до людей, і без притчі нічого Він їм не казав,
MATT|13|35|щоб справдилось те, що сказав був пророк, промовляючи: Відкрию у притчах уста Свої, розповім таємниці від почину світу!
MATT|13|36|Тоді відпустив Він народ і додому прийшов. І підійшли Його учні до Нього й сказали: Поясни нам притчу про кукіль польовий.
MATT|13|37|А Він відповів і промовив до них: Хто добре насіння посіяв був, це Син Людський,
MATT|13|38|а поле це світ, добре ж насіння це сини Царства, а кукіль сини лукавого;
MATT|13|39|а ворог, що всіяв його це диявол, жнива кінець віку, а женці Анголи.
MATT|13|40|І як збирають кукіль, і як палять в огні, так буде й наприкінці віку цього.
MATT|13|41|Пошле Людський Син Своїх Анголів, і вони позбирають із Царства Його всі спокуси, і тих, хто чинить беззаконня,
MATT|13|42|і їх повкидають до печі огненної, буде там плач і скрегіт зубів!
MATT|13|43|Тоді праведники, немов сонце, засяють у Царстві свого Отця. Хто має вуха, нехай слухає!
MATT|13|44|Царство Небесне подібне ще до захованого в полі скарбу, що людина, знайшовши, ховає його, і з радости з того йде, та й усе, що має, продає та купує те поле.
MATT|13|45|Подібне ще Царство Небесне до того купця, що пошукує перел добрих,
MATT|13|46|а як знайде одну дорогоцінну перлину, то йде, і все продає, що має, і купує її.
MATT|13|47|Подібне ще Царство Небесне до невода, у море закиненого, що зібрав він усячину.
MATT|13|48|Коли він наповниться, тягнуть на берег його, і, сівши, вибирають до посуду добре, непотріб же геть викидають.
MATT|13|49|Так буде й наприкінці віку: Анголи повиходять, і вилучать злих з-поміж праведних,
MATT|13|50|і їх повкидають до печі огненної, буде там плач і скрегіт зубів!
MATT|13|51|Чи ви зрозуміли це все? Так! відказали Йому.
MATT|13|52|І Він їм сказав: Тому кожен книжник, що навчений про Царство Небесне, подібний до того господаря, що з скарбниці своєї виносить нове та старе.
MATT|13|53|І сталось, як скінчив Ісус притчі оці, Він звідти пішов.
MATT|13|54|І прийшов Він до Своєї батьківщини, і навчав їх у їхній синагозі, так що стали вони дивуватися й питати: Звідки в Нього ця мудрість та сили чудодійні?
MATT|13|55|Чи ж Він не син теслі? Чи ж мати Його не Марією зветься, а брати Його Яків, і Йосип, і Симон та Юда?
MATT|13|56|І чи ж сестри Його не всі з нами? Звідки ж Йому все оте?
MATT|13|57|І вони спокушалися Ним. А Ісус їм сказав: Пророка нема без пошани, хіба тільки в вітчизні своїй та в домі своїм!
MATT|13|58|І Він не вчинив тут чуд багатьох через їхню невіру.
MATT|14|1|Того часу прочув Ірод чотиривласник чутки про Ісуса,
MATT|14|2|і сказав своїм слугам: Це Іван Христитель, він із мертвих воскрес, і тому чуда творяться ним...
MATT|14|3|Бо Ірод схопив був Івана, і зв'язав його, і посадив у в'язницю через Іродіяду, дружину брата свого Пилипа.
MATT|14|4|Бо до нього Іван говорив: Не годиться тобі її мати!
MATT|14|5|І хотів Ірод смерть заподіяти йому, та боявся народу, бо того за пророка вважали.
MATT|14|6|А як був день народження Ірода, танцювала посеред гостей дочка Іродіядина, та й Іродові догодила.
MATT|14|7|Тому під присягою він обіцявся їй дати, чого тільки попросить вона.
MATT|14|8|А вона, за намовою матері своєї: Дай мені проказала отут на полумиску голову Івана Христителя!...
MATT|14|9|І цар засмутився, але через клятву та тих, хто сидів при столі з ним, звелів дати.
MATT|14|10|І послав стяти Івана в в'язниці.
MATT|14|11|І принесли на полумискові його голову, та й дали дівчині, а та віднесла її своїй матері...
MATT|14|12|А учні його прибули, взяли тіло, і поховали його, та прийшли й сповістили Ісуса.
MATT|14|13|Як Ісус те почув, Він відплив звідти човном у місце пустинне й самотнє. І, прочувши, народ із міст пішов пішки за Ним.
MATT|14|14|І, як вийшов Ісус, Він побачив багато народу, і змилосердивсь над ними, і їхніх слабих уздоровив.
MATT|14|15|А коли настав вечір, підійшли Його учні до Нього й сказали: Тут місце пустинне, і година вже пізня; відпусти народ, хай по селах розійдуться, і куплять поживи собі.
MATT|14|16|А Ісус їм сказав: Непотрібно відходити їм, нагодуйте їх ви!
MATT|14|17|Вони ж кажуть Йому: Не маємо чим тут, тільки п'ятеро хліба й дві рибі.
MATT|14|18|А Він відказав: Принесіть Мені їх сюди.
MATT|14|19|І, звелівши натовпові посідати на траві, Він узяв п'ятеро хліба й дві рибі, споглянув на небо, поблагословив й поламав ті хліби, і дав учням, а учні народові.
MATT|14|20|І всі їли й наситились, а з кусків позосталих назбирали дванадцятеро повних кошів...
MATT|14|21|Їдців же було мужа тисяч із п'ять, крім жінок і дітей.
MATT|14|22|І зараз звелів Ісус учням до човна сідати, і переплисти на той бік раніше Його, аж поки народ Він відпустить.
MATT|14|23|Відпустивши ж народ, Він на гору пішов помолитися насамоті; і як вечір настав, був там Сам.
MATT|14|24|А човен вже був на середині моря, і кидали хвилі його, бо вітер зірвавсь супротивний.
MATT|14|25|А о четвертій сторожі нічній Ісус підійшов до них, ідучи по морю.
MATT|14|26|Як побачили ж учні, що йде Він по морю, то настрашилися та й казали: Мара! І від страху вони закричали...
MATT|14|27|А Ісус до них зараз озвався й сказав: Заспокойтесь, це Я, не лякайтесь!
MATT|14|28|Петро ж відповів і сказав: Коли, Господи, Ти це, то звели, щоб прийшов я до Тебе по воді.
MATT|14|29|А Він відказав йому: Іди. І, вилізши з човна, Петро став іти по воді, і пішов до Ісуса.
MATT|14|30|Але, бачачи велику бурю, злякався, і зачав потопати, і скричав: Рятуй мене, Господи!...
MATT|14|31|І зараз Ісус простяг руку й схопив його, і каже до нього: Маловірний, чого усумнився?
MATT|14|32|Як до човна ж вони ввійшли, буря вщухнула.
MATT|14|33|А приявні в човні вклонились Йому та сказали: Ти справді Син Божий!
MATT|14|34|Перепливши ж вони, прибули в землю Генісаретську.
MATT|14|35|А люди тієї місцевости, пізнавши Його, сповістили по всій тій околиці, і до Нього принесли всіх хворих.
MATT|14|36|І благали Його, щоб бодай доторкнутися краю одежі Його. А хто доторкавсь, уздоровлений був.
MATT|15|1|Тоді до Ісуса прийшли фарисеї та книжники з Єрусалиму й сказали:
MATT|15|2|Чого Твої учні ламають передання старших? Бо не миють вони своїх рук, коли хліб споживають.
MATT|15|3|А Він відповів і промовив до них: А чого й ви порушуєте Божу заповідь ради передання вашого?
MATT|15|4|Бо Бог заповів: Шануй батька та матір, та: Хто злорічить на батька чи матір, хай смертю помре.
MATT|15|5|А ви кажете: Коли скаже хто батьку чи матері: Те, чим би ви скористатись від мене хотіли, то дар Богові,
MATT|15|6|то може вже й не шанувати той батька свого або матір свою. Так ви ради передання вашого знівечили Боже Слово.
MATT|15|7|Лицеміри! Про вас добре Ісая пророкував був, говорячи:
MATT|15|8|Оці люди устами шанують Мене, серце ж їхнє далеко від Мене!
MATT|15|9|Та однак надаремне шанують Мене, бо навчають наук людських заповідей...
MATT|15|10|І Він покликав народ, і промовив до нього: Послухайте та зрозумійте!
MATT|15|11|Не те, що входить до уст, людину сквернить, але те, що виходить із уст, те людину сквернить.
MATT|15|12|Тоді учні Його приступили й сказали Йому: Чи Ти знаєш, що фарисеї, почувши це слово, спокусилися?
MATT|15|13|А Він відповів і сказав: Усяка рослина, яку насадив не Отець Мій Небесний, буде вирвана з коренем.
MATT|15|14|Залишіть ви їх: це сліпі поводатарі для сліпих. А коли сліпий водить сліпого, обоє до ями впадуть...
MATT|15|15|А Петро відповів і до Нього сказав: Поясни нам цю притчу.
MATT|15|16|А Він відказав: Чи ж і ви розуміння не маєте?
MATT|15|17|Чи ж ви не розумієте, що все те, що входить до уст, вступає в живіт, та й назовні виходить?
MATT|15|18|Що ж виходить із уст, те походить із серця, і воно опоганює людину.
MATT|15|19|Бо з серця виходять лихі думки, душогубства, перелюби, розпуста, крадіж, неправдиві засвідчення, богозневаги.
MATT|15|20|Оце те, що людину опоганює. А їсти руками невмитими, не опоганює це людини!
MATT|15|21|І, вийшовши звідти, Ісус відійшов у землі тирські й сидонські.
MATT|15|22|І ось жінка одна хананеянка, із тих околиць прийшовши, заголосила до Нього й сказала: Змилуйся надо мною, Господи, Сину Давидів, демон тяжко дочку мою мучить!
MATT|15|23|А Він їй не казав ані слова. Тоді учні Його, підійшовши, благали Його та казали: Відпусти її, бо кричить услід за нами!
MATT|15|24|А Він відповів і сказав: Я посланий тільки до овечок загинулих дому Ізраїлевого...
MATT|15|25|А вона, підійшовши, уклонилась Йому та й сказала: Господи, допоможи мені!
MATT|15|26|А Він відповів і сказав: Не годиться взяти хліб у дітей, і кинути щенятам...
MATT|15|27|Вона ж відказала: Так, Господи! Але ж і щенята їдять ті кришки, що спадають зо столу їхніх панів.
MATT|15|28|Тоді відповів і сказав їй Ісус: О жінко, твоя віра велика, нехай буде тобі, як ти хочеш! І тієї години дочка її видужала.
MATT|15|29|І, відійшовши звідти, Ісус прибув до Галілейського моря, і, зійшовши на гору, сів там.
MATT|15|30|І приступило до Нього багато народу, що мали з собою кривих, калік, сліпих, німих і інших багато, і клали їх до Ісусових ніг. І Він уздоровлював їх.
MATT|15|31|А народ не виходив із дива, бо бачив, що говорять німі, каліки стають здорові, криві ходять, і бачать сліпі, і славив він Бога Ізраїлевого!
MATT|15|32|А Ісус Своїх учнів покликав і сказав: Жаль Мені цих людей, що вже три дні зо Мною знаходяться, але їсти не мають чого; відпустити їх без їжі не хочу, щоб вони не ослабли в дорозі.
MATT|15|33|А учні Йому відказали: Де нам узяти стільки хліба в пустині, щоб нагодувати стільки народу?
MATT|15|34|А Ісус запитав їх: Скільки маєте хліба? Вони ж відказали: Семеро, та трохи рибок.
MATT|15|35|І Він ізвелів на землі посідати народові.
MATT|15|36|І, взявши сім хлібів і риби, віддавши Богу подяку, поламав і дав учням Своїм, а учні народові.
MATT|15|37|І всі їли й наситилися, а з позосталих кусків назбирали сім кошиків повних...
MATT|15|38|Їдців же було чотири тисячі мужа, окрім жінок та дітей.
MATT|15|39|І, відпустивши народ, усів Він до човна, і прибув до землі Магдалинської.
MATT|16|1|І підійшли фарисеї та саддукеї, і, випробовуючи, просили Його показати ознаку їм із неба.
MATT|16|2|А Він відповів і промовив до них: Ви звечора кажете: Буде погода, червоніє бо небо.
MATT|16|3|А ранком: Сьогодні негода, червоніє бо небо похмуре. Розпізнати небесне обличчя ви вмієте, ознак часу ж не можете!
MATT|16|4|Рід лукавий і перелюбний шукає ознаки, та ознаки йому не дадуть, окрім ознаки пророка Йони. І, їх полишивши, Він відійшов.
MATT|16|5|А учні Його, перейшовши на той бік, забули взяти хліба.
MATT|16|6|Ісус же промовив до них: Стережіться уважливо фарисейської та саддукейської розчини!
MATT|16|7|Вони ж міркували собі й говорили: Ми ж хлібів не взяли.
MATT|16|8|А Ісус, знавши те, запитав: Чого між собою міркуєте ви, маловірні, що хлібів не взяли?
MATT|16|9|Чи ж ви ще не розумієте й не пам'ятаєте про п'ять хлібів на п'ять тисяч, і скільки кошів ви зібрали?
MATT|16|10|Ані про сім хлібів на чотири тисячі, і скільки кошиків ви назбирали?
MATT|16|11|Як ви не розумієте, що Я не про хліб вам сказав? Стережіться но розчини фарисейської та саддукейської!
MATT|16|12|Тоді зрозуміли вони, що Він не казав стерегтися їм розчини хлібної, але фарисейської та саддукейської науки.
MATT|16|13|Прийшовши ж Ісус до землі Кесарії Пилипової, питав Своїх учнів і казав: За кого народ уважає Мене, Сина Людського?
MATT|16|14|Вони ж відповіли: Одні за Івана Христителя, одні за Іллю, інші ж за Єремію або за одного з пророків.
MATT|16|15|Він каже до них: А ви за кого Мене маєте?
MATT|16|16|А Симон Петро відповів і сказав: Ти Христос, Син Бога Живого!
MATT|16|17|А Ісус відповів і до нього промовив: Блаженний ти, Симоне, сину Йонин, бо не тіло і кров тобі оце виявили, але Мій Небесний Отець.
MATT|16|18|І кажу Я тобі, що ти скеля, і на скелі оцій побудую Я Церкву Свою, і сили адові не переможуть її.
MATT|16|19|І ключі тобі дам від Царства Небесного, і що на землі ти зв'яжеш, те зв'язане буде на небі, а що на землі ти розв'яжеш, те розв'язане буде на небі!
MATT|16|20|Тоді наказав Своїм учням, щоб нікому не казали, що Він Христос.
MATT|16|21|Із того часу Ісус став виказувати Своїм учням, що Він мусить іти до Єрусалиму, і постраждати багато від старших, і первосвящеників, і книжників, і вбитому бути, і воскреснути третього дня.
MATT|16|22|І, набік відвівши Його, Петро став Йому докоряти й казати: Змилуйся, Господи, такого Тобі хай не буде!
MATT|16|23|А Він обернувся й промовив Петрові: Відступися від Мене, сатано, ти спокуса Мені, бо думаєш не про Боже, а про людське!
MATT|16|24|Промовив тоді Ісус учням Своїм: Коли хоче хто йти вслід за Мною, хай зречеться самого себе, і хай візьме свого хреста, та й іде вслід за Мною.
MATT|16|25|Бо хто хоче спасти свою душу, той погубить її, хто ж за Мене свою душу погубить, той знайде її.
MATT|16|26|Яка ж користь людині, що здобуде ввесь світ, але душу свою занапастить? Або що дасть людина взамін за душу свою?
MATT|16|27|Бо прийде Син Людський у славі Свого Отця з Анголами Своїми, і тоді віддасть кожному згідно з ділами його.
MATT|16|28|Поправді кажу вам, що деякі з тут-о приявних не скуштують смерти, аж поки не побачать Сина Людського, що йде в Царстві Своїм.
MATT|17|1|А через шість день забирає Ісус Петра, і Якова, і Івана, брата його, та й веде їх осібно на гору високу.
MATT|17|2|І Він перед ними переобразився: обличчя Його, як те сонце, засяло, а одежа Його стала біла, як світло.
MATT|17|3|І ось з'явились до них Мойсей та Ілля, і розмовляли із Ним.
MATT|17|4|І озвався Петро та й сказав до Ісуса: Господи, добре бути нам тут! Коли хочеш, поставлю отут три шатрі: для Тебе одне, і одне для Мойсея, і одне для Іллі.
MATT|17|5|Як він ще говорив, ось хмара ясна заслонила їх, і ось голос із хмари почувсь, що казав: Це Син Мій Улюблений, що Його Я вподобав. Його слухайтеся!
MATT|17|6|А почувши, попадали учні долілиць, і полякалися сильно...
MATT|17|7|А Ісус підійшов, доторкнувся до них і промовив: Уставайте й не бійтесь!
MATT|17|8|Звівши ж очі свої, нікого вони не побачили, окрім Самого Ісуса.
MATT|17|9|А коли з гори сходили, заповів їм Ісус і сказав: Не кажіть нікому про цеє видіння, аж поки Син Людський із мертвих воскресне.
MATT|17|10|І запитали Його учні, говорячи: Що це книжники кажуть, ніби треба Іллі перш прийти?
MATT|17|11|А Він відповів і сказав: Ілля, правда, прийде, і все приготує.
MATT|17|12|Але кажу вам, що Ілля вже прийшов був, та його не пізнали, але з ним зробили, що тільки хотіли... Так і Син Людський має страждати від них.
MATT|17|13|Учні тоді зрозуміли, що Він їм говорив про Івана Христителя.
MATT|17|14|І як вони до народу прийшли, то до Нього один чоловік приступив, і навколішки впав перед Ним,
MATT|17|15|і сказав: Господи, змилуйсь над сином моїм, що біснується у новомісяччі, і мучиться тяжко, бо почасту падає він ув огонь, і почасту в воду.
MATT|17|16|Я його був привів до учнів Твоїх, та вони не могли вздоровити його.
MATT|17|17|А Ісус відповів і сказав: О роде невірний й розбещений, доки буду Я з вами? Доки вас Я терпітиму? Приведіть до Мене сюди його!
MATT|17|18|Потому Ісус погрозив йому, і демон вийшов із нього. І видужав хлопець тієї години!
MATT|17|19|Тоді підійшли учні насамоті до Ісуса й сказали: Чому ми не могли його вигнати?
MATT|17|20|А Він їм відповів: Через ваше невірство. Бо поправді кажу вам: коли будете ви мати віру, хоч як зерно гірчичне, і горі оцій скажете: Перейди звідси туди, то й перейде вона, і нічого не матимете неможливого!
MATT|17|21|Цей же рід не виходить інакше, як тільки молитвою й постом.
MATT|17|22|Коли пробували вони в Галілеї, то сказав їм Ісус: Людський Син буде виданий людям до рук,
MATT|17|23|і вони Його вб'ють, але третього дня Він воскресне. І тяжко вони зажурились...
MATT|17|24|Як прийшли ж вони в Капернаум, до Петра підійшли збирачі дидрахм на храм, та й сказали: Чи не заплатить ваш учитель дидрахми?
MATT|17|25|Він відказує: Так. І як він увійшов до дому, то Ісус попередив його та сказав: Як ти думаєш, Симоне: царі земні з кого беруть мито або податки: від синів своїх, чи чужих?
MATT|17|26|А як той відказав: Від чужих, то промовив до нього Ісус: Тож вільні сини!
MATT|17|27|Та щоб їх не спокусити, піди над море, та вудку закинь, і яку першу рибу ізловиш, візьми, і рота відкрий їй, і знайдеш статира; візьми ти його, і віддай їм за Мене й за себе...
MATT|18|1|Підійшли до Ісуса тоді Його учні, питаючи: Хто найбільший у Царстві Небеснім?
MATT|18|2|Він же дитину покликав, і поставив її серед них,
MATT|18|3|та й сказав: Поправді кажу вам: коли не навернетесь, і не станете, як ті діти, не ввійдете в Царство Небесне!
MATT|18|4|Отже, хто впокориться, як дитина оця, той найбільший у Царстві Небеснім.
MATT|18|5|І хто прийме таку дитину одну в Моє Ймення, той приймає Мене.
MATT|18|6|Хто ж спокусить одне з цих малих, що вірують в Мене, то краще б такому було, коли б жорно млинове на шию йому почепити, і його потопити в морській глибині...
MATT|18|7|Від спокус горе світові, бо мусять спокуси прийти; надто горе людині, що від неї приходить спокуса!
MATT|18|8|Коли тільки рука твоя, чи нога твоя спокушає тебе, відітни її й кинь від себе: краще тобі увійти в життя одноруким або одноногим, ніж з обома руками чи з обома ногами бути вкиненому в огонь вічний.
MATT|18|9|І коли твоє око тебе спокушає його вибери й кинь від себе: краще тобі однооким ввійти в життя, ніж з обома очима бути вкиненому до геєнни огненної.
MATT|18|10|Стережіться, щоб ви не погордували ані одним із малих цих; кажу бо Я вам, що їхні Анголи повсякчасно бачать у небі обличчя Мого Отця, що на небі.
MATT|18|11|Син бо Людський прийшов, щоб спасти загинуле.
MATT|18|12|Як вам здається: коли має який чоловік сто овець, а одна з них заблудить, то чи він не покине дев'ятдесятьох і дев'ятьох у горах, і не піде шукати заблудлої?
MATT|18|13|І коли пощастить відшукати її, поправді кажу вам, що радіє за неї він більше, аніж за дев'ятдесятьох і дев'ятьох незаблудлих.
MATT|18|14|Так волі нема Отця вашого, що на небі, щоб загинув один із цих малих.
MATT|18|15|А коли прогрішиться твій брат проти тебе, іди й йому викажи поміж тобою та ним самим; як тебе він послухає, ти придбав свого брата.
MATT|18|16|А коли не послухає він, то візьми з собою ще одного чи двох, щоб справа всіляка ствердилась устами двох чи трьох свідків.
MATT|18|17|А коли не послухає їх, скажи Церкві; коли ж не послухає й Церкви, хай буде тобі, як поганин і митник!
MATT|18|18|Поправді кажу вам: Що тільки зв'яжете на землі, зв'язане буде на небі, і що тільки розв'яжете на землі, розв'язане буде на небі.
MATT|18|19|Ще поправді кажу вам, що коли б двоє з вас на землі погодились про всяку річ, то коли вони будуть просити за неї, станеться їм від Мого Отця, що на небі!
MATT|18|20|Бо де двоє чи троє в Ім'я Моє зібрані, там Я серед них.
MATT|18|21|Петро приступив тоді та запитався Його: Господи, скільки разів брат мій може згрішити проти мене, а я маю прощати йому? Чи до семи раз?
MATT|18|22|Ісус промовляє до нього: Не кажу тобі до семи раз, але аж до семидесяти раз по семи!
MATT|18|23|Тим то Царство Небесне подібне одному цареві, що захотів обрахунок зробити з своїми рабами.
MATT|18|24|Коли ж він почав обраховувати, то йому привели одного, що винен був десять тисяч талантів.
MATT|18|25|А що він не мав із чого віддати, наказав пан продати його, і його дружину та діти, і все, що він мав, і заплатити.
MATT|18|26|Тоді раб той упав до ніг, і вклонявся йому та благав: Потерпи мені, я віддам тобі все!
MATT|18|27|І змилосердився пан над рабом тим, і звільнив його, і простив йому борг.
MATT|18|28|А як вийшов той раб, то спіткав він одного з своїх співтоваришів, що був винен йому сто динаріїв. І, схопивши його, він душив та казав: Віддай, що ти винен!
MATT|18|29|А товариш його впав у ноги йому, і благав його, кажучи: Потерпи мені, і я віддам тобі!
MATT|18|30|Та той не схотів, а пішов і всадив до в'язниці його, аж поки він боргу не верне.
MATT|18|31|Як побачили ж товариші його те, що сталося, то засмутилися дуже, і прийшли й розповіли своєму панові все, що було.
MATT|18|32|Тоді пан його кличе його, та й говорить до нього: Рабе лукавий, я простив був тобі ввесь той борг, бо просив ти мене.
MATT|18|33|Чи й тобі не належало змилуватись над своїм співтоваришем, як і я над тобою був змилувався?
MATT|18|34|І прогнівався пан його, і катам його видав, аж поки йому не віддасть всього боргу.
MATT|18|35|Так само й Отець Мій Небесний учинить із вами, коли кожен із вас не простить своєму братові з серця свого їхніх прогріхів.
MATT|19|1|І сталось, як Ісус закінчив ці слова, то Він вирушив із Галілеї, і прибув до країни Юдейської, на той бік Йордану.
MATT|19|2|А за Ним ішла безліч народу, і Він уздоровив їх тут.
MATT|19|3|І підійшли фарисеї до Нього, і, випробовуючи, запитали Його: Чи дозволено дружину свою відпускати з причини всякої?
MATT|19|4|А Він відповів і сказав: Чи ви не читали, що Той, Хто створив споконвіку людей, створив їх чоловіком і жінкою?
MATT|19|5|І сказав: Покине тому чоловік батька й матір, і пристане до дружини своєї, і стануть обоє вони одним тілом,
MATT|19|6|тому то немає вже двох, але одне тіло. Тож, що Бог спарував, людина нехай не розлучує!
MATT|19|7|Вони кажуть Йому: А чому ж Мойсей заповів дати листа розводового, та й відпускати?
MATT|19|8|Він говорить до них: То за ваше жорстокосердя дозволив Мойсей відпускати дружин ваших, спочатку ж так не було.
MATT|19|9|А Я вам кажу: Хто дружину відпустить свою не з причини перелюбу, і одружиться з іншою, той чинить перелюб. І хто одружиться з розведеною, той чинить перелюб.
MATT|19|10|Учні говорять Йому: Коли справа така чоловіка із дружиною, то не добре одружуватись.
MATT|19|11|А Він їм відказав: Це слово вміщають не всі, але ті, кому дано.
MATT|19|12|Бо бувають скопці, що з утроби ще матерньої народилися так; є й скопці, що їх люди оскопили, і є скопці, що самі оскопили себе ради Царства Небесного. Хто може вмістити, нехай вмістить.
MATT|19|13|Тоді привели Йому діток, щоб поклав на них руки, і за них помолився, учні ж їм докоряли.
MATT|19|14|Ісус же сказав: Пустіть діток, і не бороніть їм приходити до Мене, бо Царство Небесне належить таким.
MATT|19|15|І Він руки на них поклав, та й пішов звідтіля.
MATT|19|16|І підійшов ось один, і до Нього сказав: Учителю Добрий, що маю зробити я доброго, щоб мати життя вічне?
MATT|19|17|Він же йому відказав: Чого звеш Мене Добрим? Ніхто не є Добрий, крім Бога Самого. Коли ж хочеш ввійти до життя, то виконай заповіді.
MATT|19|18|Той питає Його: Які саме? А Ісус відказав: Не вбивай, не чини перелюбу, не кради, не свідкуй неправдиво.
MATT|19|19|Шануй батька та матір, і: Люби свого ближнього, як самого себе.
MATT|19|20|Говорить до Нього юнак: Це я виконав все. Чого ще бракує мені?
MATT|19|21|Ісус каже йому: Коли хочеш бути досконалим, піди, продай добра свої та й убогим роздай, і матимеш скарб ти на небі. Потому приходь та й іди вслід за Мною.
MATT|19|22|Почувши ж юнак таке слово, відійшов, зажурившись, бо великі маєтки він мав.
MATT|19|23|Ісус же сказав Своїм учням: Поправді кажу вам, що багатому трудно ввійти в Царство Небесне.
MATT|19|24|Іще вам кажу: Верблюдові легше пройти через голчине вушко, ніж багатому в Боже Царство ввійти!
MATT|19|25|Як учні ж Його це зачули, здивувалися дуже й сказали: Хто ж тоді може спастися?
MATT|19|26|А Ісус позирнув і сказав їм: Неможливе це людям, та можливе все Богові.
MATT|19|27|Тоді відізвався Петро та до Нього сказав: От усе ми покинули, та й пішли за Тобою слідом; що ж нам буде за це?
MATT|19|28|А Ісус відказав їм: Поправді кажу вам, що коли, при відновленні світу, Син Людський засяде на престолі слави Своєї, тоді сядете й ви, що за Мною пішли, на дванадцять престолів, щоб судити дванадцять племен Ізраїлевих.
MATT|19|29|І кожен, хто за Ймення Моє кине дім, чи братів, чи сестер, або батька, чи матір, чи діти, чи землі, той багатокротно одержить і успадкує вічне життя.
MATT|19|30|І багато-хто з перших останніми стануть, а останні першими.
MATT|20|1|Бо Царство Небесне подібне одному господареві, що вдосвіта вийшов згодити робітників у свій виноградник.
MATT|20|2|Згодившися ж він із робітниками по динарію за день, послав їх до свого виноградника.
MATT|20|3|А вийшовши коло години десь третьої, побачив він інших, що стояли без праці на ринку,
MATT|20|4|та й каже до них: Ідіть і ви до мого виноградника, і що буде належати, дам вам.
MATT|20|5|Вони ж відійшли. І вийшов він знов о годині десь шостій й дев'ятій, і те саме зробив.
MATT|20|6|А вийшовши коло години одинадцятої, знайшов інших, що стояли без праці, та й каже до них: Чого тут стоїте цілий день безробітні?
MATT|20|7|Вони кажуть до нього: Бо ніхто не найняв нас. Відказує їм: Ідіть і ви в виноградник.
MATT|20|8|Коли ж вечір настав, то говорить тоді до свого управителя пан виноградника: Поклич робітників, і дай їм заплату, почавши з останніх до перших.
MATT|20|9|І прийшли ті, що з години одинадцятої, і взяли по динарію.
MATT|20|10|Коли ж прийшли перші, то думали, що вони візьмуть більше. Та й вони по динару взяли.
MATT|20|11|А взявши, вони почали нарікати на господаря,
MATT|20|12|кажучи: Ці останні годину одну працювали, а ти прирівняв їх до нас, що витерпіли тягар дня та спекоту...
MATT|20|13|А він відповів і сказав до одного із них: Не кривджу я, друже, тебе, хіба не за динарія згодився зо мною?
MATT|20|14|Візьми ти своє та й іди. Але я хочу дати й цьому ось останньому, як і тобі.
MATT|20|15|Чи ж не вільно мені зо своїм, що я хочу, зробити? Хіба око твоє заздре від того, що я добрий?
MATT|20|16|Отак будуть останні першими, а перші останніми!
MATT|20|17|Побажавши ж піти до Єрусалиму, Ісус взяв осібно Дванадцятьох, і на дорозі їм сповістив:
MATT|20|18|Оце в Єрусалим ми йдемо, і первосвященикам і книжникам виданий буде Син Людський, і засудять на смерть Його...
MATT|20|19|І посганам Його вони видадуть на наругу та на катування, і на розп'яття, але третього дня Він воскресне!
MATT|20|20|Тоді приступила до Нього мати синів Зеведеєвих, і вклонилась, і просила від Нього чогось.
MATT|20|21|А Він їй сказав: Чого хочеш? Вона каже Йому: Скажи, щоб обидва сини мої ці сіли в Царстві Твоїм праворуч один, і ліворуч від Тебе один.
MATT|20|22|А Ісус відповів і сказав: Не знаєте, чого просите. Чи ж можете ви пити чашу, що Я її питиму або христитися хрищенням, що я ним хрищуся? Вони кажуть Йому: Можемо.
MATT|20|23|Він говорить до них: Ви питимете Мою чашу і будете христитися хрищенням, що Я ним хрищуся. А сидіти праворуч Мене та ліворуч не Моє це давати, а кому від Мого Отця те вготовано.
MATT|20|24|Як почули це десятеро, стали гніватися на обох тих братів.
MATT|20|25|А Ісус їх покликав і промовив: Ви знаєте, що князі народів панують над ними, а вельможі їх тиснуть.
MATT|20|26|Не так буде між вами, але хто великим із вас хоче бути, хай буде слугою він вам.
MATT|20|27|А хто з вас бути першим бажає, нехай буде він вам за раба.
MATT|20|28|Так само й Син Людський прийшов не на те, щоб служили Йому, а щоб послужити, і душу Свою дати на викуп за багатьох!
MATT|20|29|Як вони ж з Єрихону виходили, за Ним ішов натовп великий.
MATT|20|30|І ось двоє сліпих, що сиділи при дорозі, почувши, що переходить Ісус, стали кричати, благаючи: Змилуйсь над нами, Господи, Сину Давидів!
MATT|20|31|Народ же сварився на них, щоб мовчали, вони ж іще більше кричали, благаючи: Змилуйсь над нами, Господи, Сину Давидів!
MATT|20|32|Ісус же спинився, покликав їх та й сказав: Що хочете, щоб Я вам зробив?
MATT|20|33|Вони Йому кажуть: Господи, нехай нам розкриються очі!
MATT|20|34|І змилосердивсь Ісус, доторкнувся до їхніх очей, і зараз прозріли їм очі, і вони подалися за Ним.
MATT|21|1|А коли вони наблизились до Єрусалиму, і прийшли до Вітфагії, до гори до Оливної, тоді Ісус вислав двох учнів,
MATT|21|2|до них, кажучи: Ідіть у село, яке перед вами, і знайдете зараз ослицю прив'язану та з нею осля; відв'яжіть, і Мені приведіть їх.
MATT|21|3|А як хто вам що скаже, відкажіть, що їх потребує Господь, і він зараз пошле їх.
MATT|21|4|А це сталось, щоб справдилось те, що сказав був пророк, промовляючи:
MATT|21|5|Скажіте Сіонській доньці: Ось до тебе йде Цар твій! Він покірливий, і всів на осла, на осля, під'яремної сина.
MATT|21|6|А учні пішли та й зробили, як звелів їм Ісус.
MATT|21|7|Вони привели до Ісуса ослицю й осля, і одежу поклали на них, і Він сів на них.
MATT|21|8|І багато народу стелили одежу свою по дорозі, інші ж різали віття з дерев і стелили дорогою.
MATT|21|9|А народ, що йшов перед Ним і позаду, викрикував, кажучи: Осанна Сину Давидовому! Благословенний, хто йде у Господнє Ім'я! Осанна на висоті!
MATT|21|10|А коли увійшов Він до Єрусалиму, то здвигнулося ціле місто, питаючи: Хто це такий?
MATT|21|11|А народ говорив: Це Пророк, Ісус із Назарету Галілейського!
MATT|21|12|Потому Ісус увійшов у храм Божий, і вигнав усіх продавців і покупців у храмі, і поперевертав грошомінам столи, та ослони продавцям голубів.
MATT|21|13|І сказав їм: Написано: Дім Мій буде домом молитви, а ви робите з нього печеру розбійників.
MATT|21|14|І приступили у храмі до Нього сліпі та криві, і Він їх уздоровив.
MATT|21|15|А первосвященики й книжники, бачивши чуда, що Він учинив, і дітей, що в храмі викрикували: Осанна Сину Давидовому, обурилися,
MATT|21|16|та й сказали Йому: Чи ти чуєш, що кажуть вони? А Ісус відказав їм: Так. Чи ж ви не читали ніколи: Із уст немовлят, і тих, що ссуть, учинив Ти хвалу?
MATT|21|17|І покинувши їх, Він вийшов за місто в Віфанію, і там ніч перебув.
MATT|21|18|А вранці, до міста вертаючись, Він зголоднів.
MATT|21|19|І побачив Він при дорозі одне фіґове дерево, і до нього прийшов, та нічого, крім листя самого, на нім не знайшов. І до нього Він каже: Нехай плоду із тебе не буде ніколи повіки! І фіґове дерево зараз усохло.
MATT|21|20|А учні, побачивши це, дивувалися та говорили: Як швидко всохло це фіґове дерево!...
MATT|21|21|Ісус же промовив у відповідь їм: Поправді кажу вам: Коли б мали ви віру, і не мали сумніву, то вчинили б не тільки як із фіґовим деревом, а якби й цій горі ви сказали: Порушся та кинься до моря, то й станеться те!
MATT|21|22|І все, чого ви в молитві попросите з вірою, то одержите.
MATT|21|23|А коли Він прийшов у храм і навчав, поприходили первосвященики й старші народу до Нього й сказали: Якою Ти владою чиниш оце? І хто Тобі владу цю дав?
MATT|21|24|Ісус же промовив у відповідь їм: Запитаю й Я вас одне слово. Як про нього дасте Мені відповідь, то й Я вам скажу, якою владою Я це чиню.
MATT|21|25|Іванове хрищення звідки було: із неба, чи від людей? Вони ж міркували собі й говорили: Коли скажемо: Із неба, відкаже Він нам: Чого ж ви йому не повірили?
MATT|21|26|А як скажемо: Від людей, боїмося народу, бо Івана вважають усі за пророка.
MATT|21|27|І сказали Ісусові в відповідь: Ми не знаємо. Відказав їм і Він: То й Я вам не скажу, якою владою Я це чиню.
MATT|21|28|А як вам здається? Один чоловік мав двох синів. Прийшовши до першого, він сказав: Піди но, дитино, сьогодні, працюй у винограднику!
MATT|21|29|А той відповів і сказав: Готовий, панотче, і не пішов.
MATT|21|30|І, прийшовши до другого, так само сказав. А той відповів і сказав: Я не хочу. А потім покаявся, і пішов.
MATT|21|31|Котрий же з двох учинив волю батькову? Вони кажуть: Останній. Ісус промовляє до них: Поправді кажу вам, що митники та блудодійки випереджують вас у Боже Царство.
MATT|21|32|Бо прийшов був до вас дорогою праведности Іван, та йому не повірили ви, а митники та блудодійки йняли йому віри. А ви бачили, та проте не покаялися й опісля, щоб повірити йому.
MATT|21|33|Послухайте іншої притчі. Був господар один. Насадив виноградника він, обгородив його муром, видовбав у ньому чавило, башту поставив, і віддав його винарям, та й пішов.
MATT|21|34|Коли ж надійшов час плодів, він до винарів послав рабів своїх, щоб прийняти плоди свої.
MATT|21|35|Винарі ж рабів його похапали, і одного побили, а другого замордували, а того вкаменували.
MATT|21|36|Знов послав він інших рабів, більш як перше, та й їм учинили те саме.
MATT|21|37|Нарешті послав до них сина свого і сказав: Посоромляться сина мого.
MATT|21|38|Але винарі, як побачили сина, міркувати собі стали: Це спадкоємець; ходім, замордуймо його, і заберемо його спадщину!
MATT|21|39|І, схопивши його, вони вивели за виноградник його, та й убили.
MATT|21|40|Отож, як прибуде той пан виноградника, що зробить він тим винарям?
MATT|21|41|Вони кажуть Йому: Злочинців погубить жорстоко, виноградника ж віддасть іншим винарям, що будуть плоди віддавати йому своєчасно.
MATT|21|42|Ісус промовляє до них: Чи ви не читали ніколи в Писанні: Камінь, що його будівничі відкинули, той наріжним став каменем; від Господа сталося це, і дивне воно в очах наших!
MATT|21|43|Тому кажу вам, що від вас Царство Боже відійметься, і дасться народові, що плоди його буде приносити.
MATT|21|44|І хто впаде на цей камінь розіб'ється, а на кого він сам упаде то розчавить його.
MATT|21|45|А як первосвященики та фарисеї почули ці притчі Його, то вони зрозуміли, що про них Він говорить.
MATT|21|46|І намагались схопити Його, але побоялись людей, бо вважали Його за Пророка.
MATT|22|1|А Ісус, відповідаючи, знов почав говорити їм притчами, кажучи:
MATT|22|2|Царство Небесне подібне одному цареві, що весілля справляв був для сина свого.
MATT|22|3|І послав він своїх рабів покликати тих, хто був на весілля запрошений, та ті не хотіли прийти.
MATT|22|4|Знову послав він інших рабів, наказуючи: Скажіть запрошеним: Ось я приготував обід свій, закололи бики й відгодоване, і все готове. Ідіть на весілля!
MATT|22|5|Та вони злегковажили та порозходились, той на поле своє, а той на свій торг.
MATT|22|6|А останні, похапавши рабів його, знущалися, та й повбивали їх.
MATT|22|7|І розгнівався цар, і послав своє військо, і вигубив тих убійників, а їхнє місто спалив.
MATT|22|8|Тоді каже рабам своїм: Весілля готове, але недостойні були ті покликані.
MATT|22|9|Тож підіть на роздоріжжя, і кого тільки спіткаєте, кличте їх на весілля.
MATT|22|10|І вийшовши раби ті на роздоріжжя, зібрали всіх, кого тільки спіткали, злих і добрих. І весільна кімната гістьми переповнилась.
MATT|22|11|Як прийшов же той цар на гостей подивитись, побачив там чоловіка, в одежу весільну не вбраного,
MATT|22|12|та й каже йому: Як ти, друже, ввійшов сюди, не мавши одежі весільної? Той же мовчав.
MATT|22|13|Тоді цар сказав своїм слугам: Зв'яжіть йому ноги та руки, та й киньте до зовнішньої темряви, буде плач там і скрегіт зубів...
MATT|22|14|Бо багато покликаних, та вибраних мало.
MATT|22|15|Тоді фарисеї пішли й умовлялись, як зловити на слові Його.
MATT|22|16|І посилають до Нього своїх учнів із іродіянами, і кажуть: Учителю, знаємо ми, що Ти справедливий, і наставляєш на Божу дорогу правдиво, і не зважаєш ні на кого, бо на людське обличчя не дивишся Ти.
MATT|22|17|Скажи ж нам, як здається Тобі: чи годиться давати податок для кесаря, чи ні?
MATT|22|18|А Ісус, знавши їхнє лукавство, сказав: Чого ви, лицеміри, Мене випробовуєте?
MATT|22|19|Покажіть Мені гріш податковий. І принесли динарія Йому.
MATT|22|20|А Він каже до них: Чий це образ і напис?
MATT|22|21|Ті відказують: Кесарів. Тоді каже Він їм: Тож віддайте кесареве кесареві, а Богові Боже.
MATT|22|22|А почувши таке, вони диву далися. І, лишивши Його, відійшли.
MATT|22|23|Того дня приступили до Нього саддукеї, що твердять, ніби нема воскресення, і запитали Його,
MATT|22|24|та й сказали: Учителю, Мойсей наказав: Коли хто помре, не мавши дітей, то нехай його брат візьме вдову його, і відновить насіння для брата свого.
MATT|22|25|Було ж у нас сім братів. І перший, одружившись, умер, і, не мавши насіння, зоставив дружину свою братові своєму.
MATT|22|26|Так само і другий, і третій, аж до сьомого.
MATT|22|27|А по всіх вмерла й жінка.
MATT|22|28|Отож, у воскресенні котрому з сімох вона дружиною буде? Бо всі мали її.
MATT|22|29|Ісус же промовив у відповідь їм: Помиляєтесь ви, не знавши писання, ні Божої сили.
MATT|22|30|Бо в воскресенні ні женяться, ані заміж виходять, але як Анголи ті на небі.
MATT|22|31|А про воскресення померлих хіба не читали прореченого вам від Бога, що каже:
MATT|22|32|Я Бог Авраамів, і Бог Ісаків, і Бог Яковів; Бог не є Богом мертвих, а живих.
MATT|22|33|А народ, чувши це, дивувався науці Його.
MATT|22|34|Фарисеї ж, почувши, що Він уста замкнув саддукеям, зібралися разом.
MATT|22|35|І спитався один із них, учитель Закону, Його випробовуючи й кажучи:
MATT|22|36|Учителю, котра заповідь найбільша в Законі?
MATT|22|37|Він же промовив йому: Люби Господа Бога свого всім серцем своїм, і всією душею своєю, і всією своєю думкою.
MATT|22|38|Це найбільша й найперша заповідь.
MATT|22|39|А друга однакова з нею: Люби свого ближнього, як самого себе.
MATT|22|40|На двох оцих заповідях увесь Закон і Пророки стоять.
MATT|22|41|Коли ж фарисеї зібрались, Ісус їх запитав,
MATT|22|42|і сказав: Що ви думаєте про Христа? Чий Він син? Вони Йому кажуть: Давидів.
MATT|22|43|Він до них промовляє: Як же то силою Духа Давид Його Господом зве, коли каже:
MATT|22|44|Промовив Господь Господеві моєму: сядь праворуч Мене, доки не покладу Я Твоїх ворогів підніжком ногам Твоїм.
MATT|22|45|Тож, коли Давид зве Його Господом, як же Він йому син?
MATT|22|46|І ніхто не спромігся відповісти Йому ані слова... І ніхто з того дня не наважувався більш питати Його.
MATT|23|1|Тоді промовив Ісус до народу й до учнів Своїх,
MATT|23|2|і сказав: На сидінні Мойсеєвім усілися книжники та фарисеї.
MATT|23|3|Тож усе, що вони скажуть вам, робіть і виконуйте; та за вчинками їхніми не робіть, бо говорять вони та не роблять того!
MATT|23|4|Вони ж в'яжуть тяжкі тягарі, і кладуть їх на людські рамена, самі ж навіть пальцем своїм не хотять їх порушити...
MATT|23|5|Усі ж учинки свої вони роблять, щоб їх бачили люди, і богомілля свої розширяють, і здовжують китиці.
MATT|23|6|І люблять вони передніші місця на бенкетах, і передніші лавки в синагогах,
MATT|23|7|і привіти на ринках, і щоб звали їх люди: Учителю!
MATT|23|8|А ви вчителями не звіться, бо один вам Учитель, а ви всі брати.
MATT|23|9|І не називайте нікого отцем на землі, бо один вам Отець, що на небі.
MATT|23|10|І не звіться наставниками, бо один вам Наставник, Христос.
MATT|23|11|Хто між вами найбільший, хай слугою вам буде!
MATT|23|12|Хто бо підноситься, буде понижений, хто ж понижується, той піднесеться.
MATT|23|13|Горе ж вам, книжники та фарисеї, лицеміри, що перед людьми зачиняєте Царство Небесне, бо й самі ви не входите, ані тих, хто хоче ввійти, увійти не пускаєте!
MATT|23|14|Горе ж вам, книжники та фарисеї, лицеміри, що вдовині хати поїдаєте, і напоказ молитесь довго, через те осуд тяжчий ви приймете!
MATT|23|15|Горе вам, книжники та фарисеї, лицеміри, що обходите море та землю, щоб придбати нововірця одного; а коли те стається, то робите його сином геєнни, вдвоє гіршим від вас!
MATT|23|16|Горе вам, проводирі ви сліпі, що говорите: Коли хто поклянеться храмом, то нічого; а хто поклянеться золотом храму, то той винуватий.
MATT|23|17|Нерозумні й сліпі, що бо більше: чи золото, чи той храм, що освячує золото?
MATT|23|18|І: Коли хто поклянеться жертівником, то нічого, а хто поклянеться жертвою, що на нім, то він винуватий.
MATT|23|19|Нерозумні й сліпі, що бо більше: чи жертва, чи той жертівник, що освячує жертву?
MATT|23|20|Отож, хто клянеться жертівником, клянеться ним та всім, що на ньому.
MATT|23|21|І хто храмом клянеться, клянеться ним та Тим, Хто живе в нім.
MATT|23|22|І хто небом клянеться, клянеться Божим престолом і Тим, Хто на ньому сидить.
MATT|23|23|Горе вам, книжники та фарисеї, лицеміри, що даєте десятину із м'яти, і ганусу й кмину, але найважливіше в Законі покинули: суд, милосердя та віру; це треба робити, і того не кидати.
MATT|23|24|Проводирі ви сліпі, що відціджуєте комаря, а верблюда ковтаєте!
MATT|23|25|Горе вам, книжники та фарисеї, лицеміри, що чистите зовнішність кухля та миски, а всередині повні вони здирства й кривди!
MATT|23|26|Фарисею сліпий, очисти перше середину кухля, щоб чистий він був і назовні!
MATT|23|27|Горе вам, книжники та фарисеї, лицеміри, що подібні до гробів побілених, які гарними зверху здаються, а всередині повні трупних кісток та всякої нечистости!
MATT|23|28|Так і ви, назовні здаєтеся людям за праведних, а всередині повні лицемірства та беззаконня!
MATT|23|29|Горе вам, книжники та фарисеї, лицеміри, що пророкам надгробники ставите, і праведникам прикрашаєте пам'ятники,
MATT|23|30|та говорите: Якби ми жили за днів наших батьків, то ми не були б спільниками їхніми в крові пророків.
MATT|23|31|Тим самим на себе свідкуєте, що сини ви убивців пророків.
MATT|23|32|Доповніть і ви міру провини ваших батьків!
MATT|23|33|О змії, о роде гадючий, як ви втечете від засуду до геєнни?
MATT|23|34|І ось тому посилаю до вас Я пророків, і мудрих, і книжників; частину їх ви повбиваєте та розіпнете, а частину їх ви бичуватимете в синагогах своїх, і будете гнати з міста до міста.
MATT|23|35|Щоб спала на вас уся праведна кров, що пролита була на землі, від крови Авеля праведного, аж до крови Захарія, Варахіїного сина, що ви замордували його між храмом і жертівником!
MATT|23|36|Поправді кажу вам: Оце все спаде на рід цей!
MATT|23|37|Єрусалиме, Єрусалиме, що вбиваєш пророків та каменуєш посланих до тебе! Скільки разів Я хотів зібрати діти твої, як та квочка збирає під крила курчаток своїх, та ви не захотіли!
MATT|23|38|Ось ваш дім залишається порожній для вас!
MATT|23|39|Говорю бо Я вам: Відтепер ви Мене не побачите, аж поки не скажете: Благословенний, Хто йде у Господнє Ім'я!
MATT|24|1|І вийшов Ісус і від храму пішов. І підійшли Його учні, щоб Йому показати будинки храмові.
MATT|24|2|Він же промовив у відповідь їм: Чи бачите ви все оце? Поправді кажу вам: Не залишиться тут навіть камінь на камені, який не зруйнується!...
MATT|24|3|Коли ж Він сидів на Оливній горі, підійшли Його учні до Нього самотньо й спитали: Скажи нам, коли станеться це? І яка буде ознака приходу Твого й кінця віку?
MATT|24|4|Ісус же промовив у відповідь їм: Стережіться, щоб вас хто не звів!
MATT|24|5|Бо багато хто прийде в Ім'я Моє, кажучи: Я Христос. І зведуть багатьох.
MATT|24|6|Ви ж про війни почуєте, і про воєнні чутки, глядіть, не лякайтесь, бо статись належить тому. Але це не кінець ще.
MATT|24|7|Бо повстане народ на народ, і царство на царство, і голод, мор та землетруси настануть місцями.
MATT|24|8|А все це початок терпінь породільних.
MATT|24|9|На муки тоді видаватимуть вас, і вбиватимуть вас, і вас будуть ненавидіти всі народи за Ймення Моє.
MATT|24|10|І багато-хто в той час спокусяться, і видавати один одного будуть, і один одного будуть ненавидіти.
MATT|24|11|Постане багато фальшивих пророків, і зведуть багатьох.
MATT|24|12|І через розріст беззаконства любов багатьох охолоне.
MATT|24|13|А хто витерпить аж до кінця, той буде спасений!
MATT|24|14|І проповідана буде ця Євангелія Царства по цілому світові, на свідоцтво народам усім. І тоді прийде кінець!
MATT|24|15|Тож, коли ви побачите ту гидоту спустошення, що про неї звіщав був пророк Даниїл, на місці святому, хто читає, нехай розуміє,
MATT|24|16|тоді ті, хто в Юдеї, нехай в гори втікають.
MATT|24|17|Хто на покрівлі, нехай той не сходить узяти речі з дому свого.
MATT|24|18|І хто на полі, хай назад не вертається взяти одежу свою.
MATT|24|19|Горе ж вагітним і тим, хто годує грудьми, за днів тих!
MATT|24|20|Моліться ж, щоб ваша втеча не сталась зимою, ані в суботу.
MATT|24|21|Бо скорбота велика настане тоді, якої не було з первопочину світу аж досі й не буде.
MATT|24|22|І коли б не вкоротились ті дні, не спаслася б ніяка людина; але через вибраних дні ті вкоротяться.
MATT|24|23|Тоді, як хто скаже до вас: Ото, Христос тут чи Отам, не йміть віри.
MATT|24|24|Бо постануть христи неправдиві, і неправдиві пророки, і будуть чинити великі ознаки та чуда, що звели б, коли б можна, і вибраних.
MATT|24|25|Оце Я наперед вам сказав.
MATT|24|26|А коли скажуть вам: Ось Він у пустині не виходьте, Ось Він у криївках не вірте!
MATT|24|27|Бо як блискавка та вибігає зо сходу, і з'являється аж до заходу, так буде і прихід Сина Людського.
MATT|24|28|Бо де труп, там зберуться орли.
MATT|24|29|І зараз, по скорботі тих днів, сонце затьмиться, і місяць не дасть свого світла, і зорі попадають з неба, і сили небесні порушаться.
MATT|24|30|І того часу на небі з'явиться знак Сина Людського, і тоді заголосять всі земні племена, і побачать вони Сина Людського, що йтиме на хмарах небесних із великою потугою й славою.
MATT|24|31|І пошле Анголів Своїх Він із голосним сурмовим гуком, і зберуть Його вибраних від вітрів чотирьох, від кінців неба аж до кінців його.
MATT|24|32|Від дерева ж фіґового навчіться прикладу: коли віття його вже розпукується, і кинеться листя, то ви знаєте, що близько вже літо.
MATT|24|33|Так і ви: коли все це побачите, знайте, що близько, під дверима!
MATT|24|34|Поправді кажу вам: не перейде цей рід, аж усе оце станеться.
MATT|24|35|Небо й земля проминеться, але не минуться слова Мої!
MATT|24|36|А про день той й годину не знає ніхто: ані Анголи небесні, ані Син, лише Сам Отець.
MATT|24|37|Як було за днів Ноєвих, так буде і прихід Сина Людського.
MATT|24|38|Бо так само, як за днів до потопу всі їли й пили, женилися й заміж виходили, аж до дня, коли Ной увійшов до ковчегу,
MATT|24|39|і не знали, аж поки потоп не прийшов та й усіх не забрав, так буде і прихід Сина Людського.
MATT|24|40|Будуть двоє на полі тоді, один візьметься, а другий полишиться.
MATT|24|41|Дві будуть молоти на жорнах, одна візьметься, а друга полишиться.
MATT|24|42|Тож пильнуйте, бо не знаєте, котрого дня прийде Господь ваш.
MATT|24|43|Знайте ж це, що коли б знав господар, о котрій сторожі прийде злодій, то він пильнував би, і підкопати свого дому не дав би.
MATT|24|44|Тому будьте готові й ви, бо прийде Син Людський тієї години, коли ви не думаєте!
MATT|24|45|Хто ж вірний і мудрий раб, якого пан поставив над своїми челядниками давати своєчасно поживу для них?
MATT|24|46|Блаженний той раб, що пан його прийде та знайде, що робить він так!
MATT|24|47|Поправді кажу вам, що над цілим маєтком своїм він поставить його.
MATT|24|48|А як той злий раб скаже у серці своїм: Забариться пан мій прийти,
MATT|24|49|і зачне бити товаришів своїх, а їсти та пити з п'яницями,
MATT|24|50|то пан того раба прийде дня, якого він не сподівається, і о годині, якої не знає.
MATT|24|51|І він пополовині розітне його, і визначить долю йому з лицемірами, буде плач там і скрегіт зубів!
MATT|25|1|Тоді Царство Небесне буде подібне до десяти дів, що побрали каганці свої, та й пішли зустрічати молодого.
MATT|25|2|П'ять же з них нерозумні були, а п'ять мудрі.
MATT|25|3|Нерозумні ж, узявши каганці, не взяли із собою оливи.
MATT|25|4|А мудрі набрали оливи в посудинки разом із своїми каганцями.
MATT|25|5|А коли забаривсь молодий, то всі задрімали й поснули.
MATT|25|6|А опівночі крик залунав: Ось молодий, виходьте назустріч!
MATT|25|7|Схопились тоді всі ті діви, і каганці свої наготували.
MATT|25|8|Нерозумні ж сказали до мудрих: Дайте нам із своєї оливи, бо наші каганці ось гаснуть.
MATT|25|9|Мудрі ж відповіли та сказали: Щоб, бува, нам і вам не забракло, краще вдайтеся до продавців, і купіть собі.
MATT|25|10|І як вони купувати пішли, то прибув молодий; і готові ввійшли на весілля з ним, і замкнені двері були.
MATT|25|11|А потім прийшла й решта дів і казала: Пане, пане, відчини нам!
MATT|25|12|Він же в відповідь їм проказав: Поправді кажу вам, не знаю я вас!
MATT|25|13|Тож пильнуйте, бо не знаєте ні дня, ні години, коли прийде Син Людський!
MATT|25|14|Так само ж один чоловік, як відходив, покликав своїх рабів і передав їм добро своє.
MATT|25|15|І одному він дав п'ять талантів, а другому два, а тому один, кожному за спроможністю його. І відійшов.
MATT|25|16|А той, що взяв п'ять талантів, негайно пішов і орудував ними, і набув він п'ять інших талантів.
MATT|25|17|Так само ж і той, що взяв два і він ще два інших набув.
MATT|25|18|А той, що одного взяв, пішов та й закопав його в землю, і сховав срібло пана свого.
MATT|25|19|По довгому ж часі вернувся пан тих рабів, та й від них зажадав обрахунку.
MATT|25|20|І прийшов той, що взяв п'ять талантів, приніс іще п'ять талантів і сказав: Пане мій, п'ять талантів мені передав ти, ось я здобув інші п'ять талантів.
MATT|25|21|Сказав же йому його пан: Гаразд, рабе добрий і вірний! Ти в малому був вірний, над великим поставлю тебе, увійди до радощів пана свого!
MATT|25|22|Підійшов же й той, що взяв два таланти, і сказав: Два таланти мені передав ти, ось іще два таланти здобув я.
MATT|25|23|казав йому пан його: Гаразд, рабе добрий і вірний! Ти в малому був вірний, над великим поставлю тебе, увійди до радощів пана свого!
MATT|25|24|Підійшов же і той, що одного таланта взяв, і сказав: Я знав тебе, пане, що тверда ти людина, ти жнеш, де не сіяв, і збираєш, де не розсипав.
MATT|25|25|І я побоявся, пішов і таланта твого сховав у землю. Ото маєш своє...
MATT|25|26|І відповів його пан і сказав йому: Рабе лукавий і лінивий! Ти знав, що я жну, де не сіяв, і збираю, де не розсипав?
MATT|25|27|Тож тобі було треба віддати гроші мої грошомінам, і, вернувшись, я взяв би з прибутком своє.
MATT|25|28|Візьміть же від нього таланта, і віддайте тому, що десять талантів він має.
MATT|25|29|Бо кожному, хто має, дасться йому та й додасться, хто ж не має, забереться від нього й те, що він має.
MATT|25|30|А раба непотрібного вкиньте до зовнішньої темряви, буде плач там і скрегіт зубів!
MATT|25|31|Коли ж прийде Син Людський у славі Своїй, і всі Анголи з Ним, тоді Він засяде на престолі слави Своєї.
MATT|25|32|І перед Ним усі народи зберуться, і Він відділить одного від одного їх, як відділяє вівчар овець від козлів.
MATT|25|33|І поставить Він вівці праворуч Себе, а козлята ліворуч.
MATT|25|34|Тоді скаже Цар тим, хто праворуч Його: Прийдіть, благословенні Мого Отця, посядьте Царство, уготоване вам від закладин світу.
MATT|25|35|Бо Я голодував був і ви нагодували Мене, прагнув і ви напоїли Мене, мандрівником Я був і Мене прийняли ви.
MATT|25|36|Був нагий і Мене зодягли ви, слабував і Мене ви відвідали, у в'язниці Я був і прийшли ви до Мене.
MATT|25|37|Тоді відповідять Йому праведні й скажуть: Господи, коли то Тебе ми голодного бачили і нагодували, або спрагненого і напоїли?
MATT|25|38|Коли то Тебе мандрівником ми бачили і прийняли, чи нагим і зодягли?
MATT|25|39|Коли то Тебе ми недужого бачили, чи в в'язниці і до Тебе прийшли?
MATT|25|40|Цар відповість і промовить до них: Поправді кажу вам: що тільки вчинили ви одному з найменших братів Моїх цих, те Мені ви вчинили.
MATT|25|41|Тоді скаже й тим, хто ліворуч: Ідіть ви від Мене, прокляті, у вічний огонь, що дияволові та його посланцям приготований.
MATT|25|42|Бо Я голодував був і не нагодували Мене, прагнув і ви не напоїли Мене,
MATT|25|43|мандрівником Я був і не прийняли ви Мене, був нагий і не зодягли ви Мене, слабий і в в'язниці і Мене не відвідали ви.
MATT|25|44|Тоді відповідять і вони, промовляючи: Господи, коли то Тебе ми голодного бачили, або спрагненого, або мандрівником, чи нагого, чи недужого, чи в в'язниці і не послужили Тобі?
MATT|25|45|Тоді Він відповість їм і скаже: Поправді кажу вам: чого тільки одному з найменших цих ви не вчинили, Мені не вчинили!
MATT|25|46|І ці підуть на вічную муку, а праведники на вічне життя.
MATT|26|1|І сталось, коли закінчив Ісус усі ці слова, Він сказав Своїм учням:
MATT|26|2|Ви знаєте, що через два дні буде Пасха, і Людський Син буде виданий на розп'яття.
MATT|26|3|Тоді первосвященики, і книжники, і старші народу зібралися в домі первосвященика, званого Кайяфою,
MATT|26|4|і радилися, щоб підступом взяти Ісуса й забити.
MATT|26|5|І вони говорили: Та не в свято, щоб бува колотнеча в народі не сталась.
MATT|26|6|Коли ж Ісус був у Віфанії, у домі Симона прокаженого,
MATT|26|7|підійшла одна жінка до Нього, маючи алябастрову пляшечку дорогоцінного мира, і вилила на Його голову, як сидів при столі Він.
MATT|26|8|Як побачили ж учні це, то обурилися та й сказали: Нащо таке марнотратство?
MATT|26|9|Бо дорого можна було б це продати, і віддати убогим.
MATT|26|10|Зрозумівши Ісус, промовив до них: Чого прикрість ви робите жінці? Вона ж добрий учинок зробила Мені.
MATT|26|11|Бо вбогих ви маєте завжди з собою, а Мене не постійно ви маєте.
MATT|26|12|Бо, виливши миро оце на тіло Моє, вона те вчинила на похорон Мій.
MATT|26|13|Поправді кажу вам: де тільки оця Євангелія проповідувана буде в цілому світі, на пам'ятку їй буде сказане й те, що зробила вона!
MATT|26|14|Тоді один із Дванадцятьох, званий Юдою Іскаріотським, подався до первосвящеників,
MATT|26|15|і сказав: Що хочете дати мені, і я вам Його видам? І вони йому виплатили тридцять срібняків.
MATT|26|16|І він відтоді шукав слушного часу, щоб видати Його.
MATT|26|17|А першого дня Опрісноків учні підійшли до Ісуса й сказали Йому: Де хочеш, щоб ми приготували пасху спожити Тобі?
MATT|26|18|А Він відказав: Ідіть до такого то в місто, і перекажіть йому: каже Вчитель: час Мій близький, справлю Пасху з Своїми учнями в тебе.
MATT|26|19|І учні зробили, як звелів їм Ісус, і зачали пасху готувати.
MATT|26|20|А коли настав вечір, Він із дванадцятьма учнями сів за стіл.
MATT|26|21|І, як вони споживали, Він сказав: Поправді кажу вам, що один із вас видасть Мене...
MATT|26|22|А вони засмутилися тяжко, і кожен із них став питати Його: Чи не я то, о Господи?
MATT|26|23|А Він відповів і промовив: Хто руку свою вмочить у миску зо Мною, той видасть Мене.
MATT|26|24|Людський Син справді йде, як про Нього написано; але горе тому чоловікові, що видасть Людського Сина! Було б краще йому, коли б той чоловік не родився!
MATT|26|25|Юда ж, зрадник Його, відповів і сказав: Чи не я то, Учителю? Відказав Він йому: Ти сказав...
MATT|26|26|Як вони ж споживали, Ісус узяв хліб, і поблагословив, поламав, і давав Своїм учням, і сказав: Прийміть, споживайте, це тіло Моє.
MATT|26|27|А взявши чашу, і подяку вчинивши, Він подав їм і сказав: Пийте з неї всі,
MATT|26|28|бо це кров Моя Нового Заповіту, що за багатьох проливається на відпущення гріхів!
MATT|26|29|Кажу ж вам, що віднині не питиму Я від оцього плоду виноградного аж до дня, коли з вами його новим питиму в Царстві Мого Отця.
MATT|26|30|А коли відспівали вони, то на гору Оливну пішли.
MATT|26|31|Промовляє тоді їм Ісус: Усі ви через Мене спокуситеся ночі цієї. Бо написано: Уражу пастиря, і розпорошаться вівці отари.
MATT|26|32|По воскресенні ж Своїм Я вас випереджу в Галілеї.
MATT|26|33|А Петро відповів і сказав Йому: Якби й усі спокусились про Тебе, я не спокушуся ніколи.
MATT|26|34|Промовив до нього Ісус: Поправді кажу тобі, що ночі цієї, перше ніж заспіває півень, відречешся ти тричі від Мене...
MATT|26|35|Говорить до Нього Петро: Коли б мені навіть умерти з Тобою, я не відречуся від Тебе! Так сказали й усі учні.
MATT|26|36|Тоді з ними приходить Ісус до місцевости, званої Гефсиманія, і промовляє до учнів: Посидьте ви тут, аж поки піду й помолюся отам.
MATT|26|37|І, взявши Петра й двох синів Зеведеєвих, зачав сумувати й тужити.
MATT|26|38|Тоді промовляє до них: Обгорнена сумом смертельним душа Моя! Залишіться тут, і попильнуйте зо Мною...
MATT|26|39|І, трохи далі пройшовши, упав Він долілиць, та молився й благав: Отче Мій, коли можна, нехай обмине ця чаша Мене... Та проте, не як Я хочу, а як Ти...
MATT|26|40|І, вернувшись до учнів, знайшов їх, що спали, і промовив Петрові: Отак, не змогли ви й однієї години попильнувати зо Мною?...
MATT|26|41|Пильнуйте й моліться, щоб не впасти на спробу, бадьорий бо дух, але немічне тіло.
MATT|26|42|Відійшовши ще вдруге, Він молився й благав: Отче Мій, як ця чаша не може минути Мене, щоб не пити її, нехай станеться воля Твоя!
MATT|26|43|І, прийшовши, ізнову знайшов їх, що спали, бо зважніли їм очі були.
MATT|26|44|І, залишивши їх, знов пішов, і помолився втретє, те саме слово промовивши.
MATT|26|45|Потому приходить до учнів і їм промовляє: Ви ще далі спите й спочиваєте? Ось година наблизилась, і до рук грішникам виданий буде Син Людський...
MATT|26|46|Уставайте, ходім, ось наблизився Мій зрадник!
MATT|26|47|І коли Він іще говорив, аж ось прийшов Юда, один із Дванадцятьох, а з ним люду багато від первосвящеників і старших народу з мечами та киями.
MATT|26|48|А зрадник Його дав був знака їм, кажучи: Кого поцілую, то Він, беріть Його.
MATT|26|49|І зараз Він підійшов до Ісуса й сказав: Радій, Учителю! І поцілував Його.
MATT|26|50|Ісус же йому відказав: Чого, друже, прийшов ти? Тоді приступили та руки наклали на Ісуса, і схопили Його.
MATT|26|51|А ось один із тих, що з Ісусом були, витягнув руку, і меча свого вихопив та й рубонув раба первосвященика, і відтяв йому вухо.
MATT|26|52|Тоді промовляє до нього Ісус: Сховай свого меча в його місце, бо всі, хто візьме меча, від меча і загинуть.
MATT|26|53|Чи ти думаєш, що не можу тепер упросити Свого Отця, і Він дасть Мені зараз більше дванадцяти леґіонів Анголів?
MATT|26|54|Але як має збутись Писання, що так статися мусить?
MATT|26|55|Тієї години промовив Ісус до народу: Немов на розбійника вийшли з мечами та киями, щоб узяти Мене! Я щоденно у храмі сидів і навчав, і Мене не взяли ви.
MATT|26|56|Це ж сталось усе, щоб збулися писання пророків. Усі учні тоді залишили Його й повтікали...
MATT|26|57|А вони схопили Ісуса, і повели до первосвященика Кайяфи, де зібралися книжники й старші.
MATT|26|58|Петро ж здалека йшов услід за Ним аж до двору первосвященика, і, ввійшовши всередину, сів із службою, щоб бачити кінець.
MATT|26|59|А первосвященики та ввесь синедріон шукали на Ісуса неправдивого свідчення, щоб смерть заподіяти Йому,
MATT|26|60|і не знаходили, хоч кривосвідків багато підходило. Аж ось накінець з'явилися двоє,
MATT|26|61|і сказали: Він говорив: Я можу зруйнувати храм Божий, і за три дні збудувати його.
MATT|26|62|Тоді первосвященик устав і до Нього сказав: Ти нічого не відповідаєш на те, що свідчать супроти Тебе?
MATT|26|63|Ісус же мовчав. І первосвященик сказав Йому: Заприсягаю Тебе Живим Богом, щоб нам Ти сказав, чи Христос Ти, Син Божий?
MATT|26|64|Промовляє до нього Ісус: Ти сказав... А навіть повім вам: відтепер ви побачите Людського Сина, що сидітиме праворуч сили Божої, і на хмарах небесних приходитиме!
MATT|26|65|Тоді первосвященик роздер одежу свою та й сказав: Він богозневажив! Нащо нам іще свідки потрібні? Ось ви чули тепер Його богозневагу!
MATT|26|66|Як вам іздається? Вони ж відповіли та сказали: Повинен умерти!
MATT|26|67|Тоді стали плювати на обличчя Йому, та бити по щоках Його, інші ж киями били,
MATT|26|68|і казали: Пророкуй нам, Христе, хто то вдарив Тебе?...
MATT|26|69|А Петро перед домом сидів на подвір'ї. І приступила до нього служниця одна та й сказала: І ти був з Ісусом Галілеянином!
MATT|26|70|А він перед всіма відрікся, сказавши: Не відаю я, що ти кажеш...
MATT|26|71|А коли до воріт він підходив, побачила інша його та й сказала приявним там людям: Оцей був з Ісусом Назарянином!
MATT|26|72|І він знову відрікся та став присягатись: Не знаю Цього Чоловіка!...
MATT|26|73|Підійшли ж трохи згодом присутні й сказали Петрові: І ти справді з отих, та й мова твоя виявляє тебе.
MATT|26|74|Тоді він став клястись та божитись: Не знаю Цього Чоловіка! І заспівав півень хвилі тієї...
MATT|26|75|І згадав Петро сказане слово Ісусове: Перше ніж заспіває півень, відречешся ти тричі від Мене. І, вийшовши звідти, він гірко заплакав...
MATT|27|1|А коли настав ранок, усі первосвященики й старші народу зібрали нараду супроти Ісуса, щоб Йому заподіяти смерть.
MATT|27|2|І, зв'язавши Його, повели, та й Понтію Пилату намісникові віддали.
MATT|27|3|Тоді Юда, що видав Його, як побачив, що Його засудили, розкаявся, і вернув тридцять срібняків первосвященикам і старшим,
MATT|27|4|та й сказав: Я згрішив, невинну кров видавши. Вони ж відказали: А нам що до того? Дивись собі сам...
MATT|27|5|І, кинувши в храм срібняки, відійшов, а потому пішов, та й повісився...
MATT|27|6|А первосвященики, як взяли срібняки, то сказали: Цього не годиться покласти до сховку церковного, це ж бо заплата за кров.
MATT|27|7|А порадившись, купили на них поле ганчарське, щоб мандрівників ховати,
MATT|27|8|чому й зветься те поле полем крови аж до сьогодні.
MATT|27|9|Тоді справдилось те, що сказав був пророк Єремія, промовляючи: І взяли вони тридцять срібняків, заплату Оціненого, що Його оцінили сини Ізраїлеві,
MATT|27|10|і дали їх за поле ганчарське, як Господь наказав був мені.
MATT|27|11|Ісус же став перед намісником. І намісник Його запитав і сказав: Чи Ти Цар Юдейський? Ісус же йому відказав: Ти кажеш.
MATT|27|12|Коли ж первосвященики й старші Його винуватили, Він нічого на те не відказував.
MATT|27|13|Тоді каже до Нього Пилат: Чи не чуєш, як багато на Тебе свідкують?
MATT|27|14|А Він ні на одне слово йому не відказував, так що намісник був дуже здивований.
MATT|27|15|Мав же намісник звичай відпускати на свято народові в'язня одного, котрого хотіли вони.
MATT|27|16|Був тоді в'язень відомий, що звався Варавва.
MATT|27|17|І, як зібрались вони, то сказав їм Пилат: Котрого бажаєте, щоб я вам відпустив: Варавву, чи Ісуса, що зветься Христос?
MATT|27|18|Бо він знав, що Його через заздрощі видали.
MATT|27|19|Коли ж він сидів на суддевім сидінні, його дружина прислала сказати йому: Нічого не май з отим Праведником, бо сьогодні вві сні я багато терпіла з-за Нього...
MATT|27|20|А первосвященики й старші попідмовляли народ, щоб просити за Варавву, а Ісусові смерть заподіяти.
MATT|27|21|Намісник тоді відповів і сказав їм: Котрого ж із двох ви бажаєте, щоб я вам відпустив? Вони ж відказали: Варавву.
MATT|27|22|Пилат каже до них: А що ж маю зробити з Ісусом, що зветься Христос? Усі закричали: Нехай розп'ятий буде!...
MATT|27|23|А намісник спитав: Яке ж зло Він зробив? Вони ж зачали ще сильніше кричати й казати: Нехай розп'ятий буде!
MATT|27|24|І, як побачив Пилат, що нічого не вдіє, а неспокій ще більший стається, набрав він води, та й перед народом умив свої руки й сказав: Я невинний у крові Його! Самі ви побачите...
MATT|27|25|А ввесь народ відповів і сказав: На нас Його кров і на наших дітей!...
MATT|27|26|Тоді відпустив їм Варавву, а Ісуса, збичувавши, він видав, щоб розп'ятий був.
MATT|27|27|Тоді то намісникові вояки, до преторія взявши Ісуса, зібрали на Нього ввесь відділ.
MATT|27|28|І, роздягнувши Його, багряницю наділи на Нього.
MATT|27|29|І, сплівши з тернини вінка, поклали Йому на голову, а тростину в правицю Його. І, навколішки падаючи перед Ним, сміялися з Нього й казали: Радій, Царю Юдейський!
MATT|27|30|І, плювавши на Нього, хапали тростину, та й по голові Його били...
MATT|27|31|А коли назнущалися з Нього, зняли з Нього плаща, і зодягнули в одежу Його. І повели Його на розп'яття.
MATT|27|32|А виходячи, стріли одного кірінеянина, Симон на ймення, його змусили нести для Нього хреста.
MATT|27|33|І, прибувши на місце, що зветься Голгофа, цебто сказати Череповище,
MATT|27|34|дали Йому пити вина, із гіркотою змішаного, та, покуштувавши, Він пити не схотів.
MATT|27|35|А розп'явши Його, вони поділили одежу Його, кинувши жереба.
MATT|27|36|І, посідавши, стерегли Його там.
MATT|27|37|І напис провини Його помістили над Його головою: Це Ісус, Цар Юдейський.
MATT|27|38|Тоді розп'ято з Ним двох розбійників: одного праворуч, а одного ліворуч.
MATT|27|39|А хто побіч проходив, Його лихословили та головами своїми хитали,
MATT|27|40|і казали: Ти, що храма руйнуєш та за три дні будуєш, спаси Самого Себе! Коли Ти Божий Син, то зійди з хреста!
MATT|27|41|Так само ж і первосвященики з книжниками та старшими, насміхаючися, говорили:
MATT|27|42|Він інших спасав, а Самого Себе не може спасти! Коли Цар Він Ізраїлів, нехай зійде тепер із хреста, і ми повіримо Йому!
MATT|27|43|Покладав Він надію на Бога, нехай Той Його тепер визволить, якщо Він угодний Йому. Бо Він говорив: Я Син Божий...
MATT|27|44|Також насміхалися з Нього й розбійники, що з Ним були розп'яті.
MATT|27|45|А від години шостої аж до години дев'ятої темрява сталась по цілій землі!
MATT|27|46|А коло години дев'ятої скрикнув Ісус гучним голосом, кажучи: Елі, Елі, лама савахтані? цебто: Боже Мій, Боже Мій, нащо Мене Ти покинув?...
MATT|27|47|Дехто ж із тих, що стояли там, це почули й казали, що Він кличе Іллю.
MATT|27|48|А один із них зараз побіг і взяв губку та, оцтом її наповнивши, настромив на тростину й давав Йому пити.
MATT|27|49|Інші казали: Чекай но, побачмо, чи прийде Ілля визволяти Його.
MATT|27|50|А Ісус знову голосом гучним іскрикнув, і духа віддав...
MATT|27|51|І ось завіса у храмі роздерлась надвоє від верху аж додолу, і земля потряслася, і зачали розпадатися скелі,
MATT|27|52|і повідкривались гроби, і повставало багато тіл спочилих святих,
MATT|27|53|а з гробів повиходивши, по Його воскресенні, до міста святого ввійшли, і багатьом із'явились.
MATT|27|54|А сотник та ті, що Ісуса з ним стерегли, як землетруса побачили, і те, що там сталося, налякалися дуже й казали: Він був справді Син Божий!
MATT|27|55|Було там багато й жінок, що дивилися здалека, і що за Ісусом прийшли з Галілеї, і Йому прислуговували.
MATT|27|56|Між ними була Марія Магдалина, і Марія, мати Якова й Йосипа, і мати синів Зеведеєвих.
MATT|27|57|А коли настав вечір, то прийшов муж багатий із Ариматеї, на ім'я Йосип, що й сам був навчався в Ісуса.
MATT|27|58|Він прийшов до Пилата й просив тіла Ісусового. Пилат ізвелів тоді видати.
MATT|27|59|І взяв Йосип Ісусове тіло, обгорнув його плащаницею чистою,
MATT|27|60|і поклав його в гробі новому своїм, що був висік у скелі. До дверей гробових привалив він великого каменя, та й відійшов.
MATT|27|61|Була ж там Марія Магдалина та інша Марія, що сиділи насупроти гробу.
MATT|27|62|А наступного дня, що за п'ятницею, до Пилата зібралися первосвященики та фарисеї,
MATT|27|63|і сказали: Пригадали ми, пане, собі, що обманець отой, як живий іще був, то сказав: По трьох днях Я воскресну.
MATT|27|64|Звели ж гріб стерегти аж до третього дня, щоб учні Його не прийшли, та й не вкрали Його, і не сказали народові: Він із мертвих воскрес! І буде остання обмана гірша за першу...
MATT|27|65|Відказав їм Пилат: Сторожу ви маєте, ідіть, забезпечте, як знаєте.
MATT|27|66|І вони відійшли, і, запечатавши каменя, біля гробу сторожу поставили.
MATT|28|1|Як минула ж субота, на світанку дня першого в тижні, прийшла Марія Магдалина та інша Марія побачити гріб.
MATT|28|2|І великий ось ставсь землетрус, бо зійшов із неба Ангол Господній, і, приступивши, відвалив від гробу каменя, та й сів на ньому.
MATT|28|3|Його ж постать була, як та блискавка, а шати його були білі, як сніг.
MATT|28|4|І від страху перед ним затряслася сторожа, та й стала, як мертва.
MATT|28|5|А Ангол озвався й промовив жінкам: Не лякайтеся, бо я знаю, що Ісуса розп'ятого це ви шукаєте.
MATT|28|6|Нема Його тут, бо воскрес, як сказав. Підійдіть, подивіться на місце, де знаходився Він.
MATT|28|7|Ідіть же хутко, і скажіть Його учням, що воскрес Він із мертвих, і ото випереджує вас в Галілеї, там Його ви побачите. Ось, вам я звістив!
MATT|28|8|І пішли вони хутко від гробу, зо страхом і великою радістю, і побігли, щоб учнів Його сповістити.
MATT|28|9|Аж ось перестрів їх Ісус і сказав: Радійте! Вони ж підійшли, обняли Його ноги і вклонились Йому до землі.
MATT|28|10|Промовляє тоді їм Ісус: Не лякайтесь! Ідіть, повідомте братів Моїх, нехай вони йдуть у Галілею, там побачать Мене!
MATT|28|11|Коли ж вони йшли, ось дехто зо сторожі до міста прийшли та й первосвященикам розповіли все, що сталось.
MATT|28|12|І, зібравшись зо старшими, вони врадили раду, і дали сторожі чимало срібняків,
MATT|28|13|і сказали: Розповідайте: Його учні вночі прибули, і вкрали Його, як ми спали.
MATT|28|14|Як почує ж намісник про це, то його ми переконаємо, і від клопоту визволимо вас.
MATT|28|15|І, взявши вони срібняки, зробили, як навчено їх. І пронеслося слово оце між юдеями, і тримається аж до сьогодні.
MATT|28|16|Одинадцять же учнів пішли в Галілею на гору, куди звелів їм Ісус.
MATT|28|17|І як вони Його вгледіли, поклонились Йому до землі, а дехто вагався.
MATT|28|18|А Ісус підійшов і промовив до них та й сказав: Дана Мені всяка влада на небі й на землі.
MATT|28|19|Тож ідіть, і навчіть всі народи, христячи їх в Ім'я Отця, і Сина, і Святого Духа,
MATT|28|20|навчаючи їх зберігати все те, що Я вам заповів. І ото, Я перебуватиму з вами повсякденно аж до кінця віку! Амінь
