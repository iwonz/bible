NEH|1|1|Слова Неемии, сына Ахалиина. В месяце Кислеве, в двадцатом году, я находился в Сузах, престольном городе.
NEH|1|2|И пришел Ханани, один из братьев моих, он и [несколько] человек из Иудеи. И спросил я их об уцелевших Иудеях, которые остались от плена, и об Иерусалиме.
NEH|1|3|И сказали они мне: оставшиеся, которые остались от плена, [находятся] там, в стране [своей], в великом бедствии и в уничижении; и стена Иерусалима разрушена, и ворота его сожжены огнем.
NEH|1|4|Услышав эти слова, я сел и заплакал, и печален был несколько дней, и постился и молился пред Богом небесным
NEH|1|5|и говорил: Господи Боже небес, Боже великий и страшный, хранящий завет и милость к любящим Тебя и соблюдающим заповеди Твои!
NEH|1|6|Да будут уши Твои внимательны и очи Твои отверсты, чтобы услышать молитву раба Твоего, которою я теперь день и ночь молюсь пред Тобою о сынах Израилевых, рабах Твоих, и исповедуюсь во грехах сынов Израилевых, которыми согрешили мы пред Тобою, согрешили – и я и дом отца моего.
NEH|1|7|Мы стали преступны пред Тобою и не сохранили заповедей и уставов и определений, которые Ты заповедал Моисею, рабу Твоему.
NEH|1|8|Но помяни слово, которое Ты заповедал Моисею, рабу Твоему, говоря: [если] вы сделаетесь преступниками, то Я рассею вас по народам;
NEH|1|9|[когда] же обратитесь ко Мне и будете хранить заповеди Мои и исполнять их, то хотя бы вы изгнаны были на край неба, и оттуда соберу вас и приведу вас на место, которое избрал Я, чтобы водворить там имя Мое.
NEH|1|10|Они же рабы Твои и народ Твой, который Ты искупил силою Твоею великою и рукою Твоею могущественною.
NEH|1|11|Молю Тебя, Господи! Да будет ухо Твое внимательно к молитве раба Твоего и к молитве рабов Твоих, любящих благоговеть пред именем Твоим. И благопоспеши рабу Твоему теперь, и введи его в милость у человека сего. Я был виночерпием у царя.
NEH|2|1|В месяце Нисане, в двадцатый год царя Артаксеркса, [было] перед ним вино. И я взял вино и подал царю, и, казалось, не был печален перед ним.
NEH|2|2|Но царь сказал мне: отчего лице у тебя печально; ты не болен, этого нет, а верно печаль на сердце? Я сильно испугался
NEH|2|3|и сказал царю: да живет царь во веки! Как не быть печальным лицу моему, когда город, дом гробов отцов моих, в запустении, и ворота его сожжены огнем!
NEH|2|4|И сказал мне царь: чего же ты желаешь? Я помолился Богу небесному
NEH|2|5|и сказал царю: если царю благоугодно, и если в благоволении раб твой пред лицем твоим, то пошли меня в Иудею, в город, [где] гробы отцов моих, чтоб я обстроил его.
NEH|2|6|И сказал мне царь и царица, которая сидела подле него: сколько времени продлится путь твой, и когда возвратишься? И благоугодно было царю послать меня, после того как я назначил время.
NEH|2|7|И сказал я царю: если царю благоугодно, то дал бы мне письма к заречным областеначальникам, чтоб они давали мне пропуск, доколе я не дойду до Иудеи,
NEH|2|8|и письмо к Асафу, хранителю царских лесов, чтоб он дал мне дерев для ворот крепости, которая при доме [Божием], и для городской стены, и для дома, в котором бы мне жить. И дал мне царь, так как благодеющая рука Бога моего была надо мною.
NEH|2|9|И пришел я к заречным областеначальникам и отдал им царские письма. Послал же со мною царь воинских начальников со всадниками.
NEH|2|10|Когда услышал [сие] Санаваллат, Хоронит и Товия, Аммонитский раб, то им было весьма досадно, что пришел человек заботиться о благе сынов Израилевых.
NEH|2|11|И пришел я в Иерусалим. И пробыв там три дня,
NEH|2|12|встал я ночью с немногими людьми, [бывшими] при мне, и никому не сказал, что Бог мой положил мне на сердце сделать для Иерусалима; животного же не было со мною никакого, кроме того, на котором я ехал.
NEH|2|13|И проехал я ночью через ворота Долины перед источником Драконовым к воротам Навозным, и осмотрел я стены Иерусалима разрушенные и его ворота, сожженные огнем.
NEH|2|14|И подъехал я к воротам Источника и к царскому водоему, но [там] не было места пройти животному, которое было подо мною, –
NEH|2|15|и я поднялся назад по лощине ночью и осматривал стену, и проехав [опять] воротами Долины, возвратился.
NEH|2|16|И начальствующие не знали, куда я ходил и что я делаю: ни Иудеям, ни священникам, ни знатнейшим, ни начальствующим, ни прочим производителям работ я дотоле ничего не открывал.
NEH|2|17|И сказал я им: вы видите бедствие, в каком мы находимся; Иерусалим пуст и ворота его сожжены огнем; пойдем, построим стену Иерусалима, и не будем впредь [в таком] уничижении.
NEH|2|18|И я рассказал им о благодеявшей мне руке Бога моего, а также и слова царя, которые он говорил мне. И сказали они: будем строить, – и укрепили руки свои на благое [дело].
NEH|2|19|Услышав это, Санаваллат, Хоронит и Товия, Аммонитский раб, и Гешем Аравитянин смеялись над нами и с презрением говорили: что это за дело, которое вы делаете? уже не думаете ли возмутиться против царя?
NEH|2|20|Я дал им ответ и сказал им: Бог Небесный, Он благопоспешит нам, и мы, рабы Его, станем строить, а вам нет части и права и памяти в Иерусалиме.
NEH|3|1|И встал Елияшив, великий священник, и братья его священники и построили Овечьи ворота: они освятили их и вставили двери их, и от башни Меа освятили их до башни Хананела.
NEH|3|2|И подле него строили Иерихонцы, а подле них строил Закхур, сын Имрия.
NEH|3|3|Ворота Рыбные строили уроженцы Сенаи: они покрыли их, и вставили двери их, замки их и засовы их.
NEH|3|4|Подле них чинил [стену] Меремоф, сын Урии, сын Гаккоца; подле них чинил Мешуллам, сын Берехии, сын Мешизабела; подле них чинил Садок, сын Бааны;
NEH|3|5|подле них чинили Фекойцы; впрочем знатнейшие из них не наклонили шеи своей поработать для Господа своего.
NEH|3|6|Старые ворота чинили Иоиада, сын Пасеаха, и Мешуллам, сын Бесодии: они покрыли их и вставили двери их, и замки их и засовы их.
NEH|3|7|Подле них чинил Мелатия Гаваонитянин, и Иадон из Меронофа, с жителями Гаваона и Мицфы, подвластными заречному областеначальнику.
NEH|3|8|Подле него чинил Уззиил, сын Харгаии, серебряник, а подле него чинил Ханания, сын Гараккахима. И восстановили Иерусалим до стены широкой.
NEH|3|9|Подле них чинил Рефаия, сын Хура, начальник полуокруга Иерусалимского.
NEH|3|10|Подле них и против дома своего чинил Иедаия, сын Харумафа, а подле него чинил Хаттуш, сын Хашавнии.
NEH|3|11|На втором участке чинил Малхия, сын Харима, и Хашшув, сын Пахаф–Моава; [они же чинили] и башню Печную.
NEH|3|12|Подле них чинил Шаллум, сын Галлохеша, начальник полуокруга Иерусалимского, он и дочери его.
NEH|3|13|Ворота Долины чинил Ханун и жители Заноаха: они построили их, и вставили двери их, замки их и засовы их, и [еще чинили] они тысячу локтей стены до ворот Навозных.
NEH|3|14|А ворота Навозные чинил Малхия, сын Рехава, начальник Бефкаремского округа: он построил их и вставил двери их, замки их и засовы их.
NEH|3|15|Ворота Источника чинил Шаллум, сын Колхозея, начальник округа Мицфы: он построил их, и покрыл их, и вставил двери их, замки их и засовы их, – [он же чинил] стену у водоема Селах против царского сада и до ступеней, спускающихся из города Давидова.
NEH|3|16|За ним чинил Неемия, сын Азбука, начальник полуокруга Бефцурского, до гробниц Давидовых и до выкопанного пруда и до дома храбрых.
NEH|3|17|За ним чинили левиты: Рехум, сын Вания; подле него чинил Хашавия, начальник полуокруга Кеильского, за свой округ.
NEH|3|18|За ним чинили братья их: Баввай, сын Хенадада, начальник Кеильского полуокруга.
NEH|3|19|А подле него чинил Езер, сын Иисуса, начальник Мицфы, на втором участке, напротив всхода к оружейне на углу.
NEH|3|20|За ним ревностно чинил Варух, сын Забвая, на втором участке, от угла до дверей дома Елияшива, великого священника.
NEH|3|21|За ним чинил Меремоф, сын Урии, сын Гаккоца, на втором участке, от дверей дома Елияшивова до конца дома Елияшивова.
NEH|3|22|За ним чинили священники из окрестностей.
NEH|3|23|За ними чинил Вениамин и Хашшув, против дома своего; за ними чинил Азария, сын Маасеи, сын Анании, возле дома своего.
NEH|3|24|За ним чинил Биннуй, сын Хенадада, на втором участке, от дома Азарии до угла и поворота.
NEH|3|25|[За ним] Фалал, сын Узая, напротив угла и башни, выступающей от верхнего дома царского, которая у двора темничного. За ним Федаия, сын Пароша.
NEH|3|26|Нефинеи же, [которые] жили в Офеле, [починили] напротив Водяных ворот к востоку и до выступающей башни.
NEH|3|27|За ними чинили Фекойцы, на втором участке, от [места] напротив большой выступающей башни до стены Офела.
NEH|3|28|Далее ворот Конских чинили священники, каждый против своего дома.
NEH|3|29|За ними чинил Садок, сын Иммера, против своего дома, а за ним чинил Шемаия, сын Шехании, сторож восточных ворот.
NEH|3|30|За ним чинил Ханания, сын Шелемии, и Ханун, шестой сын Цалафа, на втором участке. За ним чинил Мешуллам, сын Берехии, против комнаты своей.
NEH|3|31|За ним чинил Малхия, сын Гацорфия, до дома нефинеев и торговцев, против ворот Гаммифкад и до угольного жилья.
NEH|3|32|А между угольным жильем до ворот Овечьих чинили серебряники и торговцы.
NEH|3|33|Когда услышал Санаваллат, что мы строим стену, он рассердился и много досадовал и издевался над Иудеями;
NEH|3|34|и говорил при братьях своих и при Самарийских военных людях, и сказал: что делают эти жалкие Иудеи? неужели им это дозволят? неужели будут они приносить жертвы? неужели они когда–либо кончат? неужели они оживят камни из груд праха, и притом пожженные?
NEH|3|35|А Товия Аммонитянин, [бывший] подле него, сказал: пусть их строят; пойдет лисица, и разрушит их каменную стену.
NEH|3|36|Услыши, Боже наш, в каком мы презрении, и обрати ругательство их на их голову, и предай их презрению в земле пленения;
NEH|3|37|и не покрой беззаконий их, и грех их да не изгладится пред лицем Твоим, потому что они огорчили строящих!
NEH|3|38|Мы однако же строили стену, и сложена была вся стена до половины ее. И у народа доставало усердия работать.
NEH|4|1|Когда услышал Санаваллат и Товия, и Аравитяне, и Аммонитяне, и Азотяне, что стены Иерусалимские восстановляются, что повреждения начали заделываться, то им было весьма досадно.
NEH|4|2|И сговорились все вместе пойти войною на Иерусалим и разрушить его.
NEH|4|3|И мы молились Богу нашему, и ставили против них стражу днем и ночью, для спасения от них.
NEH|4|4|Но Иудеи сказали: ослабела сила у носильщиков, а мусору много; мы не в состоянии строить стену.
NEH|4|5|А неприятели наши говорили: не узнают и не увидят, как [вдруг] мы войдем в средину их и перебьем их, и остановим дело.
NEH|4|6|Когда приходили Иудеи, жившие подле них, и говорили нам раз десять, со всех мест, что они нападут на нас:
NEH|4|7|тогда в низменных местах у города, за стеною, на местах сухих поставил я народ по–племенно с мечами их, с копьями их и луками их.
NEH|4|8|И осмотрел я, и стал, и сказал знатнейшим и начальствующим и прочему народу: не бойтесь их; помните Господа великого и страшного и сражайтесь за братьев своих, за сыновей своих и за дочерей своих, за жен своих и за домы свои.
NEH|4|9|Когда услышали неприятели наши, что нам известно [намерение] [их], тогда разорил Бог замысел их, и все мы возвратились к стене, каждый на свою работу.
NEH|4|10|С того дня половина молодых людей у меня занималась работою, а [другая] половина их держала копья, щиты и луки и латы; и начальствующие [находились] позади всего дома Иудина.
NEH|4|11|Строившие стену и носившие тяжести, которые налагали [на них], одною рукою производили работу, а другою держали копье.
NEH|4|12|Каждый из строивших препоясан был мечом по чреслам своим, и [так] они строили. Возле меня находился трубач.
NEH|4|13|И сказал я знатнейшим и начальствующим и прочему народу: работа велика и обширна, и мы рассеяны по стене и отдалены друг от друга;
NEH|4|14|поэтому, откуда услышите вы звук трубы, в то место собирайтесь к нам: Бог наш будет сражаться за нас.
NEH|4|15|Так производили мы работу; и половина держала копья от восхода зари до появления звезд.
NEH|4|16|Сверх сего, в то же время я сказал народу, чтобы в Иерусалиме ночевали все с рабами своими, – и будут они у нас ночью на страже, а днем на работе.
NEH|4|17|И ни я, ни братья мои, ни слуги мои, ни стражи, сопровождавшие меня, не снимали с себя одеяния своего, у каждого были под рукою меч и вода.
NEH|5|1|И сделался большой ропот в народе и у жен его на братьев своих Иудеев.
NEH|5|2|Были такие, которые говорили: нас, сыновей наших и дочерей наших много; и мы желали бы доставать хлеб и кормиться и жить.
NEH|5|3|Были и такие, которые говорили: поля свои, и виноградники свои, и домы свои мы закладываем, чтобы достать хлеба от голода.
NEH|5|4|Были и такие, которые говорили: мы занимаем серебро на подать царю [под залог] полей наших и виноградников наших;
NEH|5|5|у нас такие же тела, какие тела у братьев наших, и сыновья наши такие же, как их сыновья; а вот, мы должны отдавать сыновей наших и дочерей наших в рабы, и некоторые из дочерей наших уже находятся в порабощении. Нет никаких средств для выкупа в руках наших; и поля наши и виноградники наши у других.
NEH|5|6|Когда я услышал ропот их и такие слова, я очень рассердился.
NEH|5|7|Сердце мое возмутилось, и я строго выговорил знатнейшим и начальствующим и сказал им: вы берете лихву с братьев своих. И созвал я против них большое собрание
NEH|5|8|и сказал им: мы выкупали братьев своих, Иудеев, проданных народам, сколько было сил у нас, а вы продаете братьев своих, и они продаются нам? Они молчали и не находили ответа.
NEH|5|9|И сказал я: нехорошо вы делаете. Не в страхе ли Бога нашего должны ходить вы, дабы избегнуть поношения от народов, врагов наших?
NEH|5|10|И я также, братья мои и [служащие] при мне давали им в заем и серебро и хлеб: оставим им долг сей.
NEH|5|11|Возвратите им ныне же поля их, виноградные и масличные сады их, и домы их, и рост с серебра и хлеба, и вина и масла, за который вы ссудили их.
NEH|5|12|И сказали они: возвратим и не будем с них требовать; сделаем так, как ты говоришь. И позвал я священников и велел им дать клятву, что они так сделают.
NEH|5|13|И вытряхнул я [одежду] мою и сказал: так пусть вытряхнет Бог всякого человека, который не сдержит слова сего, из дома его и из имения его, и так да будет у него вытрясено и пусто! И сказало все собрание: аминь. И прославили Бога; и народ выполнил слово сие.
NEH|5|14|Еще: с того дня, как определен я был областеначальником их в земле Иудейской, от двадцатого года до тридцать второго года царя Артаксеркса, в продолжение двенадцати лет я и братья мои не ели хлеба областеначальнического.
NEH|5|15|А прежние областеначальники, которые [были] до меня, отягощали народ и брали с них хлеб и вино, кроме сорока сиклей серебра; даже и слуги их господствовали над народом. Я же не делал так по страху Божию.
NEH|5|16|При этом работы на стене сей я поддерживал; и полей мы не закупали, и все слуги мои собирались туда на работу.
NEH|5|17|Иудеев и начальствующих по сто пятидесяти человек [бывало] за столом у меня, кроме приходивших к нам из окрестных народов.
NEH|5|18|И [вот] что было приготовляемо на один день: один бык, шесть отборных овец и птицы приготовлялись у меня; и в десять дней [издерживалось] множество всякого вина. И при [всем] том, хлеба областеначальнического я не требовал, так как тяжелая служба [лежала] на народе сем.
NEH|5|19|Помяни, Боже мой, во благо мне все, что я сделал для народа сего!
NEH|6|1|Когда дошло до слуха Санаваллата и Товии и Гешема Аравитянина и прочих неприятелей наших, что я отстроил стену, и не оставалось в ней повреждений – впрочем до того времени я еще не ставил дверей в ворота, –
NEH|6|2|тогда прислал Санаваллат и Гешем ко мне сказать: приди, и сойдемся в одном из сел на равнине Оно. Они замышляли сделать мне зло.
NEH|6|3|Но я послал к ним послов сказать: я занят большим делом, не могу сойти; дело остановилось бы, если бы я оставил его и сошел к вам.
NEH|6|4|Четыре раза присылали они ко мне с таким же приглашением, и я отвечал им то же.
NEH|6|5|Тогда прислал ко мне Санаваллат в пятый раз своего слугу, у которого в руке было открытое письмо.
NEH|6|6|В нем было написано: слух носится у народов, и Гешем говорит, будто ты и Иудеи задумали отпасть, для чего и строишь стену и хочешь быть у них царем, по тем же слухам;
NEH|6|7|и пророков поставил ты, чтоб они разглашали о тебе в Иерусалиме и говорили: царь Иудейский! И такие речи дойдут до царя. Итак приходи, и посоветуемся вместе.
NEH|6|8|Но я послал к нему сказать: ничего такого не было, о чем ты говоришь; ты выдумал это своим умом.
NEH|6|9|Ибо все они стращали нас, думая: опустятся руки их от дела сего, и оно не состоится; но я тем более укрепил руки мои.
NEH|6|10|Пришел я в дом Шемаии, сына Делаии, сына Мегетавелова, и он заперся и сказал: пойдем в дом Божий, внутрь храма, и запрем за собою двери храма, потому что придут убить тебя, и придут убить тебя ночью.
NEH|6|11|Но я сказал: может ли бежать такой человек, как я? Может ли такой, как я, войти в храм, чтобы остаться живым? Не пойду.
NEH|6|12|Я знал, что не Бог послал его, хотя он пророчески говорил мне, но что Товия и Санаваллат подкупили его.
NEH|6|13|Для того он был подкуплен, чтоб я устрашился и сделал так и согрешил, и чтобы имели о мне худое мнение и преследовали меня за это укоризнами.
NEH|6|14|Помяни, Боже мой, Товию и Санаваллата по сим делам их, а также пророчицу Ноадию и прочих пророков, которые хотели устрашить меня!
NEH|6|15|Стена была совершена в двадцать пятый день месяца Елула, в пятьдесят два дня.
NEH|6|16|Когда услышали об этом все неприятели наши, и увидели это все народы, которые вокруг нас, тогда они очень упали в глазах своих и познали, что это дело сделано Богом нашим.
NEH|6|17|Сверх того в те дни знатнейшие Иудеи много писали писем, которые посылались к Товии, а Товиины письма приходили к ним.
NEH|6|18|Ибо многие в Иудее были в клятвенном союзе с ним, потому что он был зять Шехании, сын Арахова, а сын его Иоханан взял [за себя] дочь Мешуллама, сына Верехии.
NEH|6|19|Даже о доброте его они говорили при мне, и мои слова переносились к нему. Товия присылал письма, чтоб устрашить меня.
NEH|7|1|Когда стена была построена, и я вставил двери, и поставлены были на свое служение привратники и певцы и левиты,
NEH|7|2|тогда приказал я брату моему Ханани и начальнику Иерусалимской крепости Хананию, ибо он более многих других был человек верный и богобоязненный,
NEH|7|3|и сказал я им: пусть не отворяют ворот Иерусалимских, доколе не обогреет солнце, и доколе они стоят, пусть замыкают и запирают двери. И поставил я стражами жителей Иерусалима, каждого на свою стражу и каждого напротив дома его.
NEH|7|4|Но город был пространен и велик, а народа в нем было немного, и домы не были построены.
NEH|7|5|И положил мне Бог мой на сердце собрать знатнейших и начальствующих и народ, чтобы сделать перепись. И нашел я родословную перепись тех, которые сначала пришли, и в ней написано:
NEH|7|6|вот жители страны, которые отправились из пленников, переселенных Навуходоносором, царем Вавилонским, и возвратились в Иерусалим и Иудею, каждый в свой город, –
NEH|7|7|те, которые пошли с Зоровавелем, Иисусом, Неемиею, Азариею, Раамиею, Нахманием, Мардохеем, Билшаном, Мисферефом, Бигваем, Нехумом, Вааною. Число людей народа Израилева:
NEH|7|8|сыновей Пароша две тысячи сто семьдесят два.
NEH|7|9|Сыновей Сафатии триста семьдесят два.
NEH|7|10|Сыновей Араха шестьсот пятьдесят два.
NEH|7|11|Сыновей Пахаф–Моава, из сыновей Иисуса и Иоава, две тысячи восемьсот восемнадцать.
NEH|7|12|Сыновей Елама тысяча двести пятьдесят четыре.
NEH|7|13|Сыновей Заффу восемьсот сорок пять.
NEH|7|14|Сыновей Закхая семьсот шестьдесят.
NEH|7|15|Сыновей Биннуя шестьсот сорок восемь.
NEH|7|16|Сыновей Бевая шестьсот двадцать восемь.
NEH|7|17|Сыновей Азгада две тысячи триста двадцать два.
NEH|7|18|Сыновей Адоникама шестьсот шестьдесят семь.
NEH|7|19|Сыновей Бигвая две тысячи шестьсот семь.
NEH|7|20|Сыновей Адина шестьсот пятьдесят пять.
NEH|7|21|Сыновей Атера из [дома] Езекии девяносто восемь.
NEH|7|22|Сыновей Хашума триста двадцать восемь.
NEH|7|23|Сыновей Вецая триста двадцать четыре.
NEH|7|24|Сыновей Харифа сто двенадцать.
NEH|7|25|Уроженцев Гаваона девяносто пять.
NEH|7|26|Жителей Вифлеема и Нетофы сто восемьдесят восемь.
NEH|7|27|Жителей Анафофа сто двадцать восемь.
NEH|7|28|Жителей Беф–Азмавефа сорок два.
NEH|7|29|Жителей Кириаф–Иарима, Кефиры и Беерофа семьсот сорок три.
NEH|7|30|Жителей Рамы и Гевы шестьсот двадцать один.
NEH|7|31|Жителей Михмаса сто двадцать два.
NEH|7|32|Жителей Вефиля и Гая сто двадцать три.
NEH|7|33|Жителей Нево другого пятьдесят два.
NEH|7|34|Сыновей Елама другого тысяча двести пятьдесят четыре.
NEH|7|35|Сыновей Харима триста двадцать.
NEH|7|36|Уроженцев Иерихона триста сорок пять.
NEH|7|37|Уроженцев Лода, Хадида и Оно семьсот двадцать один.
NEH|7|38|Уроженцев Сенаи три тысячи девятьсот тридцать.
NEH|7|39|Священников, сыновей Иедаии, из дома Иисусова, девятьсот семьдесят три.
NEH|7|40|Сыновей Иммера тысяча пятьдесят два.
NEH|7|41|Сыновей Пашхура тысяча двести сорок семь.
NEH|7|42|Сыновей Харима тысяча семнадцать.
NEH|7|43|Левитов: сыновей Иисуса, из [дома] Кадмиилова, из дома сыновей Годевы, семьдесят четыре.
NEH|7|44|Певцов: сыновей Асафа сто сорок восемь.
NEH|7|45|Привратники: сыновья Шаллума, сыновья Атера, сыновья Талмона, сыновья Аккува, сыновья Хатиты, сыновья Шовая – сто тридцать восемь.
NEH|7|46|Нефинеи: сыновья Цихи, сыновья Хасуфы, сыновья Таббаофа,
NEH|7|47|сыновья Кироса, сыновья Сии, сыновья Фадона,
NEH|7|48|сыновья Леваны, сыновья Хагавы, сыновья Салмая,
NEH|7|49|сыновья Ханана, сыновья Гиддела, сыновья Гахара,
NEH|7|50|сыновья Реаии, сыновья Рецина, сыновья Некоды,
NEH|7|51|сыновья Газзама, сыновья Уззы, сыновья Пасеаха,
NEH|7|52|сыновья Весая, сыновья Меунима, сыновья Нефишсима,
NEH|7|53|сыновья Бакбука, сыновья Хакуфы, сыновья Хархура,
NEH|7|54|сыновья Бацлифа, сыновья Мехиды, сыновья Харши,
NEH|7|55|сыновья Баркоса, сыновья Сисары, сыновья Фамаха,
NEH|7|56|сыновья Нециаха, сыновья Хатифы.
NEH|7|57|Сыновья рабов Соломоновых: сыновья Сотая, сыновья Соферефа, сыновья Фериды,
NEH|7|58|сыновья Иаалы, сыновья Даркона, сыновья Гиддела,
NEH|7|59|сыновья Сафатии, сыновья Хаттила, сыновья Похереф – Гаццевайима, сыновья Амона.
NEH|7|60|Всех нефинеев и сыновей рабов Соломоновых триста девяносто два.
NEH|7|61|И вот вышедшие из Тел–Мелаха, Тел–Харши, Херув–Аддона и Иммера; но они не могли показать о поколении своем и о племени своем, от Израиля ли они.
NEH|7|62|Сыновья Делаии, сыновья Товии, сыновья Некоды – шестьсот сорок два.
NEH|7|63|И из священников: сыновья Ховаии, сыновья Гаккоца, сыновья Верзеллия, который взял жену из дочерей Верзеллия Галаадитянина и стал называться их именем.
NEH|7|64|Они искали родословной своей записи, и не нашлось, и потому исключены из священства.
NEH|7|65|И Тиршафа сказал им, чтоб они не ели великой святыни, доколе не восстанет священник с уримом и туммимом.
NEH|7|66|Все общество вместе [состояло] из сорока двух тысяч трехсот шестидесяти [человек],
NEH|7|67|кроме рабов их и рабынь их, которых было семь тысяч триста тридцать семь; и при них певцов и певиц двести сорок пять.
NEH|7|68|Коней у них было семьсот тридцать шесть, лошаков у них двести сорок пять,
NEH|7|69|верблюдов четыреста тридцать пять, ослов шесть тысяч семьсот двадцать.
NEH|7|70|Некоторые главы поколений дали вклады на производство работ. Тиршафа дал в сокровищницу золотом тысячу драхм, пятьдесят чаш, пятьсот тридцать священнических одежд.
NEH|7|71|И некоторые из глав поколений дали в сокровищницу на производство работ двадцать тысяч драхм золота и две тысячи двести мин серебра.
NEH|7|72|Прочие из народа дали двадцать тысяч драхм золота и две тысячи мин серебра и шестьдесят семь священнических одежд.
NEH|7|73|И стали жить священники и левиты, и привратники и певцы, и народ и нефинеи, и весь Израиль в городах своих.
NEH|8|1|Когда наступил седьмой месяц, и сыны Израилевы [жили] по городам своим, тогда собрался весь народ, как один человек, на площадь, которая пред Водяными воротами, и сказали книжнику Ездре, чтобы он принес книгу закона Моисеева, который заповедал Господь Израилю.
NEH|8|2|И принес священник Ездра закон пред собрание мужчин и женщин, и всех, которые могли понимать, в первый день седьмого месяца;
NEH|8|3|и читал из него на площади, которая пред Водяными воротами, от рассвета до полудня, пред мужчинами и женщинами и всеми, которые могли понимать; и уши всего народа [были приклонены] к книге закона.
NEH|8|4|Книжник Ездра стоял на деревянном возвышении, которое для сего сделали, а подле него, по правую руку его, стояли Маттифия и Шема, и Анаия и Урия, и Хелкия и Маасея, а по левую руку его Федаия и Мисаил, и Малхия и Хашум, и Хашбаддана, и Захария и Мешуллам.
NEH|8|5|И открыл Ездра книгу пред глазами всего народа, потому что он стоял выше всего народа. И когда он открыл ее, весь народ встал.
NEH|8|6|И благословил Ездра Господа Бога великого. И весь народ отвечал: аминь, аминь, поднимая вверх руки свои, – и поклонялись и повергались пред Господом лицем до земли.
NEH|8|7|Иисус, Ванаия, Шеревия, Иамин, Аккув, Шавтай, Годия, Маасея, Клита, Азария, Иозавад, Ханан, Фелаия и левиты поясняли народу закон, между тем как народ стоял на своем месте.
NEH|8|8|И читали из книги, из закона Божия, внятно, и присоединяли толкование, и [народ] понимал прочитанное.
NEH|8|9|Тогда Неемия, он же Тиршафа, и книжник Ездра, священник, и левиты, учившие народ, сказали всему народу: день сей свят Господу Богу вашему; не печальтесь и не плачьте, потому что весь народ плакал, слушая слова закона.
NEH|8|10|И сказал им: пойдите, ешьте тучное и пейте сладкое, и посылайте части тем, у кого ничего не приготовлено, потому что день сей свят Господу нашему. И не печальтесь, потому что радость пред Господом – подкрепление для вас.
NEH|8|11|И левиты успокаивали весь народ, говоря: перестаньте, ибо день сей свят, не печальтесь.
NEH|8|12|И пошел весь народ есть, и пить, и посылать части, и праздновать с великим веселием, ибо поняли слова, которые сказали им.
NEH|8|13|На другой день собрались главы поколений от всего народа, священники и левиты к книжнику Ездре, чтобы он изъяснял им слова закона.
NEH|8|14|И нашли написанное в законе, который Господь дал чрез Моисея, чтобы сыны Израилевы в седьмом месяце, в праздник, жили в кущах.
NEH|8|15|И потому объявили и провозгласили по всем городам своим и в Иерусалиме, говоря: пойдите на гору и несите ветви маслины садовой и ветви маслины дикой, и ветви миртовые и ветви пальмовые, и ветви [других] широколиственных дерев, чтобы сделать кущи по написанному.
NEH|8|16|И пошел народ, и принесли, и сделали себе кущи, каждый на своей кровле и на дворах своих, и на дворах дома Божия, и на площади у Водяных ворот, и на площади у Ефремовых ворот.
NEH|8|17|Все общество возвратившихся из плена сделало кущи и жило в кущах. От дней Иисуса, сына Навина, до этого дня не делали так сыны Израилевы. Радость была весьма великая.
NEH|8|18|И читали из книги закона Божия каждый день, от первого дня до последнего дня. И праздновали праздник семь дней, а в восьмой день попразднество по уставу.
NEH|9|1|В двадцать четвертый день этого месяца собрались все сыны Израилевы, постящиеся и во вретищах и с пеплом на головах своих.
NEH|9|2|И отделилось семя Израилево от всех инородных, и встали и исповедывались во грехах своих и в преступлениях отцов своих.
NEH|9|3|И стояли на своем месте, и четверть дня читали из книги закона Господа Бога своего, и четверть исповедывались и поклонялись Господу Богу своему.
NEH|9|4|И стали на возвышенное место левитов: Иисус, Вания, Кадмиил, Шевания, Вунний, Шеревия, Вания, Хенани, и громко взывали к Господу Богу своему.
NEH|9|5|И сказали левиты – Иисус, Кадмиил, Вания, Хашавния, Шеревия, Годия, Шевания, Петахия: встаньте, славьте Господа Бога вашего, от века и до века. Да славословят достославное и превысшее всякого славословия и хвалы имя Твое!
NEH|9|6|Ты, Господи, един, Ты создал небо, небеса небес и все воинство их, землю и все, что на ней, моря и все, что в них, и Ты живишь все сие, и небесные воинства Тебе поклоняются.
NEH|9|7|Ты Сам, Господи Боже, избрал Аврама, и вывел его из Ура Халдейского, и дал ему имя Авраама,
NEH|9|8|и нашел сердце его верным пред Тобою, и заключил с ним завет, чтобы дать семени его землю Хананеев, Хеттеев, Аморреев, Ферезеев, Иевусеев и Гергесеев. И Ты исполнил слово Свое, потому что Ты праведен.
NEH|9|9|Ты увидел бедствие отцов наших в Египте и услышал вопль их у Чермного моря,
NEH|9|10|и явил знамения и чудеса над фараоном и над всеми рабами его, и над всем народом земли его, так как Ты знал, что они надменно поступали с ними, и сделал Ты Себе имя до сего дня.
NEH|9|11|Ты рассек пред ними море, и они среди моря прошли посуху, и гнавшихся за ними Ты поверг в глубины, как камень в сильные воды.
NEH|9|12|В столпе облачном Ты вел их днем и в столпе огненном – ночью, чтоб освещать им путь, по которому идти им.
NEH|9|13|И снисшел Ты на гору Синай и говорил с ними с неба, и дал им суды справедливые, законы верные, уставы и заповеди добрые.
NEH|9|14|И указал им святую Твою субботу и заповеди, и уставы и закон преподал им чрез раба Твоего Моисея.
NEH|9|15|И хлеб с неба Ты давал им в голоде их, и воду из камня источал им в жажде их, и сказал им, чтоб они пошли и овладели землею, которую Ты, подняв руку Твою, [клялся] дать им.
NEH|9|16|Но они и отцы наши упрямствовали, и шею свою держали упруго, и не слушали заповедей Твоих;
NEH|9|17|не захотели повиноваться и не вспомнили чудных дел Твоих, которые Ты делал с ними, и держали шею свою упруго, и, по упорству своему, поставили над собою вождя, чтобы возвратиться в рабство свое. Но Ты Бог, любящий прощать, благий и милосердый, долготерпеливый и многомилостивый, и Ты не оставил их.
NEH|9|18|И хотя они сделали себе литаго тельца, и сказали: вот бог твой, который вывел тебя из Египта, и хотя делали великие оскорбления,
NEH|9|19|но Ты, по великому милосердию Твоему, не оставлял их в пустыне; столп облачный не отходил от них днем, чтобы вести их по пути, и столп огненный – ночью, чтобы светить им на пути, по которому им идти.
NEH|9|20|И Ты дал им Духа Твоего благого, чтобы наставлять их, и манну Твою не отнимал от уст их, и воду давал им для утоления жажды их.
NEH|9|21|Сорок лет Ты питал их в пустыне; они ни в чем не терпели недостатка; одежды их не ветшали, и ноги их не пухли.
NEH|9|22|И Ты дал им царства и народы и разделил им, и они овладели землею Сигона, и землею царя Есевонского, и землею Ога, царя Васанского.
NEH|9|23|И сыновей их Ты размножил, как звезды небесные, и ввел их в землю, о которой Ты говорил отцам их, что они придут владеть [ею].
NEH|9|24|И вошли сыновья их, и овладели землею. И Ты покорил им жителей земли, Хананеев, и отдал их в руки их, и царей их, и народы земли, чтобы они поступали с ними по своей воле.
NEH|9|25|И заняли они укрепленные города и тучную землю, и взяли во владение домы, наполненные всяким добром, водоемы, высеченные [из камня], виноградные и масличные сады и множество дерев [с плодами] для пищи. Они ели, насыщались, тучнели и наслаждались по великой благости Твоей;
NEH|9|26|и сделались упорны и возмутились против Тебя, и презрели закон Твой, убивали пророков Твоих, которые увещевали их обратиться к Тебе, и делали великие оскорбления.
NEH|9|27|И Ты отдал их в руки врагов их, которые теснили их. Но когда, в тесное для них время, они взывали к Тебе, Ты выслушивал их с небес и, по великому милосердию Твоему, давал им спасителей, и они спасали их от рук врагов их.
NEH|9|28|Когда же успокаивались, то снова начинали делать зло пред лицем Твоим, и Ты отдавал их в руки неприятелей их, и они господствовали над ними. Но когда они опять взывали к Тебе, Ты выслушивал их с небес и, по великому милосердию Твоему, избавлял их многократно.
NEH|9|29|Ты напоминал им обратиться к закону Твоему, но они упорствовали и не слушали заповедей Твоих, и отклонялись от уставов Твоих, которыми жил бы человек, если бы исполнял их, и хребет [свой] сделали упорным, и шею свою держали упруго, и не слушали.
NEH|9|30|Ожидая их [обращения], Ты медлил многие годы и напоминал им Духом Твоим чрез пророков Твоих, но они не слушали. И Ты предал их в руки иноземных народов.
NEH|9|31|Но, по великому милосердию Твоему, Ты не истребил их до конца, и не оставлял их, потому что Ты Бог благий и милостивый.
NEH|9|32|И ныне, Боже наш, Боже великий, сильный и страшный, хранящий завет и милость! да не будет малым пред лицем Твоим все страдание, которое постигло нас, царей наших, князей наших, и священников наших, и пророков наших, и отцов наших и весь народ Твой от дней царей Ассирийских до сего дня.
NEH|9|33|Во всем постигшем нас Ты праведен, потому что Ты делал по правде, а мы виновны.
NEH|9|34|Цари наши, князья наши, священники наши и отцы наши не исполняли закона Твоего, и не внимали заповедям Твоим и напоминаниям Твоим, которыми Ты напоминал им.
NEH|9|35|И в царстве своем, при великом добре Твоем, которое Ты давал им, и на обширной и тучной земле, которую Ты отделил им, они не служили Тебе и не обращались от злых дел своих.
NEH|9|36|И вот, мы ныне рабы; на той земле, которую Ты дал отцам нашим, чтобы питаться ее плодами и ее добром, вот, мы рабствуем.
NEH|9|37|И произведения свои она во множестве приносит для царей, которым Ты покорил нас за грехи наши. И телами нашими и скотом нашим они владеют по своему произволу, и мы в великом стеснении.
NEH|9|38|По всему этому мы даем твердое обязательство и подписываем, и на подписи печать князей наших, левитов наших и священников наших.
NEH|10|1|Приложившие печати были: Неемия–Тиршафа, сын Гахалии, и Седекия,
NEH|10|2|Сераия, Азария, Иеремия,
NEH|10|3|Пашхур, Амария, Малхия,
NEH|10|4|Хаттуш, Шевания, Маллух,
NEH|10|5|Харим, Меремоф, Овадия,
NEH|10|6|Даниил, Гиннефон, Варух,
NEH|10|7|Мешуллам, Авия, Миямин,
NEH|10|8|Маазия, Вилгай, Шемаия: это священники.
NEH|10|9|Левиты: Иисус, сын Азании, Биннуй, из сыновей Хенадада, Кадмиил,
NEH|10|10|и братья их: Шевания, Годия, Клита, Фелаия, Ханан,
NEH|10|11|Миха, Рехов, Хашавия,
NEH|10|12|Закхур, Шеревия, Шевания,
NEH|10|13|Годия, Ваний, Венинуй.
NEH|10|14|Главы народа: Парош, Пахаф–Моав, Елам, Заффу, Вания,
NEH|10|15|Вунний, Азгар, Бевай,
NEH|10|16|Адония, Бигвай, Адин,
NEH|10|17|Атер, Езекия, Азур,
NEH|10|18|Годия, Хашум, Бецай,
NEH|10|19|Хариф, Анафоф, Невай,
NEH|10|20|Магпиаш, Мешуллам, Хезир,
NEH|10|21|Мешезавел, Садок, Иаддуй,
NEH|10|22|Фелатия, Ханан, Анаия,
NEH|10|23|Осия, Ханания, Хашшув,
NEH|10|24|Лохеш, Пилха, Шовек,
NEH|10|25|Рехум, Хашавна, Маасея,
NEH|10|26|Ахия, Ханан, Анан,
NEH|10|27|Маллух, Харим, Ваана.
NEH|10|28|И прочий народ, священники, левиты, привратники, певцы, нефинеи и все, отделившиеся от народов иноземных к закону Божию, жены их, сыновья их и дочери их, все, которые могли понимать,
NEH|10|29|пристали к братьям своим, к почетнейшим из них, и вступили в обязательство с клятвою и проклятием – поступать по закону Божию, который дан рукою Моисея, раба Божия, и соблюдать и исполнять все заповеди Господа Бога нашего, и уставы Его и предписания Его,
NEH|10|30|и не отдавать дочерей своих иноземным народам, и их дочерей не брать за сыновей своих;
NEH|10|31|и когда иноземные народы будут привозить товары и все продажное в субботу, не брать у них в субботу и в священный день, и в седьмой год оставлять долги всякого рода.
NEH|10|32|И поставили мы себе в закон давать от себя по трети сикля в год на потребности для дома Бога нашего:
NEH|10|33|на хлебы предложения, на всегдашнее хлебное приношение и на всегдашнее всесожжение, на субботы, на новомесячия, на праздники, на священные вещи и на жертвы за грех для очищения Израиля, и на все, совершаемое в доме Бога нашего.
NEH|10|34|И бросили мы жребии о доставке дров, священники, левиты и народ, когда которому поколению нашему в назначенные времена, из года в год, привозить [их] к дому Бога нашего, чтоб они горели на жертвеннике Господа Бога нашего, по написанному в законе.
NEH|10|35|[И обязались мы] каждый год приносить в дом Господень начатки с земли нашей и начатки всяких плодов со всякого дерева;
NEH|10|36|также приводить в дом Бога нашего к священникам, служащим в доме Бога нашего, первенцев из сыновей наших и из скота нашего, как написано в законе, и первородное от крупного и мелкого скота нашего.
NEH|10|37|И начатки из молотого хлеба нашего и приношений наших, и плодов со всякого дерева, вина и масла мы будем доставлять священникам в кладовые при доме Бога нашего и десятину с земли нашей левитам. Они, левиты, будут брать десятину во всех городах, где у нас земледелие.
NEH|10|38|При левитах, когда они будут брать левитскую десятину, будет находиться священник, сын Аарона, чтобы левиты десятину из своих десятин отвозили в дом Бога нашего в комнаты, [отделенные] для кладовой,
NEH|10|39|потому что в эти комнаты как сыны Израилевы, так и левиты должны доставлять приносимое в дар: хлеб, вино и масло. Там священные сосуды, и служащие священники, и привратники, и певцы. И мы не оставим дома Бога нашего.
NEH|11|1|И жили начальники народа в Иерусалиме, а прочие из народа бросили жребии, чтоб одна из десяти частей их шла на жительство в святой город Иерусалим, а девять [оставались] в [прочих] городах.
NEH|11|2|И благословил народ всех, которые добровольно согласились жить в Иерусалиме.
NEH|11|3|Вот главы страны, которые жили в Иерусалиме, – а в городах Иудеи жили, всякий в своем владении, по городам своим: Израильтяне, священники, левиты и нефинеи и сыновья рабов Соломоновых; –
NEH|11|4|в Иерусалиме жили из сыновей Иуды и из сыновей Вениамина. Из сыновей Иуды: Афаия, сын Уззии, сын Захарии, сын Амарии, сын Сафатии, сын Малелеила, из сыновей Фареса,
NEH|11|5|и Маасея, сын Варуха, сын Колхозея, сын Хазаии, сын Адаии, сын Иоиарива, сын Захарии, сын Шилония.
NEH|11|6|Всех сыновей Фареса, живших в Иерусалиме, четыреста шестьдесят восемь, люди отличные.
NEH|11|7|И вот сыновья Вениамина: Саллу, сын Мешуллама, сын Иоеда, сын Федаии, сын Колаии, сын Маасеи, сын Ифиила, сын Исаии,
NEH|11|8|и за ним Габбай, Саллай – девятьсот двадцать восемь.
NEH|11|9|Иоиль, сын Зихри, был начальником над ними, а Иуда, сын Сенуи, был вторым над городом.
NEH|11|10|Из священников: Иедаия, сын Иоиарива, Иахин,
NEH|11|11|Сераия, сын Хелкии, сын Мешуллама, сын Садока, сын Мераиофа, сын Ахитува, начальствующий в доме Божием,
NEH|11|12|и братья их, отправлявшие службу в доме [Божием] – восемьсот двадцать два; и Адаия, сын Иерохама, сын Фелалии, сын Амция, сын Захарии, сын Пашхура, сын Малхии,
NEH|11|13|и братья его, главы поколений – двести сорок два; и Амашсай, сын Азариила, сын Ахзая, сын Мешиллемофа, сын Иммера,
NEH|11|14|и братья его, люди отличные – сто двадцать восемь. Начальником над ними был Завдиил, сын Гагедолима.
NEH|11|15|А из левитов: Шемаия, сын Хашшува, сын Азрикама, сын Хашавии, сын Вунния,
NEH|11|16|и Шавфай, и Иозавад, из глав левитов по внешним делам дома Божия,
NEH|11|17|и Матфания, сын Михи, сын Завдия, сын Асафа, главный начинатель славословия при молитве, и Бакбукия, второй [по нем] из братьев его, и Авда, сын Шаммуя, сын Галала, сын Идифуна.
NEH|11|18|Всех левитов во святом городе двести восемьдесят четыре.
NEH|11|19|А привратники: Аккув, Талмон и братья их, содержавшие стражу у ворот – сто семьдесят два.
NEH|11|20|Прочие Израильтяне, священники, левиты [жили] по всем городам Иудеи, каждый в своем уделе.
NEH|11|21|А нефинеи жили в Офеле; над нефинеями Циха и Гишфа.
NEH|11|22|Начальником над левитами в Иерусалиме был Уззий, сын Вания, сын Хашавии, сын Матфании, сын Михи, из сыновей Асафовых, которые были певцами при служении в доме Божием,
NEH|11|23|потому что от царя [было] о них [особое] повеление, и назначено было на каждый день для певцов определенное содержание.
NEH|11|24|И Петахия, сын Мешезавела, из сыновей Зары, сына Иуды, был доверенным от царя по всяким делам, [касающимся] до народа.
NEH|11|25|Из [живших] же в селах, на полях своих, сыновья Иуды жили в Кириаф–Арбе и зависящих от нее городах, в Дивоне и зависящих от него городах, в Иекавцеиле и селах его,
NEH|11|26|в Иешуе, в Моладе и в Беф–Палете,
NEH|11|27|в Хацар–Шуале, в Вирсавии и зависящих от нее городах,
NEH|11|28|в Секелаге, в Мехоне и зависящих от нее городах,
NEH|11|29|в Ен–Риммоне, в Цоре и в Иармуфе,
NEH|11|30|в Заноахе, Одолламе и селах их, в Лахисе и на полях его, в Азеке и зависящих от нее городах. Они расположились от Вирсавии и до долины Енномовой.
NEH|11|31|Сыновья Вениаминовы, [начиная] от Гевы, в Михмасе, Гае, в Вефиле и зависящих от него городах,
NEH|11|32|в Анафофе, Нове, Анании,
NEH|11|33|Гацоре, Раме, Гиффаиме,
NEH|11|34|Хадиде, Цевоиме, Неваллате,
NEH|11|35|Лоде, Оно, в долине Харашиме.
NEH|11|36|И левиты имели жилища свои в участках Иуды и Вениамина.
NEH|12|1|Вот священники и левиты, которые пришли с Зоровавелем, сыном Салафииловым, и с Иисусом: Сераия, Иеремия, Ездра,
NEH|12|2|Амария, Маллух, Хаттуш,
NEH|12|3|Шехания, Рехум, Меремоф,
NEH|12|4|Иддо, Гиннефой, Авия,
NEH|12|5|Миямин, Маадия, Вилга,
NEH|12|6|Шемаия, Иоиарив, Иедаия,
NEH|12|7|Саллу, Амок, Хелкия, Иедаия. Это главы священников и братья их во дни Иисуса.
NEH|12|8|А левиты: Иисус, Биннуй, Кадмиил, Шеревия, Иуда, Матфания, [главный] при славословии, он и братья его,
NEH|12|9|и Бакбукия и Унний, братья их, наряду с ними [державшие] стражу.
NEH|12|10|Иисус родил Иоакима, Иоаким родил Елиашива, Елиашив родил Иоиаду,
NEH|12|11|Иоиада родил Ионафана, Ионафан родил Иаддуя.
NEH|12|12|Во дни Иоакима были священники, главы поколений: из [дома] Сераии Мераия, из [дома] Иеремии Ханания,
NEH|12|13|из [дома] Ездры Мешуллам, из [дома] Амарии Иоханан,
NEH|12|14|из [дома] Мелиху Ионафан, из [дома] Шевании Иосиф,
NEH|12|15|из [дома] Харима Адна, из [дома] Мераиофа Хелкия,
NEH|12|16|из [дома] Иддо Захария, из [дома] Гиннефона Мешуллам,
NEH|12|17|из [дома] Авии Зихрий, из [дома] Миниамина, из [дома] Моадии Пилтай,
NEH|12|18|из [дома] Вилги Шаммуй, из [дома] Шемаии Ионафан,
NEH|12|19|из [дома] Иоиарива Мафнай, из [дома] Иедаии Уззий,
NEH|12|20|из [дома] Саллая Каллай, из [дома] Амока Евер,
NEH|12|21|из [дома] Хелкии Хашавия, из [дома] Иедаии Нафанаил.
NEH|12|22|Левиты, главы поколений, внесены в запись во дни Елиашива, Иоиады, Иоханана и Иаддуя, и также священники в царствование Дария Персидского.
NEH|12|23|Сыновья Левия, главы поколений, вписаны в летописи до дней Иоханана, сына Елиашивова.
NEH|12|24|Главы левитов: Хашавия, Шеревия, и Иисус, сын Кадмиила, и братья их, при них [поставленные] для славословия при благодарениях, по установлению Давида, человека Божия – смена за сменою.
NEH|12|25|Матфания, Бакбукия, Овадия, Мешуллам, Талмон, Аккув – стражи, привратники на страже у порогов ворот.
NEH|12|26|Они были во дни Иоакима, сына Иисусова, сына Иоседекова, и во дни областеначальника Неемии и книжника Ездры, священника.
NEH|12|27|При освящении стены Иерусалимской потребовали левитов из всех мест их, приказывая им придти в Иерусалим для совершения освящения и радостного празднества со славословиями и песнями при [звуке] кимвалов, псалтирей и гуслей.
NEH|12|28|И собрались сыновья певцов из округа Иерусалимского и из сел Нетофафских,
NEH|12|29|и из Беф–Гаггилгала, и с полей Гевы и Азмавета, потому что певцы выстроили себе села в окрестностях Иерусалима.
NEH|12|30|И очистились священники и левиты, и очистили народ и ворота, и стену.
NEH|12|31|Тогда я повел начальствующих в Иудее на стену и поставил два больших хора для шествия, и один из них шел по правой стороне стены к Навозным воротам.
NEH|12|32|За ними шел Гошаия и половина начальствующих в Иудее,
NEH|12|33|Азария, Ездра и Мешуллам,
NEH|12|34|Иуда и Вениамин, и Шемаия и Иеремия,
NEH|12|35|а из сыновей священнических с трубами: Захария, сын Ионафана, сын Шемаии, сын Матфании, сын Михея, сын Закхура, сын Асафа,
NEH|12|36|и братья его: Шемаия, Азариил, Милалай, Гилалай, Маай, Нафанаил, Иуда и Хананий с музыкальными орудиями Давида, человека Божия, и книжник Ездра впереди них.
NEH|12|37|Подле ворот Источника, против них, они взошли по ступеням города Давидова, по лестнице, ведущей на стену сверх дома Давидова до Водяных ворот к востоку.
NEH|12|38|Другой хор шел напротив них, и за ним я и половина народа, по стене от Печной башни и до широкой стены,
NEH|12|39|и от ворот Ефремовых, мимо старых ворот и ворот Рыбных, и башни Хананела, и башни Меа, к Овечьим воротам, и остановились у ворот Темничных.
NEH|12|40|Потом оба хора стали у дома Божия, и я и половина начальствующих со мною,
NEH|12|41|и священники: Елиаким, Маасея, Миниамин, Михей, Елиоенай, Захария, Ханания с трубами,
NEH|12|42|и Маасея и Шемаия, и Елеазар и Уззий, и Иоханан и Малхия, и Елам и Езер. И пели певцы громко; главным [у них был] Израхия.
NEH|12|43|И приносили в тот день большие жертвы и веселились, потому что Бог дал им великую радость. Веселились и жены и дети, и веселие Иерусалима далеко было слышно.
NEH|12|44|В тот же день приставлены были люди к кладовым комнатам для приношений начатков и десятин, чтобы собирать с полей при городах части, положенные законом для священников и левитов, потому что Иудеям радостно было [смотреть] на стоящих священников и левитов,
NEH|12|45|которые совершали службу Богу своему и дела очищения и были певцами и привратниками по установлению Давида и сына его Соломона.
NEH|12|46|Ибо издавна во дни Давида и Асафа были установлены главы певцов и песни Богу, хвалебные и благодарственные.
NEH|12|47|Все Израильтяне во дни Зоровавеля и во дни Неемии давали части певцам и привратникам на каждый день и отдавали святыни левитам, а левиты отдавали святыни сынам Аарона.
NEH|13|1|В тот день читано было из книги Моисеевой вслух народа и найдено написанное в ней: Аммонитянин и Моавитянин не может войти в общество Божие во веки,
NEH|13|2|потому что они не встретили сынов Израиля с хлебом и водою и наняли против него Валаама, чтобы проклясть его, но Бог наш обратил проклятие в благословение.
NEH|13|3|Услышав этот закон, они отделили все иноплеменное от Израиля.
NEH|13|4|А прежде того священник Елиашив, приставленный к комнатам при доме Бога нашего, близкий родственник Товии,
NEH|13|5|отделал для него большую комнату, в которую прежде клали хлебное приношение, ладан и сосуды, и десятины хлеба, вина и масла, положенные законом для левитов, певцов и привратников, и приношения для священников.
NEH|13|6|Когда все это [происходило], я не был в Иерусалиме, потому что в тридцать втором году Вавилонского царя Артаксеркса я ходил к царю, и по прошествии нескольких дней [опять] выпросился у царя.
NEH|13|7|Когда я пришел в Иерусалим и узнал о худом деле, которое сделал Елиашив, отделав для Товии комнату на дворах дома Божия,
NEH|13|8|тогда мне было весьма неприятно, и я выбросил все домашние вещи Товиины вон из комнаты
NEH|13|9|и сказал, чтобы очистили комнаты, и велел опять внести туда сосуды дома Божия, хлебное приношение и ладан.
NEH|13|10|Еще узнал я, что части левитам не отдаются, и что левиты и певцы, делавшие [свое] дело, разбежались, каждый на свое поле.
NEH|13|11|Я сделал [за это] выговор начальствующим и сказал: зачем оставлен нами дом Божий? И я собрал их и поставил их на место их.
NEH|13|12|И все Иудеи стали приносить десятины хлеба, вина и масла в кладовые.
NEH|13|13|И приставил я к кладовым Шелемию священника и Садока книжника и Федаию из левитов, и при них Ханана, сына Закхура, сына Матфании, потому что они считались верными. И на них [возложено] раздавать части братьям своим.
NEH|13|14|Помяни меня за это, Боже мой, и не изгладь усердных дел моих, которые я сделал для дома Бога моего и для служения при нем!
NEH|13|15|В те дни я увидел в Иудее, что в субботу топчут точила, возят снопы и навьючивают ослов вином, виноградом, смоквами и всяким грузом, и отвозят в субботний день в Иерусалим. И я строго выговорил [им] в тот же день, когда они продавали съестное.
NEH|13|16|И Тиряне жили в [Иудее] и привозили рыбу и всякий товар и продавали в субботу жителям Иудеи и в Иерусалиме.
NEH|13|17|И я сделал выговор знатнейшим из Иудеев и сказал им: зачем вы делаете такое зло и оскверняете день субботний?
NEH|13|18|Не так ли поступали отцы ваши, и за то Бог наш навел на нас и на город сей все это бедствие? А вы увеличиваете гнев [Его] на Израиля, оскверняя субботу.
NEH|13|19|После сего, когда смеркалось у ворот Иерусалимских, перед субботою, я велел запирать двери и сказал, чтобы не отпирали их до [утра] после субботы. И слуг моих я ставил у ворот, чтобы никакая ноша не проходила в день субботний.
NEH|13|20|И ночевали торговцы и продавцы всякого товара вне Иерусалима раз и два.
NEH|13|21|Но я строго выговорил им и сказал им: зачем вы ночуете возле стены? Если сделаете это в другой раз, я наложу руку на вас. С того времени они не приходили в субботу.
NEH|13|22|И сказал я левитам, чтобы они очистились и пришли содержать стражу у ворот, дабы святить день субботний. И за сие помяни меня, Боже мой, и пощади меня по великой милости Твоей!
NEH|13|23|Еще в те дни я видел Иудеев, которые взяли себе жен из Азотянок, Аммонитянок и Моавитянок;
NEH|13|24|и от того сыновья их в половину говорят по–азотски, или языком других народов, и не умеют говорить по–иудейски.
NEH|13|25|Я сделал за это выговор и проклинал их, и некоторых из мужей бил, рвал у них волоса и заклинал их Богом, чтобы они не отдавали дочерей своих за сыновей их и не брали дочерей их за сыновей своих и за себя.
NEH|13|26|Не из–за них ли, [говорил я,] грешил Соломон, царь Израилев? У многих народов не было такого царя, как он. Он был любим Богом своим, и Бог поставил его царем над всеми Израильтянами; и однако же чужеземные жены ввели в грех и его.
NEH|13|27|И можно ли нам слышать о вас, что вы делаете все сие великое зло, грешите пред Богом нашим, принимая в сожительство чужеземных жен?
NEH|13|28|И из сыновей Иоиады, сына великого священника Елиашива, один был зятем Санаваллата, Хоронита. Я прогнал его от себя.
NEH|13|29|Воспомяни им, Боже мой, что они опорочили священство и завет священнический и левитский!
NEH|13|30|Так очистил я их от всего чужеземного и восстановил службы священников и левитов, каждого в деле его,
NEH|13|31|и доставку дров в назначенные времена и начатки. Помяни меня, Боже мой, во благо [мне]!
