MAL|1|1|耶和華的話，藉 瑪拉基 傳給 以色列 的默示。
MAL|1|2|耶和華說：「我曾愛你們。」你們卻說：「你在何事上愛我們呢？」耶和華說：「 以掃 不是 雅各 的哥哥嗎？我卻愛 雅各 ，
MAL|1|3|惡 以掃 ，使他的山嶺荒涼，把他的地業交給曠野的野狗。」
MAL|1|4|以東 若說：「我們雖被毀壞，卻要重建荒廢之處。」萬軍之耶和華如此說：「任他們建造，我必拆毀；人必稱他們為『邪惡之境』，為『耶和華永遠惱怒之民』。」
MAL|1|5|你們必親眼看見，你們要說：「耶和華在 以色列 疆界之外必尊為大！」
MAL|1|6|萬軍之耶和華對你們說：「兒子孝敬父親，僕人敬畏主人；我既為父親，孝敬我的在哪裏呢？我既為主人，敬畏我的在哪裏呢？你們這些藐視我名的祭司啊！」你們卻說：「我們在何事上藐視你的名呢？」
MAL|1|7|「你們將不潔淨的食物獻在我的祭壇上，卻說：『我們在何事上使你不潔淨呢？』你們說，耶和華的供桌是可藐視的。
MAL|1|8|你們將瞎眼的獻為祭物，這不算為惡嗎？將瘸腿的、有病的獻上，這不算為惡嗎？那麼，請把這些獻給你的省長，他豈會悅納你 ，豈會抬舉你呢？這是萬軍之耶和華說的。」
MAL|1|9|現在我勸你們要懇求上帝，好讓他施恩給我們。這事既出於你們的手，他豈會抬舉你們任何人呢？這是萬軍之耶和華說的。
MAL|1|10|萬軍之耶和華說：「甚願你們中間有人把殿的門 關上，免得你們徒然在我壇上燒火。我不喜歡你們，也不從你們手中悅納供物。」
MAL|1|11|萬軍之耶和華說：「從日出之地到日落之處，我的名在列國中必尊為大。在各處，人必奉我的名燒香，獻潔淨的供物，因為我的名在列國中必尊為大。
MAL|1|12|你們卻褻瀆我的名，說：『主的供桌是不潔淨的，供桌上的果子和食物是可藐視的。』
MAL|1|13|你們又說：『看哪，這些事何等煩瑣！』並嗤之以鼻 。這是萬軍之耶和華說的。你們把搶來的、瘸腿的、有病的拿來獻上為祭，我豈能從你們手中悅納它呢？這是耶和華說的。
MAL|1|14|行詭詐的人是可詛咒的！他的群畜中雖有公羊，他許了願，卻將有殘疾的獻給主。因我是大君王，我的名在列國中是可畏的。這是萬軍之耶和華說的。」
MAL|2|1|現在，眾祭司啊，這誡命是給你們的。
MAL|2|2|萬軍之耶和華說：「你們若不聽，不放在心上，不將榮耀歸給我的名，我就使詛咒臨到你們，使你們的福分變為詛咒；其實我已經詛咒了你們的福分，因你們不把誡命放在心上。
MAL|2|3|看哪，我要斥責你們的後裔，把糞抹在你們臉上，就是你們祭牲 的糞。人要把你們和糞一起抬出去，
MAL|2|4|你們就知道我頒這誡命給你們，使我與 利未 所立的約可以常存。這是萬軍之耶和華說的。
MAL|2|5|我曾與他立生命和平安的約。我將這兩樣賜給他，使他存敬畏的心；他就敬畏我，懼怕我的名。
MAL|2|6|真實的訓誨在他口中，他的嘴唇中沒有不義。他以平安和正直與我同行，使許多人回轉離開罪孽。
MAL|2|7|祭司的嘴唇當守護知識，人也當從他口中尋求訓誨，因為他是萬軍之耶和華的使者。
MAL|2|8|你們卻偏離正道，使許多人在這訓誨上絆跌。你們破壞了我與 利未 人所立的約。這是萬軍之耶和華說的。
MAL|2|9|所以我使你們被眾百姓藐視，看為卑賤；因你們不遵守我的道，在律法上看人的情面 。」
MAL|2|10|我們豈不都有一位父嗎？豈不是一位上帝創造了我們嗎？為何互相行詭詐，褻瀆了上帝與我們列祖所立的約呢？
MAL|2|11|猶大 行事詭詐，在 以色列 和 耶路撒冷 中行了可憎的事；因為 猶大 人褻瀆耶和華所喜愛的聖殿，娶外邦神明的女子為妻。
MAL|2|12|凡做這事的，無論是清醒的 或回應的，即使獻供物給萬軍之耶和華，耶和華也要將他從 雅各 的帳棚中剪除。
MAL|2|13|你們又再做這樣的事，使哭泣和嘆息的眼淚遮蓋耶和華的祭壇，以致耶和華不再理會那供物，也不喜歡從你們的手中收納。
MAL|2|14|你們還說：「這是為甚麼呢？」因為耶和華在你和你年輕時所娶的妻之間作證。她雖是你的配偶，你誓約 的妻，你卻背棄她。
MAL|2|15|一個人如果還剩下一點靈性，他不會這麼做。這人在尋找甚麼呢？上帝的後裔！ 當謹守你們的靈性，誰也不可背棄年輕時所娶的妻。
MAL|2|16|耶和華－ 以色列 的上帝說：「我恨惡休妻的事和衣服外面披上暴力的人。所以當謹守你們的心，不可行詭詐。這是萬軍之耶和華說的。」
MAL|2|17|你們用言語使耶和華厭煩，卻說：「我們在何事上使他厭煩呢？」因為你們說：「凡行惡的，耶和華看為善，並且喜愛他們；」又說：「公平的上帝在哪裏呢？」
MAL|3|1|萬軍之耶和華說：「看哪，我要差遣我的使者在我前面預備道路。你們所尋求的主必忽然來到他的殿；立約的使者，就是你們所仰慕的，看哪，快要來到。」
MAL|3|2|他來的日子，誰能當得起呢？他顯現的時候，誰能立得住呢？因為他如煉金匠的火，如漂洗者的鹼。
MAL|3|3|他必坐下如煉淨銀子的人，必潔淨 利未 人，熬煉他們像金銀一樣；他們就憑公義獻供物給耶和華。
MAL|3|4|那時， 猶大 和 耶路撒冷 所獻的供物必蒙耶和華悅納，彷彿古時之日、上古之年。
MAL|3|5|萬軍之耶和華說：「我必臨近你們，施行審判。我必速速作見證，警戒那些行邪術的、犯姦淫的、起假誓的、剝削雇工工錢的、欺壓孤兒寡婦的、屈枉寄居者的和不敬畏我的人。」
MAL|3|6|「我－耶和華是不改變的；所以， 雅各 的子孫啊，你們不致滅亡。
MAL|3|7|從你們祖先的日子以來，你們就偏離我的律例而不遵守。現在你們要轉向我，我就轉向你們。這是萬軍之耶和華說的。你們卻說：『我們如何轉向呢？』
MAL|3|8|人豈可搶奪上帝呢？你們竟搶奪我！你們卻說：『我們在何事上搶奪你呢？』其實就是在你們當納的十分之一奉獻和當獻的供物上。
MAL|3|9|因你們全國上下都搶奪我的供物，詛咒就臨到你們身上。
MAL|3|10|你們要將當納的十分之一全然送入倉庫，使我家有糧，以此試試我，是否為你們敞開天上的窗戶，傾福與你們，甚至無處可容。這是萬軍之耶和華說的。
MAL|3|11|我必為你們斥責蝗蟲 ，不容牠毀壞你們的土產。你們田間的葡萄樹，果實未熟以先也不會掉落。這是萬軍之耶和華說的。
MAL|3|12|萬國必稱你們為有福的，因你們必成為喜樂之地。這是萬軍之耶和華說的。」
MAL|3|13|耶和華說：「你們用話頂撞我。」你們卻說：「我們說了甚麼話頂撞你呢？」
MAL|3|14|你們說：「事奉上帝是枉然，我們遵守上帝所吩咐的，在萬軍之耶和華面前哀痛而行，有甚麼益處呢？
MAL|3|15|現在，我們稱狂傲的人為有福，並且行惡的人得以建立；他們雖然試探上帝，卻得以逃脫。」
MAL|3|16|那時，敬畏耶和華的人彼此談論，耶和華側耳而聽，且有紀念冊在他面前，記錄那敬畏耶和華、思念他名的人。
MAL|3|17|萬軍之耶和華說：「在我所定的日子，他們必屬我，是我寶貴的產業。我必憐憫他們，如同人憐憫那服侍他的兒子。
MAL|3|18|那時你們必再一次 看出義人和惡人，事奉上帝和不事奉上帝的人有何差別。」
MAL|4|1|萬軍之耶和華說：「看哪，那日臨近，勢如燒著的火爐，凡狂傲的和行惡的都如碎秸，在那日被燒盡，根與枝條無一存留。
MAL|4|2|但是，對你們敬畏我名的人，必有公義的太陽出現，其光線 有醫治的能力。你們必出來跳躍如圈裏的牛犢。
MAL|4|3|你們必踐踏惡人；在我所定的日子，他們必成為你們腳掌下的灰塵。這是萬軍之耶和華說的。
MAL|4|4|「你們當記念我僕人 摩西 的律法，就是我在 何烈山 為 以色列 眾人所吩咐他的律例典章。
MAL|4|5|「看哪，耶和華大而可畏之日未到以前，我要差遣 以利亞 先知到你們那裏去。
MAL|4|6|他必使父親的心轉向兒女，兒女的心轉向父親，免得我來詛咒這地。」
