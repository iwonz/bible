JOEL|1|1|verbum Domini quod factum est ad Iohel filium Fatuhel
JOEL|1|2|audite hoc senes et auribus percipite omnes habitatores terrae si factum est istud in diebus vestris aut in diebus patrum vestrorum
JOEL|1|3|super hoc filiis vestris narrate et filii vestri filiis suis et filii eorum generationi alterae
JOEL|1|4|residuum erucae comedit lucusta et residuum lucustae comedit bruchus et residuum bruchi comedit rubigo
JOEL|1|5|expergescimini ebrii et flete et ululate omnes qui bibitis vinum in dulcedine quoniam periit ab ore vestro
JOEL|1|6|gens enim ascendit super terram meam fortis et innumerabilis dentes eius ut dentes leonis et molares eius ut catuli leonis
JOEL|1|7|posuit vineam meam in desertum et ficum meam decorticavit nudans spoliavit eam et proiecit albi facti sunt rami eius
JOEL|1|8|plange quasi virgo accincta sacco super virum pubertatis suae
JOEL|1|9|periit sacrificium et libatio de domo Domini luxerunt sacerdotes ministri Domini
JOEL|1|10|depopulata est regio luxit humus quoniam devastatum est triticum confusum est vinum elanguit oleum
JOEL|1|11|confusi sunt agricolae ululaverunt vinitores super frumento et hordeo quia periit messis agri
JOEL|1|12|vinea confusa est et ficus elanguit malogranatum et palma et malum et omnia ligna agri aruerunt quia confusum est gaudium a filiis hominum
JOEL|1|13|accingite vos et plangite sacerdotes ululate ministri altaris ingredimini cubate in sacco ministri Dei mei quoniam interiit de domo Dei vestri sacrificium et libatio
JOEL|1|14|sanctificate ieiunium vocate coetum congregate senes omnes habitatores terrae in domum Dei vestri et clamate ad Dominum
JOEL|1|15|a a a diei quia prope est dies Domini et quasi vastitas a potente veniet
JOEL|1|16|numquid non coram oculis vestris alimenta perierunt de domo Dei nostri laetitia et exultatio
JOEL|1|17|conputruerunt iumenta in stercore suo demolita sunt horrea dissipatae sunt apothecae quoniam confusum est triticum
JOEL|1|18|quid ingemuit animal mugierunt greges armenti quia non est pascua eis sed et greges pecorum disperierunt
JOEL|1|19|ad te Domine clamabo quia ignis comedit speciosa deserti et flamma succendit omnia ligna regionis
JOEL|1|20|sed et bestiae agri quasi area sitiens imbrem suspexerunt ad te quoniam exsiccati sunt fontes aquarum et ignis devoravit speciosa deserti
JOEL|2|1|canite tuba in Sion ululate in monte sancto meo conturbentur omnes habitatores terrae quia venit dies Domini quia prope est
JOEL|2|2|dies tenebrarum et caliginis dies nubis et turbinis quasi mane expansum super montes populus multus et fortis similis ei non fuit a principio et post eum non erit usque in annos generationis et generationis
JOEL|2|3|ante faciem eius ignis vorans et post eum exurens flamma quasi hortus voluptatis terra coram eo et post eum solitudo deserti neque est qui effugiat eum
JOEL|2|4|quasi aspectus equorum aspectus eorum et quasi equites sic current
JOEL|2|5|sicut sonitus quadrigarum super capita montium exilient sicut sonitus flammae ignis devorantis stipulam velut populus fortis praeparatus ad proelium
JOEL|2|6|a facie eius cruciabuntur populi omnes vultus redigentur in ollam
JOEL|2|7|sicut fortes current quasi viri bellatores ascendent murum vir in viis suis gradietur et non declinabunt a semitis suis
JOEL|2|8|unusquisque fratrem suum non coartabit singuli in calle suo ambulabunt sed et per fenestras cadent et non demolientur
JOEL|2|9|urbem ingredientur in muro current domos conscendent per fenestras intrabunt quasi fur
JOEL|2|10|a facie eius contremuit terra moti sunt caeli sol et luna obtenebrati sunt et stellae retraxerunt splendorem suum
JOEL|2|11|et Dominus dedit vocem suam ante faciem exercitus sui quia multa sunt nimis castra eius quia fortia et facientia verbum eius magnus enim dies Domini et terribilis valde et quis sustinebit eum
JOEL|2|12|nunc ergo dicit Dominus convertimini ad me in toto corde vestro in ieiunio et in fletu et in planctu
JOEL|2|13|et scindite corda vestra et non vestimenta vestra et convertimini ad Dominum Deum vestrum quia benignus et misericors est patiens et multae misericordiae et praestabilis super malitia
JOEL|2|14|quis scit si convertatur et ignoscat et relinquat post se benedictionem sacrificium et libamen Domino Deo nostro
JOEL|2|15|canite tuba in Sion sanctificate ieiunium vocate coetum
JOEL|2|16|congregate populum sanctificate ecclesiam coadunate senes congregate parvulos et sugentes ubera egrediatur sponsus de cubili suo et sponsa de thalamo suo
JOEL|2|17|inter vestibulum et altare plorabunt sacerdotes ministri Domini et dicent parce Domine populo tuo et ne des hereditatem tuam in obprobrium ut dominentur eis nationes quare dicunt in populis ubi est Deus eorum
JOEL|2|18|zelatus est Dominus terram suam et pepercit populo suo
JOEL|2|19|et respondit Dominus et dixit populo suo ecce ego mittam vobis frumentum et vinum et oleum et replebimini eo et non dabo vos ultra obprobrium in gentibus
JOEL|2|20|et eum qui ab aquilone est procul faciam a vobis et expellam eum in terram inviam et desertam faciem eius contra mare orientale et extremum eius ad mare novissimum et ascendet fetor eius et ascendet putredo eius quia superbe egit
JOEL|2|21|noli timere terra exulta et laetare quoniam magnificavit Dominus ut faceret
JOEL|2|22|nolite timere animalia regionis quia germinaverunt speciosa deserti quia lignum adtulit fructum suum ficus et vinea dederunt virtutem suam
JOEL|2|23|et filii Sion exultate et laetamini in Domino Deo vestro quia dedit vobis doctorem iustitiae et descendere faciet ad vos imbrem matutinum et serotinum in principio
JOEL|2|24|et implebuntur areae frumento et redundabunt torcularia vino et oleo
JOEL|2|25|et reddam vobis annos quos comedit lucusta bruchus et rubigo et eruca fortitudo mea magna quam misi in vos
JOEL|2|26|et comedetis vescentes et saturabimini et laudabitis nomen Domini Dei vestri qui fecit vobiscum mirabilia et non confundetur populus meus in sempiternum
JOEL|2|27|et scietis quia in medio Israhel ego sum et ego Dominus Deus vester et non est amplius et non confundetur populus meus in aeternum
JOEL|2|28|et erit post haec effundam spiritum meum super omnem carnem et prophetabunt filii vestri et filiae vestrae senes vestri somnia somniabunt et iuvenes vestri visiones videbunt
JOEL|2|29|sed et super servos et ancillas in diebus illis effundam spiritum meum
JOEL|2|30|et dabo prodigia in caelo et in terra sanguinem et ignem et vaporem fumi
JOEL|2|31|sol vertetur in tenebras et luna in sanguinem antequam veniat dies Domini magnus et horribilis
JOEL|2|32|et erit omnis qui invocaverit nomen Domini salvus erit quia in monte Sion et in Hierusalem erit salvatio sicut dixit Dominus et in residuis quos Dominus vocaverit
JOEL|3|1|quia ecce in diebus illis et in tempore illo cum convertero captivitatem Iuda et Hierusalem
JOEL|3|2|congregabo omnes gentes et deducam eas in valle Iosaphat et disceptabo cum eis ibi super populo meo et hereditate mea Israhel quos disperserunt in nationibus et terram meam diviserunt
JOEL|3|3|et super populum meum miserunt sortem et posuerunt puerum in prostibulum et puellam vendiderunt pro vino ut biberent
JOEL|3|4|verum quid vobis et mihi Tyrus et Sidon et omnis terminus Palestinorum numquid ultionem vos redditis mihi et si ulciscimini vos contra me cito velociter reddam vicissitudinem vobis super caput vestrum
JOEL|3|5|argentum enim meum et aurum tulistis et desiderabilia mea et pulcherrima intulistis in delubra vestra
JOEL|3|6|et filios Iuda et filios Hierusalem vendidistis filiis Graecorum ut longe faceretis eos de finibus suis
JOEL|3|7|ecce ego suscitabo eos de loco in quo vendidistis eos et convertam retributionem vestram in caput vestrum
JOEL|3|8|et vendam filios vestros et filias vestras in manibus filiorum Iuda et venundabunt eos Sabeis genti longinquae quia Dominus locutus est
JOEL|3|9|clamate hoc in gentibus sanctificate bellum suscitate robustos accedant ascendant omnes viri bellatores
JOEL|3|10|concidite aratra vestra in gladios et ligones vestros in lanceas infirmus dicat quia fortis ego sum
JOEL|3|11|erumpite et venite omnes gentes de circuitu et congregamini ibi occumbere faciet Dominus robustos tuos
JOEL|3|12|consurgant et ascendant gentes in vallem Iosaphat quia ibi sedebo ut iudicem omnes gentes in circuitu
JOEL|3|13|mittite falces quoniam maturavit messis venite et descendite quia plenum est torcular exuberant torcularia quia multiplicata est malitia eorum
JOEL|3|14|populi populi in valle concisionis quia iuxta est dies Domini in valle concisionis
JOEL|3|15|sol et luna obtenebricata sunt et stellae retraxerunt splendorem suum
JOEL|3|16|et Dominus de Sion rugiet et de Hierusalem dabit vocem suam et movebuntur caeli et terra et Dominus spes populi sui et fortitudo filiorum Israhel
JOEL|3|17|et scietis quia ego Dominus Deus vester habitans in Sion in monte sancto meo et erit Hierusalem sancta et alieni non transibunt per eam amplius
JOEL|3|18|et erit in die illa stillabunt montes dulcedinem et colles fluent lacte et per omnes rivos Iuda ibunt aquae et fons de domo Domini egredietur et inrigabit torrentem Spinarum
JOEL|3|19|Aegyptus in desolatione erit et Idumea in desertum perditionis pro eo quod inique egerint in filios Iuda et effuderint sanguinem innocentem in terra sua
JOEL|3|20|et Iudaea in aeternum habitabitur et Hierusalem in generatione et generationem
JOEL|3|21|et mundabo sanguinem eorum quem non mundaveram et Dominus commorabitur in Sion
