JONAH|1|1|И было слово Господне к Ионе, сыну Амафиину:
JONAH|1|2|встань, иди в Ниневию, город великий, и проповедуй в нем, ибо злодеяния его дошли до Меня.
JONAH|1|3|И встал Иона, чтобы бежать в Фарсис от лица Господня, и пришел в Иоппию, и нашел корабль, отправлявшийся в Фарсис, отдал плату за провоз и вошел в него, чтобы плыть с ними в Фарсис от лица Господа.
JONAH|1|4|Но Господь воздвиг на море крепкий ветер, и сделалась на море великая буря, и корабль готов был разбиться.
JONAH|1|5|И устрашились корабельщики, и взывали каждый к своему богу, и стали бросать в море кладь с корабля, чтобы облегчить его от нее; Иона же спустился во внутренность корабля, лег и крепко заснул.
JONAH|1|6|И пришел к нему начальник корабля и сказал ему: что ты спишь? встань, воззови к Богу твоему; может быть, Бог вспомнит о нас и мы не погибнем.
JONAH|1|7|И сказали друг другу: пойдем, бросим жребии, чтобы узнать, за кого постигает нас эта беда. И бросили жребии, и пал жребий на Иону.
JONAH|1|8|Тогда сказали ему: скажи нам, за кого постигла нас эта беда? какое твое занятие, и откуда идешь ты? где твоя страна, и из какого ты народа?
JONAH|1|9|И он сказал им: я Еврей, чту Господа Бога небес, сотворившего море и сушу.
JONAH|1|10|И устрашились люди страхом великим и сказали ему: для чего ты это сделал? Ибо узнали эти люди, что он бежит от лица Господня, как он сам объявил им.
JONAH|1|11|И сказали ему: что сделать нам с тобою, чтобы море утихло для нас? Ибо море не переставало волноваться.
JONAH|1|12|Тогда он сказал им: возьмите меня и бросьте меня в море, и море утихнет для вас, ибо я знаю, что ради меня постигла вас эта великая буря.
JONAH|1|13|Но эти люди начали усиленно грести, чтобы пристать к земле, но не могли, потому что море все продолжало бушевать против них.
JONAH|1|14|Тогда воззвали они к Господу и сказали: молим Тебя, Господи, да не погибнем за душу человека сего, и да не вменишь нам кровь невинную; ибо Ты, Господи, соделал, что угодно Тебе!
JONAH|1|15|И взяли Иону и бросили его в море, и утихло море от ярости своей.
JONAH|1|16|И устрашились эти люди Господа великим страхом, и принесли Господу жертву, и дали обеты.
JONAH|2|1|И повелел Господь большому киту поглотить Иону; и был Иона во чреве этого кита три дня и три ночи.
JONAH|2|2|И помолился Иона Господу Богу своему из чрева кита
JONAH|2|3|и сказал: к Господу воззвал я в скорби моей, и Он услышал меня; из чрева преисподней я возопил, и Ты услышал голос мой.
JONAH|2|4|Ты вверг меня в глубину, в сердце моря, и потоки окружили меня, все воды Твои и волны Твои проходили надо мною.
JONAH|2|5|И я сказал: отринут я от очей Твоих, однако я опять увижу святый храм Твой.
JONAH|2|6|Объяли меня воды до души моей, бездна заключила меня; морскою травою обвита была голова моя.
JONAH|2|7|До основания гор я нисшел, земля своими запорами навек заградила меня; но Ты, Господи Боже мой, изведешь душу мою из ада.
JONAH|2|8|Когда изнемогла во мне душа моя, я вспомнил о Господе, и молитва моя дошла до Тебя, до храма святаго Твоего.
JONAH|2|9|Чтущие суетных и ложных [богов] оставили Милосердаго своего,
JONAH|2|10|а я гласом хвалы принесу Тебе жертву; что обещал, исполню: у Господа спасение!
JONAH|2|11|И сказал Господь киту, и он изверг Иону на сушу.
JONAH|3|1|И было слово Господне к Ионе вторично:
JONAH|3|2|встань, иди в Ниневию, город великий, и проповедуй в ней, что Я повелел тебе.
JONAH|3|3|И встал Иона и пошел в Ниневию, по слову Господню; Ниневия же была город великий у Бога, на три дня ходьбы.
JONAH|3|4|И начал Иона ходить по городу, сколько можно пройти в один день, и проповедывал, говоря: еще сорок дней и Ниневия будет разрушена!
JONAH|3|5|И поверили Ниневитяне Богу, и объявили пост, и оделись во вретища, от большого из них до малого.
JONAH|3|6|Это слово дошло до царя Ниневии, и он встал с престола своего, и снял с себя царское облачение свое, и оделся во вретище, и сел на пепле,
JONAH|3|7|и повелел провозгласить и сказать в Ниневии от имени царя и вельмож его: "чтобы ни люди, ни скот, ни волы, ни овцы ничего не ели, не ходили на пастбище и воды не пили,
JONAH|3|8|и чтобы покрыты были вретищем люди и скот и крепко вопияли к Богу, и чтобы каждый обратился от злого пути своего и от насилия рук своих.
JONAH|3|9|Кто знает, может быть, еще Бог умилосердится и отвратит от нас пылающий гнев Свой, и мы не погибнем".
JONAH|3|10|И увидел Бог дела их, что они обратились от злого пути своего, и пожалел Бог о бедствии, о котором сказал, что наведет на них, и не навел.
JONAH|4|1|Иона сильно огорчился этим и был раздражен.
JONAH|4|2|И молился он Господу и сказал: о, Господи! не это ли говорил я, когда еще был в стране моей? Потому я и побежал в Фарсис, ибо знал, что Ты Бог благий и милосердый, долготерпеливый и многомилостивый и сожалеешь о бедствии.
JONAH|4|3|И ныне, Господи, возьми душу мою от меня, ибо лучше мне умереть, нежели жить.
JONAH|4|4|И сказал Господь: неужели это огорчило тебя так сильно?
JONAH|4|5|И вышел Иона из города, и сел с восточной стороны у города, и сделал себе там кущу, и сел под нею в тени, чтобы увидеть, что будет с городом.
JONAH|4|6|И произрастил Господь Бог растение, и оно поднялось над Ионою, чтобы над головою его была тень и чтобы избавить его от огорчения его; Иона весьма обрадовался этому растению.
JONAH|4|7|И устроил Бог так, что на другой день при появлении зари червь подточил растение, и оно засохло.
JONAH|4|8|Когда же взошло солнце, навел Бог знойный восточный ветер, и солнце стало палить голову Ионы, так что он изнемог и просил себе смерти, и сказал: лучше мне умереть, нежели жить.
JONAH|4|9|И сказал Бог Ионе: неужели так сильно огорчился ты за растение? Он сказал: очень огорчился, даже до смерти.
JONAH|4|10|Тогда сказал Господь: ты сожалеешь о растении, над которым ты не трудился и которого не растил, которое в одну ночь выросло и в одну же ночь и пропало:
JONAH|4|11|Мне ли не пожалеть Ниневии, города великого, в котором более ста двадцати тысяч человек, не умеющих отличить правой руки от левой, и множество скота?
