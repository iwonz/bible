2CHR|1|1|Confortatus est ergo Salomon filius David in regno suo, et Dominus Deus eius erat cum eo et magnificavit eum in excelsum.
2CHR|1|2|Praecepitque Salomon universo Israeli, tribunis et centurionibus et iudicibus et ducibus omnis Israel et principibus familiarum
2CHR|1|3|et abiit cum universa multitudine in excelsum Gabaon, ubi erat tabernaculum conventus Dei, quod fecit Moyses famulus Dei in solitudine.
2CHR|1|4|Arcam autem Dei adduxerat David de Cariathiarim in locum, quem praeparaverat ei et ubi fixerat illi tabernaculum, hoc est in Ierusalem;
2CHR|1|5|altare quoque aeneum, quod fabricatus fuerat Beseleel filius Uri filii Hur, ibi erat coram tabernaculo Domini; ibique requisivit eum Salomon et omnis ecclesia.
2CHR|1|6|Ascenditque ibi Salomon ad altare aeneum coram tabernaculo conventus Domini et obtulit in eo mille hostias.
2CHR|1|7|Ecce autem in ipsa nocte apparuit ei Deus dicens: " Postula, quod vis, ut dem tibi ".
2CHR|1|8|Dixitque Salomon Deo: " Tu fecisti cum David patre meo misericordiam magnam et constituisti me regem pro eo.
2CHR|1|9|Nunc ergo, Domine Deus, impleatur sermo tuus, quem pollicitus es David patri meo; tu enim me fecisti regem super populum tuum multum, qui tam innumerabilis est quam pulvis terrae.
2CHR|1|10|Da mihi sapientiam et intellegentiam, ut ingrediar et egrediar coram populo tuo; quis enim potest hunc populum tuum digne, qui tam grandis est, iudicare? ".
2CHR|1|11|Dixit autem Deus ad Salomonem: " Quia hoc magis placuit cordi tuo et non postulasti divitias et substantiam et gloriam neque animas eorum, qui te oderant, sed nec dies vitae plurimos, petisti autem sapientiam et scientiam, ut iudicare possis populum meum, super quem constitui te regem,
2CHR|1|12|sapientia et scientia data sunt tibi; divitias autem et substantiam et gloriam dabo tibi, ita ut nullus in regibus nec ante te nec post te fuerit similis tui ".
2CHR|1|13|Venit ergo Salomon ab excelso Gabaon in Ierusalem coram tabernaculo conventus et regnavit super Israel.
2CHR|1|14|Congregavitque sibi currus et equites, et facti sunt ei mille quadringenti currus et duodecim milia equitum, et fecit eos esse in urbibus quadrigarum et cum rege in Ierusalem.
2CHR|1|15|Praebuitque rex argentum et aurum in Ierusalem quasi lapides et cedros quasi sycomoros, quae nascuntur in Sephela multitudine magna.
2CHR|1|16|Adducebantur autem ei equi de Aegypto et de Coa; negotiatores regis de Coa emebant pretio
2CHR|1|17|et faciebant ascendere et exire de Aegypto quadrigam sescentis argenteis et equum centum quinquaginta; similiter universis regibus Hetthaeorum et Syriae per manus suas educebant.
2CHR|1|18|Decrevit autem Salomon aedificare domum nomini Domini et palatium sibi.
2CHR|2|1|Et numeravit septuaginta milia virorum portantium umeris et octoginta milia, qui caederent lapides in montibus, praepositosque eorum tria milia sescentos.
2CHR|2|2|Misit quoque ad Hiram regem Tyri dicens: " Sicut egisti cum David patre meo et misisti ei ligna cedrina, ut aedificaret sibi domum ad habitandum in ea,
2CHR|2|3|sic fac mecum, ut aedificem domum nomini Domini Dei mei, ut consecrem eam ad adolendum coram illo fumiganda aromata et ad propositionem panum sempiternam et ad holocautomata mane et vespere, sabbatis quoque et neomeniis et sollemnitatibus Domini Dei nostri in sempiternum, quae mandata sunt Israeli.
2CHR|2|4|Domus enim, quam aedificare cupio, magna est; magnus est enim Deus noster super omnes deos.
2CHR|2|5|Quis ergo poterit praevalere, ut aedificet ei dignam domum? Si caelum et caeli caelorum capere eum nequeunt, quantus ego sum, ut possim aedificare ei domum? Sed ad hoc tantum, ut adoleatur incensum coram illo.
2CHR|2|6|Mitte ergo mihi virum eruditum, qui noverit operari in auro et argento, aere et ferro, purpura, coccino et hyacintho, et qui sciat sculpere caelaturas cum his artificibus, quos mecum habeo in Iudaea et Ierusalem, quos praeparavit David pater meus.
2CHR|2|7|Sed et ligna cedrina mitte mihi et arceuthina et pinea de Libano; scio enim quod servi tui noverint caedere ligna de Libano, et erunt servi mei cum servis tuis,
2CHR|2|8|ut parentur mihi ligna plurima; domus enim, quam cupio aedificare, magna erit nimis et inclita.
2CHR|2|9|Praeterea operariis, qui caesuri sunt ligna, servis tuis dabo in cibaria tritici choros viginti milia et hordei choros totidem et vini viginti milia batos, olei quoque batos viginti milia ".
2CHR|2|10|Dixit autem Hiram rex Tyri per litteras, quas miserat Salomoni: " Quia dilexit Dominus populum suum, idcirco te regnare fecit super eum ".
2CHR|2|11|Et addidit dicens: " Benedictus Dominus, Deus Israel, qui fecit caelum et terram, qui dedit David regi filium sapientem et eruditum et sensatum atque prudentem, ut aedificaret domum Domino et palatium sibi.
2CHR|2|12|Misi ergo tibi virum prudentem et scientissimum Hiram magistrum meum,
2CHR|2|13|filium mulieris de filiabus Dan, cuius pater fuit Tyrius, qui novit operari in auro et argento, aere et ferro et lapidibus et lignis, in purpura quoque et hyacintho et bysso et coccino, et qui scit caelare omnem sculpturam et adinvenire prudenter, quodcumque in opere necessarium est, cum artificibus tuis et cum artificibus domini mei David patris tui.
2CHR|2|14|Triticum ergo et hordeum et oleum et vinum, quae pollicitus es, domine mi, mitte servis tuis.
2CHR|2|15|Nos autem caedemus ligna de Libano, quot necessaria habueris, et applicabimus ea ratibus per mare in Ioppe; tuum autem erit transferre ea in Ierusalem ".
2CHR|2|16|Numeravit igitur Salomon omnes viros peregrinos, qui erant in terra Israel post dinumerationem, quam dinumeravit David pater eius; et inventi sunt centum quinquaginta milia et tria milia sescenti.
2CHR|2|17|Fecitque ex eis septuaginta milia, qui umeris onera portarent, et octoginta milia, qui lapides in montibus caederent; tria autem milia et sescentos praepositos operum populi.
2CHR|3|1|Et coepit Salomon aedificare domum Domini in Ierusalem in monte Moria, qui demonstratus fuerat a David patre eius, in loco, quem paraverat David in area Ornan Iebusaei.
2CHR|3|2|Coepit autem aedificare mense secundo anno quarto regni sui.
2CHR|3|3|Et hae sunt mensurae, quas statuit Salomon, ut aedificaret domum Dei: longitudinis cubiti in mensura prima sexaginta, latitudinis cubiti viginti.
2CHR|3|4|Porticum vero ante frontem, quae tendebatur in longum, iuxta mensuram latitudinis domus, cubitorum viginti; porro altitudo centum viginti cubitorum erat. Et deauravit eam intrinsecus auro mundissimo.
2CHR|3|5|Domum quoque maiorem texit tabulis ligneis abiegnis et laminas auri obryzi affixit per totum; scalpsitque in eis palmas et quasi catenulas se invicem complectentes.
2CHR|3|6|Stravit quoque pavimentum templi pretiosissimo marmore decore multo.
2CHR|3|7|Porro aurum erat de Parvaim, de cuius laminis texit domum, et trabes eius et postes et parietes et ostia; et caelavit cherubim in parietibus.
2CHR|3|8|Fecit quoque domum sancti sanctorum: longitudinem iuxta latitudinem domus cubitorum viginti et latitudinem similiter viginti cubitorum; et laminis auri optimi texit eam quasi talentis sescentis.
2CHR|3|9|Sed et pro clavis usus est auro ponderis quinquaginta siclorum. Cenacula quoque texit auro.
2CHR|3|10|Fecit etiam in domo sancti sanctorum cherubim duos opere statuario et texit eos auro.
2CHR|3|11|Alae cherubim viginti cubitis extendebantur, ita ut una ala haberet cubitos quinque et tangeret parietem domus, et altera quinque cubitos habens alam tangeret alterius cherub.
2CHR|3|12|Similiter cherub alterius ala quinque habebat cubitos et tangebat parietem, et ala eius altera quinque cubitorum alam cherub alterius contingebat.
2CHR|3|13|Igitur alae utriusque cherubim expansae erant et extendebantur per cubitos viginti; ipsi autem stabant erectis pedibus, et facies eorum erant versae ad exteriorem domum.
2CHR|3|14|Fecit quoque velum ex hyacintho, purpura, cocco et bysso et intexuit ei cherubim.
2CHR|3|15|Ante fores etiam templi duas columnas, quae triginta et quinque cubitos habebant altitudinis; porro capita earum quinque cubitorum.
2CHR|3|16|Necnon et quasi catenulas in torque, et superposuit eas capitibus columnarum; malogranata etiam centum, quae catenulis interposuit.
2CHR|3|17|Ipsas quoque columnas posuit ante faciem templi, unam a dextris et alteram a sinistris; eam, quae a dextris erat, vocavit Iachin et, quae ad laevam, Booz.
2CHR|4|1|Fecit quoque altare aeneum viginti cubitorum longitudinis et viginti cubitorum latitudinis et decem cubitorum
2CHR|4|2|altitudinis. Mare etiam fusile decem cubitis a labio usque ad labium rotundum per circuitum; quinque cubitos habebat altitudinis, et funiculus triginta cubitorum ambiebat gyrum eius.
2CHR|4|3|Similitudo quoque boum erat subter illud, in circuitu circumdabant illud decem cubitis - duobus versibus alvum maris circuibant boves fusiles in una fusione cum mari.
2CHR|4|4|Et ipsum mare super duodecim boves impositum erat, quorum tres respiciebant aquilonem et alii tres occidentem, porro tres alii meridiem et tres, qui reliqui erant, orientem habentes mare superpositum; posteriora autem boum erant intrinsecus sub mari.
2CHR|4|5|Porro vastitas eius habebat mensuram palmi, et labium illius erat quasi labium calicis vel repandi lilii; capiebatque tria milia batos.
2CHR|4|6|Fecit quoque luteres decem et posuit quinque a dextris et quinque a sinistris, ut lavarent in eis omnia, quae in holocaustum oblaturi erant; porro in mari sacerdotes lavabantur.
2CHR|4|7|Fecit autem et candelabra aurea decem secundum speciem, qua iussa erant fieri, et posuit ea in templo quinque a dextris et quinque a sinistris.
2CHR|4|8|Necnon et mensas decem, et posuit eas in templo quinque a dextris et quinque a sinistris; phialas quoque aureas centum.
2CHR|4|9|Fecit etiam atrium sacerdotum et atrium grande et ostia in atrio, quae texit aere.
2CHR|4|10|Porro mare posuit in latere dextro contra orientem ad meridiem.
2CHR|4|11|Fecit autem Hiram lebetes et vatilla et phialas et complevit omne opus regis Salomonis in domo Dei;
2CHR|4|12|hoc est columnas duas et globos et capitella super caput columnarum duarum et serta duo, quae tegerent globos capitellorum;
2CHR|4|13|malogranata quoque quadringenta et serta duo, ita ut bini ordines malogranatorum singulis sertis iungerentur, quae protegerent globos capitellorum columnarum.
2CHR|4|14|Bases etiam fecit et luteres, quos superposuit basibus,
2CHR|4|15|mare unum, boves quoque duodecim sub mari;
2CHR|4|16|et lebetes et vatilla et fuscinulas: omnia vasa fecit regi Salomoni Hiram magister eius pro domo Domini ex aere mundissimo.
2CHR|4|17|In regione Iordanis fudit ea rex in argillosa terra inter Succoth et Saredatha.
2CHR|4|18|Fecitque Salomon multitudinem vasorum innumerabilem, ita ut ignoraretur pondus aeris.
2CHR|4|19|Fecitque Salomon omnia vasa domus Dei et altare aureum et mensas et super eas panes propositionis;
2CHR|4|20|candelabra quoque cum lucernis suis, ut lucerent ante Dabir iuxta ritum, ex auro purissimo,
2CHR|4|21|et florem et lucernas et forcipes aureos: omnia de auro perfectissimo facta sunt;
2CHR|4|22|cultros quoque et phialas et sartagines et turibula ex auro purissimo. Et ostia templi interiora in sancta sanctorum et ostia templi forinsecus aurea.
2CHR|5|1|Sicque completum est omne opus, quod fecit Salomon in do mo Domini. Intulit igitur Salomon omnia, quae voverat David pater suus, argentum et aurum, et universa vasa posuit in thesauris domus Dei.
2CHR|5|2|Post quae congregavit maiores natu Israel et cunctos principes tribuum et capita familiarum de filiis Israel in Ierusalem, ut adducerent arcam foederis Domini de civitate David, quae est Sion.
2CHR|5|3|Venerunt igitur ad regem omnes viri Israel in die sollemni mensis septimi.
2CHR|5|4|Cumque venissent cuncti seniorum Israel, portaverunt Levitae arcam
2CHR|5|5|et intulerunt eam et tabernaculum conventus et omnem paraturam tabernaculi. Porro omnia vasa sanctuarii, quae erant in tabernaculo, portaverunt sacerdotes levitici generis.
2CHR|5|6|Rex autem Salomon et universus coetus Israel, omnes, qui fuerunt congregati ad eum ante arcam, immolabant oves et boves absque ullo numero: tanta enim erat multitudo victimarum.
2CHR|5|7|Et intulerunt sacerdotes arcam foederis Domini in locum suum ad Dabir templi, in sancta sanctorum subter alas cherubim,
2CHR|5|8|ita ut cherubim expanderent alas suas super locum, in quo posita erat arca, et ipsam arcam tegerent cum vectibus suis ab alto.
2CHR|5|9|Vectium autem, quibus portabatur arca, quia paululum longiores erant, capita parebant ante Dabir; si vero quis erat extrinsecus eos videre non poterat. Fuit itaque arca ibi usque in praesentem diem.
2CHR|5|10|Nihilque erat aliud in arca, nisi duae tabulae, quas posuerat Moyses in Horeb, quando fecit Dominus foedus cum filiis Israel egredientibus ex Aegypto.
2CHR|5|11|Egressis autem sacerdotibus de sanctuario - omnes enim sacerdotes, qui ibi potuerant inveniri, sanctificati sunt, non observantes vices et ministeriorum ordinem,
2CHR|5|12|et Levitae cantores, omnes, qui sub Asaph erant et qui sub Heman et qui sub Idithun, filii et fratres eorum, vestiti byssinis, cymbalis et psalteriis et citharis stabant ad orientalem plagam altaris, et cum eis sacerdotes centum viginti canentes tubis -
2CHR|5|13|igitur cunctis pariter et tubis et voce et cymbalis et organis et diversi generis musicorum concinentibus et vocem in sublime tollentibus, cum una voce Dominum laudare coepissent et dicere: " Confitemini Domino quoniam bonus, quoniam in aeternum misericordia eius ", impleta est domus Dei nube,
2CHR|5|14|nec potuerunt sacerdotes stare et ministrare propter nubem; compleverat enim gloria Domini domum Dei.
2CHR|6|1|Tunc Salomon ait: " Dominus pollicitus est, ut habitaret in ca ligine;
2CHR|6|2|ego autem aedificavi domum in habitaculum tuum, ut habitares ibi in perpetuum ".
2CHR|6|3|Et convertit rex faciem suam et benedixit universae multitudini Israel - nam omnis turba stabat intenta - et ait:
2CHR|6|4|" Benedictus Dominus, Deus Israel, qui, quod locutus est ore suo David patri meo, opere complevit dicens:
2CHR|6|5|"A die qua eduxi populum meum de terra Aegypti non elegi civitatem de cunctis tribubus Israel, ut aedificaretur in ea domus nomini meo, neque elegi quemquam alium virum, ut esset dux in populo meo Israel,
2CHR|6|6|sed elegi Ierusalem, ut sit nomen meum in ea, et elegi David, ut constituerem eum super populum meum Israel".
2CHR|6|7|Cumque fuisset voluntatis David patris mei, ut aedificaret domum nomini Domini, Dei Israel,
2CHR|6|8|dixit Dominus ad eum: "Quia haec fuit voluntas tua, ut aedificares domum nomini meo, bene quidem fecisti huiuscemodi habere voluntatem,
2CHR|6|9|sed non tu aedificabis domum, verum filius tuus, qui egredietur de lumbis tuis, ipse aedificabit domum nomini meo".
2CHR|6|10|Complevit ergo Dominus sermonem suum, quem locutus fuerat, et ego surrexi pro David patre meo et sedi super thronum Israel, sicut locutus est Dominus, et aedificavi domum nomini Domini, Dei Israel;
2CHR|6|11|et posui in ea arcam, in qua est pactum Domini, quod pepigit cum filiis Israel ".
2CHR|6|12|Stetit ergo coram altari Domini ex adverso universae multitudinis Israel et extendit manus suas.
2CHR|6|13|Siquidem fecerat Salomon basim aeneam et posuerat eam in medio atrii habentem quinque cubitos longitudinis et quinque cubitos latitudinis et tres cubitos altitudinis, stetitque super eam; et deinceps, flexis genibus contra universam multitudinem Israel et palmis in caelum levatis,
2CHR|6|14|ait: " Domine, Deus Israel, non est similis tui Deus in caelo et in terra, qui custodis pactum et misericordiam cum servis tuis, qui ambulant coram te in toto corde suo,
2CHR|6|15|qui praestitisti servo tuo David patri meo quaecumque locutus fueras ei, et, quae ore promiseras, opere complesti, sicut et praesens tempus probat.
2CHR|6|16|Nunc ergo, Domine, Deus Israel, imple servo tuo patri meo David, quaecumque locutus es dicens: "Non deficiet ex te vir coram me, qui sedeat super thronum Israel, ita tamen si custodierint filii tui vias suas et ambulaverint in lege mea, sicut et tu ambulasti coram me".
2CHR|6|17|Et nunc, Domine, Deus Israel, firmetur sermo tuus, quem locutus es servo tuo David!
2CHR|6|18|Ergone credibile est, ut habitet Deus cum hominibus super terram? Si caelum et caeli caelorum non te capiunt, quanto magis domus ista, quam aedificavi!
2CHR|6|19|Sed respice orationem servi tui et obsecrationem eius, Domine Deus meus, et audi clamorem et preces, quas fundit famulus tuus coram te,
2CHR|6|20|ut aperias oculos tuos super domum istam diebus ac noctibus, super locum in quo pollicitus es, ut ponas nomen tuum et exaudires orationem, quam servus tuus orat in eo.
2CHR|6|21|Et exaudi preces famuli tui et populi tui Israel, qui oraverint ad locum istum; exaudi de habitaculo tuo, de caelis, exaudi et propitiare!
2CHR|6|22|Si peccaverit quispiam in proximum suum, et ille exegerit ab eo iuramentum, ut se maledicto constringat coram altari in domo ista,
2CHR|6|23|tu audies de caelo et facies iudicium servorum tuorum, ita ut reddas iniquo viam suam in caput proprium et ulciscaris iustum retribuens ei secundum iustitiam suam.
2CHR|6|24|Si superatus fuerit populus tuus Israel ab inimicis, quia peccaturi sunt tibi, et conversi egerint paenitentiam et confitentes nomini tuo oraverint et fuerint deprecati in domo ista,
2CHR|6|25|tu exaudies de caelo, et propitiare peccato populi tui Israel et reduc eos in terram, quam dedisti eis et patribus eorum.
2CHR|6|26|Si clauso caelo pluvia non fluxerit propter peccata populi, et deprecati te fuerint in loco isto et confessi nomini tuo et conversi a peccatis suis, cum eos afflixeris,
2CHR|6|27|exaudi de caelo, Domine, et dimitte peccata servorum tuorum et populi tui Israel, doce eos viam bonam, per quam ingrediantur, et da pluviam terrae, quam dedisti populo tuo ad possidendum.
2CHR|6|28|Fames si orta fuerit in terra et pestilentia, uredo et aurugo et locusta et bruchus et hostes, vastatis regionibus, portas eius obsederint, omnisque plaga et infirmitas presserit,
2CHR|6|29|si quis de populo tuo Israel fuerit deprecatus cognoscens plagam et infirmitatem suam et expanderit manus suas ad domum hanc,
2CHR|6|30|tu exaudi de caelo, de loco habitationis tuae, et propitiare et redde unicuique secundum vias suas, quia nosti cor eius; tu enim solus nosti corda filiorum hominum,
2CHR|6|31|ut timeant te et ambulent in viis tuis cunctis diebus, quibus vivunt super faciem terrae, quam dedisti patribus nostris.
2CHR|6|32|Externum quoque, qui non est de populo tuo Israel, si venerit de terra longinqua propter nomen tuum magnum et propter manum tuam robustam et brachium tuum extentum, et oraverit in loco isto,
2CHR|6|33|tu exaudies de caelo firmissimo habitaculo tuo et facies cuncta, pro quibus invocaverit te ille peregrinus, ut sciant omnes populi terrae nomen tuum et timeant te sicut populus tuus Israel et cognoscant quia nomen tuum invocatum est super domum hanc, quam aedificavi.
2CHR|6|34|Si egressus fuerit populus tuus ad bellum contra adversarios suos per viam, in qua miseris eos, et oraverint te contra viam, in qua civitas haec est, quam elegisti, et domus, quam aedificavi nomini tuo,
2CHR|6|35|tu exaudies de caelo preces eorum et obsecrationem, et facies iudicium eorum.
2CHR|6|36|Si autem peccaverint tibi - neque enim est homo, qui non peccet - et iratus fueris eis et tradideris hostibus, et captivos duxerint eos in terram longinquam vel propinquam,
2CHR|6|37|et conversi in corde suo in terra, ad quam captivi ducti fuerant, egerint paenitentiam et deprecati te fuerint in terra captivitatis suae dicentes: "Peccavimus, inique fecimus, iniuste egimus";
2CHR|6|38|et reversi fuerint ad te in toto corde suo et in tota anima sua in terra captivitatis suae, ad quam ducti sunt, et oraverint te contra viam terrae suae, quam dedisti patribus eorum, et urbis, quam elegisti, et domus, quam aedificavi nomini tuo,
2CHR|6|39|ut exaudias de caelo, de loco habitationis tuae, preces eorum et supplicationes eorum et facias iudicium et dimittas populo tuo, qui peccavit tibi;
2CHR|6|40|tu es enim Deus meus. Aperiantur, quaeso, oculi tui, et aures tuae intentae sint ad orationem, quae fit in loco isto.
2CHR|6|41|Nunc igitur consurge, Domine Deus, in requiem tuam, tu et arca fortitudinis tuae; sacerdotes tui, Domine Deus, induantur salutem, et sancti tui laetentur in bonis.
2CHR|6|42|Domine Deus, ne averteris faciem christi tui; memento misericordiarum David servi tui ".
2CHR|7|1|Cumque complesset Salomon fundens preces, ignis descendit de caelo et devoravit holocaustum et victimas, et maiestas Domini implevit domum.
2CHR|7|2|Nec poterant sacerdotes ingredi templum Domini, eo quod implesset maiestas Domini templum Domini.
2CHR|7|3|Sed et omnes filii Israel videbant descendentem ignem et gloriam Domini super domum et corruentes proni in terram super pavimentum stratum lapide adoraverunt et laudaverunt Dominum: " Quoniam bonus, quoniam in saeculum misericordia eius ".
2CHR|7|4|Rex autem et omnis populus immolabant victimas coram Domino.
2CHR|7|5|Mactavit igitur rex Salomon hostias boum viginti duo milia, ovium centum viginti milia, et dedicavit domum Dei rex et universus populus.
2CHR|7|6|Sacerdotes autem stabant in officiis suis et Levitae in organis carminum Domini, quae fecit David rex ad laudandum Dominum: " Quoniam in aeternum misericordia eius ", hymnos David canentes per manus suas. Porro sacerdotes canebant tubis ante eos, cunctusque Israel stabat.
2CHR|7|7|Sanctificavit quoque Salomon medium atrii ante templum Domini; obtulerat enim ibi holocausta et adipes pacificorum, quia altare aeneum, quod fecerat, non poterat sustinere holocausta et oblationes et adipes.
2CHR|7|8|Fecit ergo Salomon sollemnitatem in tempore illo septem diebus, et omnis Israel cum eo, ecclesia magna valde ab introitu Emath usque ad torrentem Aegypti.
2CHR|7|9|Feceruntque die octavo collectam magnam, eo quod dedicassent altare septem diebus et sollemnitatem celebrassent diebus septem.
2CHR|7|10|Igitur in die vicesimo tertio mensis septimi dimisit populum ad tabernacula sua, laetantem atque gaudentem super bono, quod fecerat Dominus Davidi et Salomoni et Israeli populo suo.
2CHR|7|11|Complevitque Salomon domum Domini et domum regis; et in omnibus, quae disposuerat in corde suo, ut faceret in domo Domini et in domo sua, prosperatus est.
2CHR|7|12|Apparuit autem ei Dominus nocte et ait: " Audivi orationem tuam et elegi locum istum mihi in domum sacrificii.
2CHR|7|13|Si clausero caelum, et pluvia non fluxerit, et mandavero et praecepero locustae, ut devoret terram, et misero pestilentiam in populum meum,
2CHR|7|14|humiliatus autem populus meus, super quos invocatum est nomen meum, deprecatus me fuerit et exquisierit faciem meam et egerit paenitentiam a viis suis pessimis, ego exaudiam de caelo et propitius ero peccatis eorum et sanabo terram eorum.
2CHR|7|15|Nunc oculi mei erunt aperti, et aures meae attentae ad orationem eius, qui in loco isto oraverit;
2CHR|7|16|elegi enim et sanctificavi locum istum, ut sit nomen meum ibi in sempiternum, et permaneant oculi mei et cor meum ibi cunctis diebus.
2CHR|7|17|Tu quoque, si ambulaveris coram me, sicut ambulavit David pater tuus, et feceris iuxta omnia, quae praecepi tibi, et decreta et iudicia mea servaveris,
2CHR|7|18|stabiliam thronum regni tui, sicut pollicitus sum David patri tuo dicens: Non auferetur de stirpe tua vir, qui sit princeps in Israel.
2CHR|7|19|Si autem aversi fueritis et dereliqueritis decreta mea et praecepta mea, quae proposui vobis, et abeuntes servieritis diis alienis et adoraveritis eos,
2CHR|7|20|evellam vos de terra mea, quam dedi vobis, et domum hanc, quam sanctificavi nomini meo, proiciam a facie mea et tradam eam in parabolam et in fabulam cunctis populis.
2CHR|7|21|Et super domo ista, quae erat excelsa, universi transeuntes stupebunt et dicent: "Quare fecit Dominus sic terrae huic et domui huic?".
2CHR|7|22|Respondebuntque: "Quia dereliquerunt Dominum, Deum patrum suorum, qui eduxit eos de terra Aegypti, et apprehenderunt deos alienos et adoraverunt eos et coluerunt, idcirco venerunt super eos universa haec mala" ".
2CHR|8|1|Expletis autem viginti annis, postquam aedificavit Salomon domum Domini et domum suam,
2CHR|8|2|civitates, quas dederat Hiram Salomoni, aedificavit et habitare ibi fecit filios Israel.
2CHR|8|3|Abiit quoque in Emath Soba et obtinuit eam.
2CHR|8|4|Et aedificavit Palmyram in deserto et omnes civitates horreorum, quas aedificavit in Emath.
2CHR|8|5|Exstruxitque Bethoron superiorem et Bethoron inferiorem, civitates munitas habentes muros et portas et vectes,
2CHR|8|6|Baalath etiam et omnes urbes horreorum, quae fuerunt Salomonis, cunctasque urbes quadrigarum et urbes equorum. Omnia quaecumque voluit Salomon atque disposuit, aedificavit in Ierusalem et in Libano et in universa terra potestatis suae.
2CHR|8|7|Omnem populum, qui derelictus fuerat de Hetthaeis et Amorraeis et Pherezaeis et Hevaeis et Iebusaeis, qui non erant de stirpe Israel,
2CHR|8|8|de filiis eorum, qui remanserant post eos in terra, quos non interfecerant filii Israel, subiugavit Salomon in tributarios usque in diem hanc.
2CHR|8|9|Porro de filiis Israel non posuit, ut servirent operibus regis; ipsi enim erant viri bellatores et principes pugnatorum eius et principes quadrigarum et equitum eius.
2CHR|8|10|Omnes autem principes praefectorum regis Salomonis fuerunt ducenti quinquaginta, qui praefuerant populo.
2CHR|8|11|Filiam vero pharaonis transtulit de civitate David in domum, quam aedificaverat ei; dixit enim rex: " Non habitabit mulier mihi in domo David regis Israel, eo quod sanctificata sit, quia ingressa est in eam arca Domini ".
2CHR|8|12|Tunc obtulit Salomon holocausta Domino super altare Domini, quod exstruxerat ante porticum,
2CHR|8|13|ut per singulos dies offerretur in eo iuxta praeceptum Moysi in sabbatis et in calendis et in festis diebus ter per annum, id est in sollemnitate Azymorum et in sollemnitate Hebdomadarum et in sollemnitate Tabernaculorum.
2CHR|8|14|Et constituit iuxta dispositionem David patris sui officia sacerdotum in ministeriis suis et Levitas in ordine suo, ut laudarent et ministrarent coram sacerdotibus iuxta ritum uniuscuiusque diei, et ianitores in divisionibus suis per portam et portam; sic enim praeceperat David homo Dei.
2CHR|8|15|Nec praetergressi sunt mandata regis de sacerdotibus et Levitis in omnibus et in custodiis thesaurorum.
2CHR|8|16|Et firmatum est totum opus Salomonis ex eo die, quo fundavit domum Domini, usque in diem, quo perfecit eam.
2CHR|8|17|Tunc abiit Salomon in Asiongaber et in Ailath ad oram maris Rubri, quae est in terra Edom.
2CHR|8|18|Misit autem ei Hiram per manus servorum suorum naves et nautas gnaros maris; et abierunt cum servis Salomonis in Ophir tuleruntque inde quadringenta quinquaginta talenta auri et attulerunt ad regem Salomonem.
2CHR|9|1|Regina quoque Saba, cum audisset famam Salomonis, venit, ut tentaret eum in aenigmatibus in Ierusalem cum magno comitatu et camelis, qui portabant aromata et auri plurimum gemmasque pretiosas. Cumque venisset ad Salomonem, locuta est ei, quaecumque erant in corde suo.
2CHR|9|2|Et exposuit ei Salomon omnia, quae proposuerat, nec quidquam fuit quod ei non perspicuum fecerit.
2CHR|9|3|Quae postquam vidit, sapientiam scilicet Salomonis et domum, quam aedificaverat,
2CHR|9|4|necnon et cibaria mensae eius et sessionem servorum et officia ministrorum eius et vestimenta eorum, pincernas quoque et vestes eorum et victimas, quas immolabat in domo Domini, non erat prae stupore ultra in ea spiritus.
2CHR|9|5|Dixitque ad regem: " Verus est sermo, quem audieram in terra mea, de rebus tuis et sapientia tua;
2CHR|9|6|non credebam narrantibus, donec ipsa venissem, et vidissent oculi mei, et probassem vix medietatem sapientiae tuae mihi fuisse narratam; vicisti famam, quam audivi.
2CHR|9|7|Beati viri tui et beati servi tui, qui assistunt coram te omni tempore et audiunt sapientiam tuam!
2CHR|9|8|Sit Dominus Deus tuus benedictus, qui voluit te ordinare super thronum suum regem Domini Dei tui! Quia diligit Deus tuus Israel et vult servare eum in aeternum, idcirco posuit te super eum regem, ut facias iudicia atque iustitiam ".
2CHR|9|9|Dedit autem regi centum viginti talenta auri et aromata multa nimis et gemmas pretiosissimas; non fuerunt aromata talia ut haec, quae dedit regina Saba regi Salomoni.
2CHR|9|10|Sed et servi Hiram cum servis Salomonis attulerunt aurum de Ophir et ligna thyina et gemmas pretiosissimas;
2CHR|9|11|et fecit rex de lignis thyinis gradus in domo Domini et in domo regia, citharas quoque et psalteria cantoribus. Numquam visa sunt in terra Iudae ligna talia.
2CHR|9|12|Rex autem Salomon dedit reginae Saba cuncta, quae voluit et quae postulavit, et multo plura quam attulerat ad eum. Quae reversa abiit in terram suam cum servis suis.
2CHR|9|13|Erat autem pondus auri, quod afferebatur Salomoni per singulos annos, sescenta sexaginta sex talenta auri,
2CHR|9|14|excepta ea summa, quae proveniebat ex tributis mercatorum et negotiatorum afferentium et omnium regum Arabiae et ducum terrae, qui comportabant aurum et argentum Salomoni.
2CHR|9|15|Fecit igitur rex Salomon ducenta scuta aurea de summa sescentorum aureorum, qui in singulis scutis expendebantur,
2CHR|9|16|trecentas quoque peltas aureas trecentorum aureorum, quibus tegebantur singulae peltae, posuitque ea rex in domo Saltus Libani.
2CHR|9|17|Fecit quoque rex solium eburneum grande et vestivit illud auro mundissimo;
2CHR|9|18|sex quoque gradus, quibus ascendebatur ad solium, et scabellum aureum et brachiola duo altrinsecus et duos leones stantes iuxta brachiola,
2CHR|9|19|sed et alios duodecim leunculos stantes super sex gradus ex utraque parte; non fuit tale solium in universis regnis.
2CHR|9|20|Omnia quoque vasa convivii regis erant aurea, et vasa domus Saltus Libani ex auro purissimo; argentum enim in diebus Salomonis pro nihilo reputabatur.
2CHR|9|21|Siquidem naves regis ibant in Tharsis cum servis Hiram; semel in annis tribus veniebant naves Tharsis portantes aurum et argentum et ebur et simias et pavos.
2CHR|9|22|Magnificatus est igitur rex Salomon super omnes reges terrae divitiis et sapientia.
2CHR|9|23|Omnesque reges terrarum desiderabant faciem videre Salomonis, ut audirent sapientiam, quam dederat Deus in corde eius,
2CHR|9|24|et deferebant ei munera, vasa argentea et aurea et vestes et arma et aromata, equos et mulos per singulos annos.
2CHR|9|25|Habuit quoque Salomon quattuor milia stabula equorum et curruum equitumque duodecim milia; constituitque eos in urbibus quadrigarum et, ubi erat rex, in Ierusalem.
2CHR|9|26|Exercuit etiam potestatem super cunctos reges, a fluvio Euphrate usque ad terram Philisthinorum et usque ad terminos Aegypti;
2CHR|9|27|tantamque copiam praebuit argenti in Ierusalem quasi lapidum, et cedrorum tantam multitudinem velut sycomororum, quae gignuntur in Sephela.
2CHR|9|28|Adducebantur autem ei equi de Aegypto cunctisque regionibus.
2CHR|9|29|Reliqua vero operum Salomonis priorum et novissimorum scripta sunt in verbis Nathan prophetae et in prophetia Ahiae Silonitis, in visione quoque Addo videntis super Ieroboam filium Nabat.
2CHR|9|30|Regnavit autem Salomon in Ierusalem super omnem Israel quadraginta annis;
2CHR|9|31|dormivitque cum patribus suis, et sepelierunt eum in civitate David patris eius. Regnavitque Roboam filius eius pro eo.
2CHR|10|1|Profectus est autem Roboam in Sichem; illuc enim cunctus Israel convenerat, ut constituerent eum regem.
2CHR|10|2|Quod cum audisset Ieroboam filius Nabat, qui erat in Aegypto - fugerat quippe illuc ante Salomonem - statim reversus est;
2CHR|10|3|vocaveruntque eum, et venit cum universo Israel, et locuti sunt ad Roboam dicentes:
2CHR|10|4|" Pater tuus durissimo iugo nos pressit; tu leviora impera patre tuo, qui nobis gravem imposuit servitutem, et paululum de onere subleva, et serviemus tibi ".
2CHR|10|5|Qui ait: " Post tres dies revertimini ad me ".Cumque abisset populus,
2CHR|10|6|iniit rex Roboam consilium cum senibus, qui steterant coram patre eius Salomone, dum adhuc viveret, dicens: " Quid datis consilii, ut respondeam populo? ".
2CHR|10|7|Qui dixerunt ei: " Si placueris populo huic et lenieris eos verbis clementibus, servient tibi omni tempore ".
2CHR|10|8|At ille reliquit consilium senum et cum iuvenibus tractare coepit, qui cum eo nutriti fuerant et erant in comitatu illius.
2CHR|10|9|Dixitque ad eos: " Quid vobis videtur, vel respondere quid debemus populo huic, qui dixit mihi: "Subleva iugum, quod imposuit nobis pater tuus"? ".
2CHR|10|10|Et responderunt iuvenes, qui nutriti fuerant cum eo, atque dixerunt: " Sic loqueris populo, qui dixit tibi: "Pater tuus aggravavit iugum nostrum, tu subleva", et sic respondebis eis: Minimus digitus meus grossior est lumbis patris mei;
2CHR|10|11|pater meus imposuit vobis iugum grave, et ego maius pondus apponam; pater meus cecidit vos flagellis, ego vero caedam scorpionibus ".
2CHR|10|12|Venit ergo Ieroboam et universus populus ad Roboam die tertio, sicut praeceperat eis rex dicens: "Revertimini ad me die tertio ".
2CHR|10|13|Responditque rex dura, derelicto consilio seniorum;
2CHR|10|14|locutusque est iuxta iuvenum voluntatem: Pater meus grave vobis imposuit iugum,quod ego gravius faciam.Pater meus cecidit vos flagellis,ego vero caedam scorpionibus ".
2CHR|10|15|Et non acquievit populi precibus. Erat enim voluntatis Dei, ut compleretur sermo eius, quem locutus fuerat per manum Ahiae Silonitis ad Ieroboam filium Nabat.
2CHR|10|16|Israel autem universus videns quod noluisset eos audire rex, locutus est ad eum: Non est nobis pars in David,neque hereditas in filio Isai!Revertere in tabernacula tua, Israel!Tu autem vide domum tuam, David! ".Et abiit Israel in tabernacula sua.
2CHR|10|17|Super filios autem Israel, qui habitabant in civitatibus Iudae, regnavit Roboam.
2CHR|10|18|Misitque rex Roboam Adoram, qui praeerat servituti, et lapidaverunt eum filii Israel, et mortuus est. Porro rex Roboam currum festinavit ascendere et fugit in Ierusalem.
2CHR|10|19|Recessitque Israel a domo David usque ad diem hanc.
2CHR|11|1|Venit autem Roboam in Ie rusalem et convocavit univer sam domum Iudae et Beniamin, centum octoginta milia electorum bellantium, ut dimicaret contra Israel et converteret ad se regnum suum.
2CHR|11|2|Factusque est sermo Domini ad Semeiam hominem Dei dicens:
2CHR|11|3|" Loquere ad Roboam filium Salomonis regem Iudae et ad universum Israel, qui est in Iuda et Beniamin:
2CHR|11|4|Haec dicit Dominus: Non ascendetis neque pugnabitis contra fratres vestros. Revertatur unusquisque in domum suam, quia mea hoc gestum est voluntate ". Qui cum audissent sermonem Domini, reversi sunt nec perrexerunt contra Ieroboam.
2CHR|11|5|Habitavit autem Roboam in Ierusalem et aedificavit civitates muratas in Iuda.
2CHR|11|6|Exstruxitque Bethlehem et Etam et Thecue,
2CHR|11|7|Bethsur quoque et Socho et Odollam
2CHR|11|8|necnon Geth et Maresa et Ziph,
2CHR|11|9|sed et Aduram et Lachis et Azeca,
2CHR|11|10|Saraa quoque et Aialon et Hebron, quae erant in Iuda et Beniamin civitates munitissimas.
2CHR|11|11|Cumque clausisset eas muris, posuit in eis principes ciborumque horrea et olei et vini.
2CHR|11|12|Sed et in singulis urbibus fecit armamentarium scutorum et hastarum firmavitque eas summa diligentia et imperavit super Iudam et Beniamin.
2CHR|11|13|Sacerdotes autem et Levitae, qui erant in universo Israel, venerunt ad eum de cunctis sedibus suis.
2CHR|11|14|Levitae relinquentes suburbana et possessiones suas transierunt ad Iudam et Ierusalem, eo quod abiecisset eos Ieroboam et posteri eius, ne sacerdotio Domini fungerentur.
2CHR|11|15|Qui constituit sibi sacerdotes excelsorum et daemoniorum vitulorumque, quos fecerat.
2CHR|11|16|Sed sequentes eos et de cunctis tribubus Israel quicumque dederant cor suum, ut quaererent Dominum, Deum Israel, venerunt Ierusalem ad immolandum victimas Domino, Deo patrum suorum.
2CHR|11|17|Et roboraverunt regnum Iudae et confirmaverunt Roboam filium Salomonis per tres annos; ambulaverunt enim in viis David et Salomonis annis tantum tribus.
2CHR|11|18|Duxit autem Roboam uxorem Mahalath filiam Ierimoth filii David et Abihail filiae Eliab filii Isai,
2CHR|11|19|quae peperit ei filios Iehus et Samariam et Zoom.
2CHR|11|20|Post hanc quoque accepit Maacha filiam Absalom, quae peperit ei Abia et Ethai et Ziza et Salomith.
2CHR|11|21|Amavit autem Roboam Maacha filiam Absalom super omnes uxores suas et concubinas; nam uxores decem et octo duxerat, concubinas autem sexaginta. Et genuit viginti octo filios et sexaginta filias.
2CHR|11|22|Constituit vero in capite Abiam filium Maacha ducem super fratres suos; ipsum enim regem facere cogitabat.
2CHR|11|23|Et sapienter filios suos dispersit in cunctis finibus Iudae et Beniamin in universis civitatibus muratis. Praebuitque eis escas plurimas et multas petivit uxores.
2CHR|12|1|Cumque roboratum fuisset regnum Roboam et conforta tum, dereliquit legem Domini, et omnis Israel cum eo.
2CHR|12|2|Anno autem quinto regni Roboam ascendit Sesac rex Aegypti in Ierusalem - quia peccaverunt Domino -
2CHR|12|3|cum mille ducentis curribus et sexaginta milibus equitum, nec erat numerus vulgi, quod venerat cum eo ex Aegypto, Libyes scilicet et Socciitae et Aethiopes.
2CHR|12|4|Cepitque civitates munitissimas in Iuda et venit usque Ierusalem.
2CHR|12|5|Semeias autem propheta ingressus est ad Roboam et principes Iudae, qui congregati fuerant in Ierusalem fugientes Sesac, dixitque ad eos: " Haec dicit Dominus: Vos reliquistis me, et ego reliqui vos in manu Sesac ".
2CHR|12|6|Humiliatique principes Israel et rex dixerunt: " Iustus est Dominus! ".
2CHR|12|7|Cumque vidisset Dominus quod humiliati essent, factus est sermo Domini ad Semeiam dicens: " Quia humiliati sunt, non disperdam eos daboque eis mox effugium, et non effundetur furor meus super Ierusalem per manum Sesac.
2CHR|12|8|Verumtamen servient ei, ut sciant distantiam servitutis meae et servitutis regni terrarum ".
2CHR|12|9|Ascendit itaque Sesac rex Aegypti in Ierusalem, sublatis thesauris domus Domini et domus regis; omniaque secum tulit et clipeos aureos, quos fecerat Salomon.
2CHR|12|10|Pro quibus fecit rex Roboam aeneos et tradidit illos principibus cursorum, qui custodiebant vestibulum palatii.
2CHR|12|11|Cumque introiret rex domum Domini, veniebant cursores et tollebant eos; iterumque referebant eos ad armamentarium suum.
2CHR|12|12|Verumtamen, quia humiliatus est, aversa est ab eo ira Domini, nec deletus est penitus; siquidem et in Iuda inventa sunt opera bona.
2CHR|12|13|Confortatus est igitur rex Roboam in Ierusalem atque regnavit. Quadraginta autem et unius anni erat, cum regnare coepisset, et decem septemque annis regnavit in Ierusalem urbe, quam elegit Dominus, ut confirmaret nomen suum ibi de cunctis tribubus Israel. Nomenque matris eius Naama Ammanitis.
2CHR|12|14|Fecit autem malum et non praeparavit cor suum, ut quaereret Dominum.
2CHR|12|15|Opera vero Roboam prima et novissima scripta sunt in verbis Semeiae prophetae et Addo videntis, genealogia quoque et bella, quae erant inter Roboam et Ieroboam cunctis diebus.
2CHR|12|16|Et dormivit Roboam cum patribus suis sepultusque est in civitate David; et regnavit Abia filius eius pro eo.
2CHR|13|1|Anno octavo decimo regis Ieroboam regnavit Abia su per Iudam.
2CHR|13|2|Tribus annis regnavit in Ierusalem. Nomenque matris eius Michaia filia Uriel de Gabaa.Et erat bellum inter Abiam et Ieroboam.
2CHR|13|3|Cumque inisset Abia certamen et haberet bellicosissimos viros electorum quadringenta milia, Ieroboam instruxit e contra aciem octingenta milia virorum, qui et ipsi electi erant et ad bella fortissimi.
2CHR|13|4|Stetit igitur Abia super montem Semaraim, qui est in monte Ephraim, et ait: " Audi, Ieroboam et omnis Israel:
2CHR|13|5|Num ignoratis quod Dominus, Deus Israel, dederit regnum David super Israel in sempiternum, ipsi et filiis eius, pactum salis?
2CHR|13|6|Et surrexit Ieroboam filius Nabat servus Salomonis filii David et rebellavit contra dominum suum;
2CHR|13|7|congregatique sunt ad eum viri vanissimi, filii Belial, et praevaluerunt contra Roboam filium Salomonis. Porro Roboam erat iuvenis et corde pavido nec potuit resistere eis.
2CHR|13|8|Nunc ergo vos dicitis quod resistere possitis regno Domini, quod possidet per filios David, habetisque grandem populi multitudinem atque vitulos aureos, quos fecit vobis Ieroboam in deos.
2CHR|13|9|Et eiecistis sacerdotes Domini filios Aaron atque Levitas et fecistis vobis sacerdotes sicut populi terrarum. Quicumque venerit et initiaverit manum suam in tauro de bobus et in arietibus septem, fit sacerdos eorum, qui non sunt dii.
2CHR|13|10|Noster autem Deus Dominus est, quem non reliquimus; sacerdotesque ministrant Domino de filiis Aaron, et Levitae sunt in ordine suo.
2CHR|13|11|Holocausta quoque offerunt Domino per singulos dies, mane et vespere, et thymiama aromatum, et proponuntur panes in mensa mundissima. Estque apud nos candelabrum aureum et lucernae eius, ut accendantur semper ad vesperam; nos quippe custodimus praecepta Domini Dei nostri, quem vos reliquistis.
2CHR|13|12|Ergo in exercitu nostro dux Deus est et sacerdotes eius, qui clangunt tubis et resonant contra vos, filii Israel; nolite pugnare contra Dominum, Deum patrum vestrorum, quia non vobis expedit ".
2CHR|13|13|Ieroboam autem retro moliebatur insidias, ut venirent post eos, et erant ante Iudam, et insidiae post eos.
2CHR|13|14|Respiciensque Iuda vidit instare bellum ex adverso et post tergum et clamavit ad Dominum, ac sacerdotes tubis canere coeperunt,
2CHR|13|15|omnesque viri Iudae vociferati sunt; et ecce, illis clamantibus, perterruit Deus Ieroboam et omnem Israel coram Abia et Iuda.
2CHR|13|16|Fugeruntque filii Israel Iudam, et tradidit eos Deus in manu eorum.
2CHR|13|17|Percussit ergo eos Abia et populus eius plaga magna; et corruerunt vulnerati ex Israel quingenta milia virorum fortium.
2CHR|13|18|Humiliatique sunt filii Israel in tempore illo, et confortati filii Iudae, eo quod sperassent in Domino, Deo patrum suorum.
2CHR|13|19|Persecutus est autem Abia fugientem Ieroboam et cepit civitates eius Bethel et filias eius et Iesana cum filiabus suis, Ephron quoque et filias eius.
2CHR|13|20|Nec invaluit ultra Ieroboam in diebus Abiae. Quem percussit Dominus, et mortuus est.
2CHR|13|21|Abia autem confortatus est et accepit sibi uxores quattuordecim procreavitque viginti duos filios et sedecim filias.
2CHR|13|22|Reliqua autem gestorum Abiae viarumque et sermonum eius scripta sunt in enarratione prophetae Addo.
2CHR|13|23|Dormivit autem Abia cum patribus suis, et sepelierunt eum in civitate David; regnavitque Asa filius eius pro eo. In cuius diebus quievit terra annis decem.
2CHR|14|1|Fecit autem Asa, quod bo num et placitum erat in con spectu Domini Dei sui, et subvertit altaria peregrini cultus et excelsa
2CHR|14|2|et confregit lapides palosque succidit
2CHR|14|3|ac praecepit Iudae, ut quaereret Dominum, Deum patrum suorum, et faceret legem et universa mandata,
2CHR|14|4|et abstulit e cunctis urbibus Iudae excelsa et thymiateria et regnavit in pace.
2CHR|14|5|Aedificavit quoque urbes munitas in Iuda, quia quievit terra, et nulla temporibus eius bella surrexerant, pacem Domino ei largiente.
2CHR|14|6|Dixit autem Iudae: " Aedificemus civitates istas et vallemus muris et roboremus turribus et portis et seris, donec a bellis quieta sunt omnia; quia quaesivimus Dominum Deum nostrum, quaesivit nos et dedit nobis pacem per gyrum ". Aedificaverunt igitur et prosperati sunt.
2CHR|14|7|Habuit autem Asa exercitum portantium scuta et hastas de Iuda trecenta milia, de Beniamin vero scutariorum et sagittariorum ducenta octoginta milia; omnes isti viri fortissimi.
2CHR|14|8|Egressus est autem contra eos Zara Aethiops cum exercitu, decies centena milia et curribus trecentis, et venit usque Maresa.
2CHR|14|9|Porro Asa perrexit obviam ei, et instruxerunt aciem ad bellum in valle, quae est ad septentrionem Maresa,
2CHR|14|10|et invocavit Asa Dominum Deum suum et ait: " Domine, non est apud te ulla distantia, utrum paucis auxilieris an pluribus; adiuva nos, Domine Deus noster. In te enim et in tuo nomine habentes fiduciam venimus contra hanc multitudinem. Domine, Deus noster tu es, non praevaleat contra te homo ".
2CHR|14|11|Exterruit itaque Dominus Aethiopes coram Asa et Iuda; fugeruntque Aethiopes.
2CHR|14|12|Et persecutus est eos Asa et populus, qui cum eo erat, usque Gerar; et ruerunt Aethiopes usque ad internecionem, quia Domino caedente contriti sunt et exercitu illius proeliante. Tulerunt ergo spolia multa
2CHR|14|13|et percusserunt omnes civitates per circuitum Gerarae; terror quippe Domini eos invaserat. Et diripuerunt omnes urbes et multam praedam asportaverunt.
2CHR|14|14|Sed et caulas ovium destruentes tulerunt pecorum infinitam multitudinem et camelorum reversique sunt Ierusalem.
2CHR|15|1|Azarias autem filius Oded, facto in se spiritu Dei,
2CHR|15|2|egressus est in occursum Asa et dixit ei: " Audite me, Asa et omnis Iuda et Beniamin! Dominus vobiscum, quia fuistis cum eo. Si quaesieritis eum, invenietur a vobis; si autem dereliqueritis eum, derelinquet vos.
2CHR|15|3|Transierunt autem multi dies in Israel absque Deo veritatis et absque sacerdote doctore et absque lege.
2CHR|15|4|Cumque reversi essent in angustia sua ad Dominum, Deum Israel, et quaesivissent eum, inventus est ab eis.
2CHR|15|5|In temporibus illis non erat pax egredienti et ingredienti sed perturbatio magna multa in cunctis habitatoribus terrarum;
2CHR|15|6|contundebatur enim gens contra gentem, et civitas contra civitatem, quia Dominus conturbabat eos in omni angustia.
2CHR|15|7|Vos autem confortamini, et non dissolvantur manus vestrae; erit enim merces operi vestro ".
2CHR|15|8|Cum audisset Asa verba haec et prophetiam, confortatus est et abstulit idola de omni terra Iudae et Beniamin et ex urbibus, quas ceperat montis Ephraim, et dedicavit altare Domini, quod erat ante porticum Domini.
2CHR|15|9|Congregavitque universum Iudam et Beniamin et advenas cum eis de Ephraim et de Manasse et de Simeon; plures enim ad eum confugerant ex Israel videntes quod Dominus Deus illius esset cum eo.
2CHR|15|10|Cumque convenissent in Ierusalem mense tertio anno quinto decimo regni Asa,
2CHR|15|11|immolaverunt Domino in die illa de manubiis, quas adduxerant: boves septingentos et oves septem milia.
2CHR|15|12|Et inierunt foedus, ut quaererent Dominum, Deum patrum suorum, in toto corde et in tota anima sua:
2CHR|15|13|si quis autem non quaesierit Dominum, Deum Israel, moriatur a minimo usque ad maximum, a viro usque ad mulierem.
2CHR|15|14|Iuraveruntque Domino voce magna in iubilo et in clangore tubarum et in sonitu bucinarum.
2CHR|15|15|Omnes, qui erant in Iuda, gavisi sunt de iuramento; in omni enim corde suo iuraverant et in tota voluntate quaesierant eum, et inventus fuerat ab eis. Praestititque eis Dominus requiem per circuitum.
2CHR|15|16|Sed et Maacham matrem Asa rex amovit, ne esset domina, eo quod fecisset simulacrum Aserae; quod contrivit Asa et in frusta comminuens combussit in torrente Cedron.
2CHR|15|17|Excelsa autem derelicta sunt in Israel; attamen cor Asa erat perfectum cunctis diebus eius.
2CHR|15|18|Ea quae voverat pater suus et ipse, intulit in domum Dei, argentum et aurum vasorumque diversam supellectilem.
2CHR|15|19|Bellum vero non fuit usque ad tricesimum quintum annum regni Asa.
2CHR|16|1|Anno autem tricesimo sexto regni eius ascendit Baasa rex Israel in Iudam; et muro circumdabat Rama, ut nullus tute posset egredi et ingredi de regno Asa.
2CHR|16|2|Protulit ergo Asa argentum et aurum de thesauris domus Domini et domus regis misitque ad Benadad regem Syriae, qui habitabat in Damasco, dicens:
2CHR|16|3|" Foedus inter me et te est et inter patrem meum et patrem tuum; quam ob rem misi tibi argentum et aurum, ut, rupto foedere, quod habes cum Baasa rege Israel, facias eum a me recedere ".
2CHR|16|4|Acquiescens Benadad regi Asa misit principes exercituum suorum ad urbes Israel, qui percusserunt Ahion et Dan et Abelmaim et universa horrea urbium Nephthali.
2CHR|16|5|Quod cum audisset Baasa, desivit aedificare Rama et intermisit opus suum.
2CHR|16|6|Porro Asa rex assumpsit universum Iudam, et tulerunt lapides Rama et ligna, quibus aedificaverat Baasa, aedificavitque ex eis Gabaa et Maspha.
2CHR|16|7|In tempore illo venit Hanani videns ad Asa regem Iudae et dixit ei: " Quia habuisti fiduciam in rege Syriae et non in Domino Deo tuo, idcirco evasit Syriae regis exercitus de manu tua.
2CHR|16|8|Nonne Aethiopes et Libyes magnus exercitus erant quadrigis et equitibus et multitudine nimia, quos, cum Domino credidisses, tradidit in manu tua?
2CHR|16|9|Oculi enim Domini contemplantur universam terram et praebent fortitudinem his, qui corde perfecto credunt in eum. Stulte igitur egisti in hoc, quia ex praesenti tempore contra te bella consurgent ".
2CHR|16|10|Iratusque Asa adversus videntem iussit eum mitti in nervum, valde quippe super hoc fuerat indignatus; et vexavit Asa quosdam de populo in tempore illo.
2CHR|16|11|Opera autem Asa prima et novissima scripta sunt in libro regum Iudae et Israel.
2CHR|16|12|Aegrotavit etiam Asa anno tricesimo nono regni sui dolore pedum vehementissimo et nec in infirmitate sua quaesivit Dominum, sed magis in medicorum arte confisus est.
2CHR|16|13|Dormivitque Asa cum patribus suis et mortuus est anno quadragesimo primo regni sui.
2CHR|16|14|Et sepelierunt eum in sepulcro suo, quod foderat sibi in civitate David; posueruntque eum super lectum plenum aromatibus et variis unguentis, quae erant pigmentariorum arte confecta, et fecerunt in exsequiis eius combustionem splendidam valde.
2CHR|17|1|Regnavit autem Iosaphat filius eius pro eo et invaluit contra Israel.
2CHR|17|2|Constituitque militum numeros in cunctis urbibus Iudae, quae erant vallatae muris; praesidiaque disposuit in terra Iudae et in civitatibus Ephraim, quas ceperat Asa pater eius.
2CHR|17|3|Et fuit Dominus cum Iosaphat, quia ambulavit in viis patris sui primis et non speravit in Baalim
2CHR|17|4|sed in Deo patris sui et perrexit in praeceptis illius et non iuxta peccata Israel.
2CHR|17|5|Confirmavitque Dominus regnum in manu eius, et dedit omnis Iuda munera Iosaphat; factaeque sunt ei infinitae divitiae et multa gloria.
2CHR|17|6|Cumque sumpsisset cor eius audaciam propter vias Domini, etiam excelsa et palos de Iuda abstulit.
2CHR|17|7|Tertio autem anno regni sui misit principes suos Benhail et Abdiam et Zachariam et Nathanael et Michaiam, ut docerent in civitatibus Iudae,
2CHR|17|8|et cum eis Levitas Semeiam et Nathaniam et Zabadiam, Asael quoque et Semiramoth et Ionathan Adoniamque et Thobiam Levitas et cum eis Elisama et Ioram sacerdotes.
2CHR|17|9|Docebantque in Iuda habentes librum legis Domini et circuibant cunctas urbes Iudae atque erudiebant populum.
2CHR|17|10|Itaque factus est pavor Domini super omnia regna terrarum, quae erant per gyrum Iudae, nec audebant bellare contra Iosaphat.
2CHR|17|11|Sed et de Philisthim Iosaphat munera deferebant et vectigal argenti; Arabes quoque adducebant pecora arietum septem milia septingenta et hircos totidem.
2CHR|17|12|Crevit ergo Iosaphat et magnificatus est usque in sublime atque aedificavit in Iuda castella urbesque horreorum.
2CHR|17|13|Et multae copiae praesto erant ei in urbibus Iudae; viri quoque bellatores et robusti erant in Ierusalem,
2CHR|17|14|quorum iste numerus per familias singulorum: in Iuda principes exercitus, Ednas dux, et cum eo robustissimorum trecenta milia;
2CHR|17|15|et ad latus eius Iohanan princeps et cum eo ducenta octoginta milia;
2CHR|17|16|ad latus quoque istius Amasias filius Zechri consecratus Domino et cum eo ducenta milia virorum fortium;
2CHR|17|17|de Beniamin autem robustus ad proelia Eliada et cum eo tenentium arcum et clipeum ducenta milia;
2CHR|17|18|et ad latus eius Iozabad et cum eo centum octoginta milia expeditorum militum.
2CHR|17|19|Hi omnes erant ad manum regis, exceptis aliis, quos posuerat in urbibus muratis in universo Iuda.
2CHR|18|1|Fuit ergo Iosaphat dives et inclitus multum et affinitate coniunctus est Achab.
2CHR|18|2|Descenditque post annos ad eum in Samariam, ad cuius adventum mactavit Achab oves et boves plurimos ipsi et populo, qui venerat cum eo; persuasitque illi, ut ascenderet in Ramoth Galaad.
2CHR|18|3|Dixitque Achab rex Israel ad Iosaphat regem Iudae: " Veni mecum in Ramoth Galaad ". Cui ille respondit: " Ut ego, et tu; sicut populus tuus, sic et populus meus, tecumque erimus in bello ".
2CHR|18|4|Dixitque Iosaphat ad regem Israel: " Consule, obsecro, impraesentiarum sermonem Domini ".
2CHR|18|5|Congregavitque rex Israel prophetarum quadringentos viros et dixit ad eos: " In Ramoth Galaad ad bellandum ire debemus an quiescere? ". At illi: Ascende, inquiunt, et tradet Deus in manu regis ".
2CHR|18|6|Dixitque Iosaphat: " Numquid non est hic et alius propheta Domini, ut ab illo etiam requiramus? ".
2CHR|18|7|Et ait rex Israel ad Iosaphat: " Adhuc est vir unus, a quo possumus quaerere Domini voluntatem; sed ego odi eum, quia non prophetat mihi bonum sed malum omni tempore: est autem Michaeas filius Iemla ". Dixitque Iosaphat: " Ne loquaris, rex, hoc modo ".
2CHR|18|8|Vocavit ergo rex Israel unum de eunuchis et dixit ei: " Voca cito Michaeam filium Iemla ".
2CHR|18|9|Porro rex Israel et Iosaphat rex Iudae uterque sedebant in solio suo vestiti cultu regio; sedebant autem in area iuxta portam Samariae, omnesque prophetae vaticinabantur coram eis.
2CHR|18|10|Sedecias vero filius Chanaana fecit sibi cornua ferrea et ait: " Haec dicit Dominus: His ventilabis Syriam, donec conteras eam ".
2CHR|18|11|Omnesque prophetae similiter prophetabant atque dicebant: " Ascende in Ramoth Galaad et prosperaberis; et tradet Dominus in manu regis ".
2CHR|18|12|Nuntius autem, qui ierat ad vocandum Michaeam, ait illi: " En verba omnium prophetarum uno ore bona regi annuntiant; quaeso ergo te, ut et sermo tuus ab eis non dissentiat, loquarisque prospera ".
2CHR|18|13|Cui respondit Michaeas: " Vivit Dominus, quia, quodcumque dixerit Deus meus, hoc loquar! ".
2CHR|18|14|Venit ergo ad regem. Cui rex ait: " Michaea, ire debemus in Ramoth Galaad ad bellandum an quiescere? ". Cui ille respondit: " Ascendite et prosperamini, ut tradantur hostes in manus vestras ".
2CHR|18|15|Dixitque rex: " Iterum atque iterum te adiuro, ut non mihi loquaris nisi, quod verum est, in nomine Domini ".
2CHR|18|16|At ille ait: Vidi universum Israeldispersum in montibussicut oves absque pastore.Et dixit Dominus:Non habent isti dominum; revertatur unusquisque in domum suam in pace" ".
2CHR|18|17|Et ait rex Israel ad Iosaphat: " Nonne dixi tibi quod non prophetaret iste mihi quidquam boni sed ea, quae mala sunt? ".
2CHR|18|18|At ille idcirco ait: " Audite verbum Domini: Vidi Dominum sedentem in solio suo et omnem exercitum caeli assistentem ei a dextris et sinistris.
2CHR|18|19|Et dixit Dominus: "Quis decipiet Achab regem Israel, ut ascendat et corruat in Ramoth Galaad?". Cumque diceret unus hoc modo et alter alio,
2CHR|18|20|processit spiritus et stetit coram Domino et ait: "Ego decipiam eum". Cui Dominus: "In quo, inquit, decipies?".
2CHR|18|21|At ille respondit: "Egrediar et ero spiritus mendax in ore omnium prophetarum eius". Dixitque Dominus: "Decipies et praevalebis; egredere et fac ita".
2CHR|18|22|Nunc igitur, ecce dedit Dominus spiritum mendacii in ore omnium prophetarum tuorum et Dominus locutus est de te mala ".
2CHR|18|23|Accessit autem Sedecias filius Chanaana et percussit Michaeae maxillam et ait: " Per quam viam transivit spiritus Domini a me, ut loqueretur tibi? ".
2CHR|18|24|Dixitque Michaeas: " Tu ipse videbis in die illo, quando ingressus fueris cubiculum intra cubiculum, ut abscondaris ".
2CHR|18|25|Praecepit autem rex Israel dicens: " Tollite Michaeam et ducite eum ad Amon principem civitatis et ad Ioas filium regis
2CHR|18|26|et dicetis: "Haec dicit rex: Mittite hunc in carcerem et date ei panis modicum et aquae pauxillum, donec revertar in pace" ".
2CHR|18|27|Dixitque Michaeas: " Si reversus fueris in pace, non est locutus Dominus in me ". Et ait: " Audite, populi omnes! ".
2CHR|18|28|Igitur ascenderunt rex Israel et Iosaphat rex Iudae in Ramoth Galaad.
2CHR|18|29|Dixitque rex Israel ad Iosaphat: " Mutabo habitum et sic ad pugnam vadam; tu autem induere vestibus tuis ". Mutatoque rex Israel habitu venit ad bellum.
2CHR|18|30|Rex autem Syriae praeceperat ducibus curruum suorum dicens: " Ne pugnetis contra minimum aut contra maximum, nisi contra solum regem Israel.
2CHR|18|31|Itaque, cum vidissent principes curruum Iosaphat, dixerunt: " Rex Israel est iste! ". Et circumdederunt eum dimicantes. At ille clamavit ad Dominum, et auxiliatus est ei atque avertit eos Deus ab illo.
2CHR|18|32|Cum enim vidissent duces curruum quod non esset rex Israel, reliquerunt eum.
2CHR|18|33|Accidit autem, ut unus e populo sagittam in incertum iaceret et percuteret regem Israel inter iuncturas et loricam. At ille aurigae suo ait: " Converte manum tuam et educ me de acie, quia vulneratus sum ".
2CHR|18|34|Et aggravata est pugna in die illo; porro rex Israel stabat in curru suo contra Syros usque ad vesperam et mortuus est occidente sole.
2CHR|19|1|Reversus est autem Iosaphat rex Iudae in domum suam pacifice in Ierusalem.
2CHR|19|2|Cui occurrit Iehu filius Hanani videns et ait ad eum: " Impio praebes auxilium et his, qui oderunt Dominum, amicitia iungeris, et idcirco iram quidem Domini merebaris;
2CHR|19|3|sed bona opera inventa sunt in te, eo quod abstuleris palos de terra et praeparaveris cor tuum, ut requireres Deum ".
2CHR|19|4|Habitavit ergo Iosaphat in Ierusalem. Rursumque egressus est ad populum de Bersabee usque ad montem Ephraim et revocavit eos ad Dominum, Deum patrum suorum.
2CHR|19|5|Constituitque iudices terrae in cunctis civitatibus Iudae munitis per singula loca.
2CHR|19|6|Et praecipiens iudicibus: " Videte, ait, quid faciatis. Non enim homini exercetis iudicium sed Domino, qui vobiscum est, quando iudicaveritis.
2CHR|19|7|Sit timor Domini, vobiscum et caute cuncta facite; non est enim apud Dominum Deum nostrum iniquitas nec personarum acceptio nec cupido munerum.
2CHR|19|8|In Ierusalem quoque constituit Iosaphat ex Levitis et sacerdotibus et principibus familiarum Israel pro iudicio Domini et pro causis habitatorum Ierusalem.
2CHR|19|9|Praecepitque eis dicens: " Sic agetis in timore Domini fideliter et corde perfecto.
2CHR|19|10|Omnem causam, quae venerit ad vos fratrum vestrorum, qui habitant in urbibus suis, ubicumque quaestio est de homicidio, de lege, de mandato, de praeceptis et de iustificationibus, commonete eos, ut non peccent in Dominum, et ne veniat ira super vos et super fratres vestros; sic ergo agetis et non peccabitis.
2CHR|19|11|Amarias autem sacerdos princeps super vos in omnibus, quae ad Deum pertinent, praesidebit; porro Zabadias filius Ismael, qui est dux in domo Iudae, super ea opera erit, quae ad regis officium pertinent; habetisque Levitas coram vobis ut scribas. Confortamini et agite diligenter, et sit Dominus cum bonis ".
2CHR|20|1|Post haec congregati sunt filii Moab et filii Ammon et cum eis de Meunitis ad Iosaphat, ut pugnarent contra eum.
2CHR|20|2|Veneruntque nuntii et indicaverunt Iosaphat dicentes: " Venit contra te multitudo magna de his locis, quae trans mare sunt, de Edom, et ecce consistunt in Asasonthamar, quae est Engaddi ".
2CHR|20|3|Iosaphat autem timore perterritus totum se contulit ad rogandum Dominum et praedicavit ieiunium universo Iudae.
2CHR|20|4|Congregatusque est Iuda ad precandum Dominum; sed et de omnibus urbibus suis venerunt ad obsecrandum eum.
2CHR|20|5|Cumque stetisset Iosaphat in medio coetu Iudae et Ierusalem in domo Domini ante atrium novum,
2CHR|20|6|ait: " Domine, Deus patrum nostrorum, tu es Deus in caelo et dominaris cunctis regnis gentium; in manu tua est fortitudo et potentia, nec quisquam tibi potest resistere.
2CHR|20|7|Nonne tu, Deus noster, expulisti habitatores terrae huius coram populo tuo Israel et dedisti eam semini Abraham amici tui in sempiternum?
2CHR|20|8|Habitaveruntque in ea et exstruxerunt in illa sanctuarium nomini tuo dicentes:
2CHR|20|9|"Si irruerint super nos mala, gladius iudicii, pestilentia et fames, stabimus coram domo hac in conspectu tuo, quia nomen tuum est in domo hac, et clamabimus ad te in tribulationibus nostris, et exaudies salvosque facies".
2CHR|20|10|Nunc igitur ecce filii Ammon et Moab et mons Seir, per quos non concessisti Israeli ut transirent, quando egrediebantur de Aegypto, sed declinaverunt ab eis et non interfecerunt illos,
2CHR|20|11|e contrario agunt et nituntur eicere nos de possessione tua, quam tradidisti nobis.
2CHR|20|12|Deus noster, ergo non iudicabis eos? In nobis quidem non tanta est fortitudo, ut possimus huic multitudini resistere, quae irruit super nos; sed, cum ignoremus quid agere debeamus, hoc solum habemus residui, ut oculos nostros dirigamus ad te ".
2CHR|20|13|Omnis vero Iuda stabat coram Domino cum parvulis et uxoribus et liberis suis.
2CHR|20|14|Erat autem Iahaziel filius Zachariae filii Banaiae filii Iehiel filii Matthaniae Levites de filiis Asaph, super quem factus est spiritus Domini in medio congregationis,
2CHR|20|15|et ait: " Attendite, omnis Iuda et qui habitatis Ierusalem et tu rex Iosaphat: Haec dicit Dominus vobis: Nolite timere nec paveatis hanc multitudinem magnam; non est enim vestra pugna sed Dei.
2CHR|20|16|Cras descendetis contra eos; ascensuri enim sunt per clivum nomine Sis, et invenietis illos in summitate torrentis, qui est contra solitudinem Ieruel.
2CHR|20|17|Non eritis vos, qui dimicabitis; sed tantummodo confidenter state et videbitis auxilium Domini super vos, o Iuda et Ierusalem. Nolite timere nec paveatis; cras egredimini contra eos, et Dominus erit vobiscum ".
2CHR|20|18|Iosaphat ergo inclinavit se super faciem suam in terra, et omnis Iuda et habitatores Ierusalem ceciderunt coram Domino et adoraverunt eum.
2CHR|20|19|Porro Levitae de filiis Caath, de filiis Core scilicet, surrexerunt et laudabant Dominum, Deum Israel, voce magna in excelsum.
2CHR|20|20|Cumque mane surrexissent, egressi sunt ad desertum Thecue; profectisque eis, stans Iosaphat in medio eorum dixit: " Audite me, Iuda et habitatores Ierusalem! Credite in Domino Deo vestro et permanebitis; credite prophetis eius, et cuncta evenient vobis prospera ".
2CHR|20|21|Habuitque consilium cum populo et statuit cantores Domini, ut laudarent eum in ornatu sancto et antecederent exercitum ac voce consona dicerent: " Confitemini Domino, quoniam in aeternum misericordia eius ".
2CHR|20|22|Cumque coepissent laudes canere, vertit Dominus insidias eorum contra filios Ammon et Moab et montem Seir, qui egressi fuerant, ut pugnarent contra Iudam, et percussi sunt.
2CHR|20|23|Et filii Ammon et Moab consurrexerunt adversum habitatores montis Seir, ut interficerent et delerent eos; cumque hoc opere perpetrassent, etiam in semetipsos versi mutuis concidere vulneribus.
2CHR|20|24|Porro Iuda, cum venisset ad speculam, quae respicit solitudinem, vidit procul omnem late regionem plenam cadaveribus, nec superesse quemquam, qui necem potuisset evadere.
2CHR|20|25|Venit ergo Iosaphat et omnis populus cum eo ad detrahenda spolia mortuorum inveneruntque iumenta multa et supellectilem, vestes quoque et vasa pretiosissima et diripuerunt, ita ut omnia portare non possent, et per tres dies spolia auferebant pro praedae magnitudine.
2CHR|20|26|Die autem quarto congregati sunt in valle Baracha; etenim, quoniam ibi benedixerant Domino, vocaverunt locum illum vallis Benedictionis usque in praesentem diem.
2CHR|20|27|Reversusque est omnis vir Iudae et Ierusalem et Iosaphat ante eos in Ierusalem cum laetitia magna, eo quod dedisset eis Dominus gaudium de inimicis suis;
2CHR|20|28|ingressique sunt Ierusalem cum psalteriis et citharis et tubis in domum Domini.
2CHR|20|29|Irruit autem pavor Dei super universa regna terrarum, cum audissent quod pugnasset Dominus contra inimicos Israel.
2CHR|20|30|Quievitque regnum Iosaphat, et praebuit ei Deus eius pacem per circuitum.
2CHR|20|31|Regnavit igitur Iosaphat super Iudam. Et erat triginta quinque annorum, cum regnare coepisset; viginti autem et quinque annis regnavit in Ierusalem. Nomen matris eius Azuba filia Selachi.
2CHR|20|32|Et ambulavit in via patris sui Asa nec declinavit ab ea, faciens quod rectum erat coram Domino.
2CHR|20|33|Verumtamen excelsa non ablata sunt; et adhuc populus non direxerat cor suum ad Deum patrum suorum.
2CHR|20|34|Reliqua autem gestorum Iosaphat, priorum et novissimorum, scripta sunt in verbis Iehu filii Hanani, quae digesta sunt in libros regum Israel.
2CHR|20|35|Post haec iniit amicitias Iosaphat rex Iudae cum Ochozia rege Israel, cuius opera fuerunt impiissima,
2CHR|20|36|et particeps fuit, ut facerent naves, quae irent in Tharsis, feceruntque classem in Asiongaber.
2CHR|20|37|Prophetavit autem Eliezer filius Dodiae de Maresa contra Iosaphat dicens: " Quia habuisti foedus cum Ochozia, percussit Dominus opera tua ". Contritaeque sunt naves nec potuerunt ire in Tharsis.
2CHR|21|1|Dormivit autem Iosaphat cum patribus suis et sepultus est cum eis in civitate David; regnavitque Ioram filius eius pro eo.
2CHR|21|2|Qui habuit fratres filios Iosaphat Azariam et Iahiel et Zachariam et Azariam et Michael et Saphatiam: omnes hi filii Iosaphat regis Israel.
2CHR|21|3|Deditque eis pater suus multa munera argenti et auri et res pretiosas cum civitatibus munitissimis in Iuda; regnum autem tradidit Ioram, eo quod esset primogenitus.
2CHR|21|4|Surrexit ergo Ioram super regnum patris sui; cumque se confirmasset, occidit omnes fratres suos gladio et quosdam de principibus Israel.
2CHR|21|5|Triginta duorum annorum erat Ioram, cum regnare coepisset, et octo annis regnavit in Ierusalem.
2CHR|21|6|Ambulavitque in viis regum Israel, sicut egerat domus Achab; filia quippe Achab erat uxor eius. Et fecit malum in conspectu Domini.
2CHR|21|7|Noluit autem Dominus disperdere domum David propter pactum, quod inierat cum eo, et quia promiserat, ut daret ei lucernam et filiis eius omni tempore.
2CHR|21|8|In diebus illis rebellavit Edom, ne esset subditus Iudae, et constituit sibi regem.
2CHR|21|9|Cumque transisset Ioram cum principibus suis et cunctis curribus, qui erant secum, surrexit nocte et percussit Edom, qui eum circumdederat, et omnes duces curruum eius.
2CHR|21|10|Attamen rebellavit Edom, ne esset sub dicione Iudae, usque ad hanc diem. Eo tempore et Lobna recessit, ne esset sub manu illius; dereliquerat enim Dominum, Deum patrum suorum.
2CHR|21|11|Insuper et excelsa fabricatus est in montibus Iudae et fornicari fecit habitatores Ierusalem et praevaricari Iudam.
2CHR|21|12|Allatae sunt autem ei litterae ab Elia propheta, in quibus scriptum erat: "Haec dicit Dominus, Deus David patris tui: Quoniam non ambulasti in viis Iosaphat patris tui et in viis Asa regis Iudae,
2CHR|21|13|sed incessisti per iter regum Israel et fornicari fecisti Iudam et habitatores Ierusalem imitatus fornicationem domus Achab, insuper et fratres tuos domum patris tui meliores te occidisti:
2CHR|21|14|ecce Dominus percutiet plaga magna populum tuum, filios et uxores tuas universamque substantiam tuam;
2CHR|21|15|tu autem aegrotabis pessimo languore uteri tui, donec egrediantur vitalia tua paulatim per singulos dies ".
2CHR|21|16|Suscitavit ergo Dominus contra Ioram spiritum Philisthinorum et Arabum, qui confines sunt Aethiopibus,
2CHR|21|17|et ascenderunt in terram Iudae et irruperunt in eam diripueruntque cunctam substantiam, quae inventa est in domo regis, insuper et filios eius et uxores, nec remansit ei filius nisi Ioachaz, qui minimus natu erat.
2CHR|21|18|Et post haec omnia percussit eum Dominus alvi languore insanabili.
2CHR|21|19|Cumque diei succederet dies, et temporum spatia volverentur, duorum annorum expletus est circulus; et sic longa consumptus tabe, ita ut egereret etiam viscera sua, languore pariter et vita caruit. Mortuusque est in infirmitate pessima, et non fecit ei populus eius secundum morem combustionis exsequias, sicut fecerat maioribus eius.
2CHR|21|20|Triginta duorum annorum fuit, cum regnare coepisset, et octo annis regnavit in Ierusalem. Obiitque nullo relicto desiderio sui; et sepelierunt eum in civitate David, verumtamen non in sepulcro regum.
2CHR|22|1|Constituerunt autem habita tores Ierusalem Ochoziam fi lium eius minimum regem pro eo; omnes enim maiores natu interfecerat turba, quae irruerat cum Arabibus in castra. Regnavitque Ochozias filius Ioram regis Iudae.
2CHR|22|2|Filius viginti duo annorum erat Ochozias, cum regnare coepisset, et uno anno regnavit in Ierusalem. Nomen matris eius Athalia filia Amri.
2CHR|22|3|Sed et ipse ingressus est per vias domus Achab; mater enim eius impulit eum, ut impie ageret.
2CHR|22|4|Fecit igitur malum in conspectu Domini sicut domus Achab; ipsi enim fuerunt ei consiliarii post mortem patris sui in interitum eius.
2CHR|22|5|Ambulavitque in consiliis eorum et perrexit cum Ioram filio Achab rege Israel in bellum contra Hazael regem Syriae in Ramoth Galaad; vulneraveruntque Syri Ioram.
2CHR|22|6|Qui reversus est, ut curaretur in Iezrahel a plagis, quas acceperat in supradicto certamine.Igitur Ochozias filius Ioram rex Iudae descendit, ut inviseret Ioram filium Achab in Iezrahel aegrotantem.
2CHR|22|7|Voluntatis quippe fuit Dei adversum Ochoziam, ut veniret ad Ioram et, cum venisset, egrederetur cum eo adversum Iehu filium Namsi, quem unxit Dominus, ut deleret domum Achab.
2CHR|22|8|Cum ergo iudicium faceret Iehu in domum Achab, invenit principes Iudae et filios fratrum Ochoziae, qui ministrabant ei, et interfecit illos.
2CHR|22|9|Ipsumque perquisivit Ochoziam, et comprehenderunt eum latentem in Samaria; adductumque ad se Iehu occidit. Et sepelierunt eum, eo quod dicebant eum esse filium Iosaphat, qui quaesierat Dominum in toto corde suo.Nec erat aliquis de stirpe Ochoziae, qui posset regnare.
2CHR|22|10|Athalia autem mater eius videns quod mortuus esset filius suus surrexit et interfecit omnem stirpem regiam domus Iudae.
2CHR|22|11|Porro Iosabeth filia regis tulit Ioas filium Ochoziae et furata est eum de medio filiorum regis, cum interficerentur, absconditque cum nutrice sua in cubiculo lectulorum. Iosabeth autem, quae absconderat eum, erat filia regis Ioram, uxor Ioiadae pontificis, soror Ochoziae; et idcirco Athalia non interfecit eum.
2CHR|22|12|Fuit ergo cum eis in domo Dei absconditus sex annis, quibus regnavit Athalia super terram.
2CHR|23|1|Anno autem septimo confor tatus Ioiada assumpsit centu riones, Azariam videlicet filium Ieroham et Ismael filium Iohanan, Azariam quoque filium Obed et Maasiam filium Adaiae et Elisaphat filium Zechri, et iniit cum eis foedus.
2CHR|23|2|Qui circumeuntes Iudam congregaverunt Levitas de cunctis urbibus Iudae et principes familiarum Israel veneruntque in Ierusalem.
2CHR|23|3|Iniit igitur omnis congregatio pactum in domo Dei cum rege. Dixitque ad eos Ioiada: " Ecce filius regis regnabit, sicut locutus est Dominus super filios David.
2CHR|23|4|Hoc est ergo, quod facietis.
2CHR|23|5|Tertia pars vestrum, qui veniunt ad sabbatum sacerdotum et Levitarum et ianitorum, erit in portis, tertia vero pars ad domum regis et tertia in porta, quae appellatur Fundamenti; omne vero reliquum vulgus sit in atriis domus Domini.
2CHR|23|6|Nec quisquam alius ingrediatur domum Domini, nisi sacerdotes et qui ministrant de Levitis; ipsi tantummodo ingrediantur, quia sanctificati sunt. Et omne reliquum vulgus observet observationem Domini.
2CHR|23|7|Levitae autem circumdent regem habentes singuli arma sua in manu. Et si quis alius ingressus fuerit templum, interficiatur. Sintque cum rege et intrante et egrediente ".
2CHR|23|8|Fecerunt igitur Levitae et universus Iuda iuxta omnia, quae praeceperat Ioiada pontifex; et assumpserunt singuli viros suos, qui veniebant sabbato cum his, qui sabbato egressuri erant: siquidem Ioiada pontifex non dimisit abire turmas, quae sibi per singulas hebdomadas succedere consueverant.
2CHR|23|9|Deditque Ioiada sacerdos centurionibus lanceas clipeosque et peltas regis David, quae erant in domo Dei.
2CHR|23|10|Constituitque omnem populum tenentium tela a parte templi dextra usque ad partem templi sinistram coram altari et templo per circuitum regis.
2CHR|23|11|Et eduxerunt filium regis et dederunt ei diadema et testimonium et constituerunt eum regem. Unxerunt quoque illum Ioiada pontifex et filii eius; imprecatique sunt ei atque dixerunt: " Vivat rex! ".
2CHR|23|12|Quod cum audisset Athalia, vocem scilicet currentium atque laudantium regem, ingressa est ad populum in templum Domini.
2CHR|23|13|Cumque vidisset regem stantem super gradum suum in introitu et principes tubasque circa eum omnemque populum terrae gaudentem atque clangentem tubis cantoresque cum diversi generis organis signum dantes ad laudandum, scidit vestimenta sua et ait: " Coniuratio, coniuratio! ".
2CHR|23|14|Praecepit autem Ioiada pontifex centurionibus, qui erant super exercitum, dicens: " Educite illam extra saepta templi! Qui autem sequetur eam, interficiatur foris gladio! ". Dixerat enim sacerdos: " Non occidetis eam in domo Domini! ".
2CHR|23|15|Et imposuerunt ei manus; cumque intrasset portam Equorum domus regis, interfecerunt eam ibi.
2CHR|23|16|Pepigit autem Ioiada foedus inter se universumque populum et regem, ut esset populus Domini.
2CHR|23|17|Itaque ingressus est omnis populus domum Baal et destruxerunt eam et altaria ac simulacra illius confregerunt; Matthan quoque sacerdotem Baal interfecerunt ante aras.
2CHR|23|18|Constituit autem Ioiada praepositos in domo Domini sub manibus sacerdotum et Levitarum, quos distribuit David in domo Domini, ut offerrent holocausta Domino, sicut scriptum est in lege Moysi, in gaudio et canticis iuxta dispositionem David.
2CHR|23|19|Constituit quoque ianitores in portis domus Domini, ut non ingrederetur eam immundus in omni re.
2CHR|23|20|Assumpsitque centuriones et fortissimos viros ac principes populi et omne vulgus terrae, et fecerunt descendere regem de domo Domini et introire per medium portae Superioris in domum regis et collocaverunt eum in solio regali.
2CHR|23|21|Laetatusque est omnis populus terrae, et urbs quievit; porro Athalia interfecta est gladio.
2CHR|24|1|Septem annorum erat Ioas, cum regnare coepisset, et quadraginta annis regnavit in Ierusalem. Nomen matris eius Sebia de Bersabee.
2CHR|24|2|Fecitque, quod bonum est coram Domino, cunctis diebus Ioiadae sacerdotis.
2CHR|24|3|Accepit autem ei Ioiada uxores duas, e quibus genuit filios et filias.
2CHR|24|4|Post quae placuit Ioas, ut instauraret domum Domini.
2CHR|24|5|Congregavitque sacerdotes et Levitas et dixit eis: " Egredimini ad civitates Iudae et colligite de universo Israel pecuniam ad sartatecta templi Dei vestri per singulos annos. Festinatoque hoc facite ". Porro Levitae non festinarunt.
2CHR|24|6|Vocavitque rex Ioiadam principem et dixit ei: " Quare non tibi fuit curae, ut cogeres Levitas inferre de Iuda et de Ierusalem pecuniam, quae constituta est a Moyse servo Domini, ut inferret eam omnis congregatio Israel in tabernaculum testimonii?
2CHR|24|7|Athalia enim impiissima et filii eius dissipaverunt domum Dei et de universis, quae sanctificata fuerant templo Domini, dedicaverunt Baalim ".
2CHR|24|8|Praecepit ergo rex, et fecerunt arcam posueruntque eam iuxta portam domus Domini forinsecus.
2CHR|24|9|Et praedicatum est in Iuda et Ierusalem, ut deferrent singuli pretium Domino, quod constituit Moyses servus Dei super Israel in deserto.
2CHR|24|10|Laetatique sunt cuncti principes et omnis populus et ingressi contulerunt in arcam atque miserunt ita, ut impleretur.
2CHR|24|11|Cumque tempus esset, ut deferrent arcam ad magistratus regis per manus Levitarum, et viderent multam esse pecuniam, ingrediebatur scriba regis et quem primus sacerdos constituerat, effundebantque pecuniam, quae erat in arca; porro arcam reportabant ad locum suum. Sicque faciebant per singula tempora, et congregata est infinita pecunia,
2CHR|24|12|quam dederunt rex et Ioiada his, qui praeerant operibus domus Domini. At illi conducebant ex ea caesores lapidum et artifices operum singulorum, ut instaurarent domum Domini, fabros quoque ferri et aeris, ut domus Dei fulciretur.
2CHR|24|13|Egeruntque operarii, et obducebatur cicatrix operi per manus eorum, ac suscitaverunt domum Domini in statum pristinum et firme eam stare fecerunt.
2CHR|24|14|Cumque haec complessent, detulerunt coram rege et Ioiada reliquam partem pecuniae, de qua facta sunt vasa templi in ministerium et ad holocausta, phialae quoque et cetera vasa aurea et argentea. Et offerebantur holocausta in domo Domini iugiter cunctis diebus Ioiadae.
2CHR|24|15|Senuit autem Ioiada plenus dierum et mortuus est cum centum triginta esset annorum.
2CHR|24|16|Sepelieruntque eum in civitate David cum regibus, eo quod fecisset bonum in Israel cum Deo et cum domo eius.
2CHR|24|17|Postquam autem obiit Ioiada, ingressi sunt principes Iudae et adoraverunt regem, qui delinitus obsequiis eorum acquievit eis.
2CHR|24|18|Et dereliquerunt templum Domini, Dei patrum suorum, servieruntque palis et sculptilibus, et facta est ira contra Iudam et Ierusalem propter hoc peccatum.
2CHR|24|19|Mittebatque eis prophetas, ut reverterentur ad Dominum, quos protestantes illi audire nolebant.
2CHR|24|20|Spiritus itaque Dei induit Zachariam filium Ioiadae sacerdotis; et stetit in conspectu populi et dixit eis: " Haec dicit Deus: Quare transgredimini praecepta Domini, quod vobis non proderit? Quia dereliquistis Dominum, ipse dereliquit vos ".
2CHR|24|21|Qui coniuraverunt adversus eum et lapidaverunt eum iuxta regis imperium in atrio domus Domini.
2CHR|24|22|Et non est recordatus Ioas rex misericordiae, quam fecerat Ioiada pater illius secum, sed interfecit filium eius. Qui cum moreretur, ait: " Videat Dominus et requirat! ".
2CHR|24|23|Cumque evolutus esset annus, ascendit contra eum exercitus Syriae venitque in Iudam et Ierusalem et exterminaverunt cunctos principes populi atque universam praedam miserunt regi Damascum.
2CHR|24|24|Et certe, cum permodicus venisset numerus Syrorum, tradidit Dominus manibus eorum exercitum magnum valde, eo quod reliquissent Dominum, Deum patrum suorum; in Ioas quoque ignominiosa exercuere iudicia.
2CHR|24|25|Et abeuntes dimiserunt eum in languoribus magnis. Coniuraverunt autem contra eum servi sui in ultionem sanguinis filii Ioiadae sacerdotis et occiderunt eum in lectulo suo, et mortuus est. Sepelieruntque eum in civitate David, sed non in sepulcris regum.
2CHR|24|26|Insidiati vero sunt ei Zabad filius Semath Ammanitidis et Iozabad filius Semarith Moabitidis.
2CHR|24|27|Porro de filiis eius, de summa tributi, quod impositum fuerat sub eo, et de instauratione domus Dei scriptum est in commentariis libri regum. Regnavitque Amasias filius eius pro eo.
2CHR|25|1|Viginti quinque annorum erat Amasias, cum regnare coepisset, et viginti novem annis regnavit in Ierusalem. Nomen matris eius Ioaden de Ierusalem.
2CHR|25|2|Fecitque bonum in conspectu Domini, verumtamen non in corde perfecto.
2CHR|25|3|Cumque roboratum sibi videret imperium, iugulavit servos suos, qui occiderant regem patrem suum,
2CHR|25|4|sed filios eorum non interfecit, sicut scriptum est in libro legis Moysi, ubi praecepit Dominus dicens: " Non occidentur patres pro filiis, neque filii pro patribus suis, sed unusquisque in suo peccato morietur ".
2CHR|25|5|Congregavit igitur Amasias Iudam et constituit eos per familias tribunosque et centuriones in universo Iuda et Beniamin. Et recensuit a viginti annis sursum invenitque trecenta milia iuvenum, qui egrederentur ad pugnam et tenerent hastam et clipeum.
2CHR|25|6|Mercede quoque conduxit de Israel centum milia robustorum centum talentis argenti.
2CHR|25|7|Venit autem homo Dei ad illum et ait: " O rex, ne egrediatur tecum exercitus Israel; non est enim Dominus cum Israel, cunctis filiis Ephraim.
2CHR|25|8|Quod si putas in robore exercitus bella consistere, superari te faciet Deus ab hostibus: Dei quippe est et adiuvare et in fugam vertere ".
2CHR|25|9|Dixitque Amasias ad hominem Dei: " Quid ergo fiet de centum talentis, quae dedi militibus Israel? ". Et respondit ei homo Dei: " Habet Dominus, unde tibi dare possit multo his plura ".
2CHR|25|10|Separavit itaque Amasias exercitum, qui venerat ad eum ex Ephraim, ut reverteretur in locum suum; at illi contra Iudam vehementer irati reversi sunt in regionem suam.
2CHR|25|11|Porro Amasias confidenter eduxit populum suum et abiit in vallem Salinarum percussitque filios Seir decem milia.
2CHR|25|12|Et alia decem milia virorum ceperunt filii Iudae et adduxerunt ad praeruptum cuiusdam petrae praecipitaveruntque eos de summo in praeceps, qui universi crepuerunt.
2CHR|25|13|At ille exercitus, quem remiserat Amasias, ne secum iret ad proelium, diffusus est in civitatibus Iudae a Samaria usque Bethoron et, interfectis tribus milibus, diripuit praedam magnam.
2CHR|25|14|Amasias vero, post caedem Idumaeorum et allatos deos filiorum Seir, statuit illos in deos sibi et adorabat eos et illis adolebat.
2CHR|25|15|Quam ob rem iratus Dominus contra Amasiam misit ad illum prophetam, qui diceret ei: " Cur adorasti deos, qui non liberaverunt populum suum de manu tua? ".
2CHR|25|16|Cumque haec ille loqueretur, respondit ei: " Num consiliarium regis fecimus te? Quiesce! Cur interficiam te? ". Discedensque propheta: " Sed scio, inquit, quod decrevit Deus occidere te, quia fecisti hoc et non acquievisti consilio meo ".
2CHR|25|17|Igitur Amasias rex Iudae, inito consilio, misit ad Ioas filium Ioachaz filii Iehu regem Israel dicens: " Veni, videamus nos mutuo! ".
2CHR|25|18|At ille remisit nuntium dicens: " Carduus, qui est in Libano, misit ad cedrum Libani dicens: "Da filiam tuam filio meo uxorem". Et ecce bestiae agri, quae erant in Libano, transierunt et conculcaverunt carduum.
2CHR|25|19|Dixisti: "Percussi Edom!". Et idcirco erigitur cor tuum in superbiam. Sede in domo tua! Cur malum adversum te provocas, ut cadas et tu et Iuda tecum? ".
2CHR|25|20|Noluit audire Amasias, eo quod Domini esset voluntas, ut traderetur in manibus hostium propter cultum deorum Edom.
2CHR|25|21|Ascendit igitur Ioas rex Israel, et mutuos sibi praebuere conspectus: ipse et Amasias rex Iudae in Bethsames Iudae.
2CHR|25|22|Corruitque Iuda coram Israel et fugit in tabernacula sua.
2CHR|25|23|Porro Amasiam regem Iudae filium Ioas filii Ioachaz cepit Ioas rex Israel in Bethsames et adduxit in Ierusalem destruxitque murum eius a porta Ephraim usque ad portam Anguli quadringentis cubitis.
2CHR|25|24|Omne quoque aurum et argentum et universa vasa, quae repererat in domo Dei et apud Obededom in thesauris etiam domus regiae, necnon et obsides reduxit Samariam.
2CHR|25|25|Vixit autem Amasias filius Ioas rex Iudae, postquam mortuus est Ioas filius Ioachaz rex Israel, quindecim annis.
2CHR|25|26|Reliqua vero gestorum Amasiae priorum et novissimorum scripta sunt in libro regum Iudae et Israel.
2CHR|25|27|Qui postquam recessit a Domino, tetenderunt ei insidias in Ierusalem; cumque fugisset Lachis, miserunt post eum in Lachis et interfecerunt eum ibi.
2CHR|25|28|Reportantesque super equos sepelierunt eum cum patribus suis in civitate David.
2CHR|26|1|Omnis autem populus Iudae Oziam annorum sedecim constituit regem pro patre suo Amasia.
2CHR|26|2|Ipse reaedificavit Ailath et restituit eam dicioni Iudae, postquam dormivit rex cum patribus suis.
2CHR|26|3|Sedecim annorum erat Ozias, cum regnare coepisset, et quinquaginta duobus annis regnavit in Ierusalem. Nomen matris eius Iechelia de Ierusalem.
2CHR|26|4|Fecitque, quod erat rectum in oculis Domini iuxta omnia, quae fecerat Amasias pater eius.
2CHR|26|5|Et exquisivit Deum in diebus Zachariae, qui erudivit eum in timore Dei; et quamdiu requirebat Dominum, eum prosperari fecit Deus.
2CHR|26|6|Denique egressus est et pugnavit contra Philisthim et destruxit murum Geth et murum Iabniae murumque Azoti. Aedificavit quoque oppida in regione Azoti et Philisthim.
2CHR|26|7|Et adiuvit eum Deus contra Philisthim et contra Arabas, qui habitabant in Gurbaal, et contra Meunitas.
2CHR|26|8|Pendebantque Ammonitae munera Oziae; et divulgatum est nomen eius usque ad introitum Aegypti, quia confortatus est in excelsum.
2CHR|26|9|Aedificavitque Ozias turres in Ierusalem super portam Anguli et super portam Vallis et super Angulum firmavitque eas.
2CHR|26|10|Exstruxit etiam turres in solitudine et fodit cisternas plurimas, eo quod haberet multa pecora tam in Sephela quam in planitie; agricolas quoque habuit et vinitores in montibus et in campis fertilibus; erat quippe homo agriculturae deditus.
2CHR|26|11|Fuit autem exercitus bellatorum eius, qui procedebant ad proelia in turmis secundum numerum census per manum Iehiel scribae Maasiaeque praefecti sub manu Hananiae, qui erat de ducibus regis.
2CHR|26|12|Omnisque numerus principum per familias virorum fortium duorum milium sescentorum.
2CHR|26|13|Et sub eis universus exercitus trecentorum et septem milium quingentorum, qui erant apti ad bella, ut pro rege contra adversarios dimicarent.
2CHR|26|14|Praeparavit quoque eis Ozias, id est cuncto exercitui, clipeos et hastas et galeas et loricas arcusque et fundas ad iaciendos lapides.
2CHR|26|15|Et fecit in Ierusalem machinas excogitatas arte, quas in turribus collocavit et in angulis murorum, ut mitterent sagittas et saxa grandia; egressumque est nomen eius procul, eo quod mirabiliter auxiliaretur ei Dominus et corroborasset illum.
2CHR|26|16|Sed, cum roboratus esset, elevatum est cor eius in interitum suum, et deliquit contra Dominum Deum suum; ingressusque templum Domini adolere voluit incensum super altare thymiamatis.
2CHR|26|17|Statimque ingressus post eum Azarias sacerdos et cum eo sacerdotes Domini octoginta viri fortissimi;
2CHR|26|18|restiterunt regi atque dixerunt: " Non est tui officii, Ozia, ut adoleas incensum Domino, sed sacerdotum, hoc est filiorum Aaron, qui consecrati sunt ad huiuscemodi ministerium. Egredere de sanctuario, quia praevaricatus es; et non reputabitur tibi in gloriam hoc a Domino Deo ".
2CHR|26|19|Iratusque est Ozias et tenens in manu turibulum, ut adoleret incensum, minabatur sacerdotibus. Statimque orta est lepra in fronte eius coram sacerdotibus in domo Domini super altare thymiamatis.
2CHR|26|20|Cumque respexisset eum Azarias pontifex et omnes reliqui sacerdotes, viderunt lepram in fronte eius et festinato expulerunt eum; sed et ipse acceleravit egredi, eo quod malo afflixisset eum Dominus.
2CHR|26|21|Fuit igitur Ozias rex leprosus usque ad diem mortis suae et habitavit in domo separata plenus lepra, eo quod abscissus fuerat de domo Domini. Porro Ioatham filius eius rexit domum regis et iudicabat populum terrae.
2CHR|26|22|Reliqua autem gestorum Oziae priorum et novissimorum scripsit Isaias filius Amos propheta.
2CHR|26|23|Dormivitque Ozias cum patribus suis, et sepelierunt eum in agro regalium sepulcrorum, eo quod dicebant: " Erat leprosus ". Regnavitque Ioatham filius eius pro eo.
2CHR|27|1|Viginti quinque annorum erat Ioatham, cum regnare coepisset, et sedecim annis regnavit in Ierusalem. Nomen matris eius Ierusa filia Sadoc.
2CHR|27|2|Fecitque, quod rectum erat coram Domino iuxta omnia, quae fecerat Ozias pater suus, excepto quod non est ingressus templum Domini, et adhuc populus delinquebat.
2CHR|27|3|Ipse aedificavit portam domus Domini Superiorem et in muro Ophel multa construxit.
2CHR|27|4|Urbes quoque aedificavit in montibus Iudae et in saltibus castella et turres.
2CHR|27|5|Ipse pugnavit contra regem filiorum Ammon et vicit eos, dederuntque ei filii Ammon in anno illo centum talenta argenti et decem milia choros tritici ac totidem choros hordei; haec ei praebuerunt filii Ammon etiam in anno secundo et tertio.
2CHR|27|6|Corroboratusque est Ioatham, eo quod direxisset vias suas coram Domino Deo suo.
2CHR|27|7|Reliqua autem gestorum Ioatham et omnes pugnae eius et viae scriptae sunt in libro regum Israel et Iudae.
2CHR|27|8|Viginti quinque annorum erat, cum regnare coepisset, et sedecim annis regnavit in Ierusalem.
2CHR|27|9|Dormivitque Ioatham cum patribus suis, et sepelierunt eum in civitate David; et regnavit Achaz filius eius pro eo.
2CHR|28|1|Viginti annorum erat Achaz, cum regnare coepis set, et sedecim annis regnavit in Ierusalem. Non fecit rectum in conspectu Domini sicut David pater eius,
2CHR|28|2|sed ambulavit in viis regum Israel. Insuper et simulacra fudit Baalim.
2CHR|28|3|Ipse est, qui adolevit in valle filii Ennom et lustravit filios suos in igne iuxta abominationes gentium, quas expulit Dominus coram filiis Israel.
2CHR|28|4|Sacrificabat quoque et thymiama succendebat in excelsis et in collibus et sub omni ligno frondoso.
2CHR|28|5|Tradiditque eum Dominus Deus eius in manu regis Syriae, qui percussit eum multosque captivos de eo cepit et adduxit in Damascum. Manibus quoque regis Israel traditus est et percussus plaga grandi.
2CHR|28|6|Occidit enim Phacee filius Romeliae de Iuda centum viginti milia in die uno, omnes viros bellatores, eo quod reliquissent Dominum, Deum patrum suorum.
2CHR|28|7|Eodem tempore occidit Zechri vir potens ex Ephraim Maasiam filium regis et Ezricam praefectum domus, Elcanam quoque secundum a rege.
2CHR|28|8|Ceperuntque filii Israel de fratribus suis ducenta milia mulierum, puerorum et puellarum, et infinitam praedam pertuleruntque eam in Samariam.
2CHR|28|9|Erat autem ibi propheta Domini nomine Oded, qui egressus obviam exercitui venienti in Samariam dixit eis: " Ecce, iratus Dominus, Deus patrum vestrorum, contra Iudam tradidit eos in manibus vestris, et occidistis eos atrociter, ita ut ad caelum pertingeret vestra crudelitas.
2CHR|28|10|Insuper filios Iudae et Ierusalem vultis vobis subicere in servos et ancillas. Attamen nonne vos ipsi estis in culpa coram Domino Deo vestro?
2CHR|28|11|Audite ergo consilium meum et reducite captivos, quos adduxistis de fratribus vestris, quia magnus furor Domini imminet vobis ".
2CHR|28|12|Steterunt itaque viri de principibus filiorum Ephraim, Azarias filius Iohanan, Barachias filius Mosollamoth, Ezechias filius Sellum et Amasa filius Adali, contra eos, qui veniebant de proelio,
2CHR|28|13|et dixerunt eis: " Non introducetis huc captivos, quia ad culpam coram Domino, quae iam est super nos, vultis adicere super peccata nostra et culpam nostram. Grandis quippe culpa est nobis, et ira furoris Domini super Israel ".
2CHR|28|14|Dimiseruntque viri bellatores captivos et universa, quae ceperant, coram principibus et omni multitudine.
2CHR|28|15|Et surrexerunt viri nominatim designati et confortaverunt captivos omnesque, qui nudi erant, vestierunt de spoliis. Cumque vestissent eos et calceassent et refecissent cibo ac potu unxissentque, deduxerunt eos sollicite, et quidem omnes vacillantes in iumentis, et adduxerunt Iericho civitatem Palmarum ad fratres eorum. Ipsique reversi sunt Samariam.
2CHR|28|16|Tempore illo misit rex Achaz ad regem Assyriorum auxilium postulans.
2CHR|28|17|Venerunt enim et Idumaei et percusserunt Iudam et ceperunt captivos.
2CHR|28|18|Philisthim quoque diffusi sunt per urbes Sephelae et Nageb Iudae ceperuntque Bethsames et Aialon et Gederoth, Socho quoque cum viculis eius et Thamnan et Gamzo cum viculis earum et habitaverunt in eis.
2CHR|28|19|Humiliaverat enim Dominus Iudam propter Achaz regem Israel, eo quod relaxasset ei frenum et contemptui habuisset Dominum.
2CHR|28|20|Venitque contra eum Theglathphalasar rex Assyriorum, qui afflixit eum, non autem confortavit.
2CHR|28|21|Achaz enim, spoliata domo Domini et domo regis et principum, dedit regi Assyriorum munera, et tamen nihil ei profuit.
2CHR|28|22|Insuper et in tempore angustiae suae auxit contemptum in Dominum. Ipse rex Achaz
2CHR|28|23|immolavit diis Damasci victimas percussoribus suis et dixit: " Dii regum Syriae auxiliantur eis; quos ego placabo hostiis, et aderunt mihi ", cum e contrario ipsi fuerint ruina ei et universo Israel.
2CHR|28|24|Direptis itaque Achaz omnibus vasis domus Dei atque confractis, clausit ianuas templi Dei et fecit sibi altaria in universis angulis Ierusalem.
2CHR|28|25|In singulis quoque urbibus Iudae exstruxit excelsa ad adolendum diis alienis atque ad iracundiam provocavit Dominum, Deum patrum suorum.
2CHR|28|26|Reliqua autem gestorum eius et omnium operum suorum priorum et novissimorum scripta sunt in libro regum Iudae et Israel.
2CHR|28|27|Dormivitque Achaz cum patribus suis, et sepelierunt eum in civitate Ierusalem; non autem posuerunt eum in sepulcra regum Israel. Regnavitque Ezechias filius eius pro eo.
2CHR|29|1|Igitur Ezechias regnare coepit, cum viginti quinque esset annorum, et viginti novem annis regnavit in Ierusalem. Nomen matris eius Abi filia Zachariae.
2CHR|29|2|Fecitque, quod erat placitum in conspectu Domini, iuxta omnia, quae fecerat David pater eius.
2CHR|29|3|Ipse anno et mense primo regni sui aperuit valvas domus Domini et instauravit eas.
2CHR|29|4|Adduxitque sacerdotes atque Levitas et congregavit eos in plateam orientalem
2CHR|29|5|dixitque ad eos: " Audite me, Levitae! Nunc sanctificamini; mundate domum Domini, Dei patrum vestrorum, et auferte omnem immunditiam de sanctuario.
2CHR|29|6|Peccaverunt patres nostri et fecerunt malum in conspectu Domini Dei nostri derelinquentes eum; averterunt facies suas a tabernaculo Domini et praebuerunt dorsum.
2CHR|29|7|Insuper clauserunt ostia, quae erant in porticu, et exstinxerunt lucernas incensumque non adoleverunt et holocausta non obtulerunt in sanctuario Deo Israel.
2CHR|29|8|Concitatus est itaque furor Domini super Iudam et Ierusalem; tradiditque eos in commotionem et in stuporem et in sibilum, sicut ipsi cernitis oculis vestris.
2CHR|29|9|En, corruerunt patres nostri gladiis, filii nostri et filiae nostrae et coniuges captivae ductae sunt propter hoc scelus.
2CHR|29|10|Nunc igitur placet mihi, ut ineam foedus cum Domino, Deo Israel, et avertat a nobis furorem irae suae.
2CHR|29|11|Filii mei, nolite neglegere; vos enim elegit Dominus, ut stetis coram eo et ministretis illi colatisque eum et adoleatis ".
2CHR|29|12|Surrexerunt ergo Levitae, Mahath filius Amasai et Ioel filius Azariae de filiis Caath; porro de filiis Merari Cis filius Abdi et Azarias filius Iallelel; de filiis autem Gerson Ioah filius Zimma et Eden filius Ioah;
2CHR|29|13|at vero de filiis Elisaphan Semri et Iehiel; de filiis quoque Asaph Zacharias et Matthanias;
2CHR|29|14|necnon de filiis Heman Iahiel et Semei; sed et de filiis Idithun Semeias et Oziel.
2CHR|29|15|Congregaveruntque fratres suos et sanctificati sunt et ingressi iuxta mandatum regis et imperium Domini, ut expiarent domum Dei.
2CHR|29|16|Sacerdotes quoque ingressi intra templum Domini, ut mundarent illud, extulerunt omnem immunditiam, quam intro reppererant in vestibulum domus Domini, quam tulerunt Levitae et asportaverunt ad torrentem Cedron foras.
2CHR|29|17|Coeperunt autem prima die mensis primi sanctificare et in die octava eiusdem mensis ingressi sunt porticum templi Domini et sanctificaverunt templum Domini diebus octo; et in die sexta decima mensis eiusdem, quod coeperant, impleverunt.
2CHR|29|18|Ingressi quoque sunt ad Ezechiam regem et dixerunt ei: " Mundavimus omnem domum Domini et altare holocausti vasaque eius necnon et mensam propositionis cum omnibus vasis suis
2CHR|29|19|cunctamque templi supellectilem, quam removerat rex Achaz in regno suo in praevaricatione sua, restituimus et sanctificavimus. Ecce exposita sunt omnia coram altari Domini ".
2CHR|29|20|Consurgensque diluculo Ezechias rex adunavit principes civitatis et ascendit domum Domini.
2CHR|29|21|Attuleruntque simul tauros septem, arietes septem, agnos septem et hircos septem pro peccato, pro regno, pro sanctuario, pro Iuda; dixit quoque sacerdotibus filiis Aaron, ut offerrent super altare Domini.
2CHR|29|22|Mactaverunt igitur tauros et susceperunt sacerdotes sanguinem et fuderunt illum super altare; mactaverunt etiam arietes et illorum sanguinem super altare fuderunt; immolaverunt agnos et fuderunt super altare sanguinem.
2CHR|29|23|Applicaverunt hircos pro peccato coram rege et universa multitudine imposueruntque manus suas super eos,
2CHR|29|24|et immolaverunt illos sacerdotes et asperserunt sanguinem eorum super altare pro piaculo universi Israelis; pro omni quippe Israel praeceperat rex, ut holocaustum fieret et pro peccato.
2CHR|29|25|Constituit quoque Levitas in domo Domini cum cymbalis et psalteriis et citharis secundum dispositionem David et Gad videntis regis et Nathan prophetae; siquidem Domini praeceptum fuit per manum prophetarum eius.
2CHR|29|26|Steteruntque Levitae tenentes organa David, et sacerdotes tubas.
2CHR|29|27|Et iussit Ezechias, ut offerrent holocaustum super altare; cumque offerretur holocaustum, coeperunt laudes canere Domino et clangere tubis atque in diversis organis David regis Israel concrepare.
2CHR|29|28|Omni autem turba adorante, cantores et ii, qui tenebant tubas, erant in officio suo, donec compleretur holocaustum.
2CHR|29|29|Cumque finita esset oblatio, incurvatus est rex et omnes, qui erant cum eo, et adoraverunt.
2CHR|29|30|Praecepitque Ezechias et principes Levitis, ut laudarent Dominum verbis David et Asaph videntis; qui laudaverunt eum magna laetitia et curvato genu adoraverunt.
2CHR|29|31|Ezechias autem etiam haec addidit: " Nunc, impletis manibus vestris Domino, accedite et afferte victimas et sacrificia pro gratiarum actione in domo Domini ". Attulit ergo universa multitudo hostias et sacrificia pro gratiarum actione, et omnis voluntarius et proni animi holocausta.
2CHR|29|32|Porro numerus holocaustorum, quae attulit multitudo, hic fuit: tauros septuaginta, arietes centum, agnos ducentos, in holocaustum Domino omnia haec.
2CHR|29|33|Sanctificaveruntque Domino boves sescentos et oves tria milia.
2CHR|29|34|Sacerdotes vero pauci erant nec poterant sufficere, ut pelles holocaustorum detraherent; unde et Levitae fratres eorum adiuverunt eos, donec impleretur opus, et sanctificarentur sacerdotes; Levitae quippe recti corde, ut sanctificarentur magis quam sacerdotes.
2CHR|29|35|Fuerunt igitur holocausta plurima, adipes pacificorum et libamina, quae pertinebant ad holocausta.Restitutus est ita cultus domus Domini.
2CHR|29|36|Laetatusque est Ezechias et omnis populus de eo, quod paravit Dominus populo; repente quippe hoc factum est.
2CHR|30|1|Misit quoque Ezechias ad omnem Israel et Iudam scri psitque et epistulas ad Ephraim et Manassen, ut venirent ad domum Domini in Ierusalem et facerent Pascha Domino, Deo Israel.
2CHR|30|2|Inito quoque consilio regis et principum et universi coetus in Ierusalem, decreverunt, ut facerent Pascha mense secundo.
2CHR|30|3|Non enim potuerant facere in tempore suo, quia sacerdotes, qui possent sufficere, sanctificati non fuerant, et populus necdum congregatus erat in Ierusalem.
2CHR|30|4|Placuit ergo sermo regi et omni multitudini,
2CHR|30|5|et decreverunt, ut mitterent nuntios in universum Israel de Bersabee usque Dan, ut venirent et facerent Pascha Domino, Deo Israel, in Ierusalem; in plurima enim multitudine non fecerant, sicut lege praescriptum est.
2CHR|30|6|Perrexeruntque cursores cum epistulis ex regis manu et principum eius in universum Israel et Iudam, iuxta quod rex iusserat, praedicantes: " Filii Israel, revertimini ad Dominum, Deum Abraham et Isaac et Israel, ut revertatur ad reliquias, quae effugerunt manum regum Assyriorum.
2CHR|30|7|Nolite fieri sicut patres vestri et fratres, qui recesserunt a Domino, Deo patrum suorum, et tradidit eos in interitum, ut ipsi cernitis.
2CHR|30|8|Nolite nunc indurare cervices vestras sicut patres vestri. Tradite manus Domino et venite ad sanctuarium eius, quod sanctificavit in aeternum; servite Domino Deo vestro, ut avertatur a vobis ira furoris eius.
2CHR|30|9|Si enim vos reversi fueritis ad Dominum, fratres vestri et filii habebunt misericordiam coram dominis suis, qui illos duxere captivos, et revertentur in terram hanc: misericors enim et clemens est Dominus Deus vester et non avertet faciem suam a vobis, si reversi fueritis ad eum ".
2CHR|30|10|Igitur cursores pergebant de civitate in civitatem per terram Ephraim et Manasse usque Zabulon, illis irridentibus et subsannantibus eos.
2CHR|30|11|Attamen quidam viri ex Aser et Manasse et Zabulon se humiliaverunt et venerunt Ierusalem.
2CHR|30|12|In Iuda quoque facta est manus Domini, ut daret eis cor unum, ut facerent praeceptum regis et principum iuxta verbum Domini.
2CHR|30|13|Congregatus est ergo in Ierusalem populus multus, ut faceret sollemnitatem Azymorum in mense secundo, ecclesia magna valde.
2CHR|30|14|Et surgentes destruxerunt altaria, quae erant in Ierusalem, atque universa thymiamateria subvertentes proiecerunt in torrentem Cedron.
2CHR|30|15|Et mactaverunt Pascha quarta decima die mensis secundi; sacerdotes autem atque Levitae confusi sanctificati sunt et attulerunt holocausta in domum Domini.
2CHR|30|16|Steteruntque in ordine suo iuxta dispositionem et legem Moysi hominis Dei, sacerdotes vero suscipiebant effundendum sanguinem de manibus Levitarum,
2CHR|30|17|eo quod multi in coetu sanctificati non essent; idcirco Levitae mactaverunt victimas Paschae omnibus, qui non erant mundi, ut sanctificarent illas Domino.
2CHR|30|18|Valde magna enim pars populi, de Ephraim et Manasse et Issachar et Zabulon, non erant mundati; et comederunt Pascha non iuxta, quod scriptum est. Et oravit pro eis Eze chias dicens: " Dominus bonus propitietur
2CHR|30|19|cunctis, qui direxerunt cor suum, ut requirerent Dominum, Deum patrum suorum, quamvis non secundum munditiam sanctuarii ".
2CHR|30|20|Quem exaudivit Dominus, et placatus est populo.
2CHR|30|21|Feceruntque filii Israel, qui inventi sunt in Ierusalem, sollemnitatem Azymorum septem diebus in laetitia magna, laudaverunt Dominum et per singulos dies Levitae et sacerdotes per organa benesonantia.
2CHR|30|22|Et locutus est Ezechias ad cor omnium Levitarum, qui habebant intellegentiam bonam super Domino; et compleverunt sollemnitatem septem dierum immolantes victimas pacificorum et laudantes Dominum, Deum patrum suorum.
2CHR|30|23|Placuitque universae multitudini, ut celebrarent etiam alios dies septem, quod et fecerunt cum ingenti gaudio.
2CHR|30|24|Ezechias enim rex Iudae praebuerat multitudini mille tauros et septem milia ovium; principes vero dederant populo tauros mille et oves decem milia; sanctificata est ergo sacerdotum plurima multitudo.
2CHR|30|25|Et hilaritate perfusa est omnis turba Iudae, tam sacerdotum et Levitarum quam universae frequentiae, quae venerat ex Israel, advenae quoque, qui venerant de terra Israel vel habitabant in Iuda.
2CHR|30|26|Factaque est grandis laetitia in Ierusalem, qualis a diebus Salomonis filii David regis Israel in ea urbe non fuerat.
2CHR|30|27|Surrexerunt autem sacerdotes levitici generis benedicentes populo; et exaudita est vox eorum, pervenitque oratio eorum in habitaculum sanctum eius in caelum.
2CHR|31|1|Cumque haec fuissent rite celebrata, egressus est omnis Israel, qui inventus fuerat in urbibus Iudae, et fregerunt simulacra succideruntque palos, demoliti sunt excelsa et altaria destruxerunt non solum de universo Iuda et Beniamin, sed et de Ephraim quoque et Manasse, donec penitus everterent. Reversique sunt omnes filii Israel in possessiones et civitates suas.
2CHR|31|2|Ezechias autem constituit turmas sacerdotales et leviticas per divisiones suas, unumquemque in officio proprio tam sacerdotum videlicet quam Levitarum, ad holocausta et pacifica, ut ministrarent et confiterentur canerentque laudes in portis castrorum Domini.
2CHR|31|3|Pars autem regis erat, ut de propria eius substantia offerretur holocaustum mane semper et vespere, sabbatis quoque et calendis et sollemnitatibus ceteris, sicut scriptum est in lege Moysi.
2CHR|31|4|Praecepit etiam populo habitanti Ierusalem, ut darent partes sacerdotibus et Levitis, ut possent vacare legi Domini.
2CHR|31|5|Quod cum percrebruisset in auribus multitudinis, plurimas obtulere primitias filii Israel frumenti, vini et olei, mellis quoque et omnium, quae gignit humus, et decimas obtulerunt de omnibus abundanter.
2CHR|31|6|Sed et filii Israel et Iudae, qui habitabant in urbibus Iudae, obtulerunt decimas boum et ovium decimasque sanctorum, quae sanctificabant Domino Deo suo; atque universa portantes fecerunt acervos plurimos.
2CHR|31|7|Mense tertio coeperunt acervorum iacere fundamenta et mense septimo compleverunt eos.
2CHR|31|8|Cumque ingressi fuissent Ezechias et principes, viderunt acervos et benedixerunt Domino ac populo Israel.
2CHR|31|9|Interrogavitque Ezechias sacerdotes et Levitas, cur ita iacerent acervi.
2CHR|31|10|Respondit illi Azarias sacerdos primus de stirpe Sadoc dicens: " Ex quo coeperunt offerre donationem in domum Domini, comedimus et saturati sumus, et remanserunt plurima, eo quod benedixerit Dominus populo suo; reliquiarum autem copia est ista, quam cernis ".
2CHR|31|11|Praecepit igitur Ezechias, ut praepararent cellas in domo Domini. Quod cum fecissent,
2CHR|31|12|intulerunt tam donationem quam decimas et quaecumque sanctificaverant fideliter. Fuit autem praefectus eorum Chonenias Levita et Semei frater eius secundus,
2CHR|31|13|post quem Iahiel et Azazias et Nahath et Asael et Ierimoth, Iozabad quoque et Eliel et Iesmachias et Mahath et Banaias praepositi sub manibus Choneniae et Semei fratris eius ex imperio Ezechiae regis et Azariae pontificis domus Dei.
2CHR|31|14|Core vero filius Iemna Levites et ianitor orientalis portae praepositus erat iis, quae sponte offerebantur Domino, ad distribuendum donationem Domini et sanctissima.
2CHR|31|15|Et sub cura eius Eden et Beniamin, Iesua et Semeias, Amarias quoque et Sechenias in civitatibus sacerdotum, ut fideliter distribuerent fratribus suis tam maioribus quam minoribus in divisionibus suis,
2CHR|31|16|dummodo recensiti essent mares ab annis tribus et supra, cuncti qui ingrediebantur templum Domini, ut singulorum dierum ministeria observarent iuxta divisiones suas.
2CHR|31|17|Sacerdotes recensiti erant per familias, et Levitae a vicesimo anno et supra per ministeria et turmas suas.
2CHR|31|18|Et recensita erat universa familia omnis turmae, tam pro uxoribus quam liberis eorum utriusque sexus, quia in fidelitate servitii ipsorum sanctificati erant omnes.
2CHR|31|19|Porro pro filiis Aaron, sacerdotibus in agris et suburbanis urbium singularum dispositi erant nominatim viri, qui partes distribuerent universo sexui masculino de sacerdotibus et omni, qui recensitus erat inter Levitas.
2CHR|31|20|Fecit ergo Ezechias secundum haec in omni Iuda operatusque est bonum et rectum et verum coram Domino Deo suo.
2CHR|31|21|Et in universo opere, quod coepit in servitio domus Dei, et iuxta legem et praeceptum volens requirere Deum suum, in toto corde suo operatus et prosperatus est.
2CHR|32|1|Post quae et huiuscemodi fidem venit Sennacherib rex Assyriorum et ingressus Iudam obsedit civitates munitas volens eas capere.
2CHR|32|2|Quod cum vidisset Ezechias, venisse scilicet Sennacherib et totum belli impetum verti contra Ierusalem,
2CHR|32|3|inito cum principibus consilio virisque fortissimis, ut obturarent capita fontium, qui erant extra urbem, et, hoc omnium decernente sententia,
2CHR|32|4|congregata est plurima multitudo, et obturaverunt cunctos fontes et rivum, qui fluebat in medio terrae, dicentes: " Ne veniant reges Assyriorum et inveniant aquarum abundantiam! ".
2CHR|32|5|Aedificavit quoque agens industrie omnem murum, qui fuerat dissipatus, et exstruxit turres desuper et forinsecus alterum murum instauravitque Mello in civitate David et fecit iacula plurima et clipeos.
2CHR|32|6|Constituitque principes belli super populum et convocavit illos ad se in platea portae civitatis ac locutus est ad cor eorum dicens:
2CHR|32|7|" Viriliter agite et confortamini! Nolite timere nec paveatis regem Assyriorum et universam multitudinem, quae est cum eo. Multo enim plures nobiscum sunt quam cum illo:
2CHR|32|8|cum illo est brachium carneum, nobiscum autem Dominus Deus noster, qui auxiliator est noster pugnatque pro nobis ". Confortatusque est populus huiuscemodi verbis Ezechiae regis Iudae.
2CHR|32|9|Quae postquam gesta sunt, misit Sennacherib rex Assyriorum servos suos Ierusalem - ipse enim cum universo exercitu obsidebat Lachis - ad Ezechiam regem Iudae et ad omnem populum, qui erat in urbe, dicens:
2CHR|32|10|" Haec dicit Sennacherib rex Assyriorum: In quo habentes fiduciam sedetis obsessi in Ierusalem?
2CHR|32|11|Nonne Ezechias decipit vos, ut tradat morti in fame et siti affirmans quod Dominus Deus vester liberet vos de manu regis Assyriorum?
2CHR|32|12|Numquid non iste est Ezechias, qui destruxit excelsa illius et altaria et praecepit Iudae et Ierusalem dicens: "Coram altari uno adorabitis et in ipso comburetis sacrificia"?
2CHR|32|13|An ignoratis quae ego fecerim et patres mei cunctis terrarum populis? Numquid praevaluerunt dii gentium terrarum liberare regionem suam de manu mea?
2CHR|32|14|Quis est de universis diis gentium, quas deleverunt patres mei, qui potuerit eruere populum suum de manu mea, ut possit etiam Deus vester eruere vos de hac manu?
2CHR|32|15|Non vos ergo decipiat Ezechias nec vana persuasione deludat, neque credatis ei! Si enim nullus potuit deus cunctarum gentium atque regnorum liberare populum suum de manu mea et de manu patrum meorum, quanto minus Deus vester poterit eruere vos de manu mea! ".
2CHR|32|16|Sed et alia multa locuti sunt servi eius contra Dominum Deum et contra Ezechiam servum eius.
2CHR|32|17|Epistulas quoque scripsit plenas blasphemiae in Dominum, Deum Israel, et locutus est adversus eum: " Sicut dii gentium terrarum non potuerunt liberare populos suos de manu mea, sic et Deus Ezechiae eruere non poterit populum suum de manu ista ".
2CHR|32|18|Insuper et clamore magno, lingua Iudaica, ad populum Ierusalem, qui sedebat in muro, personabant, ut terrerent et perturbarent eos et caperent civitatem.
2CHR|32|19|Locutusque est Sennacherib contra Deum Ierusalem sicut adversum deos populorum terrae opera manuum hominum.
2CHR|32|20|Oraverunt igitur Ezechias rex et Isaias filius Amos prophetes adversum hanc blasphemiam ac vociferati sunt in caelum.
2CHR|32|21|Et misit Dominus angelum, qui percussit omnem virum robustum et bellatorem et principem in castris regis Assyriorum; reversusque est cum ignominia in terram suam. Cumque ingressus esset domum dei sui, filii, qui egressi fuerant de visceribus eius, interfecerunt eum ibi gladio.
2CHR|32|22|Salvavit ergo Dominus Ezechiam et habitatores Ierusalem de manu Sennacherib regis Assyriorum et de manu omnium et praestitit eis quietem per circuitum.
2CHR|32|23|Multi etiam deferebant munera Domino in Ierusalem et res pretiosas Ezechiae regi Iudae, qui exaltatus est post haec coram cunctis gentibus.
2CHR|32|24|In diebus illis aegrotavit Ezechias usque ad mortem et oravit Dominum; exaudivitque eum et dedit ei signum.
2CHR|32|25|Sed non iuxta beneficia, quae acceperat, retribuit, quia elevatum est cor eius; et facta est contra eum ira et contra Iudam et Ierusalem.
2CHR|32|26|Humiliatusque est postea, eo quod exaltatum fuisset cor eius, tam ipse quam habitatores Ierusalem; et idcirco non venit super eos ira Domini in diebus Ezechiae.
2CHR|32|27|Fuit autem Ezechias dives et inclitus valde; et thesauros sibi plurimos congregavit argenti, auri et lapidis pretiosi, aromatum et clipeorum omnisque generis rerum pretiosarum.
2CHR|32|28|Apothecas quoque frumenti, vini et olei et praesepia omnium iumentorum caulasque pecoribus
2CHR|32|29|et urbes exaedificavit sibi; habebat quippe greges ovium et armentorum innumerabiles, eo quod dedisset ei Deus substantiam multam nimis.
2CHR|32|30|Ipse est Ezechias, qui obturavit superiorem exitum aquarum Gihon et avertit eas subter ad occidentem urbis David. In omnibus operibus suis prosperatus est.
2CHR|32|31|Attamen sic in legatione principum Babylonis, qui missi fuerant ad eum, ut interrogarent de portento, quod acciderat super terram, dereliquit eum Deus, ut tentaretur, et nota fierent omnia, quae erant in corde eius.
2CHR|32|32|Reliqua autem gestorum Ezechiae et misericordiarum eius scripta sunt in visione Isaiae filii Amos prophetae et in libro regum Iudae et Israel.
2CHR|32|33|Dormivitque Ezechias cum patribus suis, et sepelierunt eum in ascensu ad sepulcra filiorum David; et celebravit eius exsequias universus Iuda et omnes habitatores Ierusalem. Regnavitque Manasses filius eius pro eo.
2CHR|33|1|Duodecim annorum erat Manasses, cum regnare coe pisset, et quinquaginta quinque annis regnavit in Ierusalem.
2CHR|33|2|Fecit autem malum coram Domino iuxta abominationes gentium, quas expulit Dominus coram filiis Israel.
2CHR|33|3|Et conversus instauravit excelsa, quae demolitus fuerat Ezechias pater eius, construxitque aras Baalim et fecit palos et adoravit omnem militiam caeli et coluit eam.
2CHR|33|4|Aedificavit quoque altaria in domo Domini, de qua dixerat Dominus: " In Ierusalem erit nomen meum in aeternum ".
2CHR|33|5|Aedificavit autem ea cuncto exercitui caeli in duobus atriis domus Domini.
2CHR|33|6|Transireque fecit filios suos per ignem in valle filii Ennom. Hariolatus est, sectabatur auguria, maleficis artibus inserviebat, habebat secum pythones et aruspices; multaque mala operatus est coram Domino, ut irritaret eum.
2CHR|33|7|Posuit quoque sculptile, idolum, quod fecerat, in domo Dei, de qua locutus est Deus ad David et ad Salomonem filium eius dicens: " In domo hac et in Ierusalem, quam elegi de cunctis tribubus Israel, ponam nomen meum in sempiternum.
2CHR|33|8|Et moveri non faciam pedem Israel de terra, quam tradidi patribus eorum, ita dumtaxat si custodierint facere, quae praecepi eis, cunctamque legem et praecepta atque iudicia, per manum Moysi ".
2CHR|33|9|Igitur Manasses seduxit Iudam et habitatores Ierusalem, ut facerent malum super omnes gentes, quas subverterat Dominus a facie filiorum Israel.
2CHR|33|10|Locutusque est Dominus ad eum et ad populum illius, et attendere noluerunt.
2CHR|33|11|Idcirco superinduxit eis principes exercitus regis Assyriorum; ceperuntque Manassen compedibus et vinctum catenis duxerunt Babylonem.
2CHR|33|12|Qui, postquam coangustatus est, oravit Dominum Deum suum et egit paenitentiam valde coram Deo patrum suorum.
2CHR|33|13|Deprecatusque est eum, et placatus ei exaudivit orationem eius reduxitque eum Ierusalem in regnum suum; et cognovit Manasses quod Dominus ipse esset Deus.
2CHR|33|14|Post haec aedificavit murum extra civitatem David ad occidentem Gihon in convalle et ad introitum portae Piscium per circuitum Ophel et exaltavit illum vehementer; constituitque principes exercitus in cunctis civitatibus Iudae munitis.
2CHR|33|15|Et abstulit deos alienos et idolum de domo Domini, aras quoque, quas fecerat in monte domus Domini et in Ierusalem, et proiecit omnia extra urbem.
2CHR|33|16|Porro instauravit altare Domini et immolavit super illud victimas pacificorum et pro gratiarum actione praecepitque Iudae, ut serviret Domino, Deo Israel.
2CHR|33|17|Attamen adhuc populus immolabat in excelsis Domino Deo suo.
2CHR|33|18|Reliqua autem gestorum Manasse et obsecratio eius ad Deum suum, verba quoque videntium, qui loquebantur ad eum in nomine Domini, Dei Israel, continentur in sermonibus regum Israel.
2CHR|33|19|Oratio quoque eius et exauditio et cuncta peccata atque contemptus, loca etiam, in quibus aedificavit excelsa et fecit palos et statuas, antequam ageret paenitentiam, scripta sunt in sermonibus Hozai.
2CHR|33|20|Dormivit ergo Manasses cum patribus suis, et sepelierunt eum in domo sua. Regnavitque pro eo filius eius Amon.
2CHR|33|21|Viginti duorum annorum erat Amon, cum regnare coepisset, et duobus annis regnavit in Ierusalem.
2CHR|33|22|Fecitque malum in conspectu Domini, sicut fecerat Manasses pater eius, et cunctis idolis, quae Manasses fuerat fabricatus, immolavit atque servivit.
2CHR|33|23|Et non humiliavit se ante faciem Domini, sicut humiliaverat se Manasses pater eius, et multo maiora deliquit.
2CHR|33|24|Cumque coniurassent adversus eum servi sui, interfecerunt eum in domo sua.
2CHR|33|25|Porro populus terrae, caesis omnibus, qui conspiraverant contra regem Amon, consti tuit regem Iosiam filium eius pro eo.
2CHR|34|1|Octo annorum erat Iosias, cum regnare coepisset, et tri ginta et uno annis regnavit in Ierusalem.
2CHR|34|2|Fecitque quod erat rectum in conspectu Domini, et ambulavit in viis David patris sui; non declinavit neque ad dextram neque ad sinistram.
2CHR|34|3|Octavo autem anno regni sui, cum adhuc esset puer, coepit quaerere Deum patris sui David; et duodecimo anno coepit mundare Iudam et Ierusalem ab excelsis et palis sculptilibusque et conflatilibus.
2CHR|34|4|Destruxeruntque coram eo aras Baalim; et thymiamateria, quae eis superposita fuerant, demolitus est; palos etiam et sculptilia et conflatilia succidit atque comminuit et super tumulos eorum, qui eis immolare consueverant, fragmenta dispersit.
2CHR|34|5|Ossa praeterea sacerdotum combussit in altaribus ipsorum; mundavitque Iudam et Ierusalem,
2CHR|34|6|sed et in urbibus Manasse et Ephraim et Simeon usque Nephthali, in plateis eorum undique
2CHR|34|7|dissipavit altaria et palos et sculptilia contrivit in frusta; cunctaque thymiamateria demolitus est de universa terra Israel et reversus est Ierusalem.
2CHR|34|8|Igitur anno octavo decimo regni sui, cum mundaret terram et domum, misit Saphan filium Eseliae et Maasiam principem civitatis et Ioah filium Ioachaz a commentariis, ut instaurarent domum Domini Dei sui.
2CHR|34|9|Qui venerunt ad Helciam sacerdotem magnum acceptamque ab eo pecuniam, quae illata fuerat in domum Domini, et quam congregaverant Levitae ianitores de Manasse et Ephraim et universis reliquiis Israel ab omni quoque Iuda et Beniamin et habitatoribus Ierusalem,
2CHR|34|10|tradiderunt in manibus opificum, qui praeerant in domo Domini, et illi dederunt eam operariis, qui operabantur in domo Domini, ut instaurarent templum et infirma quaeque sarcirent;
2CHR|34|11|dederunt scilicet eam lignariis et caementariis, ut emerent lapides dolatos et ligna ad commissuras aedificii et ad contignationem domorum, quas destruxerant reges Iudae.
2CHR|34|12|Qui fideliter cuncta faciebant. Erant autem praepositi operantium Iahath et Abdias Levitae de filiis Merari, Zacharias et Mosollam de filiis Caath, qui dirigebant opus. Omnes autem Levitae scientes organis canere
2CHR|34|13|erant super eos, qui onera portabant et dirigebant omnes, qui varia opera faciebant. De Levitis quoque erant scribae et praefecti et ianitores.
2CHR|34|14|Cumque efferrent pecuniam, quae illata fuerat in templum Domini, repperit Helcias sacerdos librum legis Domini per manum Moysi
2CHR|34|15|et ait ad Saphan scribam: " Librum legis inveni in domo Domini ". Et tradidit ei.
2CHR|34|16|At ille intulit volumen ad regem et insuper nuntiavit ei dicens: " Omnia, quae dedisti in manu servorum tuorum, ecce complentur.
2CHR|34|17|Argentum, quod repertum est in domo Domini, effuderunt, datum que est praefectis et operariis ".
2CHR|34|18|Et nuntiavit Saphan scriba regi dicens: " Librum tradidit mihi Helcias sacerdos ". Et legebat illum Saphan coram rege.
2CHR|34|19|Et factum est, cum audisset rex verba legis, scidit vestimenta sua
2CHR|34|20|et praecepit Helciae et Ahicam filio Saphan et Abdon filio Micha, Saphan quoque scribae et Asaiae servo regis dicens:
2CHR|34|21|" Ite et consulite Dominum pro me et pro reliquiis Israel et Iudae super sermonibus libri, qui repertus est. Magnus enim furor Domini effusus est super nos, eo quod non custodierint patres nostri verba Domini, ut facerent iuxta omnia, quae scripta sunt in isto volumine ".
2CHR|34|22|Abiit igitur Helcias et hi, qui simul a rege missi fuerant, ad Holdam propheten uxorem Sellum filii Thecuae filii Haraas custodis vestium, quae habitabat in Ierusalem in secunda, et locuti sunt ei iuxta verba haec.
2CHR|34|23|Et illa respondit eis: " Haec dicit Dominus, Deus Israel: Dicite viro, qui misit vos ad me:
2CHR|34|24|Haec dicit Dominus: Ecce ego inducam mala super locum istum et super habitatores eius, cuncta maledicta, quae scripta sunt in libro hoc, quem legerunt coram rege Iudae,
2CHR|34|25|quia dereliquerunt me et sacrificaverunt diis alienis, ut me ad iracundiam provocarent in cunctis operibus manuum suarum; idcirco effundetur furor meus super locum istum et non exstinguetur.
2CHR|34|26|Ad regem autem Iudae, qui misit vos pro Domino consulendo, sic loquimini: Haec dicit Dominus, Deus Israel: Quoniam audisti verba voluminis,
2CHR|34|27|atque emollitum est cor tuum, et humiliatus es in conspectu Dei super his, quae dicta sunt contra locum hunc et habitatores Ierusalem, humiliatusque coram me scidisti vestimenta tua et flevisti coram me, ego quoque audivi, dicit Dominus.
2CHR|34|28|Ecce colligam te ad patres tuos, et infereris in sepulcrum tuum in pace; nec videbunt oculi tui omne malum, quod ego inducturus sum super locum istum et super habitatores eius ".Rettuleruntque itaque regi cuncta, quae dixerat.
2CHR|34|29|At ille, convocatis universis maioribus natu Iudae et Ierusalem,
2CHR|34|30|ascendit domum Domini, unaque omnes viri Iudae et habitatores Ierusalem, sacerdotes et Levitae et cunctus populus a minimo usque ad maximum. Quibus audientibus, in domo Domini legit rex omnia verba voluminis foederis inventi in domo Domini.
2CHR|34|31|Et stans in gradu suo percussit foedus coram Domino, ut ambularet post eum et custodiret praecepta et testimonia et iustificationes eius in toto corde suo et in tota anima sua faceretque verba foederis scripta in hoc libro.
2CHR|34|32|Adiuravit quoque super hoc omnes, qui reperti fuerant in Ierusalem et Beniamin; et fecerunt habitatores Ierusalem iuxta pactum Domini, Dei patrum suorum.
2CHR|34|33|Abstulit ergo Iosias cunctas abominationes de universis regionibus filiorum Israel et fecit omnes, qui inventi erant in Israel, servire Domino Deo suo. Cunctis diebus eius non recesserunt a Domino, Deo patrum suorum.
2CHR|35|1|Fecit autem Iosias in Ierusalem Pascha Domino, quod immolatum est quarta decima die mensis primi.
2CHR|35|2|Et constituit sacerdotes in officiis suis confortavitque eos, ut ministrarent in domo Domini.
2CHR|35|3|Levitis quoque, qui erudiebant omnem Israel et consecrati erant Domino, locutus est: " Ponite arcam sanctam in templum, quod aedificavit Salomon filius David rex Israel; nequaquam eam ultra umeris portabitis. Nunc ministrate Domino Deo vestro et populo eius Israel.
2CHR|35|4|Et praeparate vos per familias vestras in divisionibus singulis, sicut scripsit David rex Israel, et descripsit Salomon filius eius;
2CHR|35|5|et ministrate in sanctuario partibus familiarum fratrum vestrorum, filiorum populi, singulis pars familiae Levitarum.
2CHR|35|6|Mactate ergo Pascha et sanctificamini et praeparate vos pro fratribus vestris, ut faciatis iuxta verbum, quod locu tus est Dominus in manu Moysi.
2CHR|35|7|Dedit praeterea Iosias omni populo, qui ibi inventus fuerat pro Pascha, agnos et haedos de gregibus triginta milia, boumque tria milia; haec de regis universa substantia.
2CHR|35|8|Duces quoque eius sponte obtulerunt, tam populo quam sacerdotibus et Levitis; porro Helcias et Zacharias et Iahiel principes domus Domini dederunt sacerdotibus ad faciendum Pascha pecora commixtim duo milia sescenta et boves trecentos.
2CHR|35|9|Chonenias autem, Semeias etiam et Nathanael fratres eius necnon Hasabias et Iehiel et Iozabad principes Levitarum dederunt ceteris Levitis ad celebrandum Pascha quinque milia pecorum et boves quingentos.
2CHR|35|10|Praeparatumque est ministerium, et steterunt sacerdotes in loco suo, Levitae quoque in turmis iuxta regis imperium.
2CHR|35|11|Et mactatum est Pascha; asperseruntque sacerdotes manu sua sanguinem, et Levitae detraxerunt pelles holocaustorum
2CHR|35|12|et separaverunt holocaustum, ut darent partibus familiarum populi, et offerretur Domino, sicut scriptum est in libro Moysi. De bobus quoque fecere similiter.
2CHR|35|13|Et assaverunt Pascha super ignem, iuxta quod lege praeceptum est; pacificas vero hostias coxerunt in lebetis et caccabis et ollis et festinato distribuerunt universae plebi.
2CHR|35|14|Sibi autem et sacerdotibus postea paraverunt; nam in oblatione holocaustorum et adipum usque ad noctem sacerdotes fuerant occupati, unde Levitae et sibi et sacerdotibus filiis Aaron paraverunt novissimis.
2CHR|35|15|Porro cantores filii Asaph stabant in loco suo, iuxta praeceptum David et Asaph et Heman et Idithun prophetarum regis; ianitores vero per portas singulas observabant, ita ut ne puncto quidem discederent a ministerio, quia fratres eorum Levitae paraverunt eis cibos.
2CHR|35|16|Omnis igitur cultus Domini rite praeparatus est in die illa, ut facerent Pascha et offerrent holocausta super altare Domini, iuxta praeceptum regis Iosiae.
2CHR|35|17|Feceruntque filii Israel, qui reperti fuerant ibi, Pascha in tempore illo et sollemnitatem Azymorum septem diebus.
2CHR|35|18|Non fuit simile huic in Israel a diebus Samuelis prophetae, sed nec quisquam de cunctis regibus Israel fecit Pascha sicut Iosias cum sacerdotibus et Levitis et omni Iuda et Israel, qui repertus fuerat, et habitantibus in Ierusalem.
2CHR|35|19|Octavo decimo anno regni Iosiae hoc Pascha celebratum est.
2CHR|35|20|Postquam instauraverat Iosias templum, ascendit Nechao rex Aegypti ad pugnandum in Charchamis iuxta Euphraten. Et processit in occursum eius Iosias.
2CHR|35|21|At ille, missis ad eum nuntiis, ait: " Quid mihi et tibi est, rex Iudae? Non adversum te hodie venio, sed contra aliam pugno domum, ad quam me Deus festinato ire praecepit. Desine adversum Deum facere, qui mecum est, ne interficiat te ".
2CHR|35|22|Noluit Iosias reverti, sed audacter praeparavit contra eum bellum nec acquievit sermonibus Nechao ex ore Dei; verum perrexit, ut dimicaret in campo Mageddo.
2CHR|35|23|Ibique vulneratus a sagittariis dixit pueris suis: " Educite me de proelio, quia oppido vulneratus sum ".
2CHR|35|24|Qui transtulerunt eum de curru in alterum currum eius et asportaverunt in Ierusalem. Mortuusque est et sepultus in sepulcris patrum suorum; et universus Iuda et Ierusalem luxerunt eum.
2CHR|35|25|Ieremias fecit planctum super Iosiam; et omnes cantores atque cantrices usque in praesentem diem lamentationes super Iosia replicant, et quasi lex obtinuit in Israel; ecce scriptum fertur in Lamentationibus.
2CHR|35|26|Reliqua autem gestorum Iosiae et misericordiae eius, quae lege praecepta sunt Domini,
2CHR|35|27|gesta quoque illius prima et novissima scripta sunt in libro regum Israel et Iudae.
2CHR|36|1|Tulit ergo populus terrae Ioachaz filium Iosiae et con stituit regem pro patre suo in Ierusalem.
2CHR|36|2|Viginti trium annorum erat Ioachaz, cum regnare coepisset, et tribus mensibus regnavit in Ierusalem.
2CHR|36|3|Amovit autem eum rex Aegypti, cum venisset Ierusalem, et condemnavit terram centum talentis argenti et talento auri.
2CHR|36|4|Constituitque regem pro eo Eliachim fratrem eius super Iudam et Ierusalem et vertit nomen eius Ioachim. Ipsum vero Ioachaz tulit secum et adduxit in Aegyptum.
2CHR|36|5|Viginti quinque annorum erat Ioachim, cum regnare coepisset, et undecim annis regnavit in Ierusalem; fecitque malum coram Domino Deo suo.
2CHR|36|6|Contra hunc ascendit Nabuchodonosor rex Chaldaeorum et vinctum catenis duxit in Babylonem,
2CHR|36|7|ad quam et ex vasis Domini transtulit et posuit ea in templo suo.
2CHR|36|8|Reliqua autem gestorum Ioachim et abominationum eius, quas operatus est, et quae inventa sunt contra eum, continentur in libro regum Israel et Iudae. Regnavitque autem Ioachin filius eius pro eo.
2CHR|36|9|Decem et octo annorum erat Ioachin, cum regnare coepisset, et tribus mensibus ac decem diebus regnavit in Ierusalem; fecitque malum in conspectu Domini.
2CHR|36|10|Cumque anni circulus volveretur, misit Nabuchodonosor rex, qui adduxerunt eum in Babylonem, asportatis simul pretiosissimis vasis domus Domini; regem vero constituit Sedeciam fratrem eius super Iudam et Ierusalem.
2CHR|36|11|Viginti et unius anni erat Sedecias, cum regnare coepisset, et undecim annis regnavit in Ierusalem.
2CHR|36|12|Fecitque malum in oculis Domini Dei sui nec humiliavit se coram Ieremia propheta loquente ad se ex ore Domini.
2CHR|36|13|Contra regem quoque Nabuchodonosor rebellavit, qui adiuraverat eum per Deum, et induravit cervicem suam et cor, ut non reverteretur ad Dominum, Deum Israel.
2CHR|36|14|Sed et universi principes sacerdotum et populus multiplicaverunt praevaricationes suas iuxta universas abominationes gentium et polluerunt domum Domini, quam sanctificaverat in Ierusalem.
2CHR|36|15|Mittebat autem Dominus, Deus patrum suorum, ad illos per manum nuntiorum suorum de nocte consurgens et cotidie commonens, eo quod parceret populo et habitaculo suo.
2CHR|36|16|At illi subsannabant nuntios Dei et parvipendebant sermones eius illudebantque prophetis, donec ascenderet furor Domini in populum eius, et esset nulla curatio.
2CHR|36|17|Adduxit enim super eos regem Chaldaeorum et interfecit iuvenes eorum gladio in domo sanctuarii sui; non est misertus adulescentis et virginis et senis nec decrepiti quidem, sed omnes tradidit in manibus eius.
2CHR|36|18|Universaque vasa domus Dei tam maiora quam minora et thesauros templi et regis et principum transtulit in Babylonem.
2CHR|36|19|Incenderunt hostes domum Dei destruxeruntque murum Ierusalem, universa palatia combusserunt et, quidquid pretiosum fuerat, demoliti sunt.
2CHR|36|20|Si quis evaserat gladium, ductus in Babylonem servivit regi et filiis eius, donec imperaret rex Persarum,
2CHR|36|21|ut compleretur sermo Domini ex ore Ieremiae: donec terra acciperet sabbata sua, cunctis diebus devastationis egit sabbatum, usque dum complerentur septuaginta anni.
2CHR|36|22|Anno autem primo Cyri regis Persarum ad explendum sermonem Domini, quem locutus fuerat per os Ieremiae, suscitavit Dominus spiritum Cyri regis Persarum, qui iussit praedicari in universo regno suo etiam per scripturam dicens:
2CHR|36|23|" Haec dicit Cyrus rex Persarum: Omnia regna terrae dedit mihi Dominus, Deus caeli, et ipse praecepit mihi, ut aedificarem ei domum in Ierusalem, quae est in Iudaea. Quis ex vobis est de omni populo eius? Sit Dominus Deus suus cum eo, et ascendat ".
