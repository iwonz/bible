2TIM|1|1|Paul, an apostle of Christ Jesus by the will of God, according to the promise of life that is in Christ Jesus,
2TIM|1|2|To Timothy, my dear son: Grace, mercy and peace from God the Father and Christ Jesus our Lord.
2TIM|1|3|I thank God, whom I serve, as my forefathers did, with a clear conscience, as night and day I constantly remember you in my prayers.
2TIM|1|4|Recalling your tears, I long to see you, so that I may be filled with joy.
2TIM|1|5|I have been reminded of your sincere faith, which first lived in your grandmother Lois and in your mother Eunice and, I am persuaded, now lives in you also.
2TIM|1|6|For this reason I remind you to fan into flame the gift of God, which is in you through the laying on of my hands.
2TIM|1|7|For God did not give us a spirit of timidity, but a spirit of power, of love and of self-discipline.
2TIM|1|8|So do not be ashamed to testify about our Lord, or ashamed of me his prisoner. But join with me in suffering for the gospel, by the power of God,
2TIM|1|9|who has saved us and called us to a holy life--not because of anything we have done but because of his own purpose and grace. This grace was given us in Christ Jesus before the beginning of time,
2TIM|1|10|but it has now been revealed through the appearing of our Savior, Christ Jesus, who has destroyed death and has brought life and immortality to light through the gospel.
2TIM|1|11|And of this gospel I was appointed a herald and an apostle and a teacher.
2TIM|1|12|That is why I am suffering as I am. Yet I am not ashamed, because I know whom I have believed, and am convinced that he is able to guard what I have entrusted to him for that day.
2TIM|1|13|What you heard from me, keep as the pattern of sound teaching, with faith and love in Christ Jesus.
2TIM|1|14|Guard the good deposit that was entrusted to you--guard it with the help of the Holy Spirit who lives in us.
2TIM|1|15|You know that everyone in the province of Asia has deserted me, including Phygelus and Hermogenes.
2TIM|1|16|May the Lord show mercy to the household of Onesiphorus, because he often refreshed me and was not ashamed of my chains.
2TIM|1|17|On the contrary, when he was in Rome, he searched hard for me until he found me.
2TIM|1|18|May the Lord grant that he will find mercy from the Lord on that day! You know very well in how many ways he helped me in Ephesus.
2TIM|2|1|You then, my son, be strong in the grace that is in Christ Jesus.
2TIM|2|2|And the things you have heard me say in the presence of many witnesses entrust to reliable men who will also be qualified to teach others.
2TIM|2|3|Endure hardship with us like a good soldier of Christ Jesus.
2TIM|2|4|No one serving as a soldier gets involved in civilian affairs--he wants to please his commanding officer.
2TIM|2|5|Similarly, if anyone competes as an athlete, he does not receive the victor's crown unless he competes according to the rules.
2TIM|2|6|The hardworking farmer should be the first to receive a share of the crops.
2TIM|2|7|Reflect on what I am saying, for the Lord will give you insight into all this.
2TIM|2|8|Remember Jesus Christ, raised from the dead, descended from David. This is my gospel,
2TIM|2|9|for which I am suffering even to the point of being chained like a criminal. But God's word is not chained.
2TIM|2|10|Therefore I endure everything for the sake of the elect, that they too may obtain the salvation that is in Christ Jesus, with eternal glory.
2TIM|2|11|Here is a trustworthy saying: If we died with him, we will also live with him;
2TIM|2|12|if we endure, we will also reign with him. If we disown him, he will also disown us;
2TIM|2|13|if we are faithless, he will remain faithful, for he cannot disown himself.
2TIM|2|14|Keep reminding them of these things. Warn them before God against quarreling about words; it is of no value, and only ruins those who listen.
2TIM|2|15|Do your best to present yourself to God as one approved, a workman who does not need to be ashamed and who correctly handles the word of truth.
2TIM|2|16|Avoid godless chatter, because those who indulge in it will become more and more ungodly.
2TIM|2|17|Their teaching will spread like gangrene. Among them are Hymenaeus and Philetus,
2TIM|2|18|who have wandered away from the truth. They say that the resurrection has already taken place, and they destroy the faith of some.
2TIM|2|19|Nevertheless, God's solid foundation stands firm, sealed with this inscription: "The Lord knows those who are his," and, "Everyone who confesses the name of the Lord must turn away from wickedness."
2TIM|2|20|In a large house there are articles not only of gold and silver, but also of wood and clay; some are for noble purposes and some for ignoble.
2TIM|2|21|If a man cleanses himself from the latter, he will be an instrument for noble purposes, made holy, useful to the Master and prepared to do any good work.
2TIM|2|22|Flee the evil desires of youth, and pursue righteousness, faith, love and peace, along with those who call on the Lord out of a pure heart.
2TIM|2|23|Don't have anything to do with foolish and stupid arguments, because you know they produce quarrels.
2TIM|2|24|And the Lord's servant must not quarrel; instead, he must be kind to everyone, able to teach, not resentful.
2TIM|2|25|Those who oppose him he must gently instruct, in the hope that God will grant them repentance leading them to a knowledge of the truth,
2TIM|2|26|and that they will come to their senses and escape from the trap of the devil, who has taken them captive to do his will.
2TIM|3|1|But mark this: There will be terrible times in the last days.
2TIM|3|2|People will be lovers of themselves, lovers of money, boastful, proud, abusive, disobedient to their parents, ungrateful, unholy,
2TIM|3|3|without love, unforgiving, slanderous, without self-control, brutal, not lovers of the good,
2TIM|3|4|treacherous, rash, conceited, lovers of pleasure rather than lovers of God--
2TIM|3|5|having a form of godliness but denying its power. Have nothing to do with them.
2TIM|3|6|They are the kind who worm their way into homes and gain control over weak-willed women, who are loaded down with sins and are swayed by all kinds of evil desires,
2TIM|3|7|always learning but never able to acknowledge the truth.
2TIM|3|8|Just as Jannes and Jambres opposed Moses, so also these men oppose the truth--men of depraved minds, who, as far as the faith is concerned, are rejected.
2TIM|3|9|But they will not get very far because, as in the case of those men, their folly will be clear to everyone.
2TIM|3|10|You, however, know all about my teaching, my way of life, my purpose, faith, patience, love, endurance,
2TIM|3|11|persecutions, sufferings--what kinds of things happened to me in Antioch, Iconium and Lystra, the persecutions I endured. Yet the Lord rescued me from all of them.
2TIM|3|12|In fact, everyone who wants to live a godly life in Christ Jesus will be persecuted,
2TIM|3|13|while evil men and impostors will go from bad to worse, deceiving and being deceived.
2TIM|3|14|But as for you, continue in what you have learned and have become convinced of, because you know those from whom you learned it,
2TIM|3|15|and how from infancy you have known the holy Scriptures, which are able to make you wise for salvation through faith in Christ Jesus.
2TIM|3|16|All Scripture is God-breathed and is useful for teaching, rebuking, correcting and training in righteousness,
2TIM|3|17|so that the man of God may be thoroughly equipped for every good work.
2TIM|4|1|In the presence of God and of Christ Jesus, who will judge the living and the dead, and in view of his appearing and his kingdom, I give you this charge:
2TIM|4|2|Preach the Word; be prepared in season and out of season; correct, rebuke and encourage--with great patience and careful instruction.
2TIM|4|3|For the time will come when men will not put up with sound doctrine. Instead, to suit their own desires, they will gather around them a great number of teachers to say what their itching ears want to hear.
2TIM|4|4|They will turn their ears away from the truth and turn aside to myths.
2TIM|4|5|But you, keep your head in all situations, endure hardship, do the work of an evangelist, discharge all the duties of your ministry.
2TIM|4|6|For I am already being poured out like a drink offering, and the time has come for my departure.
2TIM|4|7|I have fought the good fight, I have finished the race, I have kept the faith.
2TIM|4|8|Now there is in store for me the crown of righteousness, which the Lord, the righteous Judge, will award to me on that day--and not only to me, but also to all who have longed for his appearing.
2TIM|4|9|Do your best to come to me quickly,
2TIM|4|10|for Demas, because he loved this world, has deserted me and has gone to Thessalonica. Crescens has gone to Galatia, and Titus to Dalmatia.
2TIM|4|11|Only Luke is with me. Get Mark and bring him with you, because he is helpful to me in my ministry.
2TIM|4|12|I sent Tychicus to Ephesus.
2TIM|4|13|When you come, bring the cloak that I left with Carpus at Troas, and my scrolls, especially the parchments.
2TIM|4|14|Alexander the metalworker did me a great deal of harm. The Lord will repay him for what he has done.
2TIM|4|15|You too should be on your guard against him, because he strongly opposed our message.
2TIM|4|16|At my first defense, no one came to my support, but everyone deserted me. May it not be held against them.
2TIM|4|17|But the Lord stood at my side and gave me strength, so that through me the message might be fully proclaimed and all the Gentiles might hear it. And I was delivered from the lion's mouth.
2TIM|4|18|The Lord will rescue me from every evil attack and will bring me safely to his heavenly kingdom. To him be glory for ever and ever. Amen.
2TIM|4|19|Greet Priscilla and Aquila and the household of Onesiphorus.
2TIM|4|20|Erastus stayed in Corinth, and I left Trophimus sick in Miletus.
2TIM|4|21|Do your best to get here before winter. Eubulus greets you, and so do Pudens, Linus, Claudia and all the brothers.
2TIM|4|22|The Lord be with your spirit. Grace be with you.
