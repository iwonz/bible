EZRA|1|1|In the first year of Cyrus king of Persia, in order to fulfill the word of the LORD spoken by Jeremiah, the LORD moved the heart of Cyrus king of Persia to make a proclamation throughout his realm and to put it in writing:
EZRA|1|2|"This is what Cyrus king of Persia says: "'The LORD, the God of heaven, has given me all the kingdoms of the earth and he has appointed me to build a temple for him at Jerusalem in Judah.
EZRA|1|3|Anyone of his people among you-may his God be with him, and let him go up to Jerusalem in Judah and build the temple of the LORD, the God of Israel, the God who is in Jerusalem.
EZRA|1|4|And the people of any place where survivors may now be living are to provide him with silver and gold, with goods and livestock, and with freewill offerings for the temple of God in Jerusalem.'"
EZRA|1|5|Then the family heads of Judah and Benjamin, and the priests and Levites-everyone whose heart God had moved-prepared to go up and build the house of the LORD in Jerusalem.
EZRA|1|6|All their neighbors assisted them with articles of silver and gold, with goods and livestock, and with valuable gifts, in addition to all the freewill offerings.
EZRA|1|7|Moreover, King Cyrus brought out the articles belonging to the temple of the LORD, which Nebuchadnezzar had carried away from Jerusalem and had placed in the temple of his god.
EZRA|1|8|Cyrus king of Persia had them brought by Mithredath the treasurer, who counted them out to Sheshbazzar the prince of Judah.
EZRA|1|9|This was the inventory: gold dishes 30 silver dishes 1,000 silver pans 29
EZRA|1|10|gold bowls 30 matching silver bowls 410 other articles 1,000
EZRA|1|11|In all, there were 5,400 articles of gold and of silver. Sheshbazzar brought all these along when the exiles came up from Babylon to Jerusalem.
EZRA|2|1|Now these are the people of the province who came up from the captivity of the exiles, whom Nebuchadnezzar king of Babylon had taken captive to Babylon (they returned to Jerusalem and Judah, each to his own town,
EZRA|2|2|in company with Zerubbabel, Jeshua, Nehemiah, Seraiah, Reelaiah, Mordecai, Bilshan, Mispar, Bigvai, Rehum and Baanah): The list of the men of the people of Israel:
EZRA|2|3|the descendants of Parosh 2,172
EZRA|2|4|of Shephatiah 372
EZRA|2|5|of Arah 775
EZRA|2|6|of Pahath-Moab (through the line of Jeshua and Joab) 2,812
EZRA|2|7|of Elam 1,254
EZRA|2|8|of Zattu 945
EZRA|2|9|of Zaccai 760
EZRA|2|10|of Bani 642
EZRA|2|11|of Bebai 623
EZRA|2|12|of Azgad 1,222
EZRA|2|13|of Adonikam 666
EZRA|2|14|of Bigvai 2,056
EZRA|2|15|of Adin 454
EZRA|2|16|of Ater (through Hezekiah) 98
EZRA|2|17|of Bezai 323
EZRA|2|18|of Jorah 112
EZRA|2|19|of Hashum 223
EZRA|2|20|of Gibbar 95
EZRA|2|21|the men of Bethlehem 123
EZRA|2|22|of Netophah 56
EZRA|2|23|of Anathoth 128
EZRA|2|24|of Azmaveth 42
EZRA|2|25|of Kiriath Jearim, Kephirah and Beeroth 743
EZRA|2|26|of Ramah and Geba 621
EZRA|2|27|of Micmash 122
EZRA|2|28|of Bethel and Ai 223
EZRA|2|29|of Nebo 52
EZRA|2|30|of Magbish 156
EZRA|2|31|of the other Elam 1,254
EZRA|2|32|of Harim 320
EZRA|2|33|of Lod, Hadid and Ono 725
EZRA|2|34|of Jericho 345
EZRA|2|35|of Senaah 3,630
EZRA|2|36|The priests: the descendants of Jedaiah (through the family of Jeshua) 973
EZRA|2|37|of Immer 1,052
EZRA|2|38|of Pashhur 1,247
EZRA|2|39|of Harim 1,017
EZRA|2|40|The Levites: the descendants of Jeshua and Kadmiel (through the line of Hodaviah) 74
EZRA|2|41|The singers: the descendants of Asaph 128
EZRA|2|42|The gatekeepers of the temple: the descendants of Shallum, Ater, Talmon, Akkub, Hatita and Shobai 139
EZRA|2|43|The temple servants: the descendants of Ziha, Hasupha, Tabbaoth,
EZRA|2|44|Keros, Siaha, Padon,
EZRA|2|45|Lebanah, Hagabah, Akkub,
EZRA|2|46|Hagab, Shalmai, Hanan,
EZRA|2|47|Giddel, Gahar, Reaiah,
EZRA|2|48|Rezin, Nekoda, Gazzam,
EZRA|2|49|Uzza, Paseah, Besai,
EZRA|2|50|Asnah, Meunim, Nephussim,
EZRA|2|51|Bakbuk, Hakupha, Harhur,
EZRA|2|52|Bazluth, Mehida, Harsha,
EZRA|2|53|Barkos, Sisera, Temah,
EZRA|2|54|Neziah and Hatipha
EZRA|2|55|The descendants of the servants of Solomon: the descendants of Sotai, Hassophereth, Peruda,
EZRA|2|56|Jaala, Darkon, Giddel,
EZRA|2|57|Shephatiah, Hattil, Pokereth-Hazzebaim and Ami
EZRA|2|58|The temple servants and the descendants of the servants of Solomon 392
EZRA|2|59|The following came up from the towns of Tel Melah, Tel Harsha, Kerub, Addon and Immer, but they could not show that their families were descended from Israel:
EZRA|2|60|The descendants of Delaiah, Tobiah and Nekoda 652
EZRA|2|61|And from among the priests: The descendants of Hobaiah, Hakkoz and Barzillai (a man who had married a daughter of Barzillai the Gileadite and was called by that name).
EZRA|2|62|These searched for their family records, but they could not find them and so were excluded from the priesthood as unclean.
EZRA|2|63|The governor ordered them not to eat any of the most sacred food until there was a priest ministering with the Urim and Thummim.
EZRA|2|64|The whole company numbered 42,360,
EZRA|2|65|besides their 7,337 menservants and maidservants; and they also had 200 men and women singers.
EZRA|2|66|They had 736 horses, 245 mules,
EZRA|2|67|435 camels and 6,720 donkeys.
EZRA|2|68|When they arrived at the house of the LORD in Jerusalem, some of the heads of the families gave freewill offerings toward the rebuilding of the house of God on its site.
EZRA|2|69|According to their ability they gave to the treasury for this work 61,000 drachmas of gold, 5,000 minas of silver and 100 priestly garments.
EZRA|2|70|The priests, the Levites, the singers, the gatekeepers and the temple servants settled in their own towns, along with some of the other people, and the rest of the Israelites settled in their towns.
EZRA|3|1|When the seventh month came and the Israelites had settled in their towns, the people assembled as one man in Jerusalem.
EZRA|3|2|Then Jeshua son of Jozadak and his fellow priests and Zerubbabel son of Shealtiel and his associates began to build the altar of the God of Israel to sacrifice burnt offerings on it, in accordance with what is written in the Law of Moses the man of God.
EZRA|3|3|Despite their fear of the peoples around them, they built the altar on its foundation and sacrificed burnt offerings on it to the LORD, both the morning and evening sacrifices.
EZRA|3|4|Then in accordance with what is written, they celebrated the Feast of Tabernacles with the required number of burnt offerings prescribed for each day.
EZRA|3|5|After that, they presented the regular burnt offerings, the New Moon sacrifices and the sacrifices for all the appointed sacred feasts of the LORD, as well as those brought as freewill offerings to the LORD.
EZRA|3|6|On the first day of the seventh month they began to offer burnt offerings to the LORD, though the foundation of the LORD's temple had not yet been laid.
EZRA|3|7|Then they gave money to the masons and carpenters, and gave food and drink and oil to the people of Sidon and Tyre, so that they would bring cedar logs by sea from Lebanon to Joppa, as authorized by Cyrus king of Persia.
EZRA|3|8|In the second month of the second year after their arrival at the house of God in Jerusalem, Zerubbabel son of Shealtiel, Jeshua son of Jozadak and the rest of their brothers (the priests and the Levites and all who had returned from the captivity to Jerusalem) began the work, appointing Levites twenty years of age and older to supervise the building of the house of the LORD.
EZRA|3|9|Jeshua and his sons and brothers and Kadmiel and his sons (descendants of Hodaviah ) and the sons of Henadad and their sons and brothers-all Levites-joined together in supervising those working on the house of God.
EZRA|3|10|When the builders laid the foundation of the temple of the LORD, the priests in their vestments and with trumpets, and the Levites (the sons of Asaph) with cymbals, took their places to praise the LORD, as prescribed by David king of Israel.
EZRA|3|11|With praise and thanksgiving they sang to the LORD: "He is good; his love to Israel endures forever." And all the people gave a great shout of praise to the LORD, because the foundation of the house of the LORD was laid.
EZRA|3|12|But many of the older priests and Levites and family heads, who had seen the former temple, wept aloud when they saw the foundation of this temple being laid, while many others shouted for joy.
EZRA|3|13|No one could distinguish the sound of the shouts of joy from the sound of weeping, because the people made so much noise. And the sound was heard far away.
EZRA|4|1|When the enemies of Judah and Benjamin heard that the exiles were building a temple for the LORD, the God of Israel,
EZRA|4|2|they came to Zerubbabel and to the heads of the families and said, "Let us help you build because, like you, we seek your God and have been sacrificing to him since the time of Esarhaddon king of Assyria, who brought us here."
EZRA|4|3|But Zerubbabel, Jeshua and the rest of the heads of the families of Israel answered, "You have no part with us in building a temple to our God. We alone will build it for the LORD, the God of Israel, as King Cyrus, the king of Persia, commanded us."
EZRA|4|4|Then the peoples around them set out to discourage the people of Judah and make them afraid to go on building.
EZRA|4|5|They hired counselors to work against them and frustrate their plans during the entire reign of Cyrus king of Persia and down to the reign of Darius king of Persia.
EZRA|4|6|At the beginning of the reign of Xerxes, they lodged an accusation against the people of Judah and Jerusalem.
EZRA|4|7|And in the days of Artaxerxes king of Persia, Bishlam, Mithredath, Tabeel and the rest of his associates wrote a letter to Artaxerxes. The letter was written in Aramaic script and in the Aramaic language.,
EZRA|4|8|Rehum the commanding officer and Shimshai the secretary wrote a letter against Jerusalem to Artaxerxes the king as follows:
EZRA|4|9|Rehum the commanding officer and Shimshai the secretary, together with the rest of their associates-the judges and officials over the men from Tripolis, Persia, Erech and Babylon, the Elamites of Susa,
EZRA|4|10|and the other people whom the great and honorable Ashurbanipal deported and settled in the city of Samaria and elsewhere in Trans-Euphrates.
EZRA|4|11|(This is a copy of the letter they sent him.) To King Artaxerxes, From your servants, the men of Trans-Euphrates:
EZRA|4|12|The king should know that the Jews who came up to us from you have gone to Jerusalem and are rebuilding that rebellious and wicked city. They are restoring the walls and repairing the foundations.
EZRA|4|13|Furthermore, the king should know that if this city is built and its walls are restored, no more taxes, tribute or duty will be paid, and the royal revenues will suffer.
EZRA|4|14|Now since we are under obligation to the palace and it is not proper for us to see the king dishonored, we are sending this message to inform the king,
EZRA|4|15|so that a search may be made in the archives of your predecessors. In these records you will find that this city is a rebellious city, troublesome to kings and provinces, a place of rebellion from ancient times. That is why this city was destroyed.
EZRA|4|16|We inform the king that if this city is built and its walls are restored, you will be left with nothing in Trans-Euphrates.
EZRA|4|17|The king sent this reply: To Rehum the commanding officer, Shimshai the secretary and the rest of their associates living in Samaria and elsewhere in Trans-Euphrates: Greetings.
EZRA|4|18|The letter you sent us has been read and translated in my presence.
EZRA|4|19|I issued an order and a search was made, and it was found that this city has a long history of revolt against kings and has been a place of rebellion and sedition.
EZRA|4|20|Jerusalem has had powerful kings ruling over the whole of Trans-Euphrates, and taxes, tribute and duty were paid to them.
EZRA|4|21|Now issue an order to these men to stop work, so that this city will not be rebuilt until I so order.
EZRA|4|22|Be careful not to neglect this matter. Why let this threat grow, to the detriment of the royal interests?
EZRA|4|23|As soon as the copy of the letter of King Artaxerxes was read to Rehum and Shimshai the secretary and their associates, they went immediately to the Jews in Jerusalem and compelled them by force to stop.
EZRA|4|24|Thus the work on the house of God in Jerusalem came to a standstill until the second year of the reign of Darius king of Persia.
EZRA|5|1|Now Haggai the prophet and Zechariah the prophet, a descendant of Iddo, prophesied to the Jews in Judah and Jerusalem in the name of the God of Israel, who was over them.
EZRA|5|2|Then Zerubbabel son of Shealtiel and Jeshua son of Jozadak set to work to rebuild the house of God in Jerusalem. And the prophets of God were with them, helping them.
EZRA|5|3|At that time Tattenai, governor of Trans-Euphrates, and Shethar-Bozenai and their associates went to them and asked, "Who authorized you to rebuild this temple and restore this structure?"
EZRA|5|4|They also asked, "What are the names of the men constructing this building?"
EZRA|5|5|But the eye of their God was watching over the elders of the Jews, and they were not stopped until a report could go to Darius and his written reply be received.
EZRA|5|6|This is a copy of the letter that Tattenai, governor of Trans-Euphrates, and Shethar-Bozenai and their associates, the officials of Trans-Euphrates, sent to King Darius.
EZRA|5|7|The report they sent him read as follows: To King Darius: Cordial greetings.
EZRA|5|8|The king should know that we went to the district of Judah, to the temple of the great God. The people are building it with large stones and placing the timbers in the walls. The work is being carried on with diligence and is making rapid progress under their direction.
EZRA|5|9|We questioned the elders and asked them, "Who authorized you to rebuild this temple and restore this structure?"
EZRA|5|10|We also asked them their names, so that we could write down the names of their leaders for your information.
EZRA|5|11|This is the answer they gave us: "We are the servants of the God of heaven and earth, and we are rebuilding the temple that was built many years ago, one that a great king of Israel built and finished.
EZRA|5|12|But because our fathers angered the God of heaven, he handed them over to Nebuchadnezzar the Chaldean, king of Babylon, who destroyed this temple and deported the people to Babylon.
EZRA|5|13|"However, in the first year of Cyrus king of Babylon, King Cyrus issued a decree to rebuild this house of God.
EZRA|5|14|He even removed from the temple of Babylon the gold and silver articles of the house of God, which Nebuchadnezzar had taken from the temple in Jerusalem and brought to the temple in Babylon. "Then King Cyrus gave them to a man named Sheshbazzar, whom he had appointed governor,
EZRA|5|15|and he told him, 'Take these articles and go and deposit them in the temple in Jerusalem. And rebuild the house of God on its site.'
EZRA|5|16|So this Sheshbazzar came and laid the foundations of the house of God in Jerusalem. From that day to the present it has been under construction but is not yet finished."
EZRA|5|17|Now if it pleases the king, let a search be made in the royal archives of Babylon to see if King Cyrus did in fact issue a decree to rebuild this house of God in Jerusalem. Then let the king send us his decision in this matter.
EZRA|6|1|King Darius then issued an order, and they searched in the archives stored in the treasury at Babylon.
EZRA|6|2|A scroll was found in the citadel of Ecbatana in the province of Media, and this was written on it: Memorandum:
EZRA|6|3|In the first year of King Cyrus, the king issued a decree concerning the temple of God in Jerusalem: Let the temple be rebuilt as a place to present sacrifices, and let its foundations be laid. It is to be ninety feet high and ninety feet wide,
EZRA|6|4|with three courses of large stones and one of timbers. The costs are to be paid by the royal treasury.
EZRA|6|5|Also, the gold and silver articles of the house of God, which Nebuchadnezzar took from the temple in Jerusalem and brought to Babylon, are to be returned to their places in the temple in Jerusalem; they are to be deposited in the house of God.
EZRA|6|6|Now then, Tattenai, governor of Trans-Euphrates, and Shethar-Bozenai and you, their fellow officials of that province, stay away from there.
EZRA|6|7|Do not interfere with the work on this temple of God. Let the governor of the Jews and the Jewish elders rebuild this house of God on its site.
EZRA|6|8|Moreover, I hereby decree what you are to do for these elders of the Jews in the construction of this house of God: The expenses of these men are to be fully paid out of the royal treasury, from the revenues of Trans-Euphrates, so that the work will not stop.
EZRA|6|9|Whatever is needed-young bulls, rams, male lambs for burnt offerings to the God of heaven, and wheat, salt, wine and oil, as requested by the priests in Jerusalem-must be given them daily without fail,
EZRA|6|10|so that they may offer sacrifices pleasing to the God of heaven and pray for the well-being of the king and his sons.
EZRA|6|11|Furthermore, I decree that if anyone changes this edict, a beam is to be pulled from his house and he is to be lifted up and impaled on it. And for this crime his house is to be made a pile of rubble.
EZRA|6|12|May God, who has caused his Name to dwell there, overthrow any king or people who lifts a hand to change this decree or to destroy this temple in Jerusalem. I Darius have decreed it. Let it be carried out with diligence.
EZRA|6|13|Then, because of the decree King Darius had sent, Tattenai, governor of Trans-Euphrates, and Shethar-Bozenai and their associates carried it out with diligence.
EZRA|6|14|So the elders of the Jews continued to build and prosper under the preaching of Haggai the prophet and Zechariah, a descendant of Iddo. They finished building the temple according to the command of the God of Israel and the decrees of Cyrus, Darius and Artaxerxes, kings of Persia.
EZRA|6|15|The temple was completed on the third day of the month Adar, in the sixth year of the reign of King Darius.
EZRA|6|16|Then the people of Israel-the priests, the Levites and the rest of the exiles-celebrated the dedication of the house of God with joy.
EZRA|6|17|For the dedication of this house of God they offered a hundred bulls, two hundred rams, four hundred male lambs and, as a sin offering for all Israel, twelve male goats, one for each of the tribes of Israel.
EZRA|6|18|And they installed the priests in their divisions and the Levites in their groups for the service of God at Jerusalem, according to what is written in the Book of Moses.
EZRA|6|19|On the fourteenth day of the first month, the exiles celebrated the Passover.
EZRA|6|20|The priests and Levites had purified themselves and were all ceremonially clean. The Levites slaughtered the Passover lamb for all the exiles, for their brothers the priests and for themselves.
EZRA|6|21|So the Israelites who had returned from the exile ate it, together with all who had separated themselves from the unclean practices of their Gentile neighbors in order to seek the LORD, the God of Israel.
EZRA|6|22|For seven days they celebrated with joy the Feast of Unleavened Bread, because the LORD had filled them with joy by changing the attitude of the king of Assyria, so that he assisted them in the work on the house of God, the God of Israel.
EZRA|7|1|After these things, during the reign of Artaxerxes king of Persia, Ezra son of Seraiah, the son of Azariah, the son of Hilkiah,
EZRA|7|2|the son of Shallum, the son of Zadok, the son of Ahitub,
EZRA|7|3|the son of Amariah, the son of Azariah, the son of Meraioth,
EZRA|7|4|the son of Zerahiah, the son of Uzzi, the son of Bukki,
EZRA|7|5|the son of Abishua, the son of Phinehas, the son of Eleazar, the son of Aaron the chief priest-
EZRA|7|6|this Ezra came up from Babylon. He was a teacher well versed in the Law of Moses, which the LORD, the God of Israel, had given. The king had granted him everything he asked, for the hand of the LORD his God was on him.
EZRA|7|7|Some of the Israelites, including priests, Levites, singers, gatekeepers and temple servants, also came up to Jerusalem in the seventh year of King Artaxerxes.
EZRA|7|8|Ezra arrived in Jerusalem in the fifth month of the seventh year of the king.
EZRA|7|9|He had begun his journey from Babylon on the first day of the first month, and he arrived in Jerusalem on the first day of the fifth month, for the gracious hand of his God was on him.
EZRA|7|10|For Ezra had devoted himself to the study and observance of the Law of the LORD, and to teaching its decrees and laws in Israel.
EZRA|7|11|This is a copy of the letter King Artaxerxes had given to Ezra the priest and teacher, a man learned in matters concerning the commands and decrees of the LORD for Israel:
EZRA|7|12|Artaxerxes, king of kings, To Ezra the priest, a teacher of the Law of the God of heaven: Greetings.
EZRA|7|13|Now I decree that any of the Israelites in my kingdom, including priests and Levites, who wish to go to Jerusalem with you, may go.
EZRA|7|14|You are sent by the king and his seven advisers to inquire about Judah and Jerusalem with regard to the Law of your God, which is in your hand.
EZRA|7|15|Moreover, you are to take with you the silver and gold that the king and his advisers have freely given to the God of Israel, whose dwelling is in Jerusalem,
EZRA|7|16|together with all the silver and gold you may obtain from the province of Babylon, as well as the freewill offerings of the people and priests for the temple of their God in Jerusalem.
EZRA|7|17|With this money be sure to buy bulls, rams and male lambs, together with their grain offerings and drink offerings, and sacrifice them on the altar of the temple of your God in Jerusalem.
EZRA|7|18|You and your brother Jews may then do whatever seems best with the rest of the silver and gold, in accordance with the will of your God.
EZRA|7|19|Deliver to the God of Jerusalem all the articles entrusted to you for worship in the temple of your God.
EZRA|7|20|And anything else needed for the temple of your God that you may have occasion to supply, you may provide from the royal treasury.
EZRA|7|21|Now I, King Artaxerxes, order all the treasurers of Trans-Euphrates to provide with diligence whatever Ezra the priest, a teacher of the Law of the God of heaven, may ask of you-
EZRA|7|22|up to a hundred talents of silver, a hundred cors of wheat, a hundred baths of wine, a hundred baths of olive oil, and salt without limit.
EZRA|7|23|Whatever the God of heaven has prescribed, let it be done with diligence for the temple of the God of heaven. Why should there be wrath against the realm of the king and of his sons?
EZRA|7|24|You are also to know that you have no authority to impose taxes, tribute or duty on any of the priests, Levites, singers, gatekeepers, temple servants or other workers at this house of God.
EZRA|7|25|And you, Ezra, in accordance with the wisdom of your God, which you possess, appoint magistrates and judges to administer justice to all the people of Trans-Euphrates-all who know the laws of your God. And you are to teach any who do not know them.
EZRA|7|26|Whoever does not obey the law of your God and the law of the king must surely be punished by death, banishment, confiscation of property, or imprisonment.
EZRA|7|27|Praise be to the LORD, the God of our fathers, who has put it into the king's heart to bring honor to the house of the LORD in Jerusalem in this way
EZRA|7|28|and who has extended his good favor to me before the king and his advisers and all the king's powerful officials. Because the hand of the LORD my God was on me, I took courage and gathered leading men from Israel to go up with me.
EZRA|8|1|These are the family heads and those registered with them who came up with me from Babylon during the reign of King Artaxerxes:
EZRA|8|2|of the descendants of Phinehas, Gershom; of the descendants of Ithamar, Daniel; of the descendants of David, Hattush
EZRA|8|3|of the descendants of Shecaniah; of the descendants of Parosh, Zechariah, and with him were registered 150 men;
EZRA|8|4|of the descendants of Pahath-Moab, Eliehoenai son of Zerahiah, and with him 200 men;
EZRA|8|5|of the descendants of Zattu, Shecaniah son of Jahaziel, and with him 300 men;
EZRA|8|6|of the descendants of Adin, Ebed son of Jonathan, and with him 50 men;
EZRA|8|7|of the descendants of Elam, Jeshaiah son of Athaliah, and with him 70 men;
EZRA|8|8|of the descendants of Shephatiah, Zebadiah son of Michael, and with him 80 men;
EZRA|8|9|of the descendants of Joab, Obadiah son of Jehiel, and with him 218 men;
EZRA|8|10|of the descendants of Bani, Shelomith son of Josiphiah, and with him 160 men;
EZRA|8|11|of the descendants of Bebai, Zechariah son of Bebai, and with him 28 men;
EZRA|8|12|of the descendants of Azgad, Johanan son of Hakkatan, and with him 110 men;
EZRA|8|13|of the descendants of Adonikam, the last ones, whose names were Eliphelet, Jeuel and Shemaiah, and with them 60 men;
EZRA|8|14|of the descendants of Bigvai, Uthai and Zaccur, and with them 70 men.
EZRA|8|15|I assembled them at the canal that flows toward Ahava, and we camped there three days. When I checked among the people and the priests, I found no Levites there.
EZRA|8|16|So I summoned Eliezer, Ariel, Shemaiah, Elnathan, Jarib, Elnathan, Nathan, Zechariah and Meshullam, who were leaders, and Joiarib and Elnathan, who were men of learning,
EZRA|8|17|and I sent them to Iddo, the leader in Casiphia. I told them what to say to Iddo and his kinsmen, the temple servants in Casiphia, so that they might bring attendants to us for the house of our God.
EZRA|8|18|Because the gracious hand of our God was on us, they brought us Sherebiah, a capable man, from the descendants of Mahli son of Levi, the son of Israel, and Sherebiah's sons and brothers, 18 men;
EZRA|8|19|and Hashabiah, together with Jeshaiah from the descendants of Merari, and his brothers and nephews, 20 men.
EZRA|8|20|They also brought 220 of the temple servants-a body that David and the officials had established to assist the Levites. All were registered by name.
EZRA|8|21|There, by the Ahava Canal, I proclaimed a fast, so that we might humble ourselves before our God and ask him for a safe journey for us and our children, with all our possessions.
EZRA|8|22|I was ashamed to ask the king for soldiers and horsemen to protect us from enemies on the road, because we had told the king, "The gracious hand of our God is on everyone who looks to him, but his great anger is against all who forsake him."
EZRA|8|23|So we fasted and petitioned our God about this, and he answered our prayer.
EZRA|8|24|Then I set apart twelve of the leading priests, together with Sherebiah, Hashabiah and ten of their brothers,
EZRA|8|25|and I weighed out to them the offering of silver and gold and the articles that the king, his advisers, his officials and all Israel present there had donated for the house of our God.
EZRA|8|26|I weighed out to them 650 talents of silver, silver articles weighing 100 talents, 100 talents of gold,
EZRA|8|27|20 bowls of gold valued at 1,000 darics, and two fine articles of polished bronze, as precious as gold.
EZRA|8|28|I said to them, "You as well as these articles are consecrated to the LORD. The silver and gold are a freewill offering to the LORD, the God of your fathers.
EZRA|8|29|Guard them carefully until you weigh them out in the chambers of the house of the LORD in Jerusalem before the leading priests and the Levites and the family heads of Israel."
EZRA|8|30|Then the priests and Levites received the silver and gold and sacred articles that had been weighed out to be taken to the house of our God in Jerusalem.
EZRA|8|31|On the twelfth day of the first month we set out from the Ahava Canal to go to Jerusalem. The hand of our God was on us, and he protected us from enemies and bandits along the way.
EZRA|8|32|So we arrived in Jerusalem, where we rested three days.
EZRA|8|33|On the fourth day, in the house of our God, we weighed out the silver and gold and the sacred articles into the hands of Meremoth son of Uriah, the priest. Eleazar son of Phinehas was with him, and so were the Levites Jozabad son of Jeshua and Noadiah son of Binnui.
EZRA|8|34|Everything was accounted for by number and weight, and the entire weight was recorded at that time.
EZRA|8|35|Then the exiles who had returned from captivity sacrificed burnt offerings to the God of Israel: twelve bulls for all Israel, ninety-six rams, seventy-seven male lambs and, as a sin offering, twelve male goats. All this was a burnt offering to the LORD.
EZRA|8|36|They also delivered the king's orders to the royal satraps and to the governors of Trans-Euphrates, who then gave assistance to the people and to the house of God.
EZRA|9|1|After these things had been done, the leaders came to me and said, "The people of Israel, including the priests and the Levites, have not kept themselves separate from the neighboring peoples with their detestable practices, like those of the Canaanites, Hittites, Perizzites, Jebusites, Ammonites, Moabites, Egyptians and Amorites.
EZRA|9|2|They have taken some of their daughters as wives for themselves and their sons, and have mingled the holy race with the peoples around them. And the leaders and officials have led the way in this unfaithfulness."
EZRA|9|3|When I heard this, I tore my tunic and cloak, pulled hair from my head and beard and sat down appalled.
EZRA|9|4|Then everyone who trembled at the words of the God of Israel gathered around me because of this unfaithfulness of the exiles. And I sat there appalled until the evening sacrifice.
EZRA|9|5|Then, at the evening sacrifice, I rose from my self-abasement, with my tunic and cloak torn, and fell on my knees with my hands spread out to the LORD my God
EZRA|9|6|and prayed: "O my God, I am too ashamed and disgraced to lift up my face to you, my God, because our sins are higher than our heads and our guilt has reached to the heavens.
EZRA|9|7|From the days of our forefathers until now, our guilt has been great. Because of our sins, we and our kings and our priests have been subjected to the sword and captivity, to pillage and humiliation at the hand of foreign kings, as it is today.
EZRA|9|8|"But now, for a brief moment, the LORD our God has been gracious in leaving us a remnant and giving us a firm place in his sanctuary, and so our God gives light to our eyes and a little relief in our bondage.
EZRA|9|9|Though we are slaves, our God has not deserted us in our bondage. He has shown us kindness in the sight of the kings of Persia: He has granted us new life to rebuild the house of our God and repair its ruins, and he has given us a wall of protection in Judah and Jerusalem.
EZRA|9|10|"But now, O our God, what can we say after this? For we have disregarded the commands
EZRA|9|11|you gave through your servants the prophets when you said: 'The land you are entering to possess is a land polluted by the corruption of its peoples. By their detestable practices they have filled it with their impurity from one end to the other.
EZRA|9|12|Therefore, do not give your daughters in marriage to their sons or take their daughters for your sons. Do not seek a treaty of friendship with them at any time, that you may be strong and eat the good things of the land and leave it to your children as an everlasting inheritance.'
EZRA|9|13|"What has happened to us is a result of our evil deeds and our great guilt, and yet, our God, you have punished us less than our sins have deserved and have given us a remnant like this.
EZRA|9|14|Shall we again break your commands and intermarry with the peoples who commit such detestable practices? Would you not be angry enough with us to destroy us, leaving us no remnant or survivor?
EZRA|9|15|O LORD, God of Israel, you are righteous! We are left this day as a remnant. Here we are before you in our guilt, though because of it not one of us can stand in your presence."
EZRA|10|1|While Ezra was praying and confessing, weeping and throwing himself down before the house of God, a large crowd of Israelites-men, women and children-gathered around him. They too wept bitterly.
EZRA|10|2|Then Shecaniah son of Jehiel, one of the descendants of Elam, said to Ezra, "We have been unfaithful to our God by marrying foreign women from the peoples around us. But in spite of this, there is still hope for Israel.
EZRA|10|3|Now let us make a covenant before our God to send away all these women and their children, in accordance with the counsel of my lord and of those who fear the commands of our God. Let it be done according to the Law.
EZRA|10|4|Rise up; this matter is in your hands. We will support you, so take courage and do it."
EZRA|10|5|So Ezra rose up and put the leading priests and Levites and all Israel under oath to do what had been suggested. And they took the oath.
EZRA|10|6|Then Ezra withdrew from before the house of God and went to the room of Jehohanan son of Eliashib. While he was there, he ate no food and drank no water, because he continued to mourn over the unfaithfulness of the exiles.
EZRA|10|7|A proclamation was then issued throughout Judah and Jerusalem for all the exiles to assemble in Jerusalem.
EZRA|10|8|Anyone who failed to appear within three days would forfeit all his property, in accordance with the decision of the officials and elders, and would himself be expelled from the assembly of the exiles.
EZRA|10|9|Within the three days, all the men of Judah and Benjamin had gathered in Jerusalem. And on the twentieth day of the ninth month, all the people were sitting in the square before the house of God, greatly distressed by the occasion and because of the rain.
EZRA|10|10|Then Ezra the priest stood up and said to them, "You have been unfaithful; you have married foreign women, adding to Israel's guilt.
EZRA|10|11|Now make confession to the LORD, the God of your fathers, and do his will. Separate yourselves from the peoples around you and from your foreign wives."
EZRA|10|12|The whole assembly responded with a loud voice: "You are right! We must do as you say.
EZRA|10|13|But there are many people here and it is the rainy season; so we cannot stand outside. Besides, this matter cannot be taken care of in a day or two, because we have sinned greatly in this thing.
EZRA|10|14|Let our officials act for the whole assembly. Then let everyone in our towns who has married a foreign woman come at a set time, along with the elders and judges of each town, until the fierce anger of our God in this matter is turned away from us."
EZRA|10|15|Only Jonathan son of Asahel and Jahzeiah son of Tikvah, supported by Meshullam and Shabbethai the Levite, opposed this.
EZRA|10|16|So the exiles did as was proposed. Ezra the priest selected men who were family heads, one from each family division, and all of them designated by name. On the first day of the tenth month they sat down to investigate the cases,
EZRA|10|17|and by the first day of the first month they finished dealing with all the men who had married foreign women.
EZRA|10|18|Among the descendants of the priests, the following had married foreign women: From the descendants of Jeshua son of Jozadak, and his brothers: Maaseiah, Eliezer, Jarib and Gedaliah.
EZRA|10|19|(They all gave their hands in pledge to put away their wives, and for their guilt they each presented a ram from the flock as a guilt offering.)
EZRA|10|20|From the descendants of Immer: Hanani and Zebadiah.
EZRA|10|21|From the descendants of Harim: Maaseiah, Elijah, Shemaiah, Jehiel and Uzziah.
EZRA|10|22|From the descendants of Pashhur: Elioenai, Maaseiah, Ishmael, Nethanel, Jozabad and Elasah.
EZRA|10|23|Among the Levites: Jozabad, Shimei, Kelaiah (that is, Kelita), Pethahiah, Judah and Eliezer.
EZRA|10|24|From the singers: Eliashib. From the gatekeepers: Shallum, Telem and Uri.
EZRA|10|25|And among the other Israelites: From the descendants of Parosh: Ramiah, Izziah, Malkijah, Mijamin, Eleazar, Malkijah and Benaiah.
EZRA|10|26|From the descendants of Elam: Mattaniah, Zechariah, Jehiel, Abdi, Jeremoth and Elijah.
EZRA|10|27|From the descendants of Zattu: Elioenai, Eliashib, Mattaniah, Jeremoth, Zabad and Aziza.
EZRA|10|28|From the descendants of Bebai: Jehohanan, Hananiah, Zabbai and Athlai.
EZRA|10|29|From the descendants of Bani: Meshullam, Malluch, Adaiah, Jashub, Sheal and Jeremoth.
EZRA|10|30|From the descendants of Pahath-Moab: Adna, Kelal, Benaiah, Maaseiah, Mattaniah, Bezalel, Binnui and Manasseh.
EZRA|10|31|From the descendants of Harim: Eliezer, Ishijah, Malkijah, Shemaiah, Shimeon,
EZRA|10|32|Benjamin, Malluch and Shemariah.
EZRA|10|33|From the descendants of Hashum: Mattenai, Mattattah, Zabad, Eliphelet, Jeremai, Manasseh and Shimei.
EZRA|10|34|From the descendants of Bani: Maadai, Amram, Uel,
EZRA|10|35|Benaiah, Bedeiah, Keluhi,
EZRA|10|36|Vaniah, Meremoth, Eliashib,
EZRA|10|37|Mattaniah, Mattenai and Jaasu.
EZRA|10|38|From the descendants of Binnui: Shimei,
EZRA|10|39|Shelemiah, Nathan, Adaiah,
EZRA|10|40|Macnadebai, Shashai, Sharai,
EZRA|10|41|Azarel, Shelemiah, Shemariah,
EZRA|10|42|Shallum, Amariah and Joseph.
EZRA|10|43|From the descendants of Nebo: Jeiel, Mattithiah, Zabad, Zebina, Jaddai, Joel and Benaiah.
EZRA|10|44|All these had married foreign women, and some of them had children by these wives.
