JONAH|1|1|Now the word of the LORD came to Jonah the son of Amittai, saying,
JONAH|1|2|"Arise, go to Nineveh, that great city, and call out against it, for their evil has come up before me."
JONAH|1|3|But Jonah rose to flee to Tarshish from the presence of the LORD. He went down to Joppa and found a ship going to Tarshish. So he paid the fare and went on board, to go with them to Tarshish, away from the presence of the LORD.
JONAH|1|4|But the LORD hurled a great wind upon the sea, and there was a mighty tempest on the sea, so that the ship threatened to break up.
JONAH|1|5|Then the mariners were afraid, and each cried out to his god. And they hurled the cargo that was in the ship into the sea to lighten it for them. But Jonah had gone down into the inner part of the ship and had lain down and was fast asleep.
JONAH|1|6|So the captain came and said to him, "What do you mean, you sleeper? Arise, call out to your god! Perhaps the god will give a thought to us, that we may not perish."
JONAH|1|7|And they said to one another, "Come, let us cast lots, that we may know on whose account this evil has come upon us." So they cast lots, and the lot fell on Jonah.
JONAH|1|8|Then they said to him, "Tell us on whose account this evil has come upon us. What is your occupation? And where do you come from? What is your country? And of what people are you?"
JONAH|1|9|And he said to them, "I am a Hebrew, and I fear the LORD, the God of heaven, who made the sea and the dry land."
JONAH|1|10|Then the men were exceedingly afraid and said to him, "What is this that you have done!" For the men knew that he was fleeing from the presence of the LORD, because he had told them.
JONAH|1|11|Then they said to him, "What shall we do to you, that the sea may quiet down for us?" For the sea grew more and more tempestuous.
JONAH|1|12|He said to them, "Pick me up and hurl me into the sea; then the sea will quiet down for you, for I know it is because of me that this great tempest has come upon you."
JONAH|1|13|Nevertheless, the men rowed hard to get back to dry land, but they could not, for the sea grew more and more tempestuous against them.
JONAH|1|14|Therefore they called out to the LORD, "O LORD, let us not perish for this man's life, and lay not on us innocent blood, for you, O LORD, have done as it pleased you."
JONAH|1|15|So they picked up Jonah and hurled him into the sea, and the sea ceased from its raging.
JONAH|1|16|Then the men feared the LORD exceedingly, and they offered a sacrifice to the LORD and made vows.
JONAH|1|17|And the LORD appointed a great fish to swallow up Jonah. And Jonah was in the belly of the fish three days and three nights.
JONAH|2|1|Then Jonah prayed to the LORD his God from the belly of the fish,
JONAH|2|2|saying, "I called out to the LORD, out of my distress, and he answered me; out of the belly of Sheol I cried, and you heard my voice.
JONAH|2|3|For you cast me into the deep, into the heart of the seas, and the flood surrounded me; all your waves and your billows passed over me.
JONAH|2|4|Then I said, 'I am driven away from your sight; Yet I shall again look upon your holy temple.'
JONAH|2|5|The waters closed in over me to take my life; the deep surrounded me; weeds were wrapped about my head
JONAH|2|6|at the roots of the mountains. I went down to the land whose bars closed upon me forever; yet you brought up my life from the pit, O LORD my God.
JONAH|2|7|When my life was fainting away, I remembered the LORD, and my prayer came to you, into your holy temple.
JONAH|2|8|Those who pay regard to vain idols forsake their hope of steadfast love.
JONAH|2|9|But I with the voice of thanksgiving will sacrifice to you; what I have vowed I will pay. Salvation belongs to the LORD!"
JONAH|2|10|And the LORD spoke to the fish, and it vomited Jonah out upon the dry land.
JONAH|3|1|Then the word of the LORD came to Jonah the second time, saying,
JONAH|3|2|"Arise, go to Nineveh, that great city, and call out against it the message that I tell you."
JONAH|3|3|So Jonah arose and went to Nineveh, according to the word of the LORD. Now Nineveh was an exceedingly great city, three days' journey in breadth.
JONAH|3|4|Jonah began to go into the city, going a day's journey. And he called out, "Yet forty days, and Nineveh shall be overthrown!"
JONAH|3|5|And the people of Nineveh believed God. They called for a fast and put on sackcloth, from the greatest of them to the least of them.
JONAH|3|6|The word reached the king of Nineveh, and he arose from his throne, removed his robe, covered himself with sackcloth, and sat in ashes.
JONAH|3|7|And he issued a proclamation and published through Nineveh, "By the decree of the king and his nobles: Let neither man nor beast, herd nor flock, taste anything. Let them not feed or drink water,
JONAH|3|8|but let man and beast be covered with sackcloth, and let them call out mightily to God. Let everyone turn from his evil way and from the violence that is in his hands.
JONAH|3|9|Who knows? God may turn and relent and turn from his fierce anger, so that we may not perish."
JONAH|3|10|When God saw what they did, how they turned from their evil way, God relented of the disaster that he had said he would do to them, and he did not do it.
JONAH|4|1|But it displeased Jonah exceedingly, and he was angry.
JONAH|4|2|And he prayed to the LORD and said, "O LORD, is not this what I said when I was yet in my country? That is why I made haste to flee to Tarshish; for I knew that you are a gracious God and merciful, slow to anger and abounding in steadfast love, and relenting from disaster.
JONAH|4|3|Therefore now, O LORD, please take my life from me, for it is better for me to die than to live."
JONAH|4|4|And the LORD said, "Do you do well to be angry?"
JONAH|4|5|Jonah went out of the city and sat to the east of the city and made a booth for himself there. He sat under it in the shade, till he should see what would become of the city.
JONAH|4|6|Now the LORD God appointed a plant and made it come up over Jonah, that it might be a shade over his head, to save him from his discomfort. So Jonah was exceedingly glad because of the plant.
JONAH|4|7|But when dawn came up the next day, God appointed a worm that attacked the plant, so that it withered.
JONAH|4|8|When the sun rose, God appointed a scorching east wind, and the sun beat down on the head of Jonah so that he was faint. And he asked that he might die and said, "It is better for me to die than to live."
JONAH|4|9|But God said to Jonah, "Do you do well to be angry for the plant?" And he said, "Yes, I do well to be angry, angry enough to die."
JONAH|4|10|And the LORD said, "You pity the plant, for which you did not labor, nor did you make it grow, which came into being in a night and perished in a night.
JONAH|4|11|And should not I pity Nineveh, that great city, in which there are more than 120,000 persons who do not know their right hand from their left, and also much cattle?"
