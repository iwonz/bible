1SAM|1|1|Now there was a certain man of Ramathaimzophim, of mount Ephraim, and his name was Elkanah, the son of Jeroham, the son of Elihu, the son of Tohu, the son of Zuph, an Ephrathite:
1SAM|1|2|And he had two wives; the name of the one was Hannah, and the name of the other Peninnah: and Peninnah had children, but Hannah had no children.
1SAM|1|3|And this man went up out of his city yearly to worship and to sacrifice unto the LORD of hosts in Shiloh. And the two sons of Eli, Hophni and Phinehas, the priests of the LORD, were there.
1SAM|1|4|And when the time was that Elkanah offered, he gave to Peninnah his wife, and to all her sons and her daughters, portions:
1SAM|1|5|But unto Hannah he gave a worthy portion; for he loved Hannah: but the LORD had shut up her womb.
1SAM|1|6|And her adversary also provoked her sore, for to make her fret, because the LORD had shut up her womb.
1SAM|1|7|And as he did so year by year, when she went up to the house of the LORD, so she provoked her; therefore she wept, and did not eat.
1SAM|1|8|Then said Elkanah her husband to her, Hannah, why weepest thou? and why eatest thou not? and why is thy heart grieved? am not I better to thee than ten sons?
1SAM|1|9|So Hannah rose up after they had eaten in Shiloh, and after they had drunk. Now Eli the priest sat upon a seat by a post of the temple of the LORD.
1SAM|1|10|And she was in bitterness of soul, and prayed unto the LORD, and wept sore.
1SAM|1|11|And she vowed a vow, and said, O LORD of hosts, if thou wilt indeed look on the affliction of thine handmaid, and remember me, and not forget thine handmaid, but wilt give unto thine handmaid a man child, then I will give him unto the LORD all the days of his life, and there shall no razor come upon his head.
1SAM|1|12|And it came to pass, as she continued praying before the LORD, that Eli marked her mouth.
1SAM|1|13|Now Hannah, she spake in her heart; only her lips moved, but her voice was not heard: therefore Eli thought she had been drunken.
1SAM|1|14|And Eli said unto her, How long wilt thou be drunken? put away thy wine from thee.
1SAM|1|15|And Hannah answered and said, No, my lord, I am a woman of a sorrowful spirit: I have drunk neither wine nor strong drink, but have poured out my soul before the LORD.
1SAM|1|16|Count not thine handmaid for a daughter of Belial: for out of the abundance of my complaint and grief have I spoken hitherto.
1SAM|1|17|Then Eli answered and said, Go in peace: and the God of Israel grant thee thy petition that thou hast asked of him.
1SAM|1|18|And she said, Let thine handmaid find grace in thy sight. So the woman went her way, and did eat, and her countenance was no more sad.
1SAM|1|19|And they rose up in the morning early, and worshipped before the LORD, and returned, and came to their house to Ramah: and Elkanah knew Hannah his wife; and the LORD remembered her.
1SAM|1|20|Wherefore it came to pass, when the time was come about after Hannah had conceived, that she bare a son, and called his name Samuel, saying, Because I have asked him of the LORD.
1SAM|1|21|And the man Elkanah, and all his house, went up to offer unto the LORD the yearly sacrifice, and his vow.
1SAM|1|22|But Hannah went not up; for she said unto her husband, I will not go up until the child be weaned, and then I will bring him, that he may appear before the LORD, and there abide for ever.
1SAM|1|23|And Elkanah her husband said unto her, Do what seemeth thee good; tarry until thou have weaned him; only the LORD establish his word. So the woman abode, and gave her son suck until she weaned him.
1SAM|1|24|And when she had weaned him, she took him up with her, with three bullocks, and one ephah of flour, and a bottle of wine, and brought him unto the house of the LORD in Shiloh: and the child was young.
1SAM|1|25|And they slew a bullock, and brought the child to Eli.
1SAM|1|26|And she said, Oh my lord, as thy soul liveth, my lord, I am the woman that stood by thee here, praying unto the LORD.
1SAM|1|27|For this child I prayed; and the LORD hath given me my petition which I asked of him:
1SAM|1|28|Therefore also I have lent him to the LORD; as long as he liveth he shall be lent to the LORD. And he worshipped the LORD there.
1SAM|2|1|And Hannah prayed, and said, My heart rejoiceth in the LORD, mine horn is exalted in the LORD: my mouth is enlarged over mine enemies; because I rejoice in thy salvation.
1SAM|2|2|There is none holy as the LORD: for there is none beside thee: neither is there any rock like our God.
1SAM|2|3|Talk no more so exceeding proudly; let not arrogancy come out of your mouth: for the LORD is a God of knowledge, and by him actions are weighed.
1SAM|2|4|The bows of the mighty men are broken, and they that stumbled are girded with strength.
1SAM|2|5|They that were full have hired out themselves for bread; and they that were hungry ceased: so that the barren hath born seven; and she that hath many children is waxed feeble.
1SAM|2|6|The LORD killeth, and maketh alive: he bringeth down to the grave, and bringeth up.
1SAM|2|7|The LORD maketh poor, and maketh rich: he bringeth low, and lifteth up.
1SAM|2|8|He raiseth up the poor out of the dust, and lifteth up the beggar from the dunghill, to set them among princes, and to make them inherit the throne of glory: for the pillars of the earth are the LORD's, and he hath set the world upon them.
1SAM|2|9|He will keep the feet of his saints, and the wicked shall be silent in darkness; for by strength shall no man prevail.
1SAM|2|10|The adversaries of the LORD shall be broken to pieces; out of heaven shall he thunder upon them: the LORD shall judge the ends of the earth; and he shall give strength unto his king, and exalt the horn of his anointed.
1SAM|2|11|And Elkanah went to Ramah to his house. And the child did minister unto the LORD before Eli the priest.
1SAM|2|12|Now the sons of Eli were sons of Belial; they knew not the LORD.
1SAM|2|13|And the priest's custom with the people was, that, when any man offered sacrifice, the priest's servant came, while the flesh was in seething, with a fleshhook of three teeth in his hand;
1SAM|2|14|And he struck it into the pan, or kettle, or caldron, or pot; all that the fleshhook brought up the priest took for himself. So they did in Shiloh unto all the Israelites that came thither.
1SAM|2|15|Also before they burnt the fat, the priest's servant came, and said to the man that sacrificed, Give flesh to roast for the priest; for he will not have sodden flesh of thee, but raw.
1SAM|2|16|And if any man said unto him, Let them not fail to burn the fat presently, and then take as much as thy soul desireth; then he would answer him, Nay; but thou shalt give it me now: and if not, I will take it by force.
1SAM|2|17|Wherefore the sin of the young men was very great before the LORD: for men abhorred the offering of the LORD.
1SAM|2|18|But Samuel ministered before the LORD, being a child, girded with a linen ephod.
1SAM|2|19|Moreover his mother made him a little coat, and brought it to him from year to year, when she came up with her husband to offer the yearly sacrifice.
1SAM|2|20|And Eli blessed Elkanah and his wife, and said, The LORD give thee seed of this woman for the loan which is lent to the LORD. And they went unto their own home.
1SAM|2|21|And the LORD visited Hannah, so that she conceived, and bare three sons and two daughters. And the child Samuel grew before the LORD.
1SAM|2|22|Now Eli was very old, and heard all that his sons did unto all Israel; and how they lay with the women that assembled at the door of the tabernacle of the congregation.
1SAM|2|23|And he said unto them, Why do ye such things? for I hear of your evil dealings by all this people.
1SAM|2|24|Nay, my sons; for it is no good report that I hear: ye make the LORD's people to transgress.
1SAM|2|25|If one man sin against another, the judge shall judge him: but if a man sin against the LORD, who shall entreat for him? Notwithstanding they hearkened not unto the voice of their father, because the LORD would slay them.
1SAM|2|26|And the child Samuel grew on, and was in favor both with the LORD, and also with men.
1SAM|2|27|And there came a man of God unto Eli, and said unto him, Thus saith the LORD, Did I plainly appear unto the house of thy father, when they were in Egypt in Pharaoh's house?
1SAM|2|28|And did I choose him out of all the tribes of Israel to be my priest, to offer upon mine altar, to burn incense, to wear an ephod before me? and did I give unto the house of thy father all the offerings made by fire of the children of Israel?
1SAM|2|29|Wherefore kick ye at my sacrifice and at mine offering, which I have commanded in my habitation; and honorest thy sons above me, to make yourselves fat with the chiefest of all the offerings of Israel my people?
1SAM|2|30|Wherefore the LORD God of Israel saith, I said indeed that thy house, and the house of thy father, should walk before me for ever: but now the LORD saith, Be it far from me; for them that honor me I will honor, and they that despise me shall be lightly esteemed.
1SAM|2|31|Behold, the days come, that I will cut off thine arm, and the arm of thy father's house, that there shall not be an old man in thine house.
1SAM|2|32|And thou shalt see an enemy in my habitation, in all the wealth which God shall give Israel: and there shall not be an old man in thine house for ever.
1SAM|2|33|And the man of thine, whom I shall not cut off from mine altar, shall be to consume thine eyes, and to grieve thine heart: and all the increase of thine house shall die in the flower of their age.
1SAM|2|34|And this shall be a sign unto thee, that shall come upon thy two sons, on Hophni and Phinehas; in one day they shall die both of them.
1SAM|2|35|And I will raise me up a faithful priest, that shall do according to that which is in mine heart and in my mind: and I will build him a sure house; and he shall walk before mine anointed for ever.
1SAM|2|36|And it shall come to pass, that every one that is left in thine house shall come and crouch to him for a piece of silver and a morsel of bread, and shall say, Put me, I pray thee, into one of the priests' offices, that I may eat a piece of bread.
1SAM|3|1|And the child Samuel ministered unto the LORD before Eli. And the word of the LORD was precious in those days; there was no open vision.
1SAM|3|2|And it came to pass at that time, when Eli was laid down in his place, and his eyes began to wax dim, that he could not see;
1SAM|3|3|And ere the lamp of God went out in the temple of the LORD, where the ark of God was, and Samuel was laid down to sleep;
1SAM|3|4|That the LORD called Samuel: and he answered, Here am I.
1SAM|3|5|And he ran unto Eli, and said, Here am I; for thou calledst me. And he said, I called not; lie down again. And he went and lay down.
1SAM|3|6|And the LORD called yet again, Samuel. And Samuel arose and went to Eli, and said, Here am I; for thou didst call me. And he answered, I called not, my son; lie down again.
1SAM|3|7|Now Samuel did not yet know the LORD, neither was the word of the LORD yet revealed unto him.
1SAM|3|8|And the LORD called Samuel again the third time. And he arose and went to Eli, and said, Here am I; for thou didst call me. And Eli perceived that the LORD had called the child.
1SAM|3|9|Therefore Eli said unto Samuel, Go, lie down: and it shall be, if he call thee, that thou shalt say, Speak, LORD; for thy servant heareth. So Samuel went and lay down in his place.
1SAM|3|10|And the LORD came, and stood, and called as at other times, Samuel, Samuel. Then Samuel answered, Speak; for thy servant heareth.
1SAM|3|11|And the LORD said to Samuel, Behold, I will do a thing in Israel, at which both the ears of every one that heareth it shall tingle.
1SAM|3|12|In that day I will perform against Eli all things which I have spoken concerning his house: when I begin, I will also make an end.
1SAM|3|13|For I have told him that I will judge his house for ever for the iniquity which he knoweth; because his sons made themselves vile, and he restrained them not.
1SAM|3|14|And therefore I have sworn unto the house of Eli, that the iniquity of Eli's house shall not be purged with sacrifice nor offering for ever.
1SAM|3|15|And Samuel lay until the morning, and opened the doors of the house of the LORD. And Samuel feared to show Eli the vision.
1SAM|3|16|Then Eli called Samuel, and said, Samuel, my son. And he answered, Here am I.
1SAM|3|17|And he said, What is the thing that the LORD hath said unto thee? I pray thee hide it not from me: God do so to thee, and more also, if thou hide any thing from me of all the things that he said unto thee.
1SAM|3|18|And Samuel told him every whit, and hid nothing from him. And he said, It is the LORD: let him do what seemeth him good.
1SAM|3|19|And Samuel grew, and the LORD was with him, and did let none of his words fall to the ground.
1SAM|3|20|And all Israel from Dan even to Beersheba knew that Samuel was established to be a prophet of the LORD.
1SAM|3|21|And the LORD appeared again in Shiloh: for the LORD revealed himself to Samuel in Shiloh by the word of the LORD.
1SAM|4|1|And the word of Samuel came to all Israel. Now Israel went out against the Philistines to battle, and pitched beside Ebenezer: and the Philistines pitched in Aphek.
1SAM|4|2|And the Philistines put themselves in array against Israel: and when they joined battle, Israel was smitten before the Philistines: and they slew of the army in the field about four thousand men.
1SAM|4|3|And when the people were come into the camp, the elders of Israel said, Wherefore hath the LORD smitten us to day before the Philistines? Let us fetch the ark of the covenant of the LORD out of Shiloh unto us, that, when it cometh among us, it may save us out of the hand of our enemies.
1SAM|4|4|So the people sent to Shiloh, that they might bring from thence the ark of the covenant of the LORD of hosts, which dwelleth between the cherubim: and the two sons of Eli, Hophni and Phinehas, were there with the ark of the covenant of God.
1SAM|4|5|And when the ark of the covenant of the LORD came into the camp, all Israel shouted with a great shout, so that the earth rang again.
1SAM|4|6|And when the Philistines heard the noise of the shout, they said, What meaneth the noise of this great shout in the camp of the Hebrews? And they understood that the ark of the LORD was come into the camp.
1SAM|4|7|And the Philistines were afraid, for they said, God is come into the camp. And they said, Woe unto us! for there hath not been such a thing heretofore.
1SAM|4|8|Woe unto us! who shall deliver us out of the hand of these mighty Gods? these are the Gods that smote the Egyptians with all the plagues in the wilderness.
1SAM|4|9|Be strong and quit yourselves like men, O ye Philistines, that ye be not servants unto the Hebrews, as they have been to you: quit yourselves like men, and fight.
1SAM|4|10|And the Philistines fought, and Israel was smitten, and they fled every man into his tent: and there was a very great slaughter; for there fell of Israel thirty thousand footmen.
1SAM|4|11|And the ark of God was taken; and the two sons of Eli, Hophni and Phinehas, were slain.
1SAM|4|12|And there ran a man of Benjamin out of the army, and came to Shiloh the same day with his clothes rent, and with earth upon his head.
1SAM|4|13|And when he came, lo, Eli sat upon a seat by the wayside watching: for his heart trembled for the ark of God. And when the man came into the city, and told it, all the city cried out.
1SAM|4|14|And when Eli heard the noise of the crying, he said, What meaneth the noise of this tumult? And the man came in hastily, and told Eli.
1SAM|4|15|Now Eli was ninety and eight years old; and his eyes were dim, that he could not see.
1SAM|4|16|And the man said unto Eli, I am he that came out of the army, and I fled to day out of the army. And he said, What is there done, my son?
1SAM|4|17|And the messenger answered and said, Israel is fled before the Philistines, and there hath been also a great slaughter among the people, and thy two sons also, Hophni and Phinehas, are dead, and the ark of God is taken.
1SAM|4|18|And it came to pass, when he made mention of the ark of God, that he fell from off the seat backward by the side of the gate, and his neck brake, and he died: for he was an old man, and heavy. And he had judged Israel forty years.
1SAM|4|19|And his daughter in law, Phinehas' wife, was with child, near to be delivered: and when she heard the tidings that the ark of God was taken, and that her father in law and her husband were dead, she bowed herself and travailed; for her pains came upon her.
1SAM|4|20|And about the time of her death the women that stood by her said unto her, Fear not; for thou hast born a son. But she answered not, neither did she regard it.
1SAM|4|21|And she named the child Ichabod, saying, The glory is departed from Israel: because the ark of God was taken, and because of her father in law and her husband.
1SAM|4|22|And she said, The glory is departed from Israel: for the ark of God is taken.
1SAM|5|1|And the Philistines took the ark of God, and brought it from Ebenezer unto Ashdod.
1SAM|5|2|When the Philistines took the ark of God, they brought it into the house of Dagon, and set it by Dagon.
1SAM|5|3|And when they of Ashdod arose early on the morrow, behold, Dagon was fallen upon his face to the earth before the ark of the LORD. And they took Dagon, and set him in his place again.
1SAM|5|4|And when they arose early on the morrow morning, behold, Dagon was fallen upon his face to the ground before the ark of the LORD; and the head of Dagon and both the palms of his hands were cut off upon the threshold; only the stump of Dagon was left to him.
1SAM|5|5|Therefore neither the priests of Dagon, nor any that come into Dagon's house, tread on the threshold of Dagon in Ashdod unto this day.
1SAM|5|6|But the hand of the LORD was heavy upon them of Ashdod, and he destroyed them, and smote them with emerods, even Ashdod and the coasts thereof.
1SAM|5|7|And when the men of Ashdod saw that it was so, they said, The ark of the God of Israel shall not abide with us: for his hand is sore upon us, and upon Dagon our god.
1SAM|5|8|They sent therefore and gathered all the lords of the Philistines unto them, and said, What shall we do with the ark of the God of Israel? And they answered, Let the ark of the God of Israel be carried about unto Gath. And they carried the ark of the God of Israel about thither.
1SAM|5|9|And it was so, that, after they had carried it about, the hand of the LORD was against the city with a very great destruction: and he smote the men of the city, both small and great, and they had emerods in their secret parts.
1SAM|5|10|Therefore they sent the ark of God to Ekron. And it came to pass, as the ark of God came to Ekron, that the Ekronites cried out, saying, They have brought about the ark of the God of Israel to us, to slay us and our people.
1SAM|5|11|So they sent and gathered together all the lords of the Philistines, and said, Send away the ark of the God of Israel, and let it go again to his own place, that it slay us not, and our people: for there was a deadly destruction throughout all the city; the hand of God was very heavy there.
1SAM|5|12|And the men that died not were smitten with the emerods: and the cry of the city went up to heaven.
1SAM|6|1|And the ark of the LORD was in the country of the Philistines seven months.
1SAM|6|2|And the Philistines called for the priests and the diviners, saying, What shall we do to the ark of the LORD? tell us wherewith we shall send it to his place.
1SAM|6|3|And they said, If ye send away the ark of the God of Israel, send it not empty; but in any wise return him a trespass offering: then ye shall be healed, and it shall be known to you why his hand is not removed from you.
1SAM|6|4|Then said they, What shall be the trespass offering which we shall return to him? They answered, Five golden emerods, and five golden mice, according to the number of the lords of the Philistines: for one plague was on you all, and on your lords.
1SAM|6|5|Wherefore ye shall make images of your emerods, and images of your mice that mar the land; and ye shall give glory unto the God of Israel: peradventure he will lighten his hand from off you, and from off your gods, and from off your land.
1SAM|6|6|Wherefore then do ye harden your hearts, as the Egyptians and Pharaoh hardened their hearts? when he had wrought wonderfully among them, did they not let the people go, and they departed?
1SAM|6|7|Now therefore make a new cart, and take two milch kine, on which there hath come no yoke, and tie the kine to the cart, and bring their calves home from them:
1SAM|6|8|And take the ark of the LORD, and lay it upon the cart; and put the jewels of gold, which ye return him for a trespass offering, in a coffer by the side thereof; and send it away, that it may go.
1SAM|6|9|And see, if it goeth up by the way of his own coast to Bethshemesh, then he hath done us this great evil: but if not, then we shall know that it is not his hand that smote us: it was a chance that happened to us.
1SAM|6|10|And the men did so; and took two milch kine, and tied them to the cart, and shut up their calves at home:
1SAM|6|11|And they laid the ark of the LORD upon the cart, and the coffer with the mice of gold and the images of their emerods.
1SAM|6|12|And the kine took the straight way to the way of Bethshemesh, and went along the highway, lowing as they went, and turned not aside to the right hand or to the left; and the lords of the Philistines went after them unto the border of Bethshemesh.
1SAM|6|13|And they of Bethshemesh were reaping their wheat harvest in the valley: and they lifted up their eyes, and saw the ark, and rejoiced to see it.
1SAM|6|14|And the cart came into the field of Joshua, a Bethshemite, and stood there, where there was a great stone: and they clave the wood of the cart, and offered the kine a burnt offering unto the LORD.
1SAM|6|15|And the Levites took down the ark of the LORD, and the coffer that was with it, wherein the jewels of gold were, and put them on the great stone: and the men of Bethshemesh offered burnt offerings and sacrificed sacrifices the same day unto the LORD.
1SAM|6|16|And when the five lords of the Philistines had seen it, they returned to Ekron the same day.
1SAM|6|17|And these are the golden emerods which the Philistines returned for a trespass offering unto the LORD; for Ashdod one, for Gaza one, for Askelon one, for Gath one, for Ekron one;
1SAM|6|18|And the golden mice, according to the number of all the cities of the Philistines belonging to the five lords, both of fenced cities, and of country villages, even unto the great stone of Abel, whereon they set down the ark of the LORD: which stone remaineth unto this day in the field of Joshua, the Bethshemite.
1SAM|6|19|And he smote the men of Bethshemesh, because they had looked into the ark of the LORD, even he smote of the people fifty thousand and threescore and ten men: and the people lamented, because the LORD had smitten many of the people with a great slaughter.
1SAM|6|20|And the men of Bethshemesh said, Who is able to stand before this holy LORD God? and to whom shall he go up from us?
1SAM|6|21|And they sent messengers to the inhabitants of Kirjathjearim, saying, The Philistines have brought again the ark of the LORD; come ye down, and fetch it up to you.
1SAM|7|1|And the men of Kirjathjearim came, and fetched up the ark of the LORD, and brought it into the house of Abinadab in the hill, and sanctified Eleazar his son to keep the ark of the LORD.
1SAM|7|2|And it came to pass, while the ark abode in Kirjathjearim, that the time was long; for it was twenty years: and all the house of Israel lamented after the LORD.
1SAM|7|3|And Samuel spake unto all the house of Israel, saying, If ye do return unto the LORD with all your hearts, then put away the strange gods and Ashtaroth from among you, and prepare your hearts unto the LORD, and serve him only: and he will deliver you out of the hand of the Philistines.
1SAM|7|4|Then the children of Israel did put away Baalim and Ashtaroth, and served the LORD only.
1SAM|7|5|And Samuel said, Gather all Israel to Mizpeh, and I will pray for you unto the LORD.
1SAM|7|6|And they gathered together to Mizpeh, and drew water, and poured it out before the LORD, and fasted on that day, and said there, We have sinned against the LORD. And Samuel judged the children of Israel in Mizpeh.
1SAM|7|7|And when the Philistines heard that the children of Israel were gathered together to Mizpeh, the lords of the Philistines went up against Israel. And when the children of Israel heard it, they were afraid of the Philistines.
1SAM|7|8|And the children of Israel said to Samuel, Cease not to cry unto the LORD our God for us, that he will save us out of the hand of the Philistines.
1SAM|7|9|And Samuel took a sucking lamb, and offered it for a burnt offering wholly unto the LORD: and Samuel cried unto the LORD for Israel; and the LORD heard him.
1SAM|7|10|And as Samuel was offering up the burnt offering, the Philistines drew near to battle against Israel: but the LORD thundered with a great thunder on that day upon the Philistines, and discomfited them; and they were smitten before Israel.
1SAM|7|11|And the men of Israel went out of Mizpeh, and pursued the Philistines, and smote them, until they came under Bethcar.
1SAM|7|12|Then Samuel took a stone, and set it between Mizpeh and Shen, and called the name of it Ebenezer, saying, Hitherto hath the LORD helped us.
1SAM|7|13|So the Philistines were subdued, and they came no more into the coast of Israel: and the hand of the LORD was against the Philistines all the days of Samuel.
1SAM|7|14|And the cities which the Philistines had taken from Israel were restored to Israel, from Ekron even unto Gath; and the coasts thereof did Israel deliver out of the hands of the Philistines. And there was peace between Israel and the Amorites.
1SAM|7|15|And Samuel judged Israel all the days of his life.
1SAM|7|16|And he went from year to year in circuit to Bethel, and Gilgal, and Mizpeh, and judged Israel in all those places.
1SAM|7|17|And his return was to Ramah; for there was his house; and there he judged Israel; and there he built an altar unto the LORD.
1SAM|8|1|And it came to pass, when Samuel was old, that he made his sons judges over Israel.
1SAM|8|2|Now the name of his firstborn was Joel; and the name of his second, Abiah: they were judges in Beersheba.
1SAM|8|3|And his sons walked not in his ways, but turned aside after lucre, and took bribes, and perverted judgment.
1SAM|8|4|Then all the elders of Israel gathered themselves together, and came to Samuel unto Ramah,
1SAM|8|5|And said unto him, Behold, thou art old, and thy sons walk not in thy ways: now make us a king to judge us like all the nations.
1SAM|8|6|But the thing displeased Samuel, when they said, Give us a king to judge us. And Samuel prayed unto the LORD.
1SAM|8|7|And the LORD said unto Samuel, Hearken unto the voice of the people in all that they say unto thee: for they have not rejected thee, but they have rejected me, that I should not reign over them.
1SAM|8|8|According to all the works which they have done since the day that I brought them up out of Egypt even unto this day, wherewith they have forsaken me, and served other gods, so do they also unto thee.
1SAM|8|9|Now therefore hearken unto their voice: howbeit yet protest solemnly unto them, and show them the manner of the king that shall reign over them.
1SAM|8|10|And Samuel told all the words of the LORD unto the people that asked of him a king.
1SAM|8|11|And he said, This will be the manner of the king that shall reign over you: He will take your sons, and appoint them for himself, for his chariots, and to be his horsemen; and some shall run before his chariots.
1SAM|8|12|And he will appoint him captains over thousands, and captains over fifties; and will set them to ear his ground, and to reap his harvest, and to make his instruments of war, and instruments of his chariots.
1SAM|8|13|And he will take your daughters to be confectionaries, and to be cooks, and to be bakers.
1SAM|8|14|And he will take your fields, and your vineyards, and your oliveyards, even the best of them, and give them to his servants.
1SAM|8|15|And he will take the tenth of your seed, and of your vineyards, and give to his officers, and to his servants.
1SAM|8|16|And he will take your menservants, and your maidservants, and your goodliest young men, and your asses, and put them to his work.
1SAM|8|17|He will take the tenth of your sheep: and ye shall be his servants.
1SAM|8|18|And ye shall cry out in that day because of your king which ye shall have chosen you; and the LORD will not hear you in that day.
1SAM|8|19|Nevertheless the people refused to obey the voice of Samuel; and they said, Nay; but we will have a king over us;
1SAM|8|20|That we also may be like all the nations; and that our king may judge us, and go out before us, and fight our battles.
1SAM|8|21|And Samuel heard all the words of the people, and he rehearsed them in the ears of the LORD.
1SAM|8|22|And the LORD said to Samuel, Hearken unto their voice, and make them a king. And Samuel said unto the men of Israel, Go ye every man unto his city.
1SAM|9|1|Now there was a man of Benjamin, whose name was Kish, the son of Abiel, the son of Zeror, the son of Bechorath, the son of Aphiah, a Benjamite, a mighty man of power.
1SAM|9|2|And he had a son, whose name was Saul, a choice young man, and a goodly: and there was not among the children of Israel a goodlier person than he: from his shoulders and upward he was higher than any of the people.
1SAM|9|3|And the asses of Kish Saul's father were lost. And Kish said to Saul his son, Take now one of the servants with thee, and arise, go seek the asses.
1SAM|9|4|And he passed through mount Ephraim, and passed through the land of Shalisha, but they found them not: then they passed through the land of Shalim, and there they were not: and he passed through the land of the Benjamites, but they found them not.
1SAM|9|5|And when they were come to the land of Zuph, Saul said to his servant that was with him, Come, and let us return; lest my father leave caring for the asses, and take thought for us.
1SAM|9|6|And he said unto him, Behold now, there is in this city a man of God, and he is an honorable man; all that he saith cometh surely to pass: now let us go thither; peradventure he can show us our way that we should go.
1SAM|9|7|Then said Saul to his servant, But, behold, if we go, what shall we bring the man? for the bread is spent in our vessels, and there is not a present to bring to the man of God: what have we?
1SAM|9|8|And the servant answered Saul again, and said, Behold, I have here at hand the fourth part of a shekel of silver: that will I give to the man of God, to tell us our way.
1SAM|9|9|(Beforetime in Israel, when a man went to inquire of God, thus he spake, Come, and let us go to the seer: for he that is now called a Prophet was beforetime called a Seer.)
1SAM|9|10|Then said Saul to his servant, Well said; come, let us go. So they went unto the city where the man of God was.
1SAM|9|11|And as they went up the hill to the city, they found young maidens going out to draw water, and said unto them, Is the seer here?
1SAM|9|12|And they answered them, and said, He is; behold, he is before you: make haste now, for he came to day to the city; for there is a sacrifice of the people to day in the high place:
1SAM|9|13|As soon as ye be come into the city, ye shall straightway find him, before he go up to the high place to eat: for the people will not eat until he come, because he doth bless the sacrifice; and afterwards they eat that be bidden. Now therefore get you up; for about this time ye shall find him.
1SAM|9|14|And they went up into the city: and when they were come into the city, behold, Samuel came out against them, for to go up to the high place.
1SAM|9|15|Now the LORD had told Samuel in his ear a day before Saul came, saying,
1SAM|9|16|To morrow about this time I will send thee a man out of the land of Benjamin, and thou shalt anoint him to be captain over my people Israel, that he may save my people out of the hand of the Philistines: for I have looked upon my people, because their cry is come unto me.
1SAM|9|17|And when Samuel saw Saul, the LORD said unto him, Behold the man whom I spake to thee of! this same shall reign over my people.
1SAM|9|18|Then Saul drew near to Samuel in the gate, and said, Tell me, I pray thee, where the seer's house is.
1SAM|9|19|And Samuel answered Saul, and said, I am the seer: go up before me unto the high place; for ye shall eat with me to day, and to morrow I will let thee go, and will tell thee all that is in thine heart.
1SAM|9|20|And as for thine asses that were lost three days ago, set not thy mind on them; for they are found. And on whom is all the desire of Israel? Is it not on thee, and on all thy father's house?
1SAM|9|21|And Saul answered and said, Am not I a Benjamite, of the smallest of the tribes of Israel? and my family the least of all the families of the tribe of Benjamin? wherefore then speakest thou so to me?
1SAM|9|22|And Samuel took Saul and his servant, and brought them into the parlor, and made them sit in the chiefest place among them that were bidden, which were about thirty persons.
1SAM|9|23|And Samuel said unto the cook, Bring the portion which I gave thee, of which I said unto thee, Set it by thee.
1SAM|9|24|And the cook took up the shoulder, and that which was upon it, and set it before Saul. And Samuel said, Behold that which is left! set it before thee, and eat: for unto this time hath it been kept for thee since I said, I have invited the people. So Saul did eat with Samuel that day.
1SAM|9|25|And when they were come down from the high place into the city, Samuel communed with Saul upon the top of the house.
1SAM|9|26|And they arose early: and it came to pass about the spring of the day, that Samuel called Saul to the top of the house, saying, Up, that I may send thee away. And Saul arose, and they went out both of them, he and Samuel, abroad.
1SAM|9|27|And as they were going down to the end of the city, Samuel said to Saul, Bid the servant pass on before us, (and he passed on), but stand thou still a while, that I may show thee the word of God.
1SAM|10|1|Then Samuel took a vial of oil, and poured it upon his head, and kissed him, and said, Is it not because the LORD hath anointed thee to be captain over his inheritance?
1SAM|10|2|When thou art departed from me to day, then thou shalt find two men by Rachel's sepulchre in the border of Benjamin at Zelzah; and they will say unto thee, The asses which thou wentest to seek are found: and, lo, thy father hath left the care of the asses, and sorroweth for you, saying, What shall I do for my son?
1SAM|10|3|Then shalt thou go on forward from thence, and thou shalt come to the plain of Tabor, and there shall meet thee three men going up to God to Bethel, one carrying three kids, and another carrying three loaves of bread, and another carrying a bottle of wine:
1SAM|10|4|And they will salute thee, and give thee two loaves of bread; which thou shalt receive of their hands.
1SAM|10|5|After that thou shalt come to the hill of God, where is the garrison of the Philistines: and it shall come to pass, when thou art come thither to the city, that thou shalt meet a company of prophets coming down from the high place with a psaltery, and a tabret, and a pipe, and a harp, before them; and they shall prophesy:
1SAM|10|6|And the Spirit of the LORD will come upon thee, and thou shalt prophesy with them, and shalt be turned into another man.
1SAM|10|7|And let it be, when these signs are come unto thee, that thou do as occasion serve thee; for God is with thee.
1SAM|10|8|And thou shalt go down before me to Gilgal; and, behold, I will come down unto thee, to offer burnt offerings, and to sacrifice sacrifices of peace offerings: seven days shalt thou tarry, till I come to thee, and show thee what thou shalt do.
1SAM|10|9|And it was so, that when he had turned his back to go from Samuel, God gave him another heart: and all those signs came to pass that day.
1SAM|10|10|And when they came thither to the hill, behold, a company of prophets met him; and the Spirit of God came upon him, and he prophesied among them.
1SAM|10|11|And it came to pass, when all that knew him beforetime saw that, behold, he prophesied among the prophets, then the people said one to another, What is this that is come unto the son of Kish? Is Saul also among the prophets?
1SAM|10|12|And one of the same place answered and said, But who is their father? Therefore it became a proverb, Is Saul also among the prophets?
1SAM|10|13|And when he had made an end of prophesying, he came to the high place.
1SAM|10|14|And Saul's uncle said unto him and to his servant, Whither went ye? And he said, To seek the asses: and when we saw that they were no where, we came to Samuel.
1SAM|10|15|And Saul's uncle said, Tell me, I pray thee, what Samuel said unto you.
1SAM|10|16|And Saul said unto his uncle, He told us plainly that the asses were found. But of the matter of the kingdom, whereof Samuel spake, he told him not.
1SAM|10|17|And Samuel called the people together unto the LORD to Mizpeh;
1SAM|10|18|And said unto the children of Israel, Thus saith the LORD God of Israel, I brought up Israel out of Egypt, and delivered you out of the hand of the Egyptians, and out of the hand of all kingdoms, and of them that oppressed you:
1SAM|10|19|And ye have this day rejected your God, who himself saved you out of all your adversities and your tribulations; and ye have said unto him, Nay, but set a king over us. Now therefore present yourselves before the LORD by your tribes, and by your thousands.
1SAM|10|20|And when Samuel had caused all the tribes of Israel to come near, the tribe of Benjamin was taken.
1SAM|10|21|When he had caused the tribe of Benjamin to come near by their families, the family of Matri was taken, and Saul the son of Kish was taken: and when they sought him, he could not be found.
1SAM|10|22|Therefore they inquired of the LORD further, if the man should yet come thither. And the LORD answered, Behold he hath hid himself among the stuff.
1SAM|10|23|And they ran and fetched him thence: and when he stood among the people, he was higher than any of the people from his shoulders and upward.
1SAM|10|24|And Samuel said to all the people, See ye him whom the LORD hath chosen, that there is none like him among all the people? And all the people shouted, and said, God save the king.
1SAM|10|25|Then Samuel told the people the manner of the kingdom, and wrote it in a book, and laid it up before the LORD. And Samuel sent all the people away, every man to his house.
1SAM|10|26|And Saul also went home to Gibeah; and there went with him a band of men, whose hearts God had touched.
1SAM|10|27|But the children of Belial said, How shall this man save us? And they despised him, and brought no presents. But he held his peace.
1SAM|11|1|Then Nahash the Ammonite came up, and encamped against Jabeshgilead: and all the men of Jabesh said unto Nahash, Make a covenant with us, and we will serve thee.
1SAM|11|2|And Nahash the Ammonite answered them, On this condition will I make a covenant with you, that I may thrust out all your right eyes, and lay it for a reproach upon all Israel.
1SAM|11|3|And the elders of Jabesh said unto him, Give us seven days' respite, that we may send messengers unto all the coasts of Israel: and then, if there be no man to save us, we will come out to thee.
1SAM|11|4|Then came the messengers to Gibeah of Saul, and told the tidings in the ears of the people: and all the people lifted up their voices, and wept.
1SAM|11|5|And, behold, Saul came after the herd out of the field; and Saul said, What aileth the people that they weep? And they told him the tidings of the men of Jabesh.
1SAM|11|6|And the Spirit of God came upon Saul when he heard those tidings, and his anger was kindled greatly.
1SAM|11|7|And he took a yoke of oxen, and hewed them in pieces, and sent them throughout all the coasts of Israel by the hands of messengers, saying, Whosoever cometh not forth after Saul and after Samuel, so shall it be done unto his oxen. And the fear of the LORD fell on the people, and they came out with one consent.
1SAM|11|8|And when he numbered them in Bezek, the children of Israel were three hundred thousand, and the men of Judah thirty thousand.
1SAM|11|9|And they said unto the messengers that came, Thus shall ye say unto the men of Jabeshgilead, To morrow, by that time the sun be hot, ye shall have help. And the messengers came and showed it to the men of Jabesh; and they were glad.
1SAM|11|10|Therefore the men of Jabesh said, To morrow we will come out unto you, and ye shall do with us all that seemeth good unto you.
1SAM|11|11|And it was so on the morrow, that Saul put the people in three companies; and they came into the midst of the host in the morning watch, and slew the Ammonites until the heat of the day: and it came to pass, that they which remained were scattered, so that two of them were not left together.
1SAM|11|12|And the people said unto Samuel, Who is he that said, Shall Saul reign over us? bring the men, that we may put them to death.
1SAM|11|13|And Saul said, There shall not a man be put to death this day: for to day the LORD hath wrought salvation in Israel.
1SAM|11|14|Then said Samuel to the people, Come, and let us go to Gilgal, and renew the kingdom there.
1SAM|11|15|And all the people went to Gilgal; and there they made Saul king before the LORD in Gilgal; and there they sacrificed sacrifices of peace offerings before the LORD; and there Saul and all the men of Israel rejoiced greatly.
1SAM|12|1|And Samuel said unto all Israel, Behold, I have hearkened unto your voice in all that ye said unto me, and have made a king over you.
1SAM|12|2|And now, behold, the king walketh before you: and I am old and grayheaded; and, behold, my sons are with you: and I have walked before you from my childhood unto this day.
1SAM|12|3|Behold, here I am: witness against me before the LORD, and before his anointed: whose ox have I taken? or whose ass have I taken? or whom have I defrauded? whom have I oppressed? or of whose hand have I received any bribe to blind mine eyes therewith? and I will restore it you.
1SAM|12|4|And they said, Thou hast not defrauded us, nor oppressed us, neither hast thou taken ought of any man's hand.
1SAM|12|5|And he said unto them, The LORD is witness against you, and his anointed is witness this day, that ye have not found ought in my hand. And they answered, He is witness.
1SAM|12|6|And Samuel said unto the people, It is the LORD that advanced Moses and Aaron, and that brought your fathers up out of the land of Egypt.
1SAM|12|7|Now therefore stand still, that I may reason with you before the LORD of all the righteous acts of the LORD, which he did to you and to your fathers.
1SAM|12|8|When Jacob was come into Egypt, and your fathers cried unto the LORD, then the LORD sent Moses and Aaron, which brought forth your fathers out of Egypt, and made them dwell in this place.
1SAM|12|9|And when they forgat the LORD their God, he sold them into the hand of Sisera, captain of the host of Hazor, and into the hand of the Philistines, and into the hand of the king of Moab, and they fought against them.
1SAM|12|10|And they cried unto the LORD, and said, We have sinned, because we have forsaken the LORD, and have served Baalim and Ashtaroth: but now deliver us out of the hand of our enemies, and we will serve thee.
1SAM|12|11|And the LORD sent Jerubbaal, and Bedan, and Jephthah, and Samuel, and delivered you out of the hand of your enemies on every side, and ye dwelled safe.
1SAM|12|12|And when ye saw that Nahash the king of the children of Ammon came against you, ye said unto me, Nay; but a king shall reign over us: when the LORD your God was your king.
1SAM|12|13|Now therefore behold the king whom ye have chosen, and whom ye have desired! and, behold, the LORD hath set a king over you.
1SAM|12|14|If ye will fear the LORD, and serve him, and obey his voice, and not rebel against the commandment of the LORD, then shall both ye and also the king that reigneth over you continue following the LORD your God:
1SAM|12|15|But if ye will not obey the voice of the LORD, but rebel against the commandment of the LORD, then shall the hand of the LORD be against you, as it was against your fathers.
1SAM|12|16|Now therefore stand and see this great thing, which the LORD will do before your eyes.
1SAM|12|17|Is it not wheat harvest to day? I will call unto the LORD, and he shall send thunder and rain; that ye may perceive and see that your wickedness is great, which ye have done in the sight of the LORD, in asking you a king.
1SAM|12|18|So Samuel called unto the LORD; and the LORD sent thunder and rain that day: and all the people greatly feared the LORD and Samuel.
1SAM|12|19|And all the people said unto Samuel, Pray for thy servants unto the LORD thy God, that we die not: for we have added unto all our sins this evil, to ask us a king.
1SAM|12|20|And Samuel said unto the people, Fear not: ye have done all this wickedness: yet turn not aside from following the LORD, but serve the LORD with all your heart;
1SAM|12|21|And turn ye not aside: for then should ye go after vain things, which cannot profit nor deliver; for they are vain.
1SAM|12|22|For the LORD will not forsake his people for his great name's sake: because it hath pleased the LORD to make you his people.
1SAM|12|23|Moreover as for me, God forbid that I should sin against the LORD in ceasing to pray for you: but I will teach you the good and the right way:
1SAM|12|24|Only fear the LORD, and serve him in truth with all your heart: for consider how great things he hath done for you.
1SAM|12|25|But if ye shall still do wickedly, ye shall be consumed, both ye and your king.
1SAM|13|1|Saul reigned one year; and when he had reigned two years over Israel,
1SAM|13|2|Saul chose him three thousand men of Israel; whereof two thousand were with Saul in Michmash and in mount Bethel, and a thousand were with Jonathan in Gibeah of Benjamin: and the rest of the people he sent every man to his tent.
1SAM|13|3|And Jonathan smote the garrison of the Philistines that was in Geba, and the Philistines heard of it. And Saul blew the trumpet throughout all the land, saying, Let the Hebrews hear.
1SAM|13|4|And all Israel heard say that Saul had smitten a garrison of the Philistines, and that Israel also was had in abomination with the Philistines. And the people were called together after Saul to Gilgal.
1SAM|13|5|And the Philistines gathered themselves together to fight with Israel, thirty thousand chariots, and six thousand horsemen, and people as the sand which is on the sea shore in multitude: and they came up, and pitched in Michmash, eastward from Bethaven.
1SAM|13|6|When the men of Israel saw that they were in a strait, (for the people were distressed,) then the people did hide themselves in caves, and in thickets, and in rocks, and in high places, and in pits.
1SAM|13|7|And some of the Hebrews went over Jordan to the land of Gad and Gilead. As for Saul, he was yet in Gilgal, and all the people followed him trembling.
1SAM|13|8|And he tarried seven days, according to the set time that Samuel had appointed: but Samuel came not to Gilgal; and the people were scattered from him.
1SAM|13|9|And Saul said, Bring hither a burnt offering to me, and peace offerings. And he offered the burnt offering.
1SAM|13|10|And it came to pass, that as soon as he had made an end of offering the burnt offering, behold, Samuel came; and Saul went out to meet him, that he might salute him.
1SAM|13|11|And Samuel said, What hast thou done? And Saul said, Because I saw that the people were scattered from me, and that thou camest not within the days appointed, and that the Philistines gathered themselves together at Michmash;
1SAM|13|12|Therefore said I, The Philistines will come down now upon me to Gilgal, and I have not made supplication unto the LORD: I forced myself therefore, and offered a burnt offering.
1SAM|13|13|And Samuel said to Saul, Thou hast done foolishly: thou hast not kept the commandment of the LORD thy God, which he commanded thee: for now would the LORD have established thy kingdom upon Israel for ever.
1SAM|13|14|But now thy kingdom shall not continue: the LORD hath sought him a man after his own heart, and the LORD hath commanded him to be captain over his people, because thou hast not kept that which the LORD commanded thee.
1SAM|13|15|And Samuel arose, and gat him up from Gilgal unto Gibeah of Benjamin. And Saul numbered the people that were present with him, about six hundred men.
1SAM|13|16|And Saul, and Jonathan his son, and the people that were present with them, abode in Gibeah of Benjamin: but the Philistines encamped in Michmash.
1SAM|13|17|And the spoilers came out of the camp of the Philistines in three companies: one company turned unto the way that leadeth to Ophrah, unto the land of Shual:
1SAM|13|18|And another company turned the way to Bethhoron: and another company turned to the way of the border that looketh to the valley of Zeboim toward the wilderness.
1SAM|13|19|Now there was no smith found throughout all the land of Israel: for the Philistines said, Lest the Hebrews make them swords or spears:
1SAM|13|20|But all the Israelites went down to the Philistines, to sharpen every man his share, and his coulter, and his axe, and his mattock.
1SAM|13|21|Yet they had a file for the mattocks, and for the coulters, and for the forks, and for the axes, and to sharpen the goads.
1SAM|13|22|So it came to pass in the day of battle, that there was neither sword nor spear found in the hand of any of the people that were with Saul and Jonathan: but with Saul and with Jonathan his son was there found.
1SAM|13|23|And the garrison of the Philistines went out to the passage of Michmash.
1SAM|14|1|Now it came to pass upon a day, that Jonathan the son of Saul said unto the young man that bare his armor, Come, and let us go over to the Philistines' garrison, that is on the other side. But he told not his father.
1SAM|14|2|And Saul tarried in the uttermost part of Gibeah under a pomegranate tree which is in Migron: and the people that were with him were about six hundred men;
1SAM|14|3|And Ahiah, the son of Ahitub, Ichabod's brother, the son of Phinehas, the son of Eli, the LORD's priest in Shiloh, wearing an ephod. And the people knew not that Jonathan was gone.
1SAM|14|4|And between the passages, by which Jonathan sought to go over unto the Philistines' garrison, there was a sharp rock on the one side, and a sharp rock on the other side: and the name of the one was Bozez, and the name of the other Seneh.
1SAM|14|5|The forefront of the one was situate northward over against Michmash, and the other southward over against Gibeah.
1SAM|14|6|And Jonathan said to the young man that bare his armor, Come, and let us go over unto the garrison of these uncircumcised: it may be that the LORD will work for us: for there is no restraint to the LORD to save by many or by few.
1SAM|14|7|And his armourbearer said unto him, Do all that is in thine heart: turn thee; behold, I am with thee according to thy heart.
1SAM|14|8|Then said Jonathan, Behold, we will pass over unto these men, and we will discover ourselves unto them.
1SAM|14|9|If they say thus unto us, Tarry until we come to you; then we will stand still in our place, and will not go up unto them.
1SAM|14|10|But if they say thus, Come up unto us; then we will go up: for the LORD hath delivered them into our hand: and this shall be a sign unto us.
1SAM|14|11|And both of them discovered themselves unto the garrison of the Philistines: and the Philistines said, Behold, the Hebrews come forth out of the holes where they had hid themselves.
1SAM|14|12|And the men of the garrison answered Jonathan and his armourbearer, and said, Come up to us, and we will show you a thing. And Jonathan said unto his armourbearer, Come up after me: for the LORD hath delivered them into the hand of Israel.
1SAM|14|13|And Jonathan climbed up upon his hands and upon his feet, and his armourbearer after him: and they fell before Jonathan; and his armourbearer slew after him.
1SAM|14|14|And that first slaughter, which Jonathan and his armourbearer made, was about twenty men, within as it were an half acre of land, which a yoke of oxen might plow.
1SAM|14|15|And there was trembling in the host, in the field, and among all the people: the garrison, and the spoilers, they also trembled, and the earth quaked: so it was a very great trembling.
1SAM|14|16|And the watchmen of Saul in Gibeah of Benjamin looked; and, behold, the multitude melted away, and they went on beating down one another.
1SAM|14|17|Then said Saul unto the people that were with him, Number now, and see who is gone from us. And when they had numbered, behold, Jonathan and his armourbearer were not there.
1SAM|14|18|And Saul said unto Ahiah, Bring hither the ark of God. For the ark of God was at that time with the children of Israel.
1SAM|14|19|And it came to pass, while Saul talked unto the priest, that the noise that was in the host of the Philistines went on and increased: and Saul said unto the priest, Withdraw thine hand.
1SAM|14|20|And Saul and all the people that were with him assembled themselves, and they came to the battle: and, behold, every man's sword was against his fellow, and there was a very great discomfiture.
1SAM|14|21|Moreover the Hebrews that were with the Philistines before that time, which went up with them into the camp from the country round about, even they also turned to be with the Israelites that were with Saul and Jonathan.
1SAM|14|22|Likewise all the men of Israel which had hid themselves in mount Ephraim, when they heard that the Philistines fled, even they also followed hard after them in the battle.
1SAM|14|23|So the LORD saved Israel that day: and the battle passed over unto Bethaven.
1SAM|14|24|And the men of Israel were distressed that day: for Saul had adjured the people, saying, Cursed be the man that eateth any food until evening, that I may be avenged on mine enemies. So none of the people tasted any food.
1SAM|14|25|And all they of the land came to a wood; and there was honey upon the ground.
1SAM|14|26|And when the people were come into the wood, behold, the honey dropped; but no man put his hand to his mouth: for the people feared the oath.
1SAM|14|27|But Jonathan heard not when his father charged the people with the oath: wherefore he put forth the end of the rod that was in his hand, and dipped it in an honeycomb, and put his hand to his mouth; and his eyes were enlightened.
1SAM|14|28|Then answered one of the people, and said, Thy father straitly charged the people with an oath, saying, Cursed be the man that eateth any food this day. And the people were faint.
1SAM|14|29|Then said Jonathan, My father hath troubled the land: see, I pray you, how mine eyes have been enlightened, because I tasted a little of this honey.
1SAM|14|30|How much more, if haply the people had eaten freely to day of the spoil of their enemies which they found? for had there not been now a much greater slaughter among the Philistines?
1SAM|14|31|And they smote the Philistines that day from Michmash to Aijalon: and the people were very faint.
1SAM|14|32|And the people flew upon the spoil, and took sheep, and oxen, and calves, and slew them on the ground: and the people did eat them with the blood.
1SAM|14|33|Then they told Saul, saying, Behold, the people sin against the LORD, in that they eat with the blood. And he said, Ye have transgressed: roll a great stone unto me this day.
1SAM|14|34|And Saul said, Disperse yourselves among the people, and say unto them, Bring me hither every man his ox, and every man his sheep, and slay them here, and eat; and sin not against the LORD in eating with the blood. And all the people brought every man his ox with him that night, and slew them there.
1SAM|14|35|And Saul built an altar unto the LORD: the same was the first altar that he built unto the LORD.
1SAM|14|36|And Saul said, Let us go down after the Philistines by night, and spoil them until the morning light, and let us not leave a man of them. And they said, Do whatsoever seemeth good unto thee. Then said the priest, Let us draw near hither unto God.
1SAM|14|37|And Saul asked counsel of God, Shall I go down after the Philistines? wilt thou deliver them into the hand of Israel? But he answered him not that day.
1SAM|14|38|And Saul said, Draw ye near hither, all the chief of the people: and know and see wherein this sin hath been this day.
1SAM|14|39|For, as the LORD liveth, which saveth Israel, though it be in Jonathan my son, he shall surely die. But there was not a man among all the people that answered him.
1SAM|14|40|Then said he unto all Israel, Be ye on one side, and I and Jonathan my son will be on the other side. And the people said unto Saul, Do what seemeth good unto thee.
1SAM|14|41|Therefore Saul said unto the LORD God of Israel, Give a perfect lot. And Saul and Jonathan were taken: but the people escaped.
1SAM|14|42|And Saul said, Cast lots between me and Jonathan my son. And Jonathan was taken.
1SAM|14|43|Then Saul said to Jonathan, Tell me what thou hast done. And Jonathan told him, and said, I did but taste a little honey with the end of the rod that was in mine hand, and, lo, I must die.
1SAM|14|44|And Saul answered, God do so and more also: for thou shalt surely die, Jonathan.
1SAM|14|45|And the people said unto Saul, Shall Jonathan die, who hath wrought this great salvation in Israel? God forbid: as the LORD liveth, there shall not one hair of his head fall to the ground; for he hath wrought with God this day. So the people rescued Jonathan, that he died not.
1SAM|14|46|Then Saul went up from following the Philistines: and the Philistines went to their own place.
1SAM|14|47|So Saul took the kingdom over Israel, and fought against all his enemies on every side, against Moab, and against the children of Ammon, and against Edom, and against the kings of Zobah, and against the Philistines: and whithersoever he turned himself, he vexed them.
1SAM|14|48|And he gathered an host, and smote the Amalekites, and delivered Israel out of the hands of them that spoiled them.
1SAM|14|49|Now the sons of Saul were Jonathan, and Ishui, and Melchishua: and the names of his two daughters were these; the name of the firstborn Merab, and the name of the younger Michal:
1SAM|14|50|And the name of Saul's wife was Ahinoam, the daughter of Ahimaaz: and the name of the captain of his host was Abner, the son of Ner, Saul's uncle.
1SAM|14|51|And Kish was the father of Saul; and Ner the father of Abner was the son of Abiel.
1SAM|14|52|And there was sore war against the Philistines all the days of Saul: and when Saul saw any strong man, or any valiant man, he took him unto him.
1SAM|15|1|Samuel also said unto Saul, The LORD sent me to anoint thee to be king over his people, over Israel: now therefore hearken thou unto the voice of the words of the LORD.
1SAM|15|2|Thus saith the LORD of hosts, I remember that which Amalek did to Israel, how he laid wait for him in the way, when he came up from Egypt.
1SAM|15|3|Now go and smite Amalek, and utterly destroy all that they have, and spare them not; but slay both man and woman, infant and suckling, ox and sheep, camel and ass.
1SAM|15|4|And Saul gathered the people together, and numbered them in Telaim, two hundred thousand footmen, and ten thousand men of Judah.
1SAM|15|5|And Saul came to a city of Amalek, and laid wait in the valley.
1SAM|15|6|And Saul said unto the Kenites, Go, depart, get you down from among the Amalekites, lest I destroy you with them: for ye showed kindness to all the children of Israel, when they came up out of Egypt. So the Kenites departed from among the Amalekites.
1SAM|15|7|And Saul smote the Amalekites from Havilah until thou comest to Shur, that is over against Egypt.
1SAM|15|8|And he took Agag the king of the Amalekites alive, and utterly destroyed all the people with the edge of the sword.
1SAM|15|9|But Saul and the people spared Agag, and the best of the sheep, and of the oxen, and of the fatlings, and the lambs, and all that was good, and would not utterly destroy them: but every thing that was vile and refuse, that they destroyed utterly.
1SAM|15|10|Then came the word of the LORD unto Samuel, saying,
1SAM|15|11|It repenteth me that I have set up Saul to be king: for he is turned back from following me, and hath not performed my commandments. And it grieved Samuel; and he cried unto the LORD all night.
1SAM|15|12|And when Samuel rose early to meet Saul in the morning, it was told Samuel, saying, Saul came to Carmel, and, behold, he set him up a place, and is gone about, and passed on, and gone down to Gilgal.
1SAM|15|13|And Samuel came to Saul: and Saul said unto him, Blessed be thou of the LORD: I have performed the commandment of the LORD.
1SAM|15|14|And Samuel said, What meaneth then this bleating of the sheep in mine ears, and the lowing of the oxen which I hear?
1SAM|15|15|And Saul said, They have brought them from the Amalekites: for the people spared the best of the sheep and of the oxen, to sacrifice unto the LORD thy God; and the rest we have utterly destroyed.
1SAM|15|16|Then Samuel said unto Saul, Stay, and I will tell thee what the LORD hath said to me this night. And he said unto him, Say on.
1SAM|15|17|And Samuel said, When thou wast little in thine own sight, wast thou not made the head of the tribes of Israel, and the LORD anointed thee king over Israel?
1SAM|15|18|And the LORD sent thee on a journey, and said, Go and utterly destroy the sinners the Amalekites, and fight against them until they be consumed.
1SAM|15|19|Wherefore then didst thou not obey the voice of the LORD, but didst fly upon the spoil, and didst evil in the sight of the LORD?
1SAM|15|20|And Saul said unto Samuel, Yea, I have obeyed the voice of the LORD, and have gone the way which the LORD sent me, and have brought Agag the king of Amalek, and have utterly destroyed the Amalekites.
1SAM|15|21|But the people took of the spoil, sheep and oxen, the chief of the things which should have been utterly destroyed, to sacrifice unto the LORD thy God in Gilgal.
1SAM|15|22|And Samuel said, Hath the LORD as great delight in burnt offerings and sacrifices, as in obeying the voice of the LORD? Behold, to obey is better than sacrifice, and to hearken than the fat of rams.
1SAM|15|23|For rebellion is as the sin of witchcraft, and stubbornness is as iniquity and idolatry. Because thou hast rejected the word of the LORD, he hath also rejected thee from being king.
1SAM|15|24|And Saul said unto Samuel, I have sinned: for I have transgressed the commandment of the LORD, and thy words: because I feared the people, and obeyed their voice.
1SAM|15|25|Now therefore, I pray thee, pardon my sin, and turn again with me, that I may worship the LORD.
1SAM|15|26|And Samuel said unto Saul, I will not return with thee: for thou hast rejected the word of the LORD, and the LORD hath rejected thee from being king over Israel.
1SAM|15|27|And as Samuel turned about to go away, he laid hold upon the skirt of his mantle, and it rent.
1SAM|15|28|And Samuel said unto him, The LORD hath rent the kingdom of Israel from thee this day, and hath given it to a neighbor of thine, that is better than thou.
1SAM|15|29|And also the Strength of Israel will not lie nor repent: for he is not a man, that he should repent.
1SAM|15|30|Then he said, I have sinned: yet honor me now, I pray thee, before the elders of my people, and before Israel, and turn again with me, that I may worship the LORD thy God.
1SAM|15|31|So Samuel turned again after Saul; and Saul worshipped the LORD.
1SAM|15|32|Then said Samuel, Bring ye hither to me Agag the king of the Amalekites. And Agag came unto him delicately. And Agag said, Surely the bitterness of death is past.
1SAM|15|33|And Samuel said, As the sword hath made women childless, so shall thy mother be childless among women. And Samuel hewed Agag in pieces before the LORD in Gilgal.
1SAM|15|34|Then Samuel went to Ramah; and Saul went up to his house to Gibeah of Saul.
1SAM|15|35|And Samuel came no more to see Saul until the day of his death: nevertheless Samuel mourned for Saul: and the LORD repented that he had made Saul king over Israel.
1SAM|16|1|And the LORD said unto Samuel, How long wilt thou mourn for Saul, seeing I have rejected him from reigning over Israel? fill thine horn with oil, and go, I will send thee to Jesse the Bethlehemite: for I have provided me a king among his sons.
1SAM|16|2|And Samuel said, How can I go? if Saul hear it, he will kill me. And the LORD said, Take an heifer with thee, and say, I am come to sacrifice to the LORD.
1SAM|16|3|And call Jesse to the sacrifice, and I will show thee what thou shalt do: and thou shalt anoint unto me him whom I name unto thee.
1SAM|16|4|And Samuel did that which the LORD spake, and came to Bethlehem. And the elders of the town trembled at his coming, and said, Comest thou peaceably?
1SAM|16|5|And he said, Peaceably: I am come to sacrifice unto the LORD: sanctify yourselves, and come with me to the sacrifice. And he sanctified Jesse and his sons, and called them to the sacrifice.
1SAM|16|6|And it came to pass, when they were come, that he looked on Eliab, and said, Surely the LORD's anointed is before him.
1SAM|16|7|But the LORD said unto Samuel, Look not on his countenance, or on the height of his stature; because I have refused him: for the LORD seeth not as man seeth; for man looketh on the outward appearance, but the LORD looketh on the heart.
1SAM|16|8|Then Jesse called Abinadab, and made him pass before Samuel. And he said, Neither hath the LORD chosen this.
1SAM|16|9|Then Jesse made Shammah to pass by. And he said, Neither hath the LORD chosen this.
1SAM|16|10|Again, Jesse made seven of his sons to pass before Samuel. And Samuel said unto Jesse, The LORD hath not chosen these.
1SAM|16|11|And Samuel said unto Jesse, Are here all thy children? And he said, There remaineth yet the youngest, and, behold, he keepeth the sheep. And Samuel said unto Jesse, Send and fetch him: for we will not sit down till he come hither.
1SAM|16|12|And he sent, and brought him in. Now he was ruddy, and withal of a beautiful countenance, and goodly to look to. And the LORD said, Arise, anoint him: for this is he.
1SAM|16|13|Then Samuel took the horn of oil, and anointed him in the midst of his brethren: and the Spirit of the LORD came upon David from that day forward. So Samuel rose up, and went to Ramah.
1SAM|16|14|But the Spirit of the LORD departed from Saul, and an evil spirit from the LORD troubled him.
1SAM|16|15|And Saul's servants said unto him, Behold now, an evil spirit from God troubleth thee.
1SAM|16|16|Let our lord now command thy servants, which are before thee, to seek out a man, who is a cunning player on an harp: and it shall come to pass, when the evil spirit from God is upon thee, that he shall play with his hand, and thou shalt be well.
1SAM|16|17|And Saul said unto his servants, Provide me now a man that can play well, and bring him to me.
1SAM|16|18|Then answered one of the servants, and said, Behold, I have seen a son of Jesse the Bethlehemite, that is cunning in playing, and a mighty valiant man, and a man of war, and prudent in matters, and a comely person, and the LORD is with him.
1SAM|16|19|Wherefore Saul sent messengers unto Jesse, and said, Send me David thy son, which is with the sheep.
1SAM|16|20|And Jesse took an ass laden with bread, and a bottle of wine, and a kid, and sent them by David his son unto Saul.
1SAM|16|21|And David came to Saul, and stood before him: and he loved him greatly; and he became his armourbearer.
1SAM|16|22|And Saul sent to Jesse, saying, Let David, I pray thee, stand before me; for he hath found favor in my sight.
1SAM|16|23|And it came to pass, when the evil spirit from God was upon Saul, that David took an harp, and played with his hand: so Saul was refreshed, and was well, and the evil spirit departed from him.
1SAM|17|1|Now the Philistines gathered together their armies to battle, and were gathered together at Shochoh, which belongeth to Judah, and pitched between Shochoh and Azekah, in Ephesdammim.
1SAM|17|2|And Saul and the men of Israel were gathered together, and pitched by the valley of Elah, and set the battle in array against the Philistines.
1SAM|17|3|And the Philistines stood on a mountain on the one side, and Israel stood on a mountain on the other side: and there was a valley between them.
1SAM|17|4|And there went out a champion out of the camp of the Philistines, named Goliath, of Gath, whose height was six cubits and a span.
1SAM|17|5|And he had an helmet of brass upon his head, and he was armed with a coat of mail; and the weight of the coat was five thousand shekels of brass.
1SAM|17|6|And he had greaves of brass upon his legs, and a target of brass between his shoulders.
1SAM|17|7|And the staff of his spear was like a weaver's beam; and his spear's head weighed six hundred shekels of iron: and one bearing a shield went before him.
1SAM|17|8|And he stood and cried unto the armies of Israel, and said unto them, Why are ye come out to set your battle in array? am not I a Philistine, and ye servants to Saul? choose you a man for you, and let him come down to me.
1SAM|17|9|If he be able to fight with me, and to kill me, then will we be your servants: but if I prevail against him, and kill him, then shall ye be our servants, and serve us.
1SAM|17|10|And the Philistine said, I defy the armies of Israel this day; give me a man, that we may fight together.
1SAM|17|11|When Saul and all Israel heard those words of the Philistine, they were dismayed, and greatly afraid.
1SAM|17|12|Now David was the son of that Ephrathite of Bethlehemjudah, whose name was Jesse; and he had eight sons: and the man went among men for an old man in the days of Saul.
1SAM|17|13|And the three eldest sons of Jesse went and followed Saul to the battle: and the names of his three sons that went to the battle were Eliab the firstborn, and next unto him Abinadab, and the third Shammah.
1SAM|17|14|And David was the youngest: and the three eldest followed Saul.
1SAM|17|15|But David went and returned from Saul to feed his father's sheep at Bethlehem.
1SAM|17|16|And the Philistine drew near morning and evening, and presented himself forty days.
1SAM|17|17|And Jesse said unto David his son, Take now for thy brethren an ephah of this parched corn, and these ten loaves, and run to the camp of thy brethren;
1SAM|17|18|And carry these ten cheeses unto the captain of their thousand, and look how thy brethren fare, and take their pledge.
1SAM|17|19|Now Saul, and they, and all the men of Israel, were in the valley of Elah, fighting with the Philistines.
1SAM|17|20|And David rose up early in the morning, and left the sheep with a keeper, and took, and went, as Jesse had commanded him; and he came to the trench, as the host was going forth to the fight, and shouted for the battle.
1SAM|17|21|For Israel and the Philistines had put the battle in array, army against army.
1SAM|17|22|And David left his carriage in the hand of the keeper of the carriage, and ran into the army, and came and saluted his brethren.
1SAM|17|23|And as he talked with them, behold, there came up the champion, the Philistine of Gath, Goliath by name, out of the armies of the Philistines, and spake according to the same words: and David heard them.
1SAM|17|24|And all the men of Israel, when they saw the man, fled from him, and were sore afraid.
1SAM|17|25|And the men of Israel said, Have ye seen this man that is come up? surely to defy Israel is he come up: and it shall be, that the man who killeth him, the king will enrich him with great riches, and will give him his daughter, and make his father's house free in Israel.
1SAM|17|26|And David spake to the men that stood by him, saying, What shall be done to the man that killeth this Philistine, and taketh away the reproach from Israel? for who is this uncircumcised Philistine, that he should defy the armies of the living God?
1SAM|17|27|And the people answered him after this manner, saying, So shall it be done to the man that killeth him.
1SAM|17|28|And Eliab his eldest brother heard when he spake unto the men; and Eliab's anger was kindled against David, and he said, Why camest thou down hither? and with whom hast thou left those few sheep in the wilderness? I know thy pride, and the naughtiness of thine heart; for thou art come down that thou mightest see the battle.
1SAM|17|29|And David said, What have I now done? Is there not a cause?
1SAM|17|30|And he turned from him toward another, and spake after the same manner: and the people answered him again after the former manner.
1SAM|17|31|And when the words were heard which David spake, they rehearsed them before Saul: and he sent for him.
1SAM|17|32|And David said to Saul, Let no man's heart fail because of him; thy servant will go and fight with this Philistine.
1SAM|17|33|And Saul said to David, Thou art not able to go against this Philistine to fight with him: for thou art but a youth, and he a man of war from his youth.
1SAM|17|34|And David said unto Saul, Thy servant kept his father's sheep, and there came a lion, and a bear, and took a lamb out of the flock:
1SAM|17|35|And I went out after him, and smote him, and delivered it out of his mouth: and when he arose against me, I caught him by his beard, and smote him, and slew him.
1SAM|17|36|Thy servant slew both the lion and the bear: and this uncircumcised Philistine shall be as one of them, seeing he hath defied the armies of the living God.
1SAM|17|37|David said moreover, The LORD that delivered me out of the paw of the lion, and out of the paw of the bear, he will deliver me out of the hand of this Philistine. And Saul said unto David, Go, and the LORD be with thee.
1SAM|17|38|And Saul armed David with his armor, and he put an helmet of brass upon his head; also he armed him with a coat of mail.
1SAM|17|39|And David girded his sword upon his armor, and he assayed to go; for he had not proved it. And David said unto Saul, I cannot go with these; for I have not proved them. And David put them off him.
1SAM|17|40|And he took his staff in his hand, and chose him five smooth stones out of the brook, and put them in a shepherd's bag which he had, even in a scrip; and his sling was in his hand: and he drew near to the Philistine.
1SAM|17|41|And the Philistine came on and drew near unto David; and the man that bare the shield went before him.
1SAM|17|42|And when the Philistine looked about, and saw David, he disdained him: for he was but a youth, and ruddy, and of a fair countenance.
1SAM|17|43|And the Philistine said unto David, Am I a dog, that thou comest to me with staves? And the Philistine cursed David by his gods.
1SAM|17|44|And the Philistine said to David, Come to me, and I will give thy flesh unto the fowls of the air, and to the beasts of the field.
1SAM|17|45|Then said David to the Philistine, Thou comest to me with a sword, and with a spear, and with a shield: but I come to thee in the name of the LORD of hosts, the God of the armies of Israel, whom thou hast defied.
1SAM|17|46|This day will the LORD deliver thee into mine hand; and I will smite thee, and take thine head from thee; and I will give the carcasses of the host of the Philistines this day unto the fowls of the air, and to the wild beasts of the earth; that all the earth may know that there is a God in Israel.
1SAM|17|47|And all this assembly shall know that the LORD saveth not with sword and spear: for the battle is the LORD's, and he will give you into our hands.
1SAM|17|48|And it came to pass, when the Philistine arose, and came, and drew nigh to meet David, that David hastened, and ran toward the army to meet the Philistine.
1SAM|17|49|And David put his hand in his bag, and took thence a stone, and slang it, and smote the Philistine in his forehead, that the stone sunk into his forehead; and he fell upon his face to the earth.
1SAM|17|50|So David prevailed over the Philistine with a sling and with a stone, and smote the Philistine, and slew him; but there was no sword in the hand of David.
1SAM|17|51|Therefore David ran, and stood upon the Philistine, and took his sword, and drew it out of the sheath thereof, and slew him, and cut off his head therewith. And when the Philistines saw their champion was dead, they fled.
1SAM|17|52|And the men of Israel and of Judah arose, and shouted, and pursued the Philistines, until thou come to the valley, and to the gates of Ekron. And the wounded of the Philistines fell down by the way to Shaaraim, even unto Gath, and unto Ekron.
1SAM|17|53|And the children of Israel returned from chasing after the Philistines, and they spoiled their tents.
1SAM|17|54|And David took the head of the Philistine, and brought it to Jerusalem; but he put his armor in his tent.
1SAM|17|55|And when Saul saw David go forth against the Philistine, he said unto Abner, the captain of the host, Abner, whose son is this youth? And Abner said, As thy soul liveth, O king, I cannot tell.
1SAM|17|56|And the king said, Inquire thou whose son the stripling is.
1SAM|17|57|And as David returned from the slaughter of the Philistine, Abner took him, and brought him before Saul with the head of the Philistine in his hand.
1SAM|17|58|And Saul said to him, Whose son art thou, thou young man? And David answered, I am the son of thy servant Jesse the Bethlehemite.
1SAM|18|1|And it came to pass, when he had made an end of speaking unto Saul, that the soul of Jonathan was knit with the soul of David, and Jonathan loved him as his own soul.
1SAM|18|2|And Saul took him that day, and would let him go no more home to his father's house.
1SAM|18|3|Then Jonathan and David made a covenant, because he loved him as his own soul.
1SAM|18|4|And Jonathan stripped himself of the robe that was upon him, and gave it to David, and his garments, even to his sword, and to his bow, and to his girdle.
1SAM|18|5|And David went out whithersoever Saul sent him, and behaved himself wisely: and Saul set him over the men of war, and he was accepted in the sight of all the people, and also in the sight of Saul's servants.
1SAM|18|6|And it came to pass as they came, when David was returned from the slaughter of the Philistine, that the women came out of all cities of Israel, singing and dancing, to meet king Saul, with tabrets, with joy, and with instruments of music.
1SAM|18|7|And the women answered one another as they played, and said, Saul hath slain his thousands, and David his ten thousands.
1SAM|18|8|And Saul was very wroth, and the saying displeased him; and he said, They have ascribed unto David ten thousands, and to me they have ascribed but thousands: and what can he have more but the kingdom?
1SAM|18|9|And Saul eyed David from that day and forward.
1SAM|18|10|And it came to pass on the morrow, that the evil spirit from God came upon Saul, and he prophesied in the midst of the house: and David played with his hand, as at other times: and there was a javelin in Saul's hand.
1SAM|18|11|And Saul cast the javelin; for he said, I will smite David even to the wall with it. And David avoided out of his presence twice.
1SAM|18|12|And Saul was afraid of David, because the LORD was with him, and was departed from Saul.
1SAM|18|13|Therefore Saul removed him from him, and made him his captain over a thousand; and he went out and came in before the people.
1SAM|18|14|And David behaved himself wisely in all his ways; and the LORD was with him.
1SAM|18|15|Wherefore when Saul saw that he behaved himself very wisely, he was afraid of him.
1SAM|18|16|But all Israel and Judah loved David, because he went out and came in before them.
1SAM|18|17|And Saul said to David, Behold my elder daughter Merab, her will I give thee to wife: only be thou valiant for me, and fight the LORD's battles. For Saul said, Let not mine hand be upon him, but let the hand of the Philistines be upon him.
1SAM|18|18|And David said unto Saul, Who am I? and what is my life, or my father's family in Israel, that I should be son in law to the king?
1SAM|18|19|But it came to pass at the time when Merab Saul's daughter should have been given to David, that she was given unto Adriel the Meholathite to wife.
1SAM|18|20|And Michal Saul's daughter loved David: and they told Saul, and the thing pleased him.
1SAM|18|21|And Saul said, I will give him her, that she may be a snare to him, and that the hand of the Philistines may be against him. Wherefore Saul said to David, Thou shalt this day be my son in law in the one of the twain.
1SAM|18|22|And Saul commanded his servants, saying, Commune with David secretly, and say, Behold, the king hath delight in thee, and all his servants love thee: now therefore be the king's son in law.
1SAM|18|23|And Saul's servants spake those words in the ears of David. And David said, Seemeth it to you a light thing to be a king's son in law, seeing that I am a poor man, and lightly esteemed?
1SAM|18|24|And the servants of Saul told him, saying, On this manner spake David.
1SAM|18|25|And Saul said, Thus shall ye say to David, The king desireth not any dowry, but an hundred foreskins of the Philistines, to be avenged of the king's enemies. But Saul thought to make David fall by the hand of the Philistines.
1SAM|18|26|And when his servants told David these words, it pleased David well to be the king's son in law: and the days were not expired.
1SAM|18|27|Wherefore David arose and went, he and his men, and slew of the Philistines two hundred men; and David brought their foreskins, and they gave them in full tale to the king, that he might be the king's son in law. And Saul gave him Michal his daughter to wife.
1SAM|18|28|And Saul saw and knew that the LORD was with David, and that Michal Saul's daughter loved him.
1SAM|18|29|And Saul was yet the more afraid of David; and Saul became David's enemy continually.
1SAM|18|30|Then the princes of the Philistines went forth: and it came to pass, after they went forth, that David behaved himself more wisely than all the servants of Saul; so that his name was much set by.
1SAM|19|1|And Saul spake to Jonathan his son, and to all his servants, that they should kill David.
1SAM|19|2|But Jonathan Saul's son delighted much in David: and Jonathan told David, saying, Saul my father seeketh to kill thee: now therefore, I pray thee, take heed to thyself until the morning, and abide in a secret place, and hide thyself:
1SAM|19|3|And I will go out and stand beside my father in the field where thou art, and I will commune with my father of thee; and what I see, that I will tell thee.
1SAM|19|4|And Jonathan spake good of David unto Saul his father, and said unto him, Let not the king sin against his servant, against David; because he hath not sinned against thee, and because his works have been to thee-ward very good:
1SAM|19|5|For he did put his life in his hand, and slew the Philistine, and the LORD wrought a great salvation for all Israel: thou sawest it, and didst rejoice: wherefore then wilt thou sin against innocent blood, to slay David without a cause?
1SAM|19|6|And Saul hearkened unto the voice of Jonathan: and Saul sware, As the LORD liveth, he shall not be slain.
1SAM|19|7|And Jonathan called David, and Jonathan showed him all those things. And Jonathan brought David to Saul, and he was in his presence, as in times past.
1SAM|19|8|And there was war again: and David went out, and fought with the Philistines, and slew them with a great slaughter; and they fled from him.
1SAM|19|9|And the evil spirit from the LORD was upon Saul, as he sat in his house with his javelin in his hand: and David played with his hand.
1SAM|19|10|And Saul sought to smite David even to the wall with the javelin: but he slipped away out of Saul's presence, and he smote the javelin into the wall: and David fled, and escaped that night.
1SAM|19|11|Saul also sent messengers unto David's house, to watch him, and to slay him in the morning: and Michal David's wife told him, saying, If thou save not thy life to night, to morrow thou shalt be slain.
1SAM|19|12|So Michal let David down through a window: and he went, and fled, and escaped.
1SAM|19|13|And Michal took an image, and laid it in the bed, and put a pillow of goats' hair for his bolster, and covered it with a cloth.
1SAM|19|14|And when Saul sent messengers to take David, she said, He is sick.
1SAM|19|15|And Saul sent the messengers again to see David, saying, Bring him up to me in the bed, that I may slay him.
1SAM|19|16|And when the messengers were come in, behold, there was an image in the bed, with a pillow of goats' hair for his bolster.
1SAM|19|17|And Saul said unto Michal, Why hast thou deceived me so, and sent away mine enemy, that he is escaped? And Michal answered Saul, He said unto me, Let me go; why should I kill thee?
1SAM|19|18|So David fled, and escaped, and came to Samuel to Ramah, and told him all that Saul had done to him. And he and Samuel went and dwelt in Naioth.
1SAM|19|19|And it was told Saul, saying, Behold, David is at Naioth in Ramah.
1SAM|19|20|And Saul sent messengers to take David: and when they saw the company of the prophets prophesying, and Samuel standing as appointed over them, the Spirit of God was upon the messengers of Saul, and they also prophesied.
1SAM|19|21|And when it was told Saul, he sent other messengers, and they prophesied likewise. And Saul sent messengers again the third time, and they prophesied also.
1SAM|19|22|Then went he also to Ramah, and came to a great well that is in Sechu: and he asked and said, Where are Samuel and David? And one said, Behold, they be at Naioth in Ramah.
1SAM|19|23|And he went thither to Naioth in Ramah: and the Spirit of God was upon him also, and he went on, and prophesied, until he came to Naioth in Ramah.
1SAM|19|24|And he stripped off his clothes also, and prophesied before Samuel in like manner, and lay down naked all that day and all that night. Wherefore they say, Is Saul also among the prophets?
1SAM|20|1|And David fled from Naioth in Ramah, and came and said before Jonathan, What have I done? what is mine iniquity? and what is my sin before thy father, that he seeketh my life?
1SAM|20|2|And he said unto him, God forbid; thou shalt not die: behold, my father will do nothing either great or small, but that he will show it me: and why should my father hide this thing from me? it is not so.
1SAM|20|3|And David sware moreover, and said, Thy father certainly knoweth that I have found grace in thine eyes; and he saith, Let not Jonathan know this, lest he be grieved: but truly as the LORD liveth, and as thy soul liveth, there is but a step between me and death.
1SAM|20|4|Then said Jonathan unto David, Whatsoever thy soul desireth, I will even do it for thee.
1SAM|20|5|And David said unto Jonathan, Behold, to morrow is the new moon, and I should not fail to sit with the king at meat: but let me go, that I may hide myself in the field unto the third day at even.
1SAM|20|6|If thy father at all miss me, then say, David earnestly asked leave of me that he might run to Bethlehem his city: for there is a yearly sacrifice there for all the family.
1SAM|20|7|If he say thus, It is well; thy servant shall have peace: but if he be very wroth, then be sure that evil is determined by him.
1SAM|20|8|Therefore thou shalt deal kindly with thy servant; for thou hast brought thy servant into a covenant of the LORD with thee: notwithstanding, if there be in me iniquity, slay me thyself; for why shouldest thou bring me to thy father?
1SAM|20|9|And Jonathan said, Far be it from thee: for if I knew certainly that evil were determined by my father to come upon thee, then would not I tell it thee?
1SAM|20|10|Then said David to Jonathan, Who shall tell me? or what if thy father answer thee roughly?
1SAM|20|11|And Jonathan said unto David, Come, and let us go out into the field. And they went out both of them into the field.
1SAM|20|12|And Jonathan said unto David, O LORD God of Israel, when I have sounded my father about to morrow any time, or the third day, and, behold, if there be good toward David, and I then send not unto thee, and show it thee;
1SAM|20|13|The LORD do so and much more to Jonathan: but if it please my father to do thee evil, then I will show it thee, and send thee away, that thou mayest go in peace: and the LORD be with thee, as he hath been with my father.
1SAM|20|14|And thou shalt not only while yet I live show me the kindness of the LORD, that I die not:
1SAM|20|15|But also thou shalt not cut off thy kindness from my house for ever: no, not when the LORD hath cut off the enemies of David every one from the face of the earth.
1SAM|20|16|So Jonathan made a covenant with the house of David, saying, Let the LORD even require it at the hand of David's enemies.
1SAM|20|17|And Jonathan caused David to swear again, because he loved him: for he loved him as he loved his own soul.
1SAM|20|18|Then Jonathan said to David, To morrow is the new moon: and thou shalt be missed, because thy seat will be empty.
1SAM|20|19|And when thou hast stayed three days, then thou shalt go down quickly, and come to the place where thou didst hide thyself when the business was in hand, and shalt remain by the stone Ezel.
1SAM|20|20|And I will shoot three arrows on the side thereof, as though I shot at a mark.
1SAM|20|21|And, behold, I will send a lad, saying, Go, find out the arrows. If I expressly say unto the lad, Behold, the arrows are on this side of thee, take them; then come thou: for there is peace to thee, and no hurt; as the LORD liveth.
1SAM|20|22|But if I say thus unto the young man, Behold, the arrows are beyond thee; go thy way: for the LORD hath sent thee away.
1SAM|20|23|And as touching the matter which thou and I have spoken of, behold, the LORD be between thee and me for ever.
1SAM|20|24|So David hid himself in the field: and when the new moon was come, the king sat him down to eat meat.
1SAM|20|25|And the king sat upon his seat, as at other times, even upon a seat by the wall: and Jonathan arose, and Abner sat by Saul's side, and David's place was empty.
1SAM|20|26|Nevertheless Saul spake not any thing that day: for he thought, Something hath befallen him, he is not clean; surely he is not clean.
1SAM|20|27|And it came to pass on the morrow, which was the second day of the month, that David's place was empty: and Saul said unto Jonathan his son, Wherefore cometh not the son of Jesse to meat, neither yesterday, nor to day?
1SAM|20|28|And Jonathan answered Saul, David earnestly asked leave of me to go to Bethlehem:
1SAM|20|29|And he said, Let me go, I pray thee; for our family hath a sacrifice in the city; and my brother, he hath commanded me to be there: and now, if I have found favor in thine eyes, let me get away, I pray thee, and see my brethren. Therefore he cometh not unto the king's table.
1SAM|20|30|Then Saul's anger was kindled against Jonathan, and he said unto him, Thou son of the perverse rebellious woman, do not I know that thou hast chosen the son of Jesse to thine own confusion, and unto the confusion of thy mother's nakedness?
1SAM|20|31|For as long as the son of Jesse liveth upon the ground, thou shalt not be established, nor thy kingdom. Wherefore now send and fetch him unto me, for he shall surely die.
1SAM|20|32|And Jonathan answered Saul his father, and said unto him, Wherefore shall he be slain? what hath he done?
1SAM|20|33|And Saul cast a javelin at him to smite him: whereby Jonathan knew that it was determined of his father to slay David.
1SAM|20|34|So Jonathan arose from the table in fierce anger, and did eat no meat the second day of the month: for he was grieved for David, because his father had done him shame.
1SAM|20|35|And it came to pass in the morning, that Jonathan went out into the field at the time appointed with David, and a little lad with him.
1SAM|20|36|And he said unto his lad, Run, find out now the arrows which I shoot. And as the lad ran, he shot an arrow beyond him.
1SAM|20|37|And when the lad was come to the place of the arrow which Jonathan had shot, Jonathan cried after the lad, and said, Is not the arrow beyond thee?
1SAM|20|38|And Jonathan cried after the lad, Make speed, haste, stay not. And Jonathan's lad gathered up the arrows, and came to his master.
1SAM|20|39|But the lad knew not any thing: only Jonathan and David knew the matter.
1SAM|20|40|And Jonathan gave his artillery unto his lad, and said unto him, Go, carry them to the city.
1SAM|20|41|And as soon as the lad was gone, David arose out of a place toward the south, and fell on his face to the ground, and bowed himself three times: and they kissed one another, and wept one with another, until David exceeded.
1SAM|20|42|And Jonathan said to David, Go in peace, forasmuch as we have sworn both of us in the name of the LORD, saying, The LORD be between me and thee, and between my seed and thy seed for ever. And he arose and departed: and Jonathan went into the city.
1SAM|21|1|Then came David to Nob to Ahimelech the priest: and Ahimelech was afraid at the meeting of David, and said unto him, Why art thou alone, and no man with thee?
1SAM|21|2|And David said unto Ahimelech the priest, The king hath commanded me a business, and hath said unto me, Let no man know any thing of the business whereabout I send thee, and what I have commanded thee: and I have appointed my servants to such and such a place.
1SAM|21|3|Now therefore what is under thine hand? give me five loaves of bread in mine hand, or what there is present.
1SAM|21|4|And the priest answered David, and said, There is no common bread under mine hand, but there is hallowed bread; if the young men have kept themselves at least from women.
1SAM|21|5|And David answered the priest, and said unto him, Of a truth women have been kept from us about these three days, since I came out, and the vessels of the young men are holy, and the bread is in a manner common, yea, though it were sanctified this day in the vessel.
1SAM|21|6|So the priest gave him hallowed bread: for there was no bread there but the showbread, that was taken from before the LORD, to put hot bread in the day when it was taken away.
1SAM|21|7|Now a certain man of the servants of Saul was there that day, detained before the LORD; and his name was Doeg, an Edomite, the chiefest of the herdmen that belonged to Saul.
1SAM|21|8|And David said unto Ahimelech, And is there not here under thine hand spear or sword? for I have neither brought my sword nor my weapons with me, because the king's business required haste.
1SAM|21|9|And the priest said, The sword of Goliath the Philistine, whom thou slewest in the valley of Elah, behold, it is here wrapped in a cloth behind the ephod: if thou wilt take that, take it: for there is no other save that here. And David said, There is none like that; give it me.
1SAM|21|10|And David arose and fled that day for fear of Saul, and went to Achish the king of Gath.
1SAM|21|11|And the servants of Achish said unto him, Is not this David the king of the land? did they not sing one to another of him in dances, saying, Saul hath slain his thousands, and David his ten thousands?
1SAM|21|12|And David laid up these words in his heart, and was sore afraid of Achish the king of Gath.
1SAM|21|13|And he changed his behavior before them, and feigned himself mad in their hands, and scrabbled on the doors of the gate, and let his spittle fall down upon his beard.
1SAM|21|14|Then said Achish unto his servants, Lo, ye see the man is mad: wherefore then have ye brought him to me?
1SAM|21|15|Have I need of mad men, that ye have brought this fellow to play the mad man in my presence? shall this fellow come into my house?
1SAM|22|1|David therefore departed thence, and escaped to the cave Adullam: and when his brethren and all his father's house heard it, they went down thither to him.
1SAM|22|2|And every one that was in distress, and every one that was in debt, and every one that was discontented, gathered themselves unto him; and he became a captain over them: and there were with him about four hundred men.
1SAM|22|3|And David went thence to Mizpeh of Moab: and he said unto the king of Moab, Let my father and my mother, I pray thee, come forth, and be with you, till I know what God will do for me.
1SAM|22|4|And he brought them before the king of Moab: and they dwelt with him all the while that David was in the hold.
1SAM|22|5|And the prophet Gad said unto David, Abide not in the hold; depart, and get thee into the land of Judah. Then David departed, and came into the forest of Hareth.
1SAM|22|6|When Saul heard that David was discovered, and the men that were with him, (now Saul abode in Gibeah under a tree in Ramah, having his spear in his hand, and all his servants were standing about him;)
1SAM|22|7|Then Saul said unto his servants that stood about him, Hear now, ye Benjamites; will the son of Jesse give every one of you fields and vineyards, and make you all captains of thousands, and captains of hundreds;
1SAM|22|8|That all of you have conspired against me, and there is none that showeth me that my son hath made a league with the son of Jesse, and there is none of you that is sorry for me, or showeth unto me that my son hath stirred up my servant against me, to lie in wait, as at this day?
1SAM|22|9|Then answered Doeg the Edomite, which was set over the servants of Saul, and said, I saw the son of Jesse coming to Nob, to Ahimelech the son of Ahitub.
1SAM|22|10|And he inquired of the LORD for him, and gave him victuals, and gave him the sword of Goliath the Philistine.
1SAM|22|11|Then the king sent to call Ahimelech the priest, the son of Ahitub, and all his father's house, the priests that were in Nob: and they came all of them to the king.
1SAM|22|12|And Saul said, Hear now, thou son of Ahitub. And he answered, Here I am, my lord.
1SAM|22|13|And Saul said unto him, Why have ye conspired against me, thou and the son of Jesse, in that thou hast given him bread, and a sword, and hast inquired of God for him, that he should rise against me, to lie in wait, as at this day?
1SAM|22|14|Then Ahimelech answered the king, and said, And who is so faithful among all thy servants as David, which is the king's son in law, and goeth at thy bidding, and is honorable in thine house?
1SAM|22|15|Did I then begin to inquire of God for him? be it far from me: let not the king impute any thing unto his servant, nor to all the house of my father: for thy servant knew nothing of all this, less or more.
1SAM|22|16|And the king said, Thou shalt surely die, Ahimelech, thou, and all thy father's house.
1SAM|22|17|And the king said unto the footmen that stood about him, Turn, and slay the priests of the LORD: because their hand also is with David, and because they knew when he fled, and did not show it to me. But the servants of the king would not put forth their hand to fall upon the priests of the LORD.
1SAM|22|18|And the king said to Doeg, Turn thou, and fall upon the priests. And Doeg the Edomite turned, and he fell upon the priests, and slew on that day fourscore and five persons that did wear a linen ephod.
1SAM|22|19|And Nob, the city of the priests, smote he with the edge of the sword, both men and women, children and sucklings, and oxen, and asses, and sheep, with the edge of the sword.
1SAM|22|20|And one of the sons of Ahimelech the son of Ahitub, named Abiathar, escaped, and fled after David.
1SAM|22|21|And Abiathar showed David that Saul had slain the LORD's priests.
1SAM|22|22|And David said unto Abiathar, I knew it that day, when Doeg the Edomite was there, that he would surely tell Saul: I have occasioned the death of all the persons of thy father's house.
1SAM|22|23|Abide thou with me, fear not: for he that seeketh my life seeketh thy life: but with me thou shalt be in safeguard.
1SAM|23|1|Then they told David, saying, Behold, the Philistines fight against Keilah, and they rob the threshingfloors.
1SAM|23|2|Therefore David inquired of the LORD, saying, Shall I go and smite these Philistines? And the LORD said unto David, Go, and smite the Philistines, and save Keilah.
1SAM|23|3|And David's men said unto him, Behold, we be afraid here in Judah: how much more then if we come to Keilah against the armies of the Philistines?
1SAM|23|4|Then David inquired of the LORD yet again. And the LORD answered him and said, Arise, go down to Keilah; for I will deliver the Philistines into thine hand.
1SAM|23|5|So David and his men went to Keilah, and fought with the Philistines, and brought away their cattle, and smote them with a great slaughter. So David saved the inhabitants of Keilah.
1SAM|23|6|And it came to pass, when Abiathar the son of Ahimelech fled to David to Keilah, that he came down with an ephod in his hand.
1SAM|23|7|And it was told Saul that David was come to Keilah. And Saul said, God hath delivered him into mine hand; for he is shut in, by entering into a town that hath gates and bars.
1SAM|23|8|And Saul called all the people together to war, to go down to Keilah, to besiege David and his men.
1SAM|23|9|And David knew that Saul secretly practiced mischief against him; and he said to Abiathar the priest, Bring hither the ephod.
1SAM|23|10|Then said David, O LORD God of Israel, thy servant hath certainly heard that Saul seeketh to come to Keilah, to destroy the city for my sake.
1SAM|23|11|Will the men of Keilah deliver me up into his hand? will Saul come down, as thy servant hath heard? O LORD God of Israel, I beseech thee, tell thy servant. And the LORD said, He will come down.
1SAM|23|12|Then said David, Will the men of Keilah deliver me and my men into the hand of Saul? And the LORD said, They will deliver thee up.
1SAM|23|13|Then David and his men, which were about six hundred, arose and departed out of Keilah, and went whithersoever they could go. And it was told Saul that David was escaped from Keilah; and he forbare to go forth.
1SAM|23|14|And David abode in the wilderness in strong holds, and remained in a mountain in the wilderness of Ziph. And Saul sought him every day, but God delivered him not into his hand.
1SAM|23|15|And David saw that Saul was come out to seek his life: and David was in the wilderness of Ziph in a wood.
1SAM|23|16|And Jonathan Saul's son arose, and went to David into the wood, and strengthened his hand in God.
1SAM|23|17|And he said unto him, Fear not: for the hand of Saul my father shall not find thee; and thou shalt be king over Israel, and I shall be next unto thee; and that also Saul my father knoweth.
1SAM|23|18|And they two made a covenant before the LORD: and David abode in the wood, and Jonathan went to his house.
1SAM|23|19|Then came up the Ziphites to Saul to Gibeah, saying, Doth not David hide himself with us in strong holds in the wood, in the hill of Hachilah, which is on the south of Jeshimon?
1SAM|23|20|Now therefore, O king, come down according to all the desire of thy soul to come down; and our part shall be to deliver him into the king's hand.
1SAM|23|21|And Saul said, Blessed be ye of the LORD; for ye have compassion on me.
1SAM|23|22|Go, I pray you, prepare yet, and know and see his place where his haunt is, and who hath seen him there: for it is told me that he dealeth very subtilly.
1SAM|23|23|See therefore, and take knowledge of all the lurking places where he hideth himself, and come ye again to me with the certainty, and I will go with you: and it shall come to pass, if he be in the land, that I will search him out throughout all the thousands of Judah.
1SAM|23|24|And they arose, and went to Ziph before Saul: but David and his men were in the wilderness of Maon, in the plain on the south of Jeshimon.
1SAM|23|25|Saul also and his men went to seek him. And they told David; wherefore he came down into a rock, and abode in the wilderness of Maon. And when Saul heard that, he pursued after David in the wilderness of Maon.
1SAM|23|26|And Saul went on this side of the mountain, and David and his men on that side of the mountain: and David made haste to get away for fear of Saul; for Saul and his men compassed David and his men round about to take them.
1SAM|23|27|But there came a messenger unto Saul, saying, Haste thee, and come; for the Philistines have invaded the land.
1SAM|23|28|Wherefore Saul returned from pursuing after David, and went against the Philistines: therefore they called that place Selahammahlekoth.
1SAM|23|29|And David went up from thence, and dwelt in strong holds at Engedi.
1SAM|24|1|And it came to pass, when Saul was returned from following the Philistines, that it was told him, saying, Behold, David is in the wilderness of Engedi.
1SAM|24|2|Then Saul took three thousand chosen men out of all Israel, and went to seek David and his men upon the rocks of the wild goats.
1SAM|24|3|And he came to the sheepcotes by the way, where was a cave; and Saul went in to cover his feet: and David and his men remained in the sides of the cave.
1SAM|24|4|And the men of David said unto him, Behold the day of which the LORD said unto thee, Behold, I will deliver thine enemy into thine hand, that thou mayest do to him as it shall seem good unto thee. Then David arose, and cut off the skirt of Saul's robe privily.
1SAM|24|5|And it came to pass afterward, that David's heart smote him, because he had cut off Saul's skirt.
1SAM|24|6|And he said unto his men, The LORD forbid that I should do this thing unto my master, the LORD's anointed, to stretch forth mine hand against him, seeing he is the anointed of the LORD.
1SAM|24|7|So David stayed his servants with these words, and suffered them not to rise against Saul. But Saul rose up out of the cave, and went on his way.
1SAM|24|8|David also arose afterward, and went out of the cave, and cried after Saul, saying, My lord the king. And when Saul looked behind him, David stooped with his face to the earth, and bowed himself.
1SAM|24|9|And David said to Saul, Wherefore hearest thou men's words, saying, Behold, David seeketh thy hurt?
1SAM|24|10|Behold, this day thine eyes have seen how that the LORD had delivered thee to day into mine hand in the cave: and some bade me kill thee: but mine eye spared thee; and I said, I will not put forth mine hand against my lord; for he is the LORD's anointed.
1SAM|24|11|Moreover, my father, see, yea, see the skirt of thy robe in my hand: for in that I cut off the skirt of thy robe, and killed thee not, know thou and see that there is neither evil nor transgression in mine hand, and I have not sinned against thee; yet thou huntest my soul to take it.
1SAM|24|12|The LORD judge between me and thee, and the LORD avenge me of thee: but mine hand shall not be upon thee.
1SAM|24|13|As saith the proverb of the ancients, Wickedness proceedeth from the wicked: but mine hand shall not be upon thee.
1SAM|24|14|After whom is the king of Israel come out? after whom dost thou pursue? after a dead dog, after a flea.
1SAM|24|15|The LORD therefore be judge, and judge between me and thee, and see, and plead my cause, and deliver me out of thine hand.
1SAM|24|16|And it came to pass, when David had made an end of speaking these words unto Saul, that Saul said, Is this thy voice, my son David? And Saul lifted up his voice, and wept.
1SAM|24|17|And he said to David, Thou art more righteous than I: for thou hast rewarded me good, whereas I have rewarded thee evil.
1SAM|24|18|And thou hast showed this day how that thou hast dealt well with me: forasmuch as when the LORD had delivered me into thine hand, thou killedst me not.
1SAM|24|19|For if a man find his enemy, will he let him go well away? wherefore the LORD reward thee good for that thou hast done unto me this day.
1SAM|24|20|And now, behold, I know well that thou shalt surely be king, and that the kingdom of Israel shall be established in thine hand.
1SAM|24|21|Swear now therefore unto me by the LORD, that thou wilt not cut off my seed after me, and that thou wilt not destroy my name out of my father's house.
1SAM|24|22|And David sware unto Saul. And Saul went home; but David and his men gat them up unto the hold.
1SAM|25|1|And Samuel died; and all the Israelites were gathered together, and lamented him, and buried him in his house at Ramah. And David arose, and went down to the wilderness of Paran.
1SAM|25|2|And there was a man in Maon, whose possessions were in Carmel; and the man was very great, and he had three thousand sheep, and a thousand goats: and he was shearing his sheep in Carmel.
1SAM|25|3|Now the name of the man was Nabal; and the name of his wife Abigail: and she was a woman of good understanding, and of a beautiful countenance: but the man was churlish and evil in his doings; and he was of the house of Caleb.
1SAM|25|4|And David heard in the wilderness that Nabal did shear his sheep.
1SAM|25|5|And David sent out ten young men, and David said unto the young men, Get you up to Carmel, and go to Nabal, and greet him in my name:
1SAM|25|6|And thus shall ye say to him that liveth in prosperity, Peace be both to thee, and peace be to thine house, and peace be unto all that thou hast.
1SAM|25|7|And now I have heard that thou hast shearers: now thy shepherds which were with us, we hurt them not, neither was there ought missing unto them, all the while they were in Carmel.
1SAM|25|8|Ask thy young men, and they will show thee. Wherefore let the young men find favor in thine eyes: for we come in a good day: give, I pray thee, whatsoever cometh to thine hand unto thy servants, and to thy son David.
1SAM|25|9|And when David's young men came, they spake to Nabal according to all those words in the name of David, and ceased.
1SAM|25|10|And Nabal answered David's servants, and said, Who is David? and who is the son of Jesse? there be many servants now a days that break away every man from his master.
1SAM|25|11|Shall I then take my bread, and my water, and my flesh that I have killed for my shearers, and give it unto men, whom I know not whence they be?
1SAM|25|12|So David's young men turned their way, and went again, and came and told him all those sayings.
1SAM|25|13|And David said unto his men, Gird ye on every man his sword. And they girded on every man his sword; and David also girded on his sword: and there went up after David about four hundred men; and two hundred abode by the stuff.
1SAM|25|14|But one of the young men told Abigail, Nabal's wife, saying, Behold, David sent messengers out of the wilderness to salute our master; and he railed on them.
1SAM|25|15|But the men were very good unto us, and we were not hurt, neither missed we any thing, as long as we were conversant with them, when we were in the fields:
1SAM|25|16|They were a wall unto us both by night and day, all the while we were with them keeping the sheep.
1SAM|25|17|Now therefore know and consider what thou wilt do; for evil is determined against our master, and against all his household: for he is such a son of Belial, that a man cannot speak to him.
1SAM|25|18|Then Abigail made haste, and took two hundred loaves, and two bottles of wine, and five sheep ready dressed, and five measures of parched corn, and an hundred clusters of raisins, and two hundred cakes of figs, and laid them on asses.
1SAM|25|19|And she said unto her servants, Go on before me; behold, I come after you. But she told not her husband Nabal.
1SAM|25|20|And it was so, as she rode on the ass, that she came down by the covert on the hill, and, behold, David and his men came down against her; and she met them.
1SAM|25|21|Now David had said, Surely in vain have I kept all that this fellow hath in the wilderness, so that nothing was missed of all that pertained unto him: and he hath requited me evil for good.
1SAM|25|22|So and more also do God unto the enemies of David, if I leave of all that pertain to him by the morning light any that pisseth against the wall.
1SAM|25|23|And when Abigail saw David, she hasted, and lighted off the ass, and fell before David on her face, and bowed herself to the ground,
1SAM|25|24|And fell at his feet, and said, Upon me, my lord, upon me let this iniquity be: and let thine handmaid, I pray thee, speak in thine audience, and hear the words of thine handmaid.
1SAM|25|25|Let not my lord, I pray thee, regard this man of Belial, even Nabal: for as his name is, so is he; Nabal is his name, and folly is with him: but I thine handmaid saw not the young men of my lord, whom thou didst send.
1SAM|25|26|Now therefore, my lord, as the LORD liveth, and as thy soul liveth, seeing the LORD hath withholden thee from coming to shed blood, and from avenging thyself with thine own hand, now let thine enemies, and they that seek evil to my lord, be as Nabal.
1SAM|25|27|And now this blessing which thine handmaid hath brought unto my lord, let it even be given unto the young men that follow my lord.
1SAM|25|28|I pray thee, forgive the trespass of thine handmaid: for the LORD will certainly make my lord a sure house; because my lord fighteth the battles of the LORD, and evil hath not been found in thee all thy days.
1SAM|25|29|Yet a man is risen to pursue thee, and to seek thy soul: but the soul of my lord shall be bound in the bundle of life with the LORD thy God; and the souls of thine enemies, them shall he sling out, as out of the middle of a sling.
1SAM|25|30|And it shall come to pass, when the LORD shall have done to my lord according to all the good that he hath spoken concerning thee, and shall have appointed thee ruler over Israel;
1SAM|25|31|That this shall be no grief unto thee, nor offense of heart unto my lord, either that thou hast shed blood causeless, or that my lord hath avenged himself: but when the LORD shall have dealt well with my lord, then remember thine handmaid.
1SAM|25|32|And David said to Abigail, Blessed be the LORD God of Israel, which sent thee this day to meet me:
1SAM|25|33|And blessed be thy advice, and blessed be thou, which hast kept me this day from coming to shed blood, and from avenging myself with mine own hand.
1SAM|25|34|For in very deed, as the LORD God of Israel liveth, which hath kept me back from hurting thee, except thou hadst hasted and come to meet me, surely there had not been left unto Nabal by the morning light any that pisseth against the wall.
1SAM|25|35|So David received of her hand that which she had brought him, and said unto her, Go up in peace to thine house; see, I have hearkened to thy voice, and have accepted thy person.
1SAM|25|36|And Abigail came to Nabal; and, behold, he held a feast in his house, like the feast of a king; and Nabal's heart was merry within him, for he was very drunken: wherefore she told him nothing, less or more, until the morning light.
1SAM|25|37|But it came to pass in the morning, when the wine was gone out of Nabal, and his wife had told him these things, that his heart died within him, and he became as a stone.
1SAM|25|38|And it came to pass about ten days after, that the LORD smote Nabal, that he died.
1SAM|25|39|And when David heard that Nabal was dead, he said, Blessed be the LORD, that hath pleaded the cause of my reproach from the hand of Nabal, and hath kept his servant from evil: for the LORD hath returned the wickedness of Nabal upon his own head. And David sent and communed with Abigail, to take her to him to wife.
1SAM|25|40|And when the servants of David were come to Abigail to Carmel, they spake unto her, saying, David sent us unto thee, to take thee to him to wife.
1SAM|25|41|And she arose, and bowed herself on her face to the earth, and said, Behold, let thine handmaid be a servant to wash the feet of the servants of my lord.
1SAM|25|42|And Abigail hasted, and arose and rode upon an ass, with five damsels of hers that went after her; and she went after the messengers of David, and became his wife.
1SAM|25|43|David also took Ahinoam of Jezreel; and they were also both of them his wives.
1SAM|25|44|But Saul had given Michal his daughter, David's wife, to Phalti the son of Laish, which was of Gallim.
1SAM|26|1|And the Ziphites came unto Saul to Gibeah, saying, Doth not David hide himself in the hill of Hachilah, which is before Jeshimon?
1SAM|26|2|Then Saul arose, and went down to the wilderness of Ziph, having three thousand chosen men of Israel with him, to seek David in the wilderness of Ziph.
1SAM|26|3|And Saul pitched in the hill of Hachilah, which is before Jeshimon, by the way. But David abode in the wilderness, and he saw that Saul came after him into the wilderness.
1SAM|26|4|David therefore sent out spies, and understood that Saul was come in very deed.
1SAM|26|5|And David arose, and came to the place where Saul had pitched: and David beheld the place where Saul lay, and Abner the son of Ner, the captain of his host: and Saul lay in the trench, and the people pitched round about him.
1SAM|26|6|Then answered David and said to Ahimelech the Hittite, and to Abishai the son of Zeruiah, brother to Joab, saying, Who will go down with me to Saul to the camp? And Abishai said, I will go down with thee.
1SAM|26|7|So David and Abishai came to the people by night: and, behold, Saul lay sleeping within the trench, and his spear stuck in the ground at his bolster: but Abner and the people lay round about him.
1SAM|26|8|Then said Abishai to David, God hath delivered thine enemy into thine hand this day: now therefore let me smite him, I pray thee, with the spear even to the earth at once, and I will not smite him the second time.
1SAM|26|9|And David said to Abishai, Destroy him not: for who can stretch forth his hand against the LORD's anointed, and be guiltless?
1SAM|26|10|David said furthermore, As the LORD liveth, the LORD shall smite him; or his day shall come to die; or he shall descend into battle, and perish.
1SAM|26|11|The LORD forbid that I should stretch forth mine hand against the LORD's anointed: but, I pray thee, take thou now the spear that is at his bolster, and the cruse of water, and let us go.
1SAM|26|12|So David took the spear and the cruse of water from Saul's bolster; and they gat them away, and no man saw it, nor knew it, neither awaked: for they were all asleep; because a deep sleep from the LORD was fallen upon them.
1SAM|26|13|Then David went over to the other side, and stood on the top of an hill afar off; a great space being between them:
1SAM|26|14|And David cried to the people, and to Abner the son of Ner, saying, Answerest thou not, Abner? Then Abner answered and said, Who art thou that criest to the king?
1SAM|26|15|And David said to Abner, Art not thou a valiant man? and who is like to thee in Israel? wherefore then hast thou not kept thy lord the king? for there came one of the people in to destroy the king thy lord.
1SAM|26|16|This thing is not good that thou hast done. As the LORD liveth, ye are worthy to die, because ye have not kept your master, the LORD's anointed. And now see where the king's spear is, and the cruse of water that was at his bolster.
1SAM|26|17|And Saul knew David's voice, and said, Is this thy voice, my son David? And David said, It is my voice, my lord, O king.
1SAM|26|18|And he said, Wherefore doth my lord thus pursue after his servant? for what have I done? or what evil is in mine hand?
1SAM|26|19|Now therefore, I pray thee, let my lord the king hear the words of his servant. If the LORD have stirred thee up against me, let him accept an offering: but if they be the children of men, cursed be they before the LORD; for they have driven me out this day from abiding in the inheritance of the LORD, saying, Go, serve other gods.
1SAM|26|20|Now therefore, let not my blood fall to the earth before the face of the LORD: for the king of Israel is come out to seek a flea, as when one doth hunt a partridge in the mountains.
1SAM|26|21|Then said Saul, I have sinned: return, my son David: for I will no more do thee harm, because my soul was precious in thine eyes this day: behold, I have played the fool, and have erred exceedingly.
1SAM|26|22|And David answered and said, Behold the king's spear! and let one of the young men come over and fetch it.
1SAM|26|23|The LORD render to every man his righteousness and his faithfulness; for the LORD delivered thee into my hand to day, but I would not stretch forth mine hand against the LORD's anointed.
1SAM|26|24|And, behold, as thy life was much set by this day in mine eyes, so let my life be much set by in the eyes of the LORD, and let him deliver me out of all tribulation.
1SAM|26|25|Then Saul said to David, Blessed be thou, my son David: thou shalt both do great things, and also shalt still prevail. So David went on his way, and Saul returned to his place.
1SAM|27|1|And David said in his heart, I shall now perish one day by the hand of Saul: there is nothing better for me than that I should speedily escape into the land of the Philistines; and Saul shall despair of me, to seek me any more in any coast of Israel: so shall I escape out of his hand.
1SAM|27|2|And David arose, and he passed over with the six hundred men that were with him unto Achish, the son of Maoch, king of Gath.
1SAM|27|3|And David dwelt with Achish at Gath, he and his men, every man with his household, even David with his two wives, Ahinoam the Jezreelitess, and Abigail the Carmelitess, Nabal's wife.
1SAM|27|4|And it was told Saul that David was fled to Gath: and he sought no more again for him.
1SAM|27|5|And David said unto Achish, If I have now found grace in thine eyes, let them give me a place in some town in the country, that I may dwell there: for why should thy servant dwell in the royal city with thee?
1SAM|27|6|Then Achish gave him Ziklag that day: wherefore Ziklag pertaineth unto the kings of Judah unto this day.
1SAM|27|7|And the time that David dwelt in the country of the Philistines was a full year and four months.
1SAM|27|8|And David and his men went up, and invaded the Geshurites, and the Gezrites, and the Amalekites: for those nations were of old the inhabitants of the land, as thou goest to Shur, even unto the land of Egypt.
1SAM|27|9|And David smote the land, and left neither man nor woman alive, and took away the sheep, and the oxen, and the asses, and the camels, and the apparel, and returned, and came to Achish.
1SAM|27|10|And Achish said, Whither have ye made a road to day? And David said, Against the south of Judah, and against the south of the Jerahmeelites, and against the south of the Kenites.
1SAM|27|11|And David saved neither man nor woman alive, to bring tidings to Gath, saying, Lest they should tell on us, saying, So did David, and so will be his manner all the while he dwelleth in the country of the Philistines.
1SAM|27|12|And Achish believed David, saying, He hath made his people Israel utterly to abhor him; therefore he shall be my servant for ever.
1SAM|28|1|And it came to pass in those days, that the Philistines gathered their armies together for warfare, to fight with Israel. And Achish said unto David, Know thou assuredly, that thou shalt go out with me to battle, thou and thy men.
1SAM|28|2|And David said to Achish, Surely thou shalt know what thy servant can do. And Achish said to David, Therefore will I make thee keeper of mine head for ever.
1SAM|28|3|Now Samuel was dead, and all Israel had lamented him, and buried him in Ramah, even in his own city. And Saul had put away those that had familiar spirits, and the wizards, out of the land.
1SAM|28|4|And the Philistines gathered themselves together, and came and pitched in Shunem: and Saul gathered all Israel together, and they pitched in Gilboa.
1SAM|28|5|And when Saul saw the host of the Philistines, he was afraid, and his heart greatly trembled.
1SAM|28|6|And when Saul inquired of the LORD, the LORD answered him not, neither by dreams, nor by Urim, nor by prophets.
1SAM|28|7|Then said Saul unto his servants, Seek me a woman that hath a familiar spirit, that I may go to her, and inquire of her. And his servants said to him, Behold, there is a woman that hath a familiar spirit at Endor.
1SAM|28|8|And Saul disguised himself, and put on other raiment, and he went, and two men with him, and they came to the woman by night: and he said, I pray thee, divine unto me by the familiar spirit, and bring me him up, whom I shall name unto thee.
1SAM|28|9|And the woman said unto him, Behold, thou knowest what Saul hath done, how he hath cut off those that have familiar spirits, and the wizards, out of the land: wherefore then layest thou a snare for my life, to cause me to die?
1SAM|28|10|And Saul sware to her by the LORD, saying, As the LORD liveth, there shall no punishment happen to thee for this thing.
1SAM|28|11|Then said the woman, Whom shall I bring up unto thee? And he said, Bring me up Samuel.
1SAM|28|12|And when the woman saw Samuel, she cried with a loud voice: and the woman spake to Saul, saying, Why hast thou deceived me? for thou art Saul.
1SAM|28|13|And the king said unto her, Be not afraid: for what sawest thou? And the woman said unto Saul, I saw gods ascending out of the earth.
1SAM|28|14|And he said unto her, What form is he of? And she said, An old man cometh up; and he is covered with a mantle. And Saul perceived that it was Samuel, and he stooped with his face to the ground, and bowed himself.
1SAM|28|15|And Samuel said to Saul, Why hast thou disquieted me, to bring me up? And Saul answered, I am sore distressed; for the Philistines make war against me, and God is departed from me, and answereth me no more, neither by prophets, nor by dreams: therefore I have called thee, that thou mayest make known unto me what I shall do.
1SAM|28|16|Then said Samuel, Wherefore then dost thou ask of me, seeing the LORD is departed from thee, and is become thine enemy?
1SAM|28|17|And the LORD hath done to him, as he spake by me: for the LORD hath rent the kingdom out of thine hand, and given it to thy neighbor, even to David:
1SAM|28|18|Because thou obeyedst not the voice of the LORD, nor executedst his fierce wrath upon Amalek, therefore hath the LORD done this thing unto thee this day.
1SAM|28|19|Moreover the LORD will also deliver Israel with thee into the hand of the Philistines: and to morrow shalt thou and thy sons be with me: the LORD also shall deliver the host of Israel into the hand of the Philistines.
1SAM|28|20|Then Saul fell straightway all along on the earth, and was sore afraid, because of the words of Samuel: and there was no strength in him; for he had eaten no bread all the day, nor all the night.
1SAM|28|21|And the woman came unto Saul, and saw that he was sore troubled, and said unto him, Behold, thine handmaid hath obeyed thy voice, and I have put my life in my hand, and have hearkened unto thy words which thou spakest unto me.
1SAM|28|22|Now therefore, I pray thee, hearken thou also unto the voice of thine handmaid, and let me set a morsel of bread before thee; and eat, that thou mayest have strength, when thou goest on thy way.
1SAM|28|23|But he refused, and said, I will not eat. But his servants, together with the woman, compelled him; and he hearkened unto their voice. So he arose from the earth, and sat upon the bed.
1SAM|28|24|And the woman had a fat calf in the house; and she hasted, and killed it, and took flour, and kneaded it, and did bake unleavened bread thereof:
1SAM|28|25|And she brought it before Saul, and before his servants; and they did eat. Then they rose up, and went away that night.
1SAM|29|1|Now the Philistines gathered together all their armies to Aphek: and the Israelites pitched by a fountain which is in Jezreel.
1SAM|29|2|And the lords of the Philistines passed on by hundreds, and by thousands: but David and his men passed on in the rearward with Achish.
1SAM|29|3|Then said the princes of the Philistines, What do these Hebrews here? And Achish said unto the princes of the Philistines, Is not this David, the servant of Saul the king of Israel, which hath been with me these days, or these years, and I have found no fault in him since he fell unto me unto this day?
1SAM|29|4|And the princes of the Philistines were wroth with him; and the princes of the Philistines said unto him, Make this fellow return, that he may go again to his place which thou hast appointed him, and let him not go down with us to battle, lest in the battle he be an adversary to us: for wherewith should he reconcile himself unto his master? should it not be with the heads of these men?
1SAM|29|5|Is not this David, of whom they sang one to another in dances, saying, Saul slew his thousands, and David his ten thousands?
1SAM|29|6|Then Achish called David, and said unto him, Surely, as the LORD liveth, thou hast been upright, and thy going out and thy coming in with me in the host is good in my sight: for I have not found evil in thee since the day of thy coming unto me unto this day: nevertheless the lords favor thee not.
1SAM|29|7|Wherefore now return, and go in peace, that thou displease not the lords of the Philistines.
1SAM|29|8|And David said unto Achish, But what have I done? and what hast thou found in thy servant so long as I have been with thee unto this day, that I may not go fight against the enemies of my lord the king?
1SAM|29|9|And Achish answered and said to David, I know that thou art good in my sight, as an angel of God: notwithstanding the princes of the Philistines have said, He shall not go up with us to the battle.
1SAM|29|10|Wherefore now rise up early in the morning with thy master's servants that are come with thee: and as soon as ye be up early in the morning, and have light, depart.
1SAM|29|11|So David and his men rose up early to depart in the morning, to return into the land of the Philistines. And the Philistines went up to Jezreel.
1SAM|30|1|And it came to pass, when David and his men were come to Ziklag on the third day, that the Amalekites had invaded the south, and Ziklag, and smitten Ziklag, and burned it with fire;
1SAM|30|2|And had taken the women captives, that were therein: they slew not any, either great or small, but carried them away, and went on their way.
1SAM|30|3|So David and his men came to the city, and, behold, it was burned with fire; and their wives, and their sons, and their daughters, were taken captives.
1SAM|30|4|Then David and the people that were with him lifted up their voice and wept, until they had no more power to weep.
1SAM|30|5|And David's two wives were taken captives, Ahinoam the Jezreelitess, and Abigail the wife of Nabal the Carmelite.
1SAM|30|6|And David was greatly distressed; for the people spake of stoning him, because the soul of all the people was grieved, every man for his sons and for his daughters: but David encouraged himself in the LORD his God.
1SAM|30|7|And David said to Abiathar the priest, Ahimelech's son, I pray thee, bring me hither the ephod. And Abiathar brought thither the ephod to David.
1SAM|30|8|And David inquired at the LORD, saying, Shall I pursue after this troop? shall I overtake them? And he answered him, Pursue: for thou shalt surely overtake them, and without fail recover all.
1SAM|30|9|So David went, he and the six hundred men that were with him, and came to the brook Besor, where those that were left behind stayed.
1SAM|30|10|But David pursued, he and four hundred men: for two hundred abode behind, which were so faint that they could not go over the brook Besor.
1SAM|30|11|And they found an Egyptian in the field, and brought him to David, and gave him bread, and he did eat; and they made him drink water;
1SAM|30|12|And they gave him a piece of a cake of figs, and two clusters of raisins: and when he had eaten, his spirit came again to him: for he had eaten no bread, nor drunk any water, three days and three nights.
1SAM|30|13|And David said unto him, To whom belongest thou? and whence art thou? And he said, I am a young man of Egypt, servant to an Amalekite; and my master left me, because three days agone I fell sick.
1SAM|30|14|We made an invasion upon the south of the Cherethites, and upon the coast which belongeth to Judah, and upon the south of Caleb; and we burned Ziklag with fire.
1SAM|30|15|And David said to him, Canst thou bring me down to this company? And he said, Swear unto me by God, that thou wilt neither kill me, nor deliver me into the hands of my master, and I will bring thee down to this company.
1SAM|30|16|And when he had brought him down, behold, they were spread abroad upon all the earth, eating and drinking, and dancing, because of all the great spoil that they had taken out of the land of the Philistines, and out of the land of Judah.
1SAM|30|17|And David smote them from the twilight even unto the evening of the next day: and there escaped not a man of them, save four hundred young men, which rode upon camels, and fled.
1SAM|30|18|And David recovered all that the Amalekites had carried away: and David rescued his two wives.
1SAM|30|19|And there was nothing lacking to them, neither small nor great, neither sons nor daughters, neither spoil, nor any thing that they had taken to them: David recovered all.
1SAM|30|20|And David took all the flocks and the herds, which they drave before those other cattle, and said, This is David's spoil.
1SAM|30|21|And David came to the two hundred men, which were so faint that they could not follow David, whom they had made also to abide at the brook Besor: and they went forth to meet David, and to meet the people that were with him: and when David came near to the people, he saluted them.
1SAM|30|22|Then answered all the wicked men and men of Belial, of those that went with David, and said, Because they went not with us, we will not give them ought of the spoil that we have recovered, save to every man his wife and his children, that they may lead them away, and depart.
1SAM|30|23|Then said David, Ye shall not do so, my brethren, with that which the LORD hath given us, who hath preserved us, and delivered the company that came against us into our hand.
1SAM|30|24|For who will hearken unto you in this matter? but as his part is that goeth down to the battle, so shall his part be that tarrieth by the stuff: they shall part alike.
1SAM|30|25|And it was so from that day forward, that he made it a statute and an ordinance for Israel unto this day.
1SAM|30|26|And when David came to Ziklag, he sent of the spoil unto the elders of Judah, even to his friends, saying, Behold a present for you of the spoil of the enemies of the LORD;
1SAM|30|27|To them which were in Bethel, and to them which were in south Ramoth, and to them which were in Jattir,
1SAM|30|28|And to them which were in Aroer, and to them which were in Siphmoth, and to them which were in Eshtemoa,
1SAM|30|29|And to them which were in Rachal, and to them which were in the cities of the Jerahmeelites, and to them which were in the cities of the Kenites,
1SAM|30|30|And to them which were in Hormah, and to them which were in Chorashan, and to them which were in Athach,
1SAM|30|31|And to them which were in Hebron, and to all the places where David himself and his men were wont to haunt.
1SAM|31|1|Now the Philistines fought against Israel: and the men of Israel fled from before the Philistines, and fell down slain in mount Gilboa.
1SAM|31|2|And the Philistines followed hard upon Saul and upon his sons; and the Philistines slew Jonathan, and Abinadab, and Melchishua, Saul's sons.
1SAM|31|3|And the battle went sore against Saul, and the archers hit him; and he was sore wounded of the archers.
1SAM|31|4|Then said Saul unto his armourbearer, Draw thy sword, and thrust me through therewith; lest these uncircumcised come and thrust me through, and abuse me. But his armourbearer would not; for he was sore afraid. Therefore Saul took a sword, and fell upon it.
1SAM|31|5|And when his armourbearer saw that Saul was dead, he fell likewise upon his sword, and died with him.
1SAM|31|6|So Saul died, and his three sons, and his armourbearer, and all his men, that same day together.
1SAM|31|7|And when the men of Israel that were on the other side of the valley, and they that were on the other side Jordan, saw that the men of Israel fled, and that Saul and his sons were dead, they forsook the cities, and fled; and the Philistines came and dwelt in them.
1SAM|31|8|And it came to pass on the morrow, when the Philistines came to strip the slain, that they found Saul and his three sons fallen in mount Gilboa.
1SAM|31|9|And they cut off his head, and stripped off his armor, and sent into the land of the Philistines round about, to publish it in the house of their idols, and among the people.
1SAM|31|10|And they put his armor in the house of Ashtaroth: and they fastened his body to the wall of Bethshan.
1SAM|31|11|And when the inhabitants of Jabeshgilead heard of that which the Philistines had done to Saul;
1SAM|31|12|All the valiant men arose, and went all night, and took the body of Saul and the bodies of his sons from the wall of Bethshan, and came to Jabesh, and burnt them there.
1SAM|31|13|And they took their bones, and buried them under a tree at Jabesh, and fasted seven days.
