JOB|1|1|Був чоловік у країні Уц, на ім'я йому Йов. І був чоловік цей невинний та праведний, і він Бога боявся, а від злого втікав.
JOB|1|2|І народилися йому семеро синів та три дочки.
JOB|1|3|А маєток його був: сім тисяч худоби дрібної, і три тисячі верблюдів, і п'ять сотень пар худоби великої, і п'ять сотень ослиць та дуже багато рабів. І був цей чоловік більший від усіх синів сходу.
JOB|1|4|А сини його ходили один до одного, і справляли гостину в домі того, чий був день. І посилали вони, і кликали трьох своїх сестер, щоб їсти та пити із ними.
JOB|1|5|І бувало, як миналося коло бенкетних днів, то Йов посилав за дітьми й освячував їх, і вставав він рано вранці, і приносив цілопалення за числом їх усіх, бо Йов казав: Може згрішили сини мої, і зневажили Бога в серці своєму. Так робив Йов по всі дні.
JOB|1|6|І сталося одного дня, і поприходили Божі сини, щоб стати при Господі. І прийшов поміж ними й сатана.
JOB|1|7|І сказав Господь до сатани: Звідки ти йдеш? А сатана відповів Господеві й сказав: Я мандрував по землі та й перейшов її.
JOB|1|8|І сказав Господь до сатани: Чи звернув ти увагу на раба Мого Йова? Бо немає такого, як він, на землі: муж він невинний та праведний, що Бога боїться, а від злого втікає.
JOB|1|9|І відповів сатана Господеві й сказав: Чи ж Йов дармо боїться Бога?
JOB|1|10|Чи ж Ти не забезпечив його, і дім його, і все, що його? Чин його рук Ти поблагословив, а маєток його поширився по краю.
JOB|1|11|Але простягни тільки руку Свою, і доторкнися до всього, що його, чи він не зневажить Тебе перед лицем Твоїм?
JOB|1|12|І сказав Господь до сатани: Ось усе, що його, у твоїй руці, тільки на нього самого не простягай своєї руки! І пішов сатана від лиця Господнього.
JOB|1|13|І сталося одного дня, коли сини його та дочки його їли та вино пили в домі свого первородженого брата,
JOB|1|14|то прибіг до Йова посланець та й сказав: Худоба велика орала, а ослиці паслися при них.
JOB|1|15|Аж тут напали сабеї й позабирали їх, а слуг повбивали вістрям меча. І втік тільки я сам, щоб донести тобі...
JOB|1|16|Він ще говорив, аж прибігає інший та й каже: З неба спав Божий огонь, і спалив отару та слуг, та й пожер їх... А втік тільки я сам, щоб донести тобі...
JOB|1|17|Він ще говорив, аж біжить ще інший та й каже: Халдеї поділилися на три відділи, і напали на верблюдів, та й позабирали їх, а слуг повбивали вістрям меча... І втік тільки я сам, щоб донести тобі...
JOB|1|18|Поки він говорив, аж надбігає ще інший та й каже: Сини твої та дочки твої їли та вино пили в домі свого первородженого брата.
JOB|1|19|Аж раптово надійшов великий вітер з боку пустині, та й ударив на чотири роги дому, і він упав на юнаків, і вони повмирали... І втік тільки я сам, щоб донести тобі...
JOB|1|20|І встав Йов, і роздер плаща свого, й обстриг свою голову, та й упав на землю, і поклонився,
JOB|1|21|та й сказав: Я вийшов нагий із утроби матері своєї, і нагий повернусь туди, в землю! Господь дав, і Господь узяв... Нехай буде благословенне Господнє Ім'я!
JOB|1|22|При всьому цьому Йов не згрішив, і не сказав на Бога нічого безумного!
JOB|2|1|І сталося одного дня, і поприходили Божі сини, щоб стати перед Господом: і прийшов також сатана поміж ними, щоб стати перед Господом.
JOB|2|2|І сказав Господь до сатани: Звідки ти йдеш? А сатана відповів Господеві й сказав:
JOB|2|3|І сказав Господь до сатани: Чи звернув ти увагу на раба Мого Йова? Бо немає такого, як він, на землі: муж він невинний та праведний, який Бога боїться, а від злого втікає. І він ще тримається міцно в своїй невинності, а ти намовляв був Мене на нього, щоб без приводу його зруйнувати...
JOB|2|4|І відповів сатана Господеві й сказав: Шкіра за шкіру, і все, що хто має, віддасть він за душу свою.
JOB|2|5|Але простягни но Ти руку Свою, і доторкнись до костей його та до тіла його, чи він не зневажить Тебе перед лицем Твоїм?
JOB|2|6|І сказав Господь до сатани: Ось він у руці твоїй, тільки душу його бережи!
JOB|2|7|І вийшов сатана від лиця Господнього, та й ударив Йова злим гнояком від стопи ноги його аж до його черепа...
JOB|2|8|А той узяв собі черепка, щоб шкребти себе. І він сидів серед попелу...
JOB|2|9|І сказала йому його жінка: Ти ще міцно тримаєшся в невинності своїй? Прокляни Бога і помреш!...
JOB|2|10|А він до неї відказав: Ти говориш отак, як говорить яка з божевільних!... Чи ж ми будем приймати від Бога добре, а злого не приймем? При всьому тому Йов не згрішив своїми устами...
JOB|2|11|І почули троє приятелів Йовових про все те нещастя, що прийшло на нього, і поприходили кожен з місця свого: теманянин Еліфаз, шух'янин Біддад та нааматянин Цофар. І вмовилися вони прийти разом, щоб похитати головою над ним та потішити його.
JOB|2|12|І звели вони здалека очі свої, і не пізнали його... І піднесли вони голос свій, та й заголосили, і роздерли кожен одежу свою, і кидали порох над своїми головами аж до неба...
JOB|2|13|І сиділи вони з ним на землі сім день та сім ночей, і ніхто не промовив до нього ні слова, бо вони бачили, що біль його вельми великий...
JOB|3|1|По цьому відкрив Йов уста свої та й прокляв був свій день народження.
JOB|3|2|І Йов заговорив та й сказав:
JOB|3|3|Хай загине той день, що я в ньому родився, і та ніч, що сказала: Зачавсь чоловік!
JOB|3|4|Нехай стане цей день темнотою, нехай Бог з висоти не згадає його, і нехай не являється світло над ним!...
JOB|3|5|Бодай темрява й морок його заступили, бодай хмара над ним пробувала, бодай темнощі денні лякали його!...
JOB|3|6|Оця ніч бодай темність її обгорнула, нехай у днях року не буде названа вона, хай не ввійде вона в число місяців!...
JOB|3|7|Тож ця ніч нехай буде самітна, хай не прийде до неї співання!
JOB|3|8|Бодай її ті проклинали, що день проклинають, що левіятана готові збудити!
JOB|3|9|Хай потемніють зорі поранку її, нехай має надію на світло й не буде його, і хай вона не побачить тремтячих повік зорі ранньої,
JOB|3|10|бо вона не замкнула дверей нутра матернього, і не сховала страждання з очей моїх!...
JOB|3|11|Чому я не згинув в утробі? Як вийшов, із нутра то чому я не вмер?
JOB|3|12|Чого прийняли ті коліна мене? І нащо ті перса, які я був ссав?
JOB|3|13|Бо тепер я лежав би спокійно, я спав би, та був би мені відпочинок
JOB|3|14|з царями та з земними радниками, що гробниці будують собі,
JOB|3|15|або із князями, що золото мали, що доми свої сріблом наповнювали!...
JOB|3|16|Або чом я не ставсь недоноском прихованим, немов ті немовлята, що світла не бачили?
JOB|3|17|Там же безбожники перестають докучати, і спочивають там змученосилі,
JOB|3|18|разом з тим мають спокій ув'язнені, вони не почують вже крику гнобителя!...
JOB|3|19|Малий та великий там рівні, а раб вільний від пана свого...
JOB|3|20|І нащо Він струдженому дає світло, і життя гіркодухим,
JOB|3|21|що вичікують смерти й немає її, що її відкопали б, як скарби заховані,
JOB|3|22|тим, що радісно тішилися б, веселились, коли б знайшли гроба,
JOB|3|23|мужчині, якому дорога закрита, що Бог тінню закрив перед ним?...
JOB|3|24|Бо зідхання моє випереджує хліб мій, а зойки мої полились, як вода,
JOB|3|25|бо страх, що його я жахався, до мене прибув, і чого я боявся прийшло те мені...
JOB|3|26|Не знав я спокою й не був втихомирений, і я не відпочив, та нещастя прийшло!...
JOB|4|1|І відповів теманянин Еліфаз та й сказав:
JOB|4|2|Коли спробувать слово до тебе, чи мука не буде ще більша? Та хто стримати зможе слова?
JOB|4|3|Таж ти багатьох був навчав, а руки ослаблі зміцняв,
JOB|4|4|того, хто спотикавсь, підіймали слова твої, а коліна тремткі ти зміцняв!
JOB|4|5|А тепер, як нещастя на тебе найшло, то ти змучився, тебе досягло воно і ти налякався...
JOB|4|6|Хіба не була богобійність твоя за надію твою, за твоє сподівання невинність доріг твоїх?
JOB|4|7|Пригадай но, чи гинув невинний, і де праведні вигублені?
JOB|4|8|Як я бачив таких, що орали були беззаконня, та сіяли кривду, то й жали її:
JOB|4|9|вони гинуть від подиху Божого, і від духу гнівного Його погибають!
JOB|4|10|Левине ричання й рик лютого лева минає, і левчукам вилущаються зуби.
JOB|4|11|Гине лев, як немає здобичі, і левенята левиці втікають.
JOB|4|12|І закрадається слово до мене, і моє ухо почуло ось дещо від нього.
JOB|4|13|у роздумуваннях над нічними видіннями, коли міцний сон обіймає людей,
JOB|4|14|спіткав мене жах та тремтіння, і багато костей моїх він струсонув,
JOB|4|15|і дух перейшов по обличчі моїм, стало дуба волосся на тілі моїм...
JOB|4|16|Він стояв, але я не пізнав його вигляду, образ навпроти очей моїх був, і тихий голос почув я:
JOB|4|17|Хіба праведніша людина за Бога, хіба чоловік за свойого Творця є чистіший?
JOB|4|18|Таж рабам Своїм Він не йме віри, і накладає вину й на Своїх Анголів!
JOB|4|19|Що ж тоді мешканці глиняних хат, що в поросі їхня основа? Як міль, вони будуть розчавлені!
JOB|4|20|Вони товчені зранку до вечора, і без помочі гинуть назавжди...
JOB|4|21|Слава їхня минається з ними, вони помирають не в мудрості!...
JOB|5|1|Ану клич, чи є хто, щоб тобі відповів? І до кого з святих ти вдасися?
JOB|5|2|Бо гнів побиває безглуздого, а заздрощі смерть завдають нерозумному!
JOB|5|3|Я бачив безумного, як він розсівся, та зараз оселя його спорохнявіла...
JOB|5|4|Від спасіння далекі сини його, вони без рятунку почавлені будуть у брамі!
JOB|5|5|Його жниво голодний поїсть, і з-між терну його забере, і спрагнені ось поковтають маєток його!
JOB|5|6|Бо нещастя виходить не з пороху, а горе росте не з землі,
JOB|5|7|бо людина народжується на страждання, як іскри, щоб угору летіти...
JOB|5|8|А я б удавався до Бога, і на Бога б поклав свою справу,
JOB|5|9|Він чинить велике та недослідиме, предивне, якому немає числа,
JOB|5|10|бо Він дає дощ на поверхню землі, і на поля посилає Він воду,
JOB|5|11|щоб поставить низьких на високе, і зміцнити спасіння засмучених.
JOB|5|12|Він розвіює задуми хитрих, і не виконують плану їх руки,
JOB|5|13|Він мудрих лукавством їх ловить, і рада крутійська марною стає,
JOB|5|14|вдень знаходять вони темноту, а в полудень мацають, мов уночі!...
JOB|5|15|І Він від меча урятовує бідного, а з міцної руки бідаря,
JOB|5|16|і стається надія нужденному, і замкнула уста свої кривда!
JOB|5|17|Тож блаженна людина, яку Бог картає, і ти не цурайсь Всемогутнього кари:
JOB|5|18|Бо Він рану завдасть і перев'яже, Він ламає й вигоюють руки Його!
JOB|5|19|В шістьох лихах спасає тебе, а в сімох не діткне тебе зло:
JOB|5|20|Викупляє тебе Він від смерти за голоду, а в бою з рук меча.
JOB|5|21|Як бич язика запанує, сховаєшся ти, і не будеш боятись руїни, як прийде вона.
JOB|5|22|З насилля та з голоду будеш сміятись, а земної звірини не бійся.
JOB|5|23|Бо з камінням на полі є в тебе умова, і звір польовий примирився з тобою.
JOB|5|24|І довідаєшся, що намет твій спокійний, і переглянеш домівку свою, і не знайдеш у ній недостатку.
JOB|5|25|І довідаєшся, що численне насіння твоє, а нащадки твої як трава на землі!
JOB|5|26|І в дозрілому віці до гробу ти зійдеш, як збіжжя доспіле ввіходить до клуні за часу свого!
JOB|5|27|Отож, дослідили ми це й воно так, послухай цього, й зрозумій собі все!
JOB|6|1|А Йов відповів та й сказав:
JOB|6|2|Коли б смуток мій вірно був зважений, а з ним разом нещастя моє підняли на вазі,
JOB|6|3|то тепер воно тяжче було б від морського піску, тому нерозважне слова мої кажуть!...
JOB|6|4|Бо в мені Всемогутнього стріли, і їхня отрута п'є духа мого, страхи Божі шикуються в бій проти мене...
JOB|6|5|Чи дикий осел над травою реве? Хіба реве віл, коли ясла повні?
JOB|6|6|Чи без соли їдять несмачне, чи є смак у білкові яйця?
JOB|6|7|Чого не хотіла торкнутись душа моя, все те стало мені за поживу в хворобі...
JOB|6|8|О, коли б же збулося прохання моє, а моє сподівання дав Бог!
JOB|6|9|О, коли б зволив Бог розчавити мене, простягнув Свою руку й мене поламав,
JOB|6|10|то була б ще потіха мені, і скакав би я в немилосердному болі, бо я не зрікався слів Святого!...
JOB|6|11|Яка сила моя, що надію я матиму? І який мій кінець, щоб продовжити життя моє це?
JOB|6|12|Чи сила камінна то сила моя? Чи тіло моє мідяне?
JOB|6|13|Чи не поміч для мене в мені, чи спасіння від мене відсунене?
JOB|6|14|Для того, хто гине, товариш то ласка, хоча б опустив того страх Всемогутнього...
JOB|6|15|Брати мої зраджують, мов той потік, мов річище потоків, минають вони,
JOB|6|16|темніші від льоду вони, в них ховається сніг.
JOB|6|17|Коли сонце їх гріє, вони висихають, у теплі гинуть з місця свого.
JOB|6|18|Каравани дорогу свою відхиляють, уходять в пустиню й щезають.
JOB|6|19|Каравани з Теми поглядають, походи з Шеви покладають надії на них.
JOB|6|20|І засоромилися, що вони сподівались; до нього прийшли та й збентежились.
JOB|6|21|Так і ви тепер стали ніщо, побачили страх і злякались!
JOB|6|22|Чи я говорив коли: Дайте мені, а з маєтку свого дайте підкуп за мене,
JOB|6|23|і врятуйте мене з руки ворога, і з рук гнобителевих мене викупіть?
JOB|6|24|Навчіть ви мене і я буду мовчати, а в чім я невмисне згрішив розтлумачте мені...
JOB|6|25|Які гострі слова справедливі, та що то доводить догана від вас?
JOB|6|26|Чи ви думаєте докоряти словами? Бо на вітер слова одчайдушного,
JOB|6|27|і на сироту нападаєте ви, і копаєте яму для друга свого!...
JOB|6|28|Та звольте поглянути на мене тепер, а я не скажу перед вами неправди.
JOB|6|29|Верніться ж, хай кривди не буде, і верніться, ще в тім моя правда!
JOB|6|30|Хіба в мене на язиці є неправда? чи ж не маю смаку, щоб розпізнати нещастя?
JOB|7|1|Хіба чоловік на землі не на службі військовій? І його дні як дні наймита!...
JOB|7|2|Як раб, спрагнений тіні, і як наймит чекає заплати за працю свою,
JOB|7|3|так місяці марности дано в спадок мені, та ночі терпіння мені відлічили...
JOB|7|4|Коли я кладусь, то кажу: Коли встану? І тягнеться вечір, і перевертання із боку на бік їм до ранку...
JOB|7|5|Зодяглось моє тіло червою та струпами в поросі, шкіра моя затверділа й бридка...
JOB|7|6|А дні мої стали швидчіші за ткацького човника, і в марнотній надії минають вони...
JOB|7|7|Пам'ятай, що життя моє вітер, моє око вже більш не побачить добра...
JOB|7|8|Не побачить мене око того, хто бачив мене, Твої очі поглянуть на мене та немає мене...
JOB|7|9|Як хмара зникає й проходить, так хто сходить в шеол, не виходить,
JOB|7|10|не вертається вже той до дому свого, та й його не пізнає вже місце його...
JOB|7|11|Тож не стримаю я своїх уст, говоритиму в утиску духа свого, нарікати я буду в гіркоті своєї душі:
JOB|7|12|Чи я море чи морська потвора, що Ти надо мною сторожу поставив?
JOB|7|13|Коли я кажу: Нехай постіль потішить мене, хай думки мої ложе моє забере,
JOB|7|14|то Ти снами лякаєш мене, і видіннями страшиш мене...
JOB|7|15|І душа моя прагне задушення, смерти хочуть мої кості.
JOB|7|16|Я обридив життям... Не повіки ж я житиму!... Відпусти ж Ти мене, бо марнота оці мої дні!...
JOB|7|17|Що таке чоловік, що його Ти підносиш, що серце Своє прикладаєш до нього?
JOB|7|18|Ти щоранку за ним назираєш, щохвилі його Ти досліджуєш...
JOB|7|19|Як довго від мене ще Ти не відвернешся, не пустиш мене проковтнути хоч слину свою?
JOB|7|20|Я згрішив... Що ж я маю робити, о Стороже людський? Чому Ти поклав мене ціллю для Себе, і я стався собі тягарем?
JOB|7|21|І чому Ти не простиш мойого гріха, і не відкинеш провини моєї? А тепер я до пороху ляжу, і Ти будеш шукати мене, та немає мене...
JOB|8|1|І заговорив шух'янин Білдад та й сказав:
JOB|8|2|Аж доки ти будеш таке теревенити? І доки слова твоїх уст будуть вітром бурхливим?
JOB|8|3|Чи Бог скривлює суд, і хіба Всемогутній викривлює правду?
JOB|8|4|Якщо твої діти згрішили Йому, то Він їх віддав в руку їх беззаконня!
JOB|8|5|Якщо ти звертатися будеш до Бога, і будеш благати Всемогутнього,
JOB|8|6|якщо чистий ти та безневинний, то тепер Він тобі Свою милість пробудить, і наповнить оселю твою справедливістю,
JOB|8|7|і хоч твій початок нужденний, але твій кінець буде вельми великий!
JOB|8|8|Поспитай в покоління давнішого, і міцно збагни батьків їхніх,
JOB|8|9|бо ми ж учорашні, й нічого не знаєм, бо тінь наші дні на землі,
JOB|8|10|отож вони навчать тебе, тобі скажуть, і з серця свойого слова подадуть:
JOB|8|11|Чи папірус росте без болота? Чи росте очерет без води?
JOB|8|12|Він іще в доспіванні своїм, не зривається, але сохне раніш за всіляку траву:
JOB|8|13|отакі то дороги всіх тих, хто забуває про Бога! І згине надія безбожного,
JOB|8|14|бо його сподівання як те павутиння, і як дім павуків його певність...
JOB|8|15|На свій дім опирається, та не встоїть, тримається міцно за нього, й не вдержиться він...
JOB|8|16|Він зеленіє на сонці, й галузки його випинаються понад садка його,
JOB|8|17|на купі каміння сплелося коріння його, воно між каміння вросло:
JOB|8|18|Якщо вирвуть його з його місця, то зречеться його: тебе я не бачило!...
JOB|8|19|Така радість дороги його, а з пороху інші ростуть.
JOB|8|20|Тож невинного Бог не цурається, і не буде тримати за руку злочинців,
JOB|8|21|аж наповнить уста твої сміхом, а губи твої криком радости...
JOB|8|22|Твої ненависники в сором зодягнуться, і намету безбожних не буде!
JOB|9|1|А Йов відповів та й сказав:
JOB|9|2|Справді пізнав я, що так... Та як оправдатись людині земній перед Богом?
JOB|9|3|Якщо вона схоче на прю стати з Ним, Він відповіді їй не дасть ні на одне із тисячі скаржень...
JOB|9|4|Він мудрого серця й могутньої сили; хто був проти Нього упертий і цілим зостався?
JOB|9|5|Він гори зриває, й не знають вони, що в гніві Своїм Він їх перевернув.
JOB|9|6|Він землю трясе з її місця, і стовпи її трусяться.
JOB|9|7|Він сонцеві скаже, й не сходить воно, і Він запечатує зорі.
JOB|9|8|Розтягує небо Він Сам, і ходить по морських висотах,
JOB|9|9|Він Воза створив, Оріона та Волосожара, та зорі південні.
JOB|9|10|Він чинить велике та недослідиме, предивне, якому немає числа!...
JOB|9|11|Ось Він надо мною проходить, та я не побачу, і Він перейде, а я не приглянусь до Нього...
JOB|9|12|Ось Він схопить кого, хто заверне Його, хто скаже Йому: що Ти робиш?
JOB|9|13|Бог гніву Свойого не спинить, під Ним гнуться Рагавові помічники,
JOB|9|14|що ж тоді відповім я Йому? Які я слова підберу проти Нього,
JOB|9|15|я, який коли б був справедливий, то не відповідав би, я, що благаю свойого Суддю?
JOB|9|16|Коли б я взивав, а Він мені відповідь дав, не повірю, що вчув би мій голос,
JOB|9|17|Він, що бурею може розтерти мене та помножити рани мої безневинно...
JOB|9|18|Не дає Він мені й звести духа мого, бо мене насичає гіркотою.
JOB|9|19|Коли ходить про силу, то Він Всемогутній, коли ж ходить про суд, хто посвідчить мені?
JOB|9|20|Якщо б справедливим я був, то осудять мене мої уста, якщо я безневинний, то вчинять мене винуватим...
JOB|9|21|Я невинний, проте своєї душі я не знаю, і не радий життям своїм я...
JOB|9|22|Це одне, а тому я кажу: невинного як і лукавого Він вигубляє...
JOB|9|23|Якщо нагло бич смерть заподіює, Він з проби невинних сміється...
JOB|9|24|У руку безбожного дана земля, та Він лиця суддів її закриває... Як не Він, тоді хто?
JOB|9|25|А дні мої стали швидкіші, як той скороход, повтікали, не бачили доброго,
JOB|9|26|проминули, немов ті човни очеретяні, мов орел, що несеться на здобич...
JOB|9|27|Якщо я скажу: Хай забуду своє нарікання, хай зміню я обличчя своє й підбадьорюся,
JOB|9|28|то боюся всіх смутків своїх, і я знаю, що Ти не очистиш мене...
JOB|9|29|Все одно буду я винуватий, то нащо надармо я мучитися буду?
JOB|9|30|Коли б я умився сніговою водою, і почистив би лугом долоні свої,
JOB|9|31|то й тоді Ти до гробу опустиш мене, і учинить бридким мене одіж моя...
JOB|9|32|Бо Він не людина, як я, й Йому відповіді я не дам, і не підемо разом на суд,
JOB|9|33|поміж нами нема посередника, що поклав би на нас на обох свою руку...
JOB|9|34|Нехай забере Він від мене Свойого бича, Його ж страх хай мене не жахає,
JOB|9|35|тоді буду казати, й не буду боятись Його, бо я не такий сам з собою!...
JOB|10|1|Життя моє стало бридке для моєї душі... Нехай нарікання своє я на себе пущу, нехай говорю я в гіркоті своєї душі!
JOB|10|2|Скажу Богові я: Не осуджуй мене! Повідом же мене, чого став Ти зо мною на прю?
JOB|10|3|Чи це добре Тобі, що Ти гнобиш мене, що погорджуєш творивом рук Своїх, а раду безбожних освітлюєш?
JOB|10|4|Хіба маєш Ти очі тілесні? Чи Ти бачиш так само, як бачить людина людину?
JOB|10|5|Хіба Твої дні як дні людські, чи літа Твої як дні мужа,
JOB|10|6|що шукаєш провини моєї й вивідуєш гріх мій,
JOB|10|7|хоч відаєш Ти, що я не беззаконник, та нема, хто б мене врятував від Твоєї руки?
JOB|10|8|Твої руки створили мене і вчинили мене, потім Ти обернувся і губиш мене...
JOB|10|9|Пам'ятай, що мов глину мене обробив Ти, і в порох мене обертаєш.
JOB|10|10|Чи не ллєш мене, мов молоко, і не згустив Ти мене, мов на сир?
JOB|10|11|Ти шкірою й тілом мене зодягаєш, і сплів Ти мене із костей та із жил.
JOB|10|12|Життя й милість подав Ти мені, а опіка Твоя стерегла мого духа.
JOB|10|13|А оце заховав Ти у серці Своєму, я знаю, що є воно в Тебе:
JOB|10|14|якщо я грішу, Ти мене стережеш, та з провини моєї мене не очищуєш...
JOB|10|15|Якщо я провинюся, то горе мені! А якщо я невинний, не смію підняти свою голову, ситий стидом та напоєний горем своїм!...
JOB|10|16|А коли піднесеться вона, то Ти ловиш мене, як той лев, і знову предивно зо мною поводишся:
JOB|10|17|поновлюєш свідків Своїх проти мене, помножуєш гнів Свій на мене, військо за військом на мене Ти шлеш...
JOB|10|18|І нащо з утроби Ти вивів мене? Я був би помер, і жоднісіньке око мене не побачило б,
JOB|10|19|як нібито не існував був би я, перейшов би з утроби до гробу...
JOB|10|20|Отож, дні мої нечисленні, перестань же, й від мене вступись, і нехай не турбуюся я бодай трохи,
JOB|10|21|поки я не піду й не вернуся! до краю темноти та смертної тіні,
JOB|10|22|до темного краю, як морок, до тьмяного краю, в якому порядків нема, і де світло, як темрява...
JOB|11|1|І заговорив нааматянин Цофар та й сказав:
JOB|11|2|Чи має зостатись без відповіді безліч слів? І хіба язиката людина невинною буде?
JOB|11|3|Чи мужі замовчать твої теревені, й не буде кому засоромити тебе?
JOB|11|4|Ось говориш ти: Чисте моє міркування, і я чистий в очах Твоїх, Боже!
JOB|11|5|О, коли б говорити став Бог, і відкрив Свої уста до тебе,
JOB|11|6|і представив тобі таємниці премудрости, бо вони як ті чуда роздумування! І знай, вимагає Бог менше від тебе, ніж провини твої того варті!
JOB|11|7|Чи ти Божу глибінь дослідиш, чи знаєш ти аж до кінця Всемогутнього?
JOB|11|8|Вона вища від неба, що зможеш зробити? І глибша вона за шеол, як пізнаєш її?
JOB|11|9|Її міра довша за землю, і ширша за море вона!
JOB|11|10|Якщо Він перейде й замкне щось, і згромадить, то хто заборонить Йому?
JOB|11|11|Бо Він знає нікчемності людські та бачить насилля, і Він не догляне?
JOB|11|12|Тож людина порожня мудрішає, хоч народжується, як те дике осля!
JOB|11|13|Якщо ти зміцниш своє серце, і свої руки до Нього простягнеш,
JOB|11|14|якщо є беззаконня в руці твоїй, то прожени ти його, і кривда в наметах твоїх нехай не пробуває,
JOB|11|15|тож тоді ти підіймеш обличчя невинне своє, і будеш міцний, і не будеш боятись!
JOB|11|16|Бо забудеш страждання, про них будеш згадувати, як про воду, яка пропливла...
JOB|11|17|Від півдня повстане життя, а темрява буде, як ранок.
JOB|11|18|І будеш ти певний, бо маєш надію, і викопаєш собі яму та й будеш безпечно лежати,
JOB|11|19|і будеш лежати, й ніхто не сполошить, і багато-хто будуть підлещуватися до обличчя твого...
JOB|11|20|А очі безбожних минуться, і згине притулок у них, а їхня надія то стогін душі!
JOB|12|1|А Йов відповів та й сказав:
JOB|12|2|Справді, то ж ви тільки люди, і мудрість із вами помре!...
JOB|12|3|Таж і я маю розум, як ви, я не нижчий від вас! І в кого немає такого, як це?
JOB|12|4|Посміховищем став я для друга свого, я, що кликав до Бога, і Він мені відповідав, посміховищем став справедливий, невинний...
JOB|12|5|Нещасливцю погорда, на думку спокійного, приготовлена для спотикання ноги!
JOB|12|6|Спокійні намети грабіжників, і безпечність у тих, хто Бога гнівить, у того, хто ніби то Бога провадить рукою своєю.
JOB|12|7|Але запитай хоч худобу і навчить тебе, і птаство небесне й тобі розповість.
JOB|12|8|Або говори до землі й вона вивчить тебе, і розкажуть тобі риби морські.
JOB|12|9|Хто б із цього всього не пізнав, що Господня рука це вчинила?
JOB|12|10|Що в Нього в руці душа всього живого й дух кожного людського тіла?
JOB|12|11|Чи ж не ухо слова розбирає, піднебіння ж смакує для себе поживу?
JOB|12|12|Мудрість у старших, бо довгість днів розум.
JOB|12|13|Мудрість та сила у Нього, Його рада та розум.
JOB|12|14|Ось Він зруйнує й не буде воно відбудоване, замкне чоловіка й не буде він випущений.
JOB|12|15|Ось Він стримає води і висохнуть, Він їх пустить то землю вони перевернуть.
JOB|12|16|В Нього сила та задум, у Нього заблуджений і той, хто призводить до блуду.
JOB|12|17|Він уводить у помилку радників, і обезумлює суддів,
JOB|12|18|Він розв'язує пута царів і приперізує пояса на їхні стегна.
JOB|12|19|Він провадить священиків босо, і потужних повалює,
JOB|12|20|Він надійним уста відіймає й забирає від старших розумність.
JOB|12|21|На достойників ллє Він погорду, а пояса можним ослаблює.
JOB|12|22|Відкриває Він речі глибокі із темряви, а темне провадить на світло.
JOB|12|23|Він робить народи потужними й знову їх нищить, Він народи поширює, й потім виводить в неволю.
JOB|12|24|Відіймає Він розум в народніх голів на землі та блукати їх змушує по бездорожній пустелі,
JOB|12|25|вони ходять навпомацки в темряві темній, і Він упроваджує їх в блуканину, мов п'яного!
JOB|13|1|Ось усе оце бачило око моє, чуло ухо моє, та й усе зауважило...
JOB|13|2|Як знаєте ви знаю й я, я не нижчий від вас,
JOB|13|3|і я говоритиму до Всемогутнього, і переконувати хочу Бога!
JOB|13|4|Та неправду куєте тут ви, лікарі непутящі ви всі!
JOB|13|5|О, коли б ви насправді мовчали, то вам це за мудрість було б!...
JOB|13|6|Послухайте но переконань моїх: і вислухайте заперечення уст моїх.
JOB|13|7|Чи будете ви говорити неправду про Бога, чи будете ви говорити оману про Нього?
JOB|13|8|Чи будете ви уважати на Нього? Чи за Бога на прю постаєте?
JOB|13|9|Чи добре, що вас Він дослідить? Чи як з людини сміються, так будете ви насміхатися з Нього?
JOB|13|10|Насправді Він вас покарає, якщо будете ви потурати таємно особі!
JOB|13|11|Чи ж велич Його не настрашує вас, і не нападає на вас Його страх?
JOB|13|12|Ваші нагадування це прислів'я із попелу, ваші башти це глиняні башти!
JOB|13|13|Мовчіть передо мною, а я говоритиму, і нехай щобудь прийде на мене!
JOB|13|14|Нащо дертиму я своє тіло зубами своїми, а душу свою покладу в свою руку?
JOB|13|15|Ось Він мене вб'є, і я надії не матиму, але перед обличчям Його про дороги свої сперечатися буду!
JOB|13|16|І це мені буде спасінням, бо перед обличчя Його не підійде безбожний.
JOB|13|17|Направду послухайте слова мого, а моє це освідчення в ваших ушах нехай буде.
JOB|13|18|Ось я суд спорядив, бо я справедливий, те знаю!
JOB|13|19|Хто той, що буде зо мною провадити прю? Бо тепер я замовк би й помер би...
JOB|13|20|Тільки двох цих речей не роби Ти зо мною, тоді від обличчя Твого я не буду ховатись:
JOB|13|21|віддали Свою руку від мене, а Твій страх хай мене не жахає!...
JOB|13|22|Тоді клич, а я відповідатиму, або я говоритиму, Ти ж мені відповідь дай!
JOB|13|23|Скільки в мене провин та гріхів? Покажи Ти мені мій переступ та гріх мій!
JOB|13|24|Чому Ти ховаєш обличчя Своє і вважаєш мене Собі ворогом?
JOB|13|25|Чи Ти будеш страхати завіяний вітром листок? Чи Ти соломину суху будеш гнати?
JOB|13|26|Бо Ти пишеш на мене гіркоти й провини мого молодечого віку даєш на спадок мені,
JOB|13|27|і в кайдани заковуєш ноги мої, і всі дороги мої стережеш, назирці ходиш за мною,
JOB|13|28|і він розпадається, мов та трухлявина, немов та одежа, що міль її з'їла!...
JOB|14|1|Людина, що від жінки народжена, короткоденна та повна печалями:
JOB|14|2|вона виходить, як квітка й зів'яне, і втікає, мов тінь, і не зостається...
JOB|14|3|І на такого Ти очі Свої відкриваєш, і водиш на суд із Собою його!
JOB|14|4|Хто чистого вивести може з нечистого? Ані один!
JOB|14|5|Якщо визначені його дні, число його місяців в Тебе, якщо Ти призначив для нього мету, що її не перейде,
JOB|14|6|відвернися від нього і він заспокоїться, і буде він тішитися своїм днем, як той наймит...
JOB|14|7|Бо дерево має надію: якщо буде стяте, то силу отримає знову, і парост його не загине;
JOB|14|8|якщо постаріє в землі його корінь і в поросі вмре його пень,
JOB|14|9|то від водного запаху знов зацвіте, і пустить галуззя, немов саджанець!
JOB|14|10|А помре чоловік і зникає, а сконає людина то де ж вона є?...
JOB|14|11|Як вода витікає із озера, а річка спадає та сохне,
JOB|14|12|так і та людина покладеться й не встане, аж до закінчення неба не збудяться люди та не прокинуться зо сну свого...
JOB|14|13|О, якби Ти в шеолі мене заховав, коли б Ти мене приховав, аж поки минеться Твій гнів, коли б час Ти призначив мені, та й про мене згадав!
JOB|14|14|Як помре чоловік, то чи він оживе? Буду мати надію по всі дні свойого життя, аж поки не прийде заміна для мене!
JOB|14|15|Кликав би Ти, то я відповів би Тобі, за чин Своїх рук сумував би,
JOB|14|16|бо кроки мої рахував би тепер, а мойого гріха не стеріг би,
JOB|14|17|провина моя була б запечатана в вузлику, і Ти закрив би моє беззаконня...
JOB|14|18|Але гора справді впаде, а скеля зсувається з місця свого,
JOB|14|19|каміння стирає вода, її злива сполощує порох землі, так надію того Ти губиш...
JOB|14|20|Ти силою схопиш назавжди його, і відходить, Ти міняєш обличчя його й відсилаєш його...
JOB|14|21|Чи сини його славні, того він не знає, чи в прикрому стані того він не відає...
JOB|14|22|Боліє він тільки тоді, коли тіло на ньому, коли в ньому душа тоді тужить..
JOB|15|1|І відповів теманянин Еліфаз та й сказав:
JOB|15|2|Чи відповідатиме мудра людина знанням вітряним, і східнім вітром наповнить утробу свою?
JOB|15|3|Буде виправдуватися тим словом, що не надається, чи тими речами, що пожитку немає від них?
JOB|15|4|Ти страх Божий руйнуєш також, і пустошиш молитву до Бога,
JOB|15|5|бо навчає провина твоя твої уста, і ти вибираєш собі язика хитрунів.
JOB|15|6|Оскаржають тебе твої уста, не я, й твої губи свідкують на тебе:
JOB|15|7|Чи ти народився людиною першою, чи раніше, ніж згір'я, ти створений?
JOB|15|8|Чи ти слухав у Божій таємній нараді, та мудрість для себе забрав?
JOB|15|9|Що ти знаєш, чого б ми не знали? Що ти зрозумів, і не з нами воно?
JOB|15|10|Поміж нами і сивий, отой і старий, старший днями від батька твого.
JOB|15|11|Чи мало для тебе потішення Божі та слово, яке Він сховав у тобі?
JOB|15|12|Чого то підносить тебе твоє серце, й які то знаки твої очі дають,
JOB|15|13|що на Бога звертаєш ти духа свого, і з своїх уст випускаєш подібні слова?
JOB|15|14|Що таке чоловік, щоб оправданим бути, і щоб був справедливим від жінки народжений?
JOB|15|15|Таж Він навіть святим Своїм не довіряє, і не оправдані в очах Його небеса,
JOB|15|16|що ж тоді чоловік той бридкий та зіпсутий, що п'є кривду, як воду?
JOB|15|17|Я тобі розповім, ти послухай мене, а що бачив, то те розкажу,
JOB|15|18|про що мудрі донесли та від батьків своїх не затаїли того,
JOB|15|19|їм самим була дана земля, і не приходив чужий поміж них.
JOB|15|20|Безбожний тремтить по всі дні, а насильникові мало років заховано.
JOB|15|21|Вереск жахів у нього в ушах, серед миру приходить на нього грабіжник.
JOB|15|22|Він не вірить, що вернеться від темноти, й він вичікується для меча.
JOB|15|23|Він мандрує за хлібом, та де він? Знає він, що для нього встановлений день темноти...
JOB|15|24|Страшать його утиск та гноблення, хапають його, немов цар, що готовий до бою,
JOB|15|25|бо руку свою простягав він на Бога, і повставав на Всемогутнього,
JOB|15|26|проти Нього твердою він шиєю бігав, товстими хребтами щитів своїх.
JOB|15|27|Бо закрив він обличчя своє своїм салом, і боки обклав своїм жиром,
JOB|15|28|і сидів у містах поруйнованих, у домах тих, що в них не сидять, що на купи каміння призначені.
JOB|15|29|Він не буде багатий, і не встоїться сила його, і по землі не поширяться їхні маєтки.
JOB|15|30|Не вступиться з темности він, полум'я висушить парост його, й духом уст Його буде він схоплений.
JOB|15|31|Хай не вірить в марноту заблуканий, бо марнотою буде заплата йому,
JOB|15|32|вона виповниться не за днів його, а його верховіття не буде зелене!
JOB|15|33|Поскидає насиллям, немов виноград, недозрілість свою, поронить він квіття своє, як оливка,
JOB|15|34|бо збори безбожних спустошені будуть, а огонь пожере дім хабарника:
JOB|15|35|він злом вагітніє, й породить марноту, й оману готує утроба його...
JOB|16|1|А Йов відповів та й сказав:
JOB|16|2|Чув я такого багато, даремні розрадники всі ви!
JOB|16|3|Чи настане кінець вітряним цим словам? Або що зміцнило тебе, що так відповідаєш?
JOB|16|4|І я говорив би, як ви, якби ви на місці моєму були, я додав би словами на вас, і головою своєю кивав би на вас,
JOB|16|5|устами своїми зміцняв би я вас, і не стримав би рух своїх губ на розраду!
JOB|16|6|Якщо я говоритиму, біль мій не стримається, а якщо перестану, що відійде від мене?
JOB|16|7|Та тепер ось Він змучив мене: Всю громаду мою Ти спустошив,
JOB|16|8|і поморщив мене, і це стало за свідчення, і змарнілість моя проти мене повстала, і очевидьки мені докоряє!
JOB|16|9|Його гнів мене шарпає та ненавидить мене, скрегоче на мене зубами своїми, мій ворог вигострює очі свої проти мене...
JOB|16|10|Вони пащі свої роззявляють на мене, б'ють ганебно по щоках мене, збираються разом на мене:
JOB|16|11|Бог злочинцеві видав мене, і кинув у руки безбожних мене...
JOB|16|12|Спокійний я був, та тремтячим мене Він зробив... І за шию вхопив Він мене й розторощив мене, та й поставив мене Собі ціллю:
JOB|16|13|Його стрільці мене оточили, розриває нирки мої Він не жалівши, мою жовч виливає на землю...
JOB|16|14|Він робить пролім на проломі в мені, Він на мене біжить, як силач...
JOB|16|15|Верету пошив я на шкіру свою та під порох знизив свою голову...
JOB|16|16|Зашарілось обличчя моє від плачу, й на повіках моїх залягла смертна тінь,
JOB|16|17|хоч насильства немає в долонях моїх, і чиста молитва моя!
JOB|16|18|Не прикрий, земле, крови моєї, і хай місця не буде для зойку мого,
JOB|16|19|бо тепер ось на небі мій Свідок, Самовидець мій на висоті...
JOB|16|20|Глузливці мої, мої друзі, моє око до Бога сльозить,
JOB|16|21|і нехай Він дозволить людині змагання із Богом, як між сином людським і ближнім його,
JOB|16|22|бо почислені роки минуть, і піду я дорогою, та й не вернусь...
JOB|17|1|Мій дух заламавсь, мої дні погасають, зостались мені самі гроби!...
JOB|17|2|Дійсно, насмішки зо мною, й моє око в розгірченні їхнім ночує...
JOB|17|3|Поклади, дай заставу за мене Ти Сам, хто ж то той, що умову зо мною заб'є по руках?
JOB|17|4|Бо від розуміння закрив Ти їх серце тому не звеличуєш їх.
JOB|17|5|Він призначує ближніх на поділ, а очі синів його темніють,
JOB|17|6|Він поставив мене за прислів'я в народів, і став я таким, на якого плюють...
JOB|17|7|З безталання потемніло око моє, а всі члени мої як та тінь...
JOB|17|8|Праведники остовпіють на це, і невинний встає на безбожного.
JOB|17|9|І праведний буде держатись дороги своєї, а хто чисторукий побільшиться в силі.
JOB|17|10|Але всі ви повернетеся, і приходьте, та я не знаходжу між вами розумного...
JOB|17|11|Мої дні проминули, порвалися думи мої, мого серця маєток,
JOB|17|12|вони мені ніч обертають на день, наближують світло при темряві!
JOB|17|13|Якщо сподіваюсь, то тільки шеолу, як дому свого, в темноті постелю своє ложе...
JOB|17|14|До гробу я кличу: О батьку ти мій! До черви: Моя мамо та сестро моя!...
JOB|17|15|Де ж тоді та надія моя? А надія моя, хто побачить її?
JOB|17|16|До шеолових засувів зійде вона, коли зійдемо разом до пороху...
JOB|18|1|І заговорив шух'янин Білдад та й сказав:
JOB|18|2|Як довго ви будете пастками класти слова? Розміркуйте, а потім собі поговоримо!
JOB|18|3|Чому пораховані ми, як худоба? Чому в ваших очах ми безумні?
JOB|18|4|О ти, що розшарпуєш душу свою в своїм гніві, чи для тебе земля опустіє, а скеля осунеться з місця свого?
JOB|18|5|Таж світильник безбожних погасне, і не буде світитися іскра огню його:
JOB|18|6|його світло стемніє в наметі, і згасне на ньому світильник його,
JOB|18|7|стануть тісні кроки сили його, і вдарить його власна рада!...
JOB|18|8|Бо він кинений в пастку ногами своїми, і на ґраті він буде ходити:
JOB|18|9|пастка схопить за стопу його, зміцниться сітка на ньому,
JOB|18|10|на нього захований шнур на землі, а пастка на нього на стежці...
JOB|18|11|Страхіття жахають його звідусіль, і женуться за ним по слідах.
JOB|18|12|Його сила голодною буде, а нещастя при боці його приготовлене.
JOB|18|13|Його шкіра поїджена буде хворобою, поїсть члени його первороджений смерти.
JOB|18|14|Відірвана буде безпека його від намету його, а Ти до царя жахів його приведеш...
JOB|18|15|Він перебуває в наметі своєму, який не його, на мешкання його буде кинена сірка.
JOB|18|16|Здолу посохнуть коріння його, а згори його віття зів'яне.
JOB|18|17|Його пам'ять загине з землі, а на вулиці ймення не буде йому.
JOB|18|18|Заженуть його з світла до темряви, і ввесь світ проганяє його.
JOB|18|19|У нього немає в народі нащадка, ні внука, і немає останку в місцях його мешкання.
JOB|18|20|На згадку про день його остовпівали останні, за волосся ж хапались давніші...
JOB|18|21|Ось такі то мешкання неправедного, і це місце того, хто Бога не знає!
JOB|19|1|А Йов відповів та й сказав:
JOB|19|2|Аж доки смутити ви будете душу мою, та душити словами мене?
JOB|19|3|Десять раз це мене ви соромите, гнобити мене не стидаєтесь!...
JOB|19|4|Якщо справді зблудив я, то мій гріх при мені позостане.
JOB|19|5|Чи ви величаєтесь справді над мною, і виказуєте мою ганьбу на мене?
JOB|19|6|Знайте тоді, що Бог скривдив мене, і тенета Свої розточив надо мною!
JOB|19|7|Ось ґвалт! я кричу, та не відповідає ніхто, голошу, та немає суду!...
JOB|19|8|Він дорогу мою оточив і я не перейду, Він поклав на стежки мої темряву!
JOB|19|9|Він стягнув з мене славу мою і вінця зняв мені з голови!
JOB|19|10|Звідусіль Він ламає мене, і я йду, надію мою, як те дерево, вивернув Він...
JOB|19|11|І на мене Свій гнів запалив, і зарахував Він мене до Своїх ворогів:
JOB|19|12|полки Його разом приходять, і торують на мене дорогу свою, і таборують навколо намету мого...
JOB|19|13|Віддалив Він від мене братів моїх, а знайомі мої почужіли для мене,
JOB|19|14|мої ближні відстали, і забули про мене знайомі мої...
JOB|19|15|Мешканці дому мого, і служниці мої за чужого вважають мене, чужаком я став в їхніх очах...
JOB|19|16|Я кличу свойого раба і він відповіді не дає, хоч своїми устами благаю його...
JOB|19|17|Мій дух став бридкий для моєї дружини, а мій запах синам моєї утроби...
JOB|19|18|Навіть діти малі зневажають мене, коли я встаю, то глузують із мене...
JOB|19|19|Мої всі повірники бридяться мною, а кого я кохав обернулись на мене...
JOB|19|20|До шкіри моєї й до тіла мого приліпилися кості мої, ще біля зубів лиш зосталася шкіра моя...
JOB|19|21|Змилуйтеся надо мною, о, змилуйтеся надо мною ви, ближні мої, бо Божа рука доторкнулась мене!...
JOB|19|22|Чого ви мене переслідуєте, немов Бог, і не насичуєтесь моїм тілом?
JOB|19|23|О, коли б записати слова мої, о, коли б були в книжці вони позазначувані,
JOB|19|24|коли б рильцем залізним та оливом в скелі навіки вони були витесані!
JOB|19|25|Та я знаю, що мій Викупитель живий, і останнього дня Він підійме із пороху
JOB|19|26|цю шкіру мою, яка розпадається, і з тіла свойого я Бога побачу,
JOB|19|27|сам я побачу Його, й мої очі побачать, а не очі чужі... Тануть нирки мої в моїм нутрі!...
JOB|19|28|Коли скажете ви: Нащо будемо гнати його, коли корень справи знаходиться в ньому!
JOB|19|29|то побійтесь меча собі ви, бо гнів за провину то меч, щоб ви знали, що є ще Суддя!...
JOB|20|1|І відповів нааматянин Цофар та й сказав:
JOB|20|2|Тому то думки мої відповідати мене навертають, і тому то в мені цей мій поспіх!
JOB|20|3|Соромливу нагану собі я почув, та дух з мого розуму відповідає мені.
JOB|20|4|Чи знаєш ти те, що від вічности, відколи людина на землі була поставлена,
JOB|20|5|то спів несправедливих короткий, а радість безбожного тільки на хвилю?
JOB|20|6|Якщо піднесеться величність його аж до неба, а його голова аж до хмари досягне,
JOB|20|7|проте він загине навіки, немов його гній, хто бачив його, запитає: де він?
JOB|20|8|Немов сон улетить і не знайдуть його, мов видіння нічне, він сполошений буде:
JOB|20|9|його бачило око, та бачити більше не буде, і вже не побачить його його місце...
JOB|20|10|Сини його запобігатимуть ласки в нужденних, а руки його позвертають маєток його...
JOB|20|11|Повні кості його молодечости, та до пороху з ним вона ляже!
JOB|20|12|Якщо в устах його зло солодке, його він таїть під своїм язиком,
JOB|20|13|над ним милосердиться та не пускає його, і тримає його в своїх устах,
JOB|20|14|то цей хліб в його нутрощах зміниться, стане він жовчю зміїною в нутрі його!...
JOB|20|15|Він маєток чужого ковтав, але його виблює: Бог виганяє його із утроби його...
JOB|20|16|Отруту зміїну він ссатиме, гадючий язик його вб'є!
JOB|20|17|Він річкових джерел не побачить, струмків меду та молока.
JOB|20|18|Позвертає він працю чужу, і її не ковтне, як і маєток, набутий з виміни своєї, жувати не буде...
JOB|20|19|Бо він переслідував, кидав убогих, він дім грабував, хоч не ставив його!
JOB|20|20|Бо спокою не знав він у нутрі своїм, і свого наймилішого не збереже.
JOB|20|21|Немає останку з обжирства його, тому нетривале добро його все:
JOB|20|22|за повні достатку його буде тісно йому, рука кожного скривдженого прийде на нього!
JOB|20|23|Хай наповнена буде утроба його, та пошле Він на нього жар гніву Свого, і буде дощити на нього недугами його...
JOB|20|24|Він буде втікати від зброї залізної, та прониже його мідний лук...
JOB|20|25|Він стане меча витягати, і вийде він із тіла, та держак його вийде із жовчі його, і перестрах на нього впаде!
JOB|20|26|При скарбах його всі нещастя заховані, його буде жерти огонь не роздмухуваний, позостале в наметі його буде знищене...
JOB|20|27|Небо відкриє його беззаконня, а земля проти нього повстане,
JOB|20|28|урожай його дому втече, розпливеться в день гніву Його...
JOB|20|29|Оце доля від Бога людині безбожній, і спадщина, обіцяна Богом для неї!
JOB|21|1|А Йов відповів та й сказав:
JOB|21|2|Уважно послухайте слово моє, і нехай буде мені це розрадою вашою!
JOB|21|3|Перетерпіть мені, а я промовлятиму, по промові ж моїй насміхатися будеш.
JOB|21|4|Хіба до людини моє нарікання? Чи не мав би чого стати нетерпеливим мій дух?
JOB|21|5|Оберніться до мене й жахніться, та руку на уста свої покладіть...
JOB|21|6|І якщо я згадаю про це, то жахаюсь, і морозом проймається тіло моє...
JOB|21|7|Чого несправедливі живуть, доживають до віку, й багатством зміцняються?
JOB|21|8|Насіння їх міцно стоїть перед ними, при них, а їхні нащадки на їхніх очах...
JOB|21|9|Доми їхні то спокій від страху, і над ними нема бича Божого.
JOB|21|10|Спинається бик його, і не даремно, зачинає корова його, й не скидає.
JOB|21|11|Вони випускають своїх молодят, як отару, а їх діти вибрикують.
JOB|21|12|Вони голос здіймають при бубні та цитрі, і веселяться при звуку сопілки.
JOB|21|13|Провадять в добрі свої дні, і сходять в спокої в шеол.
JOB|21|14|А до Бога говорять вони: Уступися від нас, ми ж доріг Твоїх знати не хочем!
JOB|21|15|Що таке Всемогутній, що будем служити Йому? І що скористаєм, як будем благати Його?
JOB|21|16|Та не в їхній руці добро їхнє, далека від мене порада безбожних...
JOB|21|17|Як часто світильник безбожним згасає, і приходить на них їх нещастя? Він приділює в гніві Своїм на них пастки!
JOB|21|18|Вони будуть, немов та солома на вітрі, і немов та полова, що буря схопила її!
JOB|21|19|Бог ховає синам його кривду Свою та нехай надолужить самому йому, і він знатиме!
JOB|21|20|Нехай його очі побачать нещастя його, й бодай сам він пив гнів Всемогутнього!
JOB|21|21|Яке бо старання його про родину по ньому, як для нього число його місяців вже перелічене?
JOB|21|22|Чи буде хто Бога навчати знання, Його, що й небесних судитиме?
JOB|21|23|Оцей в повній силі своїй помирає, увесь він спокійний та мирний,
JOB|21|24|діжки його повні були молока, а мізок костей його свіжий.
JOB|21|25|А цей помирає з душею огірченою, і доброго не споживав він,
JOB|21|26|та порохом будуть лежати обоє вони, і черва їх покриє...
JOB|21|27|Тож я знаю думки ваші й задуми, що хочете кривдити ними мене.
JOB|21|28|Бож питаєте ви: Де князів дім, і де намет пробування безбожних?
JOB|21|29|Тож спитайтеся тих, що дорогою йдуть, а їхніх ознак не затаюйте:
JOB|21|30|що буває врятований злий в день загибелі, на день гніву відводиться в захист!
JOB|21|31|Хто йому розповість у лице про дорогу його? А коли наробив, хто йому надолужить?
JOB|21|32|І на кладовище буде проваджений він, і про могилу подбають...
JOB|21|33|Скиби долини солодкі йому, і тягнеться кожна людина за ним, а тим, хто попереду нього, немає числа...
JOB|21|34|І як ви мене потішаєте марністю, коли з ваших відповідей зостається сама тільки фальш?...
JOB|22|1|І заговорив теманянин Еліфаз та й сказав:
JOB|22|2|Чи для Бога людина корисна? Бо мудрий корисний самому собі!
JOB|22|3|Хіба Всемогутній бажає, щоб ти ніби праведним був? І що за користь Йому, як дороги свої ти вважаєш невинними сам?
JOB|22|4|Чи Він буде карати, тебе боячись, і чи піде з тобою на суд?
JOB|22|5|Хіба твоє зло не велике? Таж твоїм беззаконням немає кінця!
JOB|22|6|Таж з братів своїх брав ти заставу даремно, а з нагого одежу стягав!
JOB|22|7|Не поїв ти водою знеможеного, і від голодного стримував хліб...
JOB|22|8|А сильна людина то їй оцей край, і почесний у ньому сидітиме.
JOB|22|9|Ти напорожньо вдів відсилав, і сирітські рамена гнобились,
JOB|22|10|тому пастки тебе оточили, і жахає тебе наглий страх,
JOB|22|11|твоє світло стемніло, нічого не бачиш, і велика вода закриває тебе...
JOB|22|12|Чи ж Бог не високий, як небо? Та на зорі угору поглянь, які стали високі вони!
JOB|22|13|А ти кажеш: Що відає Бог? Чи судитиме Він через млу?
JOB|22|14|Хмари завіса Йому, й Він не бачить, і ходить по крузі небесному.
JOB|22|15|Чи ти будеш триматись дороги відвічної, що нею ступали безбожні,
JOB|22|16|що невчасно були вони згублені, що річка розлита, підвалина їх,
JOB|22|17|що до Бога казали вони: Відступися від нас! та: Що зробить для нас Всемогутній?
JOB|22|18|А Він доми їхні наповнив добром!... Але віддалилась від мене порада безбожних!
JOB|22|19|Справедливі це бачать та тішаться, і насміхається з нього невинний:
JOB|22|20|Справді вигублений наш противник, а останок їх вижер огонь!
JOB|22|21|Заприязнися із Ним, та й май спокій, цим прийде на тебе добро.
JOB|22|22|Закона візьми з Його уст, а слова Його в серце своє поклади.
JOB|22|23|Якщо вернешся до Всемогутнього, будеш збудований, і віддалиш беззаконня з наметів своїх.
JOB|22|24|І викинь до пороху золото, і мов камінь з потоку офірське те золото,
JOB|22|25|і буде тобі Всемогутній за золото та за срібло блискуче тобі!
JOB|22|26|Бо тоді Всемогутнього ти покохаєш і до Бога підіймеш обличчя своє,
JOB|22|27|будеш благати Його й Він почує тебе, і ти обітниці свої надолужиш.
JOB|22|28|А що постановиш, то виповниться те тобі, й на дорогах твоїх буде сяяти світло.
JOB|22|29|Бо знижує Він спину пишного, хто ж смиренний, тому помагає.
JOB|22|30|Рятує Він і небезвинного, і той чистотою твоїх рук урятований буде.
JOB|23|1|А Йов відповів та й сказав:
JOB|23|2|Моя мова й сьогодні гірка, тяжче страждання моє за стогнання мої...
JOB|23|3|О, якби то я знав, де Його я знайду, то прийшов би до місця Його пробування!
JOB|23|4|Я б перед обличчям Його свою справу поклав, а уста свої я наповнив би доводами,
JOB|23|5|розізнав би слова, що мені відповість, і я зрозумів би, що скаже мені.
JOB|23|6|Чи зо мною на прю Він з великою силою стане? О ні, тільки б увагу звернув Він на мене!
JOB|23|7|Справедливий судився б там з Ним, я ж назавжди б звільнивсь від свойого Судді.
JOB|23|8|Та піду я на схід і немає Його, а на захід удамся Його не побачу,
JOB|23|9|на півночі шукаю Його й не вхоплю, збочу на південь і не добачаю...
JOB|23|10|А Він знає дорогу, яка при мені, хай би випробував Він мене, мов те золото, вийду!
JOB|23|11|Трималась нога моя коло стопи Його, дороги Його я держався й не збочив.
JOB|23|12|Я не відступався від заповідей Його губ, над уставу свою я ховав слова уст Його.
JOB|23|13|Але Він при одному, й хто заверне Його? Як чого зажадає душа Його, те Він учинить:
JOB|23|14|бо Він виконає, що про мене призначив, і в Нього багато такого, як це!
JOB|23|15|Тому перед обличчям Його я тремчу, розважаю й жахаюсь Його...
JOB|23|16|А Бог пом'якшив моє серце, і Всемогутній мене настрашив,
JOB|23|17|бо не знищений я від темноти, ані від обличчя свого, що темність закрила його!
JOB|24|1|Для чого часи не заховані від Всемогутнього? Ті ж, що знають Його, Його днів не побачать!
JOB|24|2|Пересовують межі безбожні, стадо грабують вони та пасуть,
JOB|24|3|займають осла в сиротини, беруть у заставу вола від удовиць,
JOB|24|4|вони бідних з дороги спихають, разом мусять ховатися збіджені краю...
JOB|24|5|Тож вони, бідарі, немов дикі осли на пустині, виходять на працю свою, здобичі шукаючи, степ йому хліба дає для дітей...
JOB|24|6|На полі вночі вони жнуть, і збирають собі виноград у безбожного,
JOB|24|7|наго ночують вони, без одежі, і не мають вкриття собі в холоді,
JOB|24|8|мокнуть від зливи гірської, а заслони не маючи, скелю вони обіймають...
JOB|24|9|Сироту відривають від перс, і в заставу беруть від убогого...
JOB|24|10|Ходять наго вони, без вбрання, і голодними носять снопи.
JOB|24|11|Хоч між мурами їхніми роблять оливу, топчуть чавила, та прагнуть вони!
JOB|24|12|Стогнуть люди із міста, і кричить душа вбиваних, а Бог на це зло не звертає уваги...
JOB|24|13|Вони проти світла бунтують, не знають доріг Його, і на стежках Його не сидять.
JOB|24|14|На світанку встає душогуб, замордовує бідного та злидаря, а ніч він проводить, як злодій...
JOB|24|15|А перелюбника око чекає смеркання, говорячи: Не побачить мене жодне око! і заслону кладе на обличчя...
JOB|24|16|Підкопуються під доми в темноті, замикаються вдень, світла не знають вони,
JOB|24|17|бо ранок для них усіх разом то темрява, і знають вони жахи темряви...
JOB|24|18|Такий легкий він на поверхні води, на землі їхня частка проклята, не вернеться він на дорогу садів-виноградів...
JOB|24|19|Як посуха та спека їдять сніжну воду, так шеол поїсть грішників!
JOB|24|20|Забуде його лоно матері, буде жерти черва його, мов солодощі, більше не буде він згадуваний, і безбожник поламаний буде, мов дерево!...
JOB|24|21|Чинить зло для бездітної він, щоб вона не родила, і вдовиці не зробить добра.
JOB|24|22|А міццю своєю він тягне могутніх, коли він встає, то ніхто вже не певний свойого життя!
JOB|24|23|Бог дає йому все на безпеку, і на те він спирається, та очі Його бачать їхні дороги:
JOB|24|24|підіймуться трохи й немає вже їх, бо понижені... Як усе, вони гинуть, і зрізуються, немов та колоскова головка...
JOB|24|25|Якщо ж ні, то хто зробить мене неправдомовцем, а слово моє на марноту оберне?
JOB|25|1|І заговорив шух'янин Білдад та й сказав:
JOB|25|2|Панування та острах у Нього, Який на висотах Своїх чинить мир.
JOB|25|3|Чи війську Його є число? І над ким Його світло не сходить?
JOB|25|4|І як може людина бути праведною перед Богом, і як може бути чистим, від жінки народжений?
JOB|25|5|Таж Йому навіть місяць не світить, і в очах Його й зорі не ясні!
JOB|25|6|Що ж тоді людина ота, червяк, чи син людський хробак?...
JOB|26|1|А Йов відповів та й сказав:
JOB|26|2|Як безсилому ти допоміг, як рамено підпер ти неможному?
JOB|26|3|Що ти радив немудрому, й яку раду подав багатьом?
JOB|26|4|Кому ти слова говорив, і чий дух вийшов з тебе?
JOB|26|5|Рефаїми тремтять під водою й всі її мешканці.
JOB|26|6|Голий шеол перед Ним, і нема покриття Аваддону.
JOB|26|7|Він над порожнечею північ простяг, на нічому Він землю повісив.
JOB|26|8|Він зав'язує воду в Своїх облаках, і не розбивається хмара під ними.
JOB|26|9|Він поставив престола Свого, розтягнув над ним хмару Свою.
JOB|26|10|На поверхні води Він зазначив межу аж до границі між світлом та темрявою.
JOB|26|11|Стовпи неба тремтять та страшаться від гніву Його.
JOB|26|12|Він міццю Своєю вспокоює море, і Своїм розумом нищить Рагава.
JOB|26|13|Своїм Духом Він небо прикрасив, рука Його в ньому створила втікаючого Скорпіона.
JOB|26|14|Таж це все самі кінці дороги Його, бо ми тільки слабке шепотіння чували про Нього, грім потуги ж Його хто його зрозуміє?...
JOB|27|1|І Йов далі вів мову свою та й казав:
JOB|27|2|Як живий Бог, відкинув Він право моє, і душу мою засмутив Всемогутній,
JOB|27|3|і як довго в мені ще душа моя, і дух Божий у ніздрях моїх,
JOB|27|4|неправди уста мої не говоритимуть, а язик мій не скаже омани!
JOB|27|5|Борони мене, Боже, признати вас за справедливих! Доки я не помру, своєї невинности я не відкину від себе,
JOB|27|6|за свою справедливість тримаюся міцно, й її не пущу, моє серце не буде ганьбити ні одного з днів моїх,
JOB|27|7|нехай буде мій ворог немов той безбожник, а хто повстає проти мене як кривдник!
JOB|27|8|Яка ж бо надія лукавому, коли відірве, коли візьме Бог душу його?
JOB|27|9|Чи Бог вислухає його крик, коли прийде на нього нещастя?
JOB|27|10|Чи буде втішатися він Всемогутнім? Буде кликати Бога за кожного часу?
JOB|27|11|Я вас буду навчати про Божую руку, що є у Всемогутнього я не сховаю,
JOB|27|12|таж самі ви це бачили всі, то чого ж нісенітниці плещете?
JOB|27|13|Така доля людини безбожної, це спадщина насильників, що отримають від Всемогутнього:
JOB|27|14|Як розмножаться діти його то хіба для меча, а нащадки його не наситяться хлібом!
JOB|27|15|Позосталих по нім моровиця сховає, і вдовиці його не заплачуть...
JOB|27|16|Якщо накопичить він срібла, немов того пороху, і наготує одежі, як глини,
JOB|27|17|то він наготує, а праведний вдягне, а срібло невинний поділить...
JOB|27|18|Він будує свій дім, як та міль, й як той сторож, що ставить собі куреня,
JOB|27|19|він лягає багатим, та більше не зробить того: свої очі відкриє й немає його...
JOB|27|20|Страхіття досягнуть його, мов вода, вночі буря украде його,
JOB|27|21|східній вітер його понесе і минеться, і бурею схопить його з його місця...
JOB|27|22|Оце все Він кине на нього, і не змилосердиться, і від руки Його мусить той спішно втікати!
JOB|27|23|Своїми долонями сплесне над ним, і свисне над ним з свого місця...
JOB|28|1|Отож, має срібло своє джерело, і є місце для золота, де його чистять,
JOB|28|2|залізо береться із пороху, з каменя мідь виплавляється.
JOB|28|3|Людина кладе для темноти кінця, і докраю досліджує все, і шукає каміння у темряві та в смертній тіні:
JOB|28|4|ламає в копальні далеко від мешканця; забуті ногою людини, висять місця, віддалені від чоловіка.
JOB|28|5|Земля хліб із неї походить, а під нею порито, немов би огнем,
JOB|28|6|місце сапфіру каміння її, й порох золота в ній.
JOB|28|7|Стежка туди не знає її хижий птах, її око орлине не бачило,
JOB|28|8|не ступала по ній молода звірина, не ходив нею лев.
JOB|28|9|Чоловік свою руку по кремінь витягує, гори від кореня перевертає,
JOB|28|10|пробиває у скелях канали, і все дороге бачить око його!
JOB|28|11|Він загачує ріки від виливу, а заховані речі виводить на світло.
JOB|28|12|Та де мудрість знаходиться, і де місце розуму?
JOB|28|13|Людина не знає ціни їй, і вона у країні живих не знаходиться.
JOB|28|14|Безодня говорить: Вона не в мені! і море звіщає: Вона не зо мною!
JOB|28|15|Щирого золота дати за неї не можна, і не важиться срібло ціною за неї.
JOB|28|16|Не важать за неї офірського золота, ні дорогого оніксу й сапфіру.
JOB|28|17|Золото й скло не рівняються в вартості їй, і її не зміняти на посуд із щирого золота.
JOB|28|18|Коралі й кришталь і не згадуються, а набуток премудрости ліпший за перли!
JOB|28|19|Не рівняється їй етіопський топаз, і не важиться золото щире за неї.
JOB|28|20|А мудрість ізвідки проходить, і де місце розуму?
JOB|28|21|Бо вона від очей усього живого захована, і від птаства небесного скрита вона.
JOB|28|22|Аваддон той і смерть промовляють: Ушима своїми ми чули про неї лиш чутку!
JOB|28|23|Тільки Бог розуміє дорогу її, й тільки Він знає місце її!
JOB|28|24|Бо Він аж на кінці землі придивляється, бачить під небом усім.
JOB|28|25|Коли Він чинив вагу вітрові, а воду утворював мірою,
JOB|28|26|коли Він уставу складав для дощу та дороги для блискавки грому,
JOB|28|27|тоді Він побачив її та про неї повів, міцно поставив її та її дослідив!
JOB|28|28|І сказав Він людині тоді: Таж страх Господній це мудрість, а відступ від злого це розум!
JOB|29|1|І Йов далі вів мову свою та й сказав:
JOB|29|2|О, коли б я був той, як за місяців давніх, як за днів тих, коли боронив мене Бог,
JOB|29|3|коли над головою моєю світився світильник Його, і при світлі його я ходив в темноті,
JOB|29|4|як був я за днів тих своєї погожої осени, коли Божа милість була над наметом моїм,
JOB|29|5|коли Всемогутній зо мною ще був, а навколо мене мої діти,
JOB|29|6|коли мої кроки купалися в маслі, а скеля оливні струмки біля мене лила!...
JOB|29|7|Коли я виходив до брами при місті, і ставив на площі сидіння своє,
JOB|29|8|як тільки вбачали мене юнаки то ховались, а старші вставали й стояли,
JOB|29|9|зверхники стримували свою мову та клали долоню на уста свої,
JOB|29|10|ховався тоді голос володарів, а їхній язик приліпав їм був до піднебіння...
JOB|29|11|Бо яке ухо чуло про мене, то звало блаженним мене, і яке око бачило, то свідкувало за мене,
JOB|29|12|бо я рятував бідаря, що про поміч кричав, і сироту та безпомічного.
JOB|29|13|Благословення гинучого на мене приходило, а серце вдовиці чинив я співаючим!
JOB|29|14|Зодягавсь я у праведність, і вона зодягала мене, немов плащ та завій було право моє.
JOB|29|15|Очима я був для сліпого, а кривому ногами я був.
JOB|29|16|Бідарям я був батьком, суперечку ж, якої не знав, я досліджував.
JOB|29|17|Й я торощив злочинцеві щелепи, і виривав із зубів його схоплене.
JOB|29|18|І я говорив: Умру я в своєму гнізді, і свої дні я помножу, немов той пісок:
JOB|29|19|для води був відкритий мій корень, а роса зоставалась на вітці моїй...
JOB|29|20|Моя слава була при мені все нова, і в руці моїй лук мій відновлював силу.
JOB|29|21|Мене слухалися й дожидали, і мовчали на раду мою.
JOB|29|22|По слові моїм уже не говорили, і падала мова моя на них краплями.
JOB|29|23|І чекали мене, як дощу, і уста свої відкривали, немов на весінній той дощик...
JOB|29|24|Коли я, бувало, сміявся до них, то не вірили, та світла обличчя мого не гасили.
JOB|29|25|Вибирав я дорогу для них і сидів на чолі, і пробував, немов цар той у війську, коли тішить засмучених він!
JOB|30|1|А тепер насміхаються з мене молодші від мене літами, ті, що їхніх батьків я бридився б покласти із псами отари моєї...
JOB|30|2|Та й сила рук їхніх для чого бувала мені? Повня сил їх минулась!
JOB|30|3|Самотні були в недостатку та голоді, ссали вони суху землю, зруйновану та опустілу!
JOB|30|4|рвали вони лободу на кущах, ялівцеве ж коріння було їхнім хлібом...
JOB|30|5|Вони були вигнані з-поміж людей, кричали на них, немов на злодіїв,
JOB|30|6|так що вони пробували в яругах долин, по ямах підземних та скелях,
JOB|30|7|ревіли вони між кущами, збирались під терням,
JOB|30|8|сини нерозумного й діти неславного, вони були вигнані з краю!
JOB|30|9|А тепер я став піснею їм, і зробився для них поговором...
JOB|30|10|Вони обридили мене, віддалились від мене, і від мойого обличчя не стримали слини,
JOB|30|11|бо Він розв'язав мого пояса й мучить мене, то й вони ось вуздечку із себе відкинули перед обличчям моїм...
JOB|30|12|По правиці встають жовтодзюбі, ноги мені підставляють, і топчуть на мене дороги нещастя свого...
JOB|30|13|Порили вони мою стежку, хочуть мати користь із мойого життя, немає кому їх затримати,
JOB|30|14|немов через вилім широкий приходять, валяються попід румовищем...
JOB|30|15|Обернулось страхіття на мене, моя слава пронеслась, як вітер, і, як хмара, минулося щастя моє...
JOB|30|16|А тепер розливається в мене душа моя, хапають мене дні нещастя!
JOB|30|17|Вночі мої кості від мене віддовбуються, а жили мої не вспокоюються...
JOB|30|18|З великої Божої сили змінилося тіло моє, і недуга мене оперізує, мов той хітон.
JOB|30|19|Він укинув мене до болота, і став я подібний до пороху й попелу.
JOB|30|20|Я кличу до Тебе, та Ти мені відповіді не даєш, я перед Тобою стою, Ти ж на мене лише придивляєшся...
JOB|30|21|Ти змінився мені на жорстокого, мене Ти женеш силою Своєї руки...
JOB|30|22|На вітер підняв Ти мене, на нього мене посадив, і робиш, щоб я розтопивсь на спустошення!
JOB|30|23|Знаю я: Ти до смерти провадиш мене, і до дому зібрання, якого призначив для всього живого...
JOB|30|24|Хіба не простягає руки потопельник, чи він у нещасті своїм не кричить?
JOB|30|25|Чи ж не плакав я за бідарем? Чи за вбогим душа моя не сумувала?
JOB|30|26|Бо чекав я добра, але лихо прийшло, сподівався я світла, та темнота прийшла...
JOB|30|27|Киплять мої нутрощі й не замовкають, зустріли мене дні нещастя,
JOB|30|28|ходжу почорнілий без сонця, на зборі встаю та кричу...
JOB|30|29|Я став братом шакалам, а струсятам товаришем,
JOB|30|30|моя шкіра зчорніла та й лупиться з мене, від спекоти спалилися кості мої...
JOB|30|31|І стала жалобою арфа моя, а сопілка моя зойком плачливим...
JOB|31|1|Умову я склав був з очима своїми, то як буду дивитись на дівчину?
JOB|31|2|І зверху яка доля від Бога, чи спадщина від Всемогутнього із висот?
JOB|31|3|Хіба не загибіль для кривдника, і хіба не нещастя злочинцям?
JOB|31|4|Хіба ж Він не бачить дороги мої, і не лічить усі мої кроки?
JOB|31|5|Якщо я ходив у марноті, і на оману спішила нога моя,
JOB|31|6|то нехай на вазі справедливости зважить мене, і невинність мою Бог пізнає!
JOB|31|7|Якщо збочує крок мій з дороги, і за очима моїми пішло моє серце, і до рук моїх нечисть приліпла,
JOB|31|8|то нехай сію я, а їсть інший, а рослинність моя нехай вирвана буде з корінням!
JOB|31|9|Якщо моє серце зваблялось до жінки чужої, і причаювався я при дверях мойого товариша,
JOB|31|10|то хай меле для іншого жінка моя, і над нею нехай нахиляються інші!
JOB|31|11|Бо гидота оце, й це провина підсудна,
JOB|31|12|бо огонь це, який буде жерти аж до Аваддону, і вирве з корінням увесь урожай мій!...
JOB|31|13|Якщо я понехтував правом свойого раба чи своєї невільниці в їх суперечці зо мною,
JOB|31|14|то що я зроблю, як підійметься Бог? А коли Він приглянеться, що Йому відповім?
JOB|31|15|Чи ж не Той, Хто мене учинив у нутрі, учинив і його, і Один утворив нас в утробі?
JOB|31|16|Чи бажання убогих я стримував, а очі вдовицям засмучував?
JOB|31|17|Чи я сам поїдав свій шматок, і з нього не їв сирота?
JOB|31|18|Таж від днів молодечих моїх виростав він у мене, як в батька, і від утроби матері моєї я провадив його!
JOB|31|19|Якщо бачив я гинучого без одежі, і вбрання не було в сіромахи,
JOB|31|20|чи ж не благословляли мене його стегна, і руном овечок моїх він не грівся?
JOB|31|21|Якщо на сироту я порушував руку свою, коли бачив у брамі собі допомогу,
JOB|31|22|хай рамено моє відпаде від свойого плеча, а рука моя від суглобу свого нехай буде відламана!
JOB|31|23|Бо острах на мене нещастя від Бога, а перед величчям Його я не можу встояти...
JOB|31|24|Чи я золото клав за надію собі, чи до щирого золота я говорив: Ти, безпеко моя?
JOB|31|25|Чи тішився я, що велике багатство моє, й що рука моя стільки надбала?
JOB|31|26|Коли бачив я сонце, як сяє воно, а місяць велично пливе,
JOB|31|27|то коли б потаємно повабилось серце моє, і цілунки рукою я їм посилав,
JOB|31|28|це так само провина підсудна була б, бо відрікся б я Бога Всевишнього!
JOB|31|29|Чи я тішивсь упадком свойого ненависника, чи порушувавсь я, коли зло спотикало його?
JOB|31|30|Таки ні, не давав я на гріх піднебіння свого, щоб прокляттям жадати душі його.
JOB|31|31|Хіба люди намету мого не казали: Хто покаже такого, хто з м'яса його не наситився?
JOB|31|32|Чужинець на вулиці не ночував, я двері свої відчиняв подорожньому.
JOB|31|33|Чи ховав свої прогріхи я, як людина, щоб у своєму нутрі затаїти провину свою?
JOB|31|34|Бо тоді я боявся б великого натовпу, і сором від родів жахав би мене, я мовчав би, й з дверей не виходив...
JOB|31|35|О, якби мене вислухав хто! Оце підпис моєї руки: Нехай Всемогутній мені відповість, а ось звій, зо скаргою, що його написав мій противник...
JOB|31|36|Чи ж я не носив би його на своєму плечі, не обвинувся б ним, як вінками?
JOB|31|37|Число кроків своїх я представлю йому; мов до князя, наближусь до нього.
JOB|31|38|Якщо проти мене голосить земля моя, й її борозни плачуть із нею,
JOB|31|39|якщо без грошей я їв плоди її, а її власника я стогнати примушував,
JOB|31|40|то замість пшениці хай виросте терен, а замість ячменю кукіль!... Слова Йова скінчилися.
JOB|32|1|І перестали ті троє мужів відповідати Йову, бо він був справедливий в очах своїх.
JOB|32|2|І запалився гнів Елігу, сина Барах'їлового, бузянина, з роду Рамового, на Йова запалився гнів його за те, що той уважав душу свою справедливішою за Бога.
JOB|32|3|Також на трьох приятелів його запалився його гнів за те, що не знайшли вони відповіді, а зробили тільки Йова винним.
JOB|32|4|А Елігу вичікував Йова та їх із словами, бо вони були старші віком за нього.
JOB|32|5|І побачив Елігу, що нема належної відповіді в устах тих трьох людей, і запалився його гнів!
JOB|32|6|І відповів бузянин Елігу, син Барах'їлів, та й сказав: Молодий я літами, ви ж старші, тому то я стримувався та боявся знання своє висловити вам.
JOB|32|7|Я подумав: Хай вік промовляє, і хай розуму вчить многоліття!
JOB|32|8|Справді, дух він у людині, та Всемогутнього подих їх мудрими чинить.
JOB|32|9|Многолітні не завжди розумні, і не все розуміються в праві старі.
JOB|32|10|Тому я кажу: Послухай мене, хай знання своє висловлю й я!
JOB|32|11|Тож слів ваших вичікував я, наставляв свої уші до вашої мудрости, поки справу ви дослідите.
JOB|32|12|І я приглядався до вас, й ось немає між вами, хто б Йову довів, хто б відповідь дав на слова його!
JOB|32|13|Щоб ви не сказали: Ми мудрість знайшли: не людина, а Бог переможе його!
JOB|32|14|Не на мене слова він скеровував, і я не відповім йому мовою вашою.
JOB|32|15|Полякались вони, вже не відповідають, не мають вже слів...
JOB|32|16|Я чекав, що не будуть вони говорити, що спинились, не відповідають уже.
JOB|32|17|Відповім також я свою частку, і висловлю й я свою думку.
JOB|32|18|Бо я повний словами, дух мойого нутра докучає мені...
JOB|32|19|Ось утроба моя, мов вино невідкрите, вона тріскається, як нові бурдюки!
JOB|32|20|Нехай я скажу й буде легше мені, нехай уста відкрию свої й відповім!
JOB|32|21|На особу не буду уваги звертати, не буду підлещуватись до людини,
JOB|32|22|бо не вмію підлещуватись! Коли ж ні, нехай зараз візьме мене мій Творець!
JOB|33|1|Але слухай но, Йове, промови мої, і візьми до ушей всі слова мої.
JOB|33|2|Ось я уста свої відкриваю, в моїх устах говорить язик мій.
JOB|33|3|Простота мого серця слова мої, і висловлять ясно знання мої уста.
JOB|33|4|Дух Божий мене учинив, й оживляє мене Всемогутнього подих.
JOB|33|5|Якщо можеш, то дай мені відповідь, вишикуйсь передо мною, постався!
JOB|33|6|Тож Божий і я, як і ти, з глини витиснений теж і я!
JOB|33|7|Ото страх мій тебе не настрашить, і не буде тяжкою рука моя на тобі.
JOB|33|8|Отож, говорив до моїх ушей ти, і я чув голос слів:
JOB|33|9|Чистий я, без гріха, я невинний, і немає провини в мені!
JOB|33|10|Оце Сам Він причини на мене знаходить, уважає мене Собі ворогом.
JOB|33|11|У кайдани закув мої ноги, усі стежки мої Він стереже...
JOB|33|12|Ось у цьому ти не справедливий! Відповім я тобі, бо більший же Бог за людину!
JOB|33|13|Чого Ти із Ним сперечаєшся, що про всі Свої справи Він відповіді не дає?
JOB|33|14|Бо Бог промовляє і раз, і два рази, та людина не бачить того:
JOB|33|15|у сні, у видінні нічному, коли міцний сон на людей нападає, в дрімотах на ложі,
JOB|33|16|тоді відкриває Він ухо людей, і настрашує їх осторогою,
JOB|33|17|щоб відвести людину від чину її, і Він гордість від мужа ховає,
JOB|33|18|щоб від гробу повстримати душу його, а живая його щоб не впала на ратище.
JOB|33|19|І карається хворістю він на постелі своїй, а в костях його сварка міцна.
JOB|33|20|І жива його бридиться хлібом, а душа його стравою влюбленою.
JOB|33|21|Гине тіло його, аж не видно його, і вистають його кості, що перше не видні були.
JOB|33|22|І до гробу душа його зближується, а живая його до померлих іде.
JOB|33|23|Якщо ж Ангол-заступник при нім, один з тисячі, щоб представити людині її правоту,
JOB|33|24|то Він буде йому милосердний та й скаже: Звільни ти його, щоб до гробу не йшов він, Я викуп знайшов.
JOB|33|25|Тоді відмолодиться тіло його, поверне до днів його юности.
JOB|33|26|Він благатиме Бога, й його Собі Він уподобає, і обличчя його буде бачити з окликом радости, і чоловікові верне його справедливість.
JOB|33|27|Він дивитиметься на людей й говоритиме: Я грішив був і правду кривив, та мені не відплачено.
JOB|33|28|Він викупив душу мою, щоб до гробу не йшла, і буде бачити світло живая моя.
JOB|33|29|Бог робить це все двічі-тричі з людиною,
JOB|33|30|щоб душу її відвернути від гробу, щоб він був освітлений світлом живих.
JOB|33|31|Уважай, Йове, слухай мене, мовчи, а я промовлятиму!
JOB|33|32|Коли маєш слова, то дай мені відповідь, говори, бо бажаю твого оправдання.
JOB|33|33|Якщо ні ти послухай мене; помовчи, й я навчу тебе мудрости!
JOB|34|1|І говорив Елігу та й сказав:
JOB|34|2|Слухайте, мудрі, слова ці мої, ви ж, розважні, почуйте мене!
JOB|34|3|Бо ухо слова випробовує, а піднебіння їжу куштує.
JOB|34|4|Виберім право собі, між собою пізнаймо, що добре.
JOB|34|5|Бо Йов говорив: Я був справедливий, та відкинув Бог право моє.
JOB|34|6|Чи буду неправду казати за право своє? Без вини небезпечна стріла моя...
JOB|34|7|Чи є такий муж, як цей Йов, що п'є глузування, як воду,
JOB|34|8|і товаришує з злочинцями, і ходить з людьми беззаконними?
JOB|34|9|Бо він каже: Нема людині користи, коли її Бог уподобає.
JOB|34|10|Тож вислухайте, ви розумні, мене: Бог далекий від несправедливости, і Всемогутній від кривди!
JOB|34|11|Бо за чином людини Він їй надолужить, і згідно з своєю дорогою знайде людина заплату!
JOB|34|12|Тож поправді, не чинить Бог несправедливого, і Всемогутній не скривлює права.
JOB|34|13|Хто землю довірив Йому, і хто на Нього вселенну поклав?
JOB|34|14|Коли б Він до Себе забрав Своє серце, Свій дух, і Свій подих до Себе забрав,
JOB|34|15|всяке тіло погинуло б вмить, а людина повернулася б на порох!...
JOB|34|16|Коли маєш ти розум, послухай же це, почуй голос оцих моїх слів:
JOB|34|17|Хіба стримувати може ненависник право? І хіба осудити ти зможеш Всеправедного?
JOB|34|18|Хіба можна сказати цареві: Негідний, а вельможним: Безбожний?
JOB|34|19|Таж Він не звертає уваги на зверхників, і не вирізнює можного перед убогим, бо всі вони чин Його рук,
JOB|34|20|за хвилину вони помирають, опівночі... Доторкнеться Він можних і гинуть вони, сильний усунений буде рукою не людською.
JOB|34|21|Бо очі Його на дорогах людини, і Він бачить всі кроки її,
JOB|34|22|немає темноти, немає і темряви, де б злочинці сховались.
JOB|34|23|Бо людині Він не призначає означений час, щоб ходила до Бога на суд.
JOB|34|24|Він сильних ламає без досліду, і ставить на місце їх інших.
JOB|34|25|Бож знає Він їхні діла, оберне вночі і почавлені будуть!
JOB|34|26|Як несправедливих уразить Він їх, на видному місці,
JOB|34|27|за те, що вони відступили від Нього, і не розуміли доріг Його всіх,
JOB|34|28|щоб зойк сіромахи спровадити до Нього, бо Він чує благання пригнічених.
JOB|34|29|Коли Він заспокоїть, то хто винуватити буде? Коли Він закриє лице, хто побачить Його? А це робиться і над народом, і над людиною разом,
JOB|34|30|щоб не панував чоловік нечестивий із тих, що правлять за пастку народові.
JOB|34|31|Бо Богові треба отак говорити: Несу я заслужене, злого робити не буду!
JOB|34|32|Чого я не бачу, навчи Ти мене; коли кривду зробив я, то більше не буду чинити!
JOB|34|33|Чи на думку твою надолужить Він це, бо відкинув ти те? Бо вибереш ти, а не я, а що знаєш, кажи!
JOB|34|34|Мені скажуть розумні та муж мудрий, який мене слухає:
JOB|34|35|Йов говорить немудро, а слова його без розуміння.
JOB|34|36|О, коли б Йов досліджений був аж навіки за відповіді, як злі люди,
JOB|34|37|бо він додає до свойого гріха ще провину, між нами він плеще в долоні та множить на Бога промови свої...
JOB|35|1|І говорив Елігу та й сказав:
JOB|35|2|Чи це полічив ти за право, як кажеш: Моя праведність більша за Божу?
JOB|35|3|Бо ти говорив: Що поможе тобі? Яку користь із цього я матиму більшу, аніж від свойого гріха?
JOB|35|4|Я тобі відповім, а з тобою і ближнім твоїм.
JOB|35|5|Подивися на небо й побач, і на хмари споглянь, вони вищі за тебе.
JOB|35|6|Як ти будеш грішити, що зробиш Йому? А стануть численні провини твої, що ти вчиниш Йому?
JOB|35|7|Коли праведним станеш, що даси ти Йому? Або що Він візьме з твоєї руки?
JOB|35|8|Для людини, як ти, беззаконня твоє, і для людського сина твоя справедливість!...
JOB|35|9|Від безлічі гноблення стогнуть вони, кричать від твердого плеча багатьох...
JOB|35|10|Та не скаже ніхто: Де ж той Бог, що мене Він створив, що вночі дає співи,
JOB|35|11|що нас над худобу земну Він навчає, і над птаство небесне вчиняє нас мудрими?
JOB|35|12|Вони там кричать, але через бундючність злочинців Він відповіді не дає.
JOB|35|13|Тільки марноти не слухає Бог, і Всемогутній не бачить її.
JOB|35|14|Що ж тоді, коли кажеш: Не бачив Його! Та є суд перед Ним, і чекай ти його!
JOB|35|15|А тепер, коли гнів Його не покарав, і не дуже пізнав про глупоту,
JOB|35|16|то намарно Йов уста свої відкриває та множить слова без знання...
JOB|36|1|І далі Елігу казав:
JOB|36|2|Почекай мені трохи, й тобі покажу, бо ще є про Бога слова.
JOB|36|3|Зачну викладати я здалека, і Творцеві своєму віддам справедливість.
JOB|36|4|Бо справді слова мої не неправдиві, я з тобою безвадний в знанні.
JOB|36|5|Таж Бог сильний, і не відкидає нікого, Він міцний в силі серця.
JOB|36|6|Не лишає безбожного Він при житті, але право для бідних дає.
JOB|36|7|Від праведного Він очей Своїх не відвертає, але їх садовить з царями на троні назавжди, і вони підвищаються.
JOB|36|8|А як тільки вони ланцюгами пов'язані, і тримаються в путах біди,
JOB|36|9|то Він їм представляє їх вчинок та їхні провини, що багато їх стало.
JOB|36|10|Відкриває Він ухо їх для остороги, та велить, щоб вернулися від беззаконня.
JOB|36|11|Якщо тільки послухаються, та стануть служити Йому, покінчать вони свої дні у добрі, а роки свої у приємнощах.
JOB|36|12|Коли ж не послухаються, то наскочать на ратище, і покінчать життя без знання.
JOB|36|13|А злосерді кладуть гнів на себе, не кричать, коли в'яже Він їх.
JOB|36|14|У молодості помирає душа їх, а їхня живая поміж блудниками.
JOB|36|15|Він визволяє убогого з горя його, а в переслідуванні відкриває їм ухо.
JOB|36|16|Також і тебе Він би вибавив був із тісноти на широкість, що в ній нема утиску, а те, що на стіл твій поклалося б, повне товщу було б.
JOB|36|17|Та правом безбожного ти переповнений, право ж та суд підпирають людину.
JOB|36|18|Отож лютість нехай не намовить тебе до плескання в долоні, а окуп великий нехай не заверне з дороги тебе.
JOB|36|19|Чи в біді допоможе твій зойк та всі зміцнення сили?
JOB|36|20|Не квапся до ночі тієї, коли вирвані будуть народи із місця свого.
JOB|36|21|Стережись, не звертайся до зла, яке замість біди ти обрав.
JOB|36|22|Отож, Бог найвищий у силі Своїй, хто навчає, як Він?
JOB|36|23|Хто дорогу Його Йому вказувати буде? І хто скаже: Ти кривду зробив?
JOB|36|24|Пам'ятай, щоб звеличувати Його вчинок, про якого виспівують люди,
JOB|36|25|що його бачить всяка людина, чоловік приглядається здалека.
JOB|36|26|Отож, Бог великий та недовідомий, і недослідиме число Його літ!
JOB|36|27|Бо стягає Він краплі води, і дощем вони падають з хмари Його,
JOB|36|28|що хмари спускають його, і спадають дощем на багато людей.
JOB|36|29|Також хто зрозуміє розтягнення хмари, грім намету Його?
JOB|36|30|Отож, розтягає Він світло Своє над Собою і морську глибінь закриває,
JOB|36|31|бо ними Він судить народи, багато поживи дає.
JOB|36|32|Він тримає в руках Своїх блискавку, і керує її проти цілі.
JOB|36|33|Її гуркіт звіщає про неї, і прихід її відчуває й худоба.
JOB|37|1|Отож, і від цього тремтить моє серце і зрушилось з місця свого.
JOB|37|2|Уважливо слухайте гук Його голосу, і грім, що несеться із уст Його,
JOB|37|3|його Він пускає попід усім небом, а світло Своє аж на кінці землі.
JOB|37|4|За Ним грім ричить левом, гримить гуком своєї величности, і його Він не стримує, почується голос Його.
JOB|37|5|Бог предивно гримить Своїм голосом, вчиняє великі діла, яких не розуміємо ми.
JOB|37|6|До снігу говорить Він: Падай на землю! а дощеві та зливі: Будьте сильні!
JOB|37|7|Він руку печатає кожній людині, щоб пізнали всі люди про діло Його.
JOB|37|8|І звір входить у сховище, і живе в своїх лігвищах.
JOB|37|9|Із кімнати південної буря приходить, а з вітру північного холод.
JOB|37|10|Від Божого подиху лід повстає, і водна широкість тужавіє.
JOB|37|11|Також Він обтяжує вільгістю тучу, і світло своє розпорошує хмара,
JOB|37|12|і вона по околицях ходить та блукає за Його проводом, щоб чинити все те, що накаже Він їй на поверхні вселенної,
JOB|37|13|він наводить її чи на кару для краю Свого, чи на милість.
JOB|37|14|Бери, Йове, оце до ушей, уставай і розваж Божі чуда!
JOB|37|15|Чи ти знаєш, що Бог накладає на них, і заяснює світло із хмари Своєї?
JOB|37|16|Чи ти знаєш, як носиться хмара в повітрі, про чуда Того, Який має безвадне знання,
JOB|37|17|ти, що шати твої стають теплі, як стишується земля з полудня?
JOB|37|18|Чи ти розтягав із Ним хмару, міцну, немов дзеркало лите?
JOB|37|19|Навчи нас, що скажем Йому? Через темність ми не впорядкуємо слова.
JOB|37|20|Чи Йому оповісться, що буду казати? Чи зміг хто сказати, що Він знищений буде?
JOB|37|21|І тепер ми не бачимо світла, щоб світило у хмарах, та вітер перейде і вичистить їх.
JOB|37|22|Із півночі приходить воно, немов золото те, та над Богом величність страшна.
JOB|37|23|Всемогутній, Його не знайшли ми, Він могутній у силі, але Він не мучить нікого судом та великою правдою.
JOB|37|24|Тому нехай люди бояться Його, бо на всіх мудросердих не дивиться Він.
JOB|38|1|Тоді відповів Господь Йову із бурі й сказав:
JOB|38|2|Хто то такий, що затемнює раду словами без розуму?
JOB|38|3|Підпережи но ти стегна свої, як мужчина, а Я буду питати тебе, ти ж Мені поясни!
JOB|38|4|Де ти був, коли землю основував Я? Розкажи, якщо маєш знання!
JOB|38|5|Хто основи її положив, чи ти знаєш? Або хто розтягнув по ній шнура?
JOB|38|6|У що підстави її позапущувані, або хто поклав камінь наріжний її,
JOB|38|7|коли разом співали всі зорі поранні та радісний окрик здіймали всі Божі сини?
JOB|38|8|І хто море воротами загородив, як воно виступало, немов би з утроби виходило,
JOB|38|9|коли хмари поклав Я за одіж йому, а імлу за його пелюшки,
JOB|38|10|і призначив йому Я границю Свою та поставив засува й ворота,
JOB|38|11|і сказав: Аж досі ти дійдеш, не далі, і тут ось межа твоїх хвиль гордовитих?
JOB|38|12|Чи за своїх днів ти наказував ранкові? Чи досвітній зорі показав її місце,
JOB|38|13|щоб хапалась за кінці землі та посипались з неї безбожні?
JOB|38|14|Земля змінюється, мов та глина печатки, і стають, немов одіж, вони!
JOB|38|15|І нехай від безбожних їх світло відійметься, а високе рамено зламається!
JOB|38|16|Чи ти сходив коли аж до морських джерел, і чи ти переходжувався дном безодні?
JOB|38|17|Чи для тебе відкриті були брами смерти, і чи бачив ти брами смертельної тіні?
JOB|38|18|Чи широкість землі ти оглянув? Розкажи, якщо знаєш це все!
JOB|38|19|Де та дорога, що світло на ній пробуває? А темрява де її місце,
JOB|38|20|щоб узяти її до границі її, і щоб знати стежки її дому?
JOB|38|21|Знаєш ти, бо тоді народився ж ти був, і велике число твоїх днів!
JOB|38|22|Чи доходив коли ти до схованок снігу, і схованки граду ти бачив,
JOB|38|23|які Я тримаю на час лихоліття, на день бою й війни?
JOB|38|24|Якою дорогою ділиться вітер, розпорошується по землі вітерець?
JOB|38|25|Хто для зливи протоку провів, а для громовиці дорогу,
JOB|38|26|щоб дощити на землю безлюдну, на пустиню, в якій чоловіка нема,
JOB|38|27|щоб пустиню та пущу насичувати, і щоб забезпечити вихід траві?
JOB|38|28|Чи є батько в доща, чи хто краплі роси породив?
JOB|38|29|Із чиєї утроби лід вийшов, а іній небесний хто його породив?
JOB|38|30|Як камінь, тужавіють води, а поверхня безодні ховається.
JOB|38|31|Чи зв'яжеш ти зав'язки Волосожару, чи розв'яжеш віжки в Оріона?
JOB|38|32|Чи виведеш часу свого Зодіяка, чи Воза з синами його попровадиш?
JOB|38|33|Чи ти знаєш устави небес? Чи ти покладеш на землі їхню владу?
JOB|38|34|Чи підіймеш свій голос до хмар, і багато води тебе вкриє?
JOB|38|35|Чи блискавки ти посилаєш, і підуть вони, й тобі скажуть Ось ми?
JOB|38|36|Хто мудрість вкладає людині в нутро? Або хто дає серцеві розум?
JOB|38|37|Хто мудрістю хмари зрахує, і хто може затримати небесні посуди,
JOB|38|38|коли порох зливається в зливки, а кавалки злипаються?
JOB|38|39|Чи здобич левиці ти зловиш, і заспокоїш життя левчуків,
JOB|38|40|як вони по леговищах туляться, на чатах сидять по кущах?
JOB|38|41|Хто готує для крука поживу його, як до Бога кричать його діти, як без їжі блукають вони?
JOB|39|1|Хіба ти пізнав час народження скельних козиць? Хіба ти пильнував час мук породу лані?
JOB|39|2|Чи на місяці лічиш, що сповнитись мусять, і відаєш час їх народження,
JOB|39|3|коли приклякають вони, випускають дітей своїх, і звільняються від болів породу?
JOB|39|4|Набираються сил їхні діти, на полі зростають, відходять і більше до них не вертаються.
JOB|39|5|Хто пустив осла дикого вільним, і хто розв'язав ослу дикому пута,
JOB|39|6|якому призначив Я степ його домом, а місцем його пробування солону пустиню?
JOB|39|7|Він сміється із галасу міста, не чує він крику погонича.
JOB|39|8|Що знаходить по горах, то паша його, і шукає він усього зеленого.
JOB|39|9|Чи захоче служити тобі одноріг? Чи при яслах твоїх ночуватиме він?
JOB|39|10|Чи ти однорога прив'яжеш до його борозни повороззям? Чи буде він боронувати за тобою долини?
JOB|39|11|Чи повіриш йому через те, що має він силу велику, і свою працю на нього попустиш?
JOB|39|12|Чи повіриш йому, що він верне насіння твоє, і збере тобі тік?
JOB|39|13|Крило струсеве радісно б'ється, чи ж крило це й пір'їна лелеки?
JOB|39|14|Бо яйця свої він на землю кладе та в поросі їх вигріває,
JOB|39|15|і забува, що нога може їх розчавити, а звір польовий може їх розтоптати.
JOB|39|16|Він жорстокий відносно дітей своїх, ніби вони не його, а що праця його може бути надаремна, того не боїться,
JOB|39|17|бо Бог учинив, щоб забув він про мудрість, і не наділив його розумом.
JOB|39|18|А за часу надходу стрільців ударяє він крильми повітря, і сміється з коня та з його верхівця!
JOB|39|19|Чи ти силу коневі даси, чи шию його ти зодягнеш у гриву?
JOB|39|20|Чи ти зробиш, що буде скакати він, мов сарана? Величне іржання його страшелезне!
JOB|39|21|Б'є ногою в долині та тішиться силою, іде він насупроти зброї,
JOB|39|22|сміється з страху й не жахається, і не вертається з-перед меча,
JOB|39|23|хоч дзвонить над ним сагайдак, вістря списове та ратище!
JOB|39|24|Він із шаленістю та лютістю землю ковтає, і не вірить, що чути гук рогу.
JOB|39|25|При кожному розі кричить він: І-га! і винюхує здалека бій, грім гетьманів та крик.
JOB|39|26|Чи яструб літає твоєю премудрістю, на південь простягує крила свої?
JOB|39|27|Чи з твойого наказу орел підіймається, і мостить кубло своє на висоті?
JOB|39|28|На скелі замешкує він та ночує, на скельнім вершку та твердині,
JOB|39|29|ізвідти визорює їжу, далеко вдивляються очі його,
JOB|39|30|а його пташенята п'ють кров. Де ж забиті, там він.
JOB|40|1|І говорив Господь Йову й сказав:
JOB|40|2|Чи буде ставати на прю з Всемогутнім огудник? Хто сперечається з Богом, хай на це відповість!
JOB|40|3|І Йов відповів Господеві й сказав:
JOB|40|4|Оце я знікчемнів, що ж маю Тобі відповісти? Я кладу свою руку на уста свої...
JOB|40|5|Я раз говорив був, і вже не скажу, а вдруге і більш не додам!...
JOB|40|6|І відповів Господь Йову із бурі й сказав:
JOB|40|7|Підпережи но ти стегна свої, як мужчина: Я буду питати тебе, ти ж пояснюй Мені!
JOB|40|8|Чи ти хочеш порушити право Моє, винуватити Мене, щоб оправданим бути?
JOB|40|9|Коли маєш рамено, як Бог, і голосом ти загримиш, немов Він,
JOB|40|10|то окрась Ти себе пишнотою й величністю, зодягнися у славу й красу!
JOB|40|11|Розпорош лютість гніву свого, і поглянь на все горде й принизь ти його!
JOB|40|12|Поглянь на все горде й його впокори, поспихай нечестивих на їхньому місці,
JOB|40|13|поховай їх у поросі разом, а їхні обличчя обвий в укритті.
JOB|40|14|Тоді й Я тебе славити буду, як правиця твоя допоможе тобі!
JOB|40|15|А ось бегемот, що його Я створив, як тебе, траву, як худоба велика, він їсть.
JOB|40|16|Ото сила його в його стегнах, його ж міцність у м'язах його живота.
JOB|40|17|Випростовує він, немов кедра, свойого хвоста, жили стегон його посплітались.
JOB|40|18|Його кості немов мідяні оті рури, костомахи його як ті пруття залізні.
JOB|40|19|Голова оце Божих доріг; і тільки Творець його може зблизити до нього меча...
JOB|40|20|Бо гори приносять поживу йому, і там грається вся звірина польова.
JOB|40|21|Під лотосами він вилежується, в укритті очерету й болота.
JOB|40|22|Лотоси тінню своєю вкривають його, тополі поточні його обгортають.
JOB|40|23|Ось підіймається річка, та він не боїться її, він безпечний, хоча б сам Йордан йому в пащу впливав!
JOB|40|24|Хто може схопити його в його очах, гаками ніздрю продіравити?
JOB|41|1|(40-25) Чи левіятана потягнеш гачком, і йому язика стягнеш шнуром?
JOB|41|2|(40-26) Чи очеретину вкладеш йому в ніздря, чи терниною щоку йому продіравиш?
JOB|41|3|(40-27) Чи він буде багато благати тебе, чи буде тобі говорити лагідне?
JOB|41|4|(40-28) Чи складе він умову з тобою, і ти візьмеш його за раба собі вічного?
JOB|41|5|(40-29) Чи ним бавитись будеш, як птахом, і прив'яжеш його для дівчаток своїх?
JOB|41|6|(40-30) Чи ним спільники торгуватимуть, чи поділять його між купців-хананеїв?
JOB|41|7|(40-31) Чи шпильками проколиш ти шкіру його, а острогою риб'ячою його голову?
JOB|41|8|(40-32) Поклади ж свою руку на нього, й згадай про війну, і більше того не чини!
JOB|41|9|(41-1) Тож надія твоя неправдива, на сам вигляд його упадеш.
JOB|41|10|(41-2) Нема смільчака, щоб його він збудив, а хто ж перед обличчям Моїм зможе стати?
JOB|41|11|(41-3) Хто вийде навпроти Мене й буде цілий? Що під небом усім це Моє!
JOB|41|12|(41-4) Не буду мовчати про члени його, про стан його сили й красу його складу.
JOB|41|13|(41-5) Хто відкриє поверхню одежі його? Хто підійде коли до двійних його щелепів?
JOB|41|14|(41-6) Двері обличчя його хто відчинить? Навколо зубів його жах!
JOB|41|15|(41-7) Його спина канали щитів, поєднання їх крем'яная печать.
JOB|41|16|(41-8) Одне до одного доходить, а вітер між ними не пройде.
JOB|41|17|(41-9) Одне до одного притверджені, сполучені, і не відділяться.
JOB|41|18|(41-10) Його чхання засвічує світло, а очі його як повіки зорі світової!
JOB|41|19|(41-11) Бухає полум'я з пащі його, вириваються іскри огненні!
JOB|41|20|(41-12) Із ніздер його валить дим, немов з того горшка, що кипить та біжить.
JOB|41|21|(41-13) Його подих розпалює вугіль, і бухає полум'я з пащі його.
JOB|41|22|(41-14) Сила ночує на шиї його, а страх перед ним утікає.
JOB|41|23|(41-15) М'ясо нутра його міцно тримається, воно в ньому тверде, не хитається.
JOB|41|24|(41-16) Його серце, мов з каменя вилите, і тверде, як те долішнє жорно!
JOB|41|25|(41-17) Як підводиться він, перелякуються силачі, та й ховаються з жаху.
JOB|41|26|(41-18) Той меч, що досягне його, не встоїть, ані спис, ані ратище й панцер.
JOB|41|27|(41-19) За солому залізо вважає, а мідь за гнилу деревину!
JOB|41|28|(41-20) Син лука, стріла, не примусит увтікати його, каміння із пращі для нього зміняється в сіно.
JOB|41|29|(41-21) Булаву уважає він за соломинку, і сміється із посвисту ратища.
JOB|41|30|(41-22) Під ним гостре череп'я, лягає на гостре, немов у болото.
JOB|41|31|(41-23) Чинить він, що кипить глибочінь, мов горня, і обертає море в окріп.
JOB|41|32|(41-24) Стежка світить за ним, а безодня здається йому сивиною.
JOB|41|33|(41-25) Немає подоби йому на землі, він безстрашним створений,
JOB|41|34|(41-26) він бачить усе, що високе, він цар над усім пишним звір'ям!
JOB|42|1|А Йов відповів Господеві й сказав:
JOB|42|2|Я знаю, що можеш Ти все, і не спиняється задум у Тебе!
JOB|42|3|Хто ж то такий, що ховає пораду немудру? Тому я говорив, але не розумів... Це чудніше від мене, й не знаю його:
JOB|42|4|Слухай же ти, а Я буду казати, запитаю тебе, ти ж Мені поясни...
JOB|42|5|Тільки послухом уха я чув був про Тебе, а тепер моє око ось бачить Тебе...
JOB|42|6|Тому я зрікаюсь говореного, і каюсь у поросі й попелі!...
JOB|42|7|І сталося по тому, як Господь промовив ці слова до Йова, сказав Господь теманянину Еліфазові: Запалився Мій гнів на тебе та на двох твоїх приятелів, бо ви не говорили слушного про Мене, як раб Мій Йов.
JOB|42|8|А тепер візьміть собі сім бичків та сім баранів, і йдіть до Мого раба Йова, і принесете цілопалення за себе, а Мій раб Йов помолиться за вас, бо тільки з ним Я буду рахуватися, щоб не вчинити вам злої речі, бо ви не говорили слушного про Мене, як раб Мій Йов.
JOB|42|9|І пішли теманянин Еліфаз, і шух'янин Білдад, та нааматянин Цофар, і зробили, як говорив їм Господь. І споглянув Господь на Йова.
JOB|42|10|І Господь привернув Йова до першого стану, коли він помолився за своїх приятелів. І помножив Господь усе, що Йов мав, удвоє.
JOB|42|11|І поприходили до нього всі брати його, і всі сестри його та всі попередні знайомі його, і їли з ним хліб у його домі. І вони головою хитали над ним, та потішали його за все зле, що Господь був спровадив на нього. І дали вони йому кожен по одній кеситі, і кожен по одній золотій обручці.
JOB|42|12|А Господь поблагословив останок днів Йова більше від початку його, і було в нього чотирнадцять тисяч дрібної худоби, і шість тисяч верблюдів, тисяча пар худоби великої та тисяча ослиць.
JOB|42|13|І було в нього семеро синів та три дочки.
JOB|42|14|І назвав він ім'я першій: Єміма, і ім'я другій: Кеція, а ім'я третій: Керен-Гаппух.
JOB|42|15|І таких вродливих жінок, як Йовові дочки, не знайшлося по всій землі. І дав їм їх батько спадщину поміж їхніми братами.
JOB|42|16|А Йов жив по тому сотню й сорок років, і побачив синів своїх та синів синів своїх, чотири поколінні.
JOB|42|17|І впокоївся Йов старим та насиченим днями.
