2PET|1|1|Simon Petrus servus et apostolus Iesu Christi his qui coaequalem nobis sortiti sunt fidem in iustitia Dei nostri et salvatoris Iesu Christi
2PET|1|2|gratia vobis et pax adimpleatur in cognitione Domini nostri
2PET|1|3|quomodo omnia nobis divinae virtutis suae quae ad vitam et pietatem donata est per cognitionem eius qui vocavit nos propria gloria et virtute
2PET|1|4|per quae maxima et pretiosa nobis promissa donavit ut per haec efficiamini divinae consortes naturae fugientes eius quae in mundo est concupiscentiae corruptionem
2PET|1|5|vos autem curam omnem subinferentes ministrate in fide vestra virtutem in virtute autem scientiam
2PET|1|6|in scientia autem abstinentiam in abstinentia autem patientiam in patientia autem pietatem
2PET|1|7|in pietate autem amorem fraternitatis in amore autem fraternitatis caritatem
2PET|1|8|haec enim vobis cum adsint et superent non vacuos nec sine fructu vos constituent in Domini nostri Iesu Christi cognitione
2PET|1|9|cui enim non praesto sunt haec caecus est et manu temptans oblivionem accipiens purgationis veterum suorum delictorum
2PET|1|10|quapropter fratres magis satagite ut per bona opera certam vestram vocationem et electionem faciatis haec enim facientes non peccabitis aliquando
2PET|1|11|sic enim abundanter ministrabitur vobis introitus in aeternum regnum Domini nostri et salvatoris Iesu Christi
2PET|1|12|propter quod incipiam vos semper commonere de his et quidem scientes et confirmatos in praesenti veritate
2PET|1|13|iustum autem arbitror quamdiu sum in hoc tabernaculo suscitare vos in commonitione
2PET|1|14|certus quod velox est depositio tabernaculi mei secundum quod et Dominus noster Iesus Christus significavit mihi
2PET|1|15|dabo autem operam et frequenter habere vos post obitum meum ut horum memoriam faciatis
2PET|1|16|non enim doctas fabulas secuti notam fecimus vobis Domini nostri Iesu Christi virtutem et praesentiam sed speculatores facti illius magnitudinis
2PET|1|17|accipiens enim a Deo Patre honorem et gloriam voce delapsa ad eum huiuscemodi a magnifica gloria hic est Filius meus dilectus in quo mihi conplacui
2PET|1|18|et hanc vocem nos audivimus de caelo adlatam cum essemus cum ipso in monte sancto
2PET|1|19|et habemus firmiorem propheticum sermonem cui bene facitis adtendentes quasi lucernae lucenti in caliginoso loco donec dies inlucescat et lucifer oriatur in cordibus vestris
2PET|1|20|hoc primum intellegentes quod omnis prophetia scripturae propria interpretatione non fit
2PET|1|21|non enim voluntate humana adlata est aliquando prophetia sed Spiritu Sancto inspirati locuti sunt sancti Dei homines
2PET|2|1|fuerunt vero et pseudoprophetae in populo sicut et in vobis erunt magistri mendaces qui introducent sectas perditionis et eum qui emit eos Dominum negant superducentes sibi celerem perditionem
2PET|2|2|et multi sequentur eorum luxurias per quos via veritatis blasphemabitur
2PET|2|3|et in avaritia fictis verbis de vobis negotiabuntur quibus iudicium iam olim non cessat et perditio eorum non dormitat
2PET|2|4|si enim Deus angelis peccantibus non pepercit sed rudentibus inferni detractos in tartarum tradidit in iudicium cruciatos reservari
2PET|2|5|et originali mundo non pepercit sed octavum Noe iustitiae praeconem custodivit diluvium mundo impiorum inducens
2PET|2|6|et civitates Sodomorum et Gomorraeorum in cinerem redigens eversione damnavit exemplum eorum qui impie acturi sunt ponens
2PET|2|7|et iustum Loth oppressum a nefandorum iniuria conversatione eruit
2PET|2|8|aspectu enim et auditu iustus erat habitans apud eos qui diem de die animam iustam iniquis operibus cruciabant
2PET|2|9|novit Dominus pios de temptatione eripere iniquos vero in diem iudicii cruciandos reservare
2PET|2|10|magis autem eos qui post carnem in concupiscentia inmunditiae ambulant dominationemque contemnunt audaces sibi placentes sectas non metuunt blasphemantes
2PET|2|11|ubi angeli fortitudine et virtute cum sint maiores non portant adversum se execrabile iudicium
2PET|2|12|hii vero velut inrationabilia pecora naturaliter in captionem et in perniciem in his quae ignorant blasphemantes in corruptione sua et peribunt
2PET|2|13|percipientes mercedem iniustitiae voluptatem existimantes diei delicias coinquinationes et maculae deliciis affluentes in conviviis suis luxuriantes vobiscum
2PET|2|14|oculos habentes plenos adulterio et incessabiles delicti pellicentes animas instabiles cor exercitatum avaritiae habentes maledictionis filii
2PET|2|15|derelinquentes rectam viam erraverunt secuti viam Balaam ex Bosor qui mercedem iniquitatis amavit
2PET|2|16|correptionem vero habuit suae vesaniae subiugale mutum in hominis voce loquens prohibuit prophetae insipientiam
2PET|2|17|hii sunt fontes sine aqua et nebulae turbinibus exagitatae quibus caligo tenebrarum reservatur
2PET|2|18|superba enim vanitatis loquentes pellicent in desideriis carnis luxuriae eos qui paululum effugiunt qui in errore conversantur
2PET|2|19|libertatem illis promittentes cum ipsi servi sint corruptionis a quo enim quis superatus est huius et servus est
2PET|2|20|si enim refugientes coinquinationes mundi in cognitione Domini nostri et salvatoris Iesu Christi his rursus inpliciti superantur facta sunt eis posteriora deteriora prioribus
2PET|2|21|melius enim erat illis non cognoscere viam iustitiae quam post agnitionem retrorsum converti ab eo quod illis traditum est sancto mandato
2PET|2|22|contigit enim eis illud veri proverbii canis reversus ad suum vomitum et sus lota in volutabro luti
2PET|3|1|hanc ecce vobis carissimi secundam scribo epistulam in quibus excito vestram in commonitione sinceram mentem
2PET|3|2|ut memores sitis eorum quae praedixi verborum a sanctis prophetis et apostolorum vestrorum praeceptorum Domini et salvatoris
2PET|3|3|hoc primum scientes quod venient in novissimis diebus in deceptione inlusores iuxta proprias concupiscentias ambulantes
2PET|3|4|dicentes ubi est promissio aut adventus eius ex quo enim patres dormierunt omnia sic perseverant ab initio creaturae
2PET|3|5|latet enim eos hoc volentes quod caeli erant prius et terra de aqua et per aquam consistens Dei verbo
2PET|3|6|per quae ille tunc mundus aqua inundatus periit
2PET|3|7|caeli autem qui nunc sunt et terra eodem verbo repositi sunt igni servati in diem iudicii et perditionis impiorum hominum
2PET|3|8|unum vero hoc non lateat vos carissimi quia unus dies apud Dominum sicut mille anni et mille anni sicut dies unus
2PET|3|9|non tardat Dominus promissi sed patienter agit propter vos nolens aliquos perire sed omnes ad paenitentiam reverti
2PET|3|10|adveniet autem dies Domini ut fur in qua caeli magno impetu transient elementa vero calore solventur
2PET|3|11|cum haec igitur omnia dissolvenda sint quales oportet esse vos in sanctis conversationibus et pietatibus
2PET|3|12|expectantes et properantes in adventum Dei diei per quam caeli ardentes solventur et elementa ignis ardore tabescent
2PET|3|13|novos vero caelos et novam terram et promissa ipsius expectamus in quibus iustitia habitat
2PET|3|14|propter quod carissimi haec expectantes satis agite inmaculati et inviolati ei inveniri in pace
2PET|3|15|et Domini nostri longanimitatem salutem arbitramini sicut et carissimus frater noster Paulus secundum datam sibi sapientiam scripsit vobis
2PET|3|16|sicut et in omnibus epistulis loquens in eis de his in quibus sunt quaedam difficilia intellectu quae indocti et instabiles depravant sicut et ceteras scripturas ad suam ipsorum perditionem
2PET|3|17|vos igitur fratres praescientes custodite ne insipientium errore transducti excidatis a propria firmitate
2PET|3|18|crescite vero in gratia et in cognitione Domini nostri et salvatoris Iesu Christi ipsi gloria et nunc et in die aeternitatis amen
