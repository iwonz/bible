EPH|1|1|Paul, an apostle of Christ Jesus by the will of God, To the saints who are in Ephesus, and are faithful in Christ Jesus:
EPH|1|2|Grace to you and peace from God our Father and the Lord Jesus Christ.
EPH|1|3|Blessed be the God and Father of our Lord Jesus Christ, who has blessed us in Christ with every spiritual blessing in the heavenly places,
EPH|1|4|even as he chose us in him before the foundation of the world, that we should be holy and blameless before him. In love
EPH|1|5|he predestined us for adoption through Jesus Christ, according to the purpose of his will,
EPH|1|6|to the praise of his glorious grace, with which he has blessed us in the Beloved.
EPH|1|7|In him we have redemption through his blood, the forgiveness of our trespasses, according to the riches of his grace,
EPH|1|8|which he lavished upon us, in all wisdom and insight
EPH|1|9|making known to us the mystery of his will, according to his purpose, which he set forth in Christ
EPH|1|10|as a plan for the fullness of time, to unite all things in him, things in heaven and things on earth.
EPH|1|11|In him we have obtained an inheritance, having been predestined according to the purpose of him who works all things according to the counsel of his will,
EPH|1|12|so that we who were the first to hope in Christ might be to the praise of his glory.
EPH|1|13|In him you also, when you heard the word of truth, the gospel of your salvation, and believed in him, were sealed with the promised Holy Spirit,
EPH|1|14|who is the guarantee of our inheritance until we acquire possession of it, to the praise of his glory.
EPH|1|15|For this reason, because I have heard of your faith in the Lord Jesus and your love toward all the saints,
EPH|1|16|I do not cease to give thanks for you, remembering you in my prayers,
EPH|1|17|that the God of our Lord Jesus Christ, the Father of glory, may give you a spirit of wisdom and of revelation in the knowledge of him,
EPH|1|18|having the eyes of your hearts enlightened, that you may know what is the hope to which he has called you, what are the riches of his glorious inheritance in the saints,
EPH|1|19|and what is the immeasurable greatness of his power toward us who believe, according to the working of his great might
EPH|1|20|that he worked in Christ when he raised him from the dead and seated him at his right hand in the heavenly places,
EPH|1|21|far above all rule and authority and power and dominion, and above every name that is named, not only in this age but also in the one to come.
EPH|1|22|And he put all things under his feet and gave him as head over all things to the church,
EPH|1|23|which is his body, the fullness of him who fills all in all.
EPH|2|1|And you were dead in the trespasses and sins
EPH|2|2|in which you once walked, following the course of this world, following the prince of the power of the air, the spirit that is now at work in the sons of disobedience-
EPH|2|3|among whom we all once lived in the passions of our flesh, carrying out the desires of the body and the mind, and were by nature children of wrath, like the rest of mankind.
EPH|2|4|But God, being rich in mercy, because of the great love with which he loved us,
EPH|2|5|even when we were dead in our trespasses, made us alive together with Christ- by grace you have been saved-
EPH|2|6|and raised us up with him and seated us with him in the heavenly places in Christ Jesus,
EPH|2|7|so that in the coming ages he might show the immeasurable riches of his grace in kindness toward us in Christ Jesus.
EPH|2|8|For by grace you have been saved through faith. And this is not your own doing; it is the gift of God,
EPH|2|9|not a result of works, so that no one may boast.
EPH|2|10|For we are his workmanship, created in Christ Jesus for good works, which God prepared beforehand, that we should walk in them.
EPH|2|11|Therefore remember that at one time you Gentiles in the flesh, called "the uncircumcision" by what is called the circumcision, which is made in the flesh by hands-
EPH|2|12|remember that you were at that time separated from Christ, alienated from the commonwealth of Israel and strangers to the covenants of promise, having no hope and without God in the world.
EPH|2|13|But now in Christ Jesus you who once were far off have been brought near by the blood of Christ.
EPH|2|14|For he himself is our peace, who has made us both one and has broken down in his flesh the dividing wall of hostility
EPH|2|15|by abolishing the law of commandments and ordinances, that he might create in himself one new man in place of the two, so making peace,
EPH|2|16|and might reconcile us both to God in one body through the cross, thereby killing the hostility.
EPH|2|17|And he came and preached peace to you who were far off and peace to those who were near.
EPH|2|18|For through him we both have access in one Spirit to the Father.
EPH|2|19|So then you are no longer strangers and aliens, but you are fellow citizens with the saints and members of the household of God,
EPH|2|20|built on the foundation of the apostles and prophets, Christ Jesus himself being the cornerstone,
EPH|2|21|in whom the whole structure, being joined together, grows into a holy temple in the Lord.
EPH|2|22|In him you also are being built together into a dwelling place for God by the Spirit.
EPH|3|1|For this reason I, Paul, a prisoner for Christ Jesus on behalf of you Gentiles-
EPH|3|2|assuming that you have heard of the stewardship of God's grace that was given to me for you,
EPH|3|3|how the mystery was made known to me by revelation, as I have written briefly.
EPH|3|4|When you read this, you can perceive my insight into the mystery of Christ,
EPH|3|5|which was not made known to the sons of men in other generations as it has now been revealed to his holy apostles and prophets by the Spirit.
EPH|3|6|This mystery is that the Gentiles are fellow heirs, members of the same body, and partakers of the promise in Christ Jesus through the gospel.
EPH|3|7|Of this gospel I was made a minister according to the gift of God's grace, which was given me by the working of his power.
EPH|3|8|To me, though I am the very least of all the saints, this grace was given, to preach to the Gentiles the unsearchable riches of Christ,
EPH|3|9|and to bring to light for everyone what is the plan of the mystery hidden for ages in God who created all things,
EPH|3|10|so that through the church the manifold wisdom of God might now be made known to the rulers and authorities in the heavenly places.
EPH|3|11|This was according to the eternal purpose that he has realized in Christ Jesus our Lord,
EPH|3|12|in whom we have boldness and access with confidence through our faith in him.
EPH|3|13|So I ask you not to lose heart over what I am suffering for you, which is your glory.
EPH|3|14|For this reason I bow my knees before the Father,
EPH|3|15|from whom every family in heaven and on earth is named,
EPH|3|16|that according to the riches of his glory he may grant you to be strengthened with power through his Spirit in your inner being,
EPH|3|17|so that Christ may dwell in your hearts through faith- that you, being rooted and grounded in love,
EPH|3|18|may have strength to comprehend with all the saints what is the breadth and length and height and depth,
EPH|3|19|and to know the love of Christ that surpasses knowledge, that you may be filled with all the fullness of God.
EPH|3|20|Now to him who is able to do far more abundantly than all that we ask or think, according to the power at work within us,
EPH|3|21|to him be glory in the church and in Christ Jesus throughout all generations, forever and ever. Amen.
EPH|4|1|I therefore, a prisoner for the Lord, urge you to walk in a manner worthy of the calling to which you have been called,
EPH|4|2|with all humility and gentleness, with patience, bearing with one another in love,
EPH|4|3|eager to maintain the unity of the Spirit in the bond of peace.
EPH|4|4|There is one body and one Spirit- just as you were called to the one hope that belongs to your call-
EPH|4|5|one Lord, one faith, one baptism,
EPH|4|6|one God and Father of all, who is over all and through all and in all.
EPH|4|7|But grace was given to each one of us according to the measure of Christ's gift.
EPH|4|8|Therefore it says, "When he ascended on high he led a host of captives, and he gave gifts to men."
EPH|4|9|(In saying, "He ascended," what does it mean but that he had also descended into the lower parts of the earth?
EPH|4|10|He who descended is the one who also ascended far above all the heavens, that he might fill all things.)
EPH|4|11|And he gave the apostles, the prophets, the evangelists, the pastors and teachers,
EPH|4|12|to equip the saints for the work of ministry, for building up the body of Christ,
EPH|4|13|until we all attain to the unity of the faith and of the knowledge of the Son of God, to mature manhood, to the measure of the stature of the fullness of Christ,
EPH|4|14|so that we may no longer be children, tossed to and fro by the waves and carried about by every wind of doctrine, by human cunning, by craftiness in deceitful schemes.
EPH|4|15|Rather, speaking the truth in love, we are to grow up in every way into him who is the head, into Christ,
EPH|4|16|from whom the whole body, joined and held together by every joint with which it is equipped, when each part is working properly, makes the body grow so that it builds itself up in love.
EPH|4|17|Now this I say and testify in the Lord, that you must no longer walk as the Gentiles do, in the futility of their minds.
EPH|4|18|They are darkened in their understanding, alienated from the life of God because of the ignorance that is in them, due to their hardness of heart.
EPH|4|19|They have become callous and have given themselves up to sensuality, greedy to practice every kind of impurity.
EPH|4|20|But that is not the way you learned Christ!-
EPH|4|21|assuming that you have heard about him and were taught in him, as the truth is in Jesus,
EPH|4|22|to put off your old self, which belongs to your former manner of life and is corrupt through deceitful desires,
EPH|4|23|and to be renewed in the spirit of your minds,
EPH|4|24|and to put on the new self, created after the likeness of God in true righteousness and holiness.
EPH|4|25|Therefore, having put away falsehood, let each one of you speak the truth with his neighbor, for we are members one of another.
EPH|4|26|Be angry and do not sin; do not let the sun go down on your anger,
EPH|4|27|and give no opportunity to the devil.
EPH|4|28|Let the thief no longer steal, but rather let him labor, doing honest work with his own hands, so that he may have something to share with anyone in need.
EPH|4|29|Let no corrupting talk come out of your mouths, but only such as is good for building up, as fits the occasion, that it may give grace to those who hear.
EPH|4|30|And do not grieve the Holy Spirit of God, by whom you were sealed for the day of redemption.
EPH|4|31|Let all bitterness and wrath and anger and clamor and slander be put away from you, along with all malice.
EPH|4|32|Be kind to one another, tenderhearted, forgiving one another, as God in Christ forgave you.
EPH|5|1|Therefore be imitators of God, as beloved children.
EPH|5|2|And walk in love, as Christ loved us and gave himself up for us, a fragrant offering and sacrifice to God.
EPH|5|3|But sexual immorality and all impurity or covetousness must not even be named among you, as is proper among saints.
EPH|5|4|Let there be no filthiness nor foolish talk nor crude joking, which are out of place, but instead let there be thanksgiving.
EPH|5|5|For you may be sure of this, that everyone who is sexually immoral or impure, or who is covetous (that is, an idolater), has no inheritance in the kingdom of Christ and God.
EPH|5|6|Let no one deceive you with empty words, for because of these things the wrath of God comes upon the sons of disobedience.
EPH|5|7|Therefore do not associate with them;
EPH|5|8|for at one time you were darkness, but now you are light in the Lord. Walk as children of light
EPH|5|9|(for the fruit of light is found in all that is good and right and true),
EPH|5|10|and try to discern what is pleasing to the Lord.
EPH|5|11|Take no part in the unfruitful works of darkness, but instead expose them.
EPH|5|12|For it is shameful even to speak of the things that they do in secret.
EPH|5|13|But when anything is exposed by the light, it becomes visible,
EPH|5|14|for anything that becomes visible is light. Therefore it says, "Awake, O sleeper, and arise from the dead, and Christ will shine on you."
EPH|5|15|Look carefully then how you walk, not as unwise but as wise,
EPH|5|16|making the best use of the time, because the days are evil.
EPH|5|17|Therefore do not be foolish, but understand what the will of the Lord is.
EPH|5|18|And do not get drunk with wine, for that is debauchery, but be filled with the Spirit,
EPH|5|19|addressing one another in psalms and hymns and spiritual songs, singing and making melody to the Lord with all your heart,
EPH|5|20|giving thanks always and for everything to God the Father in the name of our Lord Jesus Christ,
EPH|5|21|submitting to one another out of reverence for Christ.
EPH|5|22|Wives, submit to your own husbands, as to the Lord.
EPH|5|23|For the husband is the head of the wife even as Christ is the head of the church, his body, and is himself its Savior.
EPH|5|24|Now as the church submits to Christ, so also wives should submit in everything to their husbands.
EPH|5|25|Husbands, love your wives, as Christ loved the church and gave himself up for her,
EPH|5|26|that he might sanctify her, having cleansed her by the washing of water with the word,
EPH|5|27|so that he might present the church to himself in splendor, without spot or wrinkle or any such thing, that she might be holy and without blemish.
EPH|5|28|In the same way husbands should love their wives as their own bodies. He who loves his wife loves himself.
EPH|5|29|For no one ever hated his own flesh, but nourishes and cherishes it, just as Christ does the church,
EPH|5|30|because we are members of his body.
EPH|5|31|"Therefore a man shall leave his father and mother and hold fast to his wife, and the two shall become one flesh."
EPH|5|32|This mystery is profound, and I am saying that it refers to Christ and the church.
EPH|5|33|However, let each one of you love his wife as himself, and let the wife see that she respects her husband.
EPH|6|1|Children, obey your parents in the Lord, for this is right.
EPH|6|2|"Honor your father and mother" (this is the first commandment with a promise),
EPH|6|3|"that it may go well with you and that you may live long in the land."
EPH|6|4|Fathers, do not provoke your children to anger, but bring them up in the discipline and instruction of the Lord.
EPH|6|5|Slaves, obey your earthly masters with fear and trembling, with a sincere heart, as you would Christ,
EPH|6|6|not by the way of eye-service, as people-pleasers, but as servants of Christ, doing the will of God from the heart,
EPH|6|7|rendering service with a good will as to the Lord and not to man,
EPH|6|8|knowing that whatever good anyone does, this he will receive back from the Lord, whether he is a slave or free.
EPH|6|9|Masters, do the same to them, and stop your threatening, knowing that he who is both their Master and yours is in heaven, and that there is no partiality with him.
EPH|6|10|Finally, be strong in the Lord and in the strength of his might.
EPH|6|11|Put on the whole armor of God, that you may be able to stand against the schemes of the devil.
EPH|6|12|For we do not wrestle against flesh and blood, but against the rulers, against the authorities, against the cosmic powers over this present darkness, against the spiritual forces of evil in the heavenly places.
EPH|6|13|Therefore take up the whole armor of God, that you may be able to withstand in the evil day, and having done all, to stand firm.
EPH|6|14|Stand therefore, having fastened on the belt of truth, and having put on the breastplate of righteousness,
EPH|6|15|and, as shoes for your feet, having put on the readiness given by the gospel of peace.
EPH|6|16|In all circumstances take up the shield of faith, with which you can extinguish all the flaming darts of the evil one;
EPH|6|17|and take the helmet of salvation, and the sword of the Spirit, which is the word of God,
EPH|6|18|praying at all times in the Spirit, with all prayer and supplication. To that end keep alert with all perseverance, making supplication for all the saints,
EPH|6|19|and also for me, that words may be given to me in opening my mouth boldly to proclaim the mystery of the gospel,
EPH|6|20|for which I am an ambassador in chains, that I may declare it boldly, as I ought to speak.
EPH|6|21|So that you also may know how I am and what I am doing, Tychicus the beloved brother and faithful minister in the Lord will tell you everything.
EPH|6|22|I have sent him to you for this very purpose, that you may know how we are, and that he may encourage your hearts.
EPH|6|23|Peace be to the brothers, and love with faith, from God the Father and the Lord Jesus Christ.
EPH|6|24|Grace be with all who love our Lord Jesus Christ with love incorruptible.
