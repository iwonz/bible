PHIL|1|1|Paulus et Timotheus servi Iesu Christi omnibus sanctis in Christo Iesu qui sunt Philippis cum episcopis et diaconis
PHIL|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
PHIL|1|3|gratias ago Deo meo in omni memoria vestri
PHIL|1|4|semper in cunctis orationibus meis pro omnibus vobis cum gaudio deprecationem faciens
PHIL|1|5|super communicatione vestra in evangelio a prima die usque nunc
PHIL|1|6|confidens hoc ipsum quia qui coepit in vobis opus bonum perficiet usque in diem Christi Iesu
PHIL|1|7|sicut est mihi iustum hoc sentire pro omnibus vobis eo quod habeam in corde vos et in vinculis meis et in defensione et confirmatione evangelii socios gaudii mei omnes vos esse
PHIL|1|8|testis enim mihi est Deus quomodo cupiam omnes vos in visceribus Christi Iesu
PHIL|1|9|et hoc oro ut caritas vestra magis ac magis abundet in scientia et omni sensu
PHIL|1|10|ut probetis potiora ut sitis sinceres et sine offensa in diem Christi
PHIL|1|11|repleti fructu iustitiae per Christum Iesum in gloriam et laudem Dei
PHIL|1|12|scire autem vos volo fratres quia quae circa me sunt magis ad profectum venerunt evangelii
PHIL|1|13|ita ut vincula mea manifesta fierent in Christo in omni praetorio et in ceteris omnibus
PHIL|1|14|et plures e fratribus in Domino confidentes vinculis meis abundantius audere sine timore verbum Dei loqui
PHIL|1|15|quidam quidem et propter invidiam et contentionem quidam autem et propter bonam voluntatem Christum praedicant
PHIL|1|16|quidam ex caritate scientes quoniam in defensionem evangelii positus sum
PHIL|1|17|quidam autem ex contentione Christum adnuntiant non sincere existimantes pressuram se suscitare vinculis meis
PHIL|1|18|quid enim dum omni modo sive per occasionem sive per veritatem Christus adnuntiatur et in hoc gaudeo sed et gaudebo
PHIL|1|19|scio enim quia hoc mihi proveniet in salutem per vestram orationem et subministrationem Spiritus Iesu Christi
PHIL|1|20|secundum expectationem et spem meam quia in nullo confundar sed in omni fiducia sicut semper et nunc magnificabitur Christus in corpore meo sive per vitam sive per mortem
PHIL|1|21|mihi enim vivere Christus est et mori lucrum
PHIL|1|22|quod si vivere in carne hic mihi fructus operis est et quid eligam ignoro
PHIL|1|23|coartor autem e duobus desiderium habens dissolvi et cum Christo esse multo magis melius
PHIL|1|24|permanere autem in carne magis necessarium est propter vos
PHIL|1|25|et hoc confidens scio quia manebo et permanebo omnibus vobis ad profectum vestrum et gaudium fidei
PHIL|1|26|ut gratulatio vestra abundet in Christo Iesu in me per meum adventum iterum ad vos
PHIL|1|27|tantum digne evangelio Christi conversamini ut sive cum venero et videro vos sive absens audiam de vobis quia stetistis uno spiritu unianimes conlaborantes fide evangelii
PHIL|1|28|et in nullo terreamini ab adversariis quae est illis causa perditionis vobis autem salutis et hoc a Deo
PHIL|1|29|quia vobis donatum est pro Christo non solum ut in eum credatis sed ut etiam pro illo patiamini
PHIL|1|30|eundem certamen habentes qualem et vidistis in me et nunc audistis de me
PHIL|2|1|si qua ergo consolatio in Christo si quod solacium caritatis si qua societas spiritus si quid viscera et miserationes
PHIL|2|2|implete gaudium meum ut idem sapiatis eandem caritatem habentes unianimes id ipsum sentientes
PHIL|2|3|nihil per contentionem neque per inanem gloriam sed in humilitate superiores sibi invicem arbitrantes
PHIL|2|4|non quae sua sunt singuli considerantes sed et ea quae aliorum
PHIL|2|5|hoc enim sentite in vobis quod et in Christo Iesu
PHIL|2|6|qui cum in forma Dei esset non rapinam arbitratus est esse se aequalem Deo
PHIL|2|7|sed semet ipsum exinanivit formam servi accipiens in similitudinem hominum factus et habitu inventus ut homo
PHIL|2|8|humiliavit semet ipsum factus oboediens usque ad mortem mortem autem crucis
PHIL|2|9|propter quod et Deus illum exaltavit et donavit illi nomen super omne nomen
PHIL|2|10|ut in nomine Iesu omne genu flectat caelestium et terrestrium et infernorum
PHIL|2|11|et omnis lingua confiteatur quia Dominus Iesus Christus in gloria est Dei Patris
PHIL|2|12|itaque carissimi mei sicut semper oboedistis non ut in praesentia mei tantum sed multo magis nunc in absentia mea cum metu et tremore vestram salutem operamini
PHIL|2|13|Deus est enim qui operatur in vobis et velle et perficere pro bona voluntate
PHIL|2|14|omnia autem facite sine murmurationibus et haesitationibus
PHIL|2|15|ut sitis sine querella et simplices filii Dei sine reprehensione in medio nationis pravae et perversae inter quos lucetis sicut luminaria in mundo
PHIL|2|16|verbum vitae continentes ad gloriam meam in die Christi quia non in vacuum cucurri neque in vacuum laboravi
PHIL|2|17|sed et si immolor supra sacrificium et obsequium fidei vestrae gaudeo et congratulor omnibus vobis
PHIL|2|18|id ipsum autem et vos gaudete et congratulamini mihi
PHIL|2|19|spero autem in Domino Iesu Timotheum cito me mittere ad vos ut et ego bono animo sim cognitis quae circa vos sunt
PHIL|2|20|neminem enim habeo tam unianimem qui sincera affectione pro vobis sollicitus sit
PHIL|2|21|omnes enim sua quaerunt non quae sunt Christi Iesu
PHIL|2|22|experimentum autem eius cognoscite quoniam sicut patri filius mecum servivit in evangelium
PHIL|2|23|hunc igitur spero me mittere mox ut videro quae circa me sunt
PHIL|2|24|confido autem in Domino quoniam et ipse veniam ad vos cito
PHIL|2|25|necessarium autem existimavi Epafroditum fratrem et cooperatorem et commilitonem meum vestrum autem apostolum et ministrum necessitatis meae mittere ad vos
PHIL|2|26|quoniam quidem omnes vos desiderabat et maestus erat propterea quod audieratis illum infirmatum
PHIL|2|27|nam et infirmatus est usque ad mortem sed Deus misertus est eius non solum autem eius verum etiam et mei ne tristitiam super tristitiam haberem
PHIL|2|28|festinantius ergo misi illum ut viso eo iterum gaudeatis et ego sine tristitia sim
PHIL|2|29|excipite itaque illum cum omni gaudio in Domino et eiusmodi cum honore habetote
PHIL|2|30|quoniam propter opus Christi usque ad mortem accessit tradens animam suam ut impleret id quod ex vobis deerat erga meum obsequium
PHIL|3|1|de cetero fratres mei gaudete in Domino eadem vobis scribere mihi quidem non pigrum vobis autem necessarium
PHIL|3|2|videte canes videte malos operarios videte concisionem
PHIL|3|3|nos enim sumus circumcisio qui spiritu Deo servimus et gloriamur in Christo Iesu et non in carne fiduciam habentes
PHIL|3|4|quamquam ego habeam confidentiam et in carne si quis alius videtur confidere in carne ego magis
PHIL|3|5|circumcisus octava die ex genere Israhel de tribu Beniamin Hebraeus ex Hebraeis secundum legem Pharisaeus
PHIL|3|6|secundum aemulationem persequens ecclesiam Dei secundum iustitiam quae in lege est conversatus sine querella
PHIL|3|7|sed quae mihi fuerunt lucra haec arbitratus sum propter Christum detrimenta
PHIL|3|8|verumtamen existimo omnia detrimentum esse propter eminentem scientiam Iesu Christi Domini mei propter quem omnia detrimentum feci et arbitror ut stercora ut Christum lucri faciam
PHIL|3|9|et inveniar in illo non habens meam iustitiam quae ex lege est sed illam quae ex fide est Christi quae ex Deo est iustitia in fide
PHIL|3|10|ad agnoscendum illum et virtutem resurrectionis eius et societatem passionum illius configuratus morti eius
PHIL|3|11|si quo modo occurram ad resurrectionem quae est ex mortuis
PHIL|3|12|non quod iam acceperim aut iam perfectus sim sequor autem si conprehendam in quo et conprehensus sum a Christo Iesu
PHIL|3|13|fratres ego me non arbitror conprehendisse unum autem quae quidem retro sunt obliviscens ad ea vero quae sunt in priora extendens me
PHIL|3|14|ad destinatum persequor ad bravium supernae vocationis Dei in Christo Iesu
PHIL|3|15|quicumque ergo perfecti hoc sentiamus et si quid aliter sapitis et hoc vobis Deus revelabit
PHIL|3|16|verumtamen ad quod pervenimus ut idem sapiamus et in eadem permaneamus regula
PHIL|3|17|imitatores mei estote fratres et observate eos qui ita ambulant sicut habetis formam nos
PHIL|3|18|multi enim ambulant quos saepe dicebam vobis nunc autem et flens dico inimicos crucis Christi
PHIL|3|19|quorum finis interitus quorum deus venter et gloria in confusione ipsorum qui terrena sapiunt
PHIL|3|20|nostra autem conversatio in caelis est unde etiam salvatorem expectamus Dominum Iesum Christum
PHIL|3|21|qui reformabit corpus humilitatis nostrae configuratum corpori claritatis suae secundum operationem qua possit etiam subicere sibi omnia
PHIL|4|1|itaque fratres mei carissimi et desiderantissimi gaudium meum et corona mea sic state in Domino carissimi
PHIL|4|2|Euhodiam rogo et Syntychen deprecor id ipsum sapere in Domino
PHIL|4|3|etiam rogo et te germane conpar adiuva illas quae mecum laboraverunt in evangelio cum Clemente et ceteris adiutoribus meis quorum nomina sunt in libro vitae
PHIL|4|4|gaudete in Domino semper iterum dico gaudete
PHIL|4|5|modestia vestra nota sit omnibus hominibus Dominus prope
PHIL|4|6|nihil solliciti sitis sed in omni oratione et obsecratione cum gratiarum actione petitiones vestrae innotescant apud Deum
PHIL|4|7|et pax Dei quae exsuperat omnem sensum custodiat corda vestra et intellegentias vestras in Christo Iesu
PHIL|4|8|de cetero fratres quaecumque sunt vera quaecumque pudica quaecumque iusta quaecumque sancta quaecumque amabilia quaecumque bonae famae si qua virtus si qua laus haec cogitate
PHIL|4|9|quae et didicistis et accepistis et audistis et vidistis in me haec agite et Deus pacis erit vobiscum
PHIL|4|10|gavisus sum autem in Domino vehementer quoniam tandem aliquando refloruistis pro me sentire sicut et sentiebatis occupati autem eratis
PHIL|4|11|non quasi propter penuriam dico ego enim didici in quibus sum sufficiens esse
PHIL|4|12|scio et humiliari scio et abundare ubique et in omnibus institutus sum et satiari et esurire et abundare et penuriam pati
PHIL|4|13|omnia possum in eo qui me confortat
PHIL|4|14|verumtamen bene fecistis communicantes tribulationi meae
PHIL|4|15|scitis autem et vos Philippenses quod in principio evangelii quando profectus sum a Macedonia nulla mihi ecclesia communicavit in ratione dati et accepti nisi vos soli
PHIL|4|16|quia et Thessalonicam et semel et bis in usum mihi misistis
PHIL|4|17|non quia quaero datum sed requiro fructum abundantem in rationem vestram
PHIL|4|18|habeo autem omnia et abundo repletus sum acceptis ab Epafrodito quae misistis odorem suavitatis hostiam acceptam placentem Deo
PHIL|4|19|Deus autem meus impleat omne desiderium vestrum secundum divitias suas in gloria in Christo Iesu
PHIL|4|20|Deo autem et Patri nostro gloria in saecula saeculorum amen
PHIL|4|21|salutate omnem sanctum in Christo Iesu salutant vos qui mecum sunt fratres
PHIL|4|22|salutant vos omnes sancti maxime autem qui de Caesaris domo sunt
PHIL|4|23|gratia Domini Iesu Christi cum spiritu vestro amen
