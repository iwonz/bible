1PET|1|1|Peter, an apostle of Jesus Christ, To those who are elect exiles of the dispersion in Pontus, Galatia, Cappadocia, Asia, and Bithynia,
1PET|1|2|according to the foreknowledge of God the Father, in the sanctification of the Spirit, for obedience to Jesus Christ and for sprinkling with his blood: May grace and peace be multiplied to you.
1PET|1|3|Blessed be the God and Father of our Lord Jesus Christ! According to his great mercy, he has caused us to be born again to a living hope through the resurrection of Jesus Christ from the dead,
1PET|1|4|to an inheritance that is imperishable, undefiled, and unfading, kept in heaven for you,
1PET|1|5|who by God's power are being guarded through faith for a salvation ready to be revealed in the last time.
1PET|1|6|In this you rejoice, though now for a little while, as was necessary, you have been grieved by various trials,
1PET|1|7|so that the tested genuineness of your faith- more precious than gold that perishes though it is tested by fire- may be found to result in praise and glory and honor at the revelation of Jesus Christ.
1PET|1|8|Though you have not seen him, you love him. Though you do not now see him, you believe in him and rejoice with joy that is inexpressible and filled with glory,
1PET|1|9|obtaining the outcome of your faith, the salvation of your souls.
1PET|1|10|Concerning this salvation, the prophets who prophesied about the grace that was to be yours searched and inquired carefully,
1PET|1|11|inquiring what person or time the Spirit of Christ in them was indicating when he predicted the sufferings of Christ and the subsequent glories.
1PET|1|12|It was revealed to them that they were serving not themselves but you, in the things that have now been announced to you through those who preached the good news to you by the Holy Spirit sent from heaven, things into which angels long to look.
1PET|1|13|Therefore, preparing your minds for action, and being sober-minded, set your hope fully on the grace that will be brought to you at the revelation of Jesus Christ.
1PET|1|14|As obedient children, do not be conformed to the passions of your former ignorance,
1PET|1|15|but as he who called you is holy, you also be holy in all your conduct,
1PET|1|16|since it is written, "You shall be holy, for I am holy."
1PET|1|17|And if you call on him as Father who judges impartially according to each one's deeds, conduct yourselves with fear throughout the time of your exile,
1PET|1|18|knowing that you were ransomed from the futile ways inherited from your forefathers, not with perishable things such as silver or gold,
1PET|1|19|but with the precious blood of Christ, like that of a lamb without blemish or spot.
1PET|1|20|He was foreknown before the foundation of the world but was made manifest in the last times for your sake,
1PET|1|21|who through him are believers in God, who raised him from the dead and gave him glory, so that your faith and hope are in God.
1PET|1|22|Having purified your souls by your obedience to the truth for a sincere brotherly love, love one another earnestly from a pure heart,
1PET|1|23|since you have been born again, not of perishable seed but of imperishable, through the living and abiding word of God;
1PET|1|24|for "All flesh is like grass and all its glory like the flower of grass. The grass withers, and the flower falls,
1PET|1|25|but the word of the Lord remains forever." And this word is the good news that was preached to you.
1PET|2|1|So put away all malice and all deceit and hypocrisy and envy and all slander.
1PET|2|2|Like newborn infants, long for the pure spiritual milk, that by it you may grow up to salvation-
1PET|2|3|if indeed you have tasted that the Lord is good.
1PET|2|4|As you come to him, a living stone rejected by men but in the sight of God chosen and precious,
1PET|2|5|you yourselves like living stones are being built up as a spiritual house, to be a holy priesthood, to offer spiritual sacrifices acceptable to God through Jesus Christ.
1PET|2|6|For it stands in Scripture: "Behold, I am laying in Zion a stone, a cornerstone chosen and precious, and whoever believes in him will not be put to shame."
1PET|2|7|So the honor is for you who believe, but for those who do not believe, "The stone that the builders rejected has become the cornerstone,"
1PET|2|8|and "A stone of stumbling, and a rock of offense." They stumble because they disobey the word, as they were destined to do.
1PET|2|9|But you are a chosen race, a royal priesthood, a holy nation, a people for his own possession, that you may proclaim the excellencies of him who called you out of darkness into his marvelous light.
1PET|2|10|Once you were not a people, but now you are God's people; once you had not received mercy, but now you have received mercy.
1PET|2|11|Beloved, I urge you as sojourners and exiles to abstain from the passions of the flesh, which wage war against your soul.
1PET|2|12|Keep your conduct among the Gentiles honorable, so that when they speak against you as evildoers, they may see your good deeds and glorify God on the day of visitation.
1PET|2|13|Be subject for the Lord's sake to every human institution, whether it be to the emperor as supreme,
1PET|2|14|or to governors as sent by him to punish those who do evil and to praise those who do good.
1PET|2|15|For this is the will of God, that by doing good you should put to silence the ignorance of foolish people.
1PET|2|16|Live as people who are free, not using your freedom as a cover-up for evil, but living as servants of God.
1PET|2|17|Honor everyone. Love the brotherhood. Fear God. Honor the emperor.
1PET|2|18|Servants, be subject to your masters with all respect, not only to the good and gentle but also to the unjust.
1PET|2|19|For this is a gracious thing, when, mindful of God, one endures sorrows while suffering unjustly.
1PET|2|20|For what credit is it if, when you sin and are beaten for it, you endure? But if when you do good and suffer for it you endure, this is a gracious thing in the sight of God.
1PET|2|21|For to this you have been called, because Christ also suffered for you, leaving you an example, so that you might follow in his steps.
1PET|2|22|He committed no sin, neither was deceit found in his mouth.
1PET|2|23|When he was reviled, he did not revile in return; when he suffered, he did not threaten, but continued entrusting himself to him who judges justly.
1PET|2|24|He himself bore our sins in his body on the tree, that we might die to sin and live to righteousness. By his wounds you have been healed.
1PET|2|25|For you were straying like sheep, but have now returned to the Shepherd and Overseer of your souls.
1PET|3|1|Likewise, wives, be subject to your own husbands, so that even if some do not obey the word, they may be won without a word by the conduct of their wives-
1PET|3|2|when they see your respectful and pure conduct.
1PET|3|3|Do not let your adorning be external- the braiding of hair, the wearing of gold, or the putting on of clothing-
1PET|3|4|but let your adorning be the hidden person of the heart with the imperishable beauty of a gentle and quiet spirit, which in God's sight is very precious.
1PET|3|5|For this is how the holy women who hoped in God used to adorn themselves, by submitting to their husbands,
1PET|3|6|as Sarah obeyed Abraham, calling him lord. And you are her children, if you do good and do not fear anything that is frightening.
1PET|3|7|Likewise, husbands, live with your wives in an understanding way, showing honor to the woman as the weaker vessel, since they are heirs with you of the grace of life, so that your prayers may not be hindered.
1PET|3|8|Finally, all of you, have unity of mind, sympathy, brotherly love, a tender heart, and a humble mind.
1PET|3|9|Do not repay evil for evil or reviling for reviling, but on the contrary, bless, for to this you were called, that you may obtain a blessing.
1PET|3|10|For "Whoever desires to love life and see good days, let him keep his tongue from evil and his lips from speaking deceit;
1PET|3|11|let him turn away from evil and do good; let him seek peace and pursue it.
1PET|3|12|For the eyes of the Lord are on the righteous, and his ears are open to their prayer. But the face of the Lord is against those who do evil."
1PET|3|13|Now who is there to harm you if you are zealous for what is good?
1PET|3|14|But even if you should suffer for righteousness' sake, you will be blessed. Have no fear of them, nor be troubled,
1PET|3|15|but in your hearts regard Christ the Lord as holy, always being prepared to make a defense to anyone who asks you for a reason for the hope that is in you;
1PET|3|16|yet do it with gentleness and respect, having a good conscience, so that, when you are slandered, those who revile your good behavior in Christ may be put to shame.
1PET|3|17|For it is better to suffer for doing good, if that should be God's will, than for doing evil.
1PET|3|18|For Christ also suffered once for sins, the righteous for the unrighteous, that he might bring us to God, being put to death in the flesh but made alive in the spirit,
1PET|3|19|in which he went and proclaimed to the spirits in prison,
1PET|3|20|because they formerly did not obey, when God's patience waited in the days of Noah, while the ark was being prepared, in which a few, that is, eight persons, were brought safely through water.
1PET|3|21|Baptism, which corresponds to this, now saves you, not as a removal of dirt from the body but as an appeal to God for a good conscience, through the resurrection of Jesus Christ,
1PET|3|22|who has gone into heaven and is at the right hand of God, with angels, authorities, and powers having been subjected to him.
1PET|4|1|Since therefore Christ suffered in the flesh, arm yourselves with the same way of thinking, for whoever has suffered in the flesh has ceased from sin,
1PET|4|2|so as to live for the rest of the time in the flesh no longer for human passions but for the will of God.
1PET|4|3|The time that is past suffices for doing what the Gentiles want to do, living in sensuality, passions, drunkenness, orgies, drinking parties, and lawless idolatry.
1PET|4|4|With respect to this they are surprised when you do not join them in the same flood of debauchery, and they malign you;
1PET|4|5|but they will give account to him who is ready to judge the living and the dead.
1PET|4|6|For this is why the gospel was preached even to those who are dead, that though judged in the flesh the way people are, they might live in the spirit the way God does.
1PET|4|7|The end of all things is at hand; therefore be self-controlled and sober-minded for the sake of your prayers.
1PET|4|8|Above all, keep loving one another earnestly, since love covers a multitude of sins.
1PET|4|9|Show hospitality to one another without grumbling.
1PET|4|10|As each has received a gift, use it to serve one another, as good stewards of God's varied grace:
1PET|4|11|whoever speaks, as one who speaks oracles of God; whoever serves, as one who serves by the strength that God supplies- in order that in everything God may be glorified through Jesus Christ. To him belong glory and dominion forever and ever. Amen.
1PET|4|12|Beloved, do not be surprised at the fiery trial when it comes upon you to test you, as though something strange were happening to you.
1PET|4|13|But rejoice insofar as you share Christ's sufferings, that you may also rejoice and be glad when his glory is revealed.
1PET|4|14|If you are insulted for the name of Christ, you are blessed, because the Spirit of glory and of God rests upon you.
1PET|4|15|But let none of you suffer as a murderer or a thief or an evildoer or as a meddler.
1PET|4|16|Yet if anyone suffers as a Christian, let him not be ashamed, but let him glorify God in that name.
1PET|4|17|For it is time for judgment to begin at the household of God; and if it begins with us, what will be the outcome for those who do not obey the gospel of God?
1PET|4|18|And "If the righteous is scarcely saved, what will become of the ungodly and the sinner?"
1PET|4|19|Therefore let those who suffer according to God's will entrust their souls to a faithful Creator while doing good.
1PET|5|1|So I exhort the elders among you, as a fellow elder and a witness of the sufferings of Christ, as well as a partaker in the glory that is going to be revealed:
1PET|5|2|shepherd the flock of God that is among you, exercising oversight, not under compulsion, but willingly, as God would have you; not for shameful gain, but eagerly;
1PET|5|3|not domineering over those in your charge, but being examples to the flock.
1PET|5|4|And when the chief Shepherd appears, you will receive the unfading crown of glory.
1PET|5|5|Likewise, you who are younger, be subject to the elders. Clothe yourselves, all of you, with humility toward one another, for "God opposes the proud but gives grace to the humble."
1PET|5|6|Humble yourselves, therefore, under the mighty hand of God so that at the proper time he may exalt you,
1PET|5|7|casting all your anxieties on him, because he cares for you.
1PET|5|8|Be sober-minded; be watchful. Your adversary the devil prowls around like a roaring lion, seeking someone to devour.
1PET|5|9|Resist him, firm in your faith, knowing that the same kinds of suffering are being experienced by your brotherhood throughout the world.
1PET|5|10|And after you have suffered a little while, the God of all grace, who has called you to his eternal glory in Christ, will himself restore, confirm, strengthen, and establish you.
1PET|5|11|To him be the dominion forever and ever. Amen.
1PET|5|12|By Silvanus, a faithful brother as I regard him, I have written briefly to you, exhorting and declaring that this is the true grace of God. Stand firm in it.
1PET|5|13|She who is at Babylon, who is likewise chosen, sends you greetings, and so does Mark, my son.
1PET|5|14|Greet one another with the kiss of love. Peace to all of you who are in Christ.
