PS|1|1|Beatus vir, qui non abiit in consilio impiorumet in via peccatorum non stetitet in conventu derisorum non sedit,
PS|1|2|sed in lege Domini voluntas eius,et in lege eius meditatur die ac nocte.
PS|1|3|Et erit tamquam lignum plantatum secus decursus aquarum,quod fructum suum dabit in tempore suo;et folium eius non defluet,et omnia, quaecumque faciet, prosperabuntur.
PS|1|4|Non sic impii, non sic,sed tamquam pulvis, quem proicit ventus.
PS|1|5|Ideo non consurgent impii in iudicio,neque peccatores in concilio iustorum.
PS|1|6|Quoniam novit Dominus viam iustorum,et iter impiorum peribit.
PS|2|1|Quare fremuerunt gentes,et populi meditati sunt inania?
PS|2|2|Astiterunt reges terrae,et principes convenerunt in unumadversus Dominum et adversus christum eius:
PS|2|3|" Dirumpamus vincula eorumet proiciamus a nobis iugum ipsorum! ".
PS|2|4|Qui habitat in caelis, irridebit eos,Dominus subsannabit eos.
PS|2|5|Tunc loquetur ad eos in ira suaet in furore suo conturbabit eos:
PS|2|6|" Ego autem constitui regem meum super Sion, montem sanctum meum! ".
PS|2|7|Praedicabo decretum eius.Dominus dixit ad me: " Filius meus es tu;ego hodie genui te.
PS|2|8|Postula a me, et dabo tibi gentes hereditatem tuamet possessionem tuam terminos terrae.
PS|2|9|Reges eos in virga ferreaet tamquam vas figuli confringes eos ".
PS|2|10|Et nunc, reges, intellegite;erudimini, qui iudicatis terram.
PS|2|11|Servite Domino in timoreet exsultate ei cum tremore.
PS|2|12|Apprehendite disciplinam, ne quando irascatur,et pereatis de via,cum exarserit in brevi ira eius.Beati omnes, qui confidunt in eo.
PS|3|1|PSALMUS. David, cum fugit a filio suo Absalom.
PS|3|2|Domine, quid multiplicati sunt, qui tribulant me?Multi insurgunt adversum me,
PS|3|3|multi dicunt animae meae: Non est salus ipsi in Deo ".
PS|3|4|Tu autem, Domine, protector meus es,gloria mea et exaltans caput meum.
PS|3|5|Voce mea ad Dominum clamavi,et exaudivit me de monte sancto suo.
PS|3|6|Ego obdormivi et soporatus sum,exsurrexi, quia Dominus suscepit me.
PS|3|7|Non timebo milia populi circumdantis me.Exsurge, Domine salvum me fac, Deus meus;
PS|3|8|quoniam tu percussisti in maxillam omnes adversantes mihi,dentes peccatorum contrivisti.
PS|3|9|Domini est salus,et super populum tuum benedictio tua.
PS|4|1|Magistro chori. Fidibus. PSALMUS. David.
PS|4|2|Cum invocarem, exaudivit me Deus iustitiae meae.In tribulatione dilatasti mihi;miserere mei et exaudi orationem meam.
PS|4|3|Filii hominum, usquequo gravi corde?Ut quid diligitis vanitatem et quaeritis mendacium?
PS|4|4|Et scitote quoniam mirificavit Dominus sanctum suum;Dominus exaudiet, cum clamavero ad eum.
PS|4|5|Irascimini et nolite peccare;loquimini in cordibus vestris,in cubilibus vestris et conquiescite.
PS|4|6|Sacrificate sacrificium iustitiaeet sperate in Domino.
PS|4|7|Multi dicunt: " Quis ostendit nobis bona? ".Leva in signum super nos lumen vultus tui, Domine!
PS|4|8|Maiorem dedisti laetitiam in corde meo,quam cum multiplicantur frumentum et vinum eorum.
PS|4|9|In pace in idipsum dormiam et requiescam,quoniam tu, Domine, singulariter in spe constituisti me.
PS|5|1|Magistro chori. Ad tibias. PSALMUS. David.
PS|5|2|Verba mea auribus percipe, Domine;intellege gemitum meum.
PS|5|3|Intende voci clamoris mei,rex meus et Deus meus.
PS|5|4|Quoniam ad te orabo, Domine,mane exaudies vocem meam;mane astabo tibi et exspectabo.
PS|5|5|Quoniam non Deus volens iniquitatem tu es;neque habitabit iuxta te malignus,
PS|5|6|neque permanebunt iniusti ante oculos tuos.
PS|5|7|Odisti omnes, qui operantur iniquitatem,perdes omnes, qui loquuntur mendacium;virum sanguinum et dolosum abominabitur Dominus.
PS|5|8|Ego autem in multitudine misericordiae tuaeintroibo in domum tuam;adorabo ad templum sanctum tuum in timore tuo.
PS|5|9|Domine, deduc me in iustitia tua propter inimicos meos,dirige in conspectu meo viam tuam.
PS|5|10|Quoniam non est in ore eorum veritas,cor eorum fovea;sepulcrum patens est guttur eorum,molliunt linguas suas.
PS|5|11|Iudica illos, Deus; decidant a cogitationibus suis;secundum multitudinem impietatum eorum expelle eos,quoniam irritaverunt te, Domine.
PS|5|12|Et omnes, qui sperant in te,laetentur, in aeternum exsultent.Obumbrabis eis, et gloriabuntur in te,qui diligunt nomen tuum;
PS|5|13|quoniam tu benedices iusto, Domine,quasi scuto, bona voluntate coronabis eum.
PS|6|1|Magistro chori. Fidibus. Super octavam. PSALMUS. David.
PS|6|2|Domine, ne in furore tuo arguas meneque in ira tua corripias me.
PS|6|3|Miserere mei, Domine, quoniam infirmus sum;sana me, Domine, quoniam conturbata sunt ossa mea.
PS|6|4|Et anima mea turbata est valde,sed tu, Domine, usquequo?
PS|6|5|Convertere, Domine, eripe animam meam;salvum me fac propter misericordiam tuam.
PS|6|6|Quoniam non est in morte, qui memor sit tui;in inferno autem quis confitebitur tibi?
PS|6|7|Laboravi in gemitu meo,lavabam per singulas noctes lectum meum;lacrimis meis stratum meum rigabam.
PS|6|8|Turbatus est a maerore oculus meus,inveteravi inter omnes inimicos meos.
PS|6|9|Discedite a me, omnes, qui operamini iniquitatem,quoniam exaudivit Dominus vocem fletus mei.
PS|6|10|Exaudivit Dominus deprecationem meam,Dominus orationem meam suscepit.
PS|6|11|Erubescant et conturbentur vehementer omnes inimici mei;convertantur et erubescant valde velociter.
PS|7|1|Lamentatio David, quam cantavit Domino propter Chus Beniaminitam.
PS|7|2|Domine Deus meus, in te speravi;salvum me fac ex omnibus persequentibus me et libera me,
PS|7|3|ne quando rapiat ut leo animam meamdiscerpens, dum non est qui salvum faciat.
PS|7|4|Domine Deus meus, si feci istud,si est iniquitas in manibus meis,
PS|7|5|si reddidi retribuenti mihi malaet exspoliavi inimicum meum dimittens inanem,
PS|7|6|persequatur inimicus animam meam et comprehendatet conculcet in terra vitam meamet gloriam meam in pulverem deducat.
PS|7|7|Exsurge, Domine, in ira tuaet exaltare contra indignationem inimicorum meorumet exsurge, Deus meus, in iudicio, quod mandasti.
PS|7|8|Et synagoga populorum circumdabit te,et super hanc in altum regredere:
PS|7|9|Dominus iudicat populos.Iudica me, Domine, secundum iustitiam meamet secundum innocentiam meam, quae est in me.
PS|7|10|Consumatur nequitia peccatorum;et iustum confirma:scrutans corda et renes Deus iustus.
PS|7|11|Adiutorium meum apud Deum,qui salvos facit rectos corde.
PS|7|12|Deus iudex iustus,fortis, irascens per singulos dies.
PS|7|13|Nonne iterum gladium suum exacuit,arcum suum tetendit et paravit illum?
PS|7|14|Et paravit sibi vasa mortis,sagittas suas ardentes effecit.
PS|7|15|Ecce parturiit iniustitiam,concepit dolorem et peperit iniquitatem;
PS|7|16|lacum aperuit et effodit eumet incidit in foveam, quam fecit.
PS|7|17|Convertetur dolor eius in caput eius,et in verticem ipsius iniquitas eius descendet.
PS|7|18|Confitebor Domino secundum iustitiam eiuset psallam nomini Domini Altissimi.
PS|8|1|Magistro chori. Ad modum cantici " Torcularia... ". PSALMUS. David.
PS|8|2|Domine, Dominus noster,quam admirabile est nomen tuum in universa terra,quoniam elevata est magnificentia tua super caelos.
PS|8|3|Ex ore infantium et lactantium perfecisti laudempropter inimicos tuos,ut destruas inimicum et ultorem.
PS|8|4|Quando video caelos tuos, opera digitorum tuorum,lunam et stellas, quae tu fundasti,
PS|8|5|quid est homo, quod memor es eius,aut filius hominis, quoniam visitas eum?
PS|8|6|Minuisti eum paulo minus ab angelis,gloria et honore coronasti eum
PS|8|7|et constituisti eum super opera manuum tuarum.Omnia subiecisti sub pedibus eius:
PS|8|8|oves et boves universas,insuper et pecora campi,
PS|8|9|volucres caeli et pisces maris,quaecumque perambulant semitas maris.
PS|8|10|Domine, Dominus noster,quam admirabile est nomen tuum in universa terra!
PS|9|1|Magistro chori. Ad modum cantici " Mut labben ". PSALMUS. David.
PS|9|2|ALEPH. Confitebor tibi, Domine, in toto corde meo,narrabo omnia mirabilia tua.
PS|9|3|Laetabor et exsultabo in te,psallam nomini tuo, Altissime.
PS|9|4|BETH. Cum convertuntur inimici mei retrorsum,infirmantur et pereunt a facie tua.
PS|9|5|Quoniam fecisti iudicium meum et causam meam,sedisti super thronum, qui iudicas iustitiam.
PS|9|6|GHIMEL. Increpasti gentes, perdidisti impium;nomen eorum delesti in aeternum et in saeculum saeculi.
PS|9|7|Inimici defecerunt, solitudines sempiternae factae sunt;et civitates destruxisti: periit memoria eorum cum ipsis.
PS|9|8|HE. Dominus autem in aeternum sedebit,paravit in iudicium thronum suum;
PS|9|9|et ipse iudicabit orbem terrae in iustitia,iudicabit populos in aequitate.
PS|9|10|VAU. Et erit Dominus refugium oppresso,refugium in opportunitatibus, in tribulatione.
PS|9|11|Et sperent in te, qui noverunt nomen tuum,quoniam non dereliquisti quaerentes te, Domine.
PS|9|12|ZAIN. Psallite Domino, qui habitat in Sion;annuntiate inter gentes studia eius.
PS|9|13|Quoniam requirens sanguinem recordatus est eorum,non est oblitus clamorem pauperum.
PS|9|14|HETH. Miserere mei, Domine;vide afflictionem meam de inimicis meis,qui exaltas me de portis mortis,
PS|9|15|ut annuntiem omnes laudationes tuas in portis filiae Sion,exsultem in salutari tuo.
PS|9|16|TETH. Infixae sunt gentes in fovea, quam fecerunt;in laqueo isto, quem absconderunt,comprehensus est pes eorum.
PS|9|17|Manifestavit se Dominus iudicium faciens;in operibus manuum suarum comprehensus est peccator.
PS|9|18|IOD. Convertentur peccatores in infernum,omnes gentes, quae obliviscuntur Deum.
PS|9|19|CAPH. Quoniam non in finem oblivio erit pauperis;exspectatio pauperum non peribit in aeternum.
PS|9|20|Exsurge, Domine, non confortetur homo;iudicentur gentes in conspectu tuo.
PS|9|21|Constitue, Domine, terrorem super eos;sciant gentes quoniam homines sunt.
PS|10|1|LAMED. Ut quid, Domine, stas a longe,abscondis te in opportunitatibus, in tribulatione?
PS|10|2|Dum superbit, impius insequitur pauperem;comprehendantur in consiliis, quae cogitant.
PS|10|3|Quoniam gloriatur peccator in desideriis animae suae,et avarus sibi benedicit.
PS|10|4|NUN. Spernit Dominum peccator in arrogantia sua: Non requiret; non est Deus ".
PS|10|5|Hae sunt omnes cogitationes eius;prosperantur viae illius in omni tempore.Excelsa nimis iudicia tua a facie eius;omnes inimicos suos aspernatur.
PS|10|6|Dixit enim in corde suo: " Non movebor;in generationem et generationem ero sine malo ".
PS|10|7|PHE. Cuius maledictione os plenum est et fraudulentia et dolo,sub lingua eius labor et nequitia.
PS|10|8|Sedet in insidiis ad vicos,in occultis interficit innocentem.
PS|10|9|SADE. Oculi eius in pauperem respiciunt;insidiatur in abscondito quasi leo in spelunca sua.Insidiatur, ut rapiat pauperem;rapit pauperem, dum attrahit in laqueum suum.
PS|10|10|Irruit et inclinat se, et miseri caduntin fortitudine brachiorum eius.
PS|10|11|Dixit enim in corde suo: " Oblitus est Deus;avertit faciem suam, non videbit in finem ". -
PS|10|12|COPH. Exsurge, Domine Deus, exalta manum tuam,ne obliviscaris pauperum.
PS|10|13|Propter quid spernit impius Deum?Dixit enim in corde suo: " Non requires ".
PS|10|14|RES. Vidisti: tu laborem et dolorem consideras,ut tradas eos in manus tuas.Tibi derelictus est pauper,orphano tu factus es adiutor.
PS|10|15|SIN. Contere brachium peccatoris et maligni;quaeres peccatum illius et non invenies.
PS|10|16|Dominus rex in aeternum et in saeculum saeculi:perierunt gentes de terra illius.
PS|10|17|TAU. Desiderium pauperum exaudisti, Domine;confirmabis cor eorum, intendes aurem tuam
PS|10|18|iudicare pupillo et humili,ut non apponat ultra inducere timorem homo de terra.
PS|11|1|Magistro chori. David.In Domino confido, quomodo dicitis animae meae: Transmigra in montem sicut passer!
PS|11|2|Quoniam ecce peccatores intenderunt arcum,paraverunt sagittas suas super nervum,ut sagittent in obscuro rectos corde.
PS|11|3|Quando fundamenta evertuntur,iustus quid faciat? ".
PS|11|4|Dominus in templo sancto suo,Dominus, in caelo sedes eius.Oculi eius in pauperem respiciunt,palpebrae eius interrogant filios hominum.
PS|11|5|Dominus interrogat iustum et impium;qui autem diligit iniquitatem, odit anima eius.
PS|11|6|Pluet super peccatores carbones ignis et sulphur;et spiritus procellarum pars calicis eorum.
PS|11|7|Quoniam iustus Dominus et iustitias dilexit,recti videbunt vultum eius.
PS|12|1|Magistro chori. Super octavam. PSALMUS. David.
PS|12|2|Salvum me fac, Domine, quoniam defecit sanctus,quoniam deminuti sunt fideles a filiis hominum.
PS|12|3|Vana locuti sunt unusquisque ad proximum suum;in labiis dolosis, in duplici corde locuti sunt.
PS|12|4|Disperdat Dominus universa labia dolosaet linguam magniloquam.
PS|12|5|Qui dixerunt: " Lingua nostra magnificabimur,labia nostra a nobis sunt;quis noster dominus est? ".
PS|12|6|" Propter miseriam inopum et gemitum pauperum,nunc exsurgam, dicit Dominus;ponam in salutari illum, quem despiciunt ".
PS|12|7|Eloquia Domini eloquia casta,argentum igne examinatum, separatum a terra,purgatum septuplum.
PS|12|8|Tu, Domine, servabis nos et custodies nosa generatione hac in aeternum.In circuitu impii ambulant,cum exaltantur sordes inter filios hominum.
PS|13|1|Magistro chori. PSALMUS. David.
PS|13|2|Usquequo, Domine, oblivisceris me in finem?Usquequo avertes faciem tuam a me?
PS|13|3|Usquequo ponam consilia in anima mea,dolorem in corde meo per diem?Usquequo exaltabitur inimicus meus super me?
PS|13|4|Respice et exaudi me, Domine Deus meus.Illumina oculos meos, ne quando obdormiam in morte,
PS|13|5|ne quando dicat inimicus meus: " Praevalui adversus eum! ";neque exsultent, qui tribulant me, si motus fuero.
PS|13|6|Ego autem in misericordia tua speravi.Exsultabit cor meum in salutari tuo;cantabo Domino, qui bona tribuit mihi.
PS|14|1|Magistro chori. David.Dixit insipiens in corde suo: " Non est Deus ".Corrupti sunt et abominationes operati sunt;non est qui faciat bonum.
PS|14|2|Dominus de caelo prospexit super filios hominum,ut videret si est intellegens aut requirens Deum.
PS|14|3|Omnes declinaverunt, simul corrupti sunt;non est qui faciat bonum, non est usque ad unum.
PS|14|4|Nonne scient omnes, qui operantur iniquitatem,qui devorant plebem meam sicut escam panis?Dominum non invocaverunt;
PS|14|5|illic trepidaverunt timore,quoniam Deus cum generatione iusta est.
PS|14|6|Vos consilium inopis confundetis,Dominus autem spes eius est.
PS|14|7|Quis dabit ex Sion salutare Israel?Cum converterit Dominus captivitatem plebis suae,exsultabit Iacob, et laetabitur Israel.
PS|15|1|PSALMUS. David.Domine, quis habitabit in tabernaculo tuo?Quis requiescet in monte sancto tuo?
PS|15|2|Qui ingreditur sine macula et operatur iustitiam,qui loquitur veritatem in corde suo,
PS|15|3|qui non egit dolum in lingua suanec fecit proximo suo malumet opprobrium non intulit proximo suo.
PS|15|4|Ad nihilum reputatus est in conspectu eius malignus,timentes autem Dominum glorificat.Qui iuravit in detrimentum suum et non mutat,
PS|15|5|qui pecuniam suam non dedit ad usuramet munera super innocentem non accepit.Qui facit haec, non movebitur in aeternum.
PS|16|1|Miktam. David.Conserva me, Deus, quoniam speravi in te.
PS|16|2|Dixi Domino: " Dominus meus es tu, bonum mihi non est sine te ".
PS|16|3|In sanctos, qui sunt in terra, inclitos viros,omnis voluntas mea in eos.
PS|16|4|Multiplicantur dolores eorum, qui post deos alienos acceleraverunt.Non effundam libationes eorum de sanguinibusneque assumam nomina eorum in labiis meis.
PS|16|5|Dominus pars hereditatis meae et calicis mei:tu es qui detines sortem meam.
PS|16|6|Funes ceciderunt mihi in praeclaris;insuper et hereditas mea speciosa est mihi.
PS|16|7|Benedicam Dominum, qui tribuit mihi intellectum;insuper et in noctibus erudierunt me renes mei.
PS|16|8|Proponebam Dominum in conspectu meo semper;quoniam a dextris est mihi, non commovebor.
PS|16|9|Propter hoc laetatum est cor meum,et exsultaverunt praecordia mea;insuper et caro mea requiescet in spe.
PS|16|10|Quoniam non derelinques animam meam in infernonec dabis sanctum tuum videre corruptionem.
PS|16|11|Notas mihi facies vias vitae,plenitudinem laetitiae cum vultu tuo,delectationes in dextera tua usque in finem.
PS|17|1|Precatio. David.Exaudi, Domine, iustitiam meam,intende deprecationem meam.Auribus percipe orationem meam, non in labiis dolosis.
PS|17|2|De vultu tuo iudicium meum prodeat;oculi tui videant aequitates.
PS|17|3|Proba cor meum et visita nocte;igne me examina, et non invenies in me iniquitatem.
PS|17|4|Non transgreditur os meum ad opera hominum,propter verba labiorum tuorum custodivi me a viis violenti.
PS|17|5|Retine gressus meos in semitis tuis,ut non moveantur vestigia mea.
PS|17|6|Ego ad te clamavi, quoniam exaudis me, Deus;inclina aurem tuam mihi et exaudi verba mea.
PS|17|7|Mirifica misericordias tuas,qui salvos facis ab insurgentibussperantes in dextera tua.
PS|17|8|Custodi me ut pupillam oculi,sub umbra alarum tuarum protege me
PS|17|9|a facie impiorum, qui me afflixerunt.Inimici mei in furore circumdederunt me,
PS|17|10|adipem suum concluserunt;os eorum locutum est superbiam.
PS|17|11|Incedentes nunc circumdederunt me,oculos suos statuerunt prosternere in terram.
PS|17|12|Aspectus eorum quasi leonis parati ad praedamet sicut catuli leonis recubantis in abditis.
PS|17|13|Exsurge, Domine, praeveni eum, supplanta eum;eripe animam meam ab impio framea tua,
PS|17|14|a mortuis manu tua, Domine,a mortuis, quorum defecit portio vitae.De reconditis tuis adimpleas ventrem eorum,saturentur filii et dimittant reliquias parvulis suis.
PS|17|15|Ego autem in iustitia videbo faciem tuam;satiabor, cum evigilavero, conspectu tuo.
PS|18|1|Magistro chori. David, servi Domini,qui locutus est ad Dominum verba huius cantici,quando Dominus eum liberaverate potestate omnium inimicorum suorum
PS|18|2|et e manu Saul. Dixit igitur:Diligam te, Domine, fortitudo mea.
PS|18|3|Domine, firmamentum meum et refugium meum et liberator meus;Deus meus, adiutor meus, et sperabo in eum;protector meus et cornu salutis meae et susceptor meus.
PS|18|4|Laudabilem invocabo Dominum,et ab inimicis meis salvus ero.
PS|18|5|Circumdederunt me fluctus mortis,et torrentes Belial conturbaverunt me;
PS|18|6|funes inferni circumdederunt me,praeoccupaverunt me laquei mortis.
PS|18|7|In tribulatione mea invocavi Dominumet ad Deum meum clamavi;exaudivit de templo suo vocem meam,et clamor meus in conspectu eius introivit in aures eius.
PS|18|8|Commota est et contremuit terra;fundamenta montium concussa suntet commota sunt, quoniam iratus est.
PS|18|9|Ascendit fumus de naribus eius,et ignis de ore eius devorans;carbones succensi processerunt ab eo.
PS|18|10|Inclinavit caelos et descendit,et caligo sub pedibus eius.
PS|18|11|Et ascendit super cherub et volavit,ferebatur super pennas ventorum.
PS|18|12|Et posuit tenebras latibulum suum,in circuitu eius tabernaculum eius,tenebrosa aqua, nubes aeris.
PS|18|13|Prae fulgore in conspectu eius nubes transierunt,grando et carbones ignis.
PS|18|14|Et intonuit de caelo Dominus,et Altissimus dedit vocem suam:grando et carbones ignis.
PS|18|15|Et misit sagittas suas et dissipavit eos,fulgura iecit et conturbavit eos.
PS|18|16|Et apparuerunt fontes aquarum,et revelata sunt fundamenta orbis terrarumab increpatione tua, Domine,ab inspiratione spiritus irae tuae.
PS|18|17|Misit de summo et accepit meet assumpsit me de aquis multis;
PS|18|18|eripuit me de inimicis meis fortissimiset ab his, qui oderunt me,quoniam confortati sunt super me.
PS|18|19|Oppugnaverunt me in die afflictionis meae,et factus est Dominus fulcimentum meum;
PS|18|20|et eduxit me in latitudinem,salvum me fecit, quoniam voluit me.
PS|18|21|Et retribuet mihi Dominus secundum iustitiam meamet secundum puritatem manuum mearum reddet mihi,
PS|18|22|quia custodivi vias Domininec impie recessi a Deo meo.
PS|18|23|Quoniam omnia iudicia eius in conspectu meo,et iustitias eius non reppuli a me;
PS|18|24|et fui immaculatus cum eoet observavi me ab iniquitate.
PS|18|25|Et retribuit mihi Dominus secundum iustitiam meamet secundum puritatem manuum mearumin conspectu oculorum eius.
PS|18|26|Cum sancto sanctus eriset cum viro innocente innocens eris
PS|18|27|et cum electo electus eriset cum perverso callidus eris.
PS|18|28|Quoniam tu populum humilem salvum facieset oculos superborum humiliabis.
PS|18|29|Quoniam tu accendis lucernam meam, Domine;Deus meus illuminat tenebras meas.
PS|18|30|Quoniam in te aggrediar hostium turmaset in Deo meo transiliam murum.
PS|18|31|Deus, impolluta via eius,eloquia Domini igne examinata;protector est omnium sperantium in se.
PS|18|32|Quoniam quis Deus praeter Dominum?Aut quae munitio praeter Deum nostrum?
PS|18|33|Deus, qui praecinxit me virtuteet posuit immaculatam viam meam;
PS|18|34|qui perfecit pedes meos tamquam cervorumet super excelsa statuit me;
PS|18|35|qui docet manus meas ad proelium,et tendunt arcum aereum brachia mea.
PS|18|36|Et dedisti mihi scutum salutis tuae,et dextera tua suscepit me,et exauditio tua magnificavit me.
PS|18|37|Dilatasti gressus meos subtus me,et non sunt infirmata vestigia mea.
PS|18|38|Persequebar inimicos meos et comprehendebam illoset non convertebar, donec deficerent.
PS|18|39|Confringebam illos, nec poterant stare,cadebant subtus pedes meos.
PS|18|40|Et praecinxisti me virtute ad bellumet supplantasti insurgentes in me subtus me.
PS|18|41|Et inimicos meos dedisti mihi dorsumet odientes me disperdidisti.
PS|18|42|Clamaverunt, nec erat qui salvos faceret,ad Dominum, nec exaudivit eos.
PS|18|43|Et comminui eos ut pulverem ante faciem venti,ut lutum platearum contrivi eos.
PS|18|44|Eripuisti me de contradictionibus populi,constituisti me in caput gentium.Populus, quem non cognovi, servivit mihi,
PS|18|45|in auditu auris oboedivit mihi.Filii alieni blanditi sunt mihi,
PS|18|46|filii alieni inveterati sunt,contremuerunt in abditis suis.
PS|18|47|Vivit Dominus, et benedictus Adiutor meus,et exaltetur Deus salutis meae.
PS|18|48|Deus, qui das vindictas mihiet subdis populos sub me,liberator meus de inimicis meis iracundis;
PS|18|49|et ab insurgentibus in me exaltas me,a viro iniquo eripis me.
PS|18|50|Propterea confitebor tibi in nationibus, Domine,et nomini tuo psalmum dicam,
PS|18|51|magnificans salutes regis suiet faciens misericordiam christo suoDavid et semini eius usque in saeculum.
PS|19|1|Magistro chori. PSALMUS. David.
PS|19|2|Caeli enarrant gloriam Dei,et opera manuum eius annuntiat firmamentum.
PS|19|3|Dies diei eructat verbum,et nox nocti indicat scientiam.
PS|19|4|Non sunt loquelae neque sermones,quorum non intellegantur voces:
PS|19|5|in omnem terram exivit sonus eorum,et in fines orbis terrae verba eorum.
PS|19|6|Soli posuit tabernaculum in eis,et ipse, tamquam sponsus procedens de thalamo suo,exsultavit ut gigas ad currendam viam.
PS|19|7|A finibus caelorum egressio eius,et occursus eius usque ad fines eorum,nec est quod se abscondat a calore eius.
PS|19|8|Lex Domini immaculata, reficiens animam,testimonium Domini fidele, sapientiam praestans parvulis.
PS|19|9|Iustitiae Domini rectae, laetificantes corda,praeceptum Domini lucidum, illuminans oculos.
PS|19|10|Timor Domini mundus, permanens in saeculum saeculi;iudicia Domini vera, iusta omnia simul,
PS|19|11|desiderabilia super aurum et lapidem pretiosum multum,et dulciora super mel et favum stillantem.
PS|19|12|Etenim servus tuus eruditur in eis;in custodiendis illis retributio multa.
PS|19|13|Errores quis intellegit?Ab occultis munda me
PS|19|14|et a superbia custodi servum tuum, ne dominetur mei,Tunc immaculatus eroet emundabor a delicto maximo.
PS|19|15|Sint ut complaceant eloquia oris mei,et meditatio cordis mei in conspectu tuo.Domine, adiutor meus et redemptor meus.
PS|20|1|Magistro chori. PSALMUS. David.
PS|20|2|Exaudiat te Dominus in die tribulationis,protegat te nomen Dei Iacob.
PS|20|3|Mittat tibi auxilium de sanctoet de Sion tueatur te.
PS|20|4|Memor sit omnis sacrificii tuiet holocaustum tuum pingue habeat.
PS|20|5|Tribuat tibi secundum cor tuumet omne consilium tuum adimpleat.
PS|20|6|Laetabimur in salutari tuoet in nomine Dei nostri levabimus signa;impleat Dominus omnes petitiones tuas.
PS|20|7|Nunc cognovi quoniam salvum fecit Dominus christum suum:exaudivit illum de caelo sancto suo,in virtutibus salutis dexterae eius.
PS|20|8|Hi in curribus, et hi in equis,nos autem nomen Domini Dei nostri invocavimus.
PS|20|9|Ipsi incurvati sunt et ceciderunt,nos autem surreximus et erecti sumus.
PS|20|10|Domine, salvum fac regem,et exaudi nos in die, qua invocaverimus te.
PS|21|1|Magistro chori. PSALMUS. David.
PS|21|2|Domine, in virtute tua laetabitur rexet super salutare tuum exsultabit vehementer.
PS|21|3|Desiderium cordis eius tribuisti eiet voluntatem labiorum eius non denegasti.
PS|21|4|Quoniam praevenisti eum in benedictionibus dulcedinis;posuisti in capite eius coronam de auro purissimo.
PS|21|5|Vitam petiit a te, et tribuisti eilongitudinem dierum in saeculum et in saeculum saeculi.
PS|21|6|Magna est gloria eius in salutari tuo,magnificentiam et decorem impones super eum;
PS|21|7|quoniam pones eum benedictionem in saeculum saeculi,laetificabis eum in gaudio ante vultum tuum.
PS|21|8|Quoniam rex sperat in Dominoet in misericordia Altissimi non commovebitur.
PS|21|9|Inveniet manus tua omnes inimicos tuos,dextera tua inveniet, qui te oderunt.
PS|21|10|Pones eos ut clibanum ignis in tempore vultus tui:Dominus in ira sua deglutiet eos,et devorabit eos ignis.
PS|21|11|Fructum eorum de terra perdeset semen eorum de filiis hominum.
PS|21|12|Quoniam intenderunt in te mala,cogitaverunt consilia: nihil potuerunt.
PS|21|13|Quoniam pones eos dorsum,arcus tuos tendes in vultum eorum.
PS|21|14|Exaltare, Domine, in virtute tua;cantabimus et psallemus virtutes tuas.
PS|22|1|Magistro chori. Ad modum cantici " Cerva diluculo ". PSALMUS. David.
PS|22|2|Deus, Deus meus, quare me dereliquisti?Longe a salute mea verba rugitus mei.
PS|22|3|Deus meus, clamo per diem, et non exaudis,et nocte, et non est requies mihi.
PS|22|4|Tu autem sanctus es,qui habitas in laudibus Israel.
PS|22|5|In te speraverunt patres nostri,speraverunt, et liberasti eos;
PS|22|6|ad te clamaverunt et salvi facti sunt,in te speraverunt et non sunt confusi.
PS|22|7|Ego autem sum vermis et non homo,opprobrium hominum et abiectio plebis.
PS|22|8|Omnes videntes me deriserunt me;torquentes labia moverunt caput:
PS|22|9|" Speravit in Domino: eripiat eum,salvum faciat eum, quoniam vult eum ".
PS|22|10|Quoniam tu es qui extraxisti me de ventre,spes mea ad ubera matris meae.
PS|22|11|In te proiectus sum ex utero,de ventre matris meae Deus meus es tu.
PS|22|12|Ne longe fias a me,quoniam tribulatio proxima est,quoniam non est qui adiuvet.
PS|22|13|Circumdederunt me vituli multi,tauri Basan obsederunt me.
PS|22|14|Aperuerunt super me os suumsicut leo rapiens et rugiens.
PS|22|15|Sicut aqua effusus sum,et dissoluta sunt omnia ossa mea.Factum est cor meum tamquam ceraliquescens in medio ventris mei.
PS|22|16|Aruit tamquam testa palatum meum,et lingua mea adhaesit faucibus meis,et in pulverem mortis deduxisti me.
PS|22|17|Quoniam circumdederunt me canes multi,concilium malignantium obsedit me.Foderunt manus meas et pedes meos,
PS|22|18|et dinumeravi omnia ossa mea.Ipsi vero consideraverunt et inspexerunt me;
PS|22|19|diviserunt sibi vestimenta meaet super vestem meam miserunt sortem.
PS|22|20|Tu autem, Domine, ne elongaveris;fortitudo mea, ad adiuvandum me festina.
PS|22|21|Erue a framea animam meamet de manu canis unicam meam.
PS|22|22|Salva me ex ore leoniset a cornibus unicornium humilitatem meam.
PS|22|23|Narrabo nomen tuum fratribus meis,in medio ecclesiae laudabo te.
PS|22|24|Qui timetis Dominum, laudate eum;universum semen Iacob, glorificate eum.Metuat eum omne semen Israel,
PS|22|25|quoniam non sprevit neque despexit afflictionem pauperisnec avertit faciem suam ab eoet, cum clamaret ad eum, exaudivit.
PS|22|26|Apud te laus mea in ecclesia magna; vota mea reddam in conspectu timentium eum.
PS|22|27|Edent pauperes et saturabuntur;et laudabunt Dominum, qui requirunt eum: Vivant corda eorum in saeculum saeculi! ".
PS|22|28|Reminiscentur et convertentur ad Dominumuniversi fines terrae,et adorabunt in conspectu eiusuniversae familiae gentium.
PS|22|29|Quoniam Domini est regnum,et ipse dominabitur gentium.
PS|22|30|Ipsum solum adorabunt omnes, qui dormiunt in terra;in conspectu eius procident omnes, qui descendunt in pulverem.Anima autem mea illi vivet,
PS|22|31|et semen meum serviet ipsi.Narrabitur de Domino generationi venturae;
PS|22|32|et annuntiabunt iustitiam eiuspopulo, qui nascetur: " Haec fecit Dominus! ".
PS|23|1|PSALMUS. David.Dominus pascit me, et nihil mihi deerit:
PS|23|2|in pascuis virentibus me collocavit,super aquas quietis eduxit me,
PS|23|3|animam meam refecit.Deduxit me super semitas iustitiae propter nomen suum.
PS|23|4|Nam et si ambulavero in valle umbrae mortis,non timebo mala, quoniam tu mecum es.Virga tua et baculus tuus,ipsa me consolata sunt.
PS|23|5|Parasti in conspectu meo mensamadversus eos, qui tribulant me;impinguasti in oleo caput meum,et calix meus redundat.
PS|23|6|Etenim benignitas et misericordia subsequentur meomnibus diebus vitae meae,et inhabitabo in domo Dominiin longitudinem dierum.
PS|24|1|David. PSALMUS.Domini est terra, et plenitudo eius,orbis terrarum, et qui habitant in eo.
PS|24|2|Quia ipse super maria fundavit eumet super flumina firmavit eum. -
PS|24|3|Quis ascendet in montem Domini,aut quis stabit in loco sancto eius?
PS|24|4|Innocens manibus et mundo corde,qui non levavit ad vana animam suamnec iuravit in dolum.
PS|24|5|Hic accipiet benedictionem a Dominoet iustificationem a Deo salutari suo.
PS|24|6|Haec est generatio quaerentium eum,quaerentium faciem Dei Iacob.
PS|24|7|Attollite, portae, capita vestra,et elevamini, portae aeternales,et introibit rex gloriae.
PS|24|8|Quis est iste rex gloriae?Dominus fortis et potens,Dominus potens in proelio.
PS|24|9|Attollite, portae, capita vestra,et elevamini, portae aeternales,et introibit rex gloriae.
PS|24|10|Quis est iste rex gloriae?Dominus virtutum ipse est rex gloriae.
PS|25|1|David.ALEPH. Ad te, Domine, levavi animam meam,
PS|25|2|BETH. Deus meus, in te confido; non erubescam.Neque exsultent super me inimici mei,
PS|25|3|GHIMEL. etenim universi, qui sustinent te, non confundentur.Confundantur infideliter agentes propter vanitatem.
PS|25|4|DALETH. Vias tuas, Domine, demonstra mihiet semitas tuas edoce me.
PS|25|5|HE. Dirige me in veritate tua et doce me,quia tu es Deus salutis meae,VAU. et te sustinui tota die.
PS|25|6|ZAIN. Reminiscere miserationum tuarum, Domine,et misericordiarum tuarum, quoniam a saeculo sunt.
PS|25|7|HETH. Peccata iuventutis meae et delicta mea ne memineris;secundum misericordiam tuam memento mei tu,propter bonitatem tuam, Domine.
PS|25|8|TETH. Dulcis et rectus Dominus,propter hoc peccatores viam docebit;
PS|25|9|IOD. diriget mansuetos in iudicio,docebit mites vias suas.
PS|25|10|CAPH. Universae viae Domini misericordia et veritascustodientibus testamentum eius et testimonia eius.
PS|25|11|LAMED. Propter nomen tuum, Domine,propitiaberis peccato meo: multum est enim.
PS|25|12|MEM. Quis est homo, qui timet Dominum?Docebit eum viam, quam eligat.
PS|25|13|NUN. Anima eius in bonis demorabitur,et semen eius hereditabit terram.
PS|25|14|SAMECH. Familiariter aget Dominus cum timentibus eum,ut testamentum suum manifestet illis.
PS|25|15|AIN. Oculi mei semper ad Dominum,quoniam ipse evellet de laqueo pedes meos.
PS|25|16|PHE. Respice in me et miserere mei,quia unicus et pauper sum ego.
PS|25|17|SADE. Dilata angustias cordis meiet de necessitatibus meis erue me.
PS|25|18|Vide humilitatem meam et laborem meumet dimitte universa delicta mea.
PS|25|19|RES. Respice inimicos meos, quoniam multiplicati suntet odio crudeli oderunt me.
PS|25|20|SIN. Custodi animam meam et erue me;non erubescam, quoniam speravi in te.
PS|25|21|TAU. Innocentia et aequitas custodiant me,quia sustinui te.
PS|25|22|PHE. Libera, Deus, Israelex omnibus tribulationibus suis.
PS|26|1|David.Iudica me, Domine, quoniam ego in innocentia mea ingressus sumet in Domino sperans non infirmabor.
PS|26|2|Proba me, Domine, et tenta me;ure renes meos et cor meum. -
PS|26|3|Quoniam misericordia tua ante oculos meos est,et ambulavi in veritate tua.
PS|26|4|Non sedi cum viris vanitatiset cum occulte agentibus non introibo.
PS|26|5|Odivi ecclesiam malignantiumet cum impiis non sedebo.
PS|26|6|Lavabo in innocentia manus measet circumdabo altare tuum, Domine,
PS|26|7|ut auditas faciam voces laudiset enarrem universa mirabilia tua.
PS|26|8|Domine, dilexi habitaculum domus tuaeet locum habitationis gloriae tuae.
PS|26|9|Ne colligas cum impiis animam meamet cum viris sanguinum vitam meam,
PS|26|10|in quorum manibus iniquitates sunt,dextera eorum repleta est muneribus.
PS|26|11|Ego autem in innocentia mea ingressus sum;redime me et miserere mei.
PS|26|12|Pes meus stetit in directo,in ecclesiis benedicam Domino.
PS|27|1|David.Dominus illuminatio mea et salus mea; quem timebo?Dominus protector vitae meae; a quo trepidabo?
PS|27|2|Dum appropiant super me nocentes,ut edant carnes meas;qui tribulant me et inimici mei,ipsi infirmati sunt et ceciderunt.
PS|27|3|Si consistant adversum me castra,non timebit cor meum;si exsurgat adversum me proelium, in hoc ego sperabo.
PS|27|4|Unum petii a Domino, hoc requiram:ut inhabitem in domo Dominiomnibus diebus vitae meae,ut videam voluptatem Dominiet visitem templum eius.
PS|27|5|Quoniam occultabit me in tentorio suoin die malorum.Abscondet me in abscondito tabernaculi sui,in petra exaltabit me.
PS|27|6|Et nunc exaltatur caput meumsuper inimicos meos in circuitu meo.Immolabo in tabernaculo eius hostias vociferationis,cantabo et psalmum dicam Domino.
PS|27|7|Exaudi, Domine, vocem meam, qua clamavi;miserere mei et exaudi me.
PS|27|8|De te dixit cor meum: " Exquirite faciem meam! ".Faciem tuam, Domine, exquiram.
PS|27|9|Ne avertas faciem tuam a me,ne declines in ira a servo tuo.Adiutor meus es tu, ne me reiciasneque derelinquas me, Deus salutis meae.
PS|27|10|Quoniam pater meus et mater mea dereliquerunt me,Dominus autem assumpsit me.
PS|27|11|Ostende mihi, Domine, viam tuamet dirige me in semitam rectam propter inimicos meos.
PS|27|12|Ne tradideris me in animam tribulantium me,quoniam insurrexerunt in me testes iniqui,et qui violentiam spirant.
PS|27|13|Credo videre bona Domini in terra viventium.
PS|27|14|Exspecta Dominum, viriliter age,et confortetur cor tuum, et sustine Dominum.
PS|28|1|David.Ad te, Domine, clamabo;Deus meus, ne sileas a me.Ne quando taceas a me,et assimilabor descendentibus in lacum.
PS|28|2|Exaudi vocem deprecationis meae, dum clamo ad te,dum extollo manus meas ad templum sanctum tuum.
PS|28|3|Ne simul trahas me cum peccatoribuset cum operantibus iniquitatem.Qui loquuntur pacem cum proximo suo,mala autem in cordibus eorum.
PS|28|4|Da illis secundum opera eorumet secundum nequitiam adinventionum ipsorum.Secundum opus manuum eorum tribue illis,redde retributionem eorum ipsis.
PS|28|5|Quoniam non intellexerunt opera Dominiet opus manuum eius,destruet illos et non aedificabit eos.
PS|28|6|Benedictus Dominus,quoniam exaudivit vocem deprecationis meae;
PS|28|7|Dominus adiutor meus et protector meus,in ipso speravit cor meum, et adiutus sum,et exsultavit cor meum,et in cantico meo confitebor ei.
PS|28|8|Dominus fortitudo plebi suae,et refugium salvationum christi sui est.
PS|28|9|Salvum fac populum tuum et benedic hereditati tuaeet pasce eos et extolle illos usque in aeternum.
PS|29|1|PSALMUS. David.Afferte Domino, filii Dei,afferte Domino gloriam et potentiam,
PS|29|2|afferte Domino gloriam nominis eius,adorate Dominum in splendore sancto.
PS|29|3|Vox Domini super aquas;Deus maiestatis intonuit,Dominus super aquas multas.
PS|29|4|Vox Domini in virtute,vox Domini in magnificentia.
PS|29|5|Vox Domini confringentis cedros;et confringet Dominus cedros Libani.
PS|29|6|Et saltare faciet, tamquam vitulum, Libanum,et Sarion, quemadmodum filium unicornium. -
PS|29|7|Vox Domini intercidentis flammam ignis,
PS|29|8|vox Domini concutientis desertum,et concutiet Dominus desertum Cades.
PS|29|9|Vox Domini properantis partum cervarum,et denudabit condensa;et in templo eius omnes dicent gloriam.
PS|29|10|Dominus super diluvium habitat,et sedebit Dominus rex in aeternum.
PS|29|11|Dominus virtutem populo suo dabit,Dominus benedicet populo suo in pace.
PS|30|1|PSALMUS. Canticum festi Dedicationis Templi. David.
PS|30|2|Exaltabo te, Domine, quoniam extraxisti menec delectasti inimicos meos super me.
PS|30|3|Domine Deus meus, clamavi ad te, et sanasti me.
PS|30|4|Domine, eduxisti ab inferno animam meam,vivificasti me, ut non descenderem in lacum.
PS|30|5|Psallite Domino, sancti eius,et confitemini memoriae sanctitatis eius,
PS|30|6|quoniam ad momentum indignatio eius,et per vitam voluntas eius.Ad vesperum demoratur fletus,ad matutinum laetitia.
PS|30|7|Ego autem dixi in securitate mea: Non movebor in aeternum ".
PS|30|8|Domine, in voluntate tuapraestitisti decori meo virtutem;avertisti faciem tuam a me,et factus sum conturbatus.
PS|30|9|Ad te, Domine, clamabamet ad Deum meum deprecabar.
PS|30|10|Quae utilitas in sanguine meo,dum descendo in corruptionem?Numquid confitebitur tibi pulvisaut annuntiabit veritatem tuam?
PS|30|11|Audivit Dominus et misertus est mei,Dominus factus est adiutor meus.
PS|30|12|Convertisti planctum meum in choros mihi,conscidisti saccum meum et accinxisti me laetitia,
PS|30|13|ut cantet tibi gloria mea et non taceat.Domine Deus meus, in aeternum confitebor tibi.
PS|31|1|Magistro chori. PSALMUS. David.
PS|31|2|In te, Domine, speravi, non confundar in aeternum;in iustitia tua libera me.
PS|31|3|Inclina ad me aurem tuam,accelera, ut eruas me.Esto mihi in rupem praesidiiet in domum munitam, ut salvum me facias.
PS|31|4|Quoniam fortitudo mea et refugium meum es tuet propter nomen tuum deduces me et pasces me.
PS|31|5|Educes me de laqueo, quem absconderunt mihi,quoniam tu es fortitudo mea.
PS|31|6|In manus tuas commendo spiritum meum;redemisti me, Domine, Deus veritatis.
PS|31|7|Odisti observantes vanitates supervacuas,ego autem in Domino speravi.
PS|31|8|Exsultabo et laetabor in misericordia tua,quoniam respexisti humilitatem meam;agnovisti necessitates animae meae
PS|31|9|nec conclusisti me in manibus inimici;statuisti in loco spatioso pedes meos.
PS|31|10|Miserere mei, Domine, quoniam tribulor;conturbatus est in maerore oculus meus,anima mea et venter meus.
PS|31|11|Quoniam defecit in dolore vita mea,et anni mei in gemitibus;infirmata est in paupertate virtus mea,et ossa mea contabuerunt.
PS|31|12|Apud omnes inimicos meos factus sum opprobriumet vicinis meis valde et timor notis meis:qui videbant me foras, fugiebant a me.
PS|31|13|Oblivioni a corde datus sum tamquam mortuus;factus sum tamquam vas perditum.
PS|31|14|Quoniam audivi vituperationem multorum: horror in circuitu;in eo dum convenirent simul adversum me,auferre animam meam consiliati sunt.
PS|31|15|Ego autem in te speravi, Domine;dixi: " Deus meus es tu,
PS|31|16|in manibus tuis sortes meae ".Eripe me de manu inimicorum meorumet a persequentibus me;
PS|31|17|illustra faciem tuam super servum tuum,salvum me fac in misericordia tua.
PS|31|18|Domine, non confundar, quoniam invocavi te;erubescant impii et obmutescant in inferno.
PS|31|19|Muta fiant labia dolosa,quae loquuntur adversus iustum protervain superbia et in abusione.
PS|31|20|Quam magna multitudo dulcedinis tuae, Domine,quam abscondisti timentibus te.Perfecisti eis, qui sperant in te,in conspectu filiorum hominum.
PS|31|21|Abscondes eos in abscondito faciei tuaea conturbatione hominum;proteges eos in tabernaculoa contradictione linguarum.
PS|31|22|Benedictus Dominus,quoniam mirificavit misericordiam suam mihi in civitate munita.
PS|31|23|Ego autem dixi in trepidatione mea: Praecisus sum a conspectu oculorum tuorum ".Verumtamen exaudisti vocem orationis meae,dum clamarem ad te.
PS|31|24|Diligite Dominum, omnes sancti eius:fideles conservat Dominuset retribuit abundanter facientibus superbiam.
PS|31|25|Viriliter agite, et confortetur cor vestrum,omnes, qui speratis in Domino.
PS|32|1|David. Maskil.Beatus, cui remissa est iniquitas,et obtectum est peccatum.
PS|32|2|Beatus vir, cui non imputavit Dominus delictum,nec est in spiritu eius dolus.
PS|32|3|Quoniam tacui, inveteraverunt ossa mea,dum rugirem tota die.
PS|32|4|Quoniam die ac nocte gravata est super me manus tua,immutatus est vigor meus in ardoribus aestatis.
PS|32|5|Peccatum meum cognitum tibi feciet delictum meum non abscondi.Dixi: " Confitebor adversum me iniquitatem meam Domino ".Et tu remisisti impietatem peccati mei.
PS|32|6|Propter hoc orabit ad te omnis sanctus in tempore opportuno.Et in diluvio aquarum multarumad eum non approximabunt.
PS|32|7|Tu es refugium meum, a tribulatione conservabis me;exsultationibus salutis circumdabis me.
PS|32|8|Intellectum tibi dabo et instruam te in via, qua gradieris;firmabo super te oculos meos.
PS|32|9|Nolite fieri sicut equus et mulus,quibus non est intellectus;in camo et freno si accedis ad constringendum,non approximant ad te.
PS|32|10|Multi dolores impii,sperantem autem in Domino misericordia circumdabit.
PS|32|11|Laetamini in Domino et exsultate, iusti;et gloriamini, omnes recti corde.
PS|33|1|Exsultate, iusti, in Domino;rectos decet collaudatio.
PS|33|2|Confitemini Domino in cithara,in psalterio decem chordarum psallite illi.
PS|33|3|Cantate ei canticum novum,bene psallite ei in vociferatione,
PS|33|4|quia rectum est verbum Domini,et omnia opera eius in fide.
PS|33|5|Diligit iustitiam et iudicium;misericordia Domini plena est terra.
PS|33|6|Verbo Domini caeli facti sunt,et spiritu oris eius omnis virtus eorum.
PS|33|7|Congregans sicut in utre aquas maris,ponens in thesauris abyssos.
PS|33|8|Timeat Dominum omnis terra,a facie autem eius formident omnes inhabitantes orbem.
PS|33|9|Quoniam ipse dixit, et facta sunt,ipse mandavit, et creata sunt.
PS|33|10|Dominus dissipat consilia gentium,irritas facit cogitationes populorum.
PS|33|11|Consilium autem Domini in aeternum manet,cogitationes cordis eius in generatione et generationem.
PS|33|12|Beata gens, cui Dominus est Deus,populus, quem elegit in hereditatem sibi.
PS|33|13|De caelo respexit Dominus,vidit omnes filios hominum.
PS|33|14|De loco habitaculi sui respexitsuper omnes, qui habitant terram,
PS|33|15|qui finxit singillatim corda eorum,qui intellegit omnia opera eorum.
PS|33|16|Non salvatur rex per multam virtutem,et gigas non liberabitur in multitudine virtutis suae.
PS|33|17|Fallax equus ad salutem,in abundantia autem virtutis suae non salvabit.
PS|33|18|Ecce oculi Domini super metuentes eum,in eos, qui sperant super misericordia eius,
PS|33|19|ut eruat a morte animas eorumet alat eos in fame.
PS|33|20|Anima nostra sustinet Dominum,quoniam adiutor et protector noster est;
PS|33|21|quia in eo laetabitur cor nostrum,et in nomine sancto eius speravimus.
PS|33|22|Fiat misericordia tua, Domine, super nos,quemadmodum speravimus in te.
PS|34|1|David, quando se mente alienatum simulavitcoram Abimelech et, ab illo dimissus, abiit.
PS|34|2|ALEPH. Benedicam Dominum in omni tempore,semper laus eius in ore meo.
PS|34|3|BETH. In Domino gloriabitur anima mea,audiant mansueti et laetentur.
PS|34|4|GHIMEL. Magnificate Dominum mecum,et exaltemus nomen eius in idipsum.
PS|34|5|DALETH. Exquisivi Dominum, et exaudivit meet ex omnibus terroribus meis eripuit me.
PS|34|6|HE. Respicite ad eum, et illuminamini,et facies vestrae non confundentur.
PS|34|7|ZAIN. Iste pauper clamavit, et Dominus exaudivit eumet de omnibus tribulationibus eius salvavit eum.
PS|34|8|HETH. Vallabit angelus Domini in circuitu timentes eumet eripiet eos.
PS|34|9|TETH. Gustate et videte quoniam suavis est Dominus;beatus vir, qui sperat in eo.
PS|34|10|IOD. Timete Dominum, sancti eius,quoniam non est inopia timentibus eum.
PS|34|11|CAPH. Divites eguerunt et esurierunt,inquirentes autem Dominum non deficient omni bono.
PS|34|12|LAMED. Venite, filii, audite me:timorem Domini docebo vos.
PS|34|13|MEM. Quis est homo, qui vult vitam,diligit dies, ut videat bonum? -
PS|34|14|NUN. Prohibe linguam tuam a malo,et labia tua, ne loquantur dolum.
PS|34|15|SAMECH. Diverte a malo et fac bonum,inquire pacem et persequere eam.
PS|34|16|AIN. Oculi Domini super iustos,et aures eius in clamorem eorum.
PS|34|17|PHE. Vultus autem Domini super facientes mala,ut perdat de terra memoriam eorum.
PS|34|18|SADE. Clamaverunt, et Dominus exaudivitet ex omnibus tribulationibus eorum liberavit eos.
PS|34|19|COPH. Iuxta est Dominus iis, qui contrito sunt corde,et confractos spiritu salvabit.
PS|34|20|RES. Multae tribulationes iustorum,et de omnibus his liberabit eos Dominus.
PS|34|21|SIN. Custodit omnia ossa eorum,unum ex his non conteretur.
PS|34|22|TAU. Interficiet peccatorem malitia;et, qui oderunt iustum, punientur.
PS|34|23|PHE. Redimet Dominus animas servorum suorum;et non punientur omnes, qui sperant in eo.
PS|35|1|David.Iudica, Domine, iudicantes me;impugna impugnantes me.
PS|35|2|Apprehende clipeum et scutumet exsurge in adiutorium mihi.
PS|35|3|Effunde frameam et securimadversus eos, qui persequuntur me.Dic animae meae: " Salus tua ego sum ".
PS|35|4|Confundantur et revereanturquaerentes animam meam;avertantur retrorsum et confundanturcogitantes mihi mala.
PS|35|5|Fiant tamquam pulvis ante ventum,et angelus Domini impellens eos;
PS|35|6|fiat via illorum tenebrae et lubricum,et angelus Domini persequens eos.
PS|35|7|Quoniam gratis absconderunt mihi laqueum suum,gratis foderunt foveam animae meae.
PS|35|8|Veniat illi calamitas, quam ignorat,et captio, quam abscondit, apprehendat eum,et in eandem calamitatem ipse cadat.
PS|35|9|Anima autem mea exsultabit in Dominoet delectabitur super salutari suo.
PS|35|10|Omnia ossa mea dicent: Domine, quis similis tibi?Eripiens inopem de manu fortiorum eius,egenum et pauperem a diripientibus eum ".
PS|35|11|Surgentes testes iniqui,quae ignorabam, interrogabant me;
PS|35|12|retribuebant mihi mala pro bonis,desolatio est animae meae.
PS|35|13|Ego autem, cum infirmarentur,induebar cilicio,humiliabam in ieiunio animam meam;et oratio mea in sinu meo convertebatur.
PS|35|14|Quasi pro proximo et quasi pro fratre meo ambulabam,quasi lugens matrem contristatus incurvabar.
PS|35|15|Cum autem vacillarem, laetati sunt et convenerunt;convenerunt contra me percutientes, et ignoravi.
PS|35|16|Diripuerunt et non desistebant;tentaverunt me, subsannaverunt me subsannatione,frenduerunt super me dentibus suis.
PS|35|17|Domine, quamdiu aspicies?Restitue animam meam a malignitate eorum,a leonibus unicam meam.
PS|35|18|Confitebor tibi in ecclesia magna,in populo multo laudabo te.
PS|35|19|Non supergaudeant mihi inimici mei mendaces,qui oderunt me gratis et annuunt oculis.
PS|35|20|Etenim non pacifice loquebanturet contra mansuetos terrae dolos cogitabant.
PS|35|21|Et dilataverunt super me os suum;dixerunt: " Euge, euge, viderunt oculi nostri ". -
PS|35|22|Vidisti, Domine, ne sileas;Domine, ne discedas a me.
PS|35|23|Exsurge et evigila ad iudicium meum,Deus meus et Dominus meus, ad causam meam.
PS|35|24|Iudica me secundum iustitiam tuam, Domine Deus meus,et non supergaudeant mihi.
PS|35|25|Non dicant in cordibus suis: Euge animae nostrae ";nec dicant: " Devoravimus eum ".
PS|35|26|Erubescant et revereantur simul, qui gratulantur malis meis;induantur confusione et reverentia, qui magna loquuntur super me
PS|35|27|Exsultent et laetentur, qui volunt iustitiam meam,et dicant semper: " Magnificetur Dominus,qui vult pacem servi sui ".
PS|35|28|Et lingua mea meditabitur iustitiam tuam,tota die laudem tuam.
PS|36|1|Magistro chori. David, servi Domini.
PS|36|2|Susurrat iniquitas ad impium in medio cordis eius;non est timor Dei ante oculos eius.
PS|36|3|Quoniam blanditur ipsi in conspectu eius,ut non inveniat iniquitatem suam et oderit.
PS|36|4|Verba oris eius iniquitas et dolus,desiit intellegere, ut bene ageret.
PS|36|5|Iniquitatem meditatus est in cubili suo,astitit omni viae non bonae,malitiam autem non odivit.
PS|36|6|Domine, in caelo misericordia tua,et veritas tua usque ad nubes;
PS|36|7|iustitia tua sicut montes Dei,iudicia tua abyssus multa:homines et iumenta salvabis, Domine.
PS|36|8|Quam pretiosa misericordia tua, Deus!Filii autem hominum in tegmine alarum tuarum sperabunt;
PS|36|9|inebriabuntur ab ubertate domus tuae,et torrente voluptatis tuae potabis eos.
PS|36|10|Quoniam apud te est fons vitae,et in lumine tuo videbimus lumen.
PS|36|11|Praetende misericordiam tuam scientibus teet iustitiam tuam his, qui recto sunt corde.
PS|36|12|Non veniat mihi pes superbiae,et manus peccatoris non moveat me.
PS|36|13|Ibi ceciderunt, qui operantur iniquitatem,expulsi sunt nec potuerunt stare.
PS|37|1|David.ALEPH. Noli aemulari in malignantibusneque zelaveris facientes iniquitatem,
PS|37|2|quoniam tamquam fenum velociter arescentet quemadmodum herba virens decident.
PS|37|3|BETH. Spera in Domino et fac bonitatem,et inhabitabis terram et pasceris in fide.
PS|37|4|Delectare in Domino,et dabit tibi petitiones cordis tui.
PS|37|5|GHIMEL. Committe Domino viam tuam et spera in eo,et ipse faciet;
PS|37|6|et educet quasi lumen iustitiam tuamet iudicium tuum tamquam meridiem.
PS|37|7|DALETH. Quiesce in Domino et exspecta eum;noli aemulari in eo, qui prosperatur in via sua,in homine, qui molitur insidias.
PS|37|8|HE. Desine ab ira et derelinque furorem,noli aemulari, quod vertit ad malum,
PS|37|9|quoniam qui malignantur, exterminabuntur,sustinentes autem Dominum ipsi hereditabunt terram.
PS|37|10|VAU. Et adhuc pusillum et non erit peccator,et quaeres locum eius et non invenies.
PS|37|11|Mansueti autem hereditabunt terramet delectabuntur in multitudine pacis.
PS|37|12|ZAIN. Insidiabitur peccator iustoet stridebit super eum dentibus suis.
PS|37|13|Dominus autem irridebit eum,quoniam prospicit quod veniet dies eius.
PS|37|14|HETH. Gladium evaginaverunt peccatores,intenderunt arcum suum,ut deiciant pauperem et inopem,ut trucident recte ambulantes in via.
PS|37|15|Gladius eorum intrabit in corda ipsorum,et arcus eorum confringetur.
PS|37|16|TETH. Melius est modicum iustosuper divitias peccatorum multas,
PS|37|17|quoniam brachia peccatorum conterentur,confirmat autem iustos Dominus.
PS|37|18|IOD. Novit Dominus dies immaculatorum,et hereditas eorum in aeternum erit.
PS|37|19|Non confundentur in tempore maloet in diebus famis saturabuntur.
PS|37|20|CAPH. Quia peccatores peribunt,inimici vero Domini ut decor camporum deficient,quemadmodum fumus deficient.
PS|37|21|LAMED. Mutuatur peccator et non solvet,iustus autem miseretur et tribuet.
PS|37|22|Quia benedicti eius hereditabunt terram,maledicti autem eius exterminabuntur.
PS|37|23|MEM. A Domino gressus hominis confirmantur,et viam eius volet.
PS|37|24|Cum ceciderit, non collidetur,quia Dominus sustentat manum eius.
PS|37|25|NUN. Iunior fui et senuiet non vidi iustum derelictumnec semen eius quaerens panem.
PS|37|26|Tota die miseretur et commodat,et semen illius in benedictione erit.
PS|37|27|SAMECH. Declina a malo et fac bonum,et inhabitabis in saeculum saeculi,
PS|37|28|quia Dominus amat iudiciumet non derelinquet sanctos suos.AIN. Iniusti in aeternum disperibunt,et semen impiorum exterminabitur.
PS|37|29|Iusti autem hereditabunt terramet inhabitabunt in saeculum saeculi super eam.
PS|37|30|PHE. Os iusti meditabitur sapientiam,et lingua eius loquetur iudicium;
PS|37|31|lex Dei eius in corde ipsius,et non vacillabunt gressus eius.
PS|37|32|SADE. Considerat peccator iustumet quaerit mortificare eum;
PS|37|33|Dominus autem non derelinquet eum in manibus eiusnec damnabit eum, cum iudicabitur illi.
PS|37|34|COPH. Exspecta Dominum et custodi viam eius,et exaltabit te, ut hereditate capias terram;cum exterminabuntur peccatores, videbis.
PS|37|35|RES. Vidi impium superexaltatumet elevatum sicut cedrum virentem;
PS|37|36|et transivi, et ecce non erat,et quaesivi eum, et non est inventus.
PS|37|37|SIN. Observa innocentiam et vide aequitatem,quoniam est posteritas homini pacifico.
PS|37|38|Iniusti autem disperibunt simul,posteritas impiorum exterminabitur.
PS|37|39|TAU. Salus autem iustorum a Domino,et protector eorum in tempore tribulationis.
PS|37|40|Et adiuvabit eos Dominus et liberabit eoset eruet eos a peccatoribus et salvabit eos,quia speraverunt in eo.
PS|38|1|PSALMUS. David. Ad commemorandum.
PS|38|2|Domine, ne in furore tuo arguas meneque in ira tua corripias me,
PS|38|3|quoniam sagittae tuae infixae sunt mihi,et descendit super me manus tua.
PS|38|4|Non est sanitas in carne mea a facie indignationis tuae,non est pax ossibus meis a facie peccatorum meorum.
PS|38|5|Quoniam iniquitates meae supergressae sunt caput meumet sicut onus grave gravant me nimis. -
PS|38|6|Putruerunt et corrupti sunt livores meia facie insipientiae meae.
PS|38|7|Inclinatus sum et incurvatus nimis;tota die contristatus ingrediebar.
PS|38|8|Quoniam lumbi mei impleti sunt ardoribus,et non est sanitas in carne mea.
PS|38|9|Afflictus sum et humiliatus sum nimis,rugiebam a gemitu cordis mei.
PS|38|10|Domine, ante te omne desiderium meum,et gemitus meus a te non est absconditus.
PS|38|11|Palpitavit cor meum, dereliquit me virtus mea,et lumen oculorum meorum, et ipsum non est mecum.
PS|38|12|Amici mei et proximi meiprocul a plaga mea steterunt,et propinqui mei de longe steterunt.
PS|38|13|Et laqueos posuerunt, qui quaerebant animam meam;et, qui requirebant mala mihi, locuti sunt insidiaset dolos tota die meditabantur.
PS|38|14|Ego autem tamquam surdus non audiebamet sicut mutus non aperiens os suum;
PS|38|15|et factus sum sicut homo non audienset non habens in ore suo redargutiones.
PS|38|16|Quoniam in te, Domine, speravi,tu exaudies, Domine Deus meus.
PS|38|17|Quia dixi: "Ne quando supergaudeant mihi;dum commoventur pedes mei,magnificantur super me ".
PS|38|18|Quoniam ego in lapsum paratus sum,et dolor meus in conspectu meo semper.
PS|38|19|Quoniam iniquitatem meam annuntiaboet sollicitus sum de peccato meo.
PS|38|20|Inimici autem mei vivunt et confirmati sunt;et multiplicati sunt, qui oderunt me inique.
PS|38|21|Retribuentes mala pro bonis detrahebant mihi,pro eo quod sequebar bonitatem.
PS|38|22|Ne derelinquas me, Domine;Deus meus, ne discesseris a me.
PS|38|23|Festina in adiutorium meum,Domine, salus mea.
PS|39|1|Magistro chori, Idithun. PSALMUS. David.
PS|39|2|Dixi: " Custodiam vias meas,ut non delinquam in lingua mea;ponam ori meo custodiam,donec consistit peccator adversum me ".
PS|39|3|Tacens obmutui et silui absque ullo bono,et dolor meus renovatus est.
PS|39|4|Concaluit cor meum intra me,et in meditatione mea exarsit ignis.
PS|39|5|Locutus sum in lingua mea: Notum fac mihi, Domine, finem meum;et numerum dierum meorum quis est,ut sciam quam brevis sit vita mea ".
PS|39|6|Ecce paucorum palmorum fecisti dies meos,et spatium vitae meae tamquam nihilum ante te.Etenim universa vanitas omnis homo constitutus est.
PS|39|7|Etenim ut imago pertransit homo.Etenim vanitas est et concitatur;thesaurizat et ignorat quis congregabit ea.
PS|39|8|Et nunc quae est exspectatio mea, Domine?Spes mea apud te est.
PS|39|9|Ab omnibus iniquitatibus meis erue me,opprobrium insipienti ne ponas me.
PS|39|10|Obmutui et non aperiam os meum,quoniam tu fecisti.
PS|39|11|Amove a me plagas tuas:ab ictu manus tuae ego defeci.
PS|39|12|In increpationibus, propter iniquitatem, corripuisti hominem,et tabescere fecisti, sicut tinea, desiderabilia eius.Etenim vanitas omnis homo.
PS|39|13|Exaudi orationem meam, Domine,et clamorem meum auribus percipe.Ad lacrimas meas ne obsurdescas,quoniam advena ego sum apud te,peregrinus sicut omnes patres mei.
PS|39|14|Avertere a me, ut refrigerer,priusquam abeam et non sim amplius.
PS|40|1|Magistro chori. David. PSALMUS.
PS|40|2|Exspectans exspectavi Dominum,et intendit mihi.
PS|40|3|Et exaudivit clamorem meumet eduxit me de lacu miseriae et de luto faecis;et statuit super petram pedes meoset firmavit gressus meos.
PS|40|4|Et immisit in os meum canticum novum,carmen Deo nostro.Videbunt multi et timebuntet sperabunt in Domino.
PS|40|5|Beatus vir, qui posuit Dominum spem suamet non respexit superbos et declinantes in mendacium.
PS|40|6|Multa fecisti tu, Domine Deus meus, mirabilia tua,et cogitationes tuas pro nobis: non est qui similis sit tibi.Si nuntiare et eloqui voluero,multiplicabuntur super numerum.
PS|40|7|Sacrificium et oblationem noluisti,aures autem fodisti mihi.Holocaustum et pro peccato non postulasti,
PS|40|8|tunc dixi: " Ecce venio.In volumine libri scriptum est de me.
PS|40|9|Facere voluntatem tuam,Deus meus, volui;et lex tua in praecordiis meis ".
PS|40|10|Annuntiavi iustitiam tuam in ecclesia magna;ecce labia mea non prohibebo, Domine, tu scisti.
PS|40|11|Iustitiam tuam non abscondi in corde meo,veritatem tuam et salutare tuum dixi.Non abscondi misericordiam tuamet veritatem tuam ab ecclesia magna.
PS|40|12|Tu autem, Domine, ne prohibeas miserationes tuas a me;misericordia tua et veritas tua semper suscipiant me,
PS|40|13|quoniam circumdederunt me mala, quorum non est numerus;comprehenderunt me iniquitates meae,et non potui videre.Multiplicatae sunt super capillos capitis mei,et cor meum dereliquit me.
PS|40|14|Complaceat tibi, Domine, ut eruas me;Domine, ad adiuvandum me festina.
PS|40|15|Confundantur et revereantur simul,qui quaerunt animam meam, ut auferant eam.Avertantur retrorsum et erubescant,qui volunt mihi mala.
PS|40|16|Obstupescant propter confusionem suam,qui dicunt mihi: " Euge, euge ".
PS|40|17|Exsultent et laetentur in te omnes quaerentes te;et dicant semper: " Magnificetur Dominus ",qui diligunt salutare tuum.
PS|40|18|Ego autem egenus et pauper sum;Dominus sollicitus est mei.Adiutor meus et liberator meus tu es;Deus meus, ne tardaveris.
PS|41|1|Magistro chori. PSALMUS. David.
PS|41|2|Beatus, qui intellegit de egeno;in die mala liberabit eum Dominus.
PS|41|3|Dominus servabit eum et vivificabit eumet beatum faciet eum in terraet non tradet eum in animam inimicorum eius.
PS|41|4|Dominus opem feret illi super lectum doloris eius;universum stratum eius versabis in infirmitate eius.
PS|41|5|Ego dixi: " Domine, miserere mei;sana animam meam, quia peccavi tibi ".
PS|41|6|Inimici mei dixerunt mala mihi: Quando morietur, et peribit nomen eius? ".
PS|41|7|Et si ingrediebatur, ut visitaret, vana loquebatur;cor eius congregabat iniquitatem sibi,egrediebatur foras et detrahebat.
PS|41|8|Simul adversum me susurrabant omnes inimici mei;adversum me cogitabant mala mihi:
PS|41|9|" Maleficium effusum est in eo;et, qui decumbit, non adiciet ut resurgat ".
PS|41|10|Sed et homo pacis meae, in quo speravi,qui edebat panem meum, levavit contra me calcaneum.
PS|41|11|Tu autem, Domine, miserere meiet resuscita me, et retribuam eis.
PS|41|12|In hoc cognovi quoniam voluisti me,quia non gaudebit inimicus meus super me;
PS|41|13|me autem propter innocentiam suscepistiet statuisti me in conspectu tuo in aeternum.
PS|41|14|Benedictus Dominus, Deus Israel,a saeculo et usque in saeculum. Fiat, fiat.
PS|42|1|Magistro chori. Maskil. Filiorum Core.
PS|42|2|Quemadmodum desiderat cervus ad fontes aquarum,ita desiderat anima mea ad te, Deus.
PS|42|3|Sitivit anima mea ad Deum, Deum vivum;quando veniam et apparebo ante faciem Dei?
PS|42|4|Fuerunt mihi lacrimae meae panis die ac nocte,dum dicitur mihi cotidie: " Ubi est Deus tuus? ".
PS|42|5|Haec recordatus sum et effudi in me animam meam;quoniam transibam in locum tabernaculi admirabilisusque ad domum Deiin voce exsultationis et confessionismultitudinis festa celebrantis.
PS|42|6|Quare tristis es, anima mea, et quare conturbaris in me?Spera in Deo, quoniam adhuc confitebor illi,salutare vultus mei et Deus meus.
PS|42|7|In meipso anima mea contristata est;propterea memor ero tuide terra Iordanis et Hermonim, de monte Misar.
PS|42|8|Abyssus abyssum invocat in voce cataractarum tuarum;omnes gurgites tui et fluctus tui super me transierunt.
PS|42|9|In die mandavit Dominus misericordiam suam,et nocte canticum eius apud me est: oratio ad Deum vitae meae.
PS|42|10|Dicam Deo: " Susceptor meus es.Quare oblitus es mei,et quare contristatus incedo,dum affligit me inimicus? ".
PS|42|11|Dum confringuntur ossa mea,exprobraverunt mihi, qui tribulant me,dum dicunt mihi quotidie: " Ubi est Deus tuus? ". -
PS|42|12|Quare tristis es, anima mea, et quare conturbaris in me?Spera in Deo, quoniam adhuc confitebor illi,salutare vultus mei et Deus meus.
PS|43|1|Iudica me, Deus, et discerne causam meam de gente non sancta;ab homine iniquo et doloso erue me.
PS|43|2|Quia tu es Deus refugii mei;quare me reppulisti,et quare tristis incedo, dum affligit me inimicus?
PS|43|3|Emitte lucem tuam et veritatem tuam;ipsae me deducant et adducantin montem sanctum tuum et in tabernacula tua.
PS|43|4|Et introibo ad altare Dei,ad Deum laetitiae exsultationis meae.Confitebor tibi in cithara, Deus, Deus meus.
PS|43|5|Quare tristis es, anima mea, et quare conturbaris in me?Spera in Deo, quoniam adhuc confitebor illi,salutare vultus mei et Deus meus.
PS|44|1|Magistro chori. Filiorum Core. Maskil.
PS|44|2|Deus, auribus nostris audivimus;patres nostri annuntiaverunt nobisopus, quod operatus es in diebus eorum, in diebus antiquis.
PS|44|3|Tu manu tua gentes depulisti et plantasti illos,afflixisti populos et dilatasti eos.
PS|44|4|Nec enim in gladio suo possederunt terram,et brachium eorum non salvavit eos;sed dextera tua et brachium tuumet illuminatio vultus tui,quoniam complacuisti in eis.
PS|44|5|Tu es rex meus et Deus meus,qui mandas salutes Iacob.
PS|44|6|In te inimicos nostros proiecimus,et in nomine tuo conculcavimus insurgentes in nos. -
PS|44|7|Non enim in arcu meo sperabo,et gladius meus non salvabit me.
PS|44|8|Tu autem salvasti nos de affligentibus noset odientes nos confudisti.
PS|44|9|In Deo gloriabimur tota dieet in nomine tuo confitebimur in saeculum.
PS|44|10|Nunc autem reppulisti et confudisti noset non egredieris, Deus, cum virtutibus nostris.
PS|44|11|Convertisti nos retrorsum coram inimicis nostris;et, qui oderunt nos, diripuerunt sibi.
PS|44|12|Dedisti nos tamquam oves ad vescendumet in gentibus dispersisti nos.
PS|44|13|Vendidisti populum tuum sine lucronec ditior factus es in commutatione eorum.
PS|44|14|Posuisti nos opprobrium vicinis nostris,subsannationem et derisum his, qui sunt in circuitu nostro.
PS|44|15|Posuisti nos similitudinem in gentibus,commotionem capitis in populis.
PS|44|16|Tota die verecundia mea contra me est,et confusio faciei meae cooperuit me
PS|44|17|a voce exprobrantis et obloquentis,a facie inimici et ultoris.
PS|44|18|Haec omnia venerunt super nos, nec obliti sumus teet inique non egimus in testamentum tuum.
PS|44|19|Et non recessit retro cor nostrum,nec declinaverunt gressus nostri a via tua;
PS|44|20|sed humiliasti nos in loco vulpiumet operuisti nos umbra mortis.
PS|44|21|Si obliti fuerimus nomen Dei nostriet si expanderimus manus nostras ad deum alienum,
PS|44|22|nonne Deus requiret ista?Ipse enim novit abscondita cordis.
PS|44|23|Quoniam propter te mortificamur tota die,aestimati sumus sicut oves occisionis.
PS|44|24|Evigila, quare obdormis, Domine?Exsurge et ne repellas in finem.
PS|44|25|Quare faciem tuam avertis,oblivisceris inopiae nostrae et tribulationis nostrae?
PS|44|26|Quoniam humiliata est in pulvere anima nostra,conglutinatus est in terra venter noster.Exsurge, Domine, adiuva noset redime nos propter misericordiam tuam.
PS|45|1|Magistro chori. Secundum " Lilia... ". Filiorum Core.Maskil. Canticum amoris.
PS|45|2|Eructavit cor meum verbum bonum,dico ego opera mea regi.Lingua mea calamus scribae velociter scribentis.
PS|45|3|Speciosus forma es prae filiis hominum,diffusa est gratia in labiis tuis,propterea benedixit te Deus in aeternum.
PS|45|4|Accingere gladio tuo super femur tuum, potentissime,magnificentia tua et ornatu tuo.
PS|45|5|Et ornatu tuo procede, currum ascendepropter veritatem et mansuetudinem et iustitiam.Et doceat te mirabilia dextera tua:
PS|45|6|sagittae tuae acutae populi sub te cadent -in corda inimicorum regis.
PS|45|7|Sedes tua, Deus, in saeculum saeculi;sceptrum aequitatis sceptrum regni tui.
PS|45|8|Dilexisti iustitiam et odisti iniquitatem,propterea unxit te Deus, Deus tuus, oleo laetitiae prae consortibus tuis.
PS|45|9|Myrrha et aloe et casia omnia vestimenta tua;e domibus eburneis chordae delectant te.
PS|45|10|Filiae regum in pretiosis tuis;astitit regina a dextris tuis ornata auro ex Ophir. -
PS|45|11|Audi, filia, et vide et inclina aurem tuamet obliviscere populum tuum et domum patris tui;
PS|45|12|et concupiscet rex speciem tuam.Quoniam ipse est dominus tuus, et adora eum.
PS|45|13|Filia Tyri cum muneribus;vultum tuum deprecabuntur divites plebis.
PS|45|14|Gloriosa nimis filia regis intrinsecus,texturis aureis circumamicta.
PS|45|15|In vestibus variegatis adducetur regi;virgines post eam, proximae eius, afferuntur tibi.
PS|45|16|Afferuntur in laetitia et exsultatione,adducuntur in domum regis.
PS|45|17|Pro patribus tuis erunt tibi filii;constitues eos principes super omnem terram.
PS|45|18|Memor ero nominis tuiin omni generatione et generatione;propterea populi confitebuntur tibi in aeternumet in saeculum saeculi.
PS|46|1|Magistro chori. Filiorum Core. Secundum " Virgines... ". Canticum.
PS|46|2|Deus est nobis refugium et virtus,adiutorium in tribulationibus inventus est nimis.
PS|46|3|Propterea non timebimus, dum turbabitur terra,et transferentur montes in cor maris.
PS|46|4|Fremant et intumescant aquae eius, conturbentur montes in elatione eius.
PS|46|5|Fluminis rivi laetificant civitatem Dei,sancta tabernacula Altissimi.
PS|46|6|Deus in medio eius, non commovebitur;adiuvabit eam Deus mane diluculo.
PS|46|7|Fremuerunt gentes, commota sunt regna;dedit vocem suam, liquefacta est terra.
PS|46|8|Dominus virtutum nobiscum,refugium nobis Deus Iacob.
PS|46|9|Venite et videte opera Domini,quae posuit prodigia super terram.Auferet bella usque ad finem terrae,
PS|46|10|arcum conteret et confringet armaet scuta comburet igne.
PS|46|11|Vacate et videte quoniam ego sum Deus:exaltabor in gentibus et exaltabor in terra.
PS|46|12|Dominus virtutum nobiscum,refugium nobis Deus Iacob.
PS|47|1|Magistro chori. Filiorum Core. PSALMUS.
PS|47|2|Omnes gentes, plaudite manibus,iubilate Deo in voce exsultationis,
PS|47|3|quoniam Dominus Altissimus, terribilis,rex magnus super omnem terram.
PS|47|4|Subiecit populos nobiset gentes sub pedibus nostris.
PS|47|5|Elegit nobis hereditatem nostram,gloriam Iacob, quem dilexit.
PS|47|6|Ascendit Deus in iubilo,et Dominus in voce tubae.
PS|47|7|Psallite Deo, psallite;psallite regi nostro, psallite.
PS|47|8|Quoniam rex omnis terrae Deus,psallite sapienter.
PS|47|9|Regnavit Deus super gentes,Deus sedet super sedem sanctam suam.
PS|47|10|Principes populorum congregati suntcum populo Dei Abraham,quoniam Dei sunt scuta terrae:vehementer elevatus est.
PS|48|1|Canticum. PSALMUS. Filiorum Core.
PS|48|2|Magnus Dominus et laudabilis nimisin civitate Dei nostri.
PS|48|3|Mons sanctus eius collis speciosus,exsultatio universae terrae.Mons Sion, extrema aquilonis,civitas regis magni.
PS|48|4|Deus in domibus eius notusfactus est ut refugium.
PS|48|5|Quoniam ecce reges congregati sunt,convenerunt in unum.
PS|48|6|Ipsi cum viderunt, sic admirati sunt,conturbati sunt, diffugerunt;
PS|48|7|illic tremor apprehendit eos,dolores ut parturientis.
PS|48|8|In spiritu orientisconteres naves Tharsis.
PS|48|9|Sicut audivimus, sic vidimusin civitate Domini virtutum,in civitate Dei nostri;Deus fundavit eam in aeternum.
PS|48|10|Recogitamus, Deus, misericordiam tuamin medio templi tui.
PS|48|11|Secundum nomen tuum, Deus,sic et laus tua in fines terrae;iustitia plena est dextera tua.
PS|48|12|Laetetur mons Sion, et exsultent filiae Iudaepropter iudicia tua.
PS|48|13|Circumdate Sion et complectimini eam,numerate turres eius.
PS|48|14|Ponite corda vestra in virtute eiuset percurrite domos eius,ut enarretis in progenie altera.
PS|48|15|Quoniam hic est Deus, Deus nosterin aeternum et in saeculum saeculi;ipse ducet nos in saecula.
PS|49|1|Magistro chori. Filiorum Core. PSALMUS.
PS|49|2|Audite haec, omnes gentes;auribus percipite, omnes, qui habitatis orbem:
PS|49|3|quique humiles et viri nobiles,simul in unum dives et pauper!
PS|49|4|Os meum loquetur sapientiam,et meditatio cordis mei prudentiam.
PS|49|5|Inclinabo in parabolam aurem meam,aperiam in psalterio aenigma meum.
PS|49|6|Cur timebo in diebus malis,cum iniquitas supplantantium circumdabit me?
PS|49|7|Qui confidunt in virtute suaet in multitudine divitiarum suarum gloriantur.
PS|49|8|Etenim seipsum non redimet homo;non dabit Deo propitiationem suam.
PS|49|9|Nimium est pretium redemptionis animae eius:ad ultimum deficiet,
PS|49|10|ut vivat usque in finem nec videat interitum.
PS|49|11|Et videbit sapientes morientes;simul insipiens et stultus peribuntet relinquent alienis divitias suas.
PS|49|12|Sepulcra eorum domus illorum in aeternum;tabernacula eorum in progeniem et progeniem,etsi vocaverunt nominibus suis terras suas.
PS|49|13|Et homo, cum sit in honore, non permanebit;comparatus est iumentis, quae pereunt,et similis factus est illis.
PS|49|14|Haec via illorum, quorum fiducia in semetipsis,et finis eorum, qui complacent in ore suo.
PS|49|15|Sicut oves in inferno positi sunt,mors depascet eos;descendent praecipites ad sepulcrum,et figura eorum erit in consumptionem:infernus habitaculum eorum.
PS|49|16|Verumtamen Deus redimet animam meam,de manu inferi vere suscipiet me.
PS|49|17|Ne timueris, cum dives factus fuerit homo,et cum multiplicata fuerit gloria domus eius,
PS|49|18|quoniam, cum interierit, non sumet omnia,neque descendet cum eo gloria eius.
PS|49|19|Cum animae suae in vita ipsius benedixerit: Laudabunt te quod benefecisti tibi ",
PS|49|20|tamen introibit ad progeniem patrum suorum,qui in aeternum non videbunt lumen.
PS|49|21|Homo, cum in honore esset, non intellexit;comparatus est iumentis, quae pereunt,et similis factus est illis.
PS|50|1|PSALMUS. Asaph.Deus deorum, Dominus, locutus estet vocavit terram a solis ortu usque ad occasum.
PS|50|2|Ex Sion speciosa decore Deus illuxit,
PS|50|3|Deus noster veniet et non silebit:ignis consumens est in conspectu eius,et in circuitu eius tempestas valida.
PS|50|4|Advocabit caelum desursumet terram discernere populum suum:
PS|50|5|" Congregate mihi sanctos meos,qui disposuerunt testamentum meum in sacrificio ".
PS|50|6|Et annuntiabunt caeli iustitiam eius,quoniam Deus iudex est.
PS|50|7|" Audi, populus meus, et loquar,Israel, et testificabor adversum te:Deus, Deus tuus, ego sum.
PS|50|8|Non in sacrificiis tuis arguam te;holocausta enim tua in conspectu meo sunt semper.
PS|50|9|Non accipiam de domo tua vitulosneque de gregibus tuis hircos.
PS|50|10|Quoniam meae sunt omnes ferae silvarum,iumentorum mille in montibus.
PS|50|11|Cognovi omnia volatilia caeli;et, quod movetur in agro, meum est.
PS|50|12|Si esuriero non dicam tibi;meus est enim orbis terrae et plenitudo eius.
PS|50|13|Numquid manducabo carnes taurorumaut sanguinem hircorum potabo?
PS|50|14|Immola Deo sacrificium laudiset redde Altissimo vota tua;
PS|50|15|et invoca me in die tribulationis:eruam te, et honorificabis me ".
PS|50|16|Peccatori autem dixit Deus: Quare tu enarras praecepta meaet assumis testamentum meum in os tuum?
PS|50|17|Tu vero odisti disciplinamet proiecisti sermones meos retrorsum.
PS|50|18|Si videbas furem, currebas cum eo;et cum adulteris erat portio tua.
PS|50|19|Os tuum dimittebas ad malitiam,et lingua tua concinnabat dolos.
PS|50|20|Sedens adversus fratrem tuum loquebariset adversus filium matris tuae proferebas opprobrium.
PS|50|21|Haec fecisti, et tacui.Existimasti quod eram tui similis.Arguam te et statuam illa contra faciem tuam.
PS|50|22|Intellegite haec, qui obliviscimini Deum,ne quando rapiam, et non sit qui eripiat.
PS|50|23|Qui immolabit sacrificium laudis, honorificabit me;et, qui immaculatus est in via, ostendam illi salutare Dei ".
PS|51|1|Magistro chori. PSALMUS. David,
PS|51|2|cum venit ad eum Nathan propheta,postquam cum Bethsabee peccavit.
PS|51|3|Miserere mei, Deus, secundum misericordiam tuam;et secundum multitudinem miserationum tuarumdele iniquitatem meam.
PS|51|4|Amplius lava me ab iniquitate meaet a peccato meo munda me.
PS|51|5|Quoniam iniquitatem meam ego cognosco,et peccatum meum contra me est semper.
PS|51|6|Tibi, tibi soli peccavi et malum coram te feci,ut iustus inveniaris in sententia tua et aequus in iudicio tuo.
PS|51|7|Ecce enim in iniquitate generatus sum,et in peccato concepit me mater mea.
PS|51|8|Ecce enim veritatem in corde dilexistiet in occulto sapientiam manifestasti mihi.
PS|51|9|Asperges me hyssopo, et mundabor;lavabis me, et super nivem dealbabor.
PS|51|10|Audire me facies gaudium et laetitiam,et exsultabunt ossa, quae contrivisti.
PS|51|11|Averte faciem tuam a peccatis meiset omnes iniquitates meas dele.
PS|51|12|Cor mundum crea in me, Deus,et spiritum firmum innova in visceribus meis.
PS|51|13|Ne proicias me a facie tuaet spiritum sanctum tuum ne auferas a me.
PS|51|14|Redde mihi laetitiam salutaris tuiet spiritu promptissimo confirma me.
PS|51|15|Docebo iniquos vias tuas,et impii ad te convertentur.
PS|51|16|Libera me de sanguinibus, Deus, Deus salutis meae,et exsultabit lingua mea iustitiam tuam.
PS|51|17|Domine, labia mea aperies,et os meum annuntiabit laudem tuam.
PS|51|18|Non enim sacrificio delectaris;holocaustum, si offeram, non placebit.
PS|51|19|Sacrificium Deo spiritus contribulatus;cor contritum et humiliatum, Deus, non despicies.
PS|51|20|Benigne fac, Domine, in bona voluntate tua Sion,ut aedificentur muri Ierusalem.
PS|51|21|Tunc acceptabis sacrificium iustitiae, oblationes et holocausta;tunc imponent super altare tuum vitulos.
PS|52|1|Magistro chori. Maskil. David,
PS|52|2|postquam Doeg Edomita ad Saul veniteique narravit dicens: David intravit in domum Abimelech ".
PS|52|3|Quid gloriaris in malitia,qui potens es iniquitate?
PS|52|4|Tota die insidias cogitasti;lingua tua sicut novacula acuta, qui facis dolum.
PS|52|5|Dilexisti malitiam super benignitatem,mendacium magis quam loqui aequitatem.
PS|52|6|Dilexisti omnia verba perditionis, lingua dolosa.
PS|52|7|Propterea Deus destruet te in finem;evellet te et emigrabit te de tabernaculoet radicem tuam de terra viventium.
PS|52|8|Videbunt iusti et timebuntet super eum ridebunt:
PS|52|9|" Ecce homo, qui non posuit Deum refugium suum,sed speravit in multitudine divitiarum suarumet praevaluit in insidiis suis ".
PS|52|10|Ego autem sicut virens oliva in domo Dei.Speravi in misericordia Deiin aeternum et in saeculum saeculi.
PS|52|11|Confitebor tibi in saeculum, quia fecisti;et exspectabo nomen tuum,quoniam bonum est, in conspectu sanctorum tuorum.
PS|53|1|Magistro chori. Secundum " Mahalat ". Maskil. David.Dixit insipiens in corde suo: " Non est Deus ".
PS|53|2|Corrupti sunt et abominationes operati sunt;non est qui faciat bonum.
PS|53|3|Deus de caelo prospexit super filios hominum,ut videat si est intellegens, aut requirens Deum.
PS|53|4|Omnes declinaverunt, simul corrupti sunt;non est qui faciat bonum, non est usque ad unum.
PS|53|5|Nonne scient omnes, qui operantur iniquitatem,qui devorant plebem meam ut cibum panis?Deum non invocaverunt;
PS|53|6|illic trepidaverunt timore, et non erat timor.Quoniam Deus dissipavit ossa eorum, qui te obsidebant,confusi sunt, quoniam Deus sprevit eos. -
PS|53|7|Quis dabit ex Sion salutare Israel?Cum converterit Deus captivitatem plebis suae,exsultabit Iacob, et laetabitur Israel.
PS|54|1|Magistro chori. Fidibus. Maskil. David,
PS|54|2|postquam Ziphaei ad Saul venerunt dicentes: Ecce David apud nos abditus latet ".
PS|54|3|Deus, in nomine tuo salvum me facet in virtute tua iudica me.
PS|54|4|Deus, exaudi orationem meam,auribus percipe verba oris mei!
PS|54|5|Quoniam superbi insurrexerunt adversum me,et fortes quaesierunt animam meamet non proposuerunt Deum ante conspectum suum.
PS|54|6|Ecce enim Deus adiuvat me,et Dominus susceptor est animae meae.
PS|54|7|Converte mala super inimicos meos et in veritate tua disperde illos.
PS|54|8|Voluntarie sacrificabo tibi,confitebor nomini tuo, Domine, quoniam bonum est;
PS|54|9|quoniam ex omni tribulatione eripuit me,et super inimicos meos despexit oculus meus.
PS|55|1|Magistro chori. Fidibus. Maskil. David.
PS|55|2|Auribus percipe, Deus, orationem meamet ne abscondaris a deprecatione mea;
PS|55|3|intende mihi et exaudi me.Excussus sum in meditatione mea et conturbatus sum
PS|55|4|a voce inimici et a tribulatione peccatoris.Quoniam devolverunt in me iniquitatemet in ira molesti erant mihi.
PS|55|5|Cor meum torquetur intra me,et formido mortis cecidit super me.
PS|55|6|Timor et tremor venerunt super me, et contexit me pavor. -
PS|55|7|Et dixi: " Quis dabit mihi pennas sicut columbae,et volabo et requiescam?
PS|55|8|Ecce elongabo fugienset manebo in solitudine.
PS|55|9|Exspectabo eum, qui salvum me faciata spiritu procellae et tempestate ".
PS|55|10|Dissipa, Domine, divide linguas eorum,quoniam vidi violentiam et contentionem in civitate.
PS|55|11|Die ac nocte circumeunt eam super muros eius,
PS|55|12|iniquitas et labor et insidiae in medio eius;et non defecit de plateis eius fraudulentia et dolus.
PS|55|13|Quoniam si inimicus meus maledixisset mihi,sustinuissem utique;et si is qui oderat me, super me magnificatus fuisset,abscondissem me forsitan ab eo.
PS|55|14|Tu vero, homo coaequalis meus,familiaris meus et notus meus,
PS|55|15|qui simul habuimus dulce consortium:in domo Dei ambulavimus in concursu.
PS|55|16|Veniat mors super illos,et descendant in infernum viventes,quoniam nequitiae in habitaculis eorum,in medio eorum.
PS|55|17|Ego autem ad Deum clamabo,et Dominus salvabit me.
PS|55|18|Vespere et mane et meridie meditabor et ingemiscam,et exaudiet vocem meam.
PS|55|19|Redimet in pace animam meam ab his, qui impugnant me,quoniam in multis sunt adversum me.
PS|55|20|Exaudiet Deus et humiliabit illos,qui est ante saecula.Non enim est illis commutatio,et non timuerunt Deum.
PS|55|21|Extendit manum suam in socios;contaminavit foedus suum.
PS|55|22|Lene super butyrum est os eius,pugna autem cor illius:molliti sunt sermones eius super oleum,et ipsi sunt gladii destricti. -
PS|55|23|Iacta super Dominum curam tuam,et ipse te enutriet;non dabit in aeternum fluctuationem iusto.
PS|55|24|Tu vero, Deus, deduces eos in puteum interitus.Viri sanguinum et dolosi non dimidiabunt dies suos;ego autem sperabo in te, Domine.
PS|56|1|Magistro chori. Secundum " Ionat elem rehoqim ".David. Miktam. Cum Gath Philistaei eum tenerent.
PS|56|2|Miserere mei, Deus, quoniam conculcavit me homo,tota die impugnans oppressit me.
PS|56|3|Conculcaverunt me inimici mei tota die,quoniam multi pugnant adversum me, Altissime.
PS|56|4|In quacumque die timebo,ego in te sperabo.
PS|56|5|In Deo, cuius laudabo sermonem,in Deo speravi;non timebo: quid faciet mihi caro?
PS|56|6|Tota die rem meam perturbabant,adversum me omnes cogitationes eorum in malum.
PS|56|7|Concitabant iurgia, insidiabantur,ipsi calcaneum meum observabant.Sicut quaesierunt animam meam,
PS|56|8|ita pro iniquitate retribue illis,in ira populos prosterne, Deus.
PS|56|9|Peregrinationes meas tu numerasti:pone lacrimas meas in utre tuo;nonne in supputatione tua?
PS|56|10|Tunc convertentur inimici mei retrorsum,in quacumque die invocavero:ecce cognovi quoniam Deus meus es.
PS|56|11|In Deo, cuius laudabo sermonem,in Domino, cuius laudabo sermonem,
PS|56|12|in Deo speravi;non timebo: quid faciet mihi homo?
PS|56|13|Super me sunt, Deus, vota tua;reddam laudationes tibi,
PS|56|14|quoniam eripuisti animam meam de morteet pedes meos de lapsu,ut ambulem coram Deo in lumine viventium.
PS|57|1|Magistro chori. Secundum " Ne destruxeris ". David.Miktam. Quando a Saul in cavernam fugit.
PS|57|2|Miserere mei, Deus, miserere mei,quoniam in te confugit anima mea;et in umbra alarum tuarum confugiam,donec transeant insidiae.
PS|57|3|Clamabo ad Deum Altissimum,Deum, qui benefecit mihi.
PS|57|4|Mittet de caelo et liberabit me;dabit in opprobrium conculcantes me.Mittet Deus misericordiam suam et veritatem suam.
PS|57|5|Anima mea recumbit in medio catulorum leonumdevorantium filios hominum.Dentes eorum arma et sagittae,et lingua eorum gladius acutus.
PS|57|6|Exaltare super caelos, Deus,super omnem terram gloria tua.
PS|57|7|Laqueum paraverunt pedibus meis,et incurvavit se anima mea;foderunt ante faciem meam foveam,et ipsi inciderunt in eam.
PS|57|8|Paratum cor meum, Deus,paratum cor meum;
PS|57|9|cantabo et psalmum dicam.Exsurge, gloria mea;exsurge, psalterium et cithara,excitabo auroram.
PS|57|10|Confitebor tibi in populis, Domine,et psalmum dicam tibi in nationibus,
PS|57|11|quoniam magnificata est usque ad caelos misericordia tua,et usque ad nubes veritas tua.
PS|57|12|Exaltare super caelos, Deus,super omnem terram gloria tua.
PS|58|1|Magistro chori. Secundum " Ne destruxeris ".David. Miktam.
PS|58|2|Numquid vere, potentes, iustitiam loquimini,recte iudicatis filios hominum?
PS|58|3|Etenim in corde iniquitates operamini,in terra violentiam manus vestrae concinnant.
PS|58|4|Alienati sunt peccatores ab utero;erraverunt a ventre, qui loquuntur falsa.
PS|58|5|Venenum illis in similitudinem serpentis,sicut aspidis surdae et obturantis aures suas,
PS|58|6|quae non exaudiet vocem incantantiumet venefici incantantis sapienter.
PS|58|7|Deus, contere dentes eorum in ore ipsorum;molas leonum confringe, Domine.
PS|58|8|Diffluant tamquam aqua decurrens,sicut fenum conculcatum arescant.
PS|58|9|Sicut limax, quae tabescens transit, sicut abortivum mulieris, quod non vidit solem.
PS|58|10|Priusquam sentiant ollae vestrae rhamnum,sicut viventes, sicut ardor irae absorbet eos.
PS|58|11|Laetabitur iustus, cum viderit vindictam,pedes suos lavabit in sanguine peccatoris.
PS|58|12|Et dicet homo: " Utique est fructus iusto,utique est Deus iudicans eos in terra ".
PS|59|1|Magistro chori. Secundum " Ne destruxeris ".David. Miktam. Quando Saul viros misit,qui domum observarent et eum occiderent.
PS|59|2|Eripe me de inimicis meis, Deus meus,et ab insurgentibus in me protege me.
PS|59|3|Eripe me de operantibus iniquitatemet de viris sanguinum salva me.
PS|59|4|Quia ecce insidiati sunt animae meae,irruerunt in me fortes.
PS|59|5|Neque delictum neque peccatum in me est, Domine;sine iniquitate mea currunt et praeparantur.Exsurge in occursum meum et vide;
PS|59|6|et tu, Domine, Deus virtutum, Deus Israel,evigila ad visitandas omnes gentes; non miserearis omnibus, qui infideliter operantur.
PS|59|7|Revertentur ad vesperam et latrabunt ut caneset circuibunt civitatem.
PS|59|8|Ecce eructabunt ore suo,et gladius in labiis eorum: " Quis enim audit? ".
PS|59|9|Et tu, Domine, deridebis eos,subsannabis omnes gentes.
PS|59|10|Fortitudo mea, tibi attendam,quia, Deus, praesidium meum es.
PS|59|11|Deus meus, misericordia eius praeveniet me.Deus faciet, ut despiciam inimicos meos.
PS|59|12|Ne occidas eos, ne quando obliviscatur populus meus;disperge illos in virtute tuaet prosterne eos, protector meus, Domine.
PS|59|13|Peccatum oris eorum, sermo labiorum ipsorum,et comprehendantur in superbia sua.Propter exsecrationem et mendacium, quod loquuntur,
PS|59|14|consume eos in furore,consume, et non erunt;et scient quia Deus dominabitur Iacob et finium terrae.
PS|59|15|Revertentur ad vesperam et latrabunt ut caneset circuibunt civitatem.
PS|59|16|Ipsi errabunt ad manducandum;si vero non fuerint saturati, murmurabunt.
PS|59|17|Ego autem cantabo fortitudinem tuamet exsultabo mane misericordiam tuam,quia factus es praesidium meumet refugium meum in die tribulationis meae.
PS|59|18|Fortitudo mea, tibi psallam,quia, Deus, praesidium meum es:Deus meus misericordia mea.
PS|60|1|Magistro chori. Secundum " Lilium praecepti ".Miktam. David. Ad docendum.
PS|60|2|Quando contra Aram Naharaim et Aram Soba egressus est,et quando Ioab reversus devicit Edom in valle Salis:duodecim milia (hominum).
PS|60|3|Deus, reppulisti nos, destruxisti nos.Iratus es. Convertere ad nos!
PS|60|4|Concussisti terram, confregisti eam;sana contritiones eius, quia commota est.
PS|60|5|Ostendisti populo tuo dura,potasti nos vino vertiginis.
PS|60|6|Dedisti metuentibus te signum,ut fugiant a facie arcus.
PS|60|7|Ut liberentur dilecti tui,salvos fac dextera tua et exaudi nos.
PS|60|8|Deus locutus est in sancto suo: Laetabor et partibor Sichimamet convallem Succoth metibor.
PS|60|9|Meus est Galaad, et meus est Manasses,et Ephraim fortitudo capitis mei.Iuda sceptrum meum,
PS|60|10|Moab olla lavacri mei.Super Idumaeam extendam calceamentum meum,super Philistaeam vociferabor ".
PS|60|11|Quis adducet me in civitatem munitam?Quis deducet me usque in Idumaeam?
PS|60|12|Nonne tu, Deus, qui reppulisti nos;et non egredieris, Deus, in virtutibus nostris?Da nobis auxilium de tribulatione, quia vana salus hominis.
PS|60|13|In Deo faciemus virtutem,et ipse conculcabit tribulantes nos.
PS|61|1|Magistro chori. Fidibus. David.
PS|61|2|Exaudi, Deus, deprecationem meam,intende orationi meae.
PS|61|3|A finibus terrae ad te clamavi,dum anxiaretur cor meum.In petram inaccessam mihi deduc me!
PS|61|4|Quia factus es spes mea,turris fortitudinis a facie inimici.
PS|61|5|Inhabitabo in tabernaculo tuo in saecula,protegar in velamento alarum tuarum,
PS|61|6|quoniam tu, Deus meus, exaudisti vota mea,dedisti hereditatem timentium nomen tuum.
PS|61|7|Dies super dies regis adicies,annos eius usque in diem generationis et generationis.
PS|61|8|Sedeat in aeternum in conspectu Dei;misericordia et veritas servent eum.
PS|61|9|Sic psalmum dicam nomini tuo in saeculum saeculi,ut reddam vota mea de die in diem.
PS|62|1|Magistro chori. Secundum Iduthun. PSALMUS. David.
PS|62|2|In Deo tantum quiesce, anima mea,ab ipso enim salutare meum.
PS|62|3|Verumtamen ipse refugium meum et salutare meum,praesidium meum; non movebor amplius.
PS|62|4|Quousque irruitis in hominem, contunditis universi vostamquam parietem inclinatum et maceriam depulsam?
PS|62|5|Verumtamen de excelso suo cogitaverunt depellere;delectabantur mendacio.Ore suo benedicebant et corde suo maledicebant.
PS|62|6|In Deo tantum quiesce, anima mea, quoniam ab ipso patientia mea.
PS|62|7|Verumtamen ipse Deus meus et salutare meum,praesidium meum; non movebor.
PS|62|8|In Deo salutare meum et gloria mea; Deus fortitudinis meae, et refugium meum in Deo est.
PS|62|9|Sperate in eo, omnis congregatio populi,effundite coram illo corda vestra;Deus refugium nobis.
PS|62|10|Verumtamen vanitas filii Adam,mendacium filii hominum.In stateram si conscendant,super fumum leves sunt omnes.
PS|62|11|Nolite sperare in violentiaet in rapina nolite decipi;divitiae si affluant, nolite cor apponere.
PS|62|12|Semel locutus est Deus,duo haec audivi:quia potestas Deo est,
PS|62|13|et tibi, Domine, misericordia;quia tu reddes unicuique iuxta opera sua.
PS|63|1|PSALMUS. David, cum in deserto Iudae commoraretur.
PS|63|2|Deus, Deus meus es tu, ad te de luce vigilo.Sitivit in te anima mea,te desideravit caro mea.In terra deserta et arida et inaquosa,
PS|63|3|sic in sancto apparui tibi,ut viderem virtutem tuam et gloriam tuam.
PS|63|4|Quoniam melior est misericordia tua super vitas,labia mea laudabunt te.
PS|63|5|Sic benedicam te in vita meaet in nomine tuo levabo manus meas.
PS|63|6|Sicut adipe et pinguedine repleatur anima mea,et labiis exsultationis laudabit os meum.
PS|63|7|Cum memor ero tui super stratum meum,in matutinis meditabor de te,
PS|63|8|quia fuisti adiutor meus,et in velamento alarum tuarum exsultabo.
PS|63|9|Adhaesit anima mea post te,me suscepit dextera tua.
PS|63|10|Ipsi vero in ruinam quaesierunt animam meam,introibunt in inferiora terrae,
PS|63|11|tradentur in potestatem gladii,partes vulpium erunt.
PS|63|12|Rex vero laetabitur in Deo;gloriabuntur omnes, qui iurant in eo,quia obstructum est os loquentium iniqua.
PS|64|1|Magistro chori. PSALMUS. David.
PS|64|2|Exaudi, Deus, vocem meam in meditatione mea;a timore inimici custodi animam meam.
PS|64|3|Protege me a conventu malignantium,a multitudine operantium iniquitatem.
PS|64|4|Qui exacuerunt ut gladium linguas suas,intenderunt sagittas suas, venefica verba,
PS|64|5|ut sagittent in occultis immaculatum.Subito sagittabunt eum et non timebunt,
PS|64|6|firmaverunt sibi consilium nequam.Disputaverunt, ut absconderent laqueos,dixerunt: " Quis videbit eos? ".
PS|64|7|Excogitaverunt iniqua, perfecerunt excogitata consilia.Interiora hominis et cor eius abyssus.
PS|64|8|Et sagittavit illos Deus;subito factae sunt plagae eorum,
PS|64|9|et infirmavit eos lingua eorum.Caput movebunt omnes, qui videbunt eos,
PS|64|10|et timebit omnis homo;et annuntiabunt opera Deiet facta eius intellegent.
PS|64|11|Laetabitur iustus in Domino et sperabit in eo,et gloriabuntur omnes recti corde.
PS|65|1|Magistro chori. PSALMUS. David. Canticum.
PS|65|2|Te decet hymnus, Deus, in Sion;et tibi reddetur votum in Ierusalem.
PS|65|3|Qui audis orationem,ad te omnis caro veniet propter iniquitatem.
PS|65|4|Etsi praevaluerunt super nos impietates nostrae,tu propitiaberis eis.
PS|65|5|Beatus, quem elegisti et assumpsisti; inhabitabit in atriis tuis.Replebimur bonis domus tuae,sanctitate templi tui.
PS|65|6|Mirabiliter in aequitateexaudies nos, Deus salutis nostrae,spes omnium finium terrae et maris longinqui.
PS|65|7|Firmans montes in virtute tua,accinctus potentia.
PS|65|8|Compescens sonitum maris,sonitum fluctuum eiuset tumultum populorum.
PS|65|9|Et timebunt, qui habitant terminos terrae, a signis tuis;exitus orientis et occidentis delectabis.
PS|65|10|Visitasti terram et inebriasti eam;multiplicasti locupletare eam.Flumen Dei repletum est aquis;parasti frumenta illorum,quoniam ita parasti eam.
PS|65|11|Sulcos eius irrigans, glebas eius complanans;imbribus emollis eam, benedicis germini eius.
PS|65|12|Coronasti annum benignitate tua,et vestigia tua stillabunt pinguedinem.
PS|65|13|Stillabunt pascua deserti,et exsultatione colles accingentur.
PS|65|14|Induta sunt ovibus prata,et valles abundabunt frumento;clamabunt, etenim hymnum dicent.
PS|66|1|Magistro chori. Canticum. PSALMUS.Iubilate Deo, omnis terra,
PS|66|2|psalmum dicite gloriae nominis eius,glorificate laudem eius.
PS|66|3|Dicite Deo: " Quam terribilia sunt opera tua.Prae multitudine virtutis tuae blandientur tibi inimici tui.
PS|66|4|Omnis terra adoret te et psallat tibi,psalmum dicat nomini tuo ".
PS|66|5|Venite et videte opera Dei,terribilis in adinventionibus super filios hominum.
PS|66|6|Convertit mare in aridam,et in flumine pertransibunt pede;ibi laetabimur in ipso.
PS|66|7|Qui dominatur in virtute sua in aeternum,oculi eius super gentes respiciunt;rebelles non exaltentur in semetipsis.
PS|66|8|Benedicite, gentes, Deum nostrumet auditam facite vocem laudis eius;
PS|66|9|qui posuit animam nostram ad vitamet non dedit in commotionem pedes nostros.
PS|66|10|Quoniam probasti nos, Deus;igne nos examinasti, sicut examinatur argentum.
PS|66|11|Induxisti nos in laqueum,posuisti tribulationes in dorso nostro.
PS|66|12|Imposuisti homines super capita nostra,transivimus per ignem et aquam,et eduxisti nos in refrigerium.
PS|66|13|Introibo in domum tuam in holocaustis;reddam tibi vota mea,
PS|66|14|quae protulerunt labia mea,et locutum est os meum in tribulatione mea.
PS|66|15|Holocausta medullata offeram tibi cum incenso arietum,offeram tibi boves cum hircis.
PS|66|16|Venite, audite, et narrabo, omnes, qui timetis Deum,quanta fecit animae meae.
PS|66|17|Ad ipsum ore meo clamaviet exaltavi in lingua mea.
PS|66|18|Iniquitatem si aspexi in corde meo,non exaudiet Dominus.
PS|66|19|Propterea exaudivit Deus,attendit voci deprecationis meae.
PS|66|20|Benedictus Deus, qui non amovit orationem meamet misericordiam suam a me.
PS|67|1|Magistro chori. Fidibus. PSALMUS. Canticum.
PS|67|2|Deus misereatur nostri et benedicat nobis;illuminet vultum suum super nos,
PS|67|3|ut cognoscatur in terra via tua,in omnibus gentibus salutare tuum.
PS|67|4|Confiteantur tibi populi, Deus;confiteantur tibi populi omnes.
PS|67|5|Laetentur et exsultent gentes,quoniam iudicas populos in aequitateet gentes in terra dirigis.
PS|67|6|Confiteantur tibi populi, Deus;confiteantur tibi populi omnes.
PS|67|7|Terra dedit fructum suum;benedicat nos Deus, Deus noster,
PS|67|8|benedicat nos Deus,et metuant eum omnes fines terrae.
PS|68|1|Magistro chori. David. PSALMUS. Canticum.
PS|68|2|Exsurgit Deus, et dissipantur inimici eius;et fugiunt, qui oderunt eum, a facie eius.
PS|68|3|Sicut dissipatur fumus, tu dissipas;sicut fluit cera a facie ignis,sic pereunt peccatores a facie Dei.
PS|68|4|Et iusti laetentur et exsultent in conspectu Deiet delectentur in laetitia.
PS|68|5|Cantate Deo, psalmum dicite nomini eius;iter facite ei, qui fertur super nubes:Dominus nomen illi.Iubilate in conspectu eius;
PS|68|6|pater orphanorum et iudex viduarum,Deus in habitaculo sancto suo.
PS|68|7|Deus, qui inhabitare facit desolatos in domo,qui educit vinctos in prosperitatem;verumtamen rebelles habitabunt in arida terra. -
PS|68|8|Deus, cum egredereris in conspectu populi tui,cum pertransires in deserto,
PS|68|9|terra mota est, etiam caeli distillaverunta facie Dei Sinai, a facie Dei Israel.
PS|68|10|Pluviam voluntariam effundebas, Deus;hereditatem tuam infirmatam, tu refecisti eam.
PS|68|11|Animalia tua habitabant in ea,parasti in bonitate tua pauperi, Deus.
PS|68|12|Dominus dat verbum;virgines annuntiantes bona sunt agmen ingens:
PS|68|13|" Reges exercituum fugiunt, fugiunt,et species domus dividit spolia.
PS|68|14|Et vos dormitis inter medias caulas:alae columbae nitent argento,et pennae eius pallore auri.
PS|68|15|Dum dispergit Omnipotens reges super eam,nive dealbatur Selmon ".
PS|68|16|Mons Dei mons Basan,mons cacuminum mons Basan.
PS|68|17|Ut quid invidetis, montes cacuminum,monti, in quo beneplacitum est Deo inhabitare?Etenim Dominus habitabit in finem.
PS|68|18|Currus Dei decem milia milium:Dominus venit de Sinai in sancta.
PS|68|19|Ascendisti in altum, captivam duxisti captivitatem;accepisti in donum homines,ut etiam rebelles habitent apud Dominum Deum.
PS|68|20|Benedictus Dominus die cotidie;portabit nos Deus salutarium nostrorum.
PS|68|21|Deus noster, Deus ad salvandum;et Domini, Domini exitus mortis.
PS|68|22|Verumtamen Deus confringet capita inimicorum suorum,verticem capillatum perambulantium in delictis suis.
PS|68|23|Dixit Dominus: " Ex Basan reducam,reducam de profundo maris,
PS|68|24|ut intingatur pes tuus in sanguine,lingua canum tuorum ex inimicis portionem inveniat ".
PS|68|25|Viderunt ingressus tuos, Deus,ingressus Dei mei, regis mei in sancta.
PS|68|26|Praecedunt cantores, postremi veniunt psallentes.in medio iuvenculae tympanistriae.
PS|68|27|" In ecclesiis benedicite Deo,Domino, vos de fontibus Israel ".
PS|68|28|Ibi Beniamin adulescentulus ducens eos,principes Iudae cum turma sua,principes Zabulon, principesNephthali.
PS|68|29|Manda, Deus, virtuti tuae;confirma hoc, Deus, quod operatus es in nobis.
PS|68|30|A templo tuo in Ierusalemtibi afferent reges munera.
PS|68|31|Increpa feram arundinis,congregationem taurorum in vitulis populorum:prosternant se cum laminis argenti.Dissipa gentes, quae bella volunt.
PS|68|32|Venient optimates ex Aegypto,Aethiopia praeveniet manus suas Deo.
PS|68|33|Regna terrae, cantate Deo,psallite Domino, psallite Deo,
PS|68|34|qui fertur super caelum caeli ad orientem;ecce dabit vocem suam, vocem virtutis.
PS|68|35|Tribuite virtutem Deo.Super Israel magnificentia eius,et virtus eius in nubibus.
PS|68|36|Mirabilis, Deus, de sanctuario tuo!Deus Israel ipse tribuet virtutem et fortitudinem plebi suae.Benedictus Deus!
PS|69|1|Magistro chori. Secundum " Lilia... ". David.
PS|69|2|Salvum me fac, Deus,quoniam venerunt aquae usque ad guttur meum.
PS|69|3|Infixus sum in limo profundi, et non est substantia;veni in profunda aquarum, et fluctus demersit me.
PS|69|4|Laboravi clamans, raucae factae sunt fauces meae;defecerunt oculi mei, dum spero in Deum meum.
PS|69|5|Multiplicati sunt super capillos capitis mei,qui oderunt me gratis.Confortati sunt, qui persecuti sunt me inimici mei mendaces;quae non rapui, tunc exsolvebam.
PS|69|6|Deus, tu scis insipientiam meam,et delicta mea a te non sunt abscondita.
PS|69|7|Non erubescant in me, qui exspectant te,Domine, Domine virtutum.Non confundantur super me,qui quaerunt te, Deus Israel.
PS|69|8|Quoniam propter te sustinui opprobrium,operuit confusio faciem meam;
PS|69|9|extraneus factus sum fratribus meiset peregrinus filiis matris meae.
PS|69|10|Quoniam zelus domus tuae comedit me,et opprobria exprobrantium tibi ceciderunt super me.
PS|69|11|Et flevi in ieiunio animam meam,et factum est in opprobrium mihi.
PS|69|12|Et posui vestimentum meum cilicium,et factus sum illis in parabolam.
PS|69|13|Adversum me loquebantur, qui sedebant in porta,et in me canebant, qui bibebant vinum.
PS|69|14|Ego vero orationem meam ad te, Domine,in tempore beneplaciti, Deus.In multitudine misericordiae tuae exaudi me,in veritate salutis tuae.
PS|69|15|Eripe me de luto, ut non infigar,eripiar ab iis, qui oderunt me,et de profundis aquarum.
PS|69|16|Non me demergat fluctus aquarum,neque absorbeat me profundum,neque urgeat super me puteus os suum.
PS|69|17|Exaudi me, Domine, quoniam benigna est misericordia tua;secundum multitudinem miserationum tuarum respice in me.
PS|69|18|Et ne avertas faciem tuam a puero tuo;quoniam tribulor, velociter exaudi me.
PS|69|19|Accede ad animam meam, vindica eam,propter inimicos meos redime me.
PS|69|20|Tu scis opprobrium meumet confusionem meam et reverentiam meam. -In conspectu tuo sunt omnes, qui tribulant me;
PS|69|21|opprobrium contrivit cor meum, et elangui.Et sustinui, qui simul contristaretur, et non fuit,et qui consolaretur, et non inveni.
PS|69|22|Et dederunt in escam meam felet in siti mea potaverunt me aceto.
PS|69|23|Fiat mensa eorum coram ipsis in laqueumet in retributiones et in scandalum.
PS|69|24|Obscurentur oculi eorum, ne videant,et lumbos eorum semper infirma.
PS|69|25|Effunde super eos iram tuam,et furor irae tuae comprehendat eos.
PS|69|26|Fiat commoratio eorum deserta,et in tabernaculis eorum non sit qui inhabitet.
PS|69|27|Quoniam, quem tu percussisti, persecuti sunt,et super dolorem eius, quem vulnerasti, addiderunt.
PS|69|28|Appone iniquitatem super iniquitatem eorum,et non veniant ad iustitiam tuam.
PS|69|29|Deleantur de libro viventiumet cum iustis non scribantur.
PS|69|30|Ego autem sum pauper et dolens;salus tua, Deus, suscipit me.
PS|69|31|Laudabo nomen Dei cum canticoet magnificabo eum in laude.
PS|69|32|Et placebit Domino super taurum,super vitulum cornua producentem et ungulas.
PS|69|33|Videant humiles et laetentur;quaerite Deum, et vivet cor vestrum,
PS|69|34|quoniam exaudivit pauperes Dominuset vinctos suos non despexit.
PS|69|35|Laudent illum caeli et terra,maria et omnia reptilia in eis.
PS|69|36|Quoniam Deus salvam faciet Sionet aedificabit civitates Iudae;et inhabitabunt ibi et possidebunt eam.
PS|69|37|Et semen servorum eius hereditabunt eam;et, qui diligunt nomen eius, habitabunt in ea.
PS|70|1|Magistro chori. David. Ad commemorandum.
PS|70|2|Deus, in adiutorium meum intende;Domine, ad adiuvandum me festina.
PS|70|3|Confundantur et revereantur,qui quaerunt animam meam.Avertantur retrorsum et erubescant,qui volunt mihi mala.
PS|70|4|Convertantur propter confusionem suam,qui dicunt mihi: " Euge, euge ".
PS|70|5|Exsultent et laetentur in te omnes, qui quaerunt te;et dicant semper: " Magnificetur Deus ",qui diligunt salutare tuum.
PS|70|6|Ego vero egenus et pauper sum;Deus, ad me festina.Adiutor meus et liberator meus es tu;Domine, ne moreris.
PS|71|1|In te, Domine, speravi,non confundar in aeternum.
PS|71|2|In iustitia tua libera me et eripe me;inclina ad me aurem tuam et salva me.
PS|71|3|Esto mihi in rupem praesidiiet in domum munitam, ut salvum me facias,quoniam fortitudo mea et refugium meum es tu.
PS|71|4|Deus meus, eripe me de manu peccatoriset de manu contra legem agentis et iniqui.
PS|71|5|Quoniam tu es exspectatio mea, Domine;Domine, spes mea a iuventute mea.
PS|71|6|Super te innixus sum ex utero,de ventre matris meae tu es susceptor meus;in te laus mea semper.
PS|71|7|Tamquam prodigium factus sum multis,et tu adiutor fortis. -
PS|71|8|Repleatur os meum laude tua,tota die magnitudine tua.
PS|71|9|Ne proicias me in tempore senectutis;cum defecerit virtus mea, ne derelinquas me.
PS|71|10|Quia dixerunt inimici mei mihi,et, qui observabant animam meam,consilium fecerunt in unum
PS|71|11|dicentes: " Deus dereliquit eum!Persequimini et comprehenditeeum,quia non est qui eripiat ".
PS|71|12|Deus, ne elongeris a me;Deus meus, in auxilium meum festina.
PS|71|13|Confundantur et deficiant adversantes animae meae;operiantur confusione et pudore, qui quaerunt mala mihi.
PS|71|14|Ego autem semper speraboet adiciam super omnem laudem tuam.
PS|71|15|Os meum annuntiabit iustitiam tuam,tota die salutare tuum:quae dinumerare nescivi.
PS|71|16|Veniam ad potentias Domini;Domine, memorabor iustitiae tuae solius.
PS|71|17|Deus, docuisti me a iuventute mea;et usque nunc annuntiabo mirabilia tua.
PS|71|18|Et usque in senectam et senium,Deus, ne derelinquas me,donec annuntiem brachium tuumgenerationi omni, quae ventura est.Potentia tua
PS|71|19|et iustitia tua, Deus,usque in altissima, qui fecisti magnalia:Deus, quis similis tibi?
PS|71|20|Quantas ostendisti mihi tribulationes multas et malas;iterum vivificasti meet de abyssis terrae iterum reduxisti me.
PS|71|21|Multiplicabis magnitudinem meam et conversus consolaberis me.
PS|71|22|Nam et ego confitebor tibiin psalterio veritatem tuam, Deus meus;psallam tibi in cithara, Sanctus Israel.
PS|71|23|Exsultabunt labia mea, cum cantavero tibi,et anima mea, quam redemisti;
PS|71|24|sed et lingua mea tota die meditabitur iustitiam tuam,cum confusi et reveriti fuerint, qui quaerunt mala mihi.
PS|72|1|Salomonis. Deus, iudicium tuum regi daet iustitiam tuam filio regis;
PS|72|2|iudicet populum tuum in iustitiaet pauperes tuos in iudicio.
PS|72|3|Afferant montes pacem populo,et colles iustitiam.
PS|72|4|Iudicabit pauperes populiet salvos faciet filios inopiset humiliabit calumniatorem.
PS|72|5|Et permanebit cum sole et ante lunamin generatione et generationem.
PS|72|6|Descendet sicut pluvia in gramen,et sicut imber irrigans terram.
PS|72|7|Florebit in diebus eius iustitia et abundantia pacis,donec auferatur luna.
PS|72|8|Et dominabitur a mari usque ad mareet a flumine usque ad terminos orbis terrarum.
PS|72|9|Coram illo procident incolae deserti,et inimici eius terram lingent.
PS|72|10|Reges Tharsis et insulae munera offerent,reges Arabum et Saba dona adducent.
PS|72|11|Et adorabunt eum omnes reges, omnes gentes servient ei.
PS|72|12|Quia liberabit inopem clamantemet pauperem, cui non erat adiutor.
PS|72|13|Parcet pauperi et inopiet animas pauperum salvas faciet.
PS|72|14|Ex oppressione et violentia redimet animas eorum,et pretiosus erit sanguis eorum coram illo. -
PS|72|15|Et vivet, et dabitur ei de auro Arabiae, et orabunt pro ipso semper; tota die benedicent ei.
PS|72|16|Et erit ubertas frumenti in terra, in summis montium fluctuabit, sicut Libanus fructus eius;et florebunt de civitate sicut fenum terrae.
PS|72|17|Sit nomen eius benedictum in saecula,ante solem permanebit nomen eius.Et benedicentur in ipso omnes tribus terrae,omnes gentes magnificabunt eum.
PS|72|18|Benedictus Dominus Deus, Deus Israel,qui facit mirabilia solus.
PS|72|19|Et benedictum nomen maiestatis eius in aeternum;et replebitur maiestate eius omnis terra. Fiat, fiat.
PS|73|1|PSALMUS. Asaph.Quam bonus rectis est Deus,Deus his, qui mundo sunt corde!
PS|73|2|Mei autem paene moti sunt pedes,paene effusi sunt gressus mei,
PS|73|3|quia zelavi super gloriantes,pacem peccatorum videns.
PS|73|4|Quia non sunt eis impedimenta,sanus et pinguis est venter eorum.
PS|73|5|In labore mortalium non suntet cum hominibus non flagellantur.
PS|73|6|Ideo quasi torques est eis superbia,et tamquam indumentum operuit eos violentia.
PS|73|7|Prodit quasi ex adipe iniquitas eorum,erumpunt cogitationes cordis.
PS|73|8|Subsannaverunt et locuti sunt nequitiam,iniquitatem ab excelso locuti sunt.
PS|73|9|Posuerunt in caelo os suum,et lingua eorum transivit in terra.
PS|73|10|Ideo in alto sedent,et aquae plenae non pervenient ad eos.
PS|73|11|Et dixerunt: " Quomodo scit Deus,et si est scientia in Excelso? ".
PS|73|12|Ecce ipsi peccatores et abundantes in saeculomultiplicaverunt divitias.
PS|73|13|Et dixi: " Ergo sine causa mundavi cor meumet lavi in innocentia manus meas;
PS|73|14|et fui flagellatus tota die,et castigatio mea in matutinis ".
PS|73|15|Si dixissem: " Loquar ut illi ",ecce generationem filiorum tuorum prodidissem.
PS|73|16|Et cogitabam, ut cognoscerem hoc;labor erat in oculis meis,
PS|73|17|donec intravi in sanctuarium Deiet intellexi novissima eorum.
PS|73|18|Verumtamen in lubrico posuisti eos,deiecisti eos in ruinas.
PS|73|19|Quomodo facti sunt in desolationem!Subito defecerunt, perierunt prae horrore.
PS|73|20|Velut somnium evigilantis, Domine,surgens imaginem ipsorum contemnes.
PS|73|21|Quia exacerbatum est cor meum,et renes mei compuncti sunt;
PS|73|22|et ego insipiens factus sum et nescivi:ut iumentum factus sum apud te.
PS|73|23|Ego autem semper tecum;tenuisti manum dexteram meam.
PS|73|24|In consilio tuo deduces meet postea cum gloria suscipies me.
PS|73|25|Quis enim mihi est in caelo?Et tecum nihil volui super terram.
PS|73|26|Defecit caro mea et cor meum;Deus cordis mei, et pars mea Deus in aeternum.
PS|73|27|Quia ecce, qui elongant se a te, peribunt;perdidisti omnes, qui fornicantur abs te.
PS|73|28|Mihi autem adhaerere Deo bonum est,ponere in Domino Deo spem meam,ut annuntiem omnes operationes tuasin portis filiae Sion.
PS|74|1|Maskil. Asaph.Ut quid, Deus, reppulisti in finem,iratus est furor tuus super oves pascuae tuae?
PS|74|2|Memor esto congregationis tuae,quam possedisti ab initio.Redemisti virgam hereditatis tuae: mons Sion, in quo habitasti.
PS|74|3|Leva gressus tuos in ruinas sempiternas:omnia vastavit inimicus in sancto.
PS|74|4|Rugierunt, qui oderunt te,in medio congregationis tuae;posuerunt signa sua in signa.
PS|74|5|Visi sunt quasi in altum securim vibrantesin silva condensa.
PS|74|6|Exciderunt ianuas eius in idipsum;in securi et ascia deiecerunt.
PS|74|7|Incenderunt igni sanctuarium tuum,in terram polluerunt tabernaculum nominis tui;
PS|74|8|dixerunt in corde suo: " Opprimamus eos simul ".Combusserunt omnes congregationes Dei in terra.
PS|74|9|Signa nostra non vidimus;iam non est propheta,et apud nos non est qui cognoscat amplius.
PS|74|10|Usquequo, Deus, improperabit inimicus,spernet adversarius nomen tuum in finem?
PS|74|11|Ut quid avertis manum tuamet tenes dexteram tuam in medio sinu tuo?
PS|74|12|Deus autem rex noster ante saecula,operatus est salutes in medio terrae.
PS|74|13|Tu conscidisti in virtute tua mare,contribulasti capita draconum in aquis.
PS|74|14|Tu confregisti capita Leviathan,dedisti eum escam monstris maris.
PS|74|15|Tu dirupisti fontes et torrentes;tu siccasti fluvios perennes.
PS|74|16|Tuus est dies, et tua est nox,tu fabricatus es luminaria et solem.
PS|74|17|Tu statuisti omnes terminos terrae,aestatem et hiemem, tu plasmasti ea.
PS|74|18|Memor esto huius:inimicus improperavit Domino,et populus insipiens sprevit nomen tuum.
PS|74|19|Ne tradas bestiis animas confitentes tibiet animas pauperum tuorum ne obliviscaris in finem.
PS|74|20|Respice in testamentum,quia repleta sunt latibula terrae tentoriis violentiae.
PS|74|21|Ne revertatur humilis factus confusus;pauper et inops laudabunt nomen tuum.
PS|74|22|Exsurge, Deus, iudica causam tuam;memor esto improperiorum tuorum,quae ab insipiente fiunt tota die.
PS|74|23|Ne obliviscaris voces inimicorum tuorum;tumultus adversariorum tuorum ascendit semper.
PS|75|1|Magistro chori. Secundum " Ne destruxeris ".PSALMUS. Asaph. Canticum.
PS|75|2|Confitebimur tibi, Deus;confitebimur et invocabimus nomen tuum:narrabimus mirabilia tua.
PS|75|3|Cum statuero tempus,ego iustitias iudicabo.
PS|75|4|Si liquefacta est terra et omnes, qui habitant in ea,ego confirmavi columnas eius.
PS|75|5|Dixi gloriantibus: " Nolite gloriari! "et delinquentibus: "Nolite exaltare cornu!
PS|75|6|Nolite exaltare in altum cornu vestrum;nolite loqui adversus Deum proterva ".
PS|75|7|Quia neque ab oriente neque ab occidenteneque a desertis exaltatio.
PS|75|8|Quoniam Deus iudex est:hunc humiliat et hunc exaltat.
PS|75|9|Quia calix in manu Dominivini meri plenus mixto.Et inclinavit ex hoc in hoc;verumtamen usque ad faeces epotabunt,bibent omnes peccatores terrae.
PS|75|10|Ego autem annuntiabo in saeculum,cantabo Deo Iacob.
PS|75|11|Et omnia cornua peccatorum confringam,et exaltabuntur cornua iusti.
PS|76|1|Magistro chori. Fidibus. PSALMUS. Asaph. Canticum.
PS|76|2|Notus in Iudaea Deus,in Israel magnum nomen eius.
PS|76|3|Et est in Salem tabernaculum eius,et habitatio eius in Sion.
PS|76|4|Ibi confregit coruscationes arcus,scutum, gladium et bellum.
PS|76|5|Illuminans tu, Mirabilis,a montibus direptionis.
PS|76|6|Spoliati sunt potentes corde, dormierunt somnum suum,et non invenerunt omnes viri fortes manus suas.
PS|76|7|Ab increpatione tua, Deus Iacob,dormitaverunt auriga et equus.
PS|76|8|Tu terribilis es, et quis resistet tibi?Ex tunc ira tua.
PS|76|9|De caelo auditum fecisti iudicium;terra tremuit et quievit,
PS|76|10|cum exsurgeret in iudicium Deus,ut salvos faceret omnes mansuetos terrae.
PS|76|11|Quoniam furor hominis confitebitur tibi,et reliquiae furoris diem festum agent tibi.
PS|76|12|Vovete et reddite Domino Deo vestro;omnes in circuitu eius afferant munera Terribili,
PS|76|13|ei, qui aufert spiritum principum,terribili apud reges terrae.
PS|77|1|Magistro chori. Secundum Idithun. Asaph. PSALMUS.
PS|77|2|Voce mea ad Dominum clamavi;voce mea ad Deum, et intendit mihi.
PS|77|3|In die tribulationis meae Deum exquisivi,manus meae nocte expansae suntet non fatigantur.Renuit consolari anima mea;
PS|77|4|memor sum Dei et ingemisco,exerceor, et deficit spiritus meus.
PS|77|5|Vigiles tenuisti palpebras oculi mei; turbatus sum et non sum locutus.
PS|77|6|Cogitavi dies antiquoset annos aeternos in mente habui.
PS|77|7|Meditatus sum nocte cum corde meoet exercitabar et scobebam spiritum meum.
PS|77|8|Numquid in aeternum proiciet Deus,aut non apponet, ut complacitior sit adhuc?
PS|77|9|Aut deficiet in finem misericordia sua,cessabit verbum a generatione in generationem?
PS|77|10|Aut obliviscetur misereri Deus,aut continebit in ira sua misericordias suas?
PS|77|11|Et dixi: " Hoc vulnus meum:mutatio dexterae Excelsi ".
PS|77|12|Memor ero operum Domini,memor ero ab initio mirabilium tuorum.
PS|77|13|Et meditabor in omnibus operibus tuiset in adinventionibus tuis exercebor.
PS|77|14|Deus, in sancto via tua;quis deus magnus sicut Deus noster?
PS|77|15|Tu es Deus, qui facis mirabilia,notam fecisti in populis virtutem tuam.
PS|77|16|Redemisti in brachio tuo populum tuum,filios Iacob et Ioseph.
PS|77|17|Viderunt te aquae, Deus,viderunt te aquae et doluerunt;etenim commotae sunt abyssi.
PS|77|18|Effuderunt aquas nubila,vocem dederunt nubes,etenim sagittae tuae transeunt.
PS|77|19|Vox tonitrui tui in rota;illuxerunt coruscationes tuae orbi terrae,commota est et contremuit terra.
PS|77|20|In mari via tua, et semitae tuae in aquis multis;et vestigia tua non cognoscuntur.
PS|77|21|Deduxisti sicut oves populum tuumin manu Moysi et Aaron.
PS|78|1|Maskil. Asaph.Attendite, popule meus, doctrinam meam;inclinate aurem vestram in verba oris mei.
PS|78|2|Aperiam in parabolis os meum,eloquar arcana aetatis antiquae.
PS|78|3|Quanta audivimus et cognovimus ea,et patres nostri narraverunt nobis,
PS|78|4|non occultabimus a filiis eorum,generationi alteri narranteslaudes Domini et virtutes eiuset mirabilia eius, quae fecit.
PS|78|5|Constituit testimonium in Iacobet legem posuit in Israel;quanta mandaverat patribus nostrisnota facere ea filiis suis,
PS|78|6|ut cognoscat generatio altera,filii, qui nascentur.Exsurgent et narrabunt filiis suis,
PS|78|7|ut ponant in Deo spem suamet non obliviscantur operum Deiet mandata eius custodiant.
PS|78|8|Ne fiant sicut patres eorum,generatio rebellis et exasperans;generatio, quae non firmavit cor suum,et non fuit fidelis Deo spiritus eius.
PS|78|9|Filii Ephraim, intendentes et mittentes arcum,conversi sunt in die belli.
PS|78|10|Non custodierunt testamentum Deiet in lege eius renuerunt ambulare.
PS|78|11|Et obliti sunt factorum eiuset mirabilium eius, quae ostendit eis.
PS|78|12|Coram patribus eorum fecit mirabiliain terra Aegypti, in campo Taneos.
PS|78|13|Scidit mare et perduxit eoset statuit aquas quasi in utre.
PS|78|14|Et deduxit eos in nube per diemet per totam noctem in illuminatione ignis.
PS|78|15|Scidit petram in eremoet adaquavit eos velut abyssus multa.
PS|78|16|Et eduxit rivulos de petraet deduxit tamquam flumina aquas.
PS|78|17|Et apposuerunt adhuc peccare ei,in iram excitaverunt Excelsum in inaquoso.
PS|78|18|Et tentaverunt Deum in cordibus suis,petentes escas animabus suis;
PS|78|19|et contra Deum locuti sunt,dixerunt: " Numquid poterit Deus parare mensam in deserto? ".
PS|78|20|Ecce percussit petram, et fluxerunt aquae,et torrentes inundaverunt. Numquid et panem poterit dareaut parare carnes populo suo? ".
PS|78|21|Ideo audivit Dominus et exarsit,et ignis accensus est in Iacob,et ira ascendit in Israel.
PS|78|22|Quia non crediderunt in Deonec speraverunt in salutari eius.
PS|78|23|Verumtamen mandavit nubibus desuperet ianuas caeli aperuit;
PS|78|24|et pluit illis manna ad manducandumet panem caeli dedit eis:
PS|78|25|panem angelorum manducavit homo;cibaria misit eis ad abundantiam.
PS|78|26|Excitavit austrum in caeloet induxit in virtute sua africum;
PS|78|27|et pluit super eos sicut pulverem carneset sicut arenam maris volatilia pennata:
PS|78|28|et ceciderunt in medio castrorum eorum,circa tabernacula eorum.
PS|78|29|Et manducaverunt et saturati sunt nimis,et desiderium eorum attulit eis.
PS|78|30|Nondum recesserant a desiderio suo,adhuc escae eorum erant in ore ipsorum,
PS|78|31|et ira Dei ascendit super eoset occidit pingues eorumet electos Israel prostravit.
PS|78|32|In omnibus his peccaverunt adhucet non crediderunt in mirabilibus eius;
PS|78|33|et consumpsit in halitu dies eorumet annos eorum cum festinatione.
PS|78|34|Cum occideret eos, quaerebant eumet conversi veniebant diluculo ad eum;
PS|78|35|et rememorati sunt quia Deus adiutor est eorum,et Deus Excelsus redemptor eorum est.
PS|78|36|Et suaserunt ei in ore suoet lingua sua mentiti sunt ei;
PS|78|37|cor autem eorum non erat rectum cum eo,nec fideles erant in testamento eius.
PS|78|38|Ipse autem est misericorset propitiatur iniquitati et non disperdit.Saepe avertit iram suamet non accendit omnem furorem suum.
PS|78|39|Et recordatus est quia caro sunt,spiritus vadens et non rediens.
PS|78|40|Quoties exacerbaverunt eum in deserto,in iram concitaverunt eum in inaquoso!
PS|78|41|Et reversi sunt et tentaverunt Deumet Sanctum Israel exacerbaverunt.
PS|78|42|Non sunt recordati manus eius,diei, qua redemit eos de manu tribulantis.
PS|78|43|Cum posuit in Aegypto signa suaet prodigia sua in campo Taneos.
PS|78|44|Convertit in sanguinem flumina eorumet rivulos eorum, ne biberent.
PS|78|45|Misit in eos coenomyiam et comedit eos,ranam et perdidit eos.
PS|78|46|Dedit brucho fructus eorum,labores eorum locustae.
PS|78|47|Occidit in grandine vineas eorum,moros eorum in pruina.
PS|78|48|Tradidit grandini iumenta eorumet greges eorum flammae ignis.
PS|78|49|Misit in eos ardorem irae suae,indignationem et comminationem et angustiam,immissionem angelorum malorum.
PS|78|50|Complanavit semitam irae suae;non pepercit a morte animabus eorumet vitam eorum in peste conclusit.
PS|78|51|Percussit omne primogenitum in terra Aegypti,primitias roboris eorum in tabernaculis Cham.
PS|78|52|Abstulit sicut oves populum suumet perduxit eos tamquam gregem in deserto.
PS|78|53|Deduxit eos in spe, et non timuerunt,et inimicos eorum operuit mare.
PS|78|54|Et induxit eos in fines sanctificationis suae,in montem, quem acquisivit dextera eius.
PS|78|55|Et eiecit a facie eorum genteset divisit eis terram in funiculo hereditatiset habitare fecit in tabernaculis eorum tribus Israel.
PS|78|56|Et tentaverunt et exacerbaverunt Deum Excelsumet testimonia eius non custodierunt.
PS|78|57|Recesserunt et praevaricati sunt,quemadmodum patres eorum;conversi sunt retro ut arcus pravus.
PS|78|58|In iram concitaverunt eum in collibus suiset in sculptilibus suis ad aemulationem eum provocaverunt.
PS|78|59|Audivit Deus et exarsitet sprevit valde Israel.
PS|78|60|Et reppulit habitaculum Silo,tabernaculum, ubi habitavit in hominibus.
PS|78|61|Et tradidit in captivitatem virtutem suamet pulchritudinem suam in manus inimici.
PS|78|62|Et conclusit in gladio populum suumet in hereditatem suam exarsit.
PS|78|63|Iuvenes eorum comedit ignis,et virgines eorum non sunt desponsatae.
PS|78|64|Sacerdotes eorum in gladio ceciderunt,et viduae eorum non plorabantur.
PS|78|65|Et excitatus est tamquam dormiens Dominus,tamquam potens crapulatus a vino.
PS|78|66|Et percussit inimicos suos in posteriora,opprobrium sempiternum dedit illis.
PS|78|67|Et reppulit tabernaculum Iosephet tribum Ephraim non elegit,
PS|78|68|sed elegit tribum Iudae,montem Sion, quem dilexit.
PS|78|69|Et aedificavit sicut excelsum sanctuarium suum,sicut terram, quam fundavit in saecula.
PS|78|70|Et elegit David servum suumet sustulit eum de gregibus ovium,
PS|78|71|de post fetantes accepit eum:pascere Iacob populum suumet Israel hereditatem suam.
PS|78|72|Et pavit eos in innocentia cordis suiet in prudentia manuum suarum deduxit eos.
PS|79|1|PSALMUS. Asaph.Deus, venerunt gentes in hereditatem tuam,polluerunt templum sanctum tuum,posuerunt Ierusalem in ruinas.
PS|79|2|Dederunt morticina servorum tuorum escas volatilibus caeli,carnes sanctorum tuorum bestiis terrae.
PS|79|3|Effuderunt sanguinem eorum tamquam aquamin circuitu Ierusalem, et non erat qui sepeliret.
PS|79|4|Facti sumus opprobrium vicinis nostris,subsannatio et illusio his, qui in circuitu nostro sunt.
PS|79|5|Usquequo, Domine? Irasceris in finem?Accendetur velut ignis zelus tuus?
PS|79|6|Effunde iram tuam in gentes, quae te non noverunt,et in regna, quae nomen tuum non invocaverunt,
PS|79|7|quia comederunt Iacobet sedem eius desolaverunt.
PS|79|8|Ne memineris iniquitatum patrum nostrorum,cito anticipent nos misericordiae tuae,quia pauperes facti sumus nimis.
PS|79|9|Adiuva nos, Deus salutaris nostri,propter gloriam nominis tui et libera nos;et propitius esto peccatis nostris propter nomen tuum.
PS|79|10|Quare dicent in gentibus: " Ubi est Deus eorum? ".Innotescat in nationibus coram oculis nostrisultio sanguinis servorum tuorum, qui effusus est.
PS|79|11|Introeat in conspectu tuo gemitus compeditorum;secundum magnitudinem brachii tuisuperstites relinque filios mortis.
PS|79|12|Et redde vicinis nostris septuplum in sinu eorum,improperium ipsorum, quod exprobraverunt tibi, Domine.
PS|79|13|Nos autem, populus tuus et oves pascuae tuae,confitebimur tibi in saeculum;in generationem et generationem annuntiabimus laudem tuam.
PS|80|1|Magistro chori. Secundum " Lilium praecepti ".Asaph. PSALMUS.
PS|80|2|Qui pascis Israel, intende,qui deducis velut ovem Ioseph.Qui sedes super cherubim, effulge
PS|80|3|coram Ephraim, Beniamin et Manasse.Excita potentiam tuam et veni,ut salvos facias nos.
PS|80|4|Deus, converte nos,illustra faciem tuam, et salvi erimus.
PS|80|5|Domine, Deus virtutum,quousque irasceris super orationem populi tui?
PS|80|6|Cibasti nos pane lacrimarumet potum dedisti nobis in lacrimis copiose.
PS|80|7|Posuisti nos in contradictionem vicinis nostris,et inimici nostri subsannaverunt nos.
PS|80|8|Deus virtutum, converte nos,illustra faciem tuam, et salvi erimus.
PS|80|9|Vineam de Aegypto transtulisti,eiecisti gentes et plantasti eam.
PS|80|10|Purgasti locum in conspectu eius,plantasti radices eius, et implevit terram.
PS|80|11|Operti sunt montes umbra eius,et ramis eius cedri Dei;
PS|80|12|extendit palmites suos usque ad mareet usque ad flumen propagines suas.
PS|80|13|Ut quid destruxisti maceriam eius,et vindemiant eam omnes, qui praetergrediuntur viam?
PS|80|14|Exterminavit eam aper de silva,et singularis ferus depastus est eam.
PS|80|15|Deus virtutum, convertere,respice de caelo et vide et visita vineam istam.
PS|80|16|Et protege eam, quam plantavit dextera tua,et super filium hominis, quem confirmasti tibi.
PS|80|17|Incensa est igni et suffossa;ab increpatione vultus tui peribunt.
PS|80|18|Fiat manus tua super virum dexterae tuae,super filium hominis, quem confirmasti tibi.
PS|80|19|Et non discedemus a te, vivificabis nos,et nomen tuum invocabimus.
PS|80|20|Domine, Deus virtutum, converte noset illustra faciem tuam, et salvi erimus.
PS|81|1|Magistro chori. Secundum " Torcularia... ". Asaph.
PS|81|2|Exsultate Deo adiutori nostro;iubilate Deo Iacob.
PS|81|3|Sumite psalmum et date tympanum,psalterium iucundum cum cithara.
PS|81|4|Bucinate in neomenia tuba,in die plenae lunae, in sollemnitate nostra.
PS|81|5|Quia praeceptum in Israel est,et iudicium Deo Iacob.
PS|81|6|Testimonium in Ioseph posuit illud,cum exiret de terra Aegypti;sermonem, quem non noveram, audivi:
PS|81|7|" Diverti ab oneribus dorsum eius;manus eius a cophino recesserunt.
PS|81|8|In tribulatione invocasti me, et liberavi te,exaudivi te in abscondito tempestatis,probavi te apud aquam Meriba.
PS|81|9|Audi, populus meus, et contestabor te;Israel, utinam audias me!
PS|81|10|Non erit in te deus alienus,neque adorabis deum extraneum.
PS|81|11|Ego enim sum Dominus Deus tuus,qui eduxi te de terra Aegypti;dilata os tuum, et implebo illud.
PS|81|12|Et non audivit populus meus vocem meam,et Israel non intendit mihi.
PS|81|13|Et dimisi eos secundum duritiam cordis eorum,ibunt in adinventionibus suis.
PS|81|14|Si populus meus audisset me,Israel si in viis meis ambulasset!
PS|81|15|In brevi inimicos eorum humiliassemet super tribulantes eos misissem manum meam.
PS|81|16|Inimici Domini blandirentur ei,et esset sors eorum in saecula;
PS|81|17|et cibarem eos ex adipe frumentiet de petra melle saturarem eos ".
PS|82|1|PSALMUS. Asaph.Deus stetit in concilio divino,in medio deorum iudicat.
PS|82|2|" Usquequo iudicabitis iniqueet facies peccatorum sumetis?
PS|82|3|Iudicate egeno et pupillo,humilem et pauperem iustificate.
PS|82|4|Eripite pauperemet egenum de manu peccatoris liberate ".
PS|82|5|Nescierunt neque intellexerunt, in tenebris ambulant;movebuntur omnia fundamenta terrae.
PS|82|6|Ego dixi: " Dii estis,et filii Excelsi omnes ".
PS|82|7|Vos autem sicut homines morieminiet sicut unus de principibus cadetis.
PS|82|8|Surge, Deus, iudica terram,quoniam tu hereditabis in omnibus gentibus.
PS|83|1|Canticum. PSALMUS. Asaph.
PS|83|2|Deus, ne quiescas, ne taceasneque compescaris, Deus,
PS|83|3|quoniam ecce inimici tui fremuerunt,et, qui oderunt te, extulerunt caput.
PS|83|4|Adversus populum tuum malignaverunt consiliumet cogitaverunt adversus eos, quos abscondisti tibi.
PS|83|5|Dixerunt: " Venite, et disperdamus eos de gente,et non memoretur nomen Israel ultra! ".
PS|83|6|Quoniam cogitaverunt unanimiter,adversum te testamentum statuerunt:
PS|83|7|tabernacula Idumaeorum et Ismaelitae,Moab et Agareni,
PS|83|8|Gebal et Ammon et Amalec,Philistaea cum habitantibus Tyrum.
PS|83|9|Etenim Assur sociabatur cum illis;facti sunt in adiutorium filiis Lot.
PS|83|10|Fac illis sicut Madian et Sisarae,sicut Iabin in torrente Cison.
PS|83|11|Disperierunt in Endor,facti sunt ut stercus super terram.
PS|83|12|Pone duces eorum sicut Oreb et Zebet Zebee et Salmana, omnes principes eorum,
PS|83|13|qui dixerunt: Hereditate possideamus pascua Dei! ".
PS|83|14|Deus meus, pone illos ut rotamet sicut stipulam ante ventum.
PS|83|15|Sicut ignis, qui comburit silvam,et sicut flamma devorans montes,
PS|83|16|ita persequeris illos in tempestate tuaet in procella tua turbabis eos.
PS|83|17|Imple facies eorum ignominia,et quaerent nomen tuum, Domine.
PS|83|18|Erubescant et conturbentur in saeculum saeculiet confundantur et pereant;
PS|83|19|et cognoscant quia nomen tibi Dominus:tu solus Altissimus super omnem terram.
PS|84|1|Magistro chori. Secundum " Torcularia ".Filiorum Core. PSALMUS.
PS|84|2|Quam dilecta tabernacula tua, Domine virtutum!
PS|84|3|Concupiscit et deficit anima mea in atria Domini.Cor meum et caro mea exsultaverunt in Deum vivum.
PS|84|4|Etenim passer invenit sibi domum,et turtur nidum sibi, ubi ponat pullos suos:altaria tua, Domine virtutum, rex meus et Deus meus.
PS|84|5|Beati, qui habitant in domo tua:in perpetuum laudabunt te.
PS|84|6|Beatus vir, cuius est auxilium abs te,ascensiones in corde suo disposuit.
PS|84|7|Transeuntes per vallem sitientemin fontem ponent eam,etenim benedictionibus vestiet eam pluvia matutina.
PS|84|8|Ibunt de virtute in virtutem,videbitur Deus deorum in Sion.
PS|84|9|Domine, Deus virtutum, exaudi orationem meam;auribus percipe, Deus Iacob.
PS|84|10|Protector noster aspice, Deus,et respice in faciem christi tui.
PS|84|11|Quia melior est dies una in atriis tuis super milia,elegi ad limen esse in domo Dei meimagis quam habitare in tabernaculis peccatorum.
PS|84|12|Quia sol et scutum est Dominus Deus,gratiam et gloriam dabit Dominus;non privabit bonis eos,qui ambulant in innocentia.
PS|84|13|Domine virtutum, beatus homo, qui sperat in te.
PS|85|1|Magistro chori. Filiorum Core. PSALMUS.
PS|85|2|Complacuisti tibi, Domine, in terra tua,convertisti captivitatem Iacob.
PS|85|3|Remisisti iniquitatem plebis tuae,operuisti omnia peccata eorum.
PS|85|4|Contraxisti omnem iram tuam,revertisti a furore indignationis tuae.
PS|85|5|Converte nos, Deus, salutaris noster,et averte iram tuam a nobis.
PS|85|6|Numquid in aeternum irasceris nobisaut extendes iram tuam a generatione in generationem?
PS|85|7|Nonne tu conversus vivificabis nos,et plebs tua laetabitur in te?
PS|85|8|Ostende nobis, Domine, misericordiam tuamet salutare tuum da nobis.
PS|85|9|Audiam, quid loquatur Dominus Deus,quoniam loquetur pacem ad plebem suam et sanctos suoset ad eos, qui convertuntur corde.
PS|85|10|Vere prope timentes eum salutare ipsius,ut inhabitet gloria in terra nostra.
PS|85|11|Misericordia et veritas obviaverunt sibi,iustitia et pax osculatae sunt.
PS|85|12|Veritas de terra orta est,et iustitia de caelo prospexit.
PS|85|13|Etenim Dominus dabit benignitatem,et terra nostra dabit fructum suum.
PS|85|14|Iustitia ante eum ambulabitet ponet in via gressus suos.
PS|86|1|Precatio. David.Inclina, Domine, aurem tuam et exaudi me,quoniam inops et pauper sum ego.
PS|86|2|Custodi animam meam, quoniam sanctus sum;salvum fac servum tuum, Deus meus, sperantem in te
PS|86|3|Miserere mei, Domine, quoniam ad te clamavi tota die.
PS|86|4|Laetifica animam servi tui,quoniam ad te, Domine, animam meam levavi.
PS|86|5|Quoniam tu, Domine, suavis et mitiset multae misericordiae omnibus invocantibus te. -
PS|86|6|Auribus percipe, Domine, orationem meamet intende voci deprecationis meae.
PS|86|7|In die tribulationis meae clamavi ad te,quia exaudies me.
PS|86|8|Non est similis tui in diis, Domine,et nihil sicut opera tua.
PS|86|9|Omnes gentes, quascumque fecisti, venientet adorabunt coram te, Domine,et glorificabunt nomen tuum,
PS|86|10|quoniam magnus es tu et faciens mirabilia:tu es Deus solus.
PS|86|11|Doce me, Domine, viam tuam,et ingrediar in veritate tua;simplex fac cor meum,ut timeat nomen tuum.
PS|86|12|Confitebor tibi, Domine Deus meus, in toto corde meoet glorificabo nomen tuum in aeternum,
PS|86|13|quia misericordia tua magna est super me,et eruisti animam meam ex inferno inferiori.
PS|86|14|Deus, superbi insurrexerunt super me,et synagoga potentium quaesierunt animam meamet non proposuerunt te in conspectu suo.
PS|86|15|Et tu, Domine, Deus miserator et misericors,patiens et multae misericordiae et veritatis,
PS|86|16|respice in me et miserere mei;da fortitudinem tuam puero tuoet salvum fac filium ancillae tuae.
PS|86|17|Fac mecum signum in bonum,ut videant, qui oderunt me, et confundantur,quoniam tu, Domine, adiuvisti me et consolatus es me.
PS|87|1|Filiorum Core. PSALMUS. Canticum.Fundamenta eius in montibus sanctis;
PS|87|2|diligit Dominus portas Sionsuper omnia tabernacula Iacob.
PS|87|3|Gloriosa dicta sunt de te, civitas Dei! -
PS|87|4|Memor ero Rahab et Babylonis inter scientes me;ecce Philistaea et Tyrus cum Aethiopia:hi nati sunt illic.
PS|87|5|Et de Sion dicetur: " Hic et ille natus est in ea;et ipse firmavit eam Altissimus ".
PS|87|6|Dominus referet in librum populorum: Hi nati sunt illic ".
PS|87|7|Et cantant sicut choros ducentes: Omnes fontes mei in te ".
PS|88|1|Canticum. PSALMUS. Filiorum Core. Magistro chori.Secundum " Mahalat ". Ad cantandum. Maskil. Heman Ezrahitae.
PS|88|2|Domine, Deus salutis meae,in die clamavi et nocte coram te.
PS|88|3|Intret in conspectu tuo oratio mea;inclina aurem tuam ad precem meam.
PS|88|4|Quia repleta est malis anima mea,et vita mea inferno appropinquavit.
PS|88|5|Aestimatus sum cum descendentibus in lacum,factus sum sicut homo sine adiutorio.
PS|88|6|Inter mortuos liber,sicut vulnerati dormientes in sepulcris;quorum non es memor amplius,et ipsi de manu tua abscissi sunt.
PS|88|7|Posuisti me in lacu inferiori,in tenebrosis et in umbra mortis.
PS|88|8|Super me gravatus est furor tuus,et omnes fluctus tuos induxisti super me.
PS|88|9|Longe fecisti notos meos a me,posuisti me abominationem eis;conclusus sum et non egrediar.
PS|88|10|Oculi mei languerunt prae afflictione.Clamavi ad te, Domine, tota die,expandi ad te manus meas. -
PS|88|11|Numquid mortuis facies mirabilia,aut surgent umbrae et confitebuntur tibi?
PS|88|12|Numquid narrabit aliquis in sepulcro misericordiam tuamet veritatem tuam in loco perditionis?
PS|88|13|Numquid cognoscentur in tenebris mirabilia tua,et iustitia tua in terra oblivionis?
PS|88|14|Et ego ad te, Domine, clamavi,et mane oratio mea praeveniet te.
PS|88|15|Ut quid, Domine, repellis animam meam,abscondis faciem tuam a me?
PS|88|16|Pauper sum ego et moriens a iuventute mea;portavi pavores tuos et conturbatus sum.
PS|88|17|Super me transierunt irae tuae,et terrores tui exciderunt me.
PS|88|18|Circuierunt me sicut aqua tota die,circumdederunt me simul.
PS|88|19|Elongasti a me amicum et proximum,et noti mei sunt tenebrae.
PS|89|1|Maskil. Ethan Ezrahitae.
PS|89|2|Misericordias Domini in aeternum cantabo;in generationem et generationemannuntiabo veritatem tuam in ore meo.
PS|89|3|Quoniam dixisti: " In aeternum misericordia aedificabitur ",in caelis firmabitur veritas tua.
PS|89|4|" Disposui testamentum electo meo,iuravi David servo meo:
PS|89|5|Usque in aeternum confirmabo semen tuumet aedificabo in generationem et generationem sedem tuam ".
PS|89|6|Confitebuntur caeli mirabilia tua, Domine,etenim veritatem tuam in ecclesia sanctorum.
PS|89|7|Quoniam quis in nubibus aequabitur Domino,similis erit Domino in filiis Dei?
PS|89|8|Deus, metuendus in consilio sanctorum,magnus et terribilis super omnes, qui in circuitu eius sunt.
PS|89|9|Domine, Deus virtutum, quis similis tibi?Potens es, Domine, et veritas tua in circuitu tuo.
PS|89|10|Tu dominaris superbiae maris,elationes fluctuum eius tu mitigas.
PS|89|11|Tu conculcasti sicut vulneratum Rahab,in brachio virtutis tuae dispersisti inimicos tuos.
PS|89|12|Tui sunt caeli, et tua est terra,orbem terrae et plenitudinem eius tu fundasti;
PS|89|13|Aquilonem et austrum tu creasti,Thabor et Hermon in nomine tuo exsultabunt.
PS|89|14|Tibi brachium cum potentia;firma est manus tua, et exaltata dextera tua.
PS|89|15|Iustitia et iudicium firmamentum sedis tuae.Misericordia et veritas praecedent faciem tuam.
PS|89|16|Beatus populus, qui scit iubilationem.Domine, in lumine vultus tui ambulabunt
PS|89|17|et in nomine tuo exsultabunt tota die et in iustitia tua exaltabuntur,
PS|89|18|quoniam decor virtutis eorum tu es,et in beneplacito tuo exaltabitur cornu nostrum.
PS|89|19|Quia Domini est scutum nostrum,et Sancti Israel rex noster.
PS|89|20|Tunc locutus es in visione sanctis tuis et dixisti: Posui adiutorium in potenteet exaltavi electum de plebe.
PS|89|21|Inveni David servum meum;oleo sancto meo unxi eum.
PS|89|22|Manus enim mea firma erit cum eo, et brachium meum confortabit eum.
PS|89|23|Nihil proficiet inimicus in eo,et filius iniquitatis non opprimet eum.
PS|89|24|Et concidam a facie ipsius inimicos eiuset odientes eum percutiam.
PS|89|25|Et veritas mea et misericordia mea cum ipso,et in nomine meo exaltabitur cornu eius.
PS|89|26|Et ponam super mare manum eiuset super flumina dexteram eius.
PS|89|27|Ipse invocabit me: "Pater meus es tu,Deus meus et refugium salutis meae".
PS|89|28|Et ego primogenitum ponam illum,excelsum prae regibus terrae.
PS|89|29|In aeternum servabo illi misericordiam meam;et testamentum meum fidele ipsi.
PS|89|30|Et ponam in saeculum saeculi semen eius;et thronum eius sicut dies caeli.
PS|89|31|Si autem dereliquerint filii eius legem meamet in iudiciis meis non ambulaverint,
PS|89|32|si iustificationes meas profanaverintet mandata mea non custodierint,
PS|89|33|visitabo in virga delictum eorumet in verberibus iniquitatem eorum.
PS|89|34|Misericordiam autem meam non avertam ab eoneque mentiar in veritate mea.
PS|89|35|Non profanabo testamentum meum et, quae procedunt de labiis meis, non faciam irrita.
PS|89|36|Semel iuravi in sancto meo: David non mentiar.
PS|89|37|Semen eius in aeternum manebit,et thronus eius sicut sol in conspectu meo
PS|89|38|et sicut luna firmus stabit in aeternumet testis in caelo fidelis ".
PS|89|39|Tu vero reppulisti et reiecisti,iratus es contra christum tuum;
PS|89|40|evertisti testamentum servi tui,profanasti in terram diadema eius.
PS|89|41|Destruxisti omnes muros eius,posuisti munitiones eius in ruinas.
PS|89|42|Diripuerunt eum omnes transeuntes viam,factus est opprobrium vicinis suis.
PS|89|43|Exaltasti dexteram deprimentium eum,laetificasti omnes inimicos eius.
PS|89|44|Avertisti aciem gladii eiuset non es auxiliatus ei in bello.
PS|89|45|Finem posuisti splendori eiuset sedem eius in terram collisisti.
PS|89|46|Minorasti dies iuventutis eius,perfudisti eum confusione.
PS|89|47|Usquequo, Domine, absconderis in finem,exardescet sicut ignis ira tua?
PS|89|48|Memorare, quam brevis mea substantia.Ad quam vanitatem creasti omnes filios hominum?
PS|89|49|Quis est homo, qui vivet et non videbit mortem,eruet animam suam de manu inferi?
PS|89|50|Ubi sunt misericordiae tuae antiquae, Domine,sicut iurasti David in veritate tua?
PS|89|51|Memor esto, Domine, opprobrii servorum tuorum,quod continui in sinu meo, multarum gentium,
PS|89|52|quo exprobraverunt inimici tui, Domine,quo exprobraverunt vestigia christi tui.
PS|89|53|Benedictus Dominus in aeternum. Fiat, fiat.
PS|90|1|Precatio. Moysis viri Dei. Domine, refugium factus es nobisa generatione in generationem.
PS|90|2|Priusquam montes nascerentur, aut gigneretur terra et orbis,a saeculo et usque in saeculum tu es Deus.
PS|90|3|Reducis hominem in pulverem;et dixisti: " Revertimini, filii hominum ".
PS|90|4|Quoniam mille anni ante oculos tuostamquam dies hesterna, quae praeteriit,et custodia in nocte.
PS|90|5|Auferes eos, somnium erunt:
PS|90|6|mane sicut herba succrescens,mane floret et crescit,vespere decidit et arescit.
PS|90|7|Quia defecimus in ira tuaet in furore tuo turbati sumus.
PS|90|8|Posuisti iniquitates nostras in conspectu tuo,occulta nostra in illuminatione vultus tui.
PS|90|9|Quoniam omnes dies nostri evanuerunt in ira tua,consumpsimus ut suspirium annos nostros.
PS|90|10|Dies annorum nostrorum sunt septuaginta anniaut in valentibus octoginta anni,et maior pars eorum labor et dolor,quoniam cito transeunt, et avolamus.
PS|90|11|Quis novit potestatem irae tuaeet secundum timorem tuum indignationem tuam?
PS|90|12|Dinumerare dies nostros sic doce nos, ut inducamus cor ad sapientiam.
PS|90|13|Convertere, Domine, usquequo?Et deprecabilis esto super servos tuos.
PS|90|14|Reple nos mane misericordia tua,et exsultabimus et delectabimur omnibus diebus nostris.
PS|90|15|Laetifica nos pro diebus, quibus nos humiliasti,pro annis, quibus vidimus mala.
PS|90|16|Appareat servis tuis opus tuum,et decor tuus filiis eorum.
PS|90|17|Et sit splendor Domini Dei nostri super nos,et opera manuum nostrarum confirma super noset opus manuum nostrarum confirma.
PS|91|1|Qui habitat in protectione Altissimi,sub umbra Omnipotentis commorabitur.
PS|91|2|Dicet Domino: " Refugium meumet fortitudo mea, Deus meus, sperabo in eum ".
PS|91|3|Quoniam ipse liberabit te de laqueo venantiumet a verbo maligno.
PS|91|4|Alis suis obumbrabit tibi,et sub pennas eius confugies;scutum et lorica veritas eius.
PS|91|5|Non timebis a timore nocturno,a sagitta volante in die,
PS|91|6|a peste perambulante in tenebris,ab exterminio vastante in meridie.
PS|91|7|Cadent a latere tuo milleet decem milia a dextris tuis;ad te autem non appropinquabit.
PS|91|8|Verumtamen oculis tuis considerabiset retributionem peccatorum videbis.
PS|91|9|Quoniam tu es, Domine, refugium meum.Altissimum posuisti habitaculum tuum.
PS|91|10|Non accedet ad te malum,et flagellum non appropinquabit tabernaculo tuo,
PS|91|11|quoniam angelis suis mandabit de te,ut custodiant te in omnibus viis tuis.
PS|91|12|In manibus portabunt te,ne forte offendas ad lapidem pedem tuum.
PS|91|13|Super aspidem et basiliscum ambulabiset conculcabis leonem et draconem.
PS|91|14|Quoniam mihi adhaesit, liberabo eum;suscipiam eum, quoniam cognovit nomen meum.
PS|91|15|Clamabit ad me, et ego exaudiam eum;cum ipso sum in tribulatione;eripiam eum et glorificabo eum.
PS|91|16|Longitudine dierum replebo eumet ostendam illi salutare meum.
PS|92|1|PSALMUS. Canticum. Pro die Sabbati.
PS|92|2|Bonum est confiteri Dominoet psallere nomini tuo, Altissime,
PS|92|3|annuntiare mane misericordiam tuamet veritatem tuam per noctem
PS|92|4|in decachordo et psalterio,cum cantico in cithara.
PS|92|5|Quia delectasti me, Domine, in factura tua,et in operibus manuum tuarum exsultabo.
PS|92|6|Quam magnificata sunt opera tua, Domine:nimis profundae factae sunt cogitationes tuae.
PS|92|7|Vir insipiens non cognoscet,et stultus non intelleget haec.
PS|92|8|Cum germinaverint peccatores sicut fenum,et floruerint omnes, qui operantur iniquitatem,hoc tamen erit ad interitum in saeculum saeculi;
PS|92|9|tu autem altissimus in aeternum, Domine.
PS|92|10|Quoniam ecce inimici tui, Domine,quoniam ecce inimici tui peribunt,et dispergentur omnes, qui operantur iniquitatem.
PS|92|11|Exaltabis sicut unicornis cornu meum,perfusus sum oleo uberi.
PS|92|12|Et despiciet oculus meus inimicos meos,et in insurgentibus in me malignantibus audiet auris mea. -
PS|92|13|Iustus ut palma florebit,sicut cedrus Libani succrescet.
PS|92|14|Plantati in domo Domini,in atriis Dei nostri florebunt.
PS|92|15|Adhuc fructus dabunt in senecta,uberes et bene virentes erunt,
PS|92|16|ut annuntient quoniam rectus Dominus,refugium meum, et non est iniquitas in eo.
PS|93|1|Dominus regnavit! Decorem indutus est;indutus est Dominus, fortitudine praecinxit se.Etenim firmavit orbem terrae, qui non commovebitur.
PS|93|2|Firmata sedes tua ex tunc,a saeculo tu es.
PS|93|3|Elevaverunt flumina, Domine.elevaverunt flumina vocem suam,elevaverunt flumina fragorem suum.
PS|93|4|Super voces aquarum multarum,super potentes elationes maris,potens in altis Dominus.
PS|93|5|Testimonia tua credibilia facta sunt nimis;domum tuam decet sanctitudo Domine,in longitudinem dierum.
PS|94|1|Deus ultionum, Domine,Deus ultionum, effulge.
PS|94|2|Exaltare, qui iudicas terram,redde retributionem superbis.
PS|94|3|Usquequo peccatores, Domine,usquequo peccatores exsultabunt?
PS|94|4|Effabuntur et loquentur proterva,gloriabuntur omnes, qui operantur iniquitatem. -
PS|94|5|Populum tuum, Domine, humiliantet hereditatem tuam vexant.
PS|94|6|Viduam et advenam interficiuntet pupillos occidunt.
PS|94|7|Et dixerunt: " Non videbit Dominus,nec intelleget Deus Iacob ".
PS|94|8|Intellegite, insipientes in populo;et stulti, quando sapietis?
PS|94|9|Qui plantavit aurem, non audiet,aut qui finxit oculum, non respiciet?
PS|94|10|Qui corripit gentes, non arguet,qui docet hominem scientiam?
PS|94|11|Dominus scit cogitationes hominum,quoniam vanae sunt.
PS|94|12|Beatus homo, quem tu erudieris, Domine,et de lege tua docueris eum,
PS|94|13|ut mitiges ei a diebus malis,donec fodiatur peccatori fovea.
PS|94|14|Quia non repellet Dominus plebem suamet hereditatem suam non derelinquet.
PS|94|15|Quia ad iustitiam revertetur iudicium,et sequentur illam omnes, qui recto sunt corde.
PS|94|16|Quis consurget mihi adversus malignantes,aut quis stabit mecum adversus operantes iniquitatem?
PS|94|17|Nisi quia Dominus adiuvit me,paulo minus habitasset in loco silentii anima mea.
PS|94|18|Si dicebam: " Motus est pes meus ", misericordia tua, Domine, sustentabat me.
PS|94|19|In multitudine sollicitudinum mearum in corde meo,consolationes tuae laetificaverunt animam meam.
PS|94|20|Numquid sociabitur tibi sedes iniquitatis,quae fingit molestiam contra praeceptum?
PS|94|21|Irruunt in animam iustiet sanguinem innocentem condemnant.
PS|94|22|Et factus est mihi Dominus in praesidium,et Deus meus in rupem refugii mei;
PS|94|23|et reddet illis iniquitatem ipsorumet in malitia eorum disperdet eos,
PS|94|24|disperdet illos Dominus Deus noster.
PS|95|1|Venite, exsultemus Domino;iubilemus Deo salutari nostro.
PS|95|2|Praeoccupemus faciem eius in confessioneet in psalmis iubilemus ei.
PS|95|3|Quoniam Deus magnus Dominus,et rex magnus super omnes deos.
PS|95|4|Quia in manu eius sunt profunda terrae,et altitudines montium ipsius sunt.
PS|95|5|Quoniam ipsius est mare, et ipse fecit illud,et siccam manus eius formaverunt.
PS|95|6|Venite, adoremus et procidamuset genua flectamus ante Dominum, qui fecit nos,
PS|95|7|quia ipse est Deus noster,et nos populus pascuae eius et oves manus eius.
PS|95|8|Utinam hodie vocem eius audiatis: Nolite obdurare corda vestra,
PS|95|9|sicut in Meriba, secundum diem Massa in deserto,ubi tentaverunt me patres vestri:probaverunt me, etsi viderunt opera mea.
PS|95|10|Quadraginta annis taeduit me generationis illiuset dixi: Populus errantium corde sunt isti.
PS|95|11|Et ipsi non cognoverunt vias meas;ideo iuravi in ira mea:Non introibunt in requiem meam ".
PS|96|1|Cantate Domino canticum novum,cantate Domino, omnis terra.
PS|96|2|Cantate Domino, benedicite nomini eius,annuntiate de die in diem salutare eius.
PS|96|3|Annuntiate inter gentes gloriam eius,in omnibus populis mirabilia eius.
PS|96|4|Quoniam magnus Dominus et laudabilis nimis,terribilis est super omnes deos.
PS|96|5|Quoniam omnes dii gentium inania,Dominus autem caelos fecit.
PS|96|6|Magnificentia et pulchritudo in conspectu eius,potentia et decor in sanctuario eius.
PS|96|7|Afferte Domino, familiae populorum,afferte Domino gloriam et potentiam,
PS|96|8|afferte Domino gloriam nominis eius.Tollite hostias et introite in atria eius,
PS|96|9|adorate Dominum in splendore sancto.Contremiscite a facie eius, universa terra;
PS|96|10|dicite in gentibus: " Dominus regnavit! ".Etenim correxit orbem terrae, qui non commovebitur;iudicabit populos in aequitate.
PS|96|11|Laetentur caeli, et exsultet terra,sonet mare et plenitudo eius;
PS|96|12|gaudebunt campi et omnia, quae in eis sunt.Tunc exsultabunt omnia ligna silvarum
PS|96|13|a facie Domini, quia venit,quoniam venit iudicare terram.Iudicabit orbem terrae in iustitiaet populos in veritate sua.
PS|97|1|Dominus regnavit! Exsultet terra,laetentur insulae multae.
PS|97|2|Nubes et caligo in circuitu eius,iustitia et iudicium firmamentum sedis eius.
PS|97|3|Ignis ante ipsum praecedetet inflammabit in circuitu inimicos eius.
PS|97|4|Illustrarunt fulgura eius orbem terrae:vidit et contremuit terra.
PS|97|5|Montes sicut cera fluxerunt a facie Domini,a facie Domini omnis terra.
PS|97|6|Annuntiaverunt caeli iustitiam eius,et viderunt omnes populi gloriam eius.
PS|97|7|Confundantur omnes, qui adorant sculptilia,et qui gloriantur in simulacris suis.Adorate eum, omnes angeli eius.
PS|97|8|Audivit et laetata est Sion,et exsultaverunt filiae Iudaepropter iudicia tua, Domine.
PS|97|9|Quoniam tu Dominus, Altissimus super omnem terram,nimis exaltatus es super omnes deos.
PS|97|10|Qui diligitis Dominum, odite malum;custodit ipse animas sanctorum suorum,de manu peccatoris liberabit eos.
PS|97|11|Lux orta est iusto,et rectis corde laetitia.
PS|97|12|Laetamini, iusti, in Dominoet confitemini memoriae sanctitatis eius.
PS|98|1|PSALMUS.Cantate Domino canticum novum,quia mirabilia fecit.Salvavit sibi dextera eius,et brachium sanctum eius.
PS|98|2|Notum fecit Dominus salutare suum,in conspectu gentium revelavit iustitiam suam.
PS|98|3|Recordatus est misericordiae suaeet veritatis suae domui Israel.Viderunt omnes termini terraesalutare Dei nostri.
PS|98|4|Iubilate Deo, omnis terra;erumpite, exsultate et psallite.
PS|98|5|Psallite Domino in cithara,in cithara et voce psalmi;
PS|98|6|in tubis ductilibus et voce tubae corneae,iubilate in conspectu regis Domini.
PS|98|7|Sonet mare et plenitudo eius,orbis terrarum et qui habitant in eo.
PS|98|8|Flumina plaudent manu,simul montes exsultabunt
PS|98|9|a conspectu Domini, quoniam venit iudicare terram.Iudicabit orbem terrarum in iustitiaet populos in aequitate.
PS|99|1|Dominus regnavit! Commoveantur populisedet super cherubim, moveatur terra.
PS|99|2|Dominus in Sion magnuset excelsus super omnes populos.
PS|99|3|Confiteantur nomini tuo magno et terribili,quoniam sanctum est.
PS|99|4|Rex potens iudicium diligit:tu statuisti, quae recta sunt,iudicium et iustitiam in Iacob tu fecisti.
PS|99|5|Exaltate Dominum Deum nostrumet adorate ad scabellum pedum eius,quoniam sanctus est.
PS|99|6|Moyses et Aaron in sacerdotibus eius,et Samuel inter eos, qui invocant nomen eius.Invocabant Dominum, et ipse exaudiebat eos,
PS|99|7|in columna nubis loquebatur ad eos.Custodiebant testimonia eiuset praeceptum, quod dedit illis.
PS|99|8|Domine Deus noster, tu exaudiebas eos;Deus, tu propitius fuisti eis,ulciscens autem adinventiones eorum.
PS|99|9|Exaltate Dominum Deum nostrumet adorate ad montem sanctum eius,quoniam sanctus Dominus Deus noster.
PS|100|1|PSALMUS. Ad gratiarum actionem.
PS|100|2|Iubilate Domino, omnis terra,servite Domino in laetitia;introite in conspectu eius in exsultatione.
PS|100|3|Scitote quoniam Dominus ipse est Deus;ipse fecit nos, et ipsius sumus,populus eius et oves pascuae eius.
PS|100|4|Introite portas eius in confessione,atria eius in hymnis,confitemini illi, benedicite nomini eius.
PS|100|5|Quoniam suavis est Dominus;in aeternum misericordia eius,et usque in generationem et generationem veritas eius.
PS|101|1|David. PSALMUS.Misericordiam et iudicium cantabo;tibi, Domine, psallam.
PS|101|2|Intellegam in via immaculata;quando venies ad me?Perambulabo in innocentia cordis mei,in medio domus meae.
PS|101|3|Non proponam ante oculos meos rem iniustam;facientem praevaricationes odio habebo,non adhaerebit mihi.
PS|101|4|Cor pravum recedet a me,malignum non cognoscam.
PS|101|5|Detrahentem secreto proximo suo,hunc cessare faciam;superbum oculo et inflatum corde,hunc non sustinebo.
PS|101|6|Oculi mei ad fideles terrae, ut sedeant mecum;qui ambulat in via immaculata, hic mihi ministrabit.
PS|101|7|Non habitabit in medio domus meae, qui facit superbiam;qui loquitur iniqua, non stabit in conspectu oculorum meorum.
PS|101|8|In matutino cessare faciam omnes peccatores terrae,ut disperdam de civitate Domini omnes operantes iniquitatem.
PS|102|1|Preces afflicti, qui defessusangorem suum ante Dominum profundit.
PS|102|2|Domine, exaudi orationem meam,et clamor meus ad te veniat.
PS|102|3|Non abscondas faciem tuam a me;in quacumque die tribulor,inclina ad me aurem tuam.In quacumque die invocavero te,velociter exaudi me.
PS|102|4|Quia defecerunt sicut fumus dies mei,et ossa mea sicut cremium aruerunt.
PS|102|5|Percussum est ut fenum et aruit cor meum,etenim oblitus sum comedere panem meum.
PS|102|6|A voce gemitus meiadhaesit os meum carni meae.
PS|102|7|Similis factus sum pellicano solitudinis,factus sum sicut nycticorax in ruinis.
PS|102|8|Vigilavi et factus sum sicut passer solitarius in tecto.
PS|102|9|Tota die exprobrabant mihi inimici mei,exardescentes in me per me iurabant.
PS|102|10|Quia cinerem tamquam panem manducabamet potum meum cum fletu miscebam,
PS|102|11|a facie irae et increpationis tuae,quia elevans allisisti me.
PS|102|12|Dies mei sicut umbra declinaverunt,et ego sicut fenum arui.
PS|102|13|Tu autem, Domine, in aeternum permanes,et memoriale tuum in generationem et generationem.
PS|102|14|Tu exsurgens misereberis Sion,quia tempus miserendi eius,quia venit tempus,
PS|102|15|quoniam placuerunt servis tuis lapides eius,et pulveris eius miserentur.
PS|102|16|Et timebunt gentes nomen tuum, Domine,et omnes reges terrae gloriam tuam,
PS|102|17|quia aedificavit Dominus Sionet apparuit in gloria sua.
PS|102|18|Respexit in orationem inopumet non sprevit precem eorum.
PS|102|19|Scribantur haec pro generatione altera,et populus, qui creabitur, laudabit Dominum.
PS|102|20|Quia prospexit de excelso sanctuario suo,Dominus de caelo in terram aspexit,
PS|102|21|ut audiret gemitus compeditorum, ut solveret filios mortis;
PS|102|22|ut annuntient in Sion nomen Dominiet laudem eius in Ierusalem,
PS|102|23|cum congregati fuerint populi in unumet regna, ut serviant Domino.
PS|102|24|Humiliavit in via virtutem meam,abbreviavit dies meos.Dicam: " Deus meus,
PS|102|25|ne auferas me in dimidio dierum meorum;in generationem et generationem sunt anni tui.
PS|102|26|Initio terram fundasti;et opera manuum tuarum sunt caeli.
PS|102|27|Ipsi peribunt, tu autem permanes;et omnes sicut vestimentum veterascent,et sicut opertorium mutabis eos, et mutabuntur.
PS|102|28|Tu autem idem ipse es, et anni tui non deficient.
PS|102|29|Filii servorum tuorum habitabunt,et semen eorum in conspectu tuo firmabitur ".
PS|103|1|David.Benedic, anima mea, Domino,et omnia, quae intra me sunt, nomini sancto eius.
PS|103|2|Benedic, anima mea, Dominoet noli oblivisci omnes retributiones eius.
PS|103|3|Qui propitiatur omnibus iniquitatibus tuis,qui sanat omnes infirmitates tuas;
PS|103|4|qui redimit de interitu vitam tuam,qui coronat te in misericordia et miserationibus;
PS|103|5|qui replet in bonis aetatem tuam:renovabitur ut aquilae iuventus tua.
PS|103|6|Faciens iustitias Dominuset iudicium omnibus iniuriam patientibus.
PS|103|7|Notas fecit vias suas Moysi,filiis Israel adinventiones suas. -
PS|103|8|Miserator et misericors Dominus,longanimis et multae misericordiae.
PS|103|9|Non in perpetuum contendetneque in aeternum irascetur.
PS|103|10|Non secundum peccata nostra fecit nobisneque secundum iniquitates nostras retribuit nobis.
PS|103|11|Quoniam, quantum exaltatur caelum a terra,praevaluit misericordia eius super timentes eum;
PS|103|12|quantum distat ortus ab occidente,longe fecit a nobis iniquitates nostras.
PS|103|13|Quomodo miseretur pater filiorum,misertus est Dominus timentibus se.
PS|103|14|Quoniam ipse cognovit figmentum nostrum,recordatus est quoniam pulvis sumus.
PS|103|15|Homo: sicut fenum dies eius,tamquam flos agri sic efflorebit.
PS|103|16|Spirat ventus in illum, et non subsistet,et non cognoscet eum amplius locus eius.
PS|103|17|Misericordia autem Domini ab aeternoet usque in aeternum super timentes eum;et iustitia illius in filios filiorum,
PS|103|18|in eos, qui servant testamentum eiuset memores sunt mandatorum ipsius ad faciendum ea.
PS|103|19|Dominus in caelo paravit sedem suam,et regnum ipsius omnibus dominabitur.
PS|103|20|Benedicite Domino, omnes angeli eius, potentes virtute, facientes verbum illiusin audiendo vocem sermonum eius.
PS|103|21|Benedicite Domino, omnes virtutes eius,ministri eius, qui facitis voluntatem eius.
PS|103|22|Benedicite Domino, omnia opera eius,in omni loco dominationis eius.Benedic, anima mea, Domino.
PS|104|1|Benedic, anima mea, Domino.Domine Deus meus, magnificatus es vehementer!Maiestatem et decorem induisti,
PS|104|2|amictus lumine sicut vestimento.Extendens caelum sicut velum,
PS|104|3|qui exstruis in aquis cenacula tua.Qui ponis nubem ascensum tuum,qui ambulas super pennas ventorum.
PS|104|4|Qui facis angelos tuos spirituset ministros tuos ignem urentem.
PS|104|5|Qui fundasti terram super stabilitatem suam,non inclinabitur in saeculum saeculi.
PS|104|6|Abyssus sicut vestimentum operuit eam,super montes stabant aquae.
PS|104|7|Ab increpatione tua fugiunt,a voce tonitrui tui formidant.
PS|104|8|Ascendunt in montes et descendunt in valles,in locum, quem statuisti eis.
PS|104|9|Terminum posuisti, quem non transgredientur,neque convertentur operire terram.
PS|104|10|Qui emittis fontes in torrentes;inter medium montium pertransibunt,
PS|104|11|potabunt omnes bestias agri,exstinguent onagri sitim suam.
PS|104|12|Super ea volucres caeli habitabunt,de medio ramorum dabunt voces.
PS|104|13|Rigas montes de cenaculis tuis,de fructu operum tuorum satias terram.
PS|104|14|Producis fenum iumentiset herbam servituti hominum,educens panem de terra
PS|104|15|et vinum, quod laetificat cor hominis;exhilarans faciem in oleo,panis autem cor hominis confirmat.
PS|104|16|Saturabuntur ligna Dominiet cedri Libani, quas plantavit.
PS|104|17|Illic passeres nidificabunt,erodii domus in vertice earum.
PS|104|18|Montes excelsi cervis,petrae refugium hyracibus.
PS|104|19|Fecit lunam ad tempora signanda,sol cognovit occasum suum.
PS|104|20|Posuisti tenebras, et facta est nox:in ipsa reptabunt omnes bestiae silvae,
PS|104|21|catuli leonum rugientes, ut rapiantet quaerant a Deo escam sibi.
PS|104|22|Oritur sol, et congreganturet in cubilibus suis recumbunt.
PS|104|23|Exit homo ad opus suumet ad operationem suam usque ad vesperum.
PS|104|24|Quam multiplicata sunt opera tua, Domine!Omnia in sapientia fecisti,impleta est terra creatura tua.
PS|104|25|Hoc mare magnum et spatiosum et latum:illic reptilia, quorum non est numerus,animalia pusilla cum magnis;
PS|104|26|illic naves pertransibunt,Leviathan, quem formasti ad ludendum cum eo.
PS|104|27|Omnia a te exspectant,ut des illis escam in tempore suo.
PS|104|28|Dante te illis, colligent,aperiente te manum tuam, implebuntur bonis.
PS|104|29|Avertente autem te faciem, turbabuntur;auferes spiritum eorum, et deficientet in pulverem suum revertentur.
PS|104|30|Emittes spiritum tuum, et creabuntur,et renovabis faciem terrae.
PS|104|31|Sit gloria Domini in saeculum;laetetur Dominus in operibus suis.
PS|104|32|Qui respicit terram et facit eam tremere,qui tangit montes, et fumigant.
PS|104|33|Cantabo Domino in vita mea,psallam Deo meo quamdiu sum.
PS|104|34|Iucundum sit ei eloquium meum,ego vero delectabor in Domino.
PS|104|35|Deficiant peccatores a terraet iniqui, ita ut non sint.Benedic, anima mea, Domino.
PS|105|1|ALLELUIA.Confitemini Domino et invocate nomen eius,annuntiate inter gentes opera eius.
PS|105|2|Cantate ei et psallite ei,meditamini in omnibus mirabilibus eius.
PS|105|3|Laudamini in nomine sancto eius,laetetur cor quaerentium Dominum.
PS|105|4|Quaerite Dominum et potentiam eius,quaerite faciem eius semper.
PS|105|5|Mementote mirabilium eius, quae fecit,prodigia eius et iudicia oris eius,
PS|105|6|semen Abraham, servi eius,filii Iacob, electi eius.
PS|105|7|Ipse Dominus Deus noster;in universa terra iudicia eius.
PS|105|8|Memor fuit in saeculum testamenti sui,verbi, quod mandavit in mille generationes,
PS|105|9|quod disposuit cum Abraham,et iuramenti sui ad Isaac.
PS|105|10|Et statuit illud Iacob in praeceptumet Israel in testamentum aeternum
PS|105|11|dicens: " Tibi dabo terram Chanaanfuniculum hereditatis vestrae ".
PS|105|12|Cum essent numero brevi,paucissimi et peregrini in ea,
PS|105|13|et pertransirent de gente in gentemet de regno ad populum alterum,
PS|105|14|non permisit hominem nocere eiset corripuit pro eis reges:
PS|105|15|" Nolite tangere christos meoset in prophetis meis nolite malignari ".
PS|105|16|Et vocavit famem super terramet omne baculum panis contrivit.
PS|105|17|Misit ante eos virum,in servum venumdatus est Ioseph.
PS|105|18|Strinxerunt in compedibus pedes eius,in ferrum intravit collum eius,
PS|105|19|donec veniret verbum eius,eloquium Domini purgaret eum.
PS|105|20|Misit rex et solvit eum,princeps populorum, et dimisit eum;
PS|105|21|constituit eum dominum domus suaeet principem omnis possessionis suae,
PS|105|22|ut erudiret principes eius sicut semetipsumet senes eius prudentiam doceret.
PS|105|23|Et intravit Israel in Aegyptum,et Iacob peregrinus fuit in terra Cham.
PS|105|24|Et auxit populum suum vehementeret confortavit eum super inimicos eius.
PS|105|25|Convertit cor eorum, ut odirent populum eiuset dolum facerent in servos eius.
PS|105|26|Misit Moysen servum suum,Aaron, quem elegit.
PS|105|27|Posuit in eis verba signorum suorumet prodigiorum in terra Cham.
PS|105|28|Misit tenebras et obscuravit,et restiterunt sermonibus eius.
PS|105|29|Convertit aquas eorum in sanguinemet occidit pisces eorum.
PS|105|30|Edidit terra eorum ranasin penetralibus regum ipsorum.
PS|105|31|Dixit, et venit coenomyiaet scinifes in omnibus finibus eorum.
PS|105|32|Posuit pluvias eorum grandinem,ignem comburentem in terra ipsorum.
PS|105|33|Et percussit vineas eorum et ficulneas eorumet contrivit lignum finium eorum.
PS|105|34|Dixit, et venit locustaet bruchus, cuius non erat numerus,
PS|105|35|et comedit omne fenum in terra eorumet comedit fructum terrae eorum.
PS|105|36|Et percussit omne primogenitum in terra eorum,primitias omnis roboris eorum.
PS|105|37|Et eduxit eos cum argento et auro;et non erat in tribubus eorum infirmus.
PS|105|38|Laetata est Aegyptus in profectione eorum,quia incubuit timor eorum super eos.
PS|105|39|Expandit nubem in protectionemet ignem, ut luceret eis per noctem.
PS|105|40|Petierunt, et venit coturnix,et pane caeli saturavit eos.
PS|105|41|Dirupit petram, et fluxerunt aquae,abierunt in sicco flumina.
PS|105|42|Quoniam memor fuit verbi sancti suiad Abraham puerum suum.
PS|105|43|Et eduxit populum suum in exsultatione,electos suos in laetitia.
PS|105|44|Et dedit illis regiones gentium,et labores populorum possederunt,
PS|105|45|ut custodiant iustificationes eiuset leges eius servent.ALLELUIA.
PS|106|1|ALLELUIA.Confitemini Domino, quoniam bonus,quoniam in saeculum misericordia eius.
PS|106|2|Quis loquetur potentias Domini,auditas faciet omnes laudes eius?
PS|106|3|Beati, qui custodiunt iudiciumet faciunt iustitiam in omni tempore.
PS|106|4|Memento nostri, Domine, in beneplacito populi tui,visita nos in salutari tuo,
PS|106|5|ut videamus bona electorum tuorum,ut laetemur in laetitia gentis tuae,ut gloriemur cum hereditate tua.
PS|106|6|Peccavimus cum patribus nostris,iniuste egimus, iniquitatem fecimus.
PS|106|7|Patres nostri in Aegypto non intellexerunt mirabilia tua,non fuerunt memores multitudinis misericordiarum tuarumet irritaverunt ascendentes in mare, mare Rubrum.
PS|106|8|Et salvavit eos propter nomen suum,ut notam faceret potentiam suam. -
PS|106|9|Et increpuit mare Rubrum, et exsiccatum est,et deduxit eos in abyssis sicut in deserto.
PS|106|10|Et salvavit eos de manu odientiset redemit eos de manu inimici.
PS|106|11|Et operuit aqua tribulantes eos:unus ex eis non remansit.
PS|106|12|Et crediderunt verbis eiuset cantaverunt laudem eius.
PS|106|13|Cito obliti sunt operum eiuset non sustinuerunt consilium eius;
PS|106|14|et concupierunt concupiscentiam in desertoet tentaverunt Deum in inaquoso.
PS|106|15|Et dedit eis petitionem ipsorumet misit saturitatem in animas eorum.
PS|106|16|Et zelati sunt Moysen in castris,Aaron sanctum Domini.
PS|106|17|Aperta est terra et deglutivit Dathanet operuit super congregationem Abiram.
PS|106|18|Et exarsit ignis in synagoga eorum,flamma combussit peccatores.
PS|106|19|Et fecerunt vitulum in Horebet adoraverunt sculptile;
PS|106|20|et mutaverunt gloriam suamin similitudinem tauri comedentis fenum.
PS|106|21|Obliti sunt Deum, qui salvavit eos,qui fecit magnalia in Aegypto,
PS|106|22|mirabilia in terra Cham,terribilia in mari Rubro.
PS|106|23|Et dixit quia disperderet eos,nisi affuisset Moyses electus eius:stetit in confractione in conspectu eius,ut averteret iram eius, ne destrueret eos.
PS|106|24|Et pro nihilo habuerunt terram desiderabilem,non crediderunt verbo eius.
PS|106|25|Et murmuraverunt in tabernaculis suis,non exaudierunt vocem Domini.
PS|106|26|Et elevavit manum suam super eos,ut prosterneret eos in deserto
PS|106|27|et ut deiceret semen eorum in nationibuset dispergeret eos in regionibus.
PS|106|28|Et adhaeserunt Baalphegoret comederunt sacrificia mortuorum;
PS|106|29|et irritaverunt eum in adinventionibus suis,et irrupit in eos ruina.
PS|106|30|Et stetit Phinees et fecit iudicium,et cessavit quassatio,
PS|106|31|et reputatum est ei in iustitiamin generationem et generationem usque in sempiternum.
PS|106|32|Et irritaverunt eum ad aquas Meriba,et vexatus est Moyses propter eos,
PS|106|33|quia exacerbaverunt spiritum eius,et temere locutus est in labiis suis.
PS|106|34|Non disperdiderunt gentes,quas dixit Dominus illis.
PS|106|35|Et commixti sunt inter genteset didicerunt opera eorum.
PS|106|36|Et servierunt sculptilibus eorum,et factum est illis in scandalum.
PS|106|37|Et immolaverunt filios suoset filias suas daemoniis.
PS|106|38|Et effuderunt sanguinem innocentem,sanguinem filiorum suorum et filiarum suarum,quas sacrificaverunt sculptilibus Chanaan.Et infecta est terra in sanguinibus,
PS|106|39|et contaminati sunt in operibus suiset fornicati sunt in adinventionibus suis.
PS|106|40|Et exarsit ira Dominus in populum suumet abominatus est hereditatem suam
PS|106|41|et tradidit eos in manus gentium,et dominati sunt eorum, qui oderunt eos.
PS|106|42|Et tribulaverunt eos inimici eorum,et humiliati sunt sub manibus eorum.
PS|106|43|Saepe liberavit eos;ipsi autem exacerbaverunt eum in consilio suoet corruerunt in iniquitatibus suis.
PS|106|44|Et vidit tribulationem eorum,cum audivit clamorem eorum. -
PS|106|45|Et memor fuit testamenti suiet paenituit eum secundum multitudinem misericordiae suae.
PS|106|46|Et dedit eos in miserationesin conspectu omnium, qui captivos duxerant eos.
PS|106|47|Salvos nos fac, Domine Deus noster,et congrega nos de nationibus,ut confiteamur nomini sancto tuoet gloriemur in laude tua.
PS|106|48|Benedictus Dominus, Deus Israel, a saeculo et usque in saeculum.Et dicet omnis populus: "Fiat, fiat".
PS|107|1|ALLELUIA. Confitemini Domino, quoniam bonus, quoniam in saeculum misericordia eius.
PS|107|2|Dicant, qui redempti sunt a Domino,quos redemit de manu adversarii
PS|107|3|et de regionibus congregavit eos,a solis ortu et occasu,ab aquilone et mari.
PS|107|4|Erraverunt in solitudine, in inaquoso,viam civitatis habitationis non invenerunt.
PS|107|5|Esurientes et sitientes,anima eorum in ipsis defecit.
PS|107|6|Et clamaverunt ad Dominum, cum tribularentur,et de necessitatibus eorum eripuit eos.
PS|107|7|Et deduxit eos in viam rectam,ut irent in civitatem habitationis.
PS|107|8|Confiteantur Domino propter misericordiam eiuset mirabilia eius in filios hominum,
PS|107|9|quia satiavit animam sitientemet animam esurientem replevit bonis.
PS|107|10|Sedentes in tenebris et umbra mortis,vincti in mendicitate et ferro,
PS|107|11|quia exacerbaverunt eloquia Deiet consilium Altissimi spreverunt.
PS|107|12|Et humiliavit in laboribus cor eorum,infirmati sunt, nec fuit qui adiuvaret.
PS|107|13|Et clamaverunt ad Dominum, cum tribularentur,et de necessitatibus eorum liberavit eos.
PS|107|14|Et eduxit eos de tenebris et umbra mortiset vincula eorum dirupit.
PS|107|15|Confiteantur Domino propter misericordiam eiuset mirabilia eius in filios hominum,
PS|107|16|quia contrivit portas aereaset vectes ferreos confregit.
PS|107|17|Stulti facti sunt in via iniquitatis suaeet propter iniustitias suas afflicti sunt;
PS|107|18|omnem escam abominata est anima eorum,et appropinquaverunt usque ad portas mortis.
PS|107|19|Et clamaverunt ad Dominum, cum tribularentur,et de necessitatibus eorum liberavit eos.
PS|107|20|Misit verbum suum et sanavit eoset eripuit eos de interitionibus eorum.
PS|107|21|Confiteantur Domino propter misericordiam eiuset mirabilia eius in filios hominum;
PS|107|22|et sacrificent sacrificium laudiset annuntient opera eius in exsultatione.
PS|107|23|Qui descendunt mare in navibus,facientes operationem in aquis multis,
PS|107|24|ipsi viderunt opera Dominiet mirabilia eius in profundo.
PS|107|25|Dixit et excitavit spiritum procellae,et exaltati sunt fluctus eius.
PS|107|26|Ascendunt usque ad caeloset descendunt usque ad abyssos;anima eorum in malis tabescebat.
PS|107|27|Turbati sunt et moti sunt sicut ebrius,et omnis sapientia eorum devorata est.
PS|107|28|Et clamaverunt ad Dominum, cum tribularentur,et de necessitatibus eorum eduxit eos.
PS|107|29|Et statuit procellam eius in auram,et tacuerunt fluctus eius.
PS|107|30|Et laetati sunt, quia siluerunt,et deduxit eos in portum voluntatis eorum.
PS|107|31|Confiteantur Domino propter misericordiam eiuset mirabilia eius in filios hominum;
PS|107|32|et exaltent eum in ecclesia plebiset in conventu seniorum laudent eum.
PS|107|33|Posuit flumina in desertumet exitus aquarum in sitim,
PS|107|34|terram fructiferam in salsuginema malitia inhabitantium in ea.
PS|107|35|Posuit desertum in stagna aquarumet terram sine aqua in exitus aquarum.
PS|107|36|Et collocavit illic esurientes,et constituerunt civitatem habitationis.
PS|107|37|Et seminaverunt agros et plantaverunt vineas,et fecerunt fructum in proventum suum.
PS|107|38|Et benedixit eis, et multiplicati sunt nimis,et iumenta eorum non minoravit.
PS|107|39|Et pauci facti sunt et vexati sunta tribulatione malorum et dolore.
PS|107|40|Effudit contemptionem super principeset errare fecit eos in deserto invio.
PS|107|41|Et suscepit pauperem de inopiaet posuit sicut oves familias.
PS|107|42|Videbunt recti et laetabuntur,et omnis iniquitas oppilabit os suum.
PS|107|43|Quis sapiens, et custodiet haecet intelleget misericordias Domini?.
PS|108|1|Canticum. PSALMUS. David.
PS|108|2|Paratum cor meum, Deus,paratum cor meum,cantabo et psallam. Euge, gloria mea!
PS|108|3|Exsurge, psalterium et cithara,excitabo auroram.
PS|108|4|Confitebor tibi in populis, Domine,et psallam tibi in nationibus,
PS|108|5|quia magna est usque ad caelos misericordia tua,et usque ad nubes veritas tua.
PS|108|6|Exaltare super caelos, Deus,et super omnem terram gloria tua.
PS|108|7|Ut liberentur dilecti tui,salvum fac dextera tua et exaudi me.
PS|108|8|Deus locutus est in sancto suo: Exsultabo et dividam Sichimamet convallem Succoth dimetiar;
PS|108|9|meus est Galaad, et meus est Manasses,et Ephraim fortitudo capitis mei,Iuda sceptrum meum.
PS|108|10|Moab lebes lavacri mei;super Idumaeam extendam calceamentum meum,super Philistaeam vociferabor ".
PS|108|11|Quis deducet me in civitatem munitam?Quis deducet me usque in Idumaeam?.
PS|108|12|Nonne, Deus, qui reppulisti nos?Et non exibis, Deus, in virtutibus nostris?
PS|108|13|Da nobis auxilium de tribulatione,quia vana salus hominis.
PS|108|14|In Deo faciemus virtutem,et ipse conculcabit inimicos nostros.
PS|109|1|Magistro chori. David. PSALMUS.Deus laudis meae, ne tacueris,
PS|109|2|quia os peccatoris et os dolosi super me apertum est.Locuti sunt adversum me lingua dolosa
PS|109|3|et sermonibus odii circumdederunt meet expugnaverunt me gratis.
PS|109|4|Pro dilectione mea adversabantur mihi;ego autem orabam.
PS|109|5|Et posuerunt adversum me mala pro boniset odium pro dilectione mea.
PS|109|6|Constitue super eum peccatorem,et adversarius stet a dextris eius.
PS|109|7|Cum iudicatur, exeat condemnatus,et oratio eius fiat in peccatum.
PS|109|8|Fiant dies eius pauci,et ministerium eius accipiat alter.
PS|109|9|Fiant filii eius orphani,et uxor eius vidua.
PS|109|10|Instabiles vagentur filii eius et mendicentet eiciantur de ruinis suis. -
PS|109|11|Scrutetur fenerator omnem substantiam eius,et diripiant alieni labores eius.
PS|109|12|Non sit qui praebeat illi misericordiam,nec sit qui misereatur pupillis eius.
PS|109|13|Fiant nati eius in interitum,in generatione una deleatur nomen eorum.
PS|109|14|In memoriam redeat iniquitas patrum eius in conspectu Domini,et peccatum matris eius non deleatur.
PS|109|15|Fiant contra Dominum semper,et disperdat de terra memoriam eorum.
PS|109|16|Pro eo quod non est recordatus facere misericordiamet persecutus est hominem inopem et mendicumet compunctum corde, ut mortificaret.
PS|109|17|Et dilexit maledictionem: et veniat ei;et noluit benedictionem: et elongetur ab eo.
PS|109|18|Et induit maledictionem sicut vestimentum:et intret sicut aqua in interiora eius,et sicut oleum in ossa eius.
PS|109|19|Fiat ei sicut indumentum, quo operitur,et sicut zona, qua semper praecingitur.
PS|109|20|Haec retributio eorum, qui adversantur mihi apud Dominum,et qui loquuntur mala adversus animam meam.
PS|109|21|Et tu, Domine, Domine, fac mecum propter nomen tuum,quia suavis est misericordia tua;libera me,
PS|109|22|quia egenus et pauper ego sum,et cor meum vulneratum est intra me.
PS|109|23|Sicut umbra, cum declinat, pertransii,excussus sum sicut locustae.
PS|109|24|Genua mea infirmata sunt ieiunio,et caro mea contabuit absque oleo.
PS|109|25|Et ego factus sum opprobrium illis:viderunt me et moverunt capita sua.
PS|109|26|Adiuva me, Domine Deus meus,salvum me fac secundum misericordiam tuam.
PS|109|27|Et sciant quia manus tua haec:tu, Domine, hoc fecisti.
PS|109|28|Maledicant illi, et tu benedicas;qui insurgunt in me, confundantur,servus autem tuus laetabitur.
PS|109|29|Induantur, qui detrahunt mihi, pudoreet operiantur sicut diploide confusione sua.
PS|109|30|Confitebor Domino nimis in ore meoet in medio multorum laudabo eum,
PS|109|31|quia astitit a dextris pauperis,ut salvam faceret a iudicantibus animam eius.
PS|110|1|David. PSALMUS.Dixit Dominus Domino meo: " Sede a dextris meis,donec ponam inimicos tuos scabellum pedum tuorum ".
PS|110|2|Virgam potentiae tuae emittet Dominus ex Sion:dominare in medio inimicorum tuorum.
PS|110|3|Tecum principatus in die virtutis tuae,in splendoribus sanctis,ex utero ante luciferum genui te.
PS|110|4|Iuravit Dominus et non paenitebit eum: Tu es sacerdos in aeternum secundum ordinem Melchisedech ".
PS|110|5|Dominus a dextris tuis,conquassabit in die irae suae reges.
PS|110|6|Iudicabit in nationibus: cumulantur cadavera,conquassabit capita in terra spatiosa.
PS|110|7|De torrente in via bibet,propterea exaltabit caput.
PS|111|1|ALLELUIA.ALEPH. Confitebor Domino in toto corde meo,BETH. in consilio iustorum et congregatione.
PS|111|2|GHIMEL. Magna opera Domini,DALETH. exquirenda omnibus, qui cupiunt ea.
PS|111|3|HE. Decor et magnificentia opus eius,VAU. et iustitia eius manet in saeculum saeculi.
PS|111|4|ZAIN. Memoriam fecit mirabilium suorum,HETH. misericors et miserator Dominus.
PS|111|5|TETH. Escam dedit timentibus se;IOD. memor erit in saeculum testamenti sui.
PS|111|6|CAPH. Virtutem operum suorum annuntiavit populo suo,LAMED. ut det illis hereditatem gentium;
PS|111|7|MEM. opera manuum eius veritas et iudicium.NUN. Fidelia omnia mandata eius,
PS|111|8|SAMECH. confirmata in saeculum saeculi,AIN. facta in veritate et aequitate.
PS|111|9|PHE. Redemptionem misit populo suo,SADE. mandavit in aeternum testamentum suum.COPH. Sanctum et terribile nomen eius.
PS|111|10|RES. Initium sapientiae timor Domini,SIN. intellectus bonus omnibus facientibus ea;TAU. laudatio eius manet in saeculum saeculi.
PS|112|1|ALLELUIA.ALEPH. Beatus vir, qui timet Dominum,BETH. in mandatis eius cupit nimis.
PS|112|2|GHIMEL. Potens in terra erit semen eius,DALETH. generatio rectorum benedicetur.
PS|112|3|HE. Gloria et divitiae in domo eius,VAU. et iustitia eius manet in saeculum saeculi.
PS|112|4|ZAIN. Exortum est in tenebris lumen rectis,HETH. misericors et miserator et iustus.
PS|112|5|TETH. Iucundus homo, qui miseretur et commodat,IOD. disponet res suas in iudicio,
PS|112|6|CAPH. quia in aeternum non commovebitur.LAMED. In memoria aeterna erit iustus,
PS|112|7|MEM. ab auditione mala non timebit.NUN. Paratum cor eius, sperans in Domino,
PS|112|8|SAMECH. confirmatum est cor eius, non timebit,AIN. donec despiciat inimicos suos.
PS|112|9|PHE. Distribuit, dedit pauperibus;SADE. iustitia eius manet in saeculum saeculi,COPH. cornu eius exaltabitur in gloria.
PS|112|10|RES. Peccator videbit et irascetur,SIN. dentibus suis fremet et tabescet.TAU. Desiderium peccatorum peribit.
PS|113|1|ALLELUIA.Laudate, pueri Domini,laudate nomen Domini.
PS|113|2|Sit nomen Domini benedictumex hoc nunc et usque in saeculum.
PS|113|3|A solis ortu usque ad occasumlaudabile nomen Domini.
PS|113|4|Excelsus super omnes gentes Dominus,super caelos gloria eius.
PS|113|5|Quis sicut Dominus Deus noster,qui in altis habitat
PS|113|6|et se inclinat, ut respiciatin caelum et in terram?
PS|113|7|Suscitans de terra inopem,de stercore erigens pauperem,
PS|113|8|ut collocet eum cum principibus,cum principibus populi sui.
PS|113|9|Qui habitare facit sterilem in domo,matrem filiorum laetantem.
PS|114|1|ALLELUIA.In exitu Israel de Aegypto,domus Iacob de populo barbaro,
PS|114|2|factus est Iuda sanctuarium eius,Israel potestas eius.
PS|114|3|Mare vidit et fugit,Iordanis conversus est retrorsum;
PS|114|4|montes saltaverunt ut arietes,et colles sicut agni ovium. -
PS|114|5|Quid est tibi, mare, quod fugisti?Et tu, Iordanis, quia conversus es retrorsum?
PS|114|6|Montes, quod saltastis sicut arietes,et colles, sicut agni ovium?
PS|114|7|A facie Domini contremisce, terra,a facie Dei Iacob,
PS|114|8|qui convertit petram in stagna aquarumet silicem in fontes aquarum.
PS|115|1|Non nobis, Domine, non nobis,sed nomini tuo da gloriamsuper misericordia tua et veritate tua.
PS|115|2|Quare dicent gentes: Ubi est Deus eorum? ".
PS|115|3|Deus autem noster in caelo;omnia, quaecumque voluit, fecit.
PS|115|4|Simulacra gentium argentum et aurum,opera manuum hominum.
PS|115|5|Os habent et non loquentur,oculos habent et non videbunt.
PS|115|6|Aures habent et non audient,nares habent et non odorabunt.
PS|115|7|Manus habent et non palpabunt,pedes habent et non ambulabunt;non clamabunt in gutture suo.
PS|115|8|Similes illis erunt, qui faciunt ea,et omnes, qui confidunt in eis.
PS|115|9|Domus Israel speravit in Domino:adiutorium eorum et scutum eorum est.
PS|115|10|Domus Aaron speravit in Domino:adiutorium eorum et scutum eorum est.
PS|115|11|Qui timent Dominum, speraverunt in Domino:adiutorium eorum et scutum eorum est.
PS|115|12|Dominus memor fuit nostriet benedicet nobis:benedicet domui Israel,benedicet domui Aaron,
PS|115|13|benedicet omnibus, qui timent Dominum,pusillis cum maioribus.
PS|115|14|Adiciat Dominus super vos,super vos et super filios vestros.
PS|115|15|Benedicti vos a Domino,qui fecit caelum et terram.
PS|115|16|Caeli, caeli sunt Domino,terram autem dedit filiis hominum.
PS|115|17|Non mortui laudabunt te, Domine,neque omnes, qui descendunt in silentium,
PS|115|18|sed nos, qui vivimus, benedicimus Dominoex hoc nunc et usque in saeculum.
PS|116|1|ALLELUIA.Dilexi, quoniam exaudit Dominusvocem deprecationis meae.
PS|116|2|Quia inclinavit aurem suam mihi,cum in diebus meis invocabam.
PS|116|3|Circumdederunt me funes mortis,et angustiae inferni invenerunt me. Tribulationem et dolorem inveni
PS|116|4|et nomen Domini invocabam: O Domine, libera animam meam ".
PS|116|5|Misericors Dominus et iustus,et Deus noster miseretur.
PS|116|6|Custodiens parvulos Dominus;humiliatus sum, et salvum me faciet.
PS|116|7|Convertere, anima mea, in requiem tuam,quia Dominus benefecit tibi;
PS|116|8|quia eripuit animam meam de morte,oculos meos a lacrimis,pedes meos a lapsu.
PS|116|9|Ambulabo coram Dominoin regione vivorum. -
PS|116|10|Credidi, etiam cum locutus sum: " Ego humiliatus sum nimis ".
PS|116|11|Ego dixi in trepidatione mea: " Omnis homo mendax ".
PS|116|12|Quid retribuam Dominopro omnibus, quae retribuit mihi?
PS|116|13|Calicem salutaris accipiamet nomen Domini invocabo.
PS|116|14|Vota mea Domino reddamcoram omni populo eius.
PS|116|15|Pretiosa in conspectu Dominimors sanctorum eius.
PS|116|16|O Domine, ego servus tuus,ego servus tuus et filius ancillae tuae.Dirupisti vincula mea:
PS|116|17|tibi sacrificabo hostiam laudiset nomen Domini invocabo.
PS|116|18|Vota mea Domino reddamcoram omni populo eius
PS|116|19|in atriis domus Domini,in medio tui, Ierusalem.
PS|117|1|ALLELUIA.Laudate Dominum, omnes gentes;collaudate eum, omnes populi.
PS|117|2|Quoniam confirmata est super nos misericordia eius,et veritas Domini manet in aeternum.
PS|118|1|ALLELUIA.Confitemini Domino, quoniam bonus,quoniam in saeculum misericordia eius.
PS|118|2|Dicat nunc Israel, quoniam bonus,quoniam in saeculum misericordia eius.
PS|118|3|Dicat nunc domus Aaron,quoniam in saeculum misericordia eius.
PS|118|4|Dicant nunc, qui timent Dominum,quoniam in saeculum misericordia eius.
PS|118|5|De tribulatione invocavi Dominum,et exaudivit me educens in latitudinem Dominus.
PS|118|6|Dominus mecum,non timebo, quid faciat mihi homo.
PS|118|7|Dominus mecum adiutor meus,et ego despiciam inimicos meos.
PS|118|8|Bonum est confugere ad Dominumquam confidere in homine.
PS|118|9|Bonum est confugere ad Dominumquam confidere in principibus.
PS|118|10|Omnes gentes circuierunt me,et in nomine Domini excidi eos.
PS|118|11|Circumdantes circumdederunt me,et in nomine Domini excidi eos.
PS|118|12|Circumdederunt me sicut apeset exarserunt sicut ignis in spinis,et in nomine Domini excidi eos.
PS|118|13|Impellentes impulerunt me, ut caderem,et Dominus adiuvit me.
PS|118|14|Fortitudo mea et laus mea Dominuset factus est mihi in salutem.
PS|118|15|Vox iubilationis et salutisin tabernaculis iustorum: Dextera Domini fecit virtutem!
PS|118|16|Dextera Domini exaltata est;dextera Domini fecit virtutem! ".
PS|118|17|Non moriar, sed vivamet narrabo opera Domini.
PS|118|18|Castigans castigavit me Dominuset morti non tradidit me.
PS|118|19|Aperite mihi portas iustitiae;ingressus in eas confitebor Domino.
PS|118|20|Haec porta Domini;iusti intrabunt in eam. -
PS|118|21|Confitebor tibi, quoniam exaudisti meet factus es mihi in salutem.
PS|118|22|Lapidem quem reprobaverunt aedificantes,hic factus est in caput anguli;
PS|118|23|a Domino factum est istudet est mirabile in oculis nostris.
PS|118|24|Haec est dies, quam fecit Dominus:exsultemus et laetemur in ea.
PS|118|25|O Domine, salvum me fac;o Domine, da prosperitatem!
PS|118|26|Benedictus, qui venit in nomine Domini.Benedicimus vobis de domo Domini.
PS|118|27|Deus Dominus et illuxit nobis.Instruite sollemnitatem in ramis condensisusque ad cornua altaris.
PS|118|28|Deus meus es tu, et confitebor tibi,Deus meus, et exaltabo te.
PS|118|29|Confitemini Domino, quoniam bonus,quoniam in saeculum misericordia eius.
PS|119|1|ALLELUIA.ALEPH. Beati immaculati in via,qui ambulant in lege Domini.
PS|119|2|Beati, qui servant testimonia eius,in toto corde exquirunt eum.
PS|119|3|Non enim operati sunt iniquitatem,in viis eius ambulaverunt.
PS|119|4|Tu mandastimandata tua custodiri nimis.
PS|119|5|Utinam dirigantur viae meaead custodiendas iustificationes tuas!
PS|119|6|Tunc non confundar,cum perspexero in omnibus praeceptis tuis.
PS|119|7|Confitebor tibi in directione cordis,in eo quod didici iudicia iustitiae tuae.
PS|119|8|Iustificationes tuas custodiam,non me derelinquas usquequaque.
PS|119|9|BETH. In quo mundabit adulescentior viam suam?In custodiendo sermones tuos.
PS|119|10|In toto corde meo exquisivi te;ne errare me facias a praeceptis tuis.
PS|119|11|In corde meo abscondi eloquia tua,ut non peccem tibi.
PS|119|12|Benedictus es, Domine;doce me iustificationes tuas.
PS|119|13|In labiis meisnumeravi omnia iudicia oris tui.
PS|119|14|In via testimoniorum tuorum delectatus sumsicut in omnibus divitiis.
PS|119|15|In mandatis tuis exerceboret considerabo vias tuas.
PS|119|16|In iustificationibus tuis delectabor,non obliviscar sermonem tuum.
PS|119|17|GHIMEL. Benefac servo tuo, et vivamet custodiam sermonem tuum.
PS|119|18|Revela oculos meos,et considerabo mirabilia de lege tua.
PS|119|19|Incola ego sum in terra,non abscondas a me praecepta tua.
PS|119|20|Defecit anima mea in desiderando iudicia tuain omni tempore.
PS|119|21|Increpasti superbos;maledicti, qui errant a praeceptis tuis.
PS|119|22|Aufer a me opprobrium et contemptum,quia testimonia tua servavi.
PS|119|23|Etsi principes sedent et adversum me loquuntur,servus tamen tuus exercetur in iustificationibus tuis.
PS|119|24|Nam et testimonia tua delectatio mea,et consilium meum iustificationes tuae.
PS|119|25|DALETH. Adhaesit pulveri anima mea;vivifica me secundum verbum tuum.
PS|119|26|Vias meas enuntiavi, et exaudisti me;doce me iustificationes tuas.
PS|119|27|Viam mandatorum tuorum fac me intellegere,et exercebor in mirabilibus tuis.
PS|119|28|Lacrimata est anima mea prae maerore;erige me secundum verbum tuum.
PS|119|29|Viam mendacii averte a meet legem tuam da mihi benigne.
PS|119|30|Viam veritatis elegi,iudicia tua proposui mihi.
PS|119|31|Adhaesi testimoniis tuis, Domine;noli me confundere.
PS|119|32|Viam mandatorum tuorum curram,quia dilatasti cor meum.
PS|119|33|HE. Legem pone mihi, Domine, viam iustificationum tuarum,et servabo eam semper.
PS|119|34|Da mihi intellectum, et servabo legem tuamet custodiam illam in toto corde meo.
PS|119|35|Deduc me in semitam praeceptorum tuorum,quia ipsam volui.
PS|119|36|Inclina cor meum in testimonia tuaet non in avaritiam.
PS|119|37|Averte oculos meos, ne videant vanitatem;in via tua vivifica me.
PS|119|38|Suscita servo tuo eloquium tuum,quod est ad timorem tuum.
PS|119|39|Amove opprobrium meum, quod suspicatus sum,quia iudicia tua iucunda.
PS|119|40|Ecce concupivi mandata tua;in iustitia tua vivifica me.
PS|119|41|VAU. Et veniat super me misericordia tua, Domine,salutare tuum secundum eloquium tuum.
PS|119|42|Et respondebo exprobrantibus mihi verbum,quia speravi in sermonibus tuis.
PS|119|43|Et ne auferas de ore meo verbum veritatis usquequaque,quia in iudiciis tuis supersperavi.
PS|119|44|Et custodiam legem tuam semper,in saeculum et in saeculum saeculi.
PS|119|45|Et ambulabo in latitudine,quia mandata tua exquisivi.
PS|119|46|Et loquar de testimoniis tuis in conspectu regumet non confundar.
PS|119|47|Et delectabor in praeceptis tuis,quae dilexi.
PS|119|48|Et levabo manus meas ad praecepta tua, quae dilexi;et exercebor in iustificationibus tuis. -
PS|119|49|ZAIN. Memor esto verbi tui servo tuo,in quo mihi spem dedisti.
PS|119|50|Hoc me consolatum est in humiliatione mea,quia eloquium tuum vivificavit me.
PS|119|51|Superbi deriserunt me vehementer;a lege autem tua non declinavi.
PS|119|52|Memor fui iudiciorum tuorum a saeculo, Domine,et consolatus sum.
PS|119|53|Indignatio tenuit mepropter peccatores derelinquentes legem tuam.
PS|119|54|Cantica factae sunt mihi iustificationes tuaein loco peregrinationis meae.
PS|119|55|Memor fui nocte nominis tui, Domine,et custodiam legem tuam.
PS|119|56|Hoc factum est mihi,quia mandata tua servavi.
PS|119|57|HETH. Portio mea Dominus:dixi custodire verba tua.
PS|119|58|Deprecatus sum faciem tuam in toto corde meo;miserere mei secundum eloquium tuum.
PS|119|59|Cogitavi vias measet converti pedes meos in testimonia tua.
PS|119|60|Festinavi et non sum moratus,ut custodiam praecepta tua.
PS|119|61|Funes peccatorum circumplexi sunt me,et legem tuam non sum oblitus.
PS|119|62|Media nocte surgebam ad confitendum tibisuper iudicia iustitiae tuae.
PS|119|63|Particeps ego sum omnium timentium teet custodientium mandata tua.
PS|119|64|Misericordia tua, Domine, plena est terra;iustificationes tuas doce me.
PS|119|65|TETH. Bonitatem fecisti cum servo tuo, Domine,secundum verbum tuum.
PS|119|66|Bonitatem et prudentiam et scientiam doce me,quia praeceptis tuis credidi.
PS|119|67|Priusquam humiliarer ego erravi;nunc autem eloquium tuum custodiam.
PS|119|68|Bonus es tu et benefaciens,doce me iustificationes tuas.
PS|119|69|Excogitaverunt contra me dolosa superbi,ego autem in toto corde meo servabo mandata tua.
PS|119|70|Incrassatum est sicut adeps cor eorum,ego vero in lege tua delectatus sum.
PS|119|71|Bonum mihi quia humiliatus sum,ut discam iustificationes tuas.
PS|119|72|Bonum mihi lex oris tuisuper milia auri et argenti.
PS|119|73|IOD. Manus tuae fecerunt me et plasmaverunt me;da mihi intellectum, et discam praecepta tua.
PS|119|74|Qui timent te, videbunt me et laetabuntur,quia in verba tua supersperavi.
PS|119|75|Cognovi, Domine, quia aequitas iudicia tua,et in veritate humiliasti me.
PS|119|76|Fiat misericordia tua, ut consoletur me,secundum eloquium tuum servo tuo.
PS|119|77|Veniant mihi miserationes tuae, et vivam,quia lex tua delectatio mea est.
PS|119|78|Confundantur superbi, quoniam dolose incurvaverunt me,ego autem exercebor in mandatis tuis.
PS|119|79|Convertantur mihi timentes te,et qui noverunt testimonia tua.
PS|119|80|Fiat cor meum immaculatum in iustificationibus tuis,ut non confundar.
PS|119|81|CAPH. Defecit in salutare tuum anima mea,et in verbum tuum supersperavi.
PS|119|82|Defecerunt oculi mei in eloquium tuum,dicentes: " Quando consolaberis me? ".
PS|119|83|Quia factus sum sicut uter in fumo;iustificationes tuas non sum oblitus.
PS|119|84|Quot sunt dies servi tui?Quando facies de persequentibus me iudicium?
PS|119|85|Foderunt mihi foveas superbi,qui non sunt secundum legem tuam.
PS|119|86|Omnia praecepta tua veritas;dolose persecuti sunt me; adiuva me.
PS|119|87|Paulo minus consummaverunt me in terra,ego autem non dereliqui mandata tua.
PS|119|88|Secundum misericordiam tuam vivifica me,et custodiam testimonia oris tui. -
PS|119|89|LAMED. In aeternum, Domine,verbum tuum constitutum est in caelo.
PS|119|90|In generationem et generationem veritas tua;firmasti terram, et permanet.
PS|119|91|Secundum iudicia tua permanent hodie,quoniam omnia serviunt tibi.
PS|119|92|Nisi quod lex tua delectatio mea est,tunc forte periissem in humilia tione mea.
PS|119|93|In aeternum non obliviscar man data tua,quia in ipsis vivificasti me.
PS|119|94|Tuus sum ego: salvum me fac,quoniam mandata tua exqui sivi.
PS|119|95|Me exspectaverunt peccatores, ut perderent me;testimonia tua intellexi.
PS|119|96|Omni consummationi vidi finem,latum praeceptum tuum nimis.
PS|119|97|MEM. Quomodo dilexi legem tuam, Domine;tota die meditatio mea est.
PS|119|98|Super inimicos meos sapientem me fecit praeceptum tuum,quia in aeternum mihi est.
PS|119|99|Super omnes docentes me prudens factus sum,quia testimonia tua meditatio mea est.
PS|119|100|Super senes intellexi,quia mandata tua servavi.
PS|119|101|Ab omni via mala prohibui pedes meos,ut custodiam verba tua.
PS|119|102|A iudiciis tuis non declinavi,quia tu legem posuisti mihi.
PS|119|103|Quam dulcia faucibus meis eloquia tua,super mel ori meo.
PS|119|104|A mandatis tuis intellexi;propterea odivi omnem viam mendacii.
PS|119|105|NUN. Lucerna pedibus meis verbum tuumet lumen semitis meis.
PS|119|106|Iuravi et statuicustodire iudicia iustitiae tuae.
PS|119|107|Humiliatus sum usquequaque, Domine;vivifica me secundum verbum tuum.
PS|119|108|Voluntaria oris mei beneplacita sint, Domine,et iudicia tua doce me.
PS|119|109|Anima mea in manibus meis semper,et legem tuam non sum oblitus.
PS|119|110|Posuerunt peccatores laqueum mihi,et de mandatis tuis non erravi.
PS|119|111|Hereditas mea testimonia tua in aeternum,quia exsultatio cordis mei sunt.
PS|119|112|Inclinavi cor meum ad faciendas iustificationes tuasin aeternum, in finem.
PS|119|113|SAMECH. Duplices corde odio habuiet legem tuam dilexi.
PS|119|114|Tegmen et scutum meum es tu,et in verbum tuum supersperavi.
PS|119|115|Declinate a me, maligni,et servabo praecepta Dei mei.
PS|119|116|Suscipe me secundum eloquium tuum, et vivam;et non confundas me ab exspectatione mea.
PS|119|117|Sustenta me, et salvus eroet delectabor in iustificationibus tuis semper.
PS|119|118|Sprevisti omnes discedentes a iustificationibus tuis,quia mendacium cogitatio eorum.
PS|119|119|Quasi scoriam delesti omnes peccatores terrae;ideo dilexi testimonia tua.
PS|119|120|Horruit a timore tuo caro mea;a iudiciis enim tuis timui.
PS|119|121|AIN. Feci iudicium et iustitiam;non tradas me calumniantibus me.
PS|119|122|Sponde pro servo tuo in bonum;non calumnientur me superbi.
PS|119|123|Oculi mei defecerunt in desiderio salutaris tuiet eloquii iustitiae tuae.
PS|119|124|Fac cum servo tuo secundum misericordiam tuamet iustificationes tuas doce me.
PS|119|125|Servus tuus sum ego;da mihi intellectum, ut sciam testimonia tua.
PS|119|126|Tempus faciendi Domino;dissipaverunt legem tuam.
PS|119|127|Ideo dilexi praecepta tuasuper aurum et obryzum.
PS|119|128|Propterea ad omnia mandata tua dirigebar,omnem viam mendacii odio habui. -
PS|119|129|PHE. Mirabilia testimonia tua,ideo servavit ea anima mea.
PS|119|130|Declaratio sermonum tuorum illuminatet intellectum dat parvulis.
PS|119|131|Os meum aperui et attraxi spiritum,quia praecepta tua desiderabam.
PS|119|132|Convertere in me et miserere meisecundum iudicium tuum cum diligentibus nomen tuum.
PS|119|133|Gressus meos dirige secundum eloquium tuum,et non dominetur mei omnis iniquitas.
PS|119|134|Redime me a calumniis hominum,ut custodiam mandata tua.
PS|119|135|Faciem tuam illumina super servum tuumet doce me iustificationes tuas.
PS|119|136|Rivulos aquarum deduxerunt oculi mei,quia non custodierunt legem tuam.
PS|119|137|SADE. Iustus es, Domine,et rectum iudicium tuum.
PS|119|138|Mandasti in iustitia testimonia tuaet in veritate nimis.
PS|119|139|Consumpsit me zelus meus,quia obliti sunt verba tua inimici mei.
PS|119|140|Ignitum eloquium tuum vehementer,et servus tuus dilexit illud.
PS|119|141|Adulescentulus sum ego et contemptus;mandata tua non sum oblitus.
PS|119|142|Iustitia tua iustitia in aeternum,et lex tua veritas.
PS|119|143|Tribulatio et angustia invenerunt me;praecepta tua delectatio mea est.
PS|119|144|Iustitia testimonia tua in aeternum;intellectum da mihi, et vivam.
PS|119|145|COPH. Clamavi in toto corde, exaudi me, Domine;iustificationes tuas servabo.
PS|119|146|Clamavi ad te, salvum me fac,ut custodiam testimonia tua.
PS|119|147|Praeveni diluculo et clamavi,in verba tua supersperavi.
PS|119|148|Praevenerunt oculi mei vigilias,ut meditarer eloquia tua.
PS|119|149|Vocem meam audi secundum misericordiam tuam, Domine,secundum iudicium tuum vivifica me.
PS|119|150|Appropinquaverunt persequentes me in malitia,a lege autem tua longe facti sunt.
PS|119|151|Prope es tu, Domine,et omnia praecepta tua veritas.
PS|119|152|Ab initio cognovi de testimoniis tuis,quia in aeternum fundasti ea.
PS|119|153|RES. Vide humiliationem meam et eripe me,quia legem tuam non sum oblitus.
PS|119|154|Iudica causam meam et redime me;propter eloquium tuum vivifica me.
PS|119|155|Longe a peccatoribus salus,quia iustificationes tuas non exquisierunt.
PS|119|156|Misericordiae tuae multae, Domine;secundum iudicia tua vivifica me.
PS|119|157|Multi, qui persequuntur me et tribulant me;a testimoniis tuis non declinavi.
PS|119|158|Vidi praevaricantes, et taeduit me,quia eloquia tua non custodierunt.
PS|119|159|Vide quoniam mandata tua dilexi, Domine;secundum misericordiam tuam vivifica me.
PS|119|160|Principium verborum tuorum veritas,in aeternum omnia iudicia iustitiae tuae.
PS|119|161|SIN. Principes persecuti sunt me gratis,et a verbis tuis formidavit cor meum.
PS|119|162|Laetabor ego super eloquia tua,sicut qui invenit spolia multa.
PS|119|163|Mendacium odio habui et abominatus sum;legem autem tuam dilexi.
PS|119|164|Septies in die laudem dixi tibisuper iudicia iustitiae tuae.
PS|119|165|Pax multa diligentibus legem tuam, et non est illis scandalum.
PS|119|166|Exspectabam salutare tuum, Domine,et praecepta tua feci.
PS|119|167|Custodivit anima mea testimonia tua,et dilexi ea vehementer.
PS|119|168|Servavi mandata tua et testimonia tua,quia omnes viae meae in conspectu tuo.
PS|119|169|TAU. Appropinquet deprecatio mea in conspectu tuo, Domine;iuxta verbum tuum da mihi intellectum.
PS|119|170|Intret postulatio mea in conspectu tuo;secundum eloquium tuum libera me.
PS|119|171|Eructabunt labia mea hymnum,cum docueris me iustificationes tuas.
PS|119|172|Cantet lingua mea eloquium tuum,quia omnia praecepta tua iustitia.
PS|119|173|Fiat manus tua, ut adiuvet me,quoniam mandata tua elegi.
PS|119|174|Concupivi salutare tuum, Domine,et lex tua delectatio mea est.
PS|119|175|Vivet anima mea et laudabit te,et iudicia tua adiuvabunt me.
PS|119|176|Erravi sicut ovis, quae periit;quaere servum tuum, quia praecepta tua non sum oblitus.
PS|120|1|Canticum ascensionum.Ad Dominum, cum tribularer, clamavi,et exaudivit me.
PS|120|2|Domine, libera animam meam a labiis mendacii,a lingua dolosa.
PS|120|3|Quid detur tibi aut quid apponatur tibi,lingua dolosa?
PS|120|4|Sagittae potentis acutaecum carbonibus iuniperorum.
PS|120|5|Heu mihi, quia peregrinatus sum in Mosoch,habitavi ad tabernacula Cedar!
PS|120|6|Multum incola fuit anima meacum his, qui oderunt pacem.
PS|120|7|Ego eram pacificus;cum loquebar, illi impugnabant me.
PS|121|1|Canticum ascensionum.Levabo oculos meos in montes:unde veniet auxilium mihi?
PS|121|2|Auxilium meum a Domino,qui fecit caelum et terram.
PS|121|3|Non dabit in commotionem pedem tuumneque dormitabit, qui custodit te.
PS|121|4|Ecce non dormitabit neque dormiet,qui custodit Israel.
PS|121|5|Dominus custodit te,Dominus umbraculum tuumad manum dexteram tuam.
PS|121|6|Per diem sol non percutiet te,neque luna per noctem.
PS|121|7|Dominus custodiet te ab omni malo;custodiet animam tuam Dominus.
PS|121|8|Dominus custodiet introitum tuum et exitum tuumex hoc nunc et usque in saeculum.
PS|122|1|Canticum ascensionum. David.Laetatus sum in eo, quod dixerunt mihi: In domum Domini ibimus ".
PS|122|2|Stantes iam sunt pedes nostriin portis tuis, Ierusalem.
PS|122|3|Ierusalem, quae aedificata est ut civitas,sibi compacta in idipsum.
PS|122|4|Illuc enim ascenderunt tribus, tribus Domini,testimonium Israel, ad confitendum nomini Domini.
PS|122|5|Quia illic sederunt sedes ad iudicium,sedes domus David.
PS|122|6|Rogate, quae ad pacem sunt Ierusalem: Securi sint diligentes te!
PS|122|7|Fiat pax in muris tuis,et securitas in turribus tuis! ".
PS|122|8|Propter fratres meos et proximos meosloquar: " Pax in te! ".
PS|122|9|Propter domum Domini Dei nostriexquiram bona tibi.
PS|123|1|Canticum ascensionum.Ad te levavi oculos meos,qui habitas in caelis.
PS|123|2|Ecce sicut oculi servorum ad manus dominorum suorum,sicut oculi ancillae ad manus dominae suae,ita oculi nostri ad Dominum Deum nostrum,donec misereatur nostri.
PS|123|3|Miserere nostri, Domine, miserere nostri,quia multum repleti sumus despectione;
PS|123|4|quia multum repleta est anima nostraderisione abundantium et despectione superborum.
PS|124|1|Canticum ascensionum. David.Nisi quia Dominus erat in nobis,dicat nunc Israel,
PS|124|2|nisi quia Dominus erat in nobis,cum exsurgerent homines in nos:
PS|124|3|forte vivos deglutissent nos,cum irasceretur furor eorum in nos.
PS|124|4|Forsitan aqua absorbuisset nos,torrens pertransisset animam nostram;
PS|124|5|forsitan pertransissent animam nostramaquae intumescentes.
PS|124|6|Benedictus Dominus,qui non dedit nos in direptionem dentibus eorum.
PS|124|7|Anima nostra sicut passer erepta estde laqueo venantium:laqueus contritus est,et nos erepti sumus.
PS|124|8|Adiutorium nostrum in nomine Domini,qui fecit caelum et terram.
PS|125|1|Canticum ascensionum.Qui confidunt in Domino, sicut mons Sion:non commovebitur, in aeternum manet.
PS|125|2|Ierusalem, montes in circuitu eius,et Dominus in circuitu populi suiex hoc nunc et usque in saeculum.
PS|125|3|Quia non requiescet virga iniquitatis super sortem iustorum,ut non extendant iusti ad iniquitatem manus suas.
PS|125|4|Benefac, Domine, boniset rectis corde.
PS|125|5|Declinantes autem per vias pravasadducet Dominus cum operantibus iniquitatem.Pax super Israel!
PS|126|1|Canticum ascensionum.In convertendo Dominus captivitatem Sion,facti sumus quasi somniantes.
PS|126|2|Tunc repletum est gaudio os nostrum,et lingua nostra exsultatione.Tunc dicebant inter gentes: Magnificavit Dominus facere cum eis ".
PS|126|3|Magnificavit Dominus facere nobiscum;facti sumus laetantes.
PS|126|4|Converte, Domine, captivitatem nostram,sicut torrentes in austro.
PS|126|5|Qui seminant in lacrimis,in exsultatione metent.
PS|126|6|Euntes ibant et flebantsemen spargendum portantes;venientes autem venient in exsultationeportantes manipulos suos.
PS|127|1|Canticum ascensionum. Salomonis.Nisi Dominus aedificaverit domum,in vanum laborant, qui aedificant eam.Nisi Dominus custodierit civitatem,frustra vigilat, qui custodit eam.
PS|127|2|Vanum est vobis ante lucem surgere et sero quiescere,qui manducatis panem laboris,quia dabit dilectis suis somnum.
PS|127|3|Ecce hereditas Domini filii,merces fructus ventris.
PS|127|4|Sicut sagittae in manu potentis,ita filii iuventutis.
PS|127|5|Beatus vir, qui implevit pharetram suam ex ipsis:non confundetur, cum loquetur inimicis suis in porta.
PS|128|1|Canticum ascensionum.Beatus omnis, qui timet Dominum,qui ambulat in viis eius.
PS|128|2|Labores manuum tuarum manducabis,beatus es, et bene tibi erit.
PS|128|3|Uxor tua sicut vitis fructiferain lateribus domus tuae;filii tui sicut novellae olivarumin circuitu mensae tuae.
PS|128|4|Ecce sic benedicetur homo,qui timet Dominum.
PS|128|5|Benedicat tibi Dominus ex Sion,et videas bona Ierusalemomnibus diebus vitae tuae;
PS|128|6|et videas filios filiorum tuorum.Pax super Israel!
PS|129|1|Canticum ascensionum.Saepe expugnaverunt me a iuventute mea,dicat nunc Israel,
PS|129|2|saepe expugnaverunt me a iuventute mea,etenim non potuerunt adversum me.
PS|129|3|Supra dorsum meum araverunt aratores,prolongaverunt sulcos suos.
PS|129|4|Dominus autem iustusconcidit cervices peccatorum.
PS|129|5|Confundantur et convertantur retrorsumomnes, qui oderunt Sion.
PS|129|6|Fiant sicut fenum tectorum,quod, priusquam evellatur, exaruit;
PS|129|7|de quo non implevit manum suam, qui metit,et sinum suum, qui manipulos colligit.
PS|129|8|Et non dixerunt, qui praeteribant: Benedictio Domini super vos,benedicimus vobis in nomine Domini ".
PS|130|1|Canticum ascensionum.De profundis clamavi ad te, Domine;
PS|130|2|Domine, exaudi vocem meam.Fiant aures tuae intendentesin vocem deprecationis meae.
PS|130|3|Si iniquitates observaveris, Domine,Domine, quis sustinebit?
PS|130|4|Quia apud te propitiatio est,ut timeamus te.
PS|130|5|Sustinui te, Domine,sustinuit anima mea in verbo eius;speravit
PS|130|6|anima mea in Dominomagis quam custodes auroram.Magis quam custodes auroram
PS|130|7|speret Israel in Domino,quia apud Dominum misericordia,et copiosa apud eum redemptio.
PS|130|8|Et ipse redimet Israelex omnibus iniquitatibus eius.
PS|131|1|Canticum ascensionum. David.Domine, non est exaltatum cor meum,neque elati sunt oculi mei,neque ambulavi in magnisneque in mirabilibus super me.
PS|131|2|Vere pacatam et quietamfeci animam meam;sicut ablactatus in sinu matris suae,sicut ablactatus, ita in me est anima mea.
PS|131|3|Speret Israel in Dominoex hoc nunc et usque in saeculum.
PS|132|1|Canticum ascensionum.Memento, Domine, Davidet omnis mansuetudinis eius,
PS|132|2|quia iuravit Domino,votum vovit Potenti Iacob:
PS|132|3|" Non introibo in tabernaculum domus meae,non ascendam in lectum strati mei,
PS|132|4|non dabo somnum oculis meiset palpebris meis dormitationem,
PS|132|5|donec inveniam locum Domino,tabernaculum Potenti Iacob ".
PS|132|6|Ecce audivimus eam esse in Ephratha,invenimus eam in campis Iaar.
PS|132|7|Ingrediamur in tabernaculum eius,adoremus ad scabellum pedum eius. -
PS|132|8|Surge, Domine, in requiem tuam,tu et arca fortitudinis tuae.
PS|132|9|Sacerdotes tui induantur iustitiam,et sancti tui exsultent.
PS|132|10|Propter David servum tuumnon avertas faciem christi tui.
PS|132|11|Iuravit Dominus David veritatemet non recedet ab ea: De fructu ventris tuiponam super sedem tuam.
PS|132|12|Si custodierint filii tui testamentum meumet testimonia mea, quae docebo eos,filii eorum usque in saeculumsedebunt super sedem tuam ".
PS|132|13|Quoniam elegit Dominus Sion,desideravit eam in habitationem sibi:
PS|132|14|" Haec requies mea in saeculum saeculi;hic habitabo, quoniam desideravi eam.
PS|132|15|Cibaria eius benedicens benedicam,pauperes eius saturabo panibus.
PS|132|16|Sacerdotes eius induam salutari,et sancti eius exsultatione exsultabunt.
PS|132|17|Illic germinare faciam cornu David,parabo lucernam christo meo.
PS|132|18|Inimicos eius induam confusione,super ipsum autem efflorebit diadema eius ".
PS|133|1|Canticum ascensionum. David.Ecce quam bonum et quam iucundumhabitare fratres in unum:
PS|133|2|sicut unguentum optimum in capite,quod descendit in barbam, barbam Aaron,quod descendit in oram vestimenti eius;
PS|133|3|sicut ros Hermon, qui descendit in montes Sion,quoniam illic mandavit Dominus benedictionem,vitam usque in saeculum.
PS|134|1|Canticum ascensionum.Ecce benedicite Dominum,omnes servi Domini,qui statis in domo Domini per noctes.
PS|134|2|Extollite manus vestras ad sanctuariumet benedicite Dominum.
PS|134|3|Benedicat te Dominus ex Sion,qui fecit caelum et terram.
PS|135|1|ALLELUIA.Laudate nomen Domini,laudate, servi Domini,
PS|135|2|qui statis in domo Domini,in atriis domus Dei nostri.
PS|135|3|Laudate Dominum, quia bonus Dominus;psallite nomini eius, quoniam suave.
PS|135|4|Quoniam Iacob elegit sibi Dominus,Israel in peculium sibi.
PS|135|5|Quia ego cognovi quod magnus est Dominus,et Deus noster prae omnibus diis.
PS|135|6|Omnia, quaecumque voluit,Dominus fecit in caelo et in terra,in mari et in omnibus abyssis.
PS|135|7|Adducens nubes ab extremo terrae,fulgura in pluviam facit,producit ventos de thesauris suis.
PS|135|8|Qui percussit primogenita Aegyptiab homine usque ad pecus.
PS|135|9|Misit signa et prodigia in medio tui, Aegypte,in pharaonem et in omnes servos eius.
PS|135|10|Qui percussit gentes multaset occidit reges fortes:
PS|135|11|Sehon regem Amorraeorumet Og regem Basanet omnia regna Chanaan.
PS|135|12|Et dedit terram eorum hereditatem,hereditatem Israel populo suo.
PS|135|13|Domine, nomen tuum in aeternum;Domine, memoriale tuum in generationem et generationem.
PS|135|14|Quia iudicabit Dominus populum suumet servorum suorum miserebitur.
PS|135|15|Simulacra gentium argentum et aurum,opera manuum hominum.
PS|135|16|Os habent et non loquentur,oculos habent et non videbunt.
PS|135|17|Aures habent et non audient;neque enim est spiritus in ore ipsorum.
PS|135|18|Similes illis erunt, qui faciunt ea,et omnes, qui confidunt in eis.
PS|135|19|Domus Israel, benedicite Domino;domus Aaron, benedicite Domino;
PS|135|20|domus Levi, benedicite Domino;qui timetis Dominum, benedicite Domino.
PS|135|21|Benedictus Dominus ex Sion,qui habitat in Ierusalem. ALLELUIA.
PS|136|1|ALLELUIA.Confitemini Domino, quoniam bonus,quoniam in aeternum misericordia eius.
PS|136|2|Confitemini Deo deorum,quoniam in aeternum misericordia eius.
PS|136|3|Confitemini Domino dominorum,quoniam in aeternum misericordia eius.
PS|136|4|Qui facit mirabilia magna solus,quoniam in aeternum misericordia eius.
PS|136|5|Qui fecit caelos in intellectu,quoniam in aeternum misericordia eius.
PS|136|6|Qui expandit terram super aquas,quoniam in aeternum misericordia eius.
PS|136|7|Qui fecit luminaria magna,quoniam in aeternum misericordia eius:
PS|136|8|solem, ut praeesset diei,quoniam in aeternum misericordia eius;
PS|136|9|lunam et stellas, ut praeessent nocti, quoniam in aeternum misericordia eius.
PS|136|10|Qui percussit Aegyptum in primogenitis eorum,quoniam in aeternum misericordia eius.
PS|136|11|Qui eduxit Israel de medio eorum,quoniam in aeternum misericordia eius,
PS|136|12|in manu potenti et brachio extento,quoniam in aeternum misericordia eius.
PS|136|13|Qui divisit mare Rubrum in divisiones,quoniam in aeternum misericordia eius.
PS|136|14|Et traduxit Israel per medium eius,quoniam in aeternum misericordia eius.
PS|136|15|Et excussit pharaonem et virtutem eius in mari Rubro,quoniam in aeternum misericordia eius.
PS|136|16|Qui traduxit populum suum per desertum,quoniam in aeternum misericordia eius.
PS|136|17|Qui percussit reges magnos,quoniam in aeternum misericordia eius;
PS|136|18|et occidit reges potentes,quoniam in aeternum misericordia eius:
PS|136|19|Sehon regem Amorraeorum,quoniam in aeternum misericordia eius;
PS|136|20|et Og regem Basan,quoniam in aeternum misericordia eius.
PS|136|21|Et dedit terram eorum hereditatem,quoniam in aeternum misericordia eius,
PS|136|22|hereditatem Israel servo suo,quoniam in aeternum misericordia eius.
PS|136|23|Qui in humilitate nostra memor fuit nostri,quoniam in aeternum misericordia eius;
PS|136|24|et redemit nos ab inimicis nostris,quoniam in aeternum misericordia eius.
PS|136|25|Qui dat escam omni carni,quoniam ìn aeternum misericordia eius.
PS|136|26|Confitemini Deo caeli,quoniam in aeternum misericordia eius.
PS|137|1|Super flumina Babylonis,illic sedimus et flevimus,cum recordaremur Sion.
PS|137|2|In salicibus in medio eiussuspendimus citharas nostras.
PS|137|3|Quia illic rogaverunt nos,qui captivos duxerunt nos,verba cantionum,et, qui affligebant nos, laetitiam: Cantate nobis de canticis Sion ".
PS|137|4|Quomodo cantabimus canticum Dominiin terra aliena?
PS|137|5|Si oblitus fuero tui, Ierusalem,oblivioni detur dextera mea;
PS|137|6|adhaereat lingua mea faucibus meis,si non meminero tui,si non praeposuero Ierusalemin capite laetitiae meae.
PS|137|7|Memor esto, Domine, adversus filios Edomdiei Ierusalem;qui dicebant: " Exinanite, exinaniteusque ad fundamentum in ea ".
PS|137|8|Filia Babylonis devastans,beatus, qui retribuet tibi retributionem tuam,quam retribuisti nobis;
PS|137|9|beatus, qui tenebitet allidet parvulos tuos ad petram.
PS|138|1|David.Confitebor tibi, Domine, in toto corde meo,quoniam audisti verba oris mei.In conspectu angelorum psallam tibi,
PS|138|2|adorabo ad templum sanctum tuum;et confitebor nomini tuopropter misericordiam tuam et veritatem tuam,quoniam magnificasti super omne nomen eloquium tuum.
PS|138|3|In quacumque die invocavero te, exaudi me;multiplicabis in anima mea virtutem.
PS|138|4|Confitebuntur tibi, Domine, omnes reges terrae,quia audierunt eloquia oris tui.
PS|138|5|Et cantabunt vias Domini,quoniam magna est gloria Domini;
PS|138|6|quoniam excelsus Dominus et humilem respicitet superbum a longe cognoscit.
PS|138|7|Si ambulavero in medio tribulationis, vivificabis me;et contra iram inimicorum meorum extendes manum tuam,et salvum me faciet dextera tua.
PS|138|8|Dominus perficiet pro me;Domine, misericordia tua in saeculum:opera manuum tuarum ne despicias.
PS|139|1|Magistro chori. David. PSALMUS.Domine, scrutatus es et cognovisti me,
PS|139|2|tu cognovisti sessionem meam et resurrectionem meam.Intellexisti cogitationes meas de longe,
PS|139|3|semitam meam et accubitum meum investigasti.Et omnes vias meas perspexisti,
PS|139|4|quia nondum est sermo in lingua mea,et ecce, Domine, tu novisti omnia.
PS|139|5|A tergo et a fronte coartasti meet posuisti super me manum tuam.
PS|139|6|Mirabilis nimis facta est scientia tua super me,sublimis, et non attingam eam.
PS|139|7|Quo ibo a spiritu tuoet quo a facie tua fugiam?
PS|139|8|Si ascendero in caelum, tu illic es;si descendero in infernum, ades.
PS|139|9|Si sumpsero pennas auroraeet habitavero in extremis maris,
PS|139|10|etiam illuc manus tua deducet me,et tenebit me dextera tua.
PS|139|11|Si dixero: " Forsitan tenebrae compriment me,et nox illuminatio erit circa me ",
PS|139|12|etiam tenebrae non obscurabuntur a te,et nox sicut dies illuminabiturC sicut tenebrae eius ita et lumen eius -.
PS|139|13|Quia tu formasti renes meos,contexuisti me in utero matris meae.
PS|139|14|Confitebor tibi, quia mirabiliter plasmatus sum;mirabilia opera tua,et anima mea cognoscit nimis.
PS|139|15|Non sunt abscondita ossa mea a te,cum factus sum in occulto,contextus in inferioribus terrae.
PS|139|16|Imperfectum adhuc me viderunt oculi tui,et in libro tuo scripti erant omnes dies:ficti erant, et nondum erat unus ex eis.
PS|139|17|Mihi autem nimis pretiosae cogitationes tuae, Deus;nimis gravis summa earum.
PS|139|18|Si dinumerabo eas, super arenam multiplicabuntur;si ad finem pervenerim, adhuc sum tecum.
PS|139|19|Utinam occidas, Deus, peccatores;viri sanguinum, declinate a me.
PS|139|20|Qui loquuntur contra te maligne:exaltantur in vanum contra te.
PS|139|21|Nonne, qui oderunt te, Domine, oderamet insurgentes in te abhorrebam?
PS|139|22|Perfecto odio oderam illos,et inimici facti sunt mihi.
PS|139|23|Scrutare me, Deus, et scito cor meum;proba me et cognosce semitas meas
PS|139|24|et vide, si via vanitatis in me est,et deduc me in via aeterna.
PS|140|1|Magistro chori. PSALMUS. David.
PS|140|2|Eripe me, Domine, ab homine malo, a viro violentiae serva me.
PS|140|3|Qui cogitaverunt mala in corde,tota die constituebant proelia.
PS|140|4|Acuerunt linguas suas sicut serpentis, venenum aspidum sub labiis eorum.
PS|140|5|Custodi me, Domine, de manu peccatoriset a viro violentiae serva me,qui cogitaverunt supplantare gressus meos.
PS|140|6|Absconderunt superbi laqueum mihiet funes extenderunt in rete,iuxta iter offendicula posuerunt mihi.
PS|140|7|Dixi Domino: " Deus meus es tu;auribus percipe, Domine, vocem deprecationis meae ".
PS|140|8|Domine, Domine, virtus salutis meae,obumbrasti caput meum in die belli.
PS|140|9|Ne concedas, Domine, desideria impii;consilia eius ne perficias.
PS|140|10|Exaltant caput, qui circumdant me;malitia labiorum ipsorum operiat eos.
PS|140|11|Cadant super eos carbones ignis,in foveas deicias eos, et non exsurgant.
PS|140|12|Vir linguosus non firmabitur in terra,virum violentiae mala capient in interitu.
PS|140|13|Cognovi quia faciet Dominus iudicium inopiset vindictam pauperum.
PS|140|14|Verumtamen iusti confitebuntur nomini tuo,et habitabunt recti in conspectu tuo.
PS|141|1|PSALMUS. David.Domine, clamavi ad te, ad me festina;intende voci meae, cum clamo ad te.
PS|141|2|Dirigatur oratio mea sicut incensum in conspectu tuo,elevatio manuum mearum ut sacrificium vespertinum. -
PS|141|3|Pone, Domine, custodiam ori meoet vigiliam ad ostium labiorum meorum.
PS|141|4|Non declines cor meum in verbum malitiaead machinandas machinationes in impietatecum hominibus operantibus iniquitatem;et non comedam ex deliciis eorum.
PS|141|5|Percutiat me iustus in misericordia et increpet me;oleum autem peccatoris non impinguet caput meum,quoniam adhuc et oratio mea in malitiis eorum.
PS|141|6|Deiecti in manus duras iudicum eorum,audient verba mea, quoniam suavia erant.
PS|141|7|Sicut frusta dolantis et dirumpentis in terra,dissipata sunt ossa eorum ad fauces inferni.
PS|141|8|Quia ad te, Domine, Domine, oculi mei;ad te confugi, non effundas animam meam.
PS|141|9|Custodi me a laqueo, quem statuerunt mihi,et a scandalis operantium iniquitatem.
PS|141|10|Cadent in retiacula sua peccatores simul,ego autem ultra pertranseam.
PS|142|1|Maskil. David, cum esset in caverna. Precatio.
PS|142|2|Voce mea ad Dominum clamo,voce mea ad Dominum deprecor;
PS|142|3|effundo in conspectu eius lamentationem meam,et tribulationem meam ante ipsum pronuntio.
PS|142|4|Cum deficit in me spiritus meus,tu nosti semitas meas.In via, qua ambulabam,absconderunt laqueum mihi.
PS|142|5|Considerabam ad dexteram et videbam,et non erat qui cognosceret me.Periit fuga a me,et non est qui requirat animam meam. -
PS|142|6|Clamavi ad te, Domine;dixi: " Tu es refugium meum,portio mea in terra viventium.
PS|142|7|Intende ad deprecationem meam,quia humiliatus sum nimis.Libera me a persequentibus me,quia confortati sunt super me.
PS|142|8|Educ de custodia animam meamad confitendum nomini tuo;me circumdabunt iusti,cum retribueris mihi ".
PS|143|1|PSALMUS. David.Domine, exaudi orationem meam, auribus percipe obsecrationem meam in veritate tua;exaudi me in tua iustitia.
PS|143|2|Et non intres in iudicium cum servo tuo,quia non iustificabitur in conspectu tuo omnis vivens.
PS|143|3|Quia persecutus est inimicus animam meam,contrivit in terra vitam meam,collocavit me in obscuris sicut mortuos a saeculo.
PS|143|4|Et anxiatus est in me spiritus meus,in medio mei obriguit cor meum.
PS|143|5|Memor fui dierum antiquorum,meditatus sum in omnibus operibus tuis,in factis manuum tuarum recogitabam.
PS|143|6|Expandi manus meas ad te,anima mea sicut terra sine aqua tibi.
PS|143|7|Velociter exaudi me, Domine;defecit spiritus meus.Non abscondas faciem tuam a me,ne similis fiam descendentibus in lacum.
PS|143|8|Auditam fac mihi mane misericordiam tuam,quia in te speravi.Notam fac mihi viam, in qua ambulem,quia ad te levavi animam meam.
PS|143|9|Eripe me de inimicis meis,Domine, ad te confugi.
PS|143|10|Doce me facere voluntatem tuam,quia Deus meus es tu.Spiritus tuus bonus deducet me in terram rectam;
PS|143|11|propter nomen tuum, Domine, vivificabis me.In iustitia tua educes de tribulatione animam meam
PS|143|12|et in misericordia tua disperdes inimicos meos;et perdes omnes, qui tribulant animam meam,quoniam ego servus tuus sum.
PS|144|1|David.Benedictus Dominus, adiutor meus,qui docet manus meas ad proeliumet digitos meos ad bellum.
PS|144|2|Misericordia mea et fortitudo mea,refugium meum et liberator meus;scutum meum, et in ipso speravi,qui subdit populum meum sub me.
PS|144|3|Domine, quid est homo, quod agnoscis eum,aut filius hominis, quod reputas eum?
PS|144|4|Homo vanitati similis factus est,dies eius sicut umbra praeteriens.
PS|144|5|Domine, inclina caelos tuos et descende;tange montes, et fumigabunt.
PS|144|6|Fulgura coruscationem et dissipa eos;emitte sagittas tuas et conturba eos.
PS|144|7|Emitte manum tuam de alto;eripe me et libera me de aquis multis,de manu filiorum alienigenarum,
PS|144|8|quorum os locutum est vanitatem,et dextera eorum dextera mendacii.
PS|144|9|Deus, canticum novum cantabo tibi,in psalterio decachordo psallam tibi,
PS|144|10|qui das salutem regibus,qui redimis David servum tuum de gladio maligno.
PS|144|11|Eripe me et libera mede manu filiorum alienigenarum,quorum os locutum est vanitatem,et dextera eorum dextera mendacii.
PS|144|12|Filii nostri sicut novellae crescentesin iuventute sua;filiae nostrae sicut columnae angulares,sculptae ut structura templi.
PS|144|13|Promptuaria nostra plena,redundantia omnibus bonis;oves nostrae in milibusinnumerabiles in campis nostris,
PS|144|14|boves nostrae crassae.Non est ruina maceriae neque egressusneque clamor in plateis nostris.
PS|144|15|Beatus populus, cui haec sunt;beatus populus, cui Dominus est Deus.
PS|145|1|Laudes. David.ALEPH. Exaltabo te, Deus meus, rex,et benedicam nomini tuoin saeculum et in saeculum saeculi.
PS|145|2|BETH. Per singulos dies benedicam tibiet laudabo nomen tuumin saeculum et in saeculum saeculi.
PS|145|3|GHIMEL. Magnus Dominus et laudabilis nimis,et magnitudinis eius non est investigatio.
PS|145|4|DALETH. Generatio generationi laudabit opera tua,et potentiam tuam pronuntiabunt.
PS|145|5|HE. Magnificentiam gloriae maiestatis tuae loquenturet mirabilia tua enarrabunt.
PS|145|6|VAU. Et virtutem terribilium tuorum dicentet magnitudinem tuam narrabunt.
PS|145|7|ZAIN. Memoriam abundantiae suavitatis tuae eructabuntet iustitia tua exsultabunt.
PS|145|8|HETH. Miserator et misericors Dominus,longanimis et multae misericordiae.
PS|145|9|TETH. Suavis Dominus universis,et miserationes eius super omnia opera eius.
PS|145|10|IOD. Confiteantur tibi, Domine, omnia opera tua;et sancti tui benedicant tibi.
PS|145|11|CAPH. Gloriam regni tui dicantet potentiam tuam loquantur,
PS|145|12|LAMED. ut notas faciant filiis hominum potentias tuaset gloriam magnificentiae regni tui.
PS|145|13|MEM. Regnum tuum regnum omnium saeculorum,et dominatio tua in omnem generationem et generationem.NUN. Fidelis Dominus in omnibus verbis suiset sanctus in omnibus operibus suis.
PS|145|14|SAMECH. Allevat Dominus omnes, qui corruunt,et erigit omnes depressos.
PS|145|15|AIN. Oculi omnium in te sperant,et tu das illis escam in tempore opportuno.
PS|145|16|PHE. Aperis tu manum tuamet imples omne animal in beneplacito.
PS|145|17|SADE. Iustus Dominus in omnibus viis suiset sanctus in omnibus operibus suis.
PS|145|18|COPH. Prope est Dominus omnibus invocantibus eum,omnibus invocantibus eum in veritate.
PS|145|19|RES. Voluntatem timentium se facietet deprecationem eorum exaudiet et salvos faciet eos.
PS|145|20|SIN. Custodit Dominus omnes diligentes seet omnes peccatores disperdet.
PS|145|21|TAU. Laudationem Domini loquetur os meum,et benedicat omnis caro nomini sancto eiusin saeculum et in saeculum saeculi.
PS|146|1|ALLELUIA.Lauda, anima mea, Dominum;
PS|146|2|laudabo Dominum in vita mea,psallam Deo meo, quamdiu fuero.
PS|146|3|Nolite confidere in principibus,in filiis hominum, in quibus non est salus.
PS|146|4|Exibit spiritus eius, et revertetur in terram suam;in illa die peribunt cogitationes eorum.
PS|146|5|Beatus, cuius Deus Iacob est adiutor,cuius spes in Domino Deo suo,
PS|146|6|qui fecit caelum et terram,mare et omnia, quae in eis sunt;qui custodit veritatem in saeculum,
PS|146|7|facit iudicium oppressis,dat escam esurientibus.Dominus solvit compeditos,
PS|146|8|Dominus illuminat caecos,Dominus erigit depressos,Dominus diligit iustos,
PS|146|9|Dominus custodit advenas,pupillum et viduam sustentatet viam peccatorum disperdit.
PS|146|10|Regnabit Dominus in saecula,Deus tuus, Sion,in generationem et generationem.
PS|147|1|ALLELUIA.Laudate Dominum, quoniam bonum est psallere Deo nostro,quoniam iucundum est celebrare laudem.
PS|147|2|Aedificans Ierusalem Dominus,dispersos Israelis congregabit.
PS|147|3|Qui sanat contritos cordeet alligat plagas eorum;
PS|147|4|qui numerat multitudinem stellarumet omnibus eis nomina vocat.
PS|147|5|Magnus Dominus noster et magnus virtute,sapientiae eius non est numerus.
PS|147|6|Sustentat mansuetos Dominus,humilians autem peccatores usque ad terram.
PS|147|7|Praecinite Domino in confessione,psallite Deo nostro in cithara.
PS|147|8|Qui operit caelum nubibuset parat terrae pluviam.Qui producit in montibus fenumet herbam servituti hominum.
PS|147|9|Qui dat iumentis escam ipsorumet pullis corvorum invocantibus eum.
PS|147|10|Non in fortitudine equi delectatur,nec in tibiis viri beneplacitum est ei.
PS|147|11|Beneplacitum est Domino super timentes eumet in eis, qui sperant super misericordia eius.
PS|147|12|Lauda, Ierusalem, Dominum;collauda Deum tuum, Sion.
PS|147|13|Quoniam confortavit seras portarum tuarum,benedixit filiis tuis in te.
PS|147|14|Qui ponit fines tuos pacemet adipe frumenti satiat te.
PS|147|15|Qui emittit eloquium suum terrae,velociter currit verbum eius.
PS|147|16|Qui dat nivem sicut lanam,pruinam sicut cinerem spargit.
PS|147|17|Mittit crystallum suam sicut buccellas;ante faciem frigoris eius quis sustinebit?
PS|147|18|Emittet verbum suum et liquefaciet ea,flabit spiritus eius, et fluent aquae.
PS|147|19|Qui annuntiat verbum suum Iacob,iustitias et iudicia sua Israel.
PS|147|20|Non fecit taliter omni nationiet iudicia sua non manifestavit eis. ALLELUIA.
PS|148|1|ALLELUIA.Laudate Dominum de caelis,laudate eum in excelsis.
PS|148|2|Laudate eum, omnes angeli eius,laudate eum, omnes virtutes eius.
PS|148|3|Laudate eum, sol et luna,laudate eum, omnes stellae lucentes.
PS|148|4|Laudate eum, caeli caelorumet aquae omnes, quae super caelos sunt. -
PS|148|5|Laudent nomen Domini,quia ipse mandavit, et creata sunt;
PS|148|6|statuit ea in aeternum et in saeculum saeculi;praeceptum posuit, et non praeteribit.
PS|148|7|Laudate Dominum de terra,dracones et omnes abyssi,
PS|148|8|ignis, grando, nix, fumus,spiritus procellarum, qui facit verbum eius,
PS|148|9|montes et omnes colles,ligna fructifera et omnes cedri,
PS|148|10|bestiae et universa pecora,serpentes et volucres pennatae.
PS|148|11|Reges terrae et omnes populi,principes et omnes iudices terrae,
PS|148|12|iuvenes et virgines,senes cum iunioribus
PS|148|13|laudent nomen Domini,quia exaltatum est nomen eius solius.Magnificentia eius super caelum et terram,
PS|148|14|et exaltavit cornu populi sui.Hymnus omnibus sanctis eius,filiis Israel, populo, qui propinquus est ei. ALLELUIA.
PS|149|1|ALLELUIA.Cantate Domino canticum novum;laus eius in ecclesia sanctorum.
PS|149|2|Laetetur Israel in eo, qui fecit eum,et filii Sion exsultent in rege suo.
PS|149|3|Laudent nomen eius in choro,in tympano et cithara psallant ei,
PS|149|4|quia beneplacitum est Domino in populo suo,et honorabit mansuetos in salute.
PS|149|5|Iubilent sancti in gloria,laetentur in cubilibus suis.
PS|149|6|Exaltationes Dei in gutture eorum,et gladii ancipites in manibus eorum,
PS|149|7|ad faciendam vindictam in nationibus,castigationes in populis,
PS|149|8|ad alligandos reges eorum in compedibuset nobiles eorum in manicis ferreis,
PS|149|9|ad faciendum in eis iudicium conscriptum.Gloria haec est omnibus sanctis eius. ALLELUIA.
PS|150|1|ALLELUIA.Laudate Dominum in sanctuario eius,laudate eum in firmamento virtutis eius.
PS|150|2|Laudate eum in magnalibus eius,laudate eum secundum multitudinem magnitudinis eius.
PS|150|3|Laudate eum in sono tubae,laudate eum in psalterio et cithara,
PS|150|4|laudate eum in tympano et choro,laudate eum in chordis et organo,
PS|150|5|laudate eum in cymbalis benesonantibus,laudate eum in cymbalis iubilationis:omne quod spirat, laudet Dominum. ALLELUIA.
