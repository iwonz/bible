1COR|1|1|奉上帝旨意，蒙召作基督耶穌使徒的 保羅 ，同弟兄 所提尼 ，
1COR|1|2|寫信給在 哥林多 上帝的教會—就是在基督耶穌裏成聖、蒙召作聖徒的—以及所有在各處求告我主耶穌基督之名的人。基督是他們的主，也是我們的主。
1COR|1|3|願恩惠、平安 從我們的父上帝並主耶穌基督歸給你們！
1COR|1|4|我常為你們感謝我的上帝，因上帝在基督耶穌裏所賜給你們的恩惠。
1COR|1|5|因為你們在他裏面凡事富足，具有各種口才、各樣知識，
1COR|1|6|正如我為基督作的見證在你們心裏得以堅固，
1COR|1|7|以致你們在恩賜上一無欠缺，切切等候我們主耶穌基督的顯現。
1COR|1|8|他也必堅固你們到底，使你們在我們主耶穌基督 的日子無可指責。
1COR|1|9|上帝是信實的，他呼召你們好與他兒子—我們的主耶穌基督—共享團契。
1COR|1|10|弟兄們，我藉我們主耶穌基督的名勸你們說話要一致。你們中間不可分裂，只要一心一意彼此團結。
1COR|1|11|我的弟兄們， 革來 氏家裏的人曾對我提起你們，說你們中間有紛爭。
1COR|1|12|我的意思是，你們各人說：「我是屬 保羅 的」；「我是屬 亞波羅 的」；「我是屬 磯法 的」；「我是屬基督的。」
1COR|1|13|基督是分裂的嗎？ 保羅 為你們釘了十字架嗎？你們是奉 保羅 的名受了洗嗎？
1COR|1|14|我感謝上帝 ，除了 基利司布 和 該猶 以外，我沒有給你們中的任何一個人施洗，
1COR|1|15|免得有人說你們是奉我的名受洗的。
1COR|1|16|我曾為 司提法那 家施過洗；此外我已記不清有沒有給別人施過洗。
1COR|1|17|因為基督差遣我不是為施洗，而是為傳福音；並不是用智慧的言論，免得基督的十字架落了空。
1COR|1|18|因為十字架的道理，在那滅亡的人是愚拙，在我們得救的人卻是上帝的大能。
1COR|1|19|就如經上所記： 「我要摧毀智慧人的智慧， 廢棄聰明人的聰明。」
1COR|1|20|智慧人在哪裏？文士在哪裏？這世上的辯士在哪裏？上帝豈不是已使這世上的智慧變成愚拙了嗎？
1COR|1|21|既然世人憑自己的智慧不認識上帝，上帝就本著自己的智慧樂意藉著人所傳愚拙的話拯救那些信的人。
1COR|1|22|猶太 人要的是神蹟， 希臘 人求的是智慧，
1COR|1|23|我們卻是傳被釘十字架的基督，這對 猶太 人是絆腳石，對外邦人是愚拙；
1COR|1|24|但對那蒙召的，無論是 猶太 人、 希臘 人，基督總是上帝的大能，上帝的智慧。
1COR|1|25|因為，上帝的愚拙總比人智慧；上帝的軟弱總比人強壯。
1COR|1|26|弟兄們哪，想一想你們的蒙召，按著人的觀點，有智慧的不多，有能力的不多，有尊貴地位的也不多。
1COR|1|27|但是，上帝揀選了世上愚拙的，為了使有智慧的羞愧；又揀選了世上軟弱的，為了使強壯的羞愧。
1COR|1|28|上帝也揀選了世上卑賤的，被人厭惡的，以及那一無所有的，為要廢掉那樣樣都有的，
1COR|1|29|使凡血肉之軀的，在上帝面前，一個也不能自誇。
1COR|1|30|但你們得以在基督耶穌裏是本乎上帝，他使基督成為我們的智慧，成為公義、聖潔、救贖。
1COR|1|31|如經上所記：「要誇耀的，該誇耀主。」
1COR|2|1|弟兄們，從前我到你們那裏去，並沒有用高言大智對你們宣講上帝的奧祕。
1COR|2|2|因為我曾定了主意，在你們中間不知道別的，只知道耶穌基督並他釘十字架。
1COR|2|3|我在你們那裏時，又軟弱，又懼怕，又戰戰兢兢。
1COR|2|4|我說的話、講的道不是用委婉智慧的言語 ，而是以聖靈的大能來證明，
1COR|2|5|為要使你們的信不靠著人的智慧，而是靠著上帝的大能。
1COR|2|6|然而，在成熟的人中，我們也講智慧，但不是今世的智慧，也不是今世有權有位、將要滅亡的人的智慧。
1COR|2|7|我們講的是從前隱藏的、上帝奧祕的智慧，就是上帝在萬世以前預定使我們得榮耀的智慧；
1COR|2|8|這智慧，今世有權有位的人沒有一個知道，若知道，他們就不會把榮耀的主釘在十字架上了。
1COR|2|9|如經上所記： 「上帝為愛他的人所預備的 是眼睛未曾看見，耳朵未曾聽見， 人心也未曾想到的。」
1COR|2|10|只有上帝藉著聖靈把這事向我們顯明了；因為聖靈參透萬事，就是上帝深奧的事也參透了。
1COR|2|11|除了在人裏頭的靈，誰知道人的事？照樣，除了上帝的靈，也沒有人知道上帝的事。
1COR|2|12|我們所領受的並不是世上的靈，而是從上帝來的靈，為使我們知道上帝把恩賜賞給我們的事。
1COR|2|13|我們也講說這些事，不是用人的智慧所教的言語，而是用聖靈所教的言語，用屬靈的話解釋屬靈的事 。
1COR|2|14|然而，屬血氣的人不接受上帝的靈的事，他反倒以這為愚拙，並且他不能了解，因為這些事惟有屬靈的人才能領悟。
1COR|2|15|屬靈的人能看透萬事，卻沒有一人能看透他。
1COR|2|16|「誰曾知道主的心？ 誰會教導他？」 至於我們，我們有基督的心。
1COR|3|1|弟兄們，我從前對你們說話，還不能把你們當作屬靈的，只能把你們當作屬肉體的，你們在基督裏僅是嬰孩。
1COR|3|2|我用奶餵你們，沒有用飯餵你們，因為那時你們不能吃。就是如今還是不能，
1COR|3|3|因為你們仍是屬肉體的。你們中間有嫉妒、紛爭，這豈不是屬乎肉體，照著世人的樣子生活嗎？
1COR|3|4|有人說：「我是屬 保羅 的」；有人說：「我是屬 亞波羅 的」；這樣你們豈不是和世人一樣嗎？
1COR|3|5|亞波羅 算甚麼？ 保羅 算甚麼？我們都是上帝的執事，藉著我們，你們信了；這不過是照著主給各人的恩賜去做罷了。
1COR|3|6|我栽種了， 亞波羅 澆灌了，惟有上帝使它生長。
1COR|3|7|可見，栽種的算不了甚麼，澆灌的也算不了甚麼；惟有上帝能使它生長。
1COR|3|8|栽種的和澆灌的都是一樣，但將來各人要照自己的勞苦得到自己的報酬。
1COR|3|9|因為我們是上帝的同工，而你們是上帝的田地、上帝的房屋。
1COR|3|10|我照上帝所給我的恩典，好像一個聰明的工頭，立好了根基，別人在上面建造；只是各人要謹慎怎樣在上面建造。
1COR|3|11|因為，那已經立好的根基就是耶穌基督，此外沒有人能立別的根基。
1COR|3|12|若有人用金銀、寶石，草木、禾秸，在這根基上建造，
1COR|3|13|各人的工程必將顯露，因為那日子要將它顯明，有火把它暴露出來，這火要試煉各人的工程怎樣。
1COR|3|14|人在那根基上所建造的工程若能保得住，他將要得賞賜。
1COR|3|15|人的工程若被燒了，他將損失，雖然他自己將得救，卻要像從火裏經過一樣。
1COR|3|16|難道不知你們是上帝的殿，上帝的靈住在你們裏面嗎？
1COR|3|17|若有人毀壞上帝的殿，上帝一定要毀滅那人；因為上帝的殿是神聖的，這殿就是你們。
1COR|3|18|誰都不可自欺。你們中間若有人自以為在今世有智慧，倒不如變為愚拙，好成為有智慧的。
1COR|3|19|因為這世界的智慧在上帝看來是愚拙的。如經上記著： 「主使有智慧的人中了自己的詭計；」
1COR|3|20|又說： 「主知道智慧人的意念， 因為它們是虛妄的。」
1COR|3|21|所以，無論誰都不可誇耀人；因為萬有都是你們的，
1COR|3|22|或 保羅 ，或 亞波羅 ，或 磯法 ，或世界，或生，或死，或現今的事，或將來的事，全是你們的，
1COR|3|23|而你們是屬基督的，基督是屬上帝的。
1COR|4|1|人應該把我們看為基督的執事，為上帝的奧祕的管家。
1COR|4|2|所求於管家的，是要他忠心。
1COR|4|3|我被你們評斷，或被別人評斷，我都以為是極小的事；連我自己也不評斷自己。
1COR|4|4|雖然我不覺得自己有錯，卻也不能因此判為無罪；審斷我的是主。
1COR|4|5|所以，時候未到，在主來以前甚麼都不要評斷，他要照出暗中的隱情，揭發人的動機。那時，各人要從上帝那裏得著稱讚。
1COR|4|6|弟兄們，為你們的緣故，我拿這些事應用到我自己和 亞波羅 身上，讓你們從我們學到「不可過於聖經所記」這話的意思，免得你們自高自大，看重這個，看輕那個。
1COR|4|7|使你與人不同的是誰呢？你所有的有哪一個不是領受的呢？若是領受的，為何自誇，彷彿不是領受的呢？
1COR|4|8|你們已經飽足了，已經富足了，用不著我們，自己就作王了。我願意你們果真作王，讓我們也可以與你們一同作王！
1COR|4|9|我想，上帝把我們作使徒的明顯地列在末後，好像定死罪的囚犯，因為我們成了一臺戲，給世界、天使和眾人觀看。
1COR|4|10|我們為基督的緣故成為愚拙的；你們在基督裏倒是聰明的。我們軟弱，你們倒強壯；你們有榮耀，我們倒被藐視。
1COR|4|11|直到如今，我們還是又飢又渴，又赤身露體，又挨打，又到處漂泊，
1COR|4|12|並且勞碌，親手做工；被人咒罵，我們就祝福；被人迫害，我們就忍受；
1COR|4|13|被人毀謗，我們就勸導。直到如今，人還把我們看作世上的污穢，萬物中的渣滓。
1COR|4|14|我寫這些話，不是要使你們羞愧，而是要警戒你們，好像我所愛的兒女一樣。
1COR|4|15|雖然你們在基督裏有無數的導師，卻沒有許多父親，因我是在基督耶穌裏用福音生了你們。
1COR|4|16|所以，我求你們要效法我。
1COR|4|17|因此，我已差 提摩太 到你們那裏去。他在主裏面是我親愛和忠心的兒子；他要提醒你們，我在基督耶穌 裏怎樣行事為人，在各處各教會中怎樣教導人。
1COR|4|18|有些人以為我不到你們那裏去而自高自大。
1COR|4|19|但是，主若准許，我會很快到你們那裏去；我所要知道的，不是那些自高自大者的言語，而是他們的權能。
1COR|4|20|因為上帝的國不在乎言語，而在乎權能。
1COR|4|21|你們願意怎麼樣呢？要我帶著棍子到你們那裏去呢，還是帶著慈愛溫柔的心呢？
1COR|5|1|我確實聽說在你們中間有淫亂的事；這種淫亂連外邦人中也沒有，就是有人和他的繼母同居。
1COR|5|2|你們還自高自大！你們不是該覺得痛心，把做這事的人從你們中間趕出去嗎？
1COR|5|3|我人雖然不在你們那裏，心卻在你們那裏，好像親自與你們同在。我奉我們主耶穌 的名，已經判斷了做這事的人。你們聚會的時候，我的心和你們同在。你們藉著我們主耶穌的權能，
1COR|5|4|
1COR|5|5|要把這樣的人交給撒但，使他的肉體敗壞，好讓他的靈魂在主的日子可以得救。
1COR|5|6|你們這樣自誇是不好的。你們不知道一點麵酵能使全團發起來嗎？
1COR|5|7|既然你們是無酵的麵，要把舊酵除淨，好使你們成為新團；因為我們逾越節的羔羊—基督已經被殺獻為祭牲了。
1COR|5|8|所以，我們來守這節，不可用舊酵，就是不可用惡毒、邪惡的酵，只用純潔真實的無酵餅。
1COR|5|9|我先前寫信告訴過你們，不可與淫亂的人交往。
1COR|5|10|此話不是泛指這世上所有行淫亂的，或貪婪的，勒索的，或拜偶像的；若是這樣，你們非離開這世界不可。
1COR|5|11|但現在，我寫信告訴你們，若有稱為弟兄的人卻仍犯淫亂，或貪婪，或拜偶像，或辱罵，或醉酒，或勒索，這樣的人不可跟他交往，就是跟他吃飯都不可以。
1COR|5|12|因為審判教外的人與我何干？教內的人豈不是你們要審判嗎？
1COR|5|13|至於外人有上帝審判他們。如經上說：「要從你們中間把那邪惡的人趕出去。」
1COR|6|1|你們中間有彼此爭吵的事，怎敢告到不義的人面前，而不告到聖徒面前呢？
1COR|6|2|你們豈不知聖徒要審判世界嗎？若世界要受你們的審判，難道你們不配審判這最小的事嗎？
1COR|6|3|你們豈不知我們要審判天使嗎？何況今生的事呢！
1COR|6|4|既是這樣，你們若有今生當審判的事，會讓教會所輕看的人來審判嗎？
1COR|6|5|我說這話是要使你們慚愧。難道你們中間沒有一個有智慧的人能審斷弟兄中的事嗎？
1COR|6|6|你們竟然有弟兄去告弟兄，而且告到不信主的人面前。
1COR|6|7|你們彼此告狀，這已經是你們的大錯了。為甚麼不情願受冤屈呢？為甚麼不情願吃虧呢？
1COR|6|8|你們反倒去冤枉人，虧負人，況且所冤枉所虧負的就是弟兄。
1COR|6|9|你們豈不知不義的人不能承受上帝的國嗎？不要自欺！無論是淫亂的、拜偶像的、姦淫的、作娼妓 的，親男色的、
1COR|6|10|偷竊的、貪婪的、醉酒的、辱罵的、勒索的，都不能承受上帝的國。
1COR|6|11|從前你們中間也有人是這樣；但現在你們奉主耶穌基督 的名，並藉著我們上帝的靈，已經洗淨，已經成聖，已經稱義了。
1COR|6|12|「凡事我都可行」，但不是凡事都有益處。「凡事我都可行」，但無論哪一件，我都不受它的轄制。
1COR|6|13|「食物是為肚腹，肚腹是為食物」；但上帝要使這兩樣都毀壞。身體不是為淫亂，而是為主；主也是為身體。
1COR|6|14|上帝已經使主復活，也要用他自己的能力使我們復活。
1COR|6|15|你們豈不知道你們的身體是基督的肢體嗎？我可以把基督的肢體作為娼妓的肢體嗎？絕對不可！
1COR|6|16|你們豈不知道與娼妓苟合的，就是與她成為一體嗎？因為主說：「二人要成為一體。」
1COR|6|17|但與主聯合的，就是與主成為一靈。
1COR|6|18|你們要遠避淫行。人所犯的，無論甚麼罪，都在身體以外；惟有行淫的，是得罪自己的身體。
1COR|6|19|你們豈不知道你們的身體是聖靈的殿嗎？這聖靈是從上帝而來，住在你們裏面的。而且你們不是屬自己的人，
1COR|6|20|因為你們是重價買來的。所以，要在你們的身體上榮耀上帝。
1COR|7|1|關於你們信上所提的事，男人不親近女人倒好。
1COR|7|2|但為了避免淫亂的事，男人當各有自己的妻子，女人也當各有自己的丈夫。
1COR|7|3|丈夫對妻子要盡本分；妻子對丈夫也要如此。
1COR|7|4|妻子對自己的身體沒有主張的權柄，權柄在丈夫；丈夫對自己的身體也沒有主張的權柄，權柄在妻子。
1COR|7|5|夫妻不可忽略對方的需求，除非為了要專心禱告，在兩相情願下暫時分房；以後仍要同房，免得撒但趁著你們情不自禁而引誘你們。
1COR|7|6|我說這話是出於容忍，不是命令。
1COR|7|7|我願眾人像我一樣；但是各人都有來自上帝的恩賜，一個是這樣，一個是那樣。
1COR|7|8|我對沒有嫁娶的和寡婦說，他們若能維持獨身像我一樣就好。
1COR|7|9|但他們若不能自制，就應該嫁娶，與其慾火攻心，倒不如結婚為妙。
1COR|7|10|至於那已經嫁娶的，我吩咐他們—其實不是我，而是主吩咐的：妻子不可離開丈夫，
1COR|7|11|若是離開了，不可再嫁，不然要跟丈夫復和；丈夫也不可離棄妻子。
1COR|7|12|我對其餘的人說—是我，不是主說—倘若某弟兄有不信的妻子，妻子也情願和他一起生活，他就不可離棄妻子。
1COR|7|13|妻子有不信的丈夫，丈夫也情願和她一起生活，她就不可離棄丈夫。
1COR|7|14|因為不信的丈夫會因著妻子成了聖潔；不信的妻子也會因著丈夫 成了聖潔。不然，你們的兒女就不潔淨了，但現在他們是聖潔的。
1COR|7|15|倘若那不信的人要離開，就由他離開吧！無論是弟兄是姊妹，遇著這樣的事都不必拘束。上帝召你們原是要你們和睦。
1COR|7|16|你這作妻子的怎麼知道不能救你的丈夫呢？你這作丈夫的怎麼知道不能救你的妻子呢？
1COR|7|17|無論如何，要照主所分給各人的恩賜和上帝所召各人的情況生活。我在各教會裏都是這樣規定的。
1COR|7|18|有人受割禮後才蒙召，他就不必除去割禮的記號。有人未受割禮前蒙召，他就不必受割禮。
1COR|7|19|受割禮算不了甚麼，不受割禮也算不了甚麼，只要謹守上帝的誡命就是了。
1COR|7|20|各人蒙召的時候是甚麼身份，要守住這身份。
1COR|7|21|你是作奴隸時蒙召的嗎？不要介意；若能獲得自由，就爭取自由更好。
1COR|7|22|因為，蒙主呼召的奴僕是主所釋放的人；蒙主呼召的自由之人是基督的奴僕。
1COR|7|23|你們是重價買來的；不要作人的奴僕。
1COR|7|24|弟兄們，你們各人蒙召的時候是甚麼身份，要在上帝面前守住這身份。
1COR|7|25|關於未婚女子，我沒有主的命令，但我既蒙主憐憫、作為一個可信靠的人，把自己的意見告訴你們。
1COR|7|26|因現今的艱難，據我看來，人不如安於現狀。
1COR|7|27|你已經有了妻子，就不要求擺脫；你還沒有妻子，就不要想娶妻。
1COR|7|28|你若娶妻，並不是犯罪；未婚女子若出嫁，也不是犯罪。然而，這等人會遭受肉身上的苦難，我寧願你們免受這苦難。
1COR|7|29|弟兄們，我是說：時候不多了。從此以後，那有妻子的，要像沒有一樣；
1COR|7|30|哀哭的，不像在哀哭；快樂的，不像在快樂；購買的，像一無所得；
1COR|7|31|享受這世界的，不像在享受這世界；因為這世界的局面將要過去了。
1COR|7|32|我願你們一無掛慮。沒有結婚的是為主的事掛慮，想怎樣令主喜悅；
1COR|7|33|結了婚的是為世上的事掛慮，想怎樣讓妻子喜悅，
1COR|7|34|於是，他就分心了。沒有結婚的和未婚的女子是為主的事掛慮，為要身體和心靈都聖潔；已經出嫁的是為世上的事掛慮，想怎樣讓丈夫喜悅。
1COR|7|35|我說這話是為你們的益處，不是要限制你們，而是要你們做合宜的事，得以不分心地對主忠誠。
1COR|7|36|若有人認為自己待他的女兒 不合宜，女兒也過了適婚年齡 ，他可以隨意處理，不算有罪，讓兩人結婚就是了。
1COR|7|37|倘若有人心裏堅定，沒有不得已的事，並且由得自己作主，心裏又決定了不讓女兒結婚 ，這樣做也好。
1COR|7|38|這樣看來，讓自己的女兒結婚 固然是好，不讓她結婚更好。
1COR|7|39|丈夫活著的時候，妻子是受約束的；丈夫若長眠了，妻子就自由了，可以隨意再嫁，只是要嫁給主裏面的人。
1COR|7|40|然而，按我的意見，她若能守節就更有福氣。我想我自己也有上帝的靈的感動。
1COR|8|1|關於祭過偶像的食物，我們曉得「我們都有知識」，但知識使人自高自大，惟有愛心能造就人。
1COR|8|2|若有人自以為知道甚麼，他其實仍不知道他所應當知道的。
1COR|8|3|若有人愛上帝，他就是上帝所認識的人了。
1COR|8|4|關於吃祭過偶像的食物，我們知道「偶像在世上算不得甚麼」；也知道「上帝只有一位，沒有別的」。
1COR|8|5|雖然在天上或地上有許多所謂的神明，就如他們中間有許多的神明，許多的主，
1COR|8|6|但是我們只有一位上帝，就是父，萬物都出於他，我們也歸於他；並只有一位主，就是耶穌基督，萬物都是藉著他而有，我們也是藉著他而有。
1COR|8|7|可是，不是人人都有這知識。有人到現在因拜慣了偶像，仍以為所吃的是祭過偶像的食物；既然他們的良心軟弱，也就污穢了。
1COR|8|8|其實，食物不能使我們更接近上帝，因為我們不吃也無損，吃也無益。
1COR|8|9|可是，你們要謹慎，免得你們這自由竟成了軟弱人的絆腳石。
1COR|8|10|若有人見你這有知識的在偶像的廟裏坐席，而這人的良心是軟弱的，他豈不放膽去吃那祭過偶像的食物嗎？
1COR|8|11|因此，基督為他死的那軟弱弟兄，也就因你的知識沉淪了。
1COR|8|12|你們這樣得罪弟兄，傷了他們軟弱的良心，就是得罪基督。
1COR|8|13|所以，食物若使我的弟兄跌倒，我就永遠不吃肉，免得使我的弟兄跌倒了。
1COR|9|1|我不是自由的嗎？我不是使徒嗎？我不是見過我們的主耶穌嗎？你們不是我在主裏面工作的成果嗎？
1COR|9|2|假若對別人來說，我不是使徒，對你們來說，我總是使徒；因為你們在主裏正是我作使徒的印證。
1COR|9|3|對那些質問我的人，這就是我的答辯。
1COR|9|4|難道我們沒有權利靠著傳福音吃喝嗎？
1COR|9|5|難道我們沒有權利帶著信主的妻子一起出入，如同其餘的使徒，和主的兄弟們，和 磯法 一樣嗎？
1COR|9|6|只有我和 巴拿巴 沒有權利不做工嗎？
1COR|9|7|有誰當兵而自備糧餉呢？有誰栽葡萄園而不吃園裏的果子呢？有誰牧養牛羊而不喝牛羊的奶呢？
1COR|9|8|我說這些話豈是照一般人的看法？律法不也是這樣說嗎？
1COR|9|9|就如 摩西 的律法記著：「牛在踹穀的時候，不可籠住牠的嘴。」難道上帝所掛念的是牛嗎？
1COR|9|10|他不全是為我們說的嗎？的確是為我們說的！因為耕種的要存著指望去耕種；收割的也要存著分享穀物的指望去收割。
1COR|9|11|我們既然把屬靈的種子撒在你們中間，若從你們收取養生之物，這還算大事嗎？
1COR|9|12|假如別人在你們身上享有這權利，何況我們呢？ 然而，我們並沒有用過這權利，倒是凡事忍受，免得基督的福音受到阻礙。
1COR|9|13|你們豈不知在聖殿供職的人吃聖殿中的食物嗎？在祭壇伺候的人分享壇上的供物嗎？
1COR|9|14|主也是這樣命令，要傳福音的人靠著福音養生。
1COR|9|15|但這權利我全然沒有用過。我寫這些話，並非要你們這樣待我，因為我寧可死也不讓人使我所誇的落了空。
1COR|9|16|我傳福音原沒有可誇耀的，因為我是不得已的，若不傳福音，我就有禍了。
1COR|9|17|我若甘心做這事，就有賞賜；若不甘心，責任卻已經託付給我了。
1COR|9|18|這樣，我的賞賜是甚麼呢？就是我傳福音的時候，使人不花錢得福音，免得我用盡了傳福音的權利。
1COR|9|19|我雖然是自由的，不受人管轄，但我甘心作了眾人的僕人，為贏得更多的人。
1COR|9|20|對 猶太 人，我就作 猶太 人，為要贏得 猶太 人；對律法以下的人，我雖不在律法以下，還是作律法以下的人，為要贏得律法以下的人。
1COR|9|21|對沒有律法的人，我就作沒有律法的人，為要贏得沒有律法的人；其實我在上帝面前，不是沒有律法，而是在基督的律法之下。
1COR|9|22|對軟弱的人，我就作軟弱的人，為要贏得軟弱的人。對甚麼樣的人，我就作甚麼樣的人。無論如何我總要救一些人。
1COR|9|23|凡我所做的，都是為福音的緣故，為要與人共享這福音的好處。
1COR|9|24|你們不知道在運動場上賽跑的，大家都跑，但得獎賞的只有一人？你們也要這樣跑，好使你們得著獎賞。
1COR|9|25|凡參加競賽的，在各方面都要有節制，他們不過是要得會朽壞的冠冕；我們卻是要得不會朽壞的冠冕。
1COR|9|26|所以，我奔跑，不像無目標的；我鬥拳，不像打空氣的。
1COR|9|27|我克制己身，使它完全順服，免得我傳福音給別人，自己反而被淘汰了。
1COR|10|1|弟兄們，我不願意你們不知道，我們的祖宗從前都在雲下，都從海中經過，
1COR|10|2|都在雲裏、海裏受洗 歸了 摩西 ，
1COR|10|3|並且都吃了一樣的靈糧，
1COR|10|4|也都喝了一樣的靈水，所喝的是出於跟隨著他們的靈磐石；那磐石就是基督。
1COR|10|5|但他們中間多半是上帝不喜歡的人，所以倒斃在曠野裏了。
1COR|10|6|這些事都是我們的鑒戒，使我們不要貪戀惡事，像他們貪戀過的一樣。
1COR|10|7|也不要拜偶像，像他們中有些人曾經拜過。如經上所記：「百姓坐下吃喝，起來玩樂。」
1COR|10|8|我們也不可犯姦淫，像他們中有些人曾經犯過，一天就倒斃了二萬三千人。
1COR|10|9|也不可試探主 ，像他們中有些人曾試探主就被蛇咬死。
1COR|10|10|你們也不可發怨言，像他們中有些人曾經發過，就被毀滅者所滅。
1COR|10|11|這些事發生在他們身上，要作為鑒戒，而且寫下來正是要警戒我們這末世的人。
1COR|10|12|所以，自以為站得穩的人必須謹慎，免得跌倒。
1COR|10|13|你們所受的考驗無非是人所承受得了的。上帝是信實的，他不會讓你們遭受無法承受的考驗，在受考驗的時候，總會給你們開一條出路，讓你們能忍受得了。
1COR|10|14|所以，我親愛的，你們要遠避拜偶像的事。
1COR|10|15|我好像對精明人說的；你們要辨別我的話。
1COR|10|16|我們所祝謝的杯，豈不是同領基督的血嗎？我們所擘開的餅，豈不是同領基督的身體嗎？
1COR|10|17|因為餅只是一個，我們雖然人多，仍是一體，我們同享一個餅。
1COR|10|18|你們看那按肉體是 以色列 人的，那些吃祭物的人豈不是與祭壇有份嗎？
1COR|10|19|那麼，我怎麼說呢？是說祭偶像之物算得了甚麼嗎？或說偶像算得了甚麼嗎？
1COR|10|20|不，我是說，他們 所獻的祭是祭鬼，不是祭上帝；我不願意你們與鬼來往。
1COR|10|21|你們不能喝主的杯，又喝鬼的杯；不能吃主的筵席，又吃鬼的筵席。
1COR|10|22|我們要惹主的嫉恨嗎？我們比他更強嗎？
1COR|10|23|「凡事都可行」，但不都有益處。「凡事都可行」，但不都造就人。
1COR|10|24|無論甚麼人，不要求自己的益處，而要求別人的益處。
1COR|10|25|凡市場上所賣的，你們只管吃，不要為良心的緣故問甚麼，
1COR|10|26|「因為地和其中所充滿的都屬於主」。
1COR|10|27|倘若有一個不信的人請你們吃飯，而你們也願意去，凡擺在你們面前的，只管吃，不要為良心的緣故問甚麼。
1COR|10|28|若有人對你們說：「這是獻過祭的物」，那麼為了那告訴你們的人，並為了良心的緣故就不吃。
1COR|10|29|我說的良心不是你自己的，而是他的。我的自由為甚麼被別人的良心評斷呢？
1COR|10|30|我若謝恩而吃，為甚麼因我謝恩的物被人毀謗呢？
1COR|10|31|所以，你們或吃或喝，無論做甚麼，都要為榮耀上帝而做。
1COR|10|32|你們不要使 猶太 人、 希臘 人，或上帝教會中的人跌倒；
1COR|10|33|但要像我一樣，凡事都使眾人喜歡，不求自己的益處，只求眾人的益處，使他們得救。
1COR|11|1|你們該效法我，像我效法基督一樣。
1COR|11|2|我稱讚你們，因為你們凡事記得我，又堅守我所傳授給你們的。
1COR|11|3|但是我要你們知道：基督是男人的頭；男人是女人的頭 ；上帝是基督的頭。
1COR|11|4|凡男人禱告或講道 ，若蒙著頭，就是羞辱自己的頭。
1COR|11|5|凡女人禱告或講道，若不蒙著頭，就是羞辱自己的頭，因為這就如同剃了頭髮一樣。
1COR|11|6|女人若不蒙著頭，就該剪了頭髮；女人若以剪髮剃髮為羞愧，就該蒙著頭。
1COR|11|7|男人本不該蒙著頭，因為他是上帝的形像和榮耀；但女人是男人的榮耀。
1COR|11|8|起初，男人不是由女人而出，女人卻是由男人而出。
1COR|11|9|而且男人不是為女人造的，女人卻是為男人造的。
1COR|11|10|因此，女人為天使的緣故應當在頭上有服權柄的記號。
1COR|11|11|然而，照主的安排，女人不可沒有男人，男人也不可沒有女人。
1COR|11|12|因為女人原是由男人而出，男人是藉著女人而生；但萬有都是出於上帝。
1COR|11|13|你們自己要判斷，女人禱告上帝，不蒙著頭合宜嗎？
1COR|11|14|你們的本性不也教導你們，男人若留長頭髮是他的羞辱嗎？
1COR|11|15|但女人留長頭髮是她的榮耀，因為這頭髮是給她蓋頭的 。
1COR|11|16|若有人想要辯駁，我們卻沒有這樣的規矩，上帝的眾教會也沒有。
1COR|11|17|我現在吩咐你們這話不是在稱讚你們，因為你們聚會是有損無益的。
1COR|11|18|首先，我聽說你們教會聚會的時候有分裂的事，我也有些相信這話。
1COR|11|19|在你們中間必然有分門結黨的事，好使那些經得起考驗的人顯明出來。
1COR|11|20|你們聚會的時候，不是在吃主的晚餐，
1COR|11|21|因為吃的時候，各人先吃自己的飯，甚至有人飢餓，有人酒醉。
1COR|11|22|難道你們沒有家可以吃喝嗎？還是你們藐視上帝的教會，使那沒有的羞愧呢？我該對你們說甚麼呢？我要稱讚你們嗎？在這事上我絕不稱讚你們！
1COR|11|23|我當日傳給你們的是從主所領受的。主耶穌被出賣的那一夜，拿起餅來，
1COR|11|24|祝謝了，就擘開，說：「這是我的身體，為你們捨 的；你們要如此行，為的是記念我。」
1COR|11|25|飯後，他也照樣拿起杯來，說：「這杯是用我的血所立的新約；你們每逢喝的時候，要如此行，來記念我。」
1COR|11|26|你們每逢吃這餅，喝這杯，是宣告主的死，直到他來。
1COR|11|27|所以，任何不按規矩吃了主的餅，喝了主的杯，就是干犯主的身體和主的血了。
1COR|11|28|人應該省察自己，然後吃這餅，喝這杯。
1COR|11|29|因為人吃喝，若不分辨是主的身體，他的吃喝就是定自己的罪了。
1COR|11|30|因此，在你們中間有好些軟弱的與患病的，長眠了的也不少。
1COR|11|31|我們若是先省察自己，就不至於受審判。
1COR|11|32|我們受審判的時候，就是被主管教，這樣就免得和世人一同被定罪。
1COR|11|33|所以，我的弟兄們，你們聚會吃晚餐的時候，要彼此等待。
1COR|11|34|若有人餓了，要在家裏先吃，免得你們聚會，反被定罪。其餘的事等我來的時候再安排。
1COR|12|1|弟兄們，關於屬靈的恩賜 ，我不願意你們不明白。
1COR|12|2|你們知道，你們作外邦人的時候，隨事被引誘，受了迷惑去拜不會出聲的偶像。
1COR|12|3|所以，我要你們知道，被上帝的靈感動的，沒有人會說「耶穌該受詛咒」；若不是被聖靈感動的，也沒有人能說「耶穌是主」。
1COR|12|4|恩賜有許多種，卻是同一位聖靈所賜。
1COR|12|5|事奉有許多種，卻是事奉同一位主。
1COR|12|6|工作有許多種，卻是同一位上帝在萬人中運行萬事。
1COR|12|7|聖靈彰顯在各人身上，是要使人得益處。
1COR|12|8|有人藉著聖靈領受智慧的言語；有人也靠著同一位聖靈領受知識的言語；
1COR|12|9|又有人由同一位聖靈領受信心；還有人由同一位聖靈領受醫病的恩賜；
1COR|12|10|又有人能行異能，又有人能作先知，又有人能辨別諸靈，又有人能說方言 ，又有人能翻方言。
1COR|12|11|這一切都是由惟一的、同一位聖靈所運行，隨著自己的旨意分給各人的。
1COR|12|12|就如身體是一個，卻有許多肢體，身體的肢體雖多，仍是一個身體；基督也是這樣。
1COR|12|13|我們無論是 猶太 人是 希臘 人，是為奴的是自主的，都從一位聖靈受洗成了一個身體，並且共享這位聖靈。
1COR|12|14|身體原不只是一個肢體，而是許多肢體。
1COR|12|15|假如腳說：「我不是手，所以不屬於身體」，它不能因此就不屬於身體。
1COR|12|16|假如耳朵說：「我不是眼睛，所以不屬於身體」，它也不能因此就不屬於身體。
1COR|12|17|假如全身是眼睛，聽覺在哪裏呢？假如全身是耳朵，嗅覺在哪裏呢？
1COR|12|18|但現在上帝隨自己的意思把肢體一一安置在身體上了。
1COR|12|19|假如全都是一個肢體，身體在哪裏呢？
1COR|12|20|但現在肢體雖多，身體還是一個。
1COR|12|21|眼睛不能對手說：「我用不著你。」頭也不能對腳說：「我用不著你。」
1COR|12|22|不但如此，身上的肢體，人以為軟弱的，更是不可缺少的；
1COR|12|23|身上的肢體，我們認為不體面的，越發給它加上體面；我們不雅觀的，越發裝飾得雅觀。
1COR|12|24|我們雅觀的肢體自然用不著裝飾；但上帝配搭這身子，把加倍的體面給那有缺欠的肢體，
1COR|12|25|免得身體不協調，總要肢體彼此照顧。
1COR|12|26|假如一個肢體受苦，所有的肢體就一同受苦；假如一個肢體得光榮，所有的肢體就一同快樂。
1COR|12|27|你們是基督的身體，並且各自都是肢體。
1COR|12|28|上帝在教會所設立的：第一是使徒；第二是先知；第三是教師；其次是行異能的；再次是醫病的恩賜，幫助人的，治理事的，說方言的。
1COR|12|29|難道個個都是使徒嗎？難道個個都是先知嗎？難道個個都是教師嗎？難道個個都是行異能的嗎？
1COR|12|30|難道個個都是有醫病的恩賜嗎？難道個個都是說方言的嗎？難道個個都是翻方言的嗎？
1COR|12|31|你們要追求那更大的恩賜。 我現今把最妙的道指示你們。
1COR|13|1|我若能說人間的方言，甚至天使的語言，卻沒有愛，我就成為鳴的鑼、響的鈸一般。
1COR|13|2|我若有先知講道的能力，也明白各樣的奧祕，各樣的知識，而且有齊備的信心，使我能夠移山，卻沒有愛，我就算不了甚麼。
1COR|13|3|我若將所有的財產救濟窮人，又犧牲自己的身體讓人誇讚 ，卻沒有愛，仍然對我無益。
1COR|13|4|愛是恆久忍耐；又有恩慈；愛是不嫉妒；愛是不自誇，不張狂，
1COR|13|5|不做害羞的事，不求自己的益處，不輕易發怒，不計算人的惡，
1COR|13|6|不喜歡不義，只喜歡真理；
1COR|13|7|凡事包容，凡事相信，凡事盼望，凡事忍耐。
1COR|13|8|愛是永不止息。先知講道之能終必歸於無有；說方言 之能終必停止；知識也終必歸於無有。
1COR|13|9|我們現在所知道的有限，先知所講的也有限，
1COR|13|10|等那完全的來到，這有限的必消逝。
1COR|13|11|我作孩子的時候，說話像孩子，心思像孩子，意念像孩子；既長大成人，就把孩子的事丟棄了。
1COR|13|12|我們現在是對著鏡子觀看，模糊不清 ；到那時，就要面對面了。我如今所認識的有限，到那時就全認識，如同主認識我一樣。
1COR|13|13|如今常存的有信，有望，有愛這三樣，其中最大的是愛。
1COR|14|1|你們要追求愛，也要切慕屬靈的恩賜，尤其是作先知講道 。
1COR|14|2|那說方言 的，不是對人說，而是對上帝說，因為沒有人聽得懂；他是藉著聖靈說各樣的奧祕。
1COR|14|3|但作先知講道的，是對人說，要造就、安慰、勸勉人。
1COR|14|4|說方言的，是造就自己；作先知講道的，是造就教會。
1COR|14|5|我希望你們都說方言，更希望你們作先知講道；因為說方言的，若不解釋出來，使教會得造就，那作先知講道的就比他強了。
1COR|14|6|弟兄們，我到你們那裏去，若只說方言，不用啟示，或知識，或預言，或教導，給你們講解，我對你們有甚麼益處呢？
1COR|14|7|就連那有聲而沒有生命的東西，如簫，如琴，發出來的音若沒有分別，怎能知道所吹所彈的是甚麼呢？
1COR|14|8|號角吹出來的音若不清楚，誰會預備打仗呢？
1COR|14|9|你們也是如此；若用舌頭說聽不懂的信息，怎能知道所說的是甚麼呢？你們就是向空氣說話了。
1COR|14|10|世上有許多種語言，卻沒有一樣是無意思的。
1COR|14|11|我若不明白那語言的意思，說話的人必以我為未開化的人，我也以他為未開化的人。
1COR|14|12|你們也是如此，既然你們切慕屬靈的恩賜，就當追求多得造就教會的恩賜。
1COR|14|13|所以，那說方言的，就當祈求有翻方言的恩賜。
1COR|14|14|我若用方言禱告，是我的靈在禱告；但我的理智沒有效果。
1COR|14|15|我應該怎麼做呢？我要用靈禱告，也要用理智禱告；我要用靈歌唱，也要用理智歌唱。
1COR|14|16|不然，你用靈祝謝，那在座不通方言的人，既然不明白你的話，怎能在你感謝的時候說「阿們」呢？
1COR|14|17|你的感謝固然是好，不過不能造就別人。
1COR|14|18|我感謝上帝，我說方言比你們眾人還多；
1COR|14|19|但在教會中，我寧可用理智說五句教導人的話，強過說萬句方言。
1COR|14|20|弟兄們，在心志上不要作小孩子。但是，在惡事上要作嬰孩，而在心志上總要作大人。
1COR|14|21|律法上記著：「主說： 我要用外邦人的舌頭 和外邦人的嘴唇 向這百姓說話； 雖然如此，他們還是不聽從我。」
1COR|14|22|這樣看來，說方言不是為信的人作標記，而是為不信的人；作先知講道不是為不信的人作標記，而是為信的人。
1COR|14|23|所以，全教會聚在一處的時候，若都說方言，偶然有不通方言的或是不信的人進來，豈不會說你們瘋了嗎？
1COR|14|24|若個個都作先知講道，偶然有不信的或是不懂方言的人進來，就被眾人勸戒，被眾人審問，
1COR|14|25|他心裏的隱情被顯露出來，就必將臉伏地，敬拜上帝，宣告說：「上帝真的是在你們中間了。」
1COR|14|26|弟兄們，那麼，你們該怎麼做呢？你們聚會的時候，各人或有詩歌，或有教導，或有啟示，或有方言，或有翻出來，凡事都應當造就人。
1COR|14|27|若有說方言的，只可有兩個人，至多三個人，且要輪流著說，也要有一個人翻出來。
1COR|14|28|若沒有人翻，就當在會中閉口，只對自己和上帝說就是了。
1COR|14|29|至於作先知講道的，只可有兩個人或是三個人，其餘的人當慎思明辨。
1COR|14|30|假如旁邊坐著的得了啟示，那先說話的就當閉口不言。
1COR|14|31|因為你們都可以一個一個地作先知講道，使眾人都可以學習，使眾人都得勸勉。
1COR|14|32|先知的靈是順服先知的，
1COR|14|33|因為上帝不是叫人混亂，而是叫人和諧的上帝。 在聖徒的眾教會中，
1COR|14|34|婦女應該閉口不言；因為，不准她們說話，總要順服，正如律法所說的。
1COR|14|35|她們若要學甚麼，應該在家裏問自己的丈夫，因為婦女在會中說話是可恥的。
1COR|14|36|難道上帝的話是從你們出來的嗎？難道是單臨到你們的嗎？
1COR|14|37|若有人自以為是先知，或是屬靈的，就應該知道，我所寫給你們的是主的命令。
1COR|14|38|若有不理會的，你們也不必理會他。
1COR|14|39|所以，我的弟兄們，你們要切慕作先知講道的恩賜，不要禁止說方言。
1COR|14|40|凡事都要規規矩矩地按著次序行。
1COR|15|1|弟兄們，我要你們認清我先前傳給你們的福音；這福音你們領受了，又靠著它站立得住，
1COR|15|2|你們若能夠持守我傳給你們的信息，就必因這福音得救，否則你們是徒然相信。
1COR|15|3|我當日所領受又傳給你們的，最重要的就是：照聖經所說，基督為我們的罪死了，
1COR|15|4|而且埋葬了；又照聖經所說，第三天復活了，
1COR|15|5|還顯給 磯法 看，又顯給十二使徒看，
1COR|15|6|後來一次顯給五百多弟兄看，其中一大半到現在還在，卻也有已經睡了的。
1COR|15|7|以後他顯給 雅各 看，再顯給眾使徒看，
1COR|15|8|最後也顯給我看；我如同未到產期而生的人一般。
1COR|15|9|我原是使徒中最小的，不配稱為使徒，因為我曾迫害過上帝的教會。
1COR|15|10|然而，由於上帝的恩典，我才成了今日的我，並且他所賜給我的恩典不是徒然的。我比眾使徒格外勞苦；其實不是我，而是上帝的恩典與我同在。
1COR|15|11|無論是我或是其他使徒，我們都如此傳，你們也都如此信了。
1COR|15|12|既然我們傳基督是從死人中復活了，怎麼在你們中間有人說沒有死人復活的事呢？
1COR|15|13|若沒有死人復活的事，基督就沒有復活了。
1COR|15|14|基督若沒有復活，我們所傳的就是枉然，你們所信的也是枉然。
1COR|15|15|這樣，我們甚至被當作是為上帝妄作見證的，因為我們見證上帝是使基督復活了。如果死人真的沒有復活，上帝就沒有使基督復活了。
1COR|15|16|因為死人若不復活，基督也就沒有復活了。
1COR|15|17|基督若沒有復活，你們的信就是徒然，你們仍活在罪裏。
1COR|15|18|就是在基督裏睡了的人也滅亡了。
1COR|15|19|我們若靠基督只在今生有指望，就比所有的人更可憐了。
1COR|15|20|其實，基督已經從死人中復活，成為睡了之人初熟的果子。
1COR|15|21|既然死是因一人而來，死人復活也因一人而來。
1COR|15|22|在 亞當 裏眾人都死了；同樣，在基督裏眾人也都要復活。
1COR|15|23|但各人是按著自己的次序復活：初熟的果子是基督；然後在他來的時候，是那些屬於基督的。
1COR|15|24|再後，終結到了，那時基督既將一切執政的、掌權的、有權能的都毀滅了，就把國交給父上帝。
1COR|15|25|因為基督必須掌權，等上帝把一切仇敵都放在他的腳下。
1COR|15|26|他要毀滅的最後仇敵就是死亡。
1COR|15|27|因為經上說：「上帝使萬物都服在他的腳下。」既然說萬物都服了他，那使萬物屈服的，很明顯地是不在其內了。
1COR|15|28|既然萬物服了他，那時，子也要自己順服那叫萬物服他的，好使上帝在萬物之中，在萬物之上。
1COR|15|29|不然，那些為死人受洗的，能做甚麼呢？如果死人不會復活，為甚麼替他們受洗呢？
1COR|15|30|我們為甚麼要時刻冒險呢？
1COR|15|31|弟兄們 ，我在我們的主基督耶穌裏，指著你們—我所誇的極力地說，我天天冒死。
1COR|15|32|從人的觀點看來，我當日在 以弗所 同野獸搏鬥，對我有甚麼益處呢？如果死人沒有復活， 「讓我們吃吃喝喝吧！ 因為明天要死了。」
1COR|15|33|不要被欺騙了； 「濫交朋友敗壞品德。」
1COR|15|34|你們要醒悟為善，不再犯罪；因為有人不認識上帝。我說這話是要使你們羞愧。
1COR|15|35|但是有人會問：「死人怎樣復活呢？他們帶著甚麼身體來呢？」
1COR|15|36|無知的人哪，你所種的若不死就不能生。
1COR|15|37|並且你所種的不是那將來要有的形體，無論是麥子或別樣穀物，都不過是子粒。
1COR|15|38|但上帝隨自己的意思給它一個形體，並叫各樣子粒各有自己的形體。
1COR|15|39|不是所有的肉體都是同樣的：人是一個樣子，獸又是一個樣子，鳥又是一個樣子，魚又是一個樣子。
1COR|15|40|有天上的形體，也有地上的形體；但天上形體的榮光是一個樣子，地上形體的榮光又是一個樣子。
1COR|15|41|日有日的光輝，月有月的光輝，星有星的光輝；這星和那星的光輝也有區別。
1COR|15|42|死人復活也是這樣。所種的是會朽壞的，復活的是不朽壞的；
1COR|15|43|所種的是羞辱的，復活的是榮耀的；所種的是軟弱的，復活的是強壯的；
1COR|15|44|所種的是血肉的身體，復活的是靈性的身體。既有血肉的身體，也就有靈性的身體。
1COR|15|45|經上也是這樣記著說：「首先的人 亞當 成了有生命的人」；末後的 亞當 成了賜生命的靈。
1COR|15|46|但是，不是屬靈的在先，而是屬血肉的在先，然後才是屬靈的。
1COR|15|47|第一個人是出於地，是屬於塵土；第二個人是出於天。
1COR|15|48|那屬塵土的怎樣，凡屬塵土的也都怎樣；屬天的怎樣，凡屬天的也都怎樣。
1COR|15|49|就如我們既有屬塵土的形像，將來也必有屬天的形像。
1COR|15|50|弟兄們，我要告訴你們的是：血肉之軀不能承受上帝的國，必朽壞的也不能承受不朽壞的。
1COR|15|51|我如今把一件奧祕的事告訴你們：我們不是都要睡覺，而是都要改變，
1COR|15|52|就在一剎那，眨眼之間，號筒末次吹響的時候。因號筒要吹響，死人要復活成為不朽壞的，我們也要改變。
1COR|15|53|這會朽壞的必須變成 不朽壞的；這會死的總要變成不會死的。
1COR|15|54|當這會朽壞的變成不朽壞的，這會死的變成不會死的，那時經上所記「死亡已被勝利吞滅了」的話就應驗了。
1COR|15|55|「死亡啊！你得勝的權勢在哪裏？ 死亡啊！你的毒刺在哪裏？」
1COR|15|56|死亡的毒刺就是罪，罪的權勢就是律法。
1COR|15|57|感謝上帝，他使我們藉著我們的主耶穌基督得勝。
1COR|15|58|所以，我親愛的弟兄們，你們務要堅固，不可動搖，常常竭力多做主工，因為你們知道，你們在主裏的勞苦不是徒然的。
1COR|16|1|關於為聖徒捐款的事，我從前怎樣吩咐 加拉太 的眾教會，你們也該怎樣做。
1COR|16|2|每逢七日的第一日，每人要照自己的收入抽出若干，保留起來，免得我來的時候現湊。
1COR|16|3|等到我來了，你們寫信舉薦誰，我就差遣他們，把你們的款項送到 耶路撒冷 去。
1COR|16|4|如果我也該去，他們可以和我同去。
1COR|16|5|我想穿越 馬其頓 ；我經過了 馬其頓 後，就到你們那裏去，
1COR|16|6|可能會和你們同住一些時候，甚至和你們一起過冬。這樣無論我往哪裏去，你們可以給我送行。
1COR|16|7|我現在不願意在路過的時候見你們；主若允許，我就指望和你們同住一些時候。
1COR|16|8|不過我要仍舊住在 以弗所 ，直到五旬節，
1COR|16|9|因為有又寬大又有效的門為我開了，雖然反對的人也多。
1COR|16|10|若是 提摩太 來到，你們要留心照顧他，使他在你們那裏無所懼怕，因為他做主的工作像我一樣。
1COR|16|11|所以，無論誰都不可藐視他。只要送他平安前行，讓他到我這裏來，因為我等著他和弟兄們同來。
1COR|16|12|至於 亞波羅 弟兄，我再三勸他同弟兄們到你們那裏去；但現在他絕不願意去，等有機會他就會去。
1COR|16|13|你們要警醒，在信仰上要站穩，要勇敢，要剛強。
1COR|16|14|你們所做的一切都要憑愛心而做。
1COR|16|15|弟兄們，你們知道 司提法那 一家，是 亞該亞 初結的果子；他們專以服事聖徒為念。
1COR|16|16|我勸你們順服這樣的人，和一切與他同工同勞的人。
1COR|16|17|司提法那 、 福徒拿都 和 亞該古 到這裏來，我很高興，因為他們補上了你們不在我身邊的遺憾。
1COR|16|18|他們使我和你們心裏都快慰；這樣的人，你們務要敬重。
1COR|16|19|亞細亞 的眾教會向你們問安。 亞居拉 、 百基拉 ，和在他們家裏的教會，在主裏熱切地向你們問安。
1COR|16|20|眾弟兄都向你們問安。要用聖潔的吻彼此問安。
1COR|16|21|我— 保羅 親筆問安。
1COR|16|22|若有人不愛主，這人該受詛咒。主啊，願你來！
1COR|16|23|願主耶穌基督的恩常與你們眾人同在。
1COR|16|24|我在基督耶穌裏的愛與你們同在！
