JOB|1|1|There was a man in the land of Uz whose name was Job, and that man was blameless and upright, one who feared God and turned away from evil.
JOB|1|2|There were born to him seven sons and three daughters.
JOB|1|3|He possessed 7,000 sheep, 3,000 camels, 500 yoke of oxen, and 500 female donkeys, and very many servants, so that this man was the greatest of all the people of the east.
JOB|1|4|His sons used to go and hold a feast in the house of each one on his day, and they would send and invite their three sisters to eat and drink with them.
JOB|1|5|And when the days of the feast had run their course, Job would send and consecrate them, and he would rise early in the morning and offer burnt offerings according to the number of them all. For Job said, "It may be that my children have sinned, and cursed God in their hearts." Thus Job did continually.
JOB|1|6|Now there was a day when the sons of God came to present themselves before the LORD, and Satan also came among them.
JOB|1|7|The LORD said to Satan, "From where have you come?" Satan answered the LORD and said, "From going to and fro on the earth, and from walking up and down on it."
JOB|1|8|And the LORD said to Satan, "Have you considered my servant Job, that there is none like him on the earth, a blameless and upright man, who fears God and turns away from evil?"
JOB|1|9|Then Satan answered the LORD and said, "Does Job fear God for no reason?
JOB|1|10|Have you not put a hedge around him and his house and all that he has, on every side? You have blessed the work of his hands, and his possessions have increased in the land.
JOB|1|11|But stretch out your hand and touch all that he has, and he will curse you to your face."
JOB|1|12|And the LORD said to Satan, "Behold, all that he has is in your hand. Only against him do not stretch out your hand." So Satan went out from the presence of the LORD.
JOB|1|13|Now there was a day when his sons and daughters were eating and drinking wine in their oldest brother's house,
JOB|1|14|and there came a messenger to Job and said, "The oxen were plowing and the donkeys feeding beside them,
JOB|1|15|and the Sabeans fell upon them and took them and struck down the servants with the edge of the sword, and I alone have escaped to tell you."
JOB|1|16|While he was yet speaking, there came another and said, "The fire of God fell from heaven and burned up the sheep and the servants and consumed them, and I alone have escaped to tell you."
JOB|1|17|While he was yet speaking, there came another and said, "The Chaldeans formed three groups and made a raid on the camels and took them and struck down the servants with the edge of the sword, and I alone have escaped to tell you."
JOB|1|18|While he was yet speaking, there came another and said, "Your sons and daughters were eating and drinking wine in their oldest brother's house,
JOB|1|19|and behold, a great wind came across the wilderness and struck the four corners of the house, and it fell upon the young people, and they are dead, and I alone have escaped to tell you."
JOB|1|20|Then Job arose and tore his robe and shaved his head and fell on the ground and worshiped.
JOB|1|21|And he said, "Naked I came from my mother's womb, and naked shall I return. The LORD gave, and the LORD has taken away; blessed be the name of the LORD."
JOB|1|22|In all this Job did not sin or charge God with wrong.
JOB|2|1|Again there was a day when the sons of God came to present themselves before the LORD, and Satan also came among them to present himself before the LORD.
JOB|2|2|And the LORD said to Satan, "From where have you come?" Satan answered the LORD and said, "From going to and fro on the earth, and from walking up and down on it."
JOB|2|3|And the LORD said to Satan, "Have you considered my servant Job, that there is none like him on the earth, a blameless and upright man, who fears God and turns away from evil? He still holds fast his integrity, although you incited me against him to destroy him without reason."
JOB|2|4|Then Satan answered the LORD and said, "Skin for skin! All that a man has he will give for his life.
JOB|2|5|But stretch out your hand and touch his bone and his flesh, and he will curse you to your face."
JOB|2|6|And the LORD said to Satan, "Behold, he is in your hand; only spare his life."
JOB|2|7|So Satan went out from the presence of the LORD and struck Job with loathsome sores from the sole of his foot to the crown of his head.
JOB|2|8|And he took a piece of broken pottery with which to scrape himself while he sat in the ashes.
JOB|2|9|Then his wife said to him, "Do you still hold fast your integrity? Curse God and die."
JOB|2|10|But he said to her, "You speak as one of the foolish women would speak. Shall we receive good from God, and shall we not receive evil?" In all this Job did not sin with his lips.
JOB|2|11|Now when Job's three friends heard of all this evil that had come upon him, they came each from his own place, Eliphaz the Temanite, Bildad the Shuhite, and Zophar the Naamathite. They made an appointment together to come to show him sympathy and comfort him.
JOB|2|12|And when they saw him from a distance, they did not recognize him. And they raised their voices and wept, and they tore their robes and sprinkled dust on their heads toward heaven.
JOB|2|13|And they sat with him on the ground seven days and seven nights, and no one spoke a word to him, for they saw that his suffering was very great.
JOB|3|1|After this Job opened his mouth and cursed the day of his birth.
JOB|3|2|And Job said:
JOB|3|3|"Let the day perish on which I was born, and the night that said, 'A man is conceived.'
JOB|3|4|Let that day be darkness! May God above not seek it, nor light shine upon it.
JOB|3|5|Let gloom and deep darkness claim it. Let clouds dwell upon it; let the blackness of the day terrify it.
JOB|3|6|That night- let thick darkness seize it! Let it not rejoice among the days of the year; let it not come into the number of the months.
JOB|3|7|Behold, let that night be barren; let no joyful cry enter it.
JOB|3|8|Let those curse it who curse the day, who are ready to rouse up Leviathan.
JOB|3|9|Let the stars of its dawn be dark; let it hope for light, but have none, nor see the eyelids of the morning,
JOB|3|10|because it did not shut the doors of my mother's womb, nor hide trouble from my eyes.
JOB|3|11|"Why did I not die at birth, come out from the womb and expire?
JOB|3|12|Why did the knees receive me? Or why the breasts, that I should nurse?
JOB|3|13|For then I would have lain down and been quiet; I would have slept; then I would have been at rest,
JOB|3|14|with kings and counselors of the earth who rebuilt ruins for themselves,
JOB|3|15|or with princes who had gold, who filled their houses with silver.
JOB|3|16|Or why was I not as a hidden stillborn child, as infants who never see the light?
JOB|3|17|There the wicked cease from troubling, and there the weary are at rest.
JOB|3|18|There the prisoners are at ease together; they hear not the voice of the taskmaster.
JOB|3|19|The small and the great are there, and the slave is free from his master.
JOB|3|20|"Why is light given to him who is in misery, and life to the bitter in soul,
JOB|3|21|who long for death, but it comes not, and dig for it more than for hidden treasures,
JOB|3|22|who rejoice exceedingly and are glad when they find the grave?
JOB|3|23|Why is light given to a man whose way is hidden, whom God has hedged in?
JOB|3|24|For my sighing comes instead of my bread, and my groanings are poured out like water.
JOB|3|25|For the thing that I fear comes upon me, and what I dread befalls me.
JOB|3|26|I am not at ease, nor am I quiet; I have no rest, but trouble comes."
JOB|4|1|Then Eliphaz the Temanite answered and said:
JOB|4|2|"If one ventures a word with you, will you be impatient? Yet who can keep from speaking?
JOB|4|3|Behold, you have instructed many, and you have strengthened the weak hands.
JOB|4|4|Your words have upheld him who was stumbling, and you have made firm the feeble knees.
JOB|4|5|But now it has come to you, and you are impatient; it touches you, and you are dismayed.
JOB|4|6|Is not your fear of God your confidence, and the integrity of your ways your hope?
JOB|4|7|"Remember: who that was innocent ever perished? Or where were the upright cut off?
JOB|4|8|As I have seen, those who plow iniquity and sow trouble reap the same.
JOB|4|9|By the breath of God they perish, and by the blast of his anger they are consumed.
JOB|4|10|The roar of the lion, the voice of the fierce lion, the teeth of the young lions are broken.
JOB|4|11|The strong lion perishes for lack of prey, and the cubs of the lioness are scattered.
JOB|4|12|"Now a word was brought to me stealthily; my ear received the whisper of it.
JOB|4|13|Amid thoughts from visions of the night, when deep sleep falls on men,
JOB|4|14|dread came upon me, and trembling, which made all my bones shake.
JOB|4|15|A spirit glided past my face; the hair of my flesh stood up.
JOB|4|16|It stood still, but I could not discern its appearance. A form was before my eyes; there was silence, then I heard a voice:
JOB|4|17|'Can mortal man be in the right before God? Can a man be pure before his Maker?
JOB|4|18|Even in his servants he puts no trust, and his angels he charges with error;
JOB|4|19|how much more those who dwell in houses of clay, whose foundation is in the dust, who are crushed like the moth.
JOB|4|20|Between morning and evening they are beaten to pieces; they perish forever without anyone regarding it.
JOB|4|21|Is not their tent-cord plucked up within them, do they not die, and that without wisdom?'
JOB|5|1|"Call now; is there anyone who will answer you? To which of the holy ones will you turn?
JOB|5|2|Surely vexation kills the fool, and jealousy slays the simple.
JOB|5|3|I have seen the fool taking root, but suddenly I cursed his dwelling.
JOB|5|4|His children are far from safety; they are crushed in the gate, and there is no one to deliver them.
JOB|5|5|The hungry eat his harvest, and he takes it even out of thorns, and the thirsty pant after his wealth.
JOB|5|6|For affliction does not come from the dust, nor does trouble sprout from the ground,
JOB|5|7|but man is born to trouble as the sparks fly upward.
JOB|5|8|"As for me, I would seek God, and to God would I commit my cause,
JOB|5|9|who does great things and unsearchable, marvelous things without number:
JOB|5|10|he gives rain on the earth and sends waters on the fields;
JOB|5|11|he sets on high those who are lowly, and those who mourn are lifted to safety.
JOB|5|12|He frustrates the devices of the crafty, so that their hands achieve no success.
JOB|5|13|He catches the wise in their own craftiness, and the schemes of the wily are brought to a quick end.
JOB|5|14|They meet with darkness in the daytime and grope at noonday as in the night.
JOB|5|15|But he saves the needy from the sword of their mouth and from the hand of the mighty.
JOB|5|16|So the poor have hope, and injustice shuts her mouth.
JOB|5|17|"Behold, blessed is the one whom God reproves; therefore despise not the discipline of the Almighty.
JOB|5|18|For he wounds, but he binds up; he shatters, but his hands heal.
JOB|5|19|He will deliver you from six troubles; in seven no evil shall touch you.
JOB|5|20|In famine he will redeem you from death, and in war from the power of the sword.
JOB|5|21|You shall be hidden from the lash of the tongue, and shall not fear destruction when it comes.
JOB|5|22|At destruction and famine you shall laugh, and shall not fear the beasts of the earth.
JOB|5|23|For you shall be in league with the stones of the field, and the beasts of the field shall be at peace with you.
JOB|5|24|You shall know that your tent is at peace, and you shall inspect your fold and miss nothing.
JOB|5|25|You shall know also that your offspring shall be many, and your descendants as the grass of the earth.
JOB|5|26|You shall come to your grave in ripe old age, like a sheaf gathered up in its season.
JOB|5|27|Behold, this we have searched out; it is true. Hear, and know it for your good."
JOB|6|1|Then Job answered and said:
JOB|6|2|"Oh that my vexation were weighed, and all my calamity laid in the balances!
JOB|6|3|For then it would be heavier than the sand of the sea; therefore my words have been rash.
JOB|6|4|For the arrows of the Almighty are in me; my spirit drinks their poison; the terrors of God are arrayed against me.
JOB|6|5|Does the wild donkey bray when he has grass, or the ox low over his fodder?
JOB|6|6|Can that which is tasteless be eaten without salt, or is there any taste in the juice of the mallow?
JOB|6|7|My appetite refuses to touch them; they are as food that is loathsome to me.
JOB|6|8|"Oh that I might have my request, and that God would fulfill my hope,
JOB|6|9|that it would please God to crush me, that he would let loose his hand and cut me off!
JOB|6|10|This would be my comfort; I would even exult in pain unsparing, for I have not denied the words of the Holy One.
JOB|6|11|What is my strength, that I should wait? And what is my end, that I should be patient?
JOB|6|12|Is my strength the strength of stones, or is my flesh bronze?
JOB|6|13|Have I any help in me, when resource is driven from me?
JOB|6|14|"He who withholds kindness from a friend forsakes the fear of the Almighty.
JOB|6|15|My brothers are treacherous as a torrent-bed, as torrential streams that pass away,
JOB|6|16|which are dark with ice, and where the snow hides itself.
JOB|6|17|When they melt, they disappear; when it is hot, they vanish from their place.
JOB|6|18|The caravans turn aside from their course; they go up into the waste and perish.
JOB|6|19|The caravans of Tema look, the travelers of Sheba hope.
JOB|6|20|They are ashamed because they were confident; they come there and are disappointed.
JOB|6|21|For you have now become nothing; you see my calamity and are afraid.
JOB|6|22|Have I said, 'Make me a gift'? Or, 'From your wealth offer a bribe for me'?
JOB|6|23|Or, 'Deliver me from the adversary's hand'? Or, 'Redeem me from the hand of the ruthless'?
JOB|6|24|"Teach me, and I will be silent; make me understand how I have gone astray.
JOB|6|25|How forceful are upright words! But what does reproof from you reprove?
JOB|6|26|Do you think that you can reprove words, when the speech of a despairing man is wind?
JOB|6|27|You would even cast lots over the fatherless, and bargain over your friend.
JOB|6|28|"But now, be pleased to look at me, for I will not lie to your face.
JOB|6|29|Please turn; let no injustice be done. Turn now; my vindication is at stake.
JOB|6|30|Is there any injustice on my tongue? Cannot my palate discern the cause of calamity?
JOB|7|1|"Has not man a hard service on earth, and are not his days like the days of a hired hand?
JOB|7|2|Like a slave who longs for the shadow, and like a hired hand who looks for his wages,
JOB|7|3|so I am allotted months of emptiness, and nights of misery are apportioned to me.
JOB|7|4|When I lie down I say, 'When shall I arise?' But the night is long, and I am full of tossing till the dawn.
JOB|7|5|My flesh is clothed with worms and dirt; my skin hardens, then breaks out afresh.
JOB|7|6|My days are swifter than a weaver's shuttle and come to their end without hope.
JOB|7|7|"Remember that my life is a breath; my eye will never again see good.
JOB|7|8|The eye of him who sees me will behold me no more; while your eyes are on me, I shall be gone.
JOB|7|9|As the cloud fades and vanishes, so he who goes down to Sheol does not come up;
JOB|7|10|he returns no more to his house, nor does his place know him anymore.
JOB|7|11|"Therefore I will not restrain my mouth; I will speak in the anguish of my spirit; I will complain in the bitterness of my soul.
JOB|7|12|Am I the sea, or a sea monster, that you set a guard over me?
JOB|7|13|When I say, 'My bed will comfort me, my couch will ease my complaint,'
JOB|7|14|then you scare me with dreams and terrify me with visions,
JOB|7|15|so that I would choose strangling and death rather than my bones.
JOB|7|16|I loathe my life; I would not live forever. Leave me alone, for my days are a breath.
JOB|7|17|What is man, that you make so much of him, and that you set your heart on him,
JOB|7|18|visit him every morning and test him every moment?
JOB|7|19|How long will you not look away from me, nor leave me alone till I swallow my spit?
JOB|7|20|If I sin, what do I do to you, you watcher of mankind? Why have you made me your mark? Why have I become a burden to you?
JOB|7|21|Why do you not pardon my transgression and take away my iniquity? For now I shall lie in the earth; you will seek me, but I shall not be."
JOB|8|1|Then Bildad the Shuhite answered and said:
JOB|8|2|"How long will you say these things, and the words of your mouth be a great wind?
JOB|8|3|Does God pervert justice? Or does the Almighty pervert the right?
JOB|8|4|If your children have sinned against him, he has delivered them into the hand of their transgression.
JOB|8|5|If you will seek God and plead with the Almighty for mercy,
JOB|8|6|if you are pure and upright, surely then he will rouse himself for you and restore your rightful habitation.
JOB|8|7|And though your beginning was small, your latter days will be very great.
JOB|8|8|"For inquire, please, of bygone ages, and consider what the fathers have searched out.
JOB|8|9|For we are but of yesterday and know nothing, for our days on earth are a shadow.
JOB|8|10|Will they not teach you and tell you and utter words out of their understanding?
JOB|8|11|"Can papyrus grow where there is no marsh? Can reeds flourish where there is no water?
JOB|8|12|While yet in flower and not cut down, they wither before any other plant.
JOB|8|13|Such are the paths of all who forget God; the hope of the godless shall perish.
JOB|8|14|His confidence is severed, and his trust is a spider's web.
JOB|8|15|He leans against his house, but it does not stand; he lays hold of it, but it does not endure.
JOB|8|16|He is a lush plant before the sun, and his shoots spread over his garden.
JOB|8|17|His roots entwine the stone heap; he looks upon a house of stones.
JOB|8|18|If he is destroyed from his place, then it will deny him, saying, 'I have never seen you.'
JOB|8|19|Behold, this is the joy of his way, and out of the soil others will spring.
JOB|8|20|"Behold, God will not reject a blameless man, nor take the hand of evildoers.
JOB|8|21|He will yet fill your mouth with laughter, and your lips with shouting.
JOB|8|22|Those who hate you will be clothed with shame, and the tent of the wicked will be no more."
JOB|9|1|Then Job answered and said:
JOB|9|2|"Truly I know that it is so: But how can a man be in the right before God?
JOB|9|3|If one wished to contend with him, one could not answer him once in a thousand times.
JOB|9|4|He is wise in heart and mighty in strength- who has hardened himself against him, and succeeded?-
JOB|9|5|he who removes mountains, and they know it not, when he overturns them in his anger,
JOB|9|6|who shakes the earth out of its place, and its pillars tremble;
JOB|9|7|who commands the sun, and it does not rise; who seals up the stars;
JOB|9|8|who alone stretched out the heavens and trampled the waves of the sea;
JOB|9|9|who made the Bear and Orion, the Pleiades and the chambers of the south;
JOB|9|10|who does great things beyond searching out, and marvelous things beyond number.
JOB|9|11|Behold, he passes by me, and I see him not; he moves on, but I do not perceive him.
JOB|9|12|Behold, he snatches away; who can turn him back? Who will say to him, 'What are you doing?'
JOB|9|13|"God will not turn back his anger; beneath him bowed the helpers of Rahab.
JOB|9|14|How then can I answer him, choosing my words with him?
JOB|9|15|Though I am in the right, I cannot answer him; I must appeal for mercy to my accuser.
JOB|9|16|If I summoned him and he answered me, I would not believe that he was listening to my voice.
JOB|9|17|For he crushes me with a tempest and multiplies my wounds without cause;
JOB|9|18|he will not let me get my breath, but fills me with bitterness.
JOB|9|19|If it is a contest of strength, behold, he is mighty! If it is a matter of justice, who can summon him?
JOB|9|20|Though I am in the right, my own mouth would condemn me; though I am blameless, he would prove me perverse.
JOB|9|21|I am blameless; I regard not myself; I loathe my life.
JOB|9|22|It is all one; therefore I say, He destroys both the blameless and the wicked.
JOB|9|23|When disaster brings sudden death, he mocks at the calamity of the innocent.
JOB|9|24|The earth is given into the hand of the wicked; he covers the faces of its judges- if it is not he, who then is it?
JOB|9|25|"My days are swifter than a runner; they flee away; they see no good.
JOB|9|26|They go by like skiffs of reed, like an eagle swooping on the prey.
JOB|9|27|If I say, 'I will forget my complaint, I will put off my sad face, and be of good cheer,'
JOB|9|28|I become afraid of all my suffering, for I know you will not hold me innocent.
JOB|9|29|I shall be condemned; why then do I labor in vain?
JOB|9|30|If I wash myself with snow and cleanse my hands with lye,
JOB|9|31|yet you will plunge me into a pit, and my own clothes will abhor me.
JOB|9|32|For he is not a man, as I am, that I might answer him, that we should come to trial together.
JOB|9|33|There is no arbiter between us, who might lay his hand on us both.
JOB|9|34|Let him take his rod away from me, and let not dread of him terrify me.
JOB|9|35|Then I would speak without fear of him, for I am not so in myself.
JOB|10|1|"I loathe my life; I will give free utterance to my complaint; I will speak in the bitterness of my soul.
JOB|10|2|I will say to God, Do not condemn me; let me know why you contend against me.
JOB|10|3|Does it seem good to you to oppress, to despise the work of your hands and favor the designs of the wicked?
JOB|10|4|Have you eyes of flesh? Do you see as man sees?
JOB|10|5|Are your days as the days of man, or your years as a man's years,
JOB|10|6|that you seek out my iniquity and search for my sin,
JOB|10|7|although you know that I am not guilty, and there is none to deliver out of your hand?
JOB|10|8|Your hands fashioned and made me, and now you have destroyed me altogether.
JOB|10|9|Remember that you have made me like clay; and will you return me to the dust?
JOB|10|10|Did you not pour me out like milk and curdle me like cheese?
JOB|10|11|You clothed me with skin and flesh, and knit me together with bones and sinews.
JOB|10|12|You have granted me life and steadfast love, and your care has preserved my spirit.
JOB|10|13|Yet these things you hid in your heart; I know that this was your purpose.
JOB|10|14|If I sin, you watch me and do not acquit me of my iniquity.
JOB|10|15|If I am guilty, woe to me! If I am in the right, I cannot lift up my head, for I am filled with disgrace and look on my affliction.
JOB|10|16|And were my head lifted up, you would hunt me like a lion and again work wonders against me.
JOB|10|17|You renew your witnesses against me and increase your vexation toward me; you bring fresh troops against me.
JOB|10|18|"Why did you bring me out from the womb? Would that I had died before any eye had seen me
JOB|10|19|and were as though I had not been, carried from the womb to the grave.
JOB|10|20|Are not my days few? Then cease, and leave me alone, that I may find a little cheer
JOB|10|21|before I go- and I shall not return- to the land of darkness and deep shadow,
JOB|10|22|the land of gloom like thick darkness, like deep shadow without any order, where light is as thick darkness."
JOB|11|1|Then Zophar the Naamathite answered and said:
JOB|11|2|"Should a multitude of words go unanswered, and a man full of talk be judged right?
JOB|11|3|Should your babble silence men, and when you mock, shall no one shame you?
JOB|11|4|For you say, 'My doctrine is pure, and I am clean in God's eyes.'
JOB|11|5|But oh, that God would speak and open his lips to you,
JOB|11|6|and that he would tell you the secrets of wisdom! For he is manifold in understanding. Know then that God exacts of you less than your guilt deserves.
JOB|11|7|"Can you find out the deep things of God? Can you find out the limit of the Almighty?
JOB|11|8|It is higher than heaven- what can you do? Deeper than Sheol- what can you know?
JOB|11|9|Its measure is longer than the earth and broader than the sea.
JOB|11|10|If he passes through and imprisons and summons the court, who can turn him back?
JOB|11|11|For he knows worthless men; when he sees iniquity, will he not consider it?
JOB|11|12|But a stupid man will get understanding when a wild donkey's colt is born a man!
JOB|11|13|"If you prepare your heart, you will stretch out your hands toward him.
JOB|11|14|If iniquity is in your hand, put it far away, and let not injustice dwell in your tents.
JOB|11|15|Surely then you will lift up your face without blemish; you will be secure and will not fear.
JOB|11|16|You will forget your misery; you will remember it as waters that have passed away.
JOB|11|17|And your life will be brighter than the noonday; its darkness will be like the morning.
JOB|11|18|And you will feel secure, because there is hope; you will look around and take your rest in security.
JOB|11|19|You will lie down, and none will make you afraid; many will court your favor.
JOB|11|20|But the eyes of the wicked will fail; all way of escape will be lost to them, and their hope is to breathe their last."
JOB|12|1|Then Job answered and said:
JOB|12|2|"No doubt you are the people, and wisdom will die with you.
JOB|12|3|But I have understanding as well as you; I am not inferior to you. Who does not know such things as these?
JOB|12|4|I am a laughingstock to my friends; I, who called to God and he answered me, a just and blameless man, am a laughingstock.
JOB|12|5|In the thought of one who is at ease there is contempt for misfortune; it is ready for those whose feet slip.
JOB|12|6|The tents of robbers are at peace, and those who provoke God are secure, who bring their god in their hand.
JOB|12|7|"But ask the beasts, and they will teach you; the birds of the heavens, and they will tell you;
JOB|12|8|or the bushes of the earth, and they will teach you; and the fish of the sea will declare to you.
JOB|12|9|Who among all these does not know that the hand of the LORD has done this?
JOB|12|10|In his hand is the life of every living thing and the breath of all mankind.
JOB|12|11|Does not the ear test words as the palate tastes food?
JOB|12|12|Wisdom is with the aged, and understanding in length of days.
JOB|12|13|"With God are wisdom and might; he has counsel and understanding.
JOB|12|14|If he tears down, none can rebuild; if he shuts a man in, none can open.
JOB|12|15|If he withholds the waters, they dry up; if he sends them out, they overwhelm the land.
JOB|12|16|With him are strength and sound wisdom; the deceived and the deceiver are his.
JOB|12|17|He leads counselors away stripped, and judges he makes fools.
JOB|12|18|He looses the bonds of kings and binds a waistcloth on their hips.
JOB|12|19|He leads priests away stripped and overthrows the mighty.
JOB|12|20|He deprives of speech those who are trusted and takes away the discernment of the elders.
JOB|12|21|He pours contempt on princes and loosens the belt of the strong.
JOB|12|22|He uncovers the deeps out of darkness and brings deep darkness to light.
JOB|12|23|He makes nations great, and he destroys them; he enlarges nations, and leads them away.
JOB|12|24|He takes away understanding from the chiefs of the people of the earth and makes them wander in a pathless waste.
JOB|12|25|They grope in the dark without light, and he makes them stagger like a drunken man.
JOB|13|1|"Behold, my eye has seen all this, my ear has heard and understood it.
JOB|13|2|What you know, I also know; I am not inferior to you.
JOB|13|3|But I would speak to the Almighty, and I desire to argue my case with God.
JOB|13|4|As for you, you whitewash with lies; worthless physicians are you all.
JOB|13|5|Oh that you would keep silent, and it would be your wisdom!
JOB|13|6|Hear now my argument and listen to the pleadings of my lips.
JOB|13|7|Will you speak falsely for God and speak deceitfully for him?
JOB|13|8|Will you show partiality toward him? Will you plead the case for God?
JOB|13|9|Will it be well with you when he searches you out? Or can you deceive him, as one deceives a man?
JOB|13|10|He will surely rebuke you if in secret you show partiality.
JOB|13|11|Will not his majesty terrify you, and the dread of him fall upon you?
JOB|13|12|Your maxims are proverbs of ashes; your defenses are defenses of clay.
JOB|13|13|"Let me have silence, and I will speak, and let come on me what may.
JOB|13|14|Why should I take my flesh in my teeth and put my life in my hand?
JOB|13|15|Though he slay me, I will hope in him; yet I will argue my ways to his face.
JOB|13|16|This will be my salvation, that the godless shall not come before him.
JOB|13|17|Keep listening to my words, and let my declaration be in your ears.
JOB|13|18|Behold, I have prepared my case; I know that I shall be in the right.
JOB|13|19|Who is there who will contend with me? For then I would be silent and die.
JOB|13|20|Only grant me two things, then I will not hide myself from your face:
JOB|13|21|withdraw your hand far from me, and let not dread of you terrify me.
JOB|13|22|Then call, and I will answer; or let me speak, and you reply to me.
JOB|13|23|How many are my iniquities and my sins? Make me know my transgression and my sin.
JOB|13|24|Why do you hide your face and count me as your enemy?
JOB|13|25|Will you frighten a driven leaf and pursue dry chaff?
JOB|13|26|For you write bitter things against me and make me inherit the iniquities of my youth.
JOB|13|27|You put my feet in the stocks and watch all my paths; you set a limit for the soles of my feet.
JOB|13|28|Man wastes away like a rotten thing, like a garment that is moth-eaten.
JOB|14|1|"Man who is born of a woman is few of days and full of trouble.
JOB|14|2|He comes out like a flower and withers; he flees like a shadow and continues not.
JOB|14|3|And do you open your eyes on such a one and bring me into judgment with you?
JOB|14|4|Who can bring a clean thing out of an unclean? There is not one.
JOB|14|5|Since his days are determined, and the number of his months is with you, and you have appointed his limits that he cannot pass,
JOB|14|6|look away from him and leave him alone, that he may enjoy, like a hired hand, his day.
JOB|14|7|"For there is hope for a tree, if it be cut down, that it will sprout again, and that its shoots will not cease.
JOB|14|8|Though its root grow old in the earth, and its stump die in the soil,
JOB|14|9|yet at the scent of water it will bud and put out branches like a young plant.
JOB|14|10|But a man dies and is laid low; man breathes his last, and where is he?
JOB|14|11|As waters fail from a lake and a river wastes away and dries up,
JOB|14|12|so a man lies down and rises not again; till the heavens are no more he will not awake or be roused out of his sleep.
JOB|14|13|Oh that you would hide me in Sheol, that you would conceal me until your wrath be past, that you would appoint me a set time, and remember me!
JOB|14|14|If a man dies, shall he live again? All the days of my service I would wait, till my renewal should come.
JOB|14|15|You would call, and I would answer you; you would long for the work of your hands.
JOB|14|16|For then you would number my steps; you would not keep watch over my sin;
JOB|14|17|my transgression would be sealed up in a bag, and you would cover over my iniquity.
JOB|14|18|"But the mountain falls and crumbles away, and the rock is removed from its place;
JOB|14|19|the waters wear away the stones; the torrents wash away the soil of the earth; so you destroy the hope of man.
JOB|14|20|You prevail forever against him, and he passes; you change his countenance, and send him away.
JOB|14|21|His sons come to honor, and he does not know it; they are brought low, and he perceives it not.
JOB|14|22|He feels only the pain of his own body, and he mourns only for himself."
JOB|15|1|Then Eliphaz the Temanite answered and said:
JOB|15|2|"Should a wise man answer with windy knowledge, and fill his belly with the east wind?
JOB|15|3|Should he argue in unprofitable talk, or in words with which he can do no good?
JOB|15|4|But you are doing away with the fear of God and hindering meditation before God.
JOB|15|5|For your iniquity teaches your mouth, and you choose the tongue of the crafty.
JOB|15|6|Your own mouth condemns you, and not I; your own lips testify against you.
JOB|15|7|"Are you the first man who was born? Or were you brought forth before the hills?
JOB|15|8|Have you listened in the council of God? And do you limit wisdom to yourself?
JOB|15|9|What do you know that we do not know? What do you understand that is not clear to us?
JOB|15|10|Both the gray-haired and the aged are among us, older than your father.
JOB|15|11|Are the comforts of God too small for you, or the word that deals gently with you?
JOB|15|12|Why does your heart carry you away, and why do your eyes flash,
JOB|15|13|that you turn your spirit against God and bring such words out of your mouth?
JOB|15|14|What is man, that he can be pure? Or he who is born of a woman, that he can be righteous?
JOB|15|15|Behold, God puts no trust in his holy ones, and the heavens are not pure in his sight;
JOB|15|16|how much less one who is abominable and corrupt, a man who drinks injustice like water!
JOB|15|17|"I will show you; hear me, and what I have seen I will declare
JOB|15|18|(what wise men have told, without hiding it from their fathers,
JOB|15|19|to whom alone the land was given, and no stranger passed among them).
JOB|15|20|The wicked man writhes in pain all his days, through all the years that are laid up for the ruthless.
JOB|15|21|Dreadful sounds are in his ears; in prosperity the destroyer will come upon him.
JOB|15|22|He does not believe that he will return out of darkness, and he is marked for the sword.
JOB|15|23|He wanders abroad for bread, saying, 'Where is it?' He knows that a day of darkness is ready at his hand;
JOB|15|24|distress and anguish terrify him; they prevail against him, like a king ready for battle.
JOB|15|25|Because he has stretched out his hand against God and defies the Almighty,
JOB|15|26|running stubbornly against him with a thickly bossed shield;
JOB|15|27|because he has covered his face with his fat and gathered fat upon his waist
JOB|15|28|and has lived in desolate cities, in houses that none should inhabit, which were ready to become heaps of ruins;
JOB|15|29|he will not be rich, and his wealth will not endure, nor will his possessions spread over the earth;
JOB|15|30|he will not depart from darkness; the flame will dry up his shoots, and by the breath of his mouth he will depart.
JOB|15|31|Let him not trust in emptiness, deceiving himself, for emptiness will be his payment.
JOB|15|32|It will be paid in full before his time, and his branch will not be green.
JOB|15|33|He will shake off his unripe grape like the vine, and cast off his blossom like the olive tree.
JOB|15|34|For the company of the godless is barren, and fire consumes the tents of bribery.
JOB|15|35|They conceive trouble and give birth to evil, and their womb prepares deceit."
JOB|16|1|Then Job answered and said:
JOB|16|2|"I have heard many such things; miserable comforters are you all.
JOB|16|3|Shall windy words have an end? Or what provokes you that you answer?
JOB|16|4|I also could speak as you do, if you were in my place; I could join words together against you and shake my head at you.
JOB|16|5|I could strengthen you with my mouth, and the solace of my lips would assuage your pain.
JOB|16|6|"If I speak, my pain is not assuaged, and if I forbear, how much of it leaves me?
JOB|16|7|Surely now God has worn me out; he has made desolate all my company.
JOB|16|8|And he has shriveled me up, which is a witness against me, and my leanness has risen up against me; it testifies to my face.
JOB|16|9|He has torn me in his wrath and hated me; he has gnashed his teeth at me; my adversary sharpens his eyes against me.
JOB|16|10|Men have gaped at me with their mouth; they have struck me insolently on the cheek; they mass themselves together against me.
JOB|16|11|God gives me up to the ungodly and casts me into the hands of the wicked.
JOB|16|12|I was at ease, and he broke me apart; he seized me by the neck and dashed me to pieces; he set me up as his target;
JOB|16|13|his archers surround me. He slashes open my kidneys and does not spare; he pours out my gall on the ground.
JOB|16|14|He breaks me with breach upon breach; he runs upon me like a warrior.
JOB|16|15|I have sewed sackcloth upon my skin and have laid my strength in the dust.
JOB|16|16|My face is red with weeping, and on my eyelids is deep darkness,
JOB|16|17|although there is no violence in my hands, and my prayer is pure.
JOB|16|18|"O earth, cover not my blood, and let my cry find no resting place.
JOB|16|19|Even now, behold, my witness is in heaven, and he who testifies for me is on high.
JOB|16|20|My friends scorn me; my eye pours out tears to God,
JOB|16|21|that he would argue the case of a man with God, as a son of man does with his neighbor.
JOB|16|22|For when a few years have come I shall go the way from which I shall not return.
JOB|17|1|My spirit is broken; my days are extinct; the graveyard is ready for me.
JOB|17|2|Surely there are mockers about me, and my eye dwells on their provocation.
JOB|17|3|"Lay down a pledge for me with yourself; who is there who will put up security for me?
JOB|17|4|Since you have closed their hearts to understanding, therefore you will not let them triumph.
JOB|17|5|He who informs against his friends to get a share of their property- the eyes of his children will fail.
JOB|17|6|"He has made me a byword of the peoples, and I am one before whom men spit.
JOB|17|7|My eye has grown dim from vexation, and all my members are like a shadow.
JOB|17|8|The upright are appalled at this, and the innocent stirs himself up against the godless.
JOB|17|9|Yet the righteous holds to his way, and he who has clean hands grows stronger and stronger.
JOB|17|10|But you, come on again, all of you, and I shall not find a wise man among you.
JOB|17|11|My days are past; my plans are broken off, the desires of my heart.
JOB|17|12|They make night into day; 'The light,' they say, 'is near to the darkness.'
JOB|17|13|If I hope for Sheol as my house, if I make my bed in darkness,
JOB|17|14|if I say to the pit, 'You are my father,' and to the worm, 'My mother,' or 'My sister,'
JOB|17|15|where then is my hope? Who will see my hope?
JOB|17|16|Will it go down to the bars of Sheol? Shall we descend together into the dust?"
JOB|18|1|Then Bildad the Shuhite answered and said:
JOB|18|2|"How long will you hunt for words? Consider, and then we will speak.
JOB|18|3|Why are we counted as cattle? Why are we stupid in your sight?
JOB|18|4|You who tear yourself in your anger, shall the earth be forsaken for you, or the rock be removed out of its place?
JOB|18|5|"Indeed, the light of the wicked is put out, and the flame of his fire does not shine.
JOB|18|6|The light is dark in his tent, and his lamp above him is put out.
JOB|18|7|His strong steps are shortened, and his own schemes throw him down.
JOB|18|8|For he is cast into a net by his own feet, and he walks on its mesh.
JOB|18|9|A trap seizes him by the heel; a snare lays hold of him.
JOB|18|10|A rope is hidden for him in the ground, a trap for him in the path.
JOB|18|11|Terrors frighten him on every side, and chase him at his heels.
JOB|18|12|His strength is famished, and calamity is ready for his stumbling.
JOB|18|13|It consumes the parts of his skin; the firstborn of death consumes his limbs.
JOB|18|14|He is torn from the tent in which he trusted and is brought to the king of terrors.
JOB|18|15|In his tent dwells that which is none of his; sulfur is scattered over his habitation.
JOB|18|16|His roots dry up beneath, and his branches wither above.
JOB|18|17|His memory perishes from the earth, and he has no name in the street.
JOB|18|18|He is thrust from light into darkness, and driven out of the world.
JOB|18|19|He has no posterity or progeny among his people, and no survivor where he used to live.
JOB|18|20|They of the west are appalled at his day, and horror seizes them of the east.
JOB|18|21|Surely such are the dwellings of the unrighteous, such is the place of him who knows not God."
JOB|19|1|Then Job answered and said:
JOB|19|2|"How long will you torment me and break me in pieces with words?
JOB|19|3|These ten times you have cast reproach upon me; are you not ashamed to wrong me?
JOB|19|4|And even if it be true that I have erred, my error remains with myself.
JOB|19|5|If indeed you magnify yourselves against me and make my disgrace an argument against me,
JOB|19|6|know then that God has put me in the wrong and closed his net about me.
JOB|19|7|Behold, I cry out, 'Violence!' but I am not answered; I call for help, but there is no justice.
JOB|19|8|He has walled up my way, so that I cannot pass, and he has set darkness upon my paths.
JOB|19|9|He has stripped from me my glory and taken the crown from my head.
JOB|19|10|He breaks me down on every side, and I am gone, and my hope has he pulled up like a tree.
JOB|19|11|He has kindled his wrath against me and counts me as his adversary.
JOB|19|12|His troops come on together; they have cast up their siege ramp against me and encamp around my tent.
JOB|19|13|"He has put my brothers far from me, and those who knew me are wholly estranged from me.
JOB|19|14|My relatives have failed me, my close friends have forgotten me.
JOB|19|15|The guests in my house and my maidservants count me as a stranger; I have become a foreigner in their eyes.
JOB|19|16|I call to my servant, but he gives me no answer; I must plead with him with my mouth for mercy.
JOB|19|17|My breath is strange to my wife, and I am a stench to the children of my own mother.
JOB|19|18|Even young children despise me; when I rise they talk against me.
JOB|19|19|All my intimate friends abhor me, and those whom I loved have turned against me.
JOB|19|20|My bones stick to my skin and to my flesh, and I have escaped by the skin of my teeth.
JOB|19|21|Have mercy on me, have mercy on me, O you my friends, for the hand of God has touched me!
JOB|19|22|Why do you, like God, pursue me? Why are you not satisfied with my flesh?
JOB|19|23|"Oh that my words were written! Oh that they were inscribed in a book!
JOB|19|24|Oh that with an iron pen and lead they were engraved in the rock forever!
JOB|19|25|For I know that my Redeemer lives, and at the last he will stand upon the earth.
JOB|19|26|And after my skin has been thus destroyed, yet in my flesh I shall see God,
JOB|19|27|whom I shall see for myself, and my eyes shall behold, and not another. My heart faints within me!
JOB|19|28|If you say, 'How we will pursue him!' and, 'The root of the matter is found in him,'
JOB|19|29|be afraid of the sword, for wrath brings the punishment of the sword, that you may know there is a judgment."
JOB|20|1|Then Zophar the Naamathite answered and said:
JOB|20|2|"Therefore my thoughts answer me, because of my haste within me.
JOB|20|3|I hear censure that insults me, and out of my understanding a spirit answers me.
JOB|20|4|Do you not know this from of old, since man was placed on earth,
JOB|20|5|that the exulting of the wicked is short, and the joy of the godless but for a moment?
JOB|20|6|Though his height mount up to the heavens, and his head reach to the clouds,
JOB|20|7|he will perish forever like his own dung; those who have seen him will say, 'Where is he?'
JOB|20|8|He will fly away like a dream and not be found; he will be chased away like a vision of the night.
JOB|20|9|The eye that saw him will see him no more, nor will his place any more behold him.
JOB|20|10|His children will seek the favor of the poor, and his hands will give back his wealth.
JOB|20|11|His bones are full of his youthful vigor, but it will lie down with him in the dust.
JOB|20|12|"Though evil is sweet in his mouth, though he hides it under his tongue,
JOB|20|13|though he is loath to let it go and holds it in his mouth,
JOB|20|14|yet his food is turned in his stomach; it is the venom of cobras within him.
JOB|20|15|He swallows down riches and vomits them up again; God casts them out of his belly.
JOB|20|16|He will suck the poison of cobras; the tongue of a viper will kill him.
JOB|20|17|He will not look upon the rivers, the streams flowing with honey and curds.
JOB|20|18|He will give back the fruit of his toil and will not swallow it down; from the profit of his trading he will get no enjoyment.
JOB|20|19|For he has crushed and abandoned the poor; he has seized a house that he did not build.
JOB|20|20|"Because he knew no contentment in his belly, he will not let anything in which he delights escape him.
JOB|20|21|There was nothing left after he had eaten; therefore his prosperity will not endure.
JOB|20|22|In the fullness of his sufficiency he will be in distress; the hand of everyone in misery will come against him.
JOB|20|23|To fill his belly to the full God will send his burning anger against him and rain it upon him into his body.
JOB|20|24|He will flee from an iron weapon; a bronze arrow will strike him through.
JOB|20|25|It is drawn forth and comes out of his body; the glittering point comes out of his gallbladder; terrors come upon him.
JOB|20|26|Utter darkness is laid up for his treasures; a fire not fanned will devour him; what is left in his tent will be consumed.
JOB|20|27|The heavens will reveal his iniquity, and the earth will rise up against him.
JOB|20|28|The possessions of his house will be carried away, dragged off in the day of God's wrath.
JOB|20|29|This is the wicked man's portion from God, the heritage decreed for him by God."
JOB|21|1|Then Job answered and said:
JOB|21|2|"Keep listening to my words, and let this be your comfort.
JOB|21|3|Bear with me, and I will speak, and after I have spoken, mock on.
JOB|21|4|As for me, is my complaint against man? Why should I not be impatient?
JOB|21|5|Look at me and be appalled, and lay your hand over your mouth.
JOB|21|6|When I remember I am dismayed, and shuddering seizes my flesh.
JOB|21|7|Why do the wicked live, reach old age, and grow mighty in power?
JOB|21|8|Their offspring are established in their presence, and their descendants before their eyes.
JOB|21|9|Their houses are safe from fear, and no rod of God is upon them.
JOB|21|10|Their bull breeds without fail; their cow calves and does not miscarry.
JOB|21|11|They send out their little boys like a flock, and their children dance.
JOB|21|12|They sing to the tambourine and the lyre and rejoice to the sound of the pipe.
JOB|21|13|They spend their days in prosperity, and in peace they go down to Sheol.
JOB|21|14|They say to God, 'Depart from us! We do not desire the knowledge of your ways.
JOB|21|15|What is the Almighty, that we should serve him? And what profit do we get if we pray to him?'
JOB|21|16|Behold, is not their prosperity in their hand? The counsel of the wicked is far from me.
JOB|21|17|"How often is it that the lamp of the wicked is put out? That their calamity comes upon them? That God distributes pains in his anger?
JOB|21|18|That they are like straw before the wind, and like chaff that the storm carries away?
JOB|21|19|You say, 'God stores up their iniquity for their children.' Let him pay it out to them, that they may know it.
JOB|21|20|Let their own eyes see their destruction, and let them drink of the wrath of the Almighty.
JOB|21|21|For what do they care for their houses after them, when the number of their months is cut off?
JOB|21|22|Will any teach God knowledge, seeing that he judges those who are on high?
JOB|21|23|One dies in his full vigor, being wholly at ease and secure,
JOB|21|24|his pails full of milk and the marrow of his bones moist.
JOB|21|25|Another dies in bitterness of soul, never having tasted of prosperity.
JOB|21|26|They lie down alike in the dust, and the worms cover them.
JOB|21|27|"Behold, I know your thoughts and your schemes to wrong me.
JOB|21|28|For you say, 'Where is the house of the prince? Where is the tent in which the wicked lived?'
JOB|21|29|Have you not asked those who travel the roads, and do you not accept their testimony
JOB|21|30|that the evil man is spared in the day of calamity, that he is rescued in the day of wrath?
JOB|21|31|Who declares his way to his face, and who repays him for what he has done?
JOB|21|32|When he is carried to the grave, watch is kept over his tomb.
JOB|21|33|The clods of the valley are sweet to him; all mankind follows after him, and those who go before him are innumerable.
JOB|21|34|How then will you comfort me with empty nothings? There is nothing left of your answers but falsehood."
JOB|22|1|Then Eliphaz the Temanite answered and said:
JOB|22|2|"Can a man be profitable to God? Surely he who is wise is profitable to himself.
JOB|22|3|Is it any pleasure to the Almighty if you are in the right, or is it gain to him if you make your ways blameless?
JOB|22|4|Is it for your fear of him that he reproves you and enters into judgment with you?
JOB|22|5|Is not your evil abundant? There is no end to your iniquities.
JOB|22|6|For you have exacted pledges of your brothers for nothing and stripped the naked of their clothing.
JOB|22|7|You have given no water to the weary to drink, and you have withheld bread from the hungry.
JOB|22|8|The man with power possessed the land, and the favored man lived in it.
JOB|22|9|You have sent widows away empty, and the arms of the fatherless were crushed.
JOB|22|10|Therefore snares are all around you, and sudden terror overwhelms you,
JOB|22|11|or darkness, so that you cannot see, and a flood of water covers you.
JOB|22|12|"Is not God high in the heavens? See the highest stars, how lofty they are!
JOB|22|13|But you say, 'What does God know? Can he judge through the deep darkness?
JOB|22|14|Thick clouds veil him, so that he does not see, and he walks on the vault of heaven.'
JOB|22|15|Will you keep to the old way that wicked men have trod?
JOB|22|16|They were snatched away before their time; their foundation was washed away.
JOB|22|17|They said to God, 'Depart from us,' and 'What can the Almighty do to us?'
JOB|22|18|Yet he filled their houses with good things- but the counsel of the wicked is far from me.
JOB|22|19|The righteous see it and are glad; the innocent one mocks at them,
JOB|22|20|saying, 'Surely our adversaries are cut off, and what they left the fire has consumed.'
JOB|22|21|"Agree with God, and be at peace; thereby good will come to you.
JOB|22|22|Receive instruction from his mouth, and lay up his words in your heart.
JOB|22|23|If you return to the Almighty you will be built up; if you remove injustice far from your tents,
JOB|22|24|if you lay gold in the dust, and gold of Ophir among the stones of the torrent bed,
JOB|22|25|then the Almighty will be your gold and your precious silver.
JOB|22|26|For then you will delight yourself in the Almighty and lift up your face to God.
JOB|22|27|You will make your prayer to him, and he will hear you, and you will pay your vows.
JOB|22|28|You will decide on a matter, and it will be established for you, and light will shine on your ways.
JOB|22|29|For when they are humbled you say, 'It is because of pride'; but he saves the lowly.
JOB|22|30|He delivers even the one who is not innocent, who will be delivered through the cleanness of your hands."
JOB|23|1|Then Job answered and said:
JOB|23|2|"Today also my complaint is bitter; my hand is heavy on account of my groaning.
JOB|23|3|Oh, that I knew where I might find him, that I might come even to his seat!
JOB|23|4|I would lay my case before him and fill my mouth with arguments.
JOB|23|5|I would know what he would answer me and understand what he would say to me.
JOB|23|6|Would he contend with me in the greatness of his power? No; he would pay attention to me.
JOB|23|7|There an upright man could argue with him, and I would be acquitted forever by my judge.
JOB|23|8|"Behold, I go forward, but he is not there, and backward, but I do not perceive him;
JOB|23|9|on the left hand when he is working, I do not behold him; he turns to the right hand, but I do not see him.
JOB|23|10|But he knows the way that I take; when he has tried me, I shall come out as gold.
JOB|23|11|My foot has held fast to his steps; I have kept his way and have not turned aside.
JOB|23|12|I have not departed from the commandment of his lips; I have treasured the words of his mouth more than my portion of food.
JOB|23|13|But he is unchangeable, and who can turn him back? What he desires, that he does.
JOB|23|14|For he will complete what he appoints for me, and many such things are in his mind.
JOB|23|15|Therefore I am terrified at his presence; when I consider, I am in dread of him.
JOB|23|16|God has made my heart faint; the Almighty has terrified me;
JOB|23|17|yet I am not silenced because of the darkness, nor because thick darkness covers my face.
JOB|24|1|"Why are not times of judgment kept by the Almighty, and why do those who know him never see his days?
JOB|24|2|Some move landmarks; they seize flocks and pasture them.
JOB|24|3|They drive away the donkey of the fatherless; they take the widow's ox for a pledge.
JOB|24|4|They thrust the poor off the road; the poor of the earth all hide themselves.
JOB|24|5|Behold, like wild donkeys in the desert the poor go out to their toil, seeking game; the wasteland yields food for their children.
JOB|24|6|They gather their fodder in the field, and they glean the vineyard of the wicked man.
JOB|24|7|They lie all night naked, without clothing, and have no covering in the cold.
JOB|24|8|They are wet with the rain of the mountains and cling to the rock for lack of shelter.
JOB|24|9|(There are those who snatch the fatherless child from the breast, and they take a pledge against the poor.)
JOB|24|10|They go about naked, without clothing; hungry, they carry the sheaves;
JOB|24|11|among the olive rows of the wicked they make oil; they tread the winepresses, but suffer thirst.
JOB|24|12|From out of the city the dying groan, and the soul of the wounded cries for help; yet God charges no one with wrong.
JOB|24|13|"There are those who rebel against the light, who are not acquainted with its ways, and do not stay in its paths.
JOB|24|14|The murderer rises before it is light, that he may kill the poor and needy, and in the night he is like a thief.
JOB|24|15|The eye of the adulterer also waits for the twilight, saying, 'No eye will see me'; and he veils his face.
JOB|24|16|In the dark they dig through houses; by day they shut themselves up; they do not know the light.
JOB|24|17|For deep darkness is morning to all of them; for they are friends with the terrors of deep darkness.
JOB|24|18|"You say, 'Swift are they on the face of the waters; their portion is cursed in the land; no treader turns toward their vineyards.
JOB|24|19|Drought and heat snatch away the snow waters; so does Sheol those who have sinned.
JOB|24|20|The womb forgets them; the worm finds them sweet; they are no longer remembered, so wickedness is broken like a tree.'
JOB|24|21|"They wrong the barren childless woman, and do no good to the widow.
JOB|24|22|Yet God prolongs the life of the mighty by his power; they rise up when they despair of life.
JOB|24|23|He gives them security, and they are supported, and his eyes are upon their ways.
JOB|24|24|They are exalted a little while, and then are gone; they are brought low and gathered up like all others; they are cut off like the heads of grain.
JOB|24|25|If it is not so, who will prove me a liar and show that there is nothing in what I say?"
JOB|25|1|Then Bildad the Shuhite answered and said:
JOB|25|2|"Dominion and fear are with God; he makes peace in his high heaven.
JOB|25|3|Is there any number to his armies? Upon whom does his light not arise?
JOB|25|4|How then can man be in the right before God? How can he who is born of woman be pure?
JOB|25|5|Behold, even the moon is not bright, and the stars are not pure in his eyes;
JOB|25|6|how much less man, who is a maggot, and the son of man, who is a worm!"
JOB|26|1|Then Job answered and said:
JOB|26|2|"How you have helped him who has no power! How you have saved the arm that has no strength!
JOB|26|3|How you have counseled him who has no wisdom, and plentifully declared sound knowledge!
JOB|26|4|With whose help have you uttered words, and whose breath has come out from you?
JOB|26|5|The dead tremble under the waters and their inhabitants.
JOB|26|6|Sheol is naked before God, and Abaddon has no covering.
JOB|26|7|He stretches out the north over the void and hangs the earth on nothing.
JOB|26|8|He binds up the waters in his thick clouds, and the cloud is not split open under them.
JOB|26|9|He covers the face of the full moon and spreads over it his cloud.
JOB|26|10|He has inscribed a circle on the face of the waters at the boundary between light and darkness.
JOB|26|11|The pillars of heaven tremble and are astounded at his rebuke.
JOB|26|12|By his power he stilled the sea; by his understanding he shattered Rahab.
JOB|26|13|By his wind the heavens were made fair; his hand pierced the fleeing serpent.
JOB|26|14|Behold, these are but the outskirts of his ways, and how small a whisper do we hear of him! But the thunder of his power who can understand?"
JOB|27|1|And Job again took up his discourse, and said:
JOB|27|2|"As God lives, who has taken away my right, and the Almighty, who has made my soul bitter,
JOB|27|3|as long as my breath is in me, and the spirit of God is in my nostrils,
JOB|27|4|my lips will not speak falsehood, and my tongue will not utter deceit.
JOB|27|5|Far be it from me to say that you are right; till I die I will not put away my integrity from me.
JOB|27|6|I hold fast my righteousness and will not let it go; my heart does not reproach me for any of my days.
JOB|27|7|"Let my enemy be as the wicked, and let him who rises up against me be as the unrighteous.
JOB|27|8|For what is the hope of the godless when God cuts him off, when God takes away his life?
JOB|27|9|Will God hear his cry when distress comes upon him?
JOB|27|10|Will he take delight in the Almighty? Will he call upon God at all times?
JOB|27|11|I will teach you concerning the hand of God; what is with the Almighty I will not conceal.
JOB|27|12|Behold, all of you have seen it yourselves; why then have you become altogether vain?
JOB|27|13|"This is the portion of a wicked man with God, and the heritage that oppressors receive from the Almighty:
JOB|27|14|If his children are multiplied, it is for the sword, and his descendants have not enough bread.
JOB|27|15|Those who survive him the pestilence buries, and his widows do not weep.
JOB|27|16|Though he heap up silver like dust, and pile up clothing like clay,
JOB|27|17|he may pile it up, but the righteous will wear it, and the innocent will divide the silver.
JOB|27|18|He builds his house like a moth's, like a booth that a watchman makes.
JOB|27|19|He goes to bed rich, but will do so no more; he opens his eyes, and his wealth is gone.
JOB|27|20|Terrors overtake him like a flood; in the night a whirlwind carries him off.
JOB|27|21|The east wind lifts him up and he is gone; it sweeps him out of his place.
JOB|27|22|It hurls at him without pity; he flees from its power in headlong flight.
JOB|27|23|It claps its hands at him and hisses at him from its place.
JOB|28|1|"Surely there is a mine for silver, and a place for gold that they refine.
JOB|28|2|Iron is taken out of the earth, and copper is smelted from the ore.
JOB|28|3|Man puts an end to darkness and searches out to the farthest limit the ore in gloom and deep darkness.
JOB|28|4|He opens shafts in a valley away from where anyone lives; they are forgotten by travelers; they hang in the air, far away from mankind; they swing to and fro.
JOB|28|5|As for the earth, out of it comes bread, but underneath it is turned up as by fire.
JOB|28|6|Its stones are the place of sapphires, and it has dust of gold.
JOB|28|7|"That path no bird of prey knows, and the falcon's eye has not seen it.
JOB|28|8|The proud beasts have not trodden it; the lion has not passed over it.
JOB|28|9|"Man puts his hand to the flinty rock and overturns mountains by the roots.
JOB|28|10|He cuts out channels in the rocks, and his eye sees every precious thing.
JOB|28|11|He dams up the streams so that they do not trickle, and the thing that is hidden he brings out to light.
JOB|28|12|"But where shall wisdom be found? And where is the place of understanding?
JOB|28|13|Man does not know its worth, and it is not found in the land of the living.
JOB|28|14|The deep says, 'It is not in me,' and the sea says, 'It is not with me.'
JOB|28|15|It cannot be bought for gold, and silver cannot be weighed as its price.
JOB|28|16|It cannot be valued in the gold of Ophir, in precious onyx or sapphire.
JOB|28|17|Gold and glass cannot equal it, nor can it be exchanged for jewels of fine gold.
JOB|28|18|No mention shall be made of coral or of crystal; the price of wisdom is above, pearls.
JOB|28|19|The topaz of Ethiopia cannot equal it, nor can it be valued in pure gold.
JOB|28|20|"From where, then, does wisdom come? And where is the place of understanding?
JOB|28|21|It is hidden from the eyes of all living and concealed from the birds of the air.
JOB|28|22|Abaddon and Death say, 'We have heard a rumor of it with our ears.'
JOB|28|23|"God understands the way to it, and he knows its place.
JOB|28|24|For he looks to the ends of the earth and sees everything under the heavens.
JOB|28|25|When he gave to the wind its weight and apportioned the waters by measure,
JOB|28|26|when he made a decree for the rain and a way for the lightning of the thunder,
JOB|28|27|then he saw it and declared it; he established it, and searched it out.
JOB|28|28|And he said to man, 'Behold, the fear of the Lord, that is wisdom, and to turn away from evil is understanding.'"
JOB|29|1|And Job again took up his discourse, and said:
JOB|29|2|"Oh, that I were as in the months of old, as in the days when God watched over me,
JOB|29|3|when his lamp shone upon my head, and by his light I walked through darkness,
JOB|29|4|as I was in my prime, when the friendship of God was upon my tent,
JOB|29|5|when the Almighty was yet with me, when my children were all around me,
JOB|29|6|when my steps were washed with butter, and the rock poured out for me streams of oil!
JOB|29|7|When I went out to the gate of the city, when I prepared my seat in the square,
JOB|29|8|the young men saw me and withdrew, and the aged rose and stood;
JOB|29|9|the princes refrained from talking and laid their hand on their mouth;
JOB|29|10|the voice of the nobles was hushed, and their tongue stuck to the roof of their mouth.
JOB|29|11|When the ear heard, it called me blessed, and when the eye saw, it approved,
JOB|29|12|because I delivered the poor who cried for help, and the fatherless who had none to help him.
JOB|29|13|The blessing of him who was about to perish came upon me, and I caused the widow's heart to sing for joy.
JOB|29|14|I put on righteousness, and it clothed me; my justice was like a robe and a turban.
JOB|29|15|I was eyes to the blind and feet to the lame.
JOB|29|16|I was a father to the needy, and I searched out the cause of him whom I did not know.
JOB|29|17|I broke the fangs of the unrighteous and made him drop his prey from his teeth.
JOB|29|18|Then I thought, 'I shall die in my nest, and I shall multiply my days as the sand,
JOB|29|19|my roots spread out to the waters, with the dew all night on my branches,
JOB|29|20|my glory fresh with me, and my bow ever new in my hand.'
JOB|29|21|"Men listened to me and waited and kept silence for my counsel.
JOB|29|22|After I spoke they did not speak again, and my word dropped upon them.
JOB|29|23|They waited for me as for the rain, and they opened their mouths as for the spring rain.
JOB|29|24|I smiled on them when they had no confidence, and the light of my face they did not cast down.
JOB|29|25|I chose their way and sat as chief, and I lived like a king among his troops, like one who comforts mourners.
JOB|30|1|"But now they laugh at me, men who are younger than I, whose fathers I would have disdained to set with the dogs of my flock.
JOB|30|2|What could I gain from the strength of their hands, men whose vigor is gone?
JOB|30|3|Through want and hard hunger they gnaw the dry ground by night in waste and desolation;
JOB|30|4|they pick saltwort and the leaves of bushes, and the roots of the broom tree for their food.
JOB|30|5|They are driven out from human company; they shout after them as after a thief.
JOB|30|6|In the gullies of the torrents they must dwell, in holes of the earth and of the rocks.
JOB|30|7|Among the bushes they bray; under the nettles they huddle together.
JOB|30|8|A senseless, a nameless brood, they have been whipped out of the land.
JOB|30|9|"And now I have become their song; I am a byword to them.
JOB|30|10|They abhor me; they keep aloof from me; they do not hesitate to spit at the sight of me.
JOB|30|11|Because God has loosed my cord and humbled me, they have cast off restraint in my presence.
JOB|30|12|On my right hand the rabble rise; they push away my feet; they cast up against me their ways of destruction.
JOB|30|13|They break up my path; they promote my calamity; they need no one to help them.
JOB|30|14|As through a wide breach they come; amid the crash they roll on.
JOB|30|15|Terrors are turned upon me; my honor is pursued as by the wind, and my prosperity has passed away like a cloud.
JOB|30|16|"And now my soul is poured out within me; days of affliction have taken hold of me.
JOB|30|17|The night racks my bones, and the pain that gnaws me takes no rest.
JOB|30|18|With great force my garment is disfigured; it binds me about like the collar of my tunic.
JOB|30|19|God has cast me into the mire, and I have become like dust and ashes.
JOB|30|20|I cry to you for help and you do not answer me; I stand, and you only look at me.
JOB|30|21|You have turned cruel to me; with the might of your hand you persecute me.
JOB|30|22|You lift me up on the wind; you make me ride on it, and you toss me about in the roar of the storm.
JOB|30|23|For I know that you will bring me to death and to the house appointed for all living.
JOB|30|24|"Yet does not one in a heap of ruins stretch out his hand, and in his disaster cry for help?
JOB|30|25|Did not I weep for him whose day was hard? Was not my soul grieved for the needy?
JOB|30|26|But when I hoped for good, evil came, and when I waited for light, darkness came.
JOB|30|27|My inward parts are in turmoil and never still; days of affliction come to meet me.
JOB|30|28|I go about darkened, but not by the sun; I stand up in the assembly and cry for help.
JOB|30|29|I am a brother of jackals and a companion of ostriches.
JOB|30|30|My skin turns black and falls from me, and my bones burn with heat.
JOB|30|31|My lyre is turned to mourning, and my pipe to the voice of those who weep.
JOB|31|1|"I have made a covenant with my eyes; how then could I gaze at a virgin?
JOB|31|2|What would be my portion from God above and my heritage from the Almighty on high?
JOB|31|3|Is not calamity for the unrighteous, and disaster for the workers of iniquity?
JOB|31|4|Does not he see my ways and number all my steps?
JOB|31|5|"If I have walked with falsehood and my foot has hastened to deceit;
JOB|31|6|(Let me be weighed in a just balance, and let God know my integrity!)
JOB|31|7|if my step has turned aside from the way and my heart has gone after my eyes, and if any spot has stuck to my hands,
JOB|31|8|then let me sow, and another eat, and let what grows for me be rooted out.
JOB|31|9|"If my heart has been enticed toward a woman, and I have lain in wait at my neighbor's door,
JOB|31|10|then let my wife grind for another, and let others bow down on her.
JOB|31|11|For that would be a heinous crime; that would be an iniquity to be punished by the judges;
JOB|31|12|for that would be a fire that consumes as far as Abaddon, and it would burn to the root all my increase.
JOB|31|13|"If I have rejected the cause of my manservant or my maidservant, when they brought a complaint against me,
JOB|31|14|what then shall I do when God rises up? When he makes inquiry, what shall I answer him?
JOB|31|15|Did not he who made me in the womb make him? And did not one fashion us in the womb?
JOB|31|16|"If I have withheld anything that the poor desired, or have caused the eyes of the widow to fail,
JOB|31|17|or have eaten my morsel alone, and the fatherless has not eaten of it
JOB|31|18|(for from my youth the fatherless grew up with me as with a father, and from my mother's womb I guided the widow),
JOB|31|19|if I have seen anyone perish for lack of clothing, or the needy without covering,
JOB|31|20|if his body has not blessed me, and if he was not warmed with the fleece of my sheep,
JOB|31|21|if I have raised my hand against the fatherless, because I saw my help in the gate,
JOB|31|22|then let my shoulder blade fall from my shoulder, and let my arm be broken from its socket.
JOB|31|23|For I was in terror of calamity from God, and I could not have faced his majesty.
JOB|31|24|"If I have made gold my trust or called fine gold my confidence,
JOB|31|25|if I have rejoiced because my wealth was abundant or because my hand had found much,
JOB|31|26|if I have looked at the sun when it shone, or the moon moving in splendor,
JOB|31|27|and my heart has been secretly enticed, and my mouth has kissed my hand,
JOB|31|28|this also would be an iniquity to be punished by the judges, for I would have been false to God above.
JOB|31|29|"If I have rejoiced at the ruin of him who hated me, or exulted when evil overtook him
JOB|31|30|(I have not let my mouth sin by asking for his life with a curse),
JOB|31|31|if the men of my tent have not said, 'Who is there that has not been filled with his meat?'
JOB|31|32|(the sojourner has not lodged in the street; I have opened my doors to the traveler),
JOB|31|33|if I have concealed my transgressions as others do by hiding my iniquity in my bosom,
JOB|31|34|because I stood in great fear of the multitude, and the contempt of families terrified me, so that I kept silence, and did not go out of doors-
JOB|31|35|Oh, that I had one to hear me! (Here is my signature! Let the Almighty answer me!) Oh, that I had the indictment written by my adversary!
JOB|31|36|Surely I would carry it on my shoulder; I would bind it on me as a crown;
JOB|31|37|I would give him an account of all my steps; like a prince I would approach him.
JOB|31|38|"If my land has cried out against me and its furrows have wept together,
JOB|31|39|if I have eaten its yield without payment and made its owners breathe their last,
JOB|31|40|let thorns grow instead of wheat, and foul weeds instead of barley." The words of Job are ended.
JOB|32|1|So these three men ceased to answer Job, because he was righteous in his own eyes.
JOB|32|2|Then Elihu the son of Barachel the Buzite, of the family of Ram, burned with anger. He burned with anger at Job because he justified himself rather than God.
JOB|32|3|He burned with anger also at Job's three friends because they had found no answer, although they had declared Job to be in the wrong.
JOB|32|4|Now Elihu had waited to speak to Job because they were older than he.
JOB|32|5|And when Elihu saw that there was no answer in the mouth of these three men, he burned with anger.
JOB|32|6|And Elihu the son of Barachel the Buzite answered and said: "I am young in years, and you are aged; therefore I was timid and afraid to declare my opinion to you.
JOB|32|7|I said, 'Let days speak, and many years teach wisdom.'
JOB|32|8|But it is the spirit in man, the breath of the Almighty, that makes him understand.
JOB|32|9|It is not the old who are wise, nor the aged who understand what is right.
JOB|32|10|Therefore I say, 'Listen to me; let me also declare my opinion.'
JOB|32|11|"Behold, I waited for your words, I listened for your wise sayings, while you searched out what to say.
JOB|32|12|I gave you my attention, and, behold, there was none among you who refuted Job or who answered his words.
JOB|32|13|Beware lest you say, 'We have found wisdom; God may vanquish him, not a man.'
JOB|32|14|He has not directed his words against me, and I will not answer him with your speeches.
JOB|32|15|"They are dismayed; they answer no more; they have not a word to say.
JOB|32|16|And shall I wait, because they do not speak, because they stand there, and answer no more?
JOB|32|17|I also will answer with my share; I also will declare my opinion.
JOB|32|18|For I am full of words; the spirit within me constrains me.
JOB|32|19|Behold, my belly is like wine that has no vent; like new wineskins ready to burst.
JOB|32|20|I must speak, that I may find relief; I must open my lips and answer.
JOB|32|21|I will not show partiality to any man or use flattery toward any person.
JOB|32|22|For I do not know how to flatter, else my Maker would soon take me away.
JOB|33|1|"But now, hear my speech, O Job, and listen to all my words.
JOB|33|2|Behold, I open my mouth; the tongue in my mouth speaks.
JOB|33|3|My words declare the uprightness of my heart, and what my lips know they speak sincerely.
JOB|33|4|The Spirit of God has made me, and the breath of the Almighty gives me life.
JOB|33|5|Answer me, if you can; set your words in order before me; take your stand.
JOB|33|6|Behold, I am toward God as you are; I too was pinched off from a piece of clay.
JOB|33|7|Behold, no fear of me need terrify you; my pressure will not be heavy upon you.
JOB|33|8|"Surely you have spoken in my ears, and I have heard the sound of your words.
JOB|33|9|You say, 'I am pure, without transgression; I am clean, and there is no iniquity in me.
JOB|33|10|Behold, he finds occasions against me, he counts me as his enemy,
JOB|33|11|he puts my feet in the stocks and watches all my paths.'
JOB|33|12|"Behold, in this you are not right. I will answer you, for God is greater than man.
JOB|33|13|Why do you contend against him, saying, 'He will answer none of man's words'?
JOB|33|14|For God speaks in one way, and in two, though man does not perceive it.
JOB|33|15|In a dream, in a vision of the night, when deep sleep falls on men, while they slumber on their beds,
JOB|33|16|then he opens the ears of men and terrifies them with warnings,
JOB|33|17|that he may turn man aside from his deed and conceal pride from a man;
JOB|33|18|he keeps back his soul from the pit, his life from perishing by the sword.
JOB|33|19|"Man is also rebuked with pain on his bed and with continual strife in his bones,
JOB|33|20|so that his life loathes bread, and his appetite the choicest food.
JOB|33|21|His flesh is so wasted away that it cannot be seen, and his bones that were not seen stick out.
JOB|33|22|His soul draws near the pit, and his life to those who bring death.
JOB|33|23|If there be for him an angel, a mediator, one of the thousand, to declare to man what is right for him,
JOB|33|24|and he is merciful to him, and says, 'Deliver him from going down into the pit; I have found a ransom;
JOB|33|25|let his flesh become fresh with youth; let him return to the days of his youthful vigor';
JOB|33|26|then man prays to God, and he accepts him; he sees his face with a shout of joy, and he restores to man his righteousness.
JOB|33|27|He sings before men and says: 'I sinned and perverted what was right, and it was not repaid to me.
JOB|33|28|He has redeemed my soul from going down into the pit, and my life shall look upon the light.'
JOB|33|29|"Behold, God does all these things, twice, three times, with a man,
JOB|33|30|to bring back his soul from the pit, that he may be lighted with the light of life.
JOB|33|31|Pay attention, O Job, listen to me; be silent, and I will speak.
JOB|33|32|If you have any words, answer me; speak, for I desire to justify you.
JOB|33|33|If not, listen to me; be silent, and I will teach you wisdom."
JOB|34|1|Then Elihu answered and said:
JOB|34|2|"Hear my words, you wise men, and give ear to me, you who know;
JOB|34|3|for the ear tests words as the palate tastes food.
JOB|34|4|Let us choose what is right; let us know among ourselves what is good.
JOB|34|5|For Job has said, 'I am in the right, and God has taken away my right;
JOB|34|6|in spite of my right I am counted a liar; my wound is incurable, though I am without transgression.'
JOB|34|7|What man is like Job, who drinks up scoffing like water,
JOB|34|8|who travels in company with evildoers and walks with wicked men?
JOB|34|9|For he has said, 'It profits a man nothing that he should take delight in God.'
JOB|34|10|"Therefore, hear me, you men of understanding: far be it from God that he should do wickedness, and from the Almighty that he should do wrong.
JOB|34|11|For according to the work of a man he will repay him, and according to his ways he will make it befall him.
JOB|34|12|Of a truth, God will not do wickedly, and the Almighty will not pervert justice.
JOB|34|13|Who gave him charge over the earth, and who laid on him the whole world?
JOB|34|14|If he should set his heart to it and gather to himself his spirit and his breath,
JOB|34|15|all flesh would perish together, and man would return to dust.
JOB|34|16|"If you have understanding, hear this; listen to what I say.
JOB|34|17|Shall one who hates justice govern? Will you condemn him who is righteous and mighty,
JOB|34|18|who says to a king, 'Worthless one,' and to nobles, 'Wicked man,'
JOB|34|19|who shows no partiality to princes, nor regards the rich more than the poor, for they are all the work of his hands?
JOB|34|20|In a moment they die; at midnight the people are shaken and pass away, and the mighty are taken away by no human hand.
JOB|34|21|"For his eyes are on the ways of a man, and he sees all his steps.
JOB|34|22|There is no gloom or deep darkness where evildoers may hide themselves.
JOB|34|23|For God has no need to consider a man further, that he should go before God in judgment.
JOB|34|24|He shatters the mighty without investigation and sets others in their place.
JOB|34|25|Thus, knowing their works, he overturns them in the night, and they are crushed.
JOB|34|26|He strikes them for their wickedness in a place for all to see,
JOB|34|27|because they turned aside from following him and had no regard for any of his ways,
JOB|34|28|so that they caused the cry of the poor to come to him, and he heard the cry of the afflicted-
JOB|34|29|When he is quiet, who can condemn? When he hides his face, who can behold him, whether it be a nation or a man?-
JOB|34|30|that a godless man should not reign, that he should not ensnare the people.
JOB|34|31|"For has anyone said to God, 'I have borne punishment; I will not offend any more;
JOB|34|32|teach me what I do not see; if I have done iniquity, I will do it no more'?
JOB|34|33|Will he then make repayment to suit you, because you reject it? For you must choose, and not I; therefore declare what you know.
JOB|34|34|Men of understanding will say to me, and the wise man who hears me will say:
JOB|34|35|'Job speaks without knowledge; his words are without insight.'
JOB|34|36|Would that Job were tried to the end, because he answers like wicked men.
JOB|34|37|For he adds rebellion to his sin; he claps his hands among us and multiplies his words against God."
JOB|35|1|And Elihu answered and said:
JOB|35|2|"Do you think this to be just? Do you say, 'It is my right before God,'
JOB|35|3|that you ask, 'What advantage have I? How am I better off than if I had sinned?'
JOB|35|4|I will answer you and your friends with you.
JOB|35|5|Look at the heavens, and see; and behold the clouds, which are higher than you.
JOB|35|6|If you have sinned, what do you accomplish against him? And if your transgressions are multiplied, what do you do to him?
JOB|35|7|If you are righteous, what do you give to him? Or what does he receive from your hand?
JOB|35|8|Your wickedness concerns a man like yourself, and your righteousness a son of man.
JOB|35|9|"Because of the multitude of oppressions people cry out; they call for help because of the arm of the mighty.
JOB|35|10|But none says, 'Where is God my Maker, who gives songs in the night,
JOB|35|11|who teaches us more than the beasts of the earth and makes us wiser than the birds of the heavens?'
JOB|35|12|There they cry out, but he does not answer, because of the pride of evil men.
JOB|35|13|Surely God does not hear an empty cry, nor does the Almighty regard it.
JOB|35|14|How much less when you say that you do not see him, that the case is before him, and you are waiting for him!
JOB|35|15|And now, because his anger does not punish, and he does not take much note of transgression,
JOB|35|16|Job opens his mouth in empty talk; he multiplies words without knowledge."
JOB|36|1|And Elihu continued, and said:
JOB|36|2|"Bear with me a little, and I will show you, for I have yet something to say on God's behalf.
JOB|36|3|I will get my knowledge from afar and ascribe righteousness to my Maker.
JOB|36|4|For truly my words are not false; one who is perfect in knowledge is with you.
JOB|36|5|"Behold, God is mighty, and does not despise any; he is mighty in strength of understanding.
JOB|36|6|He does not keep the wicked alive, but gives the afflicted their right.
JOB|36|7|He does not withdraw his eyes from the righteous, but with kings on the throne he sets them forever, and they are exalted.
JOB|36|8|And if they are bound in chains and caught in the cords of affliction,
JOB|36|9|then he declares to them their work and their transgressions, that they are behaving arrogantly.
JOB|36|10|He opens their ears to instruction and commands that they return from iniquity.
JOB|36|11|If they listen and serve him, they complete their days in prosperity, and their years in pleasantness.
JOB|36|12|But if they do not listen, they perish by the sword and die without knowledge.
JOB|36|13|"The godless in heart cherish anger; they do not cry for help when he binds them.
JOB|36|14|They die in youth, and their life ends among the cult prostitutes.
JOB|36|15|He delivers the afflicted by their affliction and opens their ear by adversity.
JOB|36|16|He also allured you out of distress into a broad place where there was no cramping, and what was set on your table was full of fatness.
JOB|36|17|"But you are full of the judgment on the wicked; judgment and justice seize you.
JOB|36|18|Beware lest wrath entice you into scoffing, and let not the greatness of the ransom turn you aside.
JOB|36|19|Will your cry for help avail to keep you from distress, or all the force of your strength?
JOB|36|20|Do not long for the night, when peoples vanish in their place.
JOB|36|21|Take care; do not turn to iniquity, for this you have chosen rather than affliction.
JOB|36|22|Behold, God is exalted in his power; who is a teacher like him?
JOB|36|23|Who has prescribed for him his way, or who can say, 'You have done wrong'?
JOB|36|24|"Remember to extol his work, of which men have sung.
JOB|36|25|All mankind has looked on it; man beholds it from afar.
JOB|36|26|Behold, God is great, and we know him not; the number of his years is unsearchable.
JOB|36|27|For he draws up the drops of water; they distill his mist in rain,
JOB|36|28|which the skies pour down and drop on mankind abundantly.
JOB|36|29|Can anyone understand the spreading of the clouds, the thunderings of his pavilion?
JOB|36|30|Behold, he scatters his lightning about him and covers the roots of the sea.
JOB|36|31|For by these he judges peoples; he gives food in abundance.
JOB|36|32|He covers his hands with the lightning and commands it to strike the mark.
JOB|36|33|Its crashing declares his presence; the cattle also declare that he rises.
JOB|37|1|"At this also my heart trembles and leaps out of its place.
JOB|37|2|Keep listening to the thunder of his voice and the rumbling that comes from his mouth.
JOB|37|3|Under the whole heaven he lets it go, and his lightning to the corners of the earth.
JOB|37|4|After it his voice roars; he thunders with his majestic voice, and he does not restrain the lightnings when his voice is heard.
JOB|37|5|God thunders wondrously with his voice; he does great things that we cannot comprehend.
JOB|37|6|For to the snow he says, 'Fall on the earth,' likewise to the downpour, his mighty downpour.
JOB|37|7|He seals up the hand of every man, that all men whom he made may know it.
JOB|37|8|Then the beasts go into their lairs, and remain in their dens.
JOB|37|9|From its chamber comes the whirlwind, and cold from the scattering winds.
JOB|37|10|By the breath of God ice is given, and the broad waters are frozen fast.
JOB|37|11|He loads the thick cloud with moisture; the clouds scatter his lightning.
JOB|37|12|They turn around and around by his guidance, to accomplish all that he commands them on the face of the habitable world.
JOB|37|13|Whether for correction or for his land or for love, he causes it to happen.
JOB|37|14|"Hear this, O Job; stop and consider the wondrous works of God.
JOB|37|15|Do you know how God lays his command upon them and causes the lightning of his cloud to shine?
JOB|37|16|Do you know the balancings of the clouds, the wondrous works of him who is perfect in knowledge,
JOB|37|17|you whose garments are hot when the earth is still because of the south wind?
JOB|37|18|Can you, like him, spread out the skies, hard as a cast metal mirror?
JOB|37|19|Teach us what we shall say to him; we cannot draw up our case because of darkness.
JOB|37|20|Shall it be told him that I would speak? Did a man ever wish that he would be swallowed up?
JOB|37|21|"And now no one looks on the light when it is bright in the skies, when the wind has passed and cleared them.
JOB|37|22|Out of the north comes golden splendor; God is clothed with awesome majesty.
JOB|37|23|The Almighty- we cannot find him; he is great in power; justice and abundant righteousness he will not violate.
JOB|37|24|Therefore men fear him; he does not regard any who are wise in their own conceit."
JOB|38|1|Then the LORD answered Job out of the whirlwind and said:
JOB|38|2|"Who is this that darkens counsel by words without knowledge?
JOB|38|3|Dress for action like a man; I will question you, and you make it known to me.
JOB|38|4|"Where were you when I laid the foundation of the earth? Tell me, if you have understanding.
JOB|38|5|Who determined its measurements- surely you know! Or who stretched the line upon it?
JOB|38|6|On what were its bases sunk, or who laid its cornerstone,
JOB|38|7|when the morning stars sang together and all the sons of God shouted for joy?
JOB|38|8|"Or who shut in the sea with doors when it burst out from the womb,
JOB|38|9|when I made clouds its garment and thick darkness its swaddling band,
JOB|38|10|and prescribed limits for it and set bars and doors,
JOB|38|11|and said, 'Thus far shall you come, and no farther, and here shall your proud waves be stayed'?
JOB|38|12|"Have you commanded the morning since your days began, and caused the dawn to know its place,
JOB|38|13|that it might take hold of the skirts of the earth, and the wicked be shaken out of it?
JOB|38|14|It is changed like clay under the seal, and its features stand out like a garment.
JOB|38|15|From the wicked their light is withheld, and their uplifted arm is broken.
JOB|38|16|"Have you entered into the springs of the sea, or walked in the recesses of the deep?
JOB|38|17|Have the gates of death been revealed to you, or have you seen the gates of deep darkness?
JOB|38|18|Have you comprehended the expanse of the earth? Declare, if you know all this.
JOB|38|19|"Where is the way to the dwelling of light, and where is the place of darkness,
JOB|38|20|that you may take it to its territory and that you may discern the paths to its home?
JOB|38|21|You know, for you were born then, and the number of your days is great!
JOB|38|22|"Have you entered the storehouses of the snow, or have you seen the storehouses of the hail,
JOB|38|23|which I have reserved for the time of trouble, for the day of battle and war?
JOB|38|24|What is the way to the place where the light is distributed, or where the east wind is scattered upon the earth?
JOB|38|25|"Who has cleft a channel for the torrents of rain and a way for the thunderbolt,
JOB|38|26|to bring rain on a land where no man is, on the desert in which there is no man,
JOB|38|27|to satisfy the waste and desolate land, and to make the ground sprout with grass?
JOB|38|28|"Has the rain a father, or who has begotten the drops of dew?
JOB|38|29|From whose womb did the ice come forth, and who has given birth to the frost of heaven?
JOB|38|30|The waters become hard like stone, and the face of the deep is frozen.
JOB|38|31|"Can you bind the chains of the Pleiades or loose the cords of Orion?
JOB|38|32|Can you lead forth the Mazzaroth1 in their season, or can you guide the Bear with its children?
JOB|38|33|Do you know the ordinances of the heavens? Can you establish their rule on the earth?
JOB|38|34|"Can you lift up your voice to the clouds, that a flood of waters may cover you?
JOB|38|35|Can you send forth lightnings, that they may go and say to you, 'Here we are'?
JOB|38|36|Who has put wisdom in the inward parts or given understanding to the mind?
JOB|38|37|Who can number the clouds by wisdom? Or who can tilt the waterskins of the heavens,
JOB|38|38|when the dust runs into a mass and the clods stick fast together?
JOB|38|39|"Can you hunt the prey for the lion, or satisfy the appetite of the young lions,
JOB|38|40|when they crouch in their dens or lie in wait in their thicket?
JOB|38|41|Who provides for the raven its prey, when its young ones cry to God for help, and wander about for lack of food?
JOB|39|1|"Do you know when the mountain goats give birth? Do you observe the calving of the does?
JOB|39|2|Can you number the months that they fulfill, and do you know the time when they give birth,
JOB|39|3|when they crouch, bring forth their offspring, and are delivered of their young?
JOB|39|4|Their young ones become strong; they grow up in the open; they go out and do not return to them.
JOB|39|5|"Who has let the wild donkey go free? Who has loosed the bonds of the swift donkey,
JOB|39|6|to whom I have given the arid plain for his home and the salt land for his dwelling place?
JOB|39|7|He scorns the tumult of the city; he hears not the shouts of the driver.
JOB|39|8|He ranges the mountains as his pasture, and he searches after every green thing.
JOB|39|9|"Is the wild ox willing to serve you? Will he spend the night at your manger?
JOB|39|10|Can you bind him in the furrow with ropes, or will he harrow the valleys after you?
JOB|39|11|Will you depend on him because his strength is great, and will you leave to him your labor?
JOB|39|12|Do you have faith in him that he will return your grain and gather it to your threshing floor?
JOB|39|13|"The wings of the ostrich wave proudly, but are they the pinions and plumage of love?
JOB|39|14|For she leaves her eggs to the earth and lets them be warmed on the ground,
JOB|39|15|forgetting that a foot may crush them and that the wild beast may trample them.
JOB|39|16|She deals cruelly with her young, as if they were not hers; though her labor be in vain, yet she has no fear,
JOB|39|17|because God has made her forget wisdom and given her no share in understanding.
JOB|39|18|When she rouses herself to flee, she laughs at the horse and his rider.
JOB|39|19|"Do you give the horse his might? Do you clothe his neck with a mane?
JOB|39|20|Do you make him leap like the locust? His majestic snorting is terrifying.
JOB|39|21|He paws in the valley and exults in his strength; he goes out to meet the weapons.
JOB|39|22|He laughs at fear and is not dismayed; he does not turn back from the sword.
JOB|39|23|Upon him rattle the quiver, the flashing spear and the javelin.
JOB|39|24|With fierceness and rage he swallows the ground; he cannot stand still at the sound of the trumpet.
JOB|39|25|When the trumpet sounds, he says 'Aha!' He smells the battle from afar, the thunder of the captains, and the shouting.
JOB|39|26|"Is it by your understanding that the hawk soars and spreads his wings toward the south?
JOB|39|27|Is it at your command that the eagle mounts up and makes his nest on high?
JOB|39|28|On the rock he dwells and makes his home, on the rocky crag and stronghold.
JOB|39|29|From there he spies out the prey; his eyes behold it afar off.
JOB|39|30|His young ones suck up blood, and where the slain are, there is he."
JOB|40|1|And the LORD said to Job:
JOB|40|2|"Shall a faultfinder contend with the Almighty? He who argues with God, let him answer it."
JOB|40|3|Then Job answered the LORD and said:
JOB|40|4|"Behold, I am of small account; what shall I answer you? I lay my hand on my mouth.
JOB|40|5|I have spoken once, and I will not answer; twice, but I will proceed no further."
JOB|40|6|Then the LORD answered Job out of the whirlwind and said:
JOB|40|7|"Dress for action like a man; I will question you, and you make it known to me.
JOB|40|8|Will you even put me in the wrong? Will you condemn me that you may be in the right?
JOB|40|9|Have you an arm like God, and can you thunder with a voice like his?
JOB|40|10|"Adorn yourself with majesty and dignity; clothe yourself with glory and splendor.
JOB|40|11|Pour out the overflowings of your anger, and look on everyone who is proud and abase him.
JOB|40|12|Look on everyone who is proud and bring him low and tread down the wicked where they stand.
JOB|40|13|Hide them all in the dust together; bind their faces in the world below.
JOB|40|14|Then will I also acknowledge to you that your own right hand can save you.
JOB|40|15|"Behold, Behemoth, which I made as I made you; he eats grass like an ox.
JOB|40|16|Behold, his strength in his loins, and his power in the muscles of his belly.
JOB|40|17|He makes his tail stiff like a cedar; the sinews of his thighs are knit together.
JOB|40|18|His bones are tubes of bronze, his limbs like bars of iron.
JOB|40|19|"He is the first of the works of God; let him who made him bring near his sword!
JOB|40|20|For the mountains yield food for him where all the wild beasts play.
JOB|40|21|Under the lotus plants he lies, in the shelter of the reeds and in the marsh.
JOB|40|22|For his shade the lotus trees cover him; the willows of the brook surround him.
JOB|40|23|Behold, if the river is turbulent he is not frightened; he is confident though Jordan rushes against his mouth.
JOB|40|24|Can one take him by his eyes, or pierce his nose with a snare?
JOB|41|1|"Can you draw out Leviathan with a fishhook or press down his tongue with a cord?
JOB|41|2|Can you put a rope in his nose or pierce his jaw with a hook?
JOB|41|3|Will he make many pleas to you? Will he speak to you soft words?
JOB|41|4|Will he make a covenant with you to take him for your servant forever?
JOB|41|5|Will you play with him as with a bird, or will you put him on a leash for your girls?
JOB|41|6|Will traders bargain over him? Will they divide him up among the merchants?
JOB|41|7|Can you fill his skin with harpoons or his head with fishing spears?
JOB|41|8|Lay your hands on him; remember the battle- you will not do it again!
JOB|41|9|Behold, the hope of a man is false; he is laid low even at the sight of him.
JOB|41|10|No one is so fierce that he dares to stir him up. Who then is he who can stand before me?
JOB|41|11|Who has first given to me, that I should repay him? Whatever is under the whole heaven is mine.
JOB|41|12|"I will not keep silence concerning his limbs, or his mighty strength, or his goodly frame.
JOB|41|13|Who can strip off his outer garment? Who would come near him with a bridle?
JOB|41|14|Who can open the doors of his face? Around his teeth is terror.
JOB|41|15|His back is made of rows of shields, shut up closely as with a seal.
JOB|41|16|One is so near to another that no air can come between them.
JOB|41|17|They are joined one to another; they clasp each other and cannot be separated.
JOB|41|18|His sneezings flash forth light, and his eyes are like the eyelids of the dawn.
JOB|41|19|Out of his mouth go flaming torches; sparks of fire leap forth.
JOB|41|20|Out of his nostrils comes forth smoke, as from a boiling pot and burning rushes.
JOB|41|21|His breath kindles coals, and a flame comes forth from his mouth.
JOB|41|22|In his neck abides strength, and terror dances before him.
JOB|41|23|The folds of his flesh stick together, firmly cast on him and immovable.
JOB|41|24|His heart is hard as a stone, hard as the lower millstone.
JOB|41|25|When he raises himself up the mighty are afraid; at the crashing they are beside themselves.
JOB|41|26|Though the sword reaches him, it does not avail, nor the spear, the dart, or the javelin.
JOB|41|27|He counts iron as straw, and bronze as rotten wood.
JOB|41|28|The arrow cannot make him flee; for him sling stones are turned to stubble.
JOB|41|29|Clubs are counted as stubble; he laughs at the rattle of javelins.
JOB|41|30|His underparts are like sharp potsherds; he spreads himself like a threshing sledge on the mire.
JOB|41|31|He makes the deep boil like a pot; he makes the sea like a pot of ointment.
JOB|41|32|Behind him he leaves a shining wake; one would think the deep to be white-haired.
JOB|41|33|On earth there is not his like, a creature without fear.
JOB|41|34|He sees everything that is high; he is king over all the sons of pride."
JOB|42|1|Then Job answered the LORD and said:
JOB|42|2|"I know that you can do all things, and that no purpose of yours can be thwarted.
JOB|42|3|'Who is this that hides counsel without knowledge?' Therefore I have uttered what I did not understand, things too wonderful for me, which I did not know.
JOB|42|4|'Hear, and I will speak; I will question you, and you make it known to me.'
JOB|42|5|I had heard of you by the hearing of the ear, but now my eye sees you;
JOB|42|6|therefore I despise myself, and repent in dust and ashes."
JOB|42|7|After the LORD had spoken these words to Job, the LORD said to Eliphaz the Temanite: "My anger burns against you and against your two friends, for you have not spoken of me what is right, as my servant Job has.
JOB|42|8|Now therefore take seven bulls and seven rams and go to my servant Job and offer up a burnt offering for yourselves. And my servant Job shall pray for you, for I will accept his prayer not to deal with you according to your folly. For you have not spoken of me what is right, as my servant Job has."
JOB|42|9|So Eliphaz the Temanite and Bildad the Shuhite and Zophar the Naamathite went and did what the LORD had told them, and the LORD accepted Job's prayer.
JOB|42|10|And the LORD restored the fortunes of Job, when he had prayed for his friends. And the LORD gave Job twice as much as he had before.
JOB|42|11|Then came to him all his brothers and sisters and all who had known him before, and ate bread with him in his house. And they showed him sympathy and comforted him for all the evil that the LORD had brought upon him. And each of them gave him a piece of money and a ring of gold.
JOB|42|12|And the LORD blessed the latter days of Job more than his beginning. And he had 14,000 sheep, 6,000 camels, 1,000 yoke of oxen, and 1,000 female donkeys.
JOB|42|13|He had also seven sons and three daughters.
JOB|42|14|And he called the name of the first daughter Jemimah, and the name of the second Keziah, and the name of the third Keren-happuch.
JOB|42|15|And in all the land there were no women so beautiful as Job's daughters. And their father gave them an inheritance among their brothers.
JOB|42|16|And after this Job lived 140 years, and saw his sons, and his sons' sons, four generations.
JOB|42|17|And Job died, an old man, and full of days.
