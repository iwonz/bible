ROM|1|1|Paul, a servant of Christ Jesus, called to be an apostle and set apart for the gospel of God--
ROM|1|2|the gospel he promised beforehand through his prophets in the Holy Scriptures
ROM|1|3|regarding his Son, who as to his human nature was a descendant of David,
ROM|1|4|and who through the Spirit of holiness was declared with power to be the Son of God by his resurrection from the dead: Jesus Christ our Lord.
ROM|1|5|Through him and for his name's sake, we received grace and apostleship to call people from among all the Gentiles to the obedience that comes from faith.
ROM|1|6|And you also are among those who are called to belong to Jesus Christ.
ROM|1|7|To all in Rome who are loved by God and called to be saints: Grace and peace to you from God our Father and from the Lord Jesus Christ.
ROM|1|8|First, I thank my God through Jesus Christ for all of you, because your faith is being reported all over the world.
ROM|1|9|God, whom I serve with my whole heart in preaching the gospel of his Son, is my witness how constantly I remember you
ROM|1|10|in my prayers at all times; and I pray that now at last by God's will the way may be opened for me to come to you.
ROM|1|11|I long to see you so that I may impart to you some spiritual gift to make you strong--
ROM|1|12|that is, that you and I may be mutually encouraged by each other's faith.
ROM|1|13|I do not want you to be unaware, brothers, that I planned many times to come to you (but have been prevented from doing so until now) in order that I might have a harvest among you, just as I have had among the other Gentiles.
ROM|1|14|I am obligated both to Greeks and non-Greeks, both to the wise and the foolish.
ROM|1|15|That is why I am so eager to preach the gospel also to you who are at Rome.
ROM|1|16|I am not ashamed of the gospel, because it is the power of God for the salvation of everyone who believes: first for the Jew, then for the Gentile.
ROM|1|17|For in the gospel a righteousness from God is revealed, a righteousness that is by faith from first to last, just as it is written: "The righteous will live by faith."
ROM|1|18|The wrath of God is being revealed from heaven against all the godlessness and wickedness of men who suppress the truth by their wickedness,
ROM|1|19|since what may be known about God is plain to them, because God has made it plain to them.
ROM|1|20|For since the creation of the world God's invisible qualities--his eternal power and divine nature--have been clearly seen, being understood from what has been made, so that men are without excuse.
ROM|1|21|For although they knew God, they neither glorified him as God nor gave thanks to him, but their thinking became futile and their foolish hearts were darkened.
ROM|1|22|Although they claimed to be wise, they became fools
ROM|1|23|and exchanged the glory of the immortal God for images made to look like mortal man and birds and animals and reptiles.
ROM|1|24|Therefore God gave them over in the sinful desires of their hearts to sexual impurity for the degrading of their bodies with one another.
ROM|1|25|They exchanged the truth of God for a lie, and worshiped and served created things rather than the Creator--who is forever praised. Amen.
ROM|1|26|Because of this, God gave them over to shameful lusts. Even their women exchanged natural relations for unnatural ones.
ROM|1|27|In the same way the men also abandoned natural relations with women and were inflamed with lust for one another. Men committed indecent acts with other men, and received in themselves the due penalty for their perversion.
ROM|1|28|Furthermore, since they did not think it worthwhile to retain the knowledge of God, he gave them over to a depraved mind, to do what ought not to be done.
ROM|1|29|They have become filled with every kind of wickedness, evil, greed and depravity. They are full of envy, murder, strife, deceit and malice. They are gossips,
ROM|1|30|slanderers, God-haters, insolent, arrogant and boastful; they invent ways of doing evil; they disobey their parents;
ROM|1|31|they are senseless, faithless, heartless, ruthless.
ROM|1|32|Although they know God's righteous decree that those who do such things deserve death, they not only continue to do these very things but also approve of those who practice them.
ROM|2|1|You, therefore, have no excuse, you who pass judgment on someone else, for at whatever point you judge the other, you are condemning yourself, because you who pass judgment do the same things.
ROM|2|2|Now we know that God's judgment against those who do such things is based on truth.
ROM|2|3|So when you, a mere man, pass judgment on them and yet do the same things, do you think you will escape God's judgment?
ROM|2|4|Or do you show contempt for the riches of his kindness, tolerance and patience, not realizing that God's kindness leads you toward repentance?
ROM|2|5|But because of your stubbornness and your unrepentant heart, you are storing up wrath against yourself for the day of God's wrath, when his righteous judgment will be revealed.
ROM|2|6|God "will give to each person according to what he has done."
ROM|2|7|To those who by persistence in doing good seek glory, honor and immortality, he will give eternal life.
ROM|2|8|But for those who are self-seeking and who reject the truth and follow evil, there will be wrath and anger.
ROM|2|9|There will be trouble and distress for every human being who does evil: first for the Jew, then for the Gentile;
ROM|2|10|but glory, honor and peace for everyone who does good: first for the Jew, then for the Gentile.
ROM|2|11|For God does not show favoritism.
ROM|2|12|All who sin apart from the law will also perish apart from the law, and all who sin under the law will be judged by the law.
ROM|2|13|For it is not those who hear the law who are righteous in God's sight, but it is those who obey the law who will be declared righteous.
ROM|2|14|(Indeed, when Gentiles, who do not have the law, do by nature things required by the law, they are a law for themselves, even though they do not have the law,
ROM|2|15|since they show that the requirements of the law are written on their hearts, their consciences also bearing witness, and their thoughts now accusing, now even defending them.)
ROM|2|16|This will take place on the day when God will judge men's secrets through Jesus Christ, as my gospel declares.
ROM|2|17|Now you, if you call yourself a Jew; if you rely on the law and brag about your relationship to God;
ROM|2|18|if you know his will and approve of what is superior because you are instructed by the law;
ROM|2|19|if you are convinced that you are a guide for the blind, a light for those who are in the dark,
ROM|2|20|an instructor of the foolish, a teacher of infants, because you have in the law the embodiment of knowledge and truth--
ROM|2|21|you, then, who teach others, do you not teach yourself? You who preach against stealing, do you steal?
ROM|2|22|You who say that people should not commit adultery, do you commit adultery? You who abhor idols, do you rob temples?
ROM|2|23|You who brag about the law, do you dishonor God by breaking the law?
ROM|2|24|As it is written: "God's name is blasphemed among the Gentiles because of you."
ROM|2|25|Circumcision has value if you observe the law, but if you break the law, you have become as though you had not been circumcised.
ROM|2|26|If those who are not circumcised keep the law's requirements, will they not be regarded as though they were circumcised?
ROM|2|27|The one who is not circumcised physically and yet obeys the law will condemn you who, even though you have the written code and circumcision, are a lawbreaker.
ROM|2|28|A man is not a Jew if he is only one outwardly, nor is circumcision merely outward and physical.
ROM|2|29|No, a man is a Jew if he is one inwardly; and circumcision is circumcision of the heart, by the Spirit, not by the written code. Such a man's praise is not from men, but from God.
ROM|3|1|What advantage, then, is there in being a Jew, or what value is there in circumcision?
ROM|3|2|Much in every way! First of all, they have been entrusted with the very words of God.
ROM|3|3|What if some did not have faith? Will their lack of faith nullify God's faithfulness?
ROM|3|4|Not at all! Let God be true, and every man a liar. As it is written: "So that you may be proved right when you speak and prevail when you judge."
ROM|3|5|But if our unrighteousness brings out God's righteousness more clearly, what shall we say? That God is unjust in bringing his wrath on us? (I am using a human argument.)
ROM|3|6|Certainly not! If that were so, how could God judge the world?
ROM|3|7|Someone might argue, "If my falsehood enhances God's truthfulness and so increases his glory, why am I still condemned as a sinner?"
ROM|3|8|Why not say--as we are being slanderously reported as saying and as some claim that we say--"Let us do evil that good may result"? Their condemnation is deserved.
ROM|3|9|What shall we conclude then? Are we any better? Not at all! We have already made the charge that Jews and Gentiles alike are all under sin.
ROM|3|10|As it is written: "There is no one righteous, not even one;
ROM|3|11|there is no one who understands, no one who seeks God.
ROM|3|12|All have turned away, they have together become worthless; there is no one who does good, not even one."
ROM|3|13|"Their throats are open graves; their tongues practice deceit.The poison of vipers is on their lips."
ROM|3|14|"Their mouths are full of cursing and bitterness."
ROM|3|15|"Their feet are swift to shed blood;
ROM|3|16|ruin and misery mark their ways,
ROM|3|17|and the way of peace they do not know."
ROM|3|18|"There is no fear of God before their eyes."
ROM|3|19|Now we know that whatever the law says, it says to those who are under the law, so that every mouth may be silenced and the whole world held accountable to God.
ROM|3|20|Therefore no one will be declared righteous in his sight by observing the law; rather, through the law we become conscious of sin.
ROM|3|21|But now a righteousness from God, apart from law, has been made known, to which the Law and the Prophets testify.
ROM|3|22|This righteousness from God comes through faith in Jesus Christ to all who believe. There is no difference,
ROM|3|23|for all have sinned and fall short of the glory of God,
ROM|3|24|and are justified freely by his grace through the redemption that came by Christ Jesus.
ROM|3|25|God presented him as a sacrifice of atonement, through faith in his blood. He did this to demonstrate his justice, because in his forbearance he had left the sins committed beforehand unpunished--
ROM|3|26|he did it to demonstrate his justice at the present time, so as to be just and the one who justifies those who have faith in Jesus.
ROM|3|27|Where, then, is boasting? It is excluded. On what principle? On that of observing the law? No, but on that of faith.
ROM|3|28|For we maintain that a man is justified by faith apart from observing the law.
ROM|3|29|Is God the God of Jews only? Is he not the God of Gentiles too? Yes, of Gentiles too,
ROM|3|30|since there is only one God, who will justify the circumcised by faith and the uncircumcised through that same faith.
ROM|3|31|Do we, then, nullify the law by this faith? Not at all! Rather, we uphold the law.
ROM|4|1|What then shall we say that Abraham, our forefather, discovered in this matter?
ROM|4|2|If, in fact, Abraham was justified by works, he had something to boast about--but not before God.
ROM|4|3|What does the Scripture say? "Abraham believed God, and it was credited to him as righteousness."
ROM|4|4|Now when a man works, his wages are not credited to him as a gift, but as an obligation.
ROM|4|5|However, to the man who does not work but trusts God who justifies the wicked, his faith is credited as righteousness.
ROM|4|6|David says the same thing when he speaks of the blessedness of the man to whom God credits righteousness apart from works:
ROM|4|7|"Blessed are they whose transgressions are forgiven, whose sins are covered.
ROM|4|8|Blessed is the man whose sin the Lord will never count against him."
ROM|4|9|Is this blessedness only for the circumcised, or also for the uncircumcised? We have been saying that Abraham's faith was credited to him as righteousness.
ROM|4|10|Under what circumstances was it credited? Was it after he was circumcised, or before? It was not after, but before!
ROM|4|11|And he received the sign of circumcision, a seal of the righteousness that he had by faith while he was still uncircumcised. So then, he is the father of all who believe but have not been circumcised, in order that righteousness might be credited to them.
ROM|4|12|And he is also the father of the circumcised who not only are circumcised but who also walk in the footsteps of the faith that our father Abraham had before he was circumcised.
ROM|4|13|It was not through law that Abraham and his offspring received the promise that he would be heir of the world, but through the righteousness that comes by faith.
ROM|4|14|For if those who live by law are heirs, faith has no value and the promise is worthless,
ROM|4|15|because law brings wrath. And where there is no law there is no transgression.
ROM|4|16|Therefore, the promise comes by faith, so that it may be by grace and may be guaranteed to all Abraham's offspring--not only to those who are of the law but also to those who are of the faith of Abraham. He is the father of us all.
ROM|4|17|As it is written: "I have made you a father of many nations." He is our father in the sight of God, in whom he believed--the God who gives life to the dead and calls things that are not as though they were.
ROM|4|18|Against all hope, Abraham in hope believed and so became the father of many nations, just as it had been said to him, "So shall your offspring be."
ROM|4|19|Without weakening in his faith, he faced the fact that his body was as good as dead--since he was about a hundred years old--and that Sarah's womb was also dead.
ROM|4|20|Yet he did not waver through unbelief regarding the promise of God, but was strengthened in his faith and gave glory to God,
ROM|4|21|being fully persuaded that God had power to do what he had promised.
ROM|4|22|This is why "it was credited to him as righteousness."
ROM|4|23|The words "it was credited to him" were written not for him alone,
ROM|4|24|but also for us, to whom God will credit righteousness--for us who believe in him who raised Jesus our Lord from the dead.
ROM|4|25|He was delivered over to death for our sins and was raised to life for our justification.
ROM|5|1|Therefore, since we have been justified through faith, we have peace with God through our Lord Jesus Christ,
ROM|5|2|through whom we have gained access by faith into this grace in which we now stand. And we rejoice in the hope of the glory of God.
ROM|5|3|Not only so, but we also rejoice in our sufferings, because we know that suffering produces perseverance;
ROM|5|4|perseverance, character; and character, hope.
ROM|5|5|And hope does not disappoint us, because God has poured out his love into our hearts by the Holy Spirit, whom he has given us.
ROM|5|6|You see, at just the right time, when we were still powerless, Christ died for the ungodly.
ROM|5|7|Very rarely will anyone die for a righteous man, though for a good man someone might possibly dare to die.
ROM|5|8|But God demonstrates his own love for us in this: While we were still sinners, Christ died for us.
ROM|5|9|Since we have now been justified by his blood, how much more shall we be saved from God's wrath through him!
ROM|5|10|For if, when we were God's enemies, we were reconciled to him through the death of his Son, how much more, having been reconciled, shall we be saved through his life!
ROM|5|11|Not only is this so, but we also rejoice in God through our Lord Jesus Christ, through whom we have now received reconciliation.
ROM|5|12|Therefore, just as sin entered the world through one man, and death through sin, and in this way death came to all men, because all sinned--
ROM|5|13|for before the law was given, sin was in the world. But sin is not taken into account when there is no law.
ROM|5|14|Nevertheless, death reigned from the time of Adam to the time of Moses, even over those who did not sin by breaking a command, as did Adam, who was a pattern of the one to come.
ROM|5|15|But the gift is not like the trespass. For if the many died by the trespass of the one man, how much more did God's grace and the gift that came by the grace of the one man, Jesus Christ, overflow to the many!
ROM|5|16|Again, the gift of God is not like the result of the one man's sin: The judgment followed one sin and brought condemnation, but the gift followed many trespasses and brought justification.
ROM|5|17|For if, by the trespass of the one man, death reigned through that one man, how much more will those who receive God's abundant provision of grace and of the gift of righteousness reign in life through the one man, Jesus Christ.
ROM|5|18|Consequently, just as the result of one trespass was condemnation for all men, so also the result of one act of righteousness was justification that brings life for all men.
ROM|5|19|For just as through the disobedience of the one man the many were made sinners, so also through the obedience of the one man the many will be made righteous.
ROM|5|20|The law was added so that the trespass might increase. But where sin increased, grace increased all the more,
ROM|5|21|so that, just as sin reigned in death, so also grace might reign through righteousness to bring eternal life through Jesus Christ our Lord.
ROM|6|1|What shall we say, then? Shall we go on sinning so that grace may increase?
ROM|6|2|By no means! We died to sin; how can we live in it any longer?
ROM|6|3|Or don't you know that all of us who were baptized into Christ Jesus were baptized into his death?
ROM|6|4|We were therefore buried with him through baptism into death in order that, just as Christ was raised from the dead through the glory of the Father, we too may live a new life.
ROM|6|5|If we have been united with him like this in his death, we will certainly also be united with him in his resurrection.
ROM|6|6|For we know that our old self was crucified with him so that the body of sin might be done away with, that we should no longer be slaves to sin--
ROM|6|7|because anyone who has died has been freed from sin.
ROM|6|8|Now if we died with Christ, we believe that we will also live with him.
ROM|6|9|For we know that since Christ was raised from the dead, he cannot die again; death no longer has mastery over him.
ROM|6|10|The death he died, he died to sin once for all; but the life he lives, he lives to God.
ROM|6|11|In the same way, count yourselves dead to sin but alive to God in Christ Jesus.
ROM|6|12|Therefore do not let sin reign in your mortal body so that you obey its evil desires.
ROM|6|13|Do not offer the parts of your body to sin, as instruments of wickedness, but rather offer yourselves to God, as those who have been brought from death to life; and offer the parts of your body to him as instruments of righteousness.
ROM|6|14|For sin shall not be your master, because you are not under law, but under grace.
ROM|6|15|What then? Shall we sin because we are not under law but under grace? By no means!
ROM|6|16|Don't you know that when you offer yourselves to someone to obey him as slaves, you are slaves to the one whom you obey--whether you are slaves to sin, which leads to death, or to obedience, which leads to righteousness?
ROM|6|17|But thanks be to God that, though you used to be slaves to sin, you wholeheartedly obeyed the form of teaching to which you were entrusted.
ROM|6|18|You have been set free from sin and have become slaves to righteousness.
ROM|6|19|I put this in human terms because you are weak in your natural selves. Just as you used to offer the parts of your body in slavery to impurity and to ever-increasing wickedness, so now offer them in slavery to righteousness leading to holiness.
ROM|6|20|When you were slaves to sin, you were free from the control of righteousness.
ROM|6|21|What benefit did you reap at that time from the things you are now ashamed of? Those things result in death!
ROM|6|22|But now that you have been set free from sin and have become slaves to God, the benefit you reap leads to holiness, and the result is eternal life.
ROM|6|23|For the wages of sin is death, but the gift of God is eternal life in Christ Jesus our Lord.
ROM|7|1|Do you not know, brothers--for I am speaking to men who know the law--that the law has authority over a man only as long as he lives?
ROM|7|2|For example, by law a married woman is bound to her husband as long as he is alive, but if her husband dies, she is released from the law of marriage.
ROM|7|3|So then, if she marries another man while her husband is still alive, she is called an adulteress. But if her husband dies, she is released from that law and is not an adulteress, even though she marries another man.
ROM|7|4|So, my brothers, you also died to the law through the body of Christ, that you might belong to another, to him who was raised from the dead, in order that we might bear fruit to God.
ROM|7|5|For when we were controlled by the sinful nature, the sinful passions aroused by the law were at work in our bodies, so that we bore fruit for death.
ROM|7|6|But now, by dying to what once bound us, we have been released from the law so that we serve in the new way of the Spirit, and not in the old way of the written code.
ROM|7|7|What shall we say, then? Is the law sin? Certainly not! Indeed I would not have known what sin was except through the law. For I would not have known what coveting really was if the law had not said, "Do not covet."
ROM|7|8|But sin, seizing the opportunity afforded by the commandment, produced in me every kind of covetous desire. For apart from law, sin is dead.
ROM|7|9|Once I was alive apart from law; but when the commandment came, sin sprang to life and I died.
ROM|7|10|I found that the very commandment that was intended to bring life actually brought death.
ROM|7|11|For sin, seizing the opportunity afforded by the commandment, deceived me, and through the commandment put me to death.
ROM|7|12|So then, the law is holy, and the commandment is holy, righteous and good.
ROM|7|13|Did that which is good, then, become death to me? By no means! But in order that sin might be recognized as sin, it produced death in me through what was good, so that through the commandment sin might become utterly sinful.
ROM|7|14|We know that the law is spiritual; but I am unspiritual, sold as a slave to sin.
ROM|7|15|I do not understand what I do. For what I want to do I do not do, but what I hate I do.
ROM|7|16|And if I do what I do not want to do, I agree that the law is good.
ROM|7|17|As it is, it is no longer I myself who do it, but it is sin living in me.
ROM|7|18|I know that nothing good lives in me, that is, in my sinful nature. For I have the desire to do what is good, but I cannot carry it out.
ROM|7|19|For what I do is not the good I want to do; no, the evil I do not want to do--this I keep on doing.
ROM|7|20|Now if I do what I do not want to do, it is no longer I who do it, but it is sin living in me that does it.
ROM|7|21|So I find this law at work: When I want to do good, evil is right there with me.
ROM|7|22|For in my inner being I delight in God's law;
ROM|7|23|but I see another law at work in the members of my body, waging war against the law of my mind and making me a prisoner of the law of sin at work within my members.
ROM|7|24|What a wretched man I am! Who will rescue me from this body of death?
ROM|7|25|Thanks be to God--through Jesus Christ our Lord! So then, I myself in my mind am a slave to God's law, but in the sinful nature a slave to the law of sin.
ROM|8|1|Therefore, there is now no condemnation for those who are in Christ Jesus,
ROM|8|2|because through Christ Jesus the law of the Spirit of life set me free from the law of sin and death.
ROM|8|3|For what the law was powerless to do in that it was weakened by the sinful nature, God did by sending his own Son in the likeness of sinful man to be a sin offering. And so he condemned sin in sinful man,
ROM|8|4|in order that the righteous requirements of the law might be fully met in us, who do not live according to the sinful nature but according to the Spirit.
ROM|8|5|Those who live according to the sinful nature have their minds set on what that nature desires; but those who live in accordance with the Spirit have their minds set on what the Spirit desires.
ROM|8|6|The mind of sinful man is death, but the mind controlled by the Spirit is life and peace;
ROM|8|7|the sinful mind is hostile to God. It does not submit to God's law, nor can it do so.
ROM|8|8|Those controlled by the sinful nature cannot please God.
ROM|8|9|You, however, are controlled not by the sinful nature but by the Spirit, if the Spirit of God lives in you. And if anyone does not have the Spirit of Christ, he does not belong to Christ.
ROM|8|10|But if Christ is in you, your body is dead because of sin, yet your spirit is alive because of righteousness.
ROM|8|11|And if the Spirit of him who raised Jesus from the dead is living in you, he who raised Christ from the dead will also give life to your mortal bodies through his Spirit, who lives in you.
ROM|8|12|Therefore, brothers, we have an obligation--but it is not to the sinful nature, to live according to it.
ROM|8|13|For if you live according to the sinful nature, you will die; but if by the Spirit you put to death the misdeeds of the body, you will live,
ROM|8|14|because those who are led by the Spirit of God are sons of God.
ROM|8|15|For you did not receive a spirit that makes you a slave again to fear, but you received the Spirit of sonship. And by him we cry, "Abba, Father."
ROM|8|16|The Spirit himself testifies with our spirit that we are God's children.
ROM|8|17|Now if we are children, then we are heirs--heirs of God and co-heirs with Christ, if indeed we share in his sufferings in order that we may also share in his glory.
ROM|8|18|I consider that our present sufferings are not worth comparing with the glory that will be revealed in us.
ROM|8|19|The creation waits in eager expectation for the sons of God to be revealed.
ROM|8|20|For the creation was subjected to frustration, not by its own choice, but by the will of the one who subjected it, in hope
ROM|8|21|that the creation itself will be liberated from its bondage to decay and brought into the glorious freedom of the children of God.
ROM|8|22|We know that the whole creation has been groaning as in the pains of childbirth right up to the present time.
ROM|8|23|Not only so, but we ourselves, who have the firstfruits of the Spirit, groan inwardly as we wait eagerly for our adoption as sons, the redemption of our bodies.
ROM|8|24|For in this hope we were saved. But hope that is seen is no hope at all. Who hopes for what he already has?
ROM|8|25|But if we hope for what we do not yet have, we wait for it patiently.
ROM|8|26|In the same way, the Spirit helps us in our weakness. We do not know what we ought to pray for, but the Spirit himself intercedes for us with groans that words cannot express.
ROM|8|27|And he who searches our hearts knows the mind of the Spirit, because the Spirit intercedes for the saints in accordance with God's will.
ROM|8|28|And we know that in all things God works for the good of those who love him, who have been called according to his purpose.
ROM|8|29|For those God foreknew he also predestined to be conformed to the likeness of his Son, that he might be the firstborn among many brothers.
ROM|8|30|And those he predestined, he also called; those he called, he also justified; those he justified, he also glorified.
ROM|8|31|What, then, shall we say in response to this? If God is for us, who can be against us?
ROM|8|32|He who did not spare his own Son, but gave him up for us all--how will he not also, along with him, graciously give us all things?
ROM|8|33|Who will bring any charge against those whom God has chosen? It is God who justifies.
ROM|8|34|Who is he that condemns? Christ Jesus, who died--more than that, who was raised to life--is at the right hand of God and is also interceding for us.
ROM|8|35|Who shall separate us from the love of Christ? Shall trouble or hardship or persecution or famine or nakedness or danger or sword?
ROM|8|36|As it is written: "For your sake we face death all day long; we are considered as sheep to be slaughtered."
ROM|8|37|No, in all these things we are more than conquerors through him who loved us.
ROM|8|38|For I am convinced that neither death nor life, neither angels nor demons, neither the present nor the future, nor any powers,
ROM|8|39|neither height nor depth, nor anything else in all creation, will be able to separate us from the love of God that is in Christ Jesus our Lord.
ROM|9|1|I speak the truth in Christ--I am not lying, my conscience confirms it in the Holy Spirit--
ROM|9|2|I have great sorrow and unceasing anguish in my heart.
ROM|9|3|For I could wish that I myself were cursed and cut off from Christ for the sake of my brothers, those of my own race,
ROM|9|4|the people of Israel. Theirs is the adoption as sons; theirs the divine glory, the covenants, the receiving of the law, the temple worship and the promises.
ROM|9|5|Theirs are the patriarchs, and from them is traced the human ancestry of Christ, who is God over all, forever praised! Amen.
ROM|9|6|It is not as though God's word had failed. For not all who are descended from Israel are Israel.
ROM|9|7|Nor because they are his descendants are they all Abraham's children. On the contrary, "It is through Isaac that your offspring will be reckoned."
ROM|9|8|In other words, it is not the natural children who are God's children, but it is the children of the promise who are regarded as Abraham's offspring.
ROM|9|9|For this was how the promise was stated: "At the appointed time I will return, and Sarah will have a son."
ROM|9|10|Not only that, but Rebekah's children had one and the same father, our father Isaac.
ROM|9|11|Yet, before the twins were born or had done anything good or bad--in order that God's purpose in election might stand:
ROM|9|12|not by works but by him who calls--she was told, "The older will serve the younger."
ROM|9|13|Just as it is written: "Jacob I loved, but Esau I hated."
ROM|9|14|What then shall we say? Is God unjust? Not at all!
ROM|9|15|For he says to Moses, "I will have mercy on whom I have mercy, and I will have compassion on whom I have compassion."
ROM|9|16|It does not, therefore, depend on man's desire or effort, but on God's mercy.
ROM|9|17|For the Scripture says to Pharaoh: "I raised you up for this very purpose, that I might display my power in you and that my name might be proclaimed in all the earth."
ROM|9|18|Therefore God has mercy on whom he wants to have mercy, and he hardens whom he wants to harden.
ROM|9|19|One of you will say to me: "Then why does God still blame us? For who resists his will?"
ROM|9|20|But who are you, O man, to talk back to God? "Shall what is formed say to him who formed it, 'Why did you make me like this?'"
ROM|9|21|Does not the potter have the right to make out of the same lump of clay some pottery for noble purposes and some for common use?
ROM|9|22|What if God, choosing to show his wrath and make his power known, bore with great patience the objects of his wrath--prepared for destruction?
ROM|9|23|What if he did this to make the riches of his glory known to the objects of his mercy, whom he prepared in advance for glory--
ROM|9|24|even us, whom he also called, not only from the Jews but also from the Gentiles?
ROM|9|25|As he says in Hosea: "I will call them 'my people' who are not my people; and I will call her 'my loved one' who is not my loved one,"
ROM|9|26|and, "It will happen that in the very place where it was said to them, 'You are not my people,' they will be called 'sons of the living God.'"
ROM|9|27|Isaiah cries out concerning Israel: "Though the number of the Israelites be like the sand by the sea, only the remnant will be saved.
ROM|9|28|For the Lord will carry out his sentence on earth with speed and finality."
ROM|9|29|It is just as Isaiah said previously: "Unless the Lord Almighty had left us descendants, we would have become like Sodom, we would have been like Gomorrah."
ROM|9|30|What then shall we say? That the Gentiles, who did not pursue righteousness, have obtained it, a righteousness that is by faith;
ROM|9|31|but Israel, who pursued a law of righteousness, has not attained it.
ROM|9|32|Why not? Because they pursued it not by faith but as if it were by works. They stumbled over the "stumbling stone."
ROM|9|33|As it is written: "See, I lay in Zion a stone that causes men to stumble and a rock that makes them fall, and the one who trusts in him will never be put to shame."
ROM|10|1|Brothers, my heart's desire and prayer to God for the Israelites is that they may be saved.
ROM|10|2|For I can testify about them that they are zealous for God, but their zeal is not based on knowledge.
ROM|10|3|Since they did not know the righteousness that comes from God and sought to establish their own, they did not submit to God's righteousness.
ROM|10|4|Christ is the end of the law so that there may be righteousness for everyone who believes.
ROM|10|5|Moses describes in this way the righteousness that is by the law: "The man who does these things will live by them."
ROM|10|6|But the righteousness that is by faith says: "Do not say in your heart, 'Who will ascend into heaven?'" (that is, to bring Christ down)
ROM|10|7|"or 'Who will descend into the deep?'" (that is, to bring Christ up from the dead).
ROM|10|8|But what does it say? "The word is near you; it is in your mouth and in your heart," that is, the word of faith we are proclaiming:
ROM|10|9|That if you confess with your mouth, "Jesus is Lord," and believe in your heart that God raised him from the dead, you will be saved.
ROM|10|10|For it is with your heart that you believe and are justified, and it is with your mouth that you confess and are saved.
ROM|10|11|As the Scripture says, "Anyone who trusts in him will never be put to shame."
ROM|10|12|For there is no difference between Jew and Gentile--the same Lord is Lord of all and richly blesses all who call on him,
ROM|10|13|for, "Everyone who calls on the name of the Lord will be saved."
ROM|10|14|How, then, can they call on the one they have not believed in? And how can they believe in the one of whom they have not heard? And how can they hear without someone preaching to them?
ROM|10|15|And how can they preach unless they are sent? As it is written, "How beautiful are the feet of those who bring good news!"
ROM|10|16|But not all the Israelites accepted the good news. For Isaiah says, "Lord, who has believed our message?"
ROM|10|17|Consequently, faith comes from hearing the message, and the message is heard through the word of Christ.
ROM|10|18|But I ask: Did they not hear? Of course they did: "Their voice has gone out into all the earth, their words to the ends of the world."
ROM|10|19|Again I ask: Did Israel not understand? First, Moses says, "I will make you envious by those who are not a nation; I will make you angry by a nation that has no understanding."
ROM|10|20|And Isaiah boldly says, "I was found by those who did not seek me; I revealed myself to those who did not ask for me."
ROM|10|21|But concerning Israel he says, "All day long I have held out my hands to a disobedient and obstinate people."
ROM|11|1|I ask then: Did God reject his people? By no means! I am an Israelite myself, a descendant of Abraham, from the tribe of Benjamin.
ROM|11|2|God did not reject his people, whom he foreknew. Don't you know what the Scripture says in the passage about Elijah--how he appealed to God against Israel:
ROM|11|3|"Lord, they have killed your prophets and torn down your altars; I am the only one left, and they are trying to kill me"?
ROM|11|4|And what was God's answer to him? "I have reserved for myself seven thousand who have not bowed the knee to Baal."
ROM|11|5|So too, at the present time there is a remnant chosen by grace.
ROM|11|6|And if by grace, then it is no longer by works; if it were, grace would no longer be grace.
ROM|11|7|What then? What Israel sought so earnestly it did not obtain, but the elect did. The others were hardened,
ROM|11|8|as it is written: "God gave them a spirit of stupor, eyes so that they could not see and ears so that they could not hear, to this very day."
ROM|11|9|And David says: "May their table become a snare and a trap, a stumbling block and a retribution for them.
ROM|11|10|May their eyes be darkened so they cannot see, and their backs be bent forever."
ROM|11|11|Again I ask: Did they stumble so as to fall beyond recovery? Not at all! Rather, because of their transgression, salvation has come to the Gentiles to make Israel envious.
ROM|11|12|But if their transgression means riches for the world, and their loss means riches for the Gentiles, how much greater riches will their fullness bring!
ROM|11|13|I am talking to you Gentiles. Inasmuch as I am the apostle to the Gentiles, I make much of my ministry
ROM|11|14|in the hope that I may somehow arouse my own people to envy and save some of them.
ROM|11|15|For if their rejection is the reconciliation of the world, what will their acceptance be but life from the dead?
ROM|11|16|If the part of the dough offered as firstfruits is holy, then the whole batch is holy; if the root is holy, so are the branches.
ROM|11|17|If some of the branches have been broken off, and you, though a wild olive shoot, have been grafted in among the others and now share in the nourishing sap from the olive root,
ROM|11|18|do not boast over those branches. If you do, consider this: You do not support the root, but the root supports you.
ROM|11|19|You will say then, "Branches were broken off so that I could be grafted in."
ROM|11|20|Granted. But they were broken off because of unbelief, and you stand by faith. Do not be arrogant, but be afraid.
ROM|11|21|For if God did not spare the natural branches, he will not spare you either.
ROM|11|22|Consider therefore the kindness and sternness of God: sternness to those who fell, but kindness to you, provided that you continue in his kindness. Otherwise, you also will be cut off.
ROM|11|23|And if they do not persist in unbelief, they will be grafted in, for God is able to graft them in again.
ROM|11|24|After all, if you were cut out of an olive tree that is wild by nature, and contrary to nature were grafted into a cultivated olive tree, how much more readily will these, the natural branches, be grafted into their own olive tree!
ROM|11|25|I do not want you to be ignorant of this mystery, brothers, so that you may not be conceited: Israel has experienced a hardening in part until the full number of the Gentiles has come in.
ROM|11|26|And so all Israel will be saved, as it is written: "The deliverer will come from Zion; he will turn godlessness away from Jacob.
ROM|11|27|And this is my covenant with them when I take away their sins."
ROM|11|28|As far as the gospel is concerned, they are enemies on your account; but as far as election is concerned, they are loved on account of the patriarchs,
ROM|11|29|for God's gifts and his call are irrevocable.
ROM|11|30|Just as you who were at one time disobedient to God have now received mercy as a result of their disobedience,
ROM|11|31|so they too have now become disobedient in order that they too may now receive mercy as a result of God's mercy to you.
ROM|11|32|For God has bound all men over to disobedience so that he may have mercy on them all.
ROM|11|33|Oh, the depth of the riches of the wisdom and knowledge of God! How unsearchable his judgments, and his paths beyond tracing out!
ROM|11|34|"Who has known the mind of the Lord? Or who has been his counselor?"
ROM|11|35|"Who has ever given to God, that God should repay him?"
ROM|11|36|For from him and through him and to him are all things. To him be the glory forever! Amen.
ROM|12|1|Therefore, I urge you, brothers, in view of God's mercy, to offer your bodies as living sacrifices, holy and pleasing to God--this is your spiritual act of worship.
ROM|12|2|Do not conform any longer to the pattern of this world, but be transformed by the renewing of your mind. Then you will be able to test and approve what God's will is--his good, pleasing and perfect will.
ROM|12|3|For by the grace given me I say to every one of you: Do not think of yourself more highly than you ought, but rather think of yourself with sober judgment, in accordance with the measure of faith God has given you.
ROM|12|4|Just as each of us has one body with many members, and these members do not all have the same function,
ROM|12|5|so in Christ we who are many form one body, and each member belongs to all the others.
ROM|12|6|We have different gifts, according to the grace given us. If a man's gift is prophesying, let him use it in proportion to his faith.
ROM|12|7|If it is serving, let him serve; if it is teaching, let him teach;
ROM|12|8|if it is encouraging, let him encourage; if it is contributing to the needs of others, let him give generously; if it is leadership, let him govern diligently; if it is showing mercy, let him do it cheerfully.
ROM|12|9|Love must be sincere. Hate what is evil; cling to what is good.
ROM|12|10|Be devoted to one another in brotherly love. Honor one another above yourselves.
ROM|12|11|Never be lacking in zeal, but keep your spiritual fervor, serving the Lord.
ROM|12|12|Be joyful in hope, patient in affliction, faithful in prayer.
ROM|12|13|Share with God's people who are in need. Practice hospitality.
ROM|12|14|Bless those who persecute you; bless and do not curse.
ROM|12|15|Rejoice with those who rejoice; mourn with those who mourn.
ROM|12|16|Live in harmony with one another. Do not be proud, but be willing to associate with people of low position. Do not be conceited.
ROM|12|17|Do not repay anyone evil for evil. Be careful to do what is right in the eyes of everybody.
ROM|12|18|If it is possible, as far as it depends on you, live at peace with everyone.
ROM|12|19|Do not take revenge, my friends, but leave room for God's wrath, for it is written: "It is mine to avenge; I will repay," says the Lord.
ROM|12|20|On the contrary: "If your enemy is hungry, feed him; if he is thirsty, give him something to drink. In doing this, you will heap burning coals on his head."
ROM|12|21|Do not be overcome by evil, but overcome evil with good.
ROM|13|1|Everyone must submit himself to the governing authorities, for there is no authority except that which God has established. The authorities that exist have been established by God.
ROM|13|2|Consequently, he who rebels against the authority is rebelling against what God has instituted, and those who do so will bring judgment on themselves.
ROM|13|3|For rulers hold no terror for those who do right, but for those who do wrong. Do you want to be free from fear of the one in authority? Then do what is right and he will commend you.
ROM|13|4|For he is God's servant to do you good. But if you do wrong, be afraid, for he does not bear the sword for nothing. He is God's servant, an agent of wrath to bring punishment on the wrongdoer.
ROM|13|5|Therefore, it is necessary to submit to the authorities, not only because of possible punishment but also because of conscience.
ROM|13|6|This is also why you pay taxes, for the authorities are God's servants, who give their full time to governing.
ROM|13|7|Give everyone what you owe him: If you owe taxes, pay taxes; if revenue, then revenue; if respect, then respect; if honor, then honor.
ROM|13|8|Let no debt remain outstanding, except the continuing debt to love one another, for he who loves his fellowman has fulfilled the law.
ROM|13|9|The commandments, "Do not commit adultery,Do not murder,Do not steal,Do not covet," and whatever other commandment there may be, are summed up in this one rule: "Love your neighbor as yourself."
ROM|13|10|Love does no harm to its neighbor. Therefore love is the fulfillment of the law.
ROM|13|11|And do this, understanding the present time. The hour has come for you to wake up from your slumber, because our salvation is nearer now than when we first believed.
ROM|13|12|The night is nearly over; the day is almost here. So let us put aside the deeds of darkness and put on the armor of light.
ROM|13|13|Let us behave decently, as in the daytime, not in orgies and drunkenness, not in sexual immorality and debauchery, not in dissension and jealousy.
ROM|13|14|Rather, clothe yourselves with the Lord Jesus Christ, and do not think about how to gratify the desires of the sinful nature.
ROM|14|1|Accept him whose faith is weak, without passing judgment on disputable matters.
ROM|14|2|One man's faith allows him to eat everything, but another man, whose faith is weak, eats only vegetables.
ROM|14|3|The man who eats everything must not look down on him who does not, and the man who does not eat everything must not condemn the man who does, for God has accepted him.
ROM|14|4|Who are you to judge someone else's servant? To his own master he stands or falls. And he will stand, for the Lord is able to make him stand.
ROM|14|5|One man considers one day more sacred than another; another man considers every day alike. Each one should be fully convinced in his own mind.
ROM|14|6|He who regards one day as special, does so to the Lord. He who eats meat, eats to the Lord, for he gives thanks to God; and he who abstains, does so to the Lord and gives thanks to God.
ROM|14|7|For none of us lives to himself alone and none of us dies to himself alone.
ROM|14|8|If we live, we live to the Lord; and if we die, we die to the Lord. So, whether we live or die, we belong to the Lord.
ROM|14|9|For this very reason, Christ died and returned to life so that he might be the Lord of both the dead and the living.
ROM|14|10|You, then, why do you judge your brother? Or why do you look down on your brother? For we will all stand before God's judgment seat.
ROM|14|11|It is written: "'As surely as I live,' says the Lord, 'every knee will bow before me; every tongue will confess to God.'"
ROM|14|12|So then, each of us will give an account of himself to God.
ROM|14|13|Therefore let us stop passing judgment on one another. Instead, make up your mind not to put any stumbling block or obstacle in your brother's way.
ROM|14|14|As one who is in the Lord Jesus, I am fully convinced that no food is unclean in itself. But if anyone regards something as unclean, then for him it is unclean.
ROM|14|15|If your brother is distressed because of what you eat, you are no longer acting in love. Do not by your eating destroy your brother for whom Christ died.
ROM|14|16|Do not allow what you consider good to be spoken of as evil.
ROM|14|17|For the kingdom of God is not a matter of eating and drinking, but of righteousness, peace and joy in the Holy Spirit,
ROM|14|18|because anyone who serves Christ in this way is pleasing to God and approved by men.
ROM|14|19|Let us therefore make every effort to do what leads to peace and to mutual edification.
ROM|14|20|Do not destroy the work of God for the sake of food. All food is clean, but it is wrong for a man to eat anything that causes someone else to stumble.
ROM|14|21|It is better not to eat meat or drink wine or to do anything else that will cause your brother to fall.
ROM|14|22|So whatever you believe about these things keep between yourself and God. Blessed is the man who does not condemn himself by what he approves.
ROM|14|23|But the man who has doubts is condemned if he eats, because his eating is not from faith; and everything that does not come from faith is sin.
ROM|15|1|We who are strong ought to bear with the failings of the weak and not to please ourselves.
ROM|15|2|Each of us should please his neighbor for his good, to build him up.
ROM|15|3|For even Christ did not please himself but, as it is written: "The insults of those who insult you have fallen on me."
ROM|15|4|For everything that was written in the past was written to teach us, so that through endurance and the encouragement of the Scriptures we might have hope.
ROM|15|5|May the God who gives endurance and encouragement give you a spirit of unity among yourselves as you follow Christ Jesus,
ROM|15|6|so that with one heart and mouth you may glorify the God and Father of our Lord Jesus Christ.
ROM|15|7|Accept one another, then, just as Christ accepted you, in order to bring praise to God.
ROM|15|8|For I tell you that Christ has become a servant of the Jews on behalf of God's truth, to confirm the promises made to the patriarchs
ROM|15|9|so that the Gentiles may glorify God for his mercy, as it is written: "Therefore I will praise you among the Gentiles; I will sing hymns to your name."
ROM|15|10|Again, it says, "Rejoice, O Gentiles, with his people."
ROM|15|11|And again, "Praise the Lord, all you Gentiles, and sing praises to him, all you peoples."
ROM|15|12|And again, Isaiah says, "The Root of Jesse will spring up, one who will arise to rule over the nations; the Gentiles will hope in him."
ROM|15|13|May the God of hope fill you with all joy and peace as you trust in him, so that you may overflow with hope by the power of the Holy Spirit.
ROM|15|14|I myself am convinced, my brothers, that you yourselves are full of goodness, complete in knowledge and competent to instruct one another.
ROM|15|15|I have written you quite boldly on some points, as if to remind you of them again, because of the grace God gave me
ROM|15|16|to be a minister of Christ Jesus to the Gentiles with the priestly duty of proclaiming the gospel of God, so that the Gentiles might become an offering acceptable to God, sanctified by the Holy Spirit.
ROM|15|17|Therefore I glory in Christ Jesus in my service to God.
ROM|15|18|I will not venture to speak of anything except what Christ has accomplished through me in leading the Gentiles to obey God by what I have said and done--
ROM|15|19|by the power of signs and miracles, through the power of the Spirit. So from Jerusalem all the way around to Illyricum, I have fully proclaimed the gospel of Christ.
ROM|15|20|It has always been my ambition to preach the gospel where Christ was not known, so that I would not be building on someone else's foundation.
ROM|15|21|Rather, as it is written: "Those who were not told about him will see, and those who have not heard will understand."
ROM|15|22|This is why I have often been hindered from coming to you.
ROM|15|23|But now that there is no more place for me to work in these regions, and since I have been longing for many years to see you,
ROM|15|24|I plan to do so when I go to Spain. I hope to visit you while passing through and to have you assist me on my journey there, after I have enjoyed your company for a while.
ROM|15|25|Now, however, I am on my way to Jerusalem in the service of the saints there.
ROM|15|26|For Macedonia and Achaia were pleased to make a contribution for the poor among the saints in Jerusalem.
ROM|15|27|They were pleased to do it, and indeed they owe it to them. For if the Gentiles have shared in the Jews' spiritual blessings, they owe it to the Jews to share with them their material blessings.
ROM|15|28|So after I have completed this task and have made sure that they have received this fruit, I will go to Spain and visit you on the way.
ROM|15|29|I know that when I come to you, I will come in the full measure of the blessing of Christ.
ROM|15|30|I urge you, brothers, by our Lord Jesus Christ and by the love of the Spirit, to join me in my struggle by praying to God for me.
ROM|15|31|Pray that I may be rescued from the unbelievers in Judea and that my service in Jerusalem may be acceptable to the saints there,
ROM|15|32|so that by God's will I may come to you with joy and together with you be refreshed.
ROM|15|33|The God of peace be with you all. Amen.
ROM|16|1|I commend to you our sister Phoebe, a servant of the church in Cenchrea.
ROM|16|2|I ask you to receive her in the Lord in a way worthy of the saints and to give her any help she may need from you, for she has been a great help to many people, including me.
ROM|16|3|Greet Priscilla and Aquila, my fellow workers in Christ Jesus.
ROM|16|4|They risked their lives for me. Not only I but all the churches of the Gentiles are grateful to them.
ROM|16|5|Greet also the church that meets at their house. Greet my dear friend Epenetus, who was the first convert to Christ in the province of Asia.
ROM|16|6|Greet Mary, who worked very hard for you.
ROM|16|7|Greet Andronicus and Junias, my relatives who have been in prison with me. They are outstanding among the apostles, and they were in Christ before I was.
ROM|16|8|Greet Ampliatus, whom I love in the Lord.
ROM|16|9|Greet Urbanus, our fellow worker in Christ, and my dear friend Stachys.
ROM|16|10|Greet Apelles, tested and approved in Christ. Greet those who belong to the household of Aristobulus.
ROM|16|11|Greet Herodion, my relative. Greet those in the household of Narcissus who are in the Lord.
ROM|16|12|Greet Tryphena and Tryphosa, those women who work hard in the Lord. Greet my dear friend Persis, another woman who has worked very hard in the Lord.
ROM|16|13|Greet Rufus, chosen in the Lord, and his mother, who has been a mother to me, too.
ROM|16|14|Greet Asyncritus, Phlegon, Hermes, Patrobas, Hermas and the brothers with them.
ROM|16|15|Greet Philologus, Julia, Nereus and his sister, and Olympas and all the saints with them.
ROM|16|16|Greet one another with a holy kiss. All the churches of Christ send greetings.
ROM|16|17|I urge you, brothers, to watch out for those who cause divisions and put obstacles in your way that are contrary to the teaching you have learned. Keep away from them.
ROM|16|18|For such people are not serving our Lord Christ, but their own appetites. By smooth talk and flattery they deceive the minds of naive people.
ROM|16|19|Everyone has heard about your obedience, so I am full of joy over you; but I want you to be wise about what is good, and innocent about what is evil.
ROM|16|20|The God of peace will soon crush Satan under your feet. The grace of our Lord Jesus be with you.
ROM|16|21|Timothy, my fellow worker, sends his greetings to you, as do Lucius, Jason and Sosipater, my relatives.
ROM|16|22|I, Tertius, who wrote down this letter, greet you in the Lord.
ROM|16|23|Gaius, whose hospitality I and the whole church here enjoy, sends you his greetings. Erastus, who is the city's director of public works, and our brother Quartus send you their greetings.
ROM|16|24|See Footnote
ROM|16|25|Now to him who is able to establish you by my gospel and the proclamation of Jesus Christ, according to the revelation of the mystery hidden for long ages past,
ROM|16|26|but now revealed and made known through the prophetic writings by the command of the eternal God, so that all nations might believe and obey him--
ROM|16|27|to the only wise God be glory forever through Jesus Christ! Amen.
