1JOHN|1|1|论到从起初原有的生命之道，就是我们所听见、所看见、亲眼看过、亲手摸过的－
1JOHN|1|2|这生命已经显现出来，我们看见了，现在又作见证，把原与父同在，并且向我们显现过的那永远的生命传扬给你们－
1JOHN|1|3|我们把所看见、所听见的传扬给你们，为要使你们也与我们有团契，而我们的团契是与父和他儿子耶稣基督所共有的。
1JOHN|1|4|我们把这些事写给你们，使我们 的喜乐得以满足。
1JOHN|1|5|上帝就是光，在他毫无黑暗；这是我们从主所听见，又报给你们的信息。
1JOHN|1|6|我们若说，我们与上帝有团契，却仍在黑暗里行走，就是说谎话，不实行真理了。
1JOHN|1|7|我们若在光明中行走，如同上帝在光明中，就彼此有团契，他儿子耶稣的血就洗净我们一切的罪。
1JOHN|1|8|我们若说自己没有罪，就是欺骗自己，真理就不在我们里面了。
1JOHN|1|9|我们若认自己的罪，上帝是信实的，是公义的，必要赦免我们的罪，洗净我们一切的不义。
1JOHN|1|10|我们若说自己没有犯过罪，就是把上帝当作说谎的，他的道就不在我们里面了。
1JOHN|2|1|我的孩子们哪，我把这些话写给你们，是要你们不犯罪。若有人犯罪，在父那里我们有一位中保，就是那义者耶稣基督。
1JOHN|2|2|他为我们的罪作了赎罪祭，不单是为我们的罪，也是为普天下人的罪。
1JOHN|2|3|我们若遵守上帝的命令，就知道我们确实认识他。
1JOHN|2|4|人若说“我认识他”，却不遵守他的命令，就是说谎话的，真理就不在他里面了。
1JOHN|2|5|凡遵守他的道的，爱上帝的心确实地在他里面达到完全了。由此我们知道我们是在他里面。
1JOHN|2|6|凡说自己住在他里面的，就该照着他所行的去行。
1JOHN|2|7|亲爱的，我写给你们的不是一条新命令，而是你们从起初所受的旧命令；这旧命令就是你们所听过的道。
1JOHN|2|8|然而，我写给你们的是一条新命令，在基督里是真实的，在你们也是真实的，因为黑暗渐渐消逝，真光已经在照耀。
1JOHN|2|9|人若说自己在光明中，却恨他的弟兄，他到如今还是在黑暗里。
1JOHN|2|10|那爱弟兄的，就是住在光明中，他不会使人失足犯罪 。
1JOHN|2|11|惟独那恨弟兄的，是在黑暗里，也在黑暗里行走，不知道往哪里去，因为黑暗使他的眼睛瞎了。
1JOHN|2|12|孩子们哪，我写信给你们， 因为你们的罪藉着基督的名得了赦免。
1JOHN|2|13|父老们啊，我写信给你们， 因为你们认识从起初就有的那一位。 青年们哪，我写信给你们， 因为你们胜过了那恶者。
1JOHN|2|14|孩子们哪，我曾写信给你们， 因为你们认识父。 父老们啊，我曾写信给你们， 因为你们认识从起初就有的那一位。 青年们哪，我曾写信给你们， 因为你们刚强， 上帝的道常存在你们心里， 你们也胜过了那恶者。
1JOHN|2|15|不要爱世界和世界上的东西，若有人爱世界，爱父的心就不在他里面了。
1JOHN|2|16|因为凡世界上的东西，好比肉体的情欲、眼目的情欲和今生的骄傲，都不是从父来的，而是从世界来的。
1JOHN|2|17|这世界和世上的情欲都要消逝，惟独那遵行上帝旨意的人永远常存。
1JOHN|2|18|孩子们哪，如今是末世的时光了。你们曾听过那敌基督者要来，现在有好些敌基督者已经出来了；由此我们就知道，如今是末世的时光了。
1JOHN|2|19|他们从我们中间出去，却不是属我们的，若是属我们的，就必仍旧与我们同在。他们出去，这就显明他们都不是属我们的。
1JOHN|2|20|你们从那圣者受了恩膏，并且你们大家都知道 。
1JOHN|2|21|我写信给你们，不是因你们不认识真理，而是因你们认识，并且知道一切虚谎都不是从真理出来的。
1JOHN|2|22|谁是说谎话的呢？不就是那不认耶稣为基督的吗？那不认父与子的，这个人就是敌基督的。
1JOHN|2|23|凡不认子的，就没有父；宣认子的，连父也有了。
1JOHN|2|24|论到你们，务要将那从起初所听见的常存在心里；若将从起初所听见的存在心里，你们就会住在子里面，也会住在父里面。
1JOHN|2|25|基督所应许我们的就是永生。
1JOHN|2|26|我将这些话写给你们，是论到那些迷惑你们的人说的。
1JOHN|2|27|至于你们，你们从基督所受的恩膏常存在你们心里，并不用人教导你们，自有他的恩膏在凡事上教导你们。这恩膏是真的，不是假的，你们要按这恩膏的教导住在他里面。
1JOHN|2|28|孩子们哪，你们要住在基督里面。这样，他若显现，我们就可以坦然无惧；当他来临的时候，在他面前不至于惭愧。
1JOHN|2|29|你们若知道他是公义的，就知道凡行公义的人都是他所生的。
1JOHN|3|1|你们看父赐给我们的是何等的慈爱，让我们得以称为上帝的儿女；我们也真是他的儿女。世人不认识我们 的理由，是因他们未曾认识父。
1JOHN|3|2|亲爱的，我们现在是上帝的儿女，将来如何还未显明。我们所知道的是：基督显现的时候，我们会像他，因为我们将见到他的本相。
1JOHN|3|3|凡对他有这指望的，就洁净自己，像他是洁净的一样。
1JOHN|3|4|凡犯罪的，就是做违背律法的事；违背律法就是罪。
1JOHN|3|5|你们知道，基督曾显现是要除掉罪 ；在他并没有罪。
1JOHN|3|6|凡住在他里面的，不犯罪；凡犯罪的，未曾看见他，也未曾认识他。
1JOHN|3|7|孩子们哪，不要让人迷惑了你们；行义的才是义人，正如基督是义的。
1JOHN|3|8|犯罪的是出于魔鬼，因为魔鬼从起初就犯罪。上帝的儿子显现出来，是为了要毁灭魔鬼的作为。
1JOHN|3|9|凡从上帝生的，不犯罪，因上帝的道 存在他里面，他也不能犯罪，因为他是由上帝所生的。
1JOHN|3|10|这就显明谁是上帝的儿女，谁是魔鬼的儿女了。凡不行义的，不是出于上帝，不爱他弟兄的，也是如此。
1JOHN|3|11|我们要彼此相爱。这就是你们从起初所听到的信息。
1JOHN|3|12|不要像 该隐 ；他是属那邪恶者，杀了自己的弟弟。为什么杀了他呢？因为自己的行为是邪恶的，而弟弟的行为是正直的。
1JOHN|3|13|弟兄们，世人若恨你们，不要惊讶。
1JOHN|3|14|我们知道，我们已经出死入生了，因为我们爱弟兄。没有爱心的，仍住在死中。
1JOHN|3|15|凡恨自己弟兄的，就是杀人的；你们知道，凡杀人的，没有永生住在他里面。
1JOHN|3|16|基督为我们舍命，我们从此就知道何为爱；我们也当为弟兄舍命。
1JOHN|3|17|凡有世上财物的，看见弟兄缺乏，却关闭了恻隐的心，上帝的爱怎能住在他里面呢？
1JOHN|3|18|孩子们哪，我们相爱，不要只在言语或舌头上，总要以行为和真诚表现出来。
1JOHN|3|19|从这一点，我们会知道，我们是出于真理的，并且我们在上帝面前可以安心，
1JOHN|3|20|即使我们的心责备自己，上帝比我们的心大，他知道一切。
1JOHN|3|21|亲爱的，我们的心若不责备我们，在上帝面前就可以坦然无惧了。
1JOHN|3|22|我们一切所求的，就从他得着，因为我们遵守他的命令，行他所喜悦的事。
1JOHN|3|23|上帝的命令就是：我们要信他儿子耶稣基督的名，并且照他所赐给我们的命令彼此相爱。
1JOHN|3|24|遵守上帝命令的，住在上帝里面，而上帝也住在他里面。从这一点，我们知道上帝住在我们里面，这是由于他所赐给我们的圣灵。
1JOHN|4|1|亲爱的，一切的灵不可都信，总要察验那些灵是否出于上帝，因为有许多假先知已经来到世上。
1JOHN|4|2|凡宣认耶稣基督是成了肉身而来的灵就是出于上帝的，由此你们可以认出上帝的灵来；
1JOHN|4|3|凡不宣认耶稣的灵，不是出于上帝。这是那敌基督者的灵；你们从前听见他要来，现在他已经在世上了。
1JOHN|4|4|孩子们哪，你们是属上帝的，并且胜过了假先知，因为那在你们里面的比那在世界上的更大。
1JOHN|4|5|他们是属世界的，所以讲论世界的事，而世人也听从他们。
1JOHN|4|6|我们是属上帝的，认识上帝的就听从我们；不属上帝的就不听从我们。从此我们可以认出真理的灵和错谬的灵来。
1JOHN|4|7|亲爱的，我们要彼此相爱，因为爱是从上帝来的。凡有爱的都是由上帝而生，并且认识上帝。
1JOHN|4|8|没有爱的就不认识上帝，因为上帝就是爱。
1JOHN|4|9|上帝差他独一的儿子到世上来，使我们藉着他得生命；由此，上帝对我们的爱就显明了。
1JOHN|4|10|不是我们爱上帝，而是上帝爱我们，差他的儿子为我们的罪作了赎罪祭；这就是爱。
1JOHN|4|11|亲爱的，既然上帝这样爱我们，我们也要彼此相爱。
1JOHN|4|12|从来没有人见过上帝，我们若彼此相爱，上帝就住在我们里面，他的爱在我们里面得以完满了。
1JOHN|4|13|因为上帝将他的灵赐给我们，由此我们知道我们是住在他里面，而他也住在我们里面。
1JOHN|4|14|父差子作世人的救主，这是我们所看见并且作见证的。
1JOHN|4|15|凡宣认耶稣为上帝儿子的，上帝就住在他里面，而他也住在上帝里面。
1JOHN|4|16|我们知道并且深信上帝是爱我们的。 上帝就是爱，住在爱里面的就是住在上帝里面；上帝也住在他里面。
1JOHN|4|17|由此，爱在我们里面得以完满：我们可以在审判的日子坦然无惧，因为基督如何，我们在这世上也如何。
1JOHN|4|18|在爱里没有惧怕；完满的爱把惧怕驱逐出去，因为惧怕里含着惩罚，惧怕的人在爱里尚未得到完满。
1JOHN|4|19|我们爱，因为上帝先爱我们。
1JOHN|4|20|人若说“我爱上帝”，却恨他的弟兄，就是说谎了；不爱他看得见的弟兄，就不能爱看不见的上帝 。
1JOHN|4|21|爱上帝的，也要爱弟兄；这是我们从上帝所受的命令。
1JOHN|5|1|凡信耶稣是基督的，都是从上帝生的；凡爱生他之上帝的，也必爱从上帝生的 。
1JOHN|5|2|我们爱上帝，又实行 他的命令，由此就知道我们爱上帝的儿女了。
1JOHN|5|3|我们遵守上帝的命令，这就是爱他了，而且他的命令并不是难守的。
1JOHN|5|4|因为凡从上帝生的就胜过世界；使我们胜过世界的就是我们的信心。
1JOHN|5|5|胜过世界的是谁呢？不就是那信耶稣是上帝儿子的吗？
1JOHN|5|6|这藉着水和血而来的，就是耶稣基督，不是单用水，而是用水又用血，并且有圣灵作见证，因为圣灵就是真理。
1JOHN|5|7|作见证的有三：
1JOHN|5|8|就是圣灵、水与血，这三样也都是一致的。
1JOHN|5|9|既然我们领受人的见证，上帝的见证更该领受 了，因为上帝的见证是为他儿子作的。
1JOHN|5|10|信上帝儿子的，就有这见证在他心里；不信上帝的，就是把上帝当作说谎的，因为不信上帝为他儿子作的见证。
1JOHN|5|11|这见证就是：上帝赐给我们永生，而这永生是在他儿子里面的。
1JOHN|5|12|那有上帝儿子的，就有生命；没有上帝儿子的，就没有生命。
1JOHN|5|13|我把这些话写给你们信奉上帝儿子之名的人，要让你们知道自己有永生。
1JOHN|5|14|我们若照着上帝的旨意祈求，他就垂听我们；这就是我们对他所存坦然无惧的心。
1JOHN|5|15|既然我们知道他听我们一切所求的，就知道我们所求于他的，无不得着。
1JOHN|5|16|人若看见弟兄犯了不至于死的罪，就要为他祈求，上帝必将生命赐给他—有些人犯的罪是不至于死的；有的是至于死的罪，我不是说要为这罪祈求。
1JOHN|5|17|一切不义的事都是罪，但也有不至于死的罪。
1JOHN|5|18|我们知道，凡从上帝生的，必不犯罪；从上帝生的那一位，必保守他，那邪恶者无法加害于他。
1JOHN|5|19|我们知道，我们是属上帝的，而全世界都伏在那邪恶者的权势之下。
1JOHN|5|20|我们知道，上帝的儿子已经来到，并且将悟性赐给我们，使我们认识那位真实者，我们也在那位真实者里面，就是在他儿子耶稣基督里面。这是真神，也是永生。
1JOHN|5|21|孩子们哪，你们要远避偶像。
