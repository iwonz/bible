MATT|1|1|亞伯拉罕 的後裔、 大衛 的子孫 耶穌基督的家譜：
MATT|1|2|亞伯拉罕 生 以撒 ， 以撒 生 雅各 ， 雅各 生 猶大 和他的兄弟，
MATT|1|3|猶大 從 她瑪 氏生 法勒斯 和 謝拉 ， 法勒斯 生 希斯崙 ， 希斯崙 生 亞蘭 ，
MATT|1|4|亞蘭 生 亞米拿達 ， 亞米拿達 生 拿順 ， 拿順 生 撒門 ，
MATT|1|5|撒門 從 喇合 氏生 波阿斯 ， 波阿斯 從 路得 氏生 俄備得 ， 俄備得 生 耶西 ，
MATT|1|6|耶西 生 大衛 王。 大衛 從 烏利亞 的妻子生 所羅門 ，
MATT|1|7|所羅門 生 羅波安 ， 羅波安 生 亞比雅 ， 亞比雅 生 亞撒 ，
MATT|1|8|亞撒 生 約沙法 ， 約沙法 生 約蘭 ， 約蘭 生 烏西雅 ，
MATT|1|9|烏西雅 生 約坦 ， 約坦 生 亞哈斯 ， 亞哈斯 生 希西家 ，
MATT|1|10|希西家 生 瑪拿西 ， 瑪拿西 生 亞們 ， 亞們 生 約西亞 ，
MATT|1|11|百姓被遷到 巴比倫 的時候， 約西亞 生 耶哥尼雅 和他的兄弟。
MATT|1|12|遷到 巴比倫 之後， 耶哥尼雅 生 撒拉鐵 ， 撒拉鐵 生 所羅巴伯 ，
MATT|1|13|所羅巴伯 生 亞比玉 ， 亞比玉 生 以利亞敬 ， 以利亞敬 生 亞所 ，
MATT|1|14|亞所 生 撒督 ， 撒督 生 亞金 ， 亞金 生 以律 ，
MATT|1|15|以律 生 以利亞撒 ， 以利亞撒 生 馬但 ， 馬但 生 雅各 ，
MATT|1|16|雅各 生 約瑟 ，就是 馬利亞 的丈夫；那稱為基督的耶穌是從 馬利亞 生的。
MATT|1|17|這樣，從 亞伯拉罕 到 大衛 共有十四代，從 大衛 到遷至 巴比倫 的時候也有十四代，從遷至 巴比倫 的時候到基督又有十四代。
MATT|1|18|耶穌基督降生的事記在下面：他母親 馬利亞 已經許配給 約瑟 ，還沒有迎娶， 馬利亞 就從聖靈懷了孕。
MATT|1|19|她丈夫 約瑟 是個義人，不願意當眾羞辱她，想要暗地裏把她休了。
MATT|1|20|正考慮這些事的時候，忽然主的使者在 約瑟 夢中向他顯現，說：「 大衛 的子孫 約瑟 ，不要怕，把你的妻子 馬利亞 娶過來，因她所懷的孕是從聖靈來的。
MATT|1|21|她將要生一個兒子，你要給他起名叫耶穌，因他要將自己的百姓從罪惡裏救出來。」
MATT|1|22|這整件事的發生，是要應驗主藉先知所說的話：
MATT|1|23|「必有童女懷孕生子； 人要稱他的名為 以馬內利 。」 （ 以馬內利 翻出來就是「上帝與我們同在」。）
MATT|1|24|約瑟 醒來，就遵照主的使者的吩咐把妻子娶過來；
MATT|1|25|但是沒有和她同房，直到她生了兒子 ，就給他起名叫耶穌。
MATT|2|1|在 希律 作王的時候，耶穌生在 猶太 的 伯利恆 。有幾個博學之士 從東方來到 耶路撒冷 ，說：
MATT|2|2|「那生下來作 猶太 人之王的在哪裏？我們在東方看見他的星，特來拜他。」
MATT|2|3|希律 王聽見了，就心裏不安； 耶路撒冷 全城的人也都不安。
MATT|2|4|他就召集了祭司長和民間的文士，問他們：「基督該生在哪裏？」
MATT|2|5|他們說：「在 猶太 的 伯利恆 。因為有先知記著：
MATT|2|6|『 猶大 地的 伯利恆 啊， 你在 猶大 諸城中並不是最小的； 因為將來有一位統治者要從你那裏出來， 牧養我 以色列 民。』」
MATT|2|7|於是， 希律 暗地裏召了博學之士來，查問那星是甚麼時候出現的，
MATT|2|8|就派他們往 伯利恆 去，說：「你們去仔細尋訪那小孩子，找到了就來報信，我也好去拜他。」
MATT|2|9|他們聽了王的話就去了。忽然，在東方所看到的那顆星在前面引領他們，一直行到小孩子所在地方的上方就停住了。
MATT|2|10|他們看見那星，就非常歡喜；
MATT|2|11|進了房子，看見小孩子和他母親 馬利亞 ，就俯伏拜那小孩子，揭開寶盒，拿出黃金、乳香、沒藥，作為禮物獻給他。
MATT|2|12|因為在夢中得到主的指示，不要回去見 希律 ，他們就從別的路回自己的家鄉去了。
MATT|2|13|他們走後，忽然主的使者在 約瑟 夢中向他顯現，說：「起來！帶著小孩子和他母親逃往 埃及 ，住在那裏，等我的指示；因為 希律 要搜尋那小孩子來殺害他。」
MATT|2|14|約瑟 就起來，連夜帶著小孩子和他母親往 埃及 去，
MATT|2|15|住在那裏，直到 希律 死了。這是要應驗主藉先知所說的話：「我從 埃及 召我的兒子出來。」
MATT|2|16|希律 見自己被博學之士愚弄，極其憤怒，差人將 伯利恆 城裏和四境所有的男孩，根據他向博學之士仔細查問到的時間，凡兩歲以內的，都殺盡了。
MATT|2|17|這就應驗了 耶利米 先知所說的話：
MATT|2|18|「在 拉瑪 聽見號咷大哭的聲音， 是 拉結 哭她兒女； 她不肯受安慰， 因為他們都不在了。」
MATT|2|19|希律 死了以後，在 埃及 ，忽然主的使者在 約瑟 夢中向他顯現，
MATT|2|20|說：「起來，帶著小孩子和他母親回 以色列 地去！因為要殺害這小孩子的人已經死了。」
MATT|2|21|約瑟 就起來，帶著小孩子和他母親進入 以色列 地去。
MATT|2|22|但是他因聽見 亞基老 繼承他父親 希律 作了 猶太 王，怕到那裏去；又在夢中得到主的指示，就往 加利利 境內去了。
MATT|2|23|他們到了一座城，名叫 拿撒勒 ，就住在那裏。這是要應驗先知所說的話：「他將稱為 拿撒勒 人。」
MATT|3|1|在那些日子，施洗的 約翰 出來，在 猶太 的曠野宣講：
MATT|3|2|「你們要悔改！因為天國近了。」
MATT|3|3|這人就是 以賽亞 先知所說的： 「在曠野有聲音呼喊著： 預備主的道， 修直他的路。」
MATT|3|4|這 約翰 身穿駱駝毛的衣服，腰束皮帶，吃的是蝗蟲和野蜜。
MATT|3|5|那時， 耶路撒冷 、全 猶太 和全 約旦河 地區的人，都到 約翰 那裏去，
MATT|3|6|承認他們的罪，在 約旦河 裏受他的洗。
MATT|3|7|約翰 看見許多法利賽人和撒都該人也來受洗，就對他們說：「毒蛇的孽種啊，誰指示你們逃避那將要來的憤怒呢？
MATT|3|8|你們要結出果子來，和悔改的心相稱。
MATT|3|9|不要自己心裏說：『我們有 亞伯拉罕 為祖宗。』我告訴你們，上帝能從這些石頭中給 亞伯拉罕 興起子孫來。
MATT|3|10|現在斧子已經放在樹根上，凡不結好果子的樹就砍下來，丟在火裏。
MATT|3|11|我是用水給你們施洗，叫你們悔改；但那在我以後來的，能力比我更大，我就是給他提鞋子也不配，他要用聖靈與火給你們施洗。
MATT|3|12|他手裏拿著簸箕，要揚淨他的穀物，把麥子收在倉裏，把糠用不滅的火燒盡。」
MATT|3|13|當時，耶穌從 加利利 來到 約旦河 ，到了 約翰 那裏，請 約翰 為他施洗。
MATT|3|14|約翰 想要阻止他，說：「我應該受你的洗，你怎麼到我這裏來呢？」
MATT|3|15|耶穌回答他：「暫且這樣做吧，因為我們理當這樣履行全部的義 。」於是 約翰 就依了他。
MATT|3|16|耶穌受了洗，隨即從水裏上來。天忽然為他 開了，他看見上帝的靈降下，彷彿鴿子落在他身上。
MATT|3|17|這時，天上有聲音說：「這是我的愛子，我所喜愛的。」
MATT|4|1|當時，耶穌被聖靈引到曠野，受魔鬼的試探。
MATT|4|2|他禁食四十晝夜，後來就餓了。
MATT|4|3|那試探者進前來對他說：「你若是上帝的兒子，叫這些石頭變成食物吧。」
MATT|4|4|耶穌卻回答說：「經上記著： 『人活著，不是單靠食物， 乃是靠上帝口裏所出的一切話。』」
MATT|4|5|魔鬼就帶他進了聖城，叫他站在聖殿頂上，
MATT|4|6|對他說：「你若是上帝的兒子，就跳下去！因為經上記著： 『主要為你命令他的使者， 用手托住你， 免得你的腳碰在石頭上。』」
MATT|4|7|耶穌對他說：「經上又記著：『不可試探主—你的上帝。』」
MATT|4|8|魔鬼又帶他上了一座很高的山，將世上的萬國和萬國的榮華都指給他看，
MATT|4|9|對他說：「你若俯伏拜我，我就把這一切賜給你。」
MATT|4|10|耶穌說：「撒但 ，退去！因為經上記著： 『要拜主—你的上帝， 惟獨事奉他。』」
MATT|4|11|於是，魔鬼離開了耶穌，立刻有天使來伺候他。
MATT|4|12|耶穌聽見 約翰 下了監，就退到 加利利 去；
MATT|4|13|後來離開 拿撒勒 ，往 迦百農 去，住在那裏。那地方靠海，在 西布倫 和 拿弗他利 地區。
MATT|4|14|這是要應驗 以賽亞 先知所說的話：
MATT|4|15|「 西布倫 ， 拿弗他利 ， 沿海的路， 約旦河 的東邊， 外邦人的 加利利 —
MATT|4|16|那坐在黑暗裏的百姓 看見了大光； 坐在死蔭之地的人 有光照耀他們。」
MATT|4|17|從那時候，耶穌開始宣講，說：「你們要悔改！因為天國近了。」
MATT|4|18|耶穌沿著 加利利 海邊行走，看見兩兄弟，就是那叫 彼得 的 西門 和他弟弟 安得烈 ，正往海裏撒網；他們本是打魚的。
MATT|4|19|耶穌對他們說：「來跟從我，我要叫你們得人如得魚一樣。」
MATT|4|20|他們立刻捨了網，跟從他。
MATT|4|21|耶穌從那裏往前走，看見另外兩兄弟，就是 西庇太 的兒子 雅各 和他弟弟 約翰 ，同他們的父親 西庇太 在船上補網，耶穌就呼召他們。
MATT|4|22|他們立刻捨了船，辭別父親，跟從了耶穌。
MATT|4|23|耶穌走遍 加利利 ，在各會堂裏教導人，宣講天國的福音，醫治百姓各樣的疾病。
MATT|4|24|他的名聲傳遍了 敘利亞 。那裏的人把一切病人，就是有各樣疾病和疼痛的、被鬼附的、癲癇的、癱瘓的，都帶了來，耶穌就治好了他們。
MATT|4|25|當時，有一大群人從 加利利 、 低加坡里 、 耶路撒冷 、 猶太 、 約旦河 的東邊，來跟從他。
MATT|5|1|耶穌看見這一群人，就上了山，坐下後，門徒到他跟前來，
MATT|5|2|他開口教導他們說：
MATT|5|3|「心靈貧窮的人有福了！ 因為天國是他們的。
MATT|5|4|哀慟的人有福了！ 因為他們必得安慰。
MATT|5|5|謙和的人有福了！ 因為他們必承受土地。
MATT|5|6|飢渴慕義的人有福了！ 因為他們必得飽足。
MATT|5|7|憐憫人的人有福了！ 因為他們必蒙憐憫。
MATT|5|8|清心的人有福了！ 因為他們必得見上帝。
MATT|5|9|締造和平的人有福了！ 因為他們必稱為上帝的兒子。
MATT|5|10|為義受迫害的人有福了！ 因為天國是他們的。
MATT|5|11|「人若因我辱罵你們，迫害你們，捏造各樣壞話毀謗你們 ，你們就有福了！
MATT|5|12|要歡喜快樂，因為你們在天上的賞賜是很多的。在你們以前的先知，人也是這樣迫害他們。」
MATT|5|13|「你們是地上的鹽。鹽若失了味，怎能叫它再鹹呢？它不再有用，只好被丟在外面，任人踐踏。
MATT|5|14|你們是世上的光。城造在山上是不能隱藏的。
MATT|5|15|人點燈，不放在斗底下，而是放在燈臺上，就照亮一家的人。
MATT|5|16|你們的光也要這樣照在人前，叫他們看見你們的好行為，把榮耀歸給你們在天上的父。」
MATT|5|17|「不要以為我來是要廢掉律法和先知。我來不是要廢掉，而是要成全。
MATT|5|18|我實在告訴你們，就是到天地都廢去，律法的一點一畫也不能廢去，直到一切都實現。
MATT|5|19|所以，無論誰廢掉這誡命中最小的一條，又教導人也這樣做，他在天國裏要稱為最小的。但無論誰遵行並如此教導人的，他在天國裏要稱為大。
MATT|5|20|我告訴你們，你們的義若不勝過文士和法利賽人的義，絕不能進天國。」
MATT|5|21|「你們聽過有對古人說：『不可殺人』；『凡殺人的，必須受審判。』
MATT|5|22|但是我告訴你們：凡向弟兄動怒的，必須受審判；凡罵弟兄是廢物的，必須受議會的審判；凡罵弟兄是白痴的，必須遭受地獄的火。
MATT|5|23|所以，你在祭壇上獻祭物的時候，若想起有弟兄對你懷恨，
MATT|5|24|就要把祭物留在壇前，先去跟弟兄和好，然後來獻祭物。
MATT|5|25|你同告你的冤家還在路上，就要趕快與他講和，免得他把你送交給法官，法官交給警衛，你就下在監裏了。
MATT|5|26|我實在告訴你，就是有一個大文錢 還沒有還清，你也絕不能從那裏出來。」
MATT|5|27|「你們聽過有話說：『不可姦淫。』
MATT|5|28|但是我告訴你們：凡看見婦女就動淫念的，這人心裏已經與她犯姦淫了。
MATT|5|29|若是你的右眼使你跌倒，就把它挖出來，丟掉。寧可失去身體中的一部分，也不讓整個身體被扔進地獄。
MATT|5|30|若是你的右手使你跌倒，就把它砍下來，丟掉。寧可失去身體中的一部分，也不讓整個身體下地獄。」
MATT|5|31|「又有話說：『無論誰休妻，都要給她休書。』
MATT|5|32|但是我告訴你們：凡休妻的，除非是因不貞的緣故，否則就是使她犯姦淫了；人若娶被休的婦人，也是犯姦淫了。」
MATT|5|33|「你們又聽過有對古人說：『不可背誓，所起的誓總要向主謹守。』
MATT|5|34|但是我告訴你們：甚麼誓都不可起。不可指著天起誓，因為天是上帝的寶座。
MATT|5|35|不可指著地起誓，因為地是他的腳凳；也不可指著 耶路撒冷 起誓，因為 耶路撒冷 是大君王的京城。
MATT|5|36|又不可指著你的頭起誓，因為你不能使一根頭髮變黑變白。
MATT|5|37|你們的話，是，就說是；不是，就說不是。若再多說，就是出於那惡者。」
MATT|5|38|「你們聽過有話說：『以眼還眼，以牙還牙。』
MATT|5|39|但是我告訴你們：不要與惡人作對。有人打你的右臉，連另一邊也轉過去由他打。
MATT|5|40|有人想要告你，要拿你的裏衣，連外衣也由他拿去。
MATT|5|41|有人強迫你走一里 路，你就跟他走二里。
MATT|5|42|有求你的，就給他；有向你借貸的，不可推辭。」
MATT|5|43|「你們聽過有話說：『要愛你的鄰舍，恨你的仇敵。』
MATT|5|44|但是我告訴你們：要愛你們的仇敵，為那迫害你們的禱告。
MATT|5|45|這樣，你們就可以作天父的兒女了。因為他叫太陽照好人，也照壞人；降雨給義人，也給不義的人。
MATT|5|46|你們若只愛那愛你們的人，有甚麼賞賜呢？就是稅吏不也是這樣做嗎？
MATT|5|47|你們若只請你弟兄的安，有甚麼比別人強呢？就是外邦人不也是這樣做嗎？
MATT|5|48|所以，你們要完全，如同你們的天父是完全的。」
MATT|6|1|「你們要謹慎，不可故意在人面前表現虔誠，叫他們看見，若是這樣，就不能得你們天父的賞賜了。
MATT|6|2|「所以，你施捨的時候，不可叫人在你前面吹號，像那假冒為善的人在會堂裏和街道上所做的，故意要得人的稱讚。我實在告訴你們，他們已經得了他們的賞賜。
MATT|6|3|你施捨的時候，不要讓左手知道右手所做的，
MATT|6|4|好使你隱祕地施捨；你父在隱祕中察看，必然賞賜你。」
MATT|6|5|「你們禱告的時候，不可像那假冒為善的人，愛站在會堂裏和十字路口禱告，故意讓人看見。我實在告訴你們，他們已經得了他們的賞賜。
MATT|6|6|你禱告的時候，要進入內室，關上門，向那在隱祕中的父禱告；你父在隱祕中察看，必將賞賜你。
MATT|6|7|你們禱告，不可像外邦人那樣重複一些空話，他們以為話多了必蒙垂聽。
MATT|6|8|你們不可效法他們。因為在你們祈求以前，你們所需要的，你們的父早已知道了。」
MATT|6|9|「所以，你們要這樣禱告： 『我們在天上的父： 願人都尊你的名為聖。
MATT|6|10|願你的國降臨； 願你的旨意行在地上， 如同行在天上。
MATT|6|11|我們日用的飲食，今日賜給我們。
MATT|6|12|免我們的債， 如同我們免了人的債。
MATT|6|13|不叫我們陷入試探； 救我們脫離那惡者。 因為國度、權柄、榮耀，全是你的， 直到永遠。阿們！ 』
MATT|6|14|「你們若饒恕人的過犯，你們的天父也必饒恕你們；
MATT|6|15|你們若不饒恕人 ，你們的天父也必不饒恕你們的過犯。」
MATT|6|16|「你們禁食的時候，不可像那假冒為善的人，臉上帶著愁容；因為他們蓬頭垢面，故意讓人看出他們在禁食。我實在告訴你們，他們已經得了他們的賞賜。
MATT|6|17|你禁食的時候，要梳頭洗臉，
MATT|6|18|不要讓人看出你在禁食，只讓你隱祕中的父看見；你父在隱祕中察看，必然賞賜你。」
MATT|6|19|「不要為自己在地上積蓄財寶；地上有蟲子咬，能銹壞，也有賊挖洞來偷。
MATT|6|20|要在天上積蓄財寶；天上沒有蟲子咬，不會銹壞，也沒有賊挖洞來偷。
MATT|6|21|因為你的財寶在哪裏，你的心也在哪裏。」
MATT|6|22|「眼睛是身體的燈。你的眼睛若明亮，全身就光明；
MATT|6|23|你的眼睛若昏花，全身就黑暗。你裏面的光若黑暗了，那黑暗是何等大呢！」
MATT|6|24|「一個人不能服侍兩個主；他不是恨這個愛那個，就是重這個輕那個。你們不能又服侍上帝，又服侍 瑪門 。」
MATT|6|25|「所以，我告訴你們，不要為你們的生命憂慮吃甚麼喝甚麼 ，或為你們的身體憂慮穿甚麼。生命不勝於飲食嗎？身體不勝於衣裳嗎？
MATT|6|26|你們看一看那天上的飛鳥，也不種也不收，也不在倉裏存糧，你們的天父尚且養活牠們。你們不比飛鳥貴重得多嗎？
MATT|6|27|你們哪一個能藉著憂慮使壽數多加一刻呢 ？
MATT|6|28|何必為衣裳憂慮呢？你們想一想野地裏的百合花是怎麼長起來的：它也不勞動也不紡線。
MATT|6|29|然而我告訴你們，就是 所羅門 極榮華的時候，他所穿戴的還不如這些花的一朵呢！
MATT|6|30|你們這小信的人哪！野地裏的草今天還在，明天就丟在爐裏，上帝還給它這樣的妝飾，何況你們呢？
MATT|6|31|所以，不要憂慮，說：『我們吃甚麼？喝甚麼？穿甚麼？』
MATT|6|32|這都是外邦人所求的。你們需要這一切東西，你們的天父都知道。
MATT|6|33|你們要先求上帝的國和他的義，這些東西都要加給你們了。
MATT|6|34|所以，不要為明天憂慮，因為明天自有明天的憂慮；一天的難處一天當就夠了。」
MATT|7|1|「你們不要評斷別人，免得你們被審判。
MATT|7|2|因為你們怎樣評斷別人，也必怎樣被審判；你們用甚麼量器量給人，也必用甚麼量器量給你們。
MATT|7|3|為甚麼看見你弟兄眼中有刺，卻不想自己眼中有梁木呢？
MATT|7|4|你自己眼中有梁木，怎能對你弟兄說『讓我去掉你眼中的刺』呢？
MATT|7|5|你這假冒為善的人！先去掉自己眼中的梁木，然後才能看得清楚，好去掉你弟兄眼中的刺。
MATT|7|6|不要把聖物給狗，也不要把你們的珍珠丟在豬面前，恐怕牠們踐踏了珍珠，轉過來咬你們。」
MATT|7|7|「你們祈求，就給你們；尋找，就找到；叩門，就給你們開門。
MATT|7|8|因為凡祈求的，就得著；尋找的，就找到；叩門的，就給他開門。
MATT|7|9|你們中間誰有兒子求餅，反給他石頭呢？
MATT|7|10|求魚，反給他蛇呢？
MATT|7|11|你們雖然不好，尚且知道拿好東西給兒女，何況你們在天上的父，他豈不更要把好東西賜給求他的人嗎？
MATT|7|12|所以，無論何事，你們想要人怎樣待你們，你們也要怎樣待人，因為這就是律法和先知的道理。」
MATT|7|13|「你們要進窄門。因為通往滅亡的門是寬的，路是大的，進去的人也多；
MATT|7|14|通往生命的門是窄的，路是小的，找到的人也少。」
MATT|7|15|「你們要防備假先知。他們到你們這裏來，外面披著羊皮，裏面卻是殘暴的狼。
MATT|7|16|豈能在荊棘上摘葡萄呢？豈能在蒺藜裏摘無花果呢？憑著他們的果子，就可以認出他們來。
MATT|7|17|這樣，凡好樹都結好果子，而壞樹結壞果子。
MATT|7|18|好樹不能結壞果子，壞樹也不能結好果子。
MATT|7|19|凡不結好果子的樹就砍下來，丟在火裏。
MATT|7|20|所以，憑著他們的果子就可以認出他們來。」
MATT|7|21|「不是每一個稱呼我『主啊，主啊』的人都能進天國；惟有遵行我天父旨意的人才能進去。
MATT|7|22|在那日必有許多人對我說：『主啊，主啊，我們不是奉你的名傳道，奉你的名趕鬼，奉你的名行許多異能嗎？』
MATT|7|23|我要向他們宣告：『我從來不認識你們，你們這些作惡的人，給我走開！』」
MATT|7|24|「所以，凡聽了我這些話又去做的，好比一個聰明人把房子蓋在磐石上。
MATT|7|25|風吹，雨打，水沖，撞擊那房子，房子總不倒塌，因為根基立在磐石上。
MATT|7|26|凡聽了我這些話而不去做的，好比一個無知的人把房子蓋在沙土上。
MATT|7|27|風吹，雨打，水沖，撞擊那房子，房子就倒塌了，並且倒塌得很厲害。」
MATT|7|28|耶穌講完了這些話，眾人對他的教導都感到驚奇，
MATT|7|29|因為他教導他們正像有權柄的人，不像他們的文士。
MATT|8|1|耶穌下了山，有一大群人跟著他。
MATT|8|2|這時，一個痲瘋病人前來拜他，說：「主啊，你若肯，你能使我潔淨。」
MATT|8|3|耶穌伸手摸他，說：「我肯，你潔淨了吧！」他的痲瘋病立刻就潔淨了。
MATT|8|4|耶穌對他說：「你要注意，不可告訴任何人，只要去，讓祭司為你檢查，並獻上 摩西 所吩咐的祭物，作為證據給眾人看。」
MATT|8|5|耶穌進了 迦百農 ，有一個百夫長進前來，求他，
MATT|8|6|說：「主啊，我的僮僕癱瘓了，躺在家裏，非常痛苦。」
MATT|8|7|耶穌說：「我去醫治他。」
MATT|8|8|百夫長回答：「主啊，你到舍下來，我不敢當；只要你說一句話，我的僮僕就會痊癒。
MATT|8|9|因為我在人的權下，也有兵在我以下。我對這個說：『去！』他就去；對那個說：『來！』他就來；對我的僕人說：『做這事！』他就去做。」
MATT|8|10|耶穌聽了就很驚訝，對跟從的人說：「我實在告訴你們，這麼大的信心，就是在 以色列 ，我也沒有見過。
MATT|8|11|我又告訴你們，從東從西，將有許多人來，在天國裏與 亞伯拉罕 、 以撒 、 雅各 一同坐席；
MATT|8|12|本國的子民反而被趕到外邊黑暗裏去，在那裏要哀哭切齒了。」
MATT|8|13|耶穌對百夫長說：「你回去吧！照你的信心成全你了。」就在那時，他的僮僕好了。
MATT|8|14|耶穌到了 彼得 家裏，見 彼得 的岳母正發燒躺著。
MATT|8|15|耶穌一摸她的手，燒就退了，於是她起來服事耶穌。
MATT|8|16|傍晚的時候，有人帶著許多被鬼附的來到耶穌跟前，他只用一句話就把邪靈都趕出去，並且治好了一切有病的人。
MATT|8|17|這是要應驗 以賽亞 先知所說的話： 「他代替了我們的軟弱， 擔當了我們的疾病。」
MATT|8|18|耶穌見許多人圍著他，就吩咐渡到對岸去。
MATT|8|19|有一個文士進前來對他說：「老師，你無論往哪裏去，我都要跟從你。」
MATT|8|20|耶穌說：「狐狸有洞，天空的飛鳥有窩，人子卻沒有枕頭的地方。」
MATT|8|21|又有一個門徒對耶穌說：「主啊，容許我先回去埋葬我的父親。」
MATT|8|22|耶穌說：「讓死人埋葬他們的死人。你跟從我吧！」
MATT|8|23|耶穌上了船，門徒跟著他。
MATT|8|24|海裏忽然起了猛烈的風暴，以致船幾乎被波浪淹沒，耶穌卻睡著了。
MATT|8|25|門徒去叫醒他，說：「主啊，救命啊，我們快沒命啦！」
MATT|8|26|耶穌說：「你們這些小信的人哪，為甚麼膽怯呢？」於是他起來，斥責風和海，風和海就大大平靜了。
MATT|8|27|眾人驚訝地說：「這是怎樣的一個人？連風和海都聽從他。」
MATT|8|28|耶穌渡到對岸去，到 加大拉 人 的地區，有兩個被鬼附的人從墳墓迎著他走來。他們極其兇猛，甚至沒有人敢從那條路經過。
MATT|8|29|他們喊著說：「上帝的兒子，你為甚麼干擾我們？時候還沒有到，你就上這裏來叫我們受苦嗎？」
MATT|8|30|離他們很遠，有一大群豬正在吃食。
MATT|8|31|鬼就央求耶穌，說：「若要把我們趕出去，就打發我們進入豬群吧！」
MATT|8|32|耶穌對他們說：「去吧！」鬼就出來，進入豬群。一轉眼，整群豬都闖下山崖，投進海裏，淹死了。
MATT|8|33|放豬的就逃進城去，把這一切事和被鬼附的人所遭遇的都告訴眾人。
MATT|8|34|全城的人都出來迎見耶穌，見了他以後，就央求他離開他們的地區。
MATT|9|1|耶穌上了船，渡過海，來到自己的城裏。
MATT|9|2|有人用褥子抬著一個癱子到耶穌跟前來。耶穌見他們的信心，就對癱子說：「孩子，放心吧，你的罪赦了。」
MATT|9|3|這時，有幾個文士心裏說：「這個人說褻瀆的話了。」
MATT|9|4|耶穌知道他們的心思，就說：「你們心裏為甚麼懷著惡念呢？
MATT|9|5|說『你的罪赦了』，或說『你起來行走』，哪一樣容易呢？
MATT|9|6|但要讓你們知道，人子在地上有赦罪的權柄」，於是對癱子說：「起來！拿你的褥子回家去吧。」
MATT|9|7|那人就起來，回家去了。
MATT|9|8|眾人看見都畏懼，歸榮耀給上帝，因為他把這樣的權柄賜給人。
MATT|9|9|耶穌從那裏往前走，看見一個人名叫 馬太 ，在稅關坐著，就對他說：「來跟從我！」他就起來跟從耶穌。
MATT|9|10|耶穌在屋裏坐席的時候，有好些稅吏和罪人來，與耶穌和他的門徒一同坐席。
MATT|9|11|法利賽人看見，就對耶穌的門徒說：「你們的老師為甚麼與稅吏和罪人一同吃飯呢？」
MATT|9|12|耶穌聽見，就說：「健康的人用不著醫生；有病的人才用得著。
MATT|9|13|經上說：『我喜愛憐憫，不喜愛祭祀。』這句話的意思，你們去揣摩。我不是來召義人，而是召罪人。」
MATT|9|14|那時， 約翰 的門徒來見耶穌，說：「我們和法利賽人常常 禁食，你的門徒卻不禁食，這是為甚麼呢？」
MATT|9|15|耶穌對他們說：「新郎和賓客在一起的時候，賓客怎麼能哀慟呢？但日子將到，新郎要被帶走，那時候他們就要禁食了。
MATT|9|16|沒有人把新布補在舊衣服上；因為所補上的會撕破那衣服，裂口就更大了。
MATT|9|17|也沒有人把新酒裝在舊皮袋裏，若是這樣，皮袋會脹破，酒就漏出來，皮袋也糟蹋了。相反地，把新酒裝在新皮袋裏，兩樣就都保全了。」
MATT|9|18|耶穌說這些話的時候，有一個會堂主管來，向他下跪，說：「我女兒剛死了，求你去按手在她身上，她就會活過來。」
MATT|9|19|耶穌就起來跟他去；門徒也跟了去。
MATT|9|20|這時，有一個女人，患了經血不止的病有十二年，來到耶穌背後，摸他的衣裳繸子；
MATT|9|21|因為她心裏說：「我只要摸他的衣裳，就會痊癒。」
MATT|9|22|耶穌轉過來，看見她，就說：「女兒，放心！你的信救了你。」從那時起，這女人就痊癒了。
MATT|9|23|耶穌到了會堂主管的家裏，看見吹鼓手和亂哄哄的一群人，
MATT|9|24|就說：「退去吧！這女孩不是死了，而是睡著了。」他們就嘲笑他。
MATT|9|25|眾人被趕出後，耶穌就進去，拉著女孩的手，女孩就起來了。
MATT|9|26|於是這消息傳遍了那地方。
MATT|9|27|耶穌從那裏往前走，有兩個盲人跟著他，喊叫說：「 大衛 之子，可憐我們吧！」
MATT|9|28|耶穌進了屋子，盲人就來到他跟前。耶穌說：「你們信我能做這事嗎？」他們說：「主啊，我們信。」
MATT|9|29|耶穌就摸他們的眼睛，說：「照著你們的信心成全你們吧。」
MATT|9|30|他們的眼睛就開了。耶穌嚴嚴地叮囑他們說：「要小心，不可讓人知道。」
MATT|9|31|他們出去，竟把他的名聲傳遍了那地方。
MATT|9|32|他們出去的時候，有人把一個被鬼附的啞巴帶到耶穌跟前來。
MATT|9|33|鬼被趕出去，啞巴就說出話來。眾人都很驚訝，說：「在 以色列 ，從來沒有見過這樣的事。」
MATT|9|34|法利賽人卻說：「他是靠著鬼王趕鬼的。」
MATT|9|35|耶穌走遍各城各鄉，在他們的會堂裏教導人，宣講天國的福音，又醫治各樣的病症。
MATT|9|36|他看見一大群人，就憐憫他們；因為他們困苦無助，如同羊沒有牧人一樣。
MATT|9|37|於是他對門徒說：「要收的莊稼多，做工的人少。
MATT|9|38|所以，你們要求莊稼的主差遣做工的人出去收他的莊稼。」
MATT|10|1|耶穌叫了十二個門徒來，給他們權柄，能驅趕污靈和醫治各樣的疾病。
MATT|10|2|這十二使徒的名字如下：頭一個叫 西門 （又稱 彼得 ），還有他弟弟 安得烈 ， 西庇太 的兒子 雅各 和 雅各 的弟弟 約翰 ，
MATT|10|3|腓力 和 巴多羅買 ， 多馬 和稅吏 馬太 ， 亞勒腓 的兒子 雅各 ，和 達太 ，
MATT|10|4|激進黨的 西門 ，還有出賣耶穌的 加略 人 猶大 。
MATT|10|5|耶穌差遣這十二個人出去，吩咐他們說：「外邦人的路，你們不要走； 撒瑪利亞 人的城，你們不要進；
MATT|10|6|寧可往 以色列 家迷失的羊那裏去。
MATT|10|7|要邊走邊傳，說『天國近了』。
MATT|10|8|要醫治病人，使死人復活，使痲瘋病人潔淨，把鬼趕出去。你們白白地得來，也要白白地給人。
MATT|10|9|腰袋裏不要帶金銀銅錢；
MATT|10|10|途中不要帶行囊，不要帶兩件內衣，也不要帶鞋子和手杖，因為工人得飲食是應當的。
MATT|10|11|你們無論進哪一城、哪一村，要打聽那裏誰是合適的人，就住在他家，直住到離開的時候。
MATT|10|12|進他家時，要向那家請安。
MATT|10|13|那家若配得平安，你們所求的平安就臨到那家；若不配得，你們所求的平安仍歸你們。
MATT|10|14|凡不接待你們，不聽你們話的人，你們離開那家，或是那城的時候，要跺掉你們腳上的塵土。
MATT|10|15|我實在告訴你們，在審判的日子， 所多瑪 和 蛾摩拉 地方所受的，比那城還容易受呢！」
MATT|10|16|「看哪！我差你們出去，如同羊進入狼群，所以你們要機警如蛇，純真如鴿。
MATT|10|17|你們要防備那些人，因為他們要把你們交給議會，也要在會堂裏鞭打你們。
MATT|10|18|你們要為我的緣故被送到統治者和君王面前，對他們和外邦人作見證。
MATT|10|19|當人把你們交出時，不要擔心怎樣說話，或說甚麼話。到那時候，必賜給你們該說的話，
MATT|10|20|因為不是你們自己說的，而是你們父的靈在你們裏面說的。
MATT|10|21|兄弟要把兄弟、父親要把兒女置於死地；兒女要起來與父母為敵，害死他們。
MATT|10|22|而且你們要為我的名被眾人憎恨。但堅忍到底的終必得救。
MATT|10|23|有人在這城迫害你們，就逃到另一城去。 我實在告訴你們， 以色列 的城鎮，你們還沒有走遍，人子就要來臨。
MATT|10|24|「學生不高過老師，僕人不高過主人。
MATT|10|25|學生所遭遇的與老師一樣，僕人所遭遇的與主人一樣，也就夠了。既然有人罵一家的主人是『 別西卜 』 ，更何況他的家人呢？」
MATT|10|26|「所以，不要怕他們，因為掩蓋的事沒有不顯露出來的，隱藏的事也沒有不被知道的。
MATT|10|27|我在暗中告訴你們的，你們要在明處說出來；你們耳中所聽的，要在屋頂上宣揚出來。
MATT|10|28|那殺人身體但不能滅人靈魂的，不要怕他們；惟有那能在地獄裏毀滅身體和靈魂的，才要怕他。
MATT|10|29|兩隻麻雀不是賣一銅錢 嗎？你們的父若不許，一隻也不會掉在地上。
MATT|10|30|就是你們的頭髮也都數過了。
MATT|10|31|所以，不要懼怕，你們比許多的麻雀還貴重！」
MATT|10|32|「所以，凡在人面前認我的，我在我天上的父面前也必認他；
MATT|10|33|凡在人面前不認我的，我在我天上的父面前也必不認他。」
MATT|10|34|「你們不要以為我來是帶給地上和平，我來並不是帶來和平，而是刀劍。
MATT|10|35|因為我來是要叫 『人與父親對立， 女兒與母親對立， 媳婦與婆婆對立。
MATT|10|36|人的仇敵就是自己家裏的人。』
MATT|10|37|愛父母勝過愛我的，不配作我的門徒；愛兒女勝過愛我的，不配作我的門徒。
MATT|10|38|不背自己的十字架跟從我的，不配作我的門徒。
MATT|10|39|得著性命的，要喪失性命；為我喪失性命的，要得著性命。」
MATT|10|40|「接納你們的就是接納我；接納我的就是接納差遣我來的那位。
MATT|10|41|把先知當作先知接納的，必得先知的賞賜；把義人當作義人接納的，必得義人的賞賜。
MATT|10|42|無論誰，只因門徒的名，就算把一杯涼水給這些小子中的一個喝，我實在告訴你們，他一定會得到賞賜。」
MATT|11|1|耶穌吩咐完了十二個門徒，就離開那裏，往各城去傳道，教導人。
MATT|11|2|約翰 在監獄裏聽見基督所做的事，就派他的門徒去，
MATT|11|3|問耶穌：「將要來的那位就是你嗎？還是我們要等候另一位呢？」
MATT|11|4|耶穌回答他們：「你們去，把所聽見、所看見的告訴 約翰 ：
MATT|11|5|就是盲人看見，瘸子行走，痲瘋病人得潔淨，聾子聽見，死人復活，窮人聽到福音。
MATT|11|6|凡不因我跌倒的有福了！」
MATT|11|7|他們一走，耶穌就對眾人談到 約翰 ，說：「你們從前到曠野去，是要看甚麼呢？看風吹動的蘆葦嗎？
MATT|11|8|你們出去到底是要看甚麼？看穿細軟衣服的人嗎？那穿細軟衣服的人是在王宮裏。
MATT|11|9|你們出去究竟是要看甚麼？是先知嗎？是的，我告訴你們，他比先知大多了。
MATT|11|10|這個人就是經上所說的： 『看哪，我要差遣我的使者在你面前， 他要在你前面為你預備道路。』
MATT|11|11|我實在告訴你們，凡女子所生的，沒有一個比施洗 約翰 大；但在天國裏，最小的比他還大。
MATT|11|12|從施洗 約翰 的日子到今天，天國受到強烈的攻擊，強者奪取它 。
MATT|11|13|眾先知和律法，直到 約翰 為止，都說了預言。
MATT|11|14|如果你們願意接受，這人就是那要來的 以利亞 。
MATT|11|15|有耳的，就應當聽！
MATT|11|16|「我該用甚麼來比這世代呢？這正像孩童坐在街市上向同伴呼喊：
MATT|11|17|『我們為你們吹笛，你們不跳舞； 我們唱哀歌，你們不捶胸。』
MATT|11|18|約翰 來了，既不吃也不喝，人們就說他是被鬼附的；
MATT|11|19|人子來了，也吃也喝，他們又說這人貪食好酒，是稅吏和罪人的朋友。而智慧是由它的果子來證實的 。」
MATT|11|20|那時，耶穌在一些城行了許多異能。因為城裏的人不肯悔改，他就責備那些城說：
MATT|11|21|「 哥拉汛 哪，你有禍了！ 伯賽大 啊，你有禍了！因為在你們中間所行的異能若行在 推羅 、 西頓 ，他們早已披麻蒙灰悔改了。
MATT|11|22|但我告訴你們，在審判的日子， 推羅 和 西頓 所受的，比你們還容易受呢！
MATT|11|23|迦百農 啊， 你以為要被舉到天上嗎？ 你要被推下陰間！ 因為在你那裏所行的異能，若行在 所多瑪 ，它還可以存留到今日。
MATT|11|24|但我告訴你們，在審判的日子， 所多瑪 地方所受的，比你們還容易受呢！」
MATT|11|25|那時，耶穌說：「父啊，天地的主，我感謝你！因為你把這些事向聰明智慧的人隱藏起來，而向嬰孩啟示出來。
MATT|11|26|父啊，是的，因為你的美意本是如此。
MATT|11|27|一切都是我父交給我的；除了父，沒有人知道子；除了子和子所願意啟示的人，沒有人知道父。
MATT|11|28|凡勞苦擔重擔的人都到我這裏來，我要使你們得安息。
MATT|11|29|我心裏柔和謙卑，你們當負我的軛，向我學習；這樣，你們的心靈就必得安息。
MATT|11|30|因為我的軛是容易的，我的擔子是輕省的。」
MATT|12|1|那時，耶穌在安息日從麥田經過。他的門徒餓了，就摘麥穗來吃。
MATT|12|2|法利賽人看見，對耶穌說：「看哪，你的門徒在安息日做不合法的事了。」
MATT|12|3|耶穌對他們說：「 大衛 和跟從他的人飢餓時所做的事，你們沒有念過嗎？
MATT|12|4|他怎麼進了上帝的居所，吃了供餅呢？這餅是他和跟從他的人不可以吃的，惟獨祭司才可以吃。
MATT|12|5|再者，律法上所記的，在安息日，祭司在聖殿裏犯了安息日也不算有罪，你們沒有念過嗎？
MATT|12|6|但我告訴你們，比聖殿更大的在這裏。
MATT|12|7|『我喜愛憐憫，不喜愛祭祀。』你們若明白這話的意思，就不將無罪的當作有罪了。
MATT|12|8|因為人子是安息日的主。」
MATT|12|9|耶穌離開那地方，進了 猶太 人的會堂；
MATT|12|10|那裏有個一隻手萎縮了的人。有人為了要控告耶穌，就問他：「安息日治病合不合法？」
MATT|12|11|耶穌對他們說：「你們中間誰有一隻羊在安息日掉在坑裏，不抓住牠，把牠拉上來呢？
MATT|12|12|人比羊貴重得多了！所以，在安息日做善事是合法的。」
MATT|12|13|於是對那人說：「伸出手來！」他把手一伸，手就復原了，和另一隻一樣。
MATT|12|14|法利賽人出去，商議怎樣除掉耶穌。
MATT|12|15|耶穌知道了，就離開那裏，有一大群人跟著他。他把所有的病人都治好了，
MATT|12|16|又囑咐他們不要把他宣揚出去。
MATT|12|17|這是要應驗 以賽亞 先知所說的話：
MATT|12|18|「看哪，我所揀選的僕人， 我所親愛，心所喜悅的； 我要將我的靈賜給他， 他必將公理傳給外邦。
MATT|12|19|他不爭吵，不喧嚷， 街上也沒有人聽見他的聲音。
MATT|12|20|壓傷的蘆葦，他不折斷， 將殘的燈火，他不吹滅， 直到他使公理得勝。
MATT|12|21|外邦人都要仰望他的名。」
MATT|12|22|當時，有人把一個被鬼附，又盲又啞的人帶到耶穌那裏，耶穌醫治他，那啞巴就能說話，又能看見。
MATT|12|23|眾人都驚奇，說：「這不是 大衛 之子嗎？」
MATT|12|24|但法利賽人聽見，就說：「這個人趕鬼，無非是靠著鬼王 別西卜 罷了。」
MATT|12|25|耶穌知道他們的心思，就對他們說：「一國自相紛爭，必定荒蕪；一城一家自相紛爭，必立不住。
MATT|12|26|若撒但趕出撒但，就是自相紛爭，他的國怎能立得住呢？
MATT|12|27|我若靠著 別西卜 趕鬼，你們的子弟趕鬼又靠著誰呢？這樣，他們要作你們的判官。
MATT|12|28|我若靠著上帝的靈趕鬼，那麼，上帝的國就已臨到你們了。
MATT|12|29|人怎能進壯士家裏搶奪他的東西呢？除非先綁住那壯士，否則無法搶奪他的家。
MATT|12|30|不跟我一起的，就是反對我；不與我一起收聚的，就是在拆散。
MATT|12|31|所以我告訴你們，人一切的罪和褻瀆的話都可得赦免，但是褻瀆聖靈，總不得赦免。
MATT|12|32|凡說話干犯人子的，還可得赦免；但是說話干犯聖靈的，今世來世總不得赦免。」
MATT|12|33|「你們知道樹好，果子也好；又知道樹壞，果子也壞；因為看果子就可以知道樹。
MATT|12|34|毒蛇的孽種啊，你們既是惡人，怎能說出好話來呢？因為心裏所充滿的，口裏就說出來。
MATT|12|35|善人從他所存的善發出善來；惡人從他所存的惡發出惡來。
MATT|12|36|我告訴你們，凡是人所說的閒話，在審判的日子，要句句供出來；
MATT|12|37|因為要憑你的話定你為義，也要憑你的話定你有罪。」
MATT|12|38|當時，有幾個文士和法利賽人對耶穌說：「老師，我們想請你顯個神蹟給我們看看。」
MATT|12|39|耶穌回答他們：「邪惡淫亂的世代求看神蹟，除了先知 約拿 的神蹟以外，再沒有神蹟給他們看了。
MATT|12|40|約拿 三日三夜在大魚肚腹中，同樣，人子也要三日三夜在地裏面。
MATT|12|41|在審判的時候， 尼尼微 人要起來定這世代的罪，因為 尼尼微 人聽了 約拿 所傳的就悔改了。看哪，比 約拿 更大的在這裏！
MATT|12|42|在審判的時候，南方的女王要起來定這世代的罪，因為她從地極而來，要聽 所羅門 智慧的話。看哪，比 所羅門 更大的在這裏！」
MATT|12|43|「污靈離了人身，走遍無水之地尋找安歇之處，卻找不到。
MATT|12|44|於是他說：『我要回到我原來的屋裏去。』他到了，看見裏面空著，打掃乾淨，修飾好了，
MATT|12|45|就去另帶了七個比自己更惡的靈來，都進去住在那裏。那人後來的景況比先前更壞了。這邪惡的世代也要如此。」
MATT|12|46|耶穌還在對眾人說話的時候，不料，他母親和他兄弟站在外邊想要跟他說話。
MATT|12|47|有人告訴他：「看哪！你母親和你兄弟站在外邊，想要跟你說話。」
MATT|12|48|他卻回答那對他說話的人，說：「誰是我的母親？誰是我的兄弟？」
MATT|12|49|於是他伸手指著門徒，說：「看哪，我的母親，我的兄弟！
MATT|12|50|凡遵行我天父旨意的人就是我的兄弟、姊妹和母親。」
MATT|13|1|就在那天，耶穌從房子裏出來，坐在海邊。
MATT|13|2|有一大群人到他那裏聚集，他只好上船坐下，眾人都站在岸上。
MATT|13|3|他用比喻對他們講了許多話。他說：「有一個撒種的出去撒種。
MATT|13|4|他撒的時候，有的落在路旁，飛鳥來把它們吃掉了。
MATT|13|5|有的落在土淺的石頭地上，因為土不深，很快就長出苗來，
MATT|13|6|太陽出來一曬，因為沒有根就枯乾了。
MATT|13|7|有的落在荊棘裏，荊棘長起來，把它擠住了。
MATT|13|8|又有的落在好土裏，就結出果實，有一百倍的，有六十倍的，有三十倍的。
MATT|13|9|有耳的，就應當聽！」
MATT|13|10|門徒進前來問耶穌：「對眾人講話，為甚麼用比喻呢？」
MATT|13|11|耶穌回答他們說：「因為天國的奧祕只讓你們知道，不讓他們知道。
MATT|13|12|凡有的，還要給他，讓他有餘；凡沒有的，連他所有的也要奪去。
MATT|13|13|我之所以用比喻對他們講，是因為 他們看卻看不清， 聽卻聽不見，也不明白。
MATT|13|14|在他們身上，正應驗了 以賽亞 的預言： 『你們聽了又聽，卻不明白， 看了又看，卻看不清。
MATT|13|15|因為這百姓的心麻木， 耳朵發沉， 眼睛閉著， 免得眼睛看見， 耳朵聽見， 心裏明白，回轉過來， 我會醫治他們。』
MATT|13|16|但你們的眼睛是有福的，因為看得見；你們的耳朵也是有福的，因為聽得見。
MATT|13|17|我實在告訴你們，從前有許多先知和義人要看你們所看的，卻沒有看見；要聽你們所聽的，卻沒有聽見。」
MATT|13|18|「所以，你們要聽這撒種的比喻。
MATT|13|19|凡聽見天國的道而不明白的，那惡者就來，把撒在他心裏的奪了去；這就是撒在路旁的了。
MATT|13|20|撒在石頭地上的，就是人聽了道，立刻歡喜領受，
MATT|13|21|只因心裏沒有根，不過是暫時的，一旦為道遭受患難或迫害，立刻就跌倒。
MATT|13|22|撒在荊棘裏的，就是人聽了道，後來有世上的憂慮、錢財的迷惑把道擠住了，結不出果實。
MATT|13|23|撒在好土裏的，就是人聽了道，明白了，後來結了果實，有一百倍的，有六十倍的，有三十倍的。」
MATT|13|24|耶穌又設個比喻對他們說：「天國好比人撒好種在田裏，
MATT|13|25|在人睡覺的時候，他的仇敵來，把雜草撒在麥子裏就走了。
MATT|13|26|到長苗吐穗的時候，雜草也顯出來。
MATT|13|27|地主的僕人進前來對他說：『主人，你不是撒好種在田裏嗎？哪裏來的雜草呢？』
MATT|13|28|主人回答他們：『這是仇敵做的。』僕人對他說：『你要我們去拔掉嗎？』
MATT|13|29|主人說：『不必，恐怕拔雜草，也把麥子連根拔出來。
MATT|13|30|讓這兩樣一起長，等到收割。當收割的時候，我會對收割的人說，先把雜草拔出來，捆成捆，留著燒，把麥子收在我的倉裏。』」
MATT|13|31|他又設個比喻對他們說：「天國好比一粒芥菜種，有人拿去種在田裏。
MATT|13|32|它原比所有的種子都小，等到長起來，卻比各樣的菜都大，且成了樹，以致天上的飛鳥來在它的枝上築巢。」
MATT|13|33|他又對他們講另一個比喻：「天國好比麵酵，有婦人拿來放進三斗麵裏，直到全團都發起來。」
MATT|13|34|這都是耶穌用比喻對眾人說的話，不用比喻，他就不對他們說甚麼。
MATT|13|35|這是要應驗先知 所說的話： 「我要開口說比喻， 說出從創世以來所隱藏的事。」
MATT|13|36|當時，耶穌離開眾人，進了屋子。他的門徒進前來，說：「請把田間雜草的比喻講給我們聽。」
MATT|13|37|他回答：「那撒好種的就是人子，
MATT|13|38|田地就是世界，好種就是天國之子，雜草就是那惡者之子，
MATT|13|39|撒雜草的仇敵就是魔鬼，收割的時候就是世代的終結，收割的人就是天使。
MATT|13|40|正如把雜草拔出來用火焚燒，世代的終結也要如此。
MATT|13|41|人子要差遣他的使者，把一切使人跌倒的和作惡的從他國裏挑出來，
MATT|13|42|丟在火爐裏，在那裏要哀哭切齒了。
MATT|13|43|那時，義人要在他們父的國裏發出光來，像太陽一樣。有耳的，就應當聽！」
MATT|13|44|「天國好比寶貝藏在地裏，人發現了就把它藏起來，歡歡喜喜地去變賣一切所有的，買這塊地。
MATT|13|45|「天國又好比商人尋找好的珍珠，
MATT|13|46|發現一顆貴重的珍珠，就去變賣他一切所有的，買下這顆珍珠。」
MATT|13|47|「天國又好比網撒在海裏，聚攏各種魚類，
MATT|13|48|網一滿，人們就把它拉上岸，坐下來，揀好的收在桶裏，不好的丟掉。
MATT|13|49|世代的終結也要這樣：天使要出來，把惡人從義人中分別出來，
MATT|13|50|丟在火爐裏，在那裏要哀哭切齒了。」
MATT|13|51|耶穌說：「這一切的話你們都明白了嗎？」他們對他說：「明白了。」
MATT|13|52|他對他們說：「凡文士學習作天國的門徒，就像一個家的主人從他庫裏拿出新的和舊的東西來。」
MATT|13|53|耶穌說完了這些比喻，就離開那裏，
MATT|13|54|來到自己的家鄉，在會堂裏教導人，以致他們都很驚奇，說：「這人哪來這樣的智慧和異能呢？
MATT|13|55|這不是那木匠的兒子嗎？他母親不是叫 馬利亞 嗎？他兄弟們不是叫 雅各 、 約瑟 、 西門 、 猶大 嗎？
MATT|13|56|他姊妹們不是都在我們這裏嗎？他這一切是從哪裏來的呢？」
MATT|13|57|他們就厭棄他。耶穌對他們說：「先知除了在本鄉和自己的家之外，沒有不被尊敬的。」
MATT|13|58|耶穌因為他們不信，沒有在那裏行很多異能。
MATT|14|1|那時， 希律 分封王聽見耶穌的名聲，
MATT|14|2|就對臣僕說：「這是施洗的 約翰 從死人中復活，因此才有這些異能在他裏面運行。」
MATT|14|3|原來， 希律 為他兄弟 腓力 的妻子 希羅底 的緣故，把 約翰 抓住綁了，關進監獄，
MATT|14|4|因為 約翰 曾對他說：「你佔有這婦人是不合法的。」
MATT|14|5|希律 就想要殺他，可是怕民眾，因為他們認為 約翰 是先知。
MATT|14|6|到了 希律 的生日， 希羅底 的女兒在眾人面前跳舞，使 希律 歡喜，
MATT|14|7|於是 希律 發誓許諾隨她所求的給她。
MATT|14|8|女兒被母親指使，就說：「請把施洗 約翰 的頭放在盤子裏，拿來給我。」
MATT|14|9|王就憂愁，然而因他所發的誓，又因同席的人，就下令給她；
MATT|14|10|於是打發人去，在監獄裏斬了 約翰 ，
MATT|14|11|把頭放在盤子裏，拿來給那女孩，她拿去給她母親。
MATT|14|12|約翰 的門徒來，把屍體領去埋葬了，又去告訴耶穌。
MATT|14|13|耶穌聽到了，就從那裏上船，私下退到荒野的地方去。眾人聽到後，從各城來，步行跟隨他。
MATT|14|14|耶穌出來，見有一大群人，就憐憫他們，治好了他們的病人。
MATT|14|15|傍晚的時候，門徒進前來，說：「這地方偏僻，而且時候已經晚了，請叫眾人散去，他們好進村子，自己買些食物。」
MATT|14|16|耶穌對他們說：「不用他們去，你們給他們吃吧！」
MATT|14|17|門徒說：「我們這裏只有五個餅、兩條魚。」
MATT|14|18|耶穌說：「拿過來給我。」
MATT|14|19|於是他吩咐眾人坐在草地上，就拿著這五個餅和兩條魚，望著天祝福，擘開餅，遞給門徒，門徒又遞給眾人。
MATT|14|20|他們都吃，並且吃飽了。門徒把剩下的碎屑收拾起來，裝滿了十二個籃子。
MATT|14|21|吃的人中，男的約有五千，還不算婦女和孩子。
MATT|14|22|耶穌隨即催門徒上船，先渡到對岸，等他叫眾人散去。
MATT|14|23|疏散了眾人以後，他獨自上山去禱告。到了晚上，只有他一人在那裏。
MATT|14|24|那時船已離岸好幾里 ，因風不順，被浪顛簸。
MATT|14|25|天快亮的時候，耶穌在海面上走，往門徒那裏去。
MATT|14|26|但門徒看見他在海面上走，就驚慌了，說：「是個鬼怪！」他們害怕得喊叫起來。
MATT|14|27|耶穌連忙對他們說：「放心！是我，不要怕！」
MATT|14|28|彼得 回答他說：「主啊，如果是你，請叫我從水面上走到你那裏去。」
MATT|14|29|耶穌說：「你來吧！」 彼得 就從船上下去，在水面上走，往耶穌那裏去；
MATT|14|30|只因見風很強 ，害怕起來，將要沉下去，就喊著說：「主啊，救我！」
MATT|14|31|耶穌立刻伸手拉住他，說：「你這小信的人哪，為甚麼疑惑呢？」
MATT|14|32|他們一上船，風就停了。
MATT|14|33|在船上的人都拜他，說：「你真是上帝的兒子。」
MATT|14|34|他們渡過了海，在 革尼撒勒 上岸。
MATT|14|35|那裏的人認出耶穌，就打發人到整個周圍地區去，把所有的病人帶到他那裏，
MATT|14|36|求耶穌讓他們只摸一摸他的衣裳繸子，摸著的人就都好了。
MATT|15|1|那時，有法利賽人和文士從 耶路撒冷 來見耶穌，說：
MATT|15|2|「你的門徒為甚麼違反古人的傳統？因為他們吃飯的時候不洗手。」
MATT|15|3|耶穌回答他們：「你們為甚麼因你們的傳統而違反上帝的誡命呢？
MATT|15|4|上帝說：『當孝敬父母』；又說：『咒罵父母的，必須處死。』
MATT|15|5|你們倒說：『無論誰對父母說：我所當供奉你的已經作了奉獻，
MATT|15|6|就可以不孝敬他的父親 。』這就是你們藉著傳統，廢了上帝的話。
MATT|15|7|假冒為善的人哪！ 以賽亞 指著你們所預言的說得好：
MATT|15|8|『這百姓用嘴唇尊敬我， 他們的心卻遠離我。
MATT|15|9|他們把人的規條當作教義教導人； 他們拜我也是枉然。』」
MATT|15|10|耶穌叫了眾人來，對他們說：「你們要聽，也要明白。
MATT|15|11|從口裏進去的不玷污人，從口裏出來的才玷污人。」
MATT|15|12|當時，門徒進前來對他說：「法利賽人聽見這話很反感，你知道嗎？」
MATT|15|13|耶穌回答：「一切植物，若不是我天父栽植的，都要連根拔出來。
MATT|15|14|由他們吧！他們是瞎子作瞎子的嚮導 ；若是瞎子領瞎子，兩個人都要掉在坑裏。」
MATT|15|15|彼得 回應他說：「請將這比喻講解給我們聽。」
MATT|15|16|耶穌說：「連你們也還不明白嗎？
MATT|15|17|難道你們不了解，凡進到口裏的，是經過肚子，又排入廁所嗎？
MATT|15|18|然而口裏出來的是出於心裏，這才玷污人。
MATT|15|19|因為出於心裏的有種種惡念，如兇殺、姦淫、淫亂、偷盜、偽證、毀謗。
MATT|15|20|這些才玷污人。至於不洗手吃飯，那並不玷污人。」
MATT|15|21|耶穌離開那裏，退到 推羅 、 西頓 境內。
MATT|15|22|有一個 迦南 婦人從那地方出來，喊著說：「主啊， 大衛 之子，可憐我！我女兒被鬼纏得很苦。」
MATT|15|23|耶穌卻一言不答。門徒進前來，求他說：「這婦人在我們後頭喊叫，請打發她走吧。」
MATT|15|24|耶穌回答：「我奉差遣只到 以色列 家迷失的羊那裏去。」
MATT|15|25|那婦人來拜他，說：「主啊，幫幫我！」
MATT|15|26|他回答：「拿孩子的餅丟給小狗吃是不妥的。」
MATT|15|27|婦人說：「主啊，不錯，可是小狗也吃牠主人桌上掉下來的碎屑。」
MATT|15|28|於是耶穌回答她說：「婦人，你的信心很大！照你所要的成全你吧。」從那時起，她的女兒就好了。
MATT|15|29|耶穌離開那地方，來到靠近 加利利 的海邊，就上山坐下。
MATT|15|30|有一大群人到他那裏，帶著瘸子、盲人、肢殘的、聾啞的，和好些別的病人，都放在他腳前，他就治好了他們。
MATT|15|31|於是眾人都驚訝，因為看見聾啞的說話，肢殘的痊癒，瘸子行走，盲人看見，他們就歸榮耀給 以色列 的上帝。
MATT|15|32|耶穌叫門徒來，說：「我憐憫這群人，因為他們同我在這裏已經三天，沒有吃的東西了。我不願意叫他們餓著回去，恐怕他們在路上餓昏了。」
MATT|15|33|門徒說：「我們在這野地，哪裏有這麼多的餅讓這許多人吃飽呢？」
MATT|15|34|耶穌對他們說：「你們有多少餅？」他們說：「有七個，還有幾條小魚。」
MATT|15|35|他就吩咐眾人坐在地上，
MATT|15|36|拿著這七個餅和幾條魚，祝謝了，擘開，遞給門徒；門徒又遞給眾人。
MATT|15|37|他們都吃，並且吃飽了，收拾剩下的碎屑，裝滿了七個筐子。
MATT|15|38|吃的人中，男的有四千，還不算婦女和孩子。
MATT|15|39|耶穌叫眾人散去，就上船，來到 馬加丹 境內。
MATT|16|1|法利賽人和撒都該人來試探耶穌，請他顯個來自天上的神蹟給他們看。
MATT|16|2|耶穌回答他們：「傍晚天發紅，你們就說：『明日天晴。』
MATT|16|3|早晨天色又紅又暗，你們就說：『今日有風雨。』你們知道分辨天上的氣象，倒不能分辨這個時代的神蹟 。
MATT|16|4|邪惡淫亂的世代求看神蹟，除了 約拿 的神蹟以外，再沒有神蹟給他們看了。」於是耶穌離開他們走了。
MATT|16|5|門徒渡到對岸，忘了帶餅。
MATT|16|6|耶穌對他們說：「你們要謹慎，要防備法利賽人和撒都該人的酵。」
MATT|16|7|門徒彼此議論說：「這是因為我們沒有帶餅吧。」
MATT|16|8|耶穌知道了，就說：「你們這小信的人，為甚麼因為沒有餅就彼此議論呢？
MATT|16|9|你們還不明白嗎？不記得那五個餅分給五千人，你們收拾了多少籃子的碎屑嗎？
MATT|16|10|也不記得那七個餅分給四千人，你們又收拾了多少筐子的碎屑嗎？
MATT|16|11|我對你們說『要防備法利賽人和撒都該人的酵』，這話不是指著餅說的，你們怎麼不明白呢？」
MATT|16|12|門徒這才明白他所說的不是要他們防備餅的酵 ，而是要防備法利賽人和撒都該人的教訓。
MATT|16|13|耶穌到了 凱撒利亞．腓立比 的境內，就問門徒：「人們說人子是誰？」
MATT|16|14|他們說：「有人說是施洗的 約翰 ；有人說是 以利亞 ；又有人說是 耶利米 或是先知中的一位。」
MATT|16|15|耶穌問他們：「你們說我是誰？」
MATT|16|16|西門．彼得 回答說：「你是基督，是永生上帝的兒子。」
MATT|16|17|耶穌回答他說：「 約拿 的兒子 西門 ，你是有福的！因為這不是屬血肉的啟示你的，而是我在天上的父啟示的。
MATT|16|18|我還告訴你，你是 彼得 ，我要把我的教會建造在這磐石上，陰間的權柄不能勝過它。
MATT|16|19|我要把天國的鑰匙給你，凡你在地上所捆綁的，在天上也要捆綁；凡你在地上所釋放的，在天上也要釋放。」
MATT|16|20|當時，耶穌囑咐門徒不可對任何人說他是基督。
MATT|16|21|從那時起，耶穌才向門徒明說，他必須上 耶路撒冷 去，受長老、祭司長和文士許多的苦，並且被殺，第三天復活。
MATT|16|22|彼得 就拉著他，責備他說：「主啊，千萬不可如此！這事絕不可臨到你身上。」
MATT|16|23|耶穌轉過來，對 彼得 說：「撒但，退到我後邊去！你是我的絆腳石，因為你不體會上帝的心意，而是體會人的意思。」
MATT|16|24|於是耶穌對門徒說：「若有人要跟從我，就當捨己，背起自己的十字架來跟從我。
MATT|16|25|因為凡要救自己生命的，要喪失生命；凡為我喪失生命的，要得著生命。
MATT|16|26|人若賺得全世界，賠上自己的生命，有甚麼益處呢？人還能拿甚麼換生命呢？
MATT|16|27|人子要在他父的榮耀裏與他的眾使者一起來臨，那時候，他要照各人的行為報應各人。
MATT|16|28|我實在告訴你們，站在這裏的，有人在沒經歷死亡以前，必定看見人子來到他的國裏。」
MATT|17|1|過了六天，耶穌帶著 彼得 、 雅各 和 雅各 的弟弟 約翰 ，領他們悄悄地上了高山。
MATT|17|2|他在他們面前變了形像，他的臉明亮如太陽，衣裳潔白如光。
MATT|17|3|忽然，有 摩西 和 以利亞 向他們顯現，與耶穌說話。
MATT|17|4|彼得 回應，對耶穌說：「主啊，我們在這裏真好！你若願意，我就在這裏搭三座棚，一座為你，一座為 摩西 ，一座為 以利亞 。」
MATT|17|5|說話之間，忽然有一朵明亮的雲彩遮蓋他們，又有聲音從雲彩裏出來，說：「這是我的愛子，我所喜愛的。你們要聽從他！」
MATT|17|6|門徒聽見，就俯伏在地，極其害怕。
MATT|17|7|耶穌進前來，拍拍他們，說：「起來，不要害怕！」
MATT|17|8|他們舉目，不見一人，只見耶穌獨自一人。
MATT|17|9|下山的時候，耶穌囑咐他們說：「人子還沒有從死人中復活，你們不要把所看到的告訴人。」
MATT|17|10|門徒問耶穌：「那麼，文士為甚麼說 以利亞 必須先來？」
MATT|17|11|耶穌回答：「 以利亞 的確要來，並要復興萬事；
MATT|17|12|可是我告訴你們， 以利亞 已經來了，人不認識他，反倒任意待他。人子也將這樣受他們的苦。」
MATT|17|13|門徒這才明白耶穌所說的是指施洗的 約翰 。
MATT|17|14|耶穌和門徒到了眾人那裏，有一個人來見耶穌，跪下，
MATT|17|15|說：「主啊，可憐我的兒子。他害癲癇病很苦，屢次跌進火裏，屢次跌進水裏。
MATT|17|16|我帶他到你門徒那裏，他們卻不能醫治他。」
MATT|17|17|耶穌回答：「唉！這又不信又悖謬的世代啊，我和你們在一起要到幾時呢？我忍耐你們要到幾時呢？把他帶到我這裏來！」
MATT|17|18|耶穌斥責那鬼，鬼就出來；從那時起，孩子就痊癒了。
MATT|17|19|門徒私下進前來問耶穌：「我們為甚麼不能趕出那鬼呢？」
MATT|17|20|耶穌對他們說：「是因你們的信心小。我實在告訴你們，你們若有信心像一粒芥菜種，就是對這座山說：『你從這邊移到那邊』，它也會移過去，並且你們沒有一件不能做的事了。 」
MATT|17|21|
MATT|17|22|他們聚集在 加利利 的時候，耶穌對門徒說：「人子將要被交在人手裏。
MATT|17|23|他們要殺害他，第三天他要復活。」門徒就非常憂愁。
MATT|17|24|他們到了 迦百農 ，收聖殿稅 的人來見 彼得 ，說：「你們的老師不納聖殿稅嗎？」
MATT|17|25|彼得 說：「納。」他進了屋子，耶穌先對他說：「 西門 ，你的意見如何？世上的君王向誰徵收關稅或丁稅？是向自己的兒子呢？還是向外人呢？」
MATT|17|26|彼得 說：「是向外人。」耶穌對他說：「既然如此，兒子就可以免了。
MATT|17|27|但恐怕觸犯他們，你往海邊去釣魚，把先釣上來的魚拿起來，開了牠的口，會發現一個司塔特 ，可以拿去給他們，作你我的稅錢。」
MATT|18|1|當時，門徒前來問耶穌：「天國裏誰是最大的？」
MATT|18|2|耶穌叫一個小孩子來，讓他站在他們當中，
MATT|18|3|說：「我實在告訴你們，你們若不回轉，變成像小孩子一樣，絕不能進天國。
MATT|18|4|所以，凡自己謙卑像這小孩子的，他在天國裏就是最大的。
MATT|18|5|凡為我的名接納一個像這小孩子的，就是接納我。」
MATT|18|6|「凡使這些信我的小子中的一個跌倒的，倒不如把大磨石拴在這人的頸項上，沉在深海裏。
MATT|18|7|這世界有禍了，因為它使人跌倒；絆倒人的事是免不了的，但那絆倒人的有禍了！
MATT|18|8|如果你一隻手或是一隻腳使你跌倒，就把它砍下來扔掉。你缺一隻手或是一隻腳進入永生，比有兩手兩腳被扔進永火裏還好。
MATT|18|9|如果你一隻眼使你跌倒，就把它挖出來扔掉。你只有一隻眼進入永生，比有兩隻眼被扔進地獄的火裏還好。」
MATT|18|10|「你們要小心，不可輕看這些小子中的一個；我告訴你們，他們的天使在天上，常見我天父的面。
MATT|18|11|
MATT|18|12|「一個人若有一百隻羊，其中一隻走迷了路，你們的意見如何？他豈不留下這九十九隻在山上，去找那隻迷路的羊嗎？
MATT|18|13|若是找到了，我實在告訴你們，他為這一隻羊歡喜，比為那沒有迷路的九十九隻歡喜還大呢！
MATT|18|14|你們 在天上的父也是這樣，不願意失去這些小子中的一個。」
MATT|18|15|「若是你的弟兄得罪你 ，你要去，趁著只有他和你在一起的時候，指出他的錯來。他若聽你，你就贏得了你的弟兄；
MATT|18|16|他若不聽，你就另外帶一個或兩個人同去，因為『任何指控都要憑兩個或三個證人的口述才能成立』。
MATT|18|17|他若是不聽他們，就去告訴教會；若是不聽教會，就把他看作外邦人和稅吏。
MATT|18|18|「我實在告訴你們，凡你們在地上所捆綁的，在天上也要捆綁；凡你們在地上所釋放的，在天上也要釋放。
MATT|18|19|我又實在 告訴你們，若是你們中間有兩個人在地上同心合意地求甚麼事，我在天上的父必為他們成全。
MATT|18|20|因為，哪裏有兩三個人奉我的名聚會，哪裏就有我在他們中間。」
MATT|18|21|那時， 彼得 進前來，對耶穌說：「主啊，我弟兄得罪我，我當饒恕他幾次呢？到七次夠嗎？」
MATT|18|22|耶穌說：「我告訴你，不是到七次，而是到七十個七次。
MATT|18|23|因為天國好像一個王要和他僕人算賬。
MATT|18|24|他開始算的時候，有人帶了一個欠一萬他連得的僕人來。
MATT|18|25|因為他沒有甚麼償還之物，主人下令把他和他妻子兒女，以及一切所有的都賣了來償還。
MATT|18|26|那僕人就俯伏向他叩頭，說：『寬容我吧，我都會還你的。』
MATT|18|27|那僕人的主人就動了慈心，把他釋放了，並且免了他的債。
MATT|18|28|那僕人出來，遇見一個欠他一百個銀幣的同伴，就揪著他，扼住他的喉嚨，說：『把你所欠的還我！』
MATT|18|29|他的同伴就俯伏央求他，說：『寬容我吧，我會還你的。』
MATT|18|30|他不肯，卻把他下在監裏，直到他還了所欠的債。
MATT|18|31|同伴們看見他所做的事就很悲憤，把這一切的事都告訴了主人。
MATT|18|32|於是主人叫了他來，對他說：『你這惡奴才！你央求我，我就把你所欠的都免了；
MATT|18|33|你不應該憐憫你的同伴，像我憐憫你嗎？』
MATT|18|34|主人就大怒，把他交給司刑的，直到他還清了所欠的債。
MATT|18|35|你們各人若不從心裏饒恕你的弟兄，我天父也要這樣待你們。」
MATT|19|1|耶穌說完了這些話，就離開 加利利 ，來到 猶太 的境內、 約旦河 的東邊。
MATT|19|2|有一大群人跟著他，他就在那裏治好了他們。
MATT|19|3|有些法利賽人來試探耶穌說：「無論甚麼緣故，人休妻都合法嗎？」
MATT|19|4|耶穌回答：「那起初造人的，是造男造女，並且說：『因此，人要離開父母，與妻子結合，二人成為一體。』這經文你們沒有念過嗎？
MATT|19|5|
MATT|19|6|既然如此，夫妻不再是兩個人，而是一體的了。所以，上帝配合的，人不可分開。」
MATT|19|7|法利賽人說：「這樣， 摩西 為甚麼吩咐給妻子休書就可以休她呢？」
MATT|19|8|耶穌說：「 摩西 因為你們的心硬，所以准許你們休妻，但起初並不是這樣。
MATT|19|9|我告訴你們，凡休妻另娶的，若不是為不貞的緣故，就是犯姦淫了。 」
MATT|19|10|門徒對耶穌說：「丈夫和妻子的關係既是這樣，倒不如不娶。」
MATT|19|11|耶穌對他們說：「這話不是人人都能領受的，惟獨賜給誰，誰才能領受。
MATT|19|12|因為有人從母腹裏就是不宜結婚的，也有因人為的緣故不宜結婚的，並有為天國的緣故自己不結婚的 。這話誰能領受，就領受吧。」
MATT|19|13|那時，有人帶著小孩子來見耶穌，要他給他們按手禱告，門徒就責備那些人。
MATT|19|14|耶穌說：「讓小孩子到我這裏來，不要阻止他們，因為在天國的正是這樣的人。」
MATT|19|15|耶穌給他們按手，然後離開那地方。
MATT|19|16|有一個人進前來問耶穌：「老師，我該做甚麼善事才能得永生？」
MATT|19|17|耶穌對他說：「你為甚麼問我關於善的事呢？只有一位是善良的。你若要進入永生，就該遵守誡命。」
MATT|19|18|他說：「哪些誡命？」耶穌說：「就是不可殺人；不可姦淫；不可偷盜；不可作假見證；
MATT|19|19|當孝敬父母；又當愛鄰 如己。」
MATT|19|20|那青年說：「這一切我都遵守了，還缺少甚麼呢？」
MATT|19|21|耶穌說：「你若願意作完全人，去變賣你所擁有的，分給窮人，就必有財寶在天上；然後來跟從我。」
MATT|19|22|那青年聽見這話，就憂憂愁愁地走了，因為他的產業很多。
MATT|19|23|耶穌對門徒說：「我實在告訴你們，財主進天國是難的。
MATT|19|24|我再告訴你們，駱駝穿過針眼比財主進上帝的國還容易呢！」
MATT|19|25|門徒聽見這話，就非常驚奇，說：「這樣，誰能得救呢？」
MATT|19|26|耶穌看著他們，說：「在人這是不能，在上帝凡事都能。」
MATT|19|27|於是 彼得 回應，對他說：「看哪，我們已經撇下一切跟從你了，我們會得到甚麼呢？」
MATT|19|28|耶穌對他們說：「我實在告訴你們，你們這些跟從我的人，到了萬物更新、人子坐在他榮耀寶座上的時候，你們也要坐在十二個寶座上，審判 以色列 十二個支派。
MATT|19|29|凡為我的名撇下房屋，或是兄弟、姊妹、父親、母親、 兒女、田地的，將得著百倍，並且承受永生。
MATT|19|30|然而，有許多在前的，將要在後；在後的，將要在前。」
MATT|20|1|「因為天國好比一家的主人清早去雇人進他的葡萄園做工。
MATT|20|2|他和工人講定一天一個銀幣 ，就打發他們進葡萄園去。
MATT|20|3|約在上午九點鐘出去，看見市場上還有閒站的人，
MATT|20|4|就對那些人說：『你們也進葡萄園去，我會給你們合理的工錢。』
MATT|20|5|他們也進去了。約在正午和下午三點鐘又出去，他也是這麼做。
MATT|20|6|約在下午五點鐘出去，他看見還有人站在那裏，就問他們：『你們為甚麼整天在這裏閒站呢？』
MATT|20|7|他們說：『因為沒有人雇我們。』他說：『你們也進葡萄園去。』
MATT|20|8|到了晚上，園主對工頭說：『叫工人都來，給他們工錢，從後來的起，到先來的為止。』
MATT|20|9|約在下午五點鐘雇的人來了，各人領了一個銀幣。
MATT|20|10|那些最先雇的來了，以為可以多領，誰知也是各領一個銀幣。
MATT|20|11|他們領了工錢，就埋怨那家的主人說：
MATT|20|12|『我們整天勞苦受熱，那些後來的只做了一小時，你竟待他們和我們一樣嗎？』
MATT|20|13|主人回答其中的一人說：『朋友，我沒虧待你，你與我講定的不是一個銀幣嗎？
MATT|20|14|拿你的錢走吧！我樂意給那後來的和給你的一樣，
MATT|20|15|難道我的東西不可隨我的意思用嗎？因為我作好人，你就眼紅了嗎？』
MATT|20|16|這樣，那在後的，將要在前；在前的，將要在後了。」
MATT|20|17|耶穌上 耶路撒冷 去的時候，在路上把十二個門徒帶到一邊，對他們說：
MATT|20|18|「看哪，我們上 耶路撒冷 去，人子將被交給祭司長和文士；他們要定他死罪，
MATT|20|19|把他交給外邦人戲弄，鞭打，釘在十字架上；第三天他要復活。」
MATT|20|20|那時， 西庇太 兒子的母親和她兩個兒子上前來，向耶穌叩頭，求他一件事。
MATT|20|21|耶穌問她：「你要甚麼呢？」她對耶穌說：「在你的國裏，請讓我這兩個兒子一個坐在你右邊，一個坐在你左邊。」
MATT|20|22|耶穌回答：「你們不知道所求的是甚麼。我將要喝的杯，你們能喝嗎？」他們對他說：「我們能。」
MATT|20|23|耶穌說：「我所喝的杯，你們要喝。可是坐在我的左右，不是我可以賜的，而是我父為誰預備就賜給誰。」
MATT|20|24|其餘十個門徒聽見，就對他們兄弟二人很生氣。
MATT|20|25|耶穌叫了他們來，說：「你們知道，外邦人有君王作主治理他們，有大臣操權管轄他們。
MATT|20|26|但是在你們中間，不可這樣。你們中間誰願為大，就要作你們的用人；
MATT|20|27|誰願為首，就要作你們的僕人。
MATT|20|28|正如人子來，不是要受人的服事，乃是要服事人，並且要捨命，作多人的贖價。」
MATT|20|29|他們出 耶利哥 的時候，有一大群人跟隨耶穌。
MATT|20|30|有兩個盲人坐在路旁，聽說是耶穌經過，就喊著說：「主啊 ， 大衛 之子，可憐我們吧！」
MATT|20|31|眾人責備他們，不許他們作聲，他們卻越發喊著說：「主啊 ， 大衛 之子，可憐我們吧！」
MATT|20|32|耶穌就站住，叫他們來，說：「你們要我為你們做甚麼？」
MATT|20|33|他們說：「主啊，讓我們的眼睛能看見。」
MATT|20|34|耶穌動了慈心，摸了他們的眼睛，他們立刻看得見，就跟從耶穌。
MATT|21|1|耶穌和門徒快到 耶路撒冷 ，進了 橄欖山 的 伯法其 時，打發兩個門徒，
MATT|21|2|對他們說：「你們往對面村子裏去，會立刻看見一匹驢拴在那裏，還有驢駒同在一處，解開牠們，牽到我這裏來。
MATT|21|3|若有人對你們說甚麼，你們就說：『主要用牠們。』那人會立刻讓你們牽來。」
MATT|21|4|這事發生是要應驗先知所說的話：
MATT|21|5|「要對 錫安 的兒女 說： 看哪，你的王來到你這裏， 謙和地騎著驢， 騎著小驢—驢的駒子。」
MATT|21|6|門徒就照耶穌所吩咐的去做，
MATT|21|7|牽了驢和驢駒來，把他們的衣服搭在上面，耶穌就騎上。
MATT|21|8|許許多多的人把自己的衣服鋪在路上，還有人砍下樹枝來鋪在路上。
MATT|21|9|前呼後擁的人群喊著說： 「和散那 歸於 大衛 之子！ 奉主名來的是應當稱頌的！ 至高無上的，和散那！」
MATT|21|10|耶穌進了 耶路撒冷 ，全城都驚動了，說：「這是誰？」
MATT|21|11|眾人說：「這是從 加利利 的 拿撒勒 來的先知耶穌。」
MATT|21|12|耶穌進了聖殿 ，趕出聖殿裏所有在做買賣的人，推倒兌換銀錢之人的桌子和賣鴿子之人的凳子，
MATT|21|13|對他們說：「經上記著： 『我的殿要稱為禱告的殿， 你們倒使它成為賊窩了。』」
MATT|21|14|在聖殿裏有盲人和瘸子到耶穌跟前，他就治好了他們。
MATT|21|15|祭司長和文士看見耶穌所行的奇事，又見小孩子在聖殿裏喊著說：「和散那歸於 大衛 之子！」就很生氣，
MATT|21|16|對他說：「這些人所喊的，你聽到了嗎？」耶穌對他們說：「聽到了。經上說：『你藉孩童和吃奶的口發出完全的讚美』，你們沒有念過嗎？」
MATT|21|17|於是他離開他們，出城到 伯大尼 去，在那裏過夜。
MATT|21|18|早晨回城的時候，他餓了，
MATT|21|19|看見路旁有一棵無花果樹，就走到跟前，在樹上找不到甚麼，只有葉子，就對樹說：「從今以後，你永不結果子！」那無花果樹立刻枯乾了。
MATT|21|20|門徒看見了，驚訝地說：「無花果樹怎麼立刻枯乾了呢？」
MATT|21|21|耶穌回答他們：「我實在告訴你們，你們若有信心，不疑惑，不但能行我對無花果樹所行的事，就是對這座山說：『離開此地，投在海裏！』也會實現。
MATT|21|22|你們禱告，無論求甚麼，只要信，就必得著。」
MATT|21|23|耶穌進了聖殿，正教導人的時候，祭司長和百姓的長老來問他：「你仗著甚麼權柄做這些事？給你這權柄的是誰呢？」
MATT|21|24|耶穌回答他們說：「我也要問你們一句話，你們若告訴我，我就告訴你們我仗著甚麼權柄做這些事。
MATT|21|25|約翰 的洗禮是從哪裏來的？是從天上來的，還是從人間來的呢？」他們彼此商議說：「我們若說『從天上來的』，他會對我們說：『這樣，你們為甚麼不信他呢？』
MATT|21|26|若說『從人間來的』，我們又怕眾人，因為大家都認為 約翰 是先知。」
MATT|21|27|於是他們回答耶穌：「我們不知道。」耶穌也對他們說：「我也不告訴你們，我仗著甚麼權柄做這些事。」
MATT|21|28|「有一件事，你們的意見如何？一個人有兩個兒子。他來對大兒子說：『孩子，今天到葡萄園裏做工去。』
MATT|21|29|他回答：『我不去』，以後自己懊悔，就去了。
MATT|21|30|他來對小兒子也是這樣說。他回答：『父親大人，我去』，卻不去。
MATT|21|31|這兩個兒子是哪一個照著父親的意願做了呢？」他們說：「大兒子。」耶穌說：「我實在告訴你們，稅吏和娼妓倒比你們先進上帝的國。
MATT|21|32|因為 約翰 到你們這裏來指引你們走義路，你們卻不信他，稅吏和娼妓倒信了他。你們看見了以後，還是不悔悟去信他。」
MATT|21|33|「你們再聽一個比喻：有一個家的主人開墾了一個葡萄園，四周圍上籬笆，裏面挖了一個榨酒池，蓋了一座守望樓，租給園戶，就出外遠行去了。
MATT|21|34|收果子的時候快到了，他打發僕人到園戶那裏去收果子。
MATT|21|35|園戶拿住僕人，打了一個，殺了一個，用石頭打死了一個。
MATT|21|36|主人又打發別的僕人去，比先前更多；園戶還是照樣對待他們。
MATT|21|37|最後他打發自己的兒子到他們那裏去，說：『他們會尊敬我的兒子。』
MATT|21|38|可是，園戶看見他兒子，彼此說：『這是承受產業的。來，我們殺了他，佔他的產業！』
MATT|21|39|於是他們拿住他，把他扔出葡萄園外，殺了。
MATT|21|40|葡萄園的主人來的時候，要怎樣處置那些園戶呢？」
MATT|21|41|他們說：「要狠狠地除滅那些惡人，將葡萄園轉租給那些按時候交果子的園戶。」
MATT|21|42|耶穌對他們說： 「『匠人所丟棄的石頭 已作了房角的頭塊石頭。 這是主所做的， 在我們眼中看為奇妙。』 這段經文你們從來沒有念過嗎？
MATT|21|43|所以我告訴你們，上帝的國必從你們奪去，賜給那能結果子的民。
MATT|21|44|誰跌在這石頭上，一定會跌得粉碎；這石頭掉在誰的身上，就要把誰壓得稀爛。 」
MATT|21|45|祭司長和法利賽人聽見他的比喻，就看出他是指著他們說的。
MATT|21|46|他們想要捉拿他，但是懼怕眾人，因為眾人認為他是先知。
MATT|22|1|耶穌又用比喻對他們說：
MATT|22|2|「天國好比一個王為他兒子擺設娶親的宴席。
MATT|22|3|他打發僕人去，請那些被邀的人來赴宴，他們卻不肯來。
MATT|22|4|王又打發別的僕人，說：『你們去告訴那被邀的人，我的宴席已經預備好了，牛和肥畜已經宰了，各樣都齊備，請你們來赴宴。』
MATT|22|5|那些人不理就走了，一個到自己田裏去，一個做買賣去。
MATT|22|6|其餘的抓住僕人，凌辱他們，把他們殺了。
MATT|22|7|王就大怒，發兵除滅那些兇手，燒燬他們的城。
MATT|22|8|於是王對僕人說：『喜宴已經齊備，只是所邀的人不配。
MATT|22|9|所以你們要往岔路口上去，凡遇見的，都邀來赴宴。』
MATT|22|10|那些僕人就出去，到大路上，凡遇見的，不論善惡都招聚了來，宴席上就坐滿了客人。
MATT|22|11|王進來見賓客，看到那裏有一個沒有穿禮服的，
MATT|22|12|就對他說：『朋友，你到這裏來怎麼不穿禮服呢？』那人無言可答。
MATT|22|13|於是王對侍從說：『捆起他的手腳，把他扔在外邊的黑暗裏；在那裏他要哀哭切齒了。』
MATT|22|14|因為被召的人多，選上的人少。」
MATT|22|15|於是，法利賽人出去商議，怎樣找話柄來陷害耶穌，
MATT|22|16|就打發他們的門徒同 希律 黨人去見耶穌，說：「老師，我們知道你是誠實的，並且誠誠實實傳上帝的道，無論誰你都一視同仁，因為你不看人的面子。
MATT|22|17|請告訴我們，你的意見如何？納稅給凱撒合不合法？」
MATT|22|18|耶穌看出他們的惡意，就說：「假冒為善的人哪，為甚麼試探我？
MATT|22|19|拿一個納稅的錢給我看！」他們就拿一個銀幣來給他。
MATT|22|20|耶穌問他們：「這像和這名號是誰的？」
MATT|22|21|他們說：「是凱撒的。」於是耶穌說：「這樣，凱撒的歸凱撒；上帝的歸上帝。」
MATT|22|22|他們聽了十分驚訝，就離開他走了。
MATT|22|23|那天，撒都該人來見耶穌。他們說沒有復活這回事，於是問耶穌：
MATT|22|24|「老師， 摩西 說：『某人若死了，沒有孩子，他弟弟該娶他的妻子，為哥哥生子立後。』
MATT|22|25|從前，在我們這裏有兄弟七人，第一個娶了妻，死了，沒有孩子，撇下妻子給弟弟。
MATT|22|26|第二、第三，直到第七個，都是如此。
MATT|22|27|後來，那婦人也死了。
MATT|22|28|那麼，在復活的時候，她是七個人中哪一個的妻子呢？因為他們都娶過她。」
MATT|22|29|耶穌回答他們說：「你們錯了，因為不明白聖經，也不知道上帝的大能。
MATT|22|30|在復活的時候，人也不娶也不嫁，而是像天上的天使一樣。
MATT|22|31|論到死人復活，上帝向你們所說的話，你們沒有念過嗎？
MATT|22|32|他說：『我是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。』上帝不是死人的上帝，而是活人的上帝。」
MATT|22|33|眾人聽見這話，對他的教導非常驚訝。
MATT|22|34|法利賽人聽見耶穌堵住了撒都該人的口，他們就聚集在一起。
MATT|22|35|其中有一個人是律法師 ，要試探耶穌，就問他：
MATT|22|36|「老師，律法上的誡命哪一條是最大的呢？」
MATT|22|37|耶穌對他說：「你要盡心、盡性、盡意愛主—你的上帝。
MATT|22|38|這是最大的，且是第一條誡命。
MATT|22|39|第二條也如此，就是要愛鄰 如己。
MATT|22|40|這兩條誡命是一切律法和先知書的總綱。」
MATT|22|41|法利賽人聚集的時候，耶穌問他們：
MATT|22|42|「論到基督，你們的意見如何？他是誰的後裔呢？」他們說：「是 大衛 的。」
MATT|22|43|耶穌說：「這樣， 大衛 被聖靈感動，怎麼還稱他為主，說：
MATT|22|44|『主對我主說： 你坐在我的右邊， 等我把你的仇敵放在你腳下？』
MATT|22|45|大衛 既稱他為主，他怎麼又是 大衛 的後裔呢？」
MATT|22|46|沒有一個人能回答一句話，從那日以後沒有人敢再問他甚麼。
MATT|23|1|那時，耶穌對眾人和門徒講論，
MATT|23|2|說：「文士和法利賽人坐在 摩西 的位上，
MATT|23|3|所以凡他們所吩咐你們的，你們都要謹守遵行。但不要效法他們的行為，因為他們能說不能行。
MATT|23|4|他們把難挑的 重擔捆起來，擱在人的肩上，但自己一個指頭也不肯動。
MATT|23|5|他們所做的一切事都是要讓人看見，所以把佩戴的經匣 加寬了，衣裳的繸子加長了，
MATT|23|6|喜愛宴席上的首座、會堂裏的高位，
MATT|23|7|又喜歡人們在街市上向他們問安，稱呼他們拉比 。
MATT|23|8|但你們不要接受拉比的稱呼，因為只有一位是你們的老師；你們都是弟兄。
MATT|23|9|也不要稱呼地上的人為父，因為只有一位是你們的父，就是在天上的父。
MATT|23|10|不要接受師傅的稱呼，因為只有一位是你們的師傅，就是基督。
MATT|23|11|你們中間誰為大，誰就要作你們的用人。
MATT|23|12|凡自高的，必降為卑；自甘卑微的，必升為高。
MATT|23|13|「你們這假冒為善的文士和法利賽人有禍了！因為你們當著人的面把天國的門關了，自己不進去，要進去的人，你們也不容他們進去。
MATT|23|14|
MATT|23|15|「你們這假冒為善的文士和法利賽人有禍了！因為你們走遍海洋陸地，說服一個人入教，既入了教，卻使他成為比你們加倍壞的地獄之子。
MATT|23|16|「你們這瞎眼的嚮導有禍了！你們說：『凡指著聖所起誓的算不得甚麼；但是凡指著聖所中的金子起誓的，他就該謹守。』
MATT|23|17|你們這無知的瞎子啊，哪個更大呢？是金子，還是使金子成聖的聖所呢？
MATT|23|18|你們又說：『凡指著祭壇起誓的算不得甚麼；但是凡指著壇上祭物起誓的，他就該謹守。』
MATT|23|19|你們這些瞎子啊，哪個更大呢？是祭物，還是使祭物成聖的壇呢？
MATT|23|20|所以，人指著祭壇起誓，就是指著壇和壇上一切所有的起誓；
MATT|23|21|人指著聖所起誓，就是指著聖所和那住在聖所裏的起誓；
MATT|23|22|人指著天起誓，就是指著上帝的寶座和那坐在上面的起誓。
MATT|23|23|「你們這假冒為善的文士和法利賽人有禍了！因為你們將薄荷、大茴香、小茴香獻上十分之一，那律法上更重要的事，就是公義、憐憫、信實，你們反倒不做；這原是你們該做的－至於那些奉獻也不可廢棄。
MATT|23|24|你們這瞎眼的嚮導，蠓蟲你們就濾出來，駱駝你們倒吞下去。
MATT|23|25|「你們這假冒為善的文士和法利賽人有禍了！因為你們洗淨杯盤的外面，裏面卻滿了貪婪和放蕩。
MATT|23|26|你這瞎眼的法利賽人，先洗淨杯子 的裏面，好使外面也乾淨了。
MATT|23|27|「你們這假冒為善的文士和法利賽人有禍了！因為你們好像粉飾了的墳墓，外面好看，裏面卻滿了死人的骨頭和一切的污穢。
MATT|23|28|你們也是如此，外面對人顯出公義，裏面卻滿了虛偽和不法的事。
MATT|23|29|「你們這假冒為善的文士和法利賽人有禍了！因為你們建造先知的墳，裝修義人的墓，
MATT|23|30|說：『若是我們在先祖的時代，必不和他們一同流先知的血。』
MATT|23|31|這樣，你們就證明自己是殺害先知的人的子孫了。
MATT|23|32|你們去充滿你們祖宗的惡貫吧！
MATT|23|33|你們這些蛇啊，毒蛇的孽種啊，怎能逃脫地獄的懲罰呢？
MATT|23|34|所以，我差遣先知、智慧人和文士到你們這裏來，有的你們要殺害，要釘十字架；有的你們要在會堂裏鞭打，從這城追逼到那城，
MATT|23|35|如此，地上所有義人流的血都歸到你們身上，從義人 亞伯 的血起，直到你們在聖所和祭壇中間所殺的 巴拉加 的兒子 撒迦利亞 的血為止。
MATT|23|36|我實在告訴你們，這一切的罪都要歸到這世代了。」
MATT|23|37|「 耶路撒冷 啊， 耶路撒冷 啊，你常殺害先知，又用石頭打死那奉差遣到你這裏來的人。我多少次想聚集你的兒女，好像母雞把小雞聚集在翅膀底下，但是你們不願意。
MATT|23|38|看吧，你們的家要被廢棄成為荒蕪。
MATT|23|39|我告訴你們，從今以後，你們絕不會再見到我，直到你們說：『奉主名來的是應當稱頌的！』」
MATT|24|1|耶穌出了聖殿，正離開的時候，門徒前來，把聖殿的建築指給他看。
MATT|24|2|耶穌回應他們說：「你們不是看見這一切嗎？我實在告訴你們，這裏將沒有一塊石頭會留在另一塊石頭上，而不被拆毀的。」
MATT|24|3|耶穌在 橄欖山 上坐著，門徒私下進前來問他：「請告訴我們，甚麼時候有這些事呢？你來臨和世代的終結有甚麼預兆呢？」
MATT|24|4|耶穌回答他們：「你們要謹慎，免得有人迷惑你們。
MATT|24|5|因為將有好些人冒我的名來，說『我是基督』，並且要迷惑許多人。
MATT|24|6|你們也將聽見打仗和打仗的風聲。注意，不要驚慌！因為這些事必須發生，但這還不是終結。
MATT|24|7|民要攻打民，國要攻打國，多處必有饑荒、地震。
MATT|24|8|這都是災難 的起頭。
MATT|24|9|那時，人要使你們陷在患難裏，也要殺害你們；你們又要為我的名被萬民憎恨。
MATT|24|10|那時，會有許多人跌倒，也會彼此陷害，彼此憎恨；
MATT|24|11|且有好些假先知起來，迷惑許多人。
MATT|24|12|因為不法的事增多，許多人的愛心漸漸冷淡了。
MATT|24|13|但堅忍到底的終必得救。
MATT|24|14|這天國的福音要傳遍天下，對萬民作見證，然後終結才來到。」
MATT|24|15|「當你們看見先知 但以理 所說的那『施行毀滅的褻瀆者』站在聖地（讀這經的人要會意），
MATT|24|16|那時，在 猶太 的，應當逃到山上；
MATT|24|17|在屋頂上的，不要下來拿家裏的東西；
MATT|24|18|在田裏的，不要回去取衣裳。
MATT|24|19|在那些日子，懷孕的和奶孩子的就苦了。
MATT|24|20|你們要祈求，好讓你們逃走的時候，不遇見冬天或安息日。
MATT|24|21|因為那時必有大災難，自從世界的起頭直到如今，從沒有這樣的災難，將來也不會有。
MATT|24|22|若不減少那些日子，凡血肉之軀的，就沒有一個能得救；可是為了選民，那些日子將減少。
MATT|24|23|那時，若有人對你們說：『看哪，基督在這裏！』或『在那裏！』你們不要信。
MATT|24|24|因為假基督和假先知將要起來，顯大神蹟、大奇事，如果可能，要把選民也迷惑了。
MATT|24|25|看哪，我已經預先告訴你們了。
MATT|24|26|若有人對你們說：『看哪，基督在曠野裏！』你們不要出去；或說：『看哪，基督在內室中！』你們不要信。
MATT|24|27|好像閃電從東邊發出，直照到西邊，人子來臨也要這樣。
MATT|24|28|屍首在哪裏，鷹也會聚在哪裏。」
MATT|24|29|「那些日子的災難一過去， 太陽要變黑， 月亮也不放光， 眾星要從天上墜落， 天上的萬象都要震動。
MATT|24|30|那時，人子的預兆要顯在天上，地上的萬族都要哀哭。他們要看見人子帶著能力和大榮耀，駕著天上的雲來臨。
MATT|24|31|他要差遣天使，用大聲的號筒，從四方，從天這邊直到天那邊，召集他的選民。」
MATT|24|32|「你們要從無花果樹學習功課：當樹枝發芽長葉的時候，你們就知道夏天近了。
MATT|24|33|同樣，當你們看見這一切，就知道那時候近了，就在門口了。
MATT|24|34|我實在告訴你們，這世代還沒有過去，這一切都要發生。
MATT|24|35|天地要廢去，我的話卻絕不廢去。」
MATT|24|36|「但那日子，那時辰，沒有人知道，連天上的天使也不知道，子也不知道，惟有父知道。
MATT|24|37|挪亞 的日子怎樣，人子來臨也要怎樣。
MATT|24|38|在洪水以前的那些日子，人照常吃喝嫁娶，直到 挪亞 進方舟的那日，
MATT|24|39|不知不覺洪水來了，把他們全都沖去。人子來臨也要這樣。
MATT|24|40|那時，兩個人在田裏，一個被接去，一個被撇下。
MATT|24|41|兩個女人推磨，一個被接去，一個被撇下。
MATT|24|42|所以，你們要警醒，因為不知道你們的主哪一天來到。
MATT|24|43|你們要知道，一家的主人若知道晚上甚麼時候有賊來，就必警醒，不讓賊挖穿房屋。
MATT|24|44|所以，你們也要預備，因為在你們想不到的時候，人子就來了。」
MATT|24|45|「那麼，誰是那忠心又精明的僕人，主人派他管理自己的家僕、按時分糧給他們的呢？
MATT|24|46|主人來到，看見僕人這樣做，那僕人就有福了。
MATT|24|47|我實在告訴你們，主人要派他管理所有的財產。
MATT|24|48|如果那惡僕心裏說：『我的主人會來得遲』，
MATT|24|49|就動手打他的同伴，又和醉酒的人一同吃喝，
MATT|24|50|在想不到的日子，不知道的時候，那僕人的主人要來，
MATT|24|51|重重地懲罰他 ，定他和假冒為善的人同罪，在那裏他要哀哭切齒了。」
MATT|25|1|「那時，天國好比十個童女拿著燈出去迎接新郎。
MATT|25|2|其中有五個是愚拙的，五個是聰明的。
MATT|25|3|愚拙的拿著燈，卻沒有帶油；
MATT|25|4|聰明的拿著燈，又盛了油在器皿裏。
MATT|25|5|新郎遲延的時候，她們都打盹，睡著了。
MATT|25|6|半夜有人喊：『看，新郎來了，你們出來迎接他。』
MATT|25|7|那些童女就都起來挑亮她們的燈。
MATT|25|8|愚拙的對聰明的說：『請分點油給我們，因為我們的燈要滅了。』
MATT|25|9|聰明的回答：『恐怕不夠你我用的；你們還是自己到賣油的那裏去買吧。』
MATT|25|10|她們去買的時候，新郎到了。那預備好了的，與他進去共赴婚宴，門就關了。
MATT|25|11|其餘的童女隨後也來了，說：『主啊，主啊，給我們開門！』
MATT|25|12|他卻回答：『我實在告訴你們，我不認識你們。』
MATT|25|13|所以，你們要警醒，因為那日子，那時辰，你們不知道。」
MATT|25|14|「天國又好比一個人要出外遠行，就叫了僕人來，把他的家業交給他們。
MATT|25|15|他按著各人的才幹，給他們銀子：一個給了五千 ，一個給了二千 ，一個給了一千 ，就出外遠行去了。
MATT|25|16|那領五千的立刻拿去做買賣，另外賺了五千。
MATT|25|17|那領二千的也照樣另賺了二千。
MATT|25|18|但那領一千的去掘開地，把主人的銀子埋藏了。
MATT|25|19|過了許久，那些僕人的主人來了，和他們算賬。
MATT|25|20|那領五千的又帶著另外的五千來，說：『主啊，你交給我五千。請看，我又賺了五千。』
MATT|25|21|主人說：『好，你這又善良又忠心的僕人，你在少許的事上忠心，我要派你管理許多的事，進來享受你主人的快樂吧！』
MATT|25|22|那領二千的也進前來，說：『主啊，你交給我二千。請看，我又賺了二千。』
MATT|25|23|主人說：『好，你這又善良又忠心的僕人，你在少許的事上忠心，我要派你管理許多的事，進來享受你主人的快樂吧！』
MATT|25|24|那領一千的也進前來，說：『主啊，我知道你，你是個嚴厲的人：沒有種的地方也要收割，沒有播的地方也要收穫，
MATT|25|25|我就害怕，去把你的一千銀子埋藏在地裏。請看，你的銀子在這裏。』
MATT|25|26|他的主人回答他說：『你這又惡又懶的僕人，你既知道我沒有種的地方也要收割，沒有播的地方也要收穫，
MATT|25|27|就該把我的銀子放給兌換銀錢的人，到我來的時候可以連本帶利收回。
MATT|25|28|把他這一千奪過來，給那有一萬 的。
MATT|25|29|因為凡有的，還要加給他，叫他有餘；沒有的，連他所有的也要奪過來。
MATT|25|30|把這無用的僕人丟在外面黑暗裏，在那裏他要哀哭切齒了。』」
MATT|25|31|「當人子在他榮耀裏，同著眾天使來臨的時候，要坐在他榮耀的寶座上。
MATT|25|32|萬民都要聚集在他面前。他要把他們分別出來，好像牧人分別綿羊、山羊一般，
MATT|25|33|把綿羊安置在右邊，山羊在左邊。
MATT|25|34|於是王要向他右邊的說：『你們這蒙我父賜福的，可來承受那創世以來為你們所預備的國。
MATT|25|35|因為我餓了，你們給我吃；渴了，你們給我喝；我流浪在外，你們留我住；
MATT|25|36|我赤身露體，你們給我穿；我病了，你們看顧我；我在監獄裏，你們來看我。』
MATT|25|37|義人就回答：『主啊，我們甚麼時候見你餓了，給你吃；渴了，給你喝？
MATT|25|38|甚麼時候見你流浪在外，留你住；或是赤身露體，給你穿？
MATT|25|39|又甚麼時候見你病了，或是在監獄裏，來看你呢？』
MATT|25|40|王回答他們說：『我實在告訴你們，這些事你們做在我弟兄中一個最小的身上，就是做在我身上了。』
MATT|25|41|「王又要向那左邊的說：『你們這被詛咒的人，離開我！進入那為魔鬼和他的使者所預備的永火裏去！
MATT|25|42|因為我餓了，你們沒有給我吃；渴了，你們沒有給我喝；
MATT|25|43|我流浪在外，你們沒有留我住；我赤身露體，你們沒有給我穿；我病了，我在監獄裏，你們沒有來看顧我。』
MATT|25|44|他們也要回答：『主啊，我們甚麼時候見你餓了，或渴了，或流浪在外，或赤身露體，或病了，或在監獄裏，沒有伺候你呢？』
MATT|25|45|王要回答：『我實在告訴你們，這些事你們沒有做在任何一個最小的弟兄身上，就是沒有做在我身上了。』
MATT|25|46|這些人要往永刑裏去；那些義人要往永生裏去。」
MATT|26|1|耶穌說完了這一切的話，就對門徒說：
MATT|26|2|「你們知道，過兩天是逾越節，人子將要被出賣，釘在十字架上。」
MATT|26|3|那時，祭司長和百姓的長老聚集在那稱為 該亞法 的大祭司的院裏。
MATT|26|4|大家商議要設計捉拿耶穌，把他殺掉。
MATT|26|5|可是他們說：「不可在過節的日子，恐怕百姓生亂。」
MATT|26|6|耶穌在 伯大尼 的痲瘋病人 西門 家裏，
MATT|26|7|有一個女人拿著一玉瓶極貴的香膏來，趁耶穌坐席的時候，澆在他的頭上。
MATT|26|8|門徒看見就很不高興，說：「何必這樣浪費呢！
MATT|26|9|這香膏可以賣許多錢，賙濟窮人。」
MATT|26|10|耶穌看出他們的意思，就說：「為甚麼難為這女人呢？她在我身上做的是一件美事。
MATT|26|11|因為常有窮人和你們在一起，但是你們不常有我。
MATT|26|12|她把這香膏澆在我身上是為我安葬作準備的。
MATT|26|13|我實在告訴你們，普天之下，無論在甚麼地方傳這福音，都要述說這女人所做的，來記念她。」
MATT|26|14|當時，十二使徒中有一個叫 加略 人 猶大 的，去見祭司長，
MATT|26|15|說：「我把他交給你們，你們願意給我多少錢？」他們給了他三十塊銀錢。
MATT|26|16|從那時候起，他就找機會要把耶穌交給他們。
MATT|26|17|除酵節的第一天，門徒來問耶穌：「你要我們在哪裏給你預備吃逾越節的宴席呢？」
MATT|26|18|耶穌說：「你們進城去，到某人那裏，對他說：『老師說：我的時候快到了，我要和我的門徒在你家裏守逾越節。』」
MATT|26|19|門徒遵照耶穌所吩咐的去預備了逾越節的宴席。
MATT|26|20|到了晚上，耶穌和十二使徒坐席。
MATT|26|21|他們吃的時候，耶穌說：「我實在告訴你們，你們中間有一個人要出賣我。」
MATT|26|22|他們就非常憂愁，一個一個地問他：「主，該不是我吧？」
MATT|26|23|耶穌回答說：「同我蘸手在盤子裏的，就是要出賣我的。
MATT|26|24|人子要去了，正如經上所寫有關他的；但出賣人子的人有禍了！那人沒有出生倒好。」
MATT|26|25|出賣耶穌的 猶大 回答他說：「拉比，該不是我吧？」耶穌說：「你自己說了。」
MATT|26|26|他們吃的時候，耶穌拿起餅來，祝福了，就擘開，遞給門徒，說：「你們拿去，吃吧。這是我的身體。」
MATT|26|27|他又拿起杯來，祝謝了，遞給他們，說：「你們都喝這個，
MATT|26|28|因為這是我立約的血，為許多人流出來，使罪得赦。
MATT|26|29|但我告訴你們，從今以後，我不再喝這葡萄汁，直到我在我父的國裏與你們同喝新的那日子。」
MATT|26|30|他們唱了詩，就出來往 橄欖山 去。
MATT|26|31|那時，耶穌對他們說：「今夜，你們為我的緣故都要跌倒。因為經上記著： 『我要擊打牧人， 羊就分散了。』
MATT|26|32|但我復活以後，要在你們之前往 加利利 去。」
MATT|26|33|彼得 回答他說：「即使眾人為你的緣故跌倒，我也絕不跌倒。」
MATT|26|34|耶穌說：「我實在告訴你，今夜雞叫以前，你要三次不認我。」
MATT|26|35|彼得 說：「我就是必須和你同死，也絕不會不認你。」所有的門徒都是這樣說。
MATT|26|36|耶穌和門徒來到一個地方，名叫 客西馬尼 。他對他們說：「你們坐在這裏，我到那邊去禱告。」
MATT|26|37|於是他帶著 彼得 和 西庇太 的兩個兒子同去。他憂愁起來，極其難過，
MATT|26|38|就對他們說：「我心裏非常憂傷，幾乎要死；你們留在這裏，和我一同警醒。」
MATT|26|39|他就稍往前走，俯伏在地，禱告說：「我父啊，如果可能，求你使這杯離開我。然而，不是照我所願的，而是照你所願的。」
MATT|26|40|他回到門徒那裏，見他們睡著了，就對 彼得 說：「怎麼樣？你們不能同我警醒一小時嗎？
MATT|26|41|總要警醒禱告，免得陷入試探。你們心靈固然願意，肉體卻軟弱了。」
MATT|26|42|他第二次又去禱告說：「我父啊，這杯若不能離開我，必須我喝，就願你的旨意成全。」
MATT|26|43|他又來，見他們睡著了，因為他們的眼睛困倦。
MATT|26|44|耶穌又離開他們，第三次去禱告，說的話跟先前一樣。
MATT|26|45|然後他來到門徒那裏，對他們說：「現在你們仍在睡覺安歇嗎？看哪，時候到了，人子被出賣在罪人手裏了。
MATT|26|46|起來，我們走吧！看哪，那出賣我的人快來了。」
MATT|26|47|耶穌還在說話的時候，十二使徒之一的 猶大 來了，還有一大群人帶著刀棒，從祭司長和百姓的長老那裏跟他同來。
MATT|26|48|那出賣耶穌的給了他們一個暗號，說：「我親誰，誰就是。你們把他抓住。」
MATT|26|49|猶大 立刻進前來對耶穌說：「拉比，你好！」就跟他親吻。
MATT|26|50|耶穌對他說：「朋友，你來要做的事，就做吧。 」於是那些人上前，下手抓住耶穌。
MATT|26|51|忽然，有一個和耶穌一起的人伸手拔出刀來，把大祭司的僕人砍了一刀，削掉了他一隻耳朵。
MATT|26|52|耶穌對他說：「收刀入鞘吧！凡動刀的，必死在刀下。
MATT|26|53|你想我不能求我父，現在為我差遣比十二營還多的天使來嗎？
MATT|26|54|若是這樣，經上所說事情必須如此發生的話怎麼應驗呢？」
MATT|26|55|就在那時，耶穌對眾人說：「你們帶著刀棒出來抓我，如同拿強盜嗎？我天天坐在聖殿裏教導人，你們並沒有抓我。
MATT|26|56|但這整件事的發生，是要應驗先知書上的話。」那時，門徒都離開他，逃走了。
MATT|26|57|抓耶穌的人把他帶到大祭司 該亞法 那裏去，文士和長老已經在那裏聚集。
MATT|26|58|彼得 遠遠地跟著耶穌，直到大祭司的院子，進到裏面，就和警衛同坐，要看結局怎樣。
MATT|26|59|祭司長和全議會尋找假見證控告耶穌，要處死他。
MATT|26|60|雖然有好些人來作假見證，總找不到實據。最後有兩個人前來，
MATT|26|61|說：「這個人曾說：『我能拆毀上帝的殿，三日內又建造起來。』」
MATT|26|62|大祭司就站起來，對耶穌說：「這些人作證告你的事，你甚麼都不回答嗎？」
MATT|26|63|耶穌卻不言語。大祭司對他說：「我指著永生上帝命令你起誓告訴我們，你是不是基督—上帝的兒子？」
MATT|26|64|耶穌對他說：「你自己說了。然而，我告訴你們， 此後你們要看見人子 坐在權能者的右邊， 駕著天上的雲來臨。」
MATT|26|65|大祭司就撕裂衣服，說：「他說了褻瀆的話，我們何必再要證人呢？現在你們已經聽見他這褻瀆的話了。
MATT|26|66|你們的意見如何？」他們回答：「他該處死。」
MATT|26|67|他們就吐唾沫在他臉上，用拳頭打他，也有打他耳光的，
MATT|26|68|說：「基督啊，向我們說預言吧！打你的是誰？」
MATT|26|69|彼得 在外面院子裏坐著，有一個使女進前來，說：「你素來也是同那 加利利 人耶穌一起的。」
MATT|26|70|彼得 在眾人面前卻不承認，說：「我不知道你說的是甚麼！」
MATT|26|71|他出去，到了門口，又有一個使女看見他，就對那裏的人說：「這個人是同 拿撒勒 人耶穌一起的。」
MATT|26|72|彼得 又不承認，起誓說：「我不認得那個人。」
MATT|26|73|過了不久，旁邊站著的人前來，對 彼得 說：「你的確是他們一夥的，你的口音把你顯露出來了。」
MATT|26|74|彼得 就賭咒發誓說：「我不認得那個人。」立刻雞就叫了。
MATT|26|75|彼得 想起耶穌所說的話：「雞叫以前，你要三次不認我。」他就出去痛哭。
MATT|27|1|到了早晨，眾祭司長和百姓的長老商議要處死耶穌，
MATT|27|2|就把他綁著，解去，交給 彼拉多 總督。
MATT|27|3|這時，出賣耶穌的 猶大 看見耶穌已經定了罪，就後悔，把那三十塊銀錢拿回來給祭司長和長老，
MATT|27|4|說：「我出賣了無辜人的血有罪了。」他們說：「那跟我們有甚麼相干？你自己承當吧！」
MATT|27|5|猶大 就把那銀錢丟在殿裏，出去吊死了。
MATT|27|6|祭司長拾起銀錢來，說：「這是血價，不可放在聖殿的銀庫裏。」
MATT|27|7|他們商議，就用那銀錢買了窯戶的一塊田，用來埋葬外鄉人。
MATT|27|8|所以，那塊田直到今日還叫做「血田」。
MATT|27|9|這就應驗了先知 耶利米 所說的話：「他們用那三十塊銀錢，就是 以色列 人給那被估定的人所估定的價錢，
MATT|27|10|買了窯戶的一塊田；這是照著主所吩咐我的。」
MATT|27|11|耶穌站在總督面前，總督問他：「你是 猶太 人的王嗎？」耶穌說：「是你說的。」
MATT|27|12|他被祭司長和長老控告的時候，甚麼都不回答。
MATT|27|13|彼拉多 就對他說：「他們作證告你這麼多的事，你沒有聽見嗎？」
MATT|27|14|耶穌仍不回答，連一句話也不說，以致總督覺得非常驚訝。
MATT|27|15|總督有一個常例，每逢這節期，隨眾人的意願釋放一個囚犯給他們。
MATT|27|16|當時有一個出名的囚犯叫 巴拉巴 。
MATT|27|17|眾人聚集的時候， 彼拉多 就對他們說：「你們要我釋放哪一個給你們？是 巴拉巴 呢？是稱為基督的耶穌呢？」
MATT|27|18|總督原知道他們是因為嫉妒才把他解了來。
MATT|27|19|正坐堂的時候，他的夫人打發人來說：「這義人的事，你一點不可管，因為我今天在夢中因他受了許多的苦。」
MATT|27|20|祭司長和長老挑唆眾人，要求釋放 巴拉巴 ，除掉耶穌。
MATT|27|21|總督回答他們說：「這兩個人，你們要我釋放哪一個給你們呢？」他們說：「 巴拉巴 。」
MATT|27|22|彼拉多 說：「這樣，那稱為基督的耶穌我怎麼辦他呢？」他們都說：「把他釘十字架！」
MATT|27|23|總督說：「為甚麼？他做了甚麼惡事呢？」他們更加喊著說：「把他釘十字架！」
MATT|27|24|彼拉多 見說也無濟於事，反要生亂，就拿水在眾人面前洗手，說：「流這人 的血，罪不在我，你們承當吧。」
MATT|27|25|眾人都回答：「他的血歸到我們和我們的子孫身上！」
MATT|27|26|於是 彼拉多 釋放 巴拉巴 給他們，把耶穌鞭打後交給人釘十字架。
MATT|27|27|總督的兵把耶穌帶進總督府，把全營的兵都聚集在耶穌那裏。
MATT|27|28|他們脫了他的衣服，穿上一件朱紅色的袍子，
MATT|27|29|用荊棘編了冠冕，戴在他頭上，拿一根蘆葦稈放在他右手裏，跪在他面前，戲弄他，說：「萬歲， 猶太 人的王！」
MATT|27|30|他們又向他吐唾沫，拿蘆葦稈打他的頭。
MATT|27|31|他們戲弄完了，就給他脫了袍子，又穿上他自己的衣服，帶他出去，要釘十字架。
MATT|27|32|他們出去的時候，遇見一個 古利奈 人，名叫 西門 ，就強迫他同去，好背耶穌的十字架。
MATT|27|33|他們到了一個地方，名叫 各各他 ，就是「髑髏地」。
MATT|27|34|士兵拿苦膽調和的酒給耶穌喝。他嘗了，不肯喝。
MATT|27|35|他們把他釘在十字架上，然後抽籤分了他的衣服，
MATT|27|36|又坐在那裏看守他。
MATT|27|37|他們在他頭上方安了一個罪狀牌，寫著：「這是 猶太 人的王耶穌。」
MATT|27|38|當時，有兩個強盜和他同釘十字架，一個在右邊，一個在左邊。
MATT|27|39|從那裏經過的人譏笑他，搖著頭，
MATT|27|40|說：「你這拆毀殿、三日又建造起來的，救救你自己吧！如果你是上帝的兒子，就從十字架上下來呀！」
MATT|27|41|眾祭司長、文士和長老也同樣嘲笑他，說：
MATT|27|42|「他救了別人，不能救自己。他是 以色列 的王，現在從十字架上下來，我們就信他。
MATT|27|43|他倚靠上帝，上帝若願意，現在就來救他，因為他曾說『我是上帝的兒子』。」
MATT|27|44|和他同釘的強盜也這樣譏諷他。
MATT|27|45|從正午到下午三點鐘，遍地都黑暗了。
MATT|27|46|約在下午三點鐘，耶穌大聲高呼，說：「以利！以利！拉馬撒巴各大尼？」就是說：「我的上帝！我的上帝！為甚麼離棄我？」
MATT|27|47|站在那裏的人，有的聽見就說：「這個人呼叫 以利亞 呢！」
MATT|27|48|其中有一個人立刻跑去，拿海綿蘸滿了醋，綁在蘆葦稈上，送給他喝。
MATT|27|49|其餘的人說：「且等著，看 以利亞 來不來救他。」
MATT|27|50|耶穌又大喊一聲，氣就斷了。
MATT|27|51|忽然，殿的幔子從上到下裂為兩半，地震動，磐石崩裂，
MATT|27|52|墳墓也開了，有許多已睡了的聖徒的身體也復活了。
MATT|27|53|耶穌復活以後，他們從墳墓裏出來，進了聖城，向許多人顯現。
MATT|27|54|百夫長和跟他一同看守耶穌的人看見地震和所經歷的事，非常害怕，說：「他真是上帝的兒子！」
MATT|27|55|有好些婦女在那裏，遠遠地觀看，她們是從 加利利 跟隨耶穌，來服事他的；
MATT|27|56|其中有 抹大拉 的 馬利亞 ，又有 雅各 和 約瑟 的母親 馬利亞 ，並有 西庇太 兩個兒子的母親。
MATT|27|57|到了晚上，有一個財主，名叫 約瑟 ，是 亞利馬太 來的，他也是耶穌的門徒。
MATT|27|58|這人去見 彼拉多 ，請求要耶穌的身體， 彼拉多 就吩咐給他。
MATT|27|59|約瑟 取了身體，用乾淨的細麻布裹好，
MATT|27|60|然後把他安放在自己的新墓穴裏，就是他鑿在巖石裏的。他又把大石頭滾到墓門口，然後離開。
MATT|27|61|有 抹大拉 的 馬利亞 和另一個 馬利亞 在那裏，對著墳墓坐著。
MATT|27|62|次日，就是預備日的第二天，祭司長和法利賽人聚集來見 彼拉多 ，
MATT|27|63|說：「大人，我們記得那迷惑人的還活著的時候曾說：『三天後我要復活。』
MATT|27|64|因此，請吩咐人將墳墓把守妥當，直到第三天，恐怕他的門徒來把他偷了去，就告訴百姓說：『他從死人中復活了。』這樣的話，那後來的迷惑就比先前的更厲害了。」
MATT|27|65|彼拉多 說：「你們有看守的兵，去吧！盡你們所能的把守妥當。」
MATT|27|66|他們就帶著看守的兵同去，封了石頭，將墳墓把守妥當。
MATT|28|1|安息日過後，七日的第一日，天快亮的時候， 抹大拉 的 馬利亞 和另一個 馬利亞 來看墳墓。
MATT|28|2|忽然，地大震動；因為有主的一個使者從天上下來，把石頭滾開，坐在上面。
MATT|28|3|他的相貌如同閃電，衣服潔白如雪。
MATT|28|4|看守的人嚇得渾身顫抖，甚至和死人一樣。
MATT|28|5|天使回應婦女說：「不要害怕！我知道你們是尋找那釘十字架的耶穌。
MATT|28|6|他不在這裏，照他所說的，他已經復活了。你們來！看看安放他的地方。
MATT|28|7|快去告訴他的門徒，說他已從死人中復活了，並且要比你們先到 加利利 去，在那裏你們會看見他。看哪！我已經告訴你們了。」
MATT|28|8|婦女們急忙離開墳墓，又害怕，又大為歡喜，跑去告訴他的門徒。
MATT|28|9|忽然，耶穌迎上她們，說：「平安！」她們就上前抱住他的腳拜他。
MATT|28|10|耶穌對她們說：「不要害怕！你們去告訴我的弟兄，叫他們往 加利利 去，在那裏會見到我。」
MATT|28|11|她們去的時候，看守的兵有幾個進城去，把所發生的事都報告祭司長。
MATT|28|12|祭司長和長老聚集商議，就拿許多銀錢給士兵，
MATT|28|13|說：「你們要這樣說：『夜間我們睡覺的時候，他的門徒來把他偷去了。』
MATT|28|14|若是這話被總督聽見，有我們勸他，保你們無事。」
MATT|28|15|士兵收了銀錢，就照所囑咐他們的去做。這話就在 猶太 人中間流傳，直到今日。
MATT|28|16|十一個門徒往 加利利 去，到了耶穌指定他們去的山上。
MATT|28|17|他們見了耶穌就拜他，然而還有人疑惑。
MATT|28|18|耶穌進前來，對他們說：「天上地下所有的權柄都賜給我了。
MATT|28|19|所以，你們要去，使萬民作我的門徒，奉父、子、聖靈的名給他們施洗 ，
MATT|28|20|凡我所吩咐你們的，都教導他們遵守。看哪，我天天與你們同在，直到世代的終結。」
