ZECH|1|1|В восьмом месяце, во второй год Дария, было слово Господне к Захарии, сыну Варахиину, сыну Аддову, пророку:
ZECH|1|2|прогневался Господь на отцов ваших великим гневом,
ZECH|1|3|и ты скажи им: так говорит Господь Саваоф: обратитесь ко Мне, говорит Господь Саваоф, и Я обращусь к вам, говорит Господь Саваоф.
ZECH|1|4|Не будьте такими, как отцы ваши, к которым взывали прежде бывшие пророки, говоря: "так говорит Господь Саваоф: обратитесь от злых путей ваших и от злых дел ваших"; но они не слушались и не внимали Мне, говорит Господь.
ZECH|1|5|Отцы ваши – где они? да и пророки, будут ли они вечно жить?
ZECH|1|6|Но слова Мои и определения Мои, которые заповедал Я рабам Моим, пророкам, разве не постигли отцов ваших? и они обращались и говорили: "как определил Господь Саваоф поступить с нами по нашим путям и по нашим делам, так и поступил с нами".
ZECH|1|7|В двадцать четвертый день одиннадцатого месяца, – это месяц Шеват, – во второй год Дария, было слово Господне к Захарии, сыну Варахиину, сыну Аддову, пророку:
ZECH|1|8|видел я ночью: вот, муж на рыжем коне стоит между миртами, которые в углублении, а позади него кони рыжие, пегие и белые, –
ZECH|1|9|и сказал я: кто они, господин мой? И сказал мне Ангел, говоривший со мною: я покажу тебе, кто они.
ZECH|1|10|И отвечал муж, который стоял между миртами, и сказал: это те, которых Господь послал обойти землю.
ZECH|1|11|И они отвечали Ангелу Господню, стоявшему между миртами, и сказали: обошли мы землю, и вот, вся земля населена и спокойна.
ZECH|1|12|И отвечал Ангел Господень и сказал: Господи Вседержителю! Доколе Ты не умилосердишься над Иерусалимом и над городами Иуды, на которые Ты гневаешься вот уже семьдесят лет?
ZECH|1|13|Тогда в ответ Ангелу, говорившему со мною, изрек Господь слова благие, слова утешительные.
ZECH|1|14|И сказал мне Ангел, говоривший со мною: провозгласи и скажи: так говорит Господь Саваоф: возревновал Я о Иерусалиме и о Сионе ревностью великою;
ZECH|1|15|и великим негодованием негодую на народы, живущие в покое; ибо, когда Я мало прогневался, они усилили зло.
ZECH|1|16|Посему так говорит Господь: Я обращаюсь к Иерусалиму с милосердием; в нем соорудится дом Мой, говорит Господь Саваоф, и землемерная вервь протянется по Иерусалиму.
ZECH|1|17|Еще провозгласи и скажи: так говорит Господь Саваоф: снова переполнятся города Мои добром, и утешит Господь Сион, и снова изберет Иерусалим.
ZECH|1|18|И поднял я глаза мои и увидел: вот четыре рога.
ZECH|1|19|И сказал я Ангелу, говорившему со мною: что это? И он ответил мне: это роги, которые разбросали Иуду, Израиля и Иерусалим.
ZECH|1|20|Потом показал мне Господь четырех рабочих.
ZECH|1|21|И сказал я: что они идут делать? Он сказал мне так: эти роги разбросали Иуду, так что никто не может поднять головы своей; а сии пришли устрашить их, сбить роги народов, поднявших рог свой против земли Иуды, чтобы рассеять ее.
ZECH|2|1|И снова я поднял глаза мои и увидел: вот муж, у которого в руке землемерная вервь.
ZECH|2|2|Я спросил: куда ты идешь? и он сказал мне: измерять Иерусалим, чтобы видеть, какая широта его и какая длина его.
ZECH|2|3|И вот Ангел, говоривший со мною, выходит, а другой Ангел идет навстречу ему,
ZECH|2|4|и сказал он этому: иди скорее, скажи этому юноше: Иерусалим заселит окрестности по причине множества людей и скота в нем.
ZECH|2|5|И Я буду для него, говорит Господь, огненною стеною вокруг него и прославлюсь посреди него.
ZECH|2|6|Эй, эй! бегите из северной страны, говорит Господь: ибо по четырем ветрам небесным Я рассеял вас, говорит Господь.
ZECH|2|7|Спасайся, Сион, обитающий у дочери Вавилона.
ZECH|2|8|Ибо так говорит Господь Саваоф: для славы Он послал Меня к народам, грабившим вас, ибо касающийся вас касается зеницы ока Его.
ZECH|2|9|И вот, Я подниму руку Мою на них, и они сделаются добычею рабов своих, и тогда узнаете, что Господь Саваоф послал Меня.
ZECH|2|10|Ликуй и веселись, дщерь Сиона! Ибо вот, Я приду и поселюсь посреди тебя, говорит Господь.
ZECH|2|11|И прибегнут к Господу многие народы в тот день, и будут Моим народом; и Я поселюсь посреди тебя, и узнаешь, что Господь Саваоф послал Меня к тебе.
ZECH|2|12|Тогда Господь возьмет во владение Иуду, Свой удел на святой земле, и снова изберет Иерусалим.
ZECH|2|13|Да молчит всякая плоть пред лицем Господа! Ибо Он поднимается от святаго жилища Своего.
ZECH|3|1|И показал он мне Иисуса, великого иерея, стоящего перед Ангелом Господним, и сатану, стоящего по правую руку его, чтобы противодействовать ему.
ZECH|3|2|И сказал Господь сатане: Господь да запретит тебе, сатана, да запретит тебе Господь, избравший Иерусалим! не головня ли он, исторгнутая из огня?
ZECH|3|3|Иисус же одет был в запятнанные одежды и стоял перед Ангелом,
ZECH|3|4|который отвечал и сказал стоявшим перед ним так: снимите с него запятнанные одежды. А ему самому сказал: смотри, Я снял с тебя вину твою и облекаю тебя в одежды торжественные.
ZECH|3|5|И сказал: возложите на голову его чистый кидар. И возложили чистый кидар на голову его и облекли его в одежду; Ангел же Господень стоял.
ZECH|3|6|И засвидетельствовал Ангел Господень и сказал Иисусу:
ZECH|3|7|так говорит Господь Саваоф: если ты будешь ходить по Моим путям и если будешь на страже Моей, то будешь судить дом Мой и наблюдать за дворами Моими. Я дам тебе ходить между сими, стоящими здесь.
ZECH|3|8|Выслушай же, Иисус, иерей великий, ты и собратия твои, сидящие перед тобою, мужи знаменательные: вот, Я привожу раба Моего, ОТРАСЛЬ.
ZECH|3|9|Ибо вот тот камень, который Я полагаю перед Иисусом; на этом одном камне семь очей; вот, Я вырежу на нем начертания его, говорит Господь Саваоф, и изглажу грех земли сей в один день.
ZECH|3|10|В тот день, говорит Господь Саваоф, будете друг друга приглашать под виноград и под смоковницу.
ZECH|4|1|И возвратился тот Ангел, который говорил со мною, и пробудил меня, как пробуждают человека от сна его.
ZECH|4|2|И сказал он мне: что ты видишь? И отвечал я: вижу, вот светильник весь из золота, и чашечка для елея наверху его, и семь лампад на нем, и по семи трубочек у лампад, которые наверху его;
ZECH|4|3|и две маслины на нем, одна с правой стороны чашечки, другая с левой стороны ее.
ZECH|4|4|И отвечал я и сказал Ангелу, говорившему со мною: что это, господин мой?
ZECH|4|5|И Ангел, говоривший со мною, отвечал и сказал мне: ты не знаешь, что это? И сказал я: не знаю, господин мой.
ZECH|4|6|Тогда отвечал он и сказал мне так: это слово Господа к Зоровавелю, выражающее: не воинством и не силою, но Духом Моим, говорит Господь Саваоф.
ZECH|4|7|Кто ты, великая гора, перед Зоровавелем? ты – равнина, и вынесет он краеугольный камень при шумных восклицаниях: "благодать, благодать на нем!"
ZECH|4|8|И было ко мне слово Господне:
ZECH|4|9|руки Зоровавеля положили основание дому сему; его руки и окончат его, и узнаешь, что Господь Саваоф послал Меня к вам.
ZECH|4|10|Ибо кто может считать день сей маловажным, когда радостно смотрят на строительный отвес в руках Зоровавеля те семь, – это очи Господа, которые объемлют взором всю землю?
ZECH|4|11|Тогда отвечал я и сказал ему: что значат те две маслины с правой стороны светильника и с левой стороны его?
ZECH|4|12|Вторично стал я говорить и сказал ему: что значат две масличные ветви, которые через две золотые трубочки изливают из себя золото?
ZECH|4|13|И сказал он мне: ты не знаешь, что это? Я отвечал: не знаю, господин мой.
ZECH|4|14|И сказал он: это два помазанные елеем, предстоящие Господу всей земли.
ZECH|5|1|И опять поднял я глаза мои и увидел: вот летит свиток.
ZECH|5|2|И сказал он мне: что видишь ты? Я отвечал: вижу летящий свиток; длина его двадцать локтей, а ширина его десять локтей.
ZECH|5|3|Он сказал мне: это проклятие, исходящее на лице всей земли; ибо всякий, кто крадет, будет истреблен, как написано на одной стороне, и всякий, клянущийся ложно, истреблен будет, как написано на другой стороне.
ZECH|5|4|Я навел его, говорит Господь Саваоф, и оно войдет в дом татя и в дом клянущегося Моим именем ложно, и пребудет в доме его, и истребит его, и дерева его, и камни его.
ZECH|5|5|И вышел Ангел, говоривший со мною, и сказал мне: подними еще глаза твои и посмотри, что это выходит?
ZECH|5|6|Когда же я сказал: что это? Он отвечал: это выходит ефа, и сказал: это образ их по всей земле.
ZECH|5|7|И вот, кусок свинца поднялся, и там сидела одна женщина посреди ефы.
ZECH|5|8|И сказал он: эта [женщина] – само нечестие, и бросил ее в средину ефы, а на отверстие ее бросил свинцовый кусок.
ZECH|5|9|И поднял я глаза мои и увидел: вот, появились две женщины, и ветер был в крыльях их, и крылья у них как крылья аиста; и подняли они ефу и понесли ее между землею и небом.
ZECH|5|10|И сказал я Ангелу, говорившему со мною: куда несут они эту ефу?
ZECH|5|11|Тогда сказал он мне: чтобы устроить для нее дом в земле Сеннаар, и когда будет все приготовлено, то она поставится там на своей основе.
ZECH|6|1|И опять поднял я глаза мои и вижу: вот, четыре колесницы выходят из ущелья между двумя горами; и горы те [были] горы медные.
ZECH|6|2|В первой колеснице кони рыжие, а во второй колеснице кони вороные;
ZECH|6|3|в третьей колеснице кони белые, а в четвертой колеснице кони пегие, сильные.
ZECH|6|4|И, начав речь, я сказал Ангелу, говорившему со мною: что это, господин мой?
ZECH|6|5|И отвечал Ангел и сказал мне: это выходят четыре духа небесных, которые предстоят пред Господом всей земли.
ZECH|6|6|Вороные кони там выходят к стране северной и белые идут за ними, а пегие идут к стране полуденной.
ZECH|6|7|И сильные вышли и стремились идти, чтобы пройти землю; и он сказал: идите, пройдите землю, – и они прошли землю.
ZECH|6|8|Тогда позвал он меня и сказал мне так: смотри, вышедшие в землю северную успокоили дух Мой на земле северной.
ZECH|6|9|И было слово Господне ко мне:
ZECH|6|10|возьми у пришедших из плена, у Хелдая, у Товии и у Иедая, и пойди в тот самый день, пойди в дом Иосии, сына Софониева, куда они пришли из Вавилона,
ZECH|6|11|возьми [у них] серебро и золото и сделай венцы, и возложи на голову Иисуса, сына Иоседекова, иерея великого,
ZECH|6|12|и скажи ему: так говорит Господь Саваоф: вот Муж, – имя Ему ОТРАСЛЬ, Он произрастет из Своего корня и создаст храм Господень.
ZECH|6|13|Он создаст храм Господень и примет славу, и воссядет, и будет владычествовать на престоле Своем; будет и священником на престоле Своем, и совет мира будет между тем и другим.
ZECH|6|14|А венцы те будут Хелему и Товии, Иедаю и Хену, сыну Софониеву, на память в храме Господнем.
ZECH|6|15|И издали придут, и примут участие в построении храма Господня, и вы узнаете, что Господь Саваоф послал меня к вам, и это будет, если вы усердно будете слушаться гласа Господа Бога вашего.
ZECH|7|1|В четвертый год царя Дария было слово Господне к Захарии, в четвертый день девятого месяца, Хаслева,
ZECH|7|2|когда Вефиль послал Сарецера и Регем–Мелеха и спутников его помолиться пред лицем Господа
ZECH|7|3|и спросить у священников, которые в доме Господа Саваофа, и у пророков, говоря: "плакать ли мне в пятый месяц и поститься, как я делал это уже много лет?"
ZECH|7|4|И было ко мне слово Господа Саваофа:
ZECH|7|5|скажи всему народу земли сей и священникам так: когда вы постились и плакали в пятом и седьмом месяце, притом уже семьдесят лет, для Меня ли вы постились? для Меня ли?
ZECH|7|6|И когда вы едите и когда пьете, не для себя ли вы едите, не для себя ли вы пьете?
ZECH|7|7|Не те же ли слова провозглашал Господь через прежних пророков, когда еще Иерусалим был населен и покоен, и города вокруг него, южная страна и низменность, были населены?
ZECH|7|8|И было слово Господне к Захарии:
ZECH|7|9|так говорил тогда Господь Саваоф: производите суд справедливый и оказывайте милость и сострадание каждый брату своему;
ZECH|7|10|вдовы и сироты, пришельца и бедного не притесняйте и зла друг против друга не мыслите в сердце вашем.
ZECH|7|11|Но они не хотели внимать, отворотились от Меня, и уши свои отяготили, чтобы не слышать.
ZECH|7|12|И сердце свое окаменили, чтобы не слышать закона и слов, которые посылал Господь Саваоф Духом Своим через прежних пророков; за то и постиг их великий гнев Господа Саваофа.
ZECH|7|13|И было: как Он взывал, а они не слушали, так и они взывали, а Я не слушал, говорит Господь Саваоф.
ZECH|7|14|И Я развеял их по всем народам, которых они не знали, и земля сия опустела после них, так что никто не ходил по ней ни взад, ни вперед, и они сделали вожделенную страну пустынею.
ZECH|8|1|И было слово Господа Саваофа:
ZECH|8|2|так говорит Господь Саваоф: возревновал Я о Сионе ревностью великою, и с великим гневом возревновал Я о нем.
ZECH|8|3|Так говорит Господь: обращусь Я к Сиону и буду жить в Иерусалиме, и будет называться Иерусалим городом истины, и гора Господа Саваофа – горою святыни.
ZECH|8|4|Так говорит Господь Саваоф: опять старцы и старицы будут сидеть на улицах в Иерусалиме, каждый с посохом в руке, от множества дней.
ZECH|8|5|И улицы города сего наполнятся отроками и отроковицами, играющими на улицах его.
ZECH|8|6|Так говорит Господь Саваоф: если это в глазах оставшегося народа покажется дивным во дни сии, то неужели оно дивно и в Моих очах? говорит Господь Саваоф.
ZECH|8|7|Так говорит Господь Саваоф: вот, Я спасу народ Мой из страны востока и из страны захождения солнца;
ZECH|8|8|и приведу их, и будут они жить в Иерусалиме, и будут Моим народом, и Я буду их Богом, в истине и правде.
ZECH|8|9|Так говорит Господь Саваоф: укрепите руки ваши вы, слышащие ныне слова сии из уст пророков, бывших при основании дома Господа Саваофа, для создания храма.
ZECH|8|10|Ибо прежде дней тех не было возмездия для человека, ни возмездия за труд животных; ни уходящему, ни приходящему не было покоя от врага; и попускал Я всякого человека враждовать против другого.
ZECH|8|11|А ныне для остатка этого народа Я не такой, как в прежние дни, говорит Господь Саваоф.
ZECH|8|12|Ибо посев будет в мире; виноградная лоза даст плод свой, и земля даст произведения свои, и небеса будут давать росу свою, и все это Я отдам во владение оставшемуся народу сему.
ZECH|8|13|И будет: как вы, дом Иудин и дом Израилев, были проклятием у народов, так Я спасу вас, и вы будете благословением; не бойтесь; да укрепятся руки ваши!
ZECH|8|14|Ибо так говорит Господь Саваоф; как Я определил наказать вас, когда отцы ваши прогневали Меня, говорит Господь Саваоф, и не отменил,
ZECH|8|15|так опять Я определил в эти дни соделать доброе Иерусалиму и дому Иудину; не бойтесь!
ZECH|8|16|Вот дела, которые вы должны делать: говорите истину друг другу; по истине и миролюбно судите у ворот ваших.
ZECH|8|17|Никто из вас да не мыслит в сердце своем зла против ближнего своего, и ложной клятвы не любите, ибо все это Я ненавижу, говорит Господь.
ZECH|8|18|И было ко мне слово Господа Саваофа:
ZECH|8|19|так говорит Господь Саваоф: пост четвертого месяца и пост пятого, и пост седьмого, и пост десятого соделается для дома Иудина радостью и веселым торжеством; только любите истину и мир.
ZECH|8|20|Так говорит Господь Саваоф: еще будут приходить народы и жители многих городов;
ZECH|8|21|и пойдут жители одного города к жителям другого и скажут: пойдем молиться лицу Господа и взыщем Господа Саваофа; [и каждый] [скажет]: пойду и я.
ZECH|8|22|И будут приходить многие племена и сильные народы, чтобы взыскать Господа Саваофа в Иерусалиме и помолиться лицу Господа.
ZECH|8|23|Так говорит Господь Саваоф: будет в те дни, возьмутся десять человек из всех разноязычных народов, возьмутся за полу Иудея и будут говорить: мы пойдем с тобою, ибо мы слышали, что с вами Бог.
ZECH|9|1|Пророческое слово Господа на землю Хадрах, и на Дамаске оно остановится, – ибо око Господа на всех людей, как и на все колена Израилевы, –
ZECH|9|2|и на Емаф, смежный с ним, на Тир и Сидон, ибо он очень умудрился.
ZECH|9|3|И устроил себе Тир крепость, накопил серебра, как пыли, и золота, как уличной грязи.
ZECH|9|4|Вот, Господь сделает его бедным и поразит силу его в море, и сам он будет истреблен огнем.
ZECH|9|5|Увидит это Аскалон и ужаснется, и Газа, и вострепещет сильно, и Екрон; ибо посрамится надежда его: не станет царя в Газе, и Аскалон будет необитаем.
ZECH|9|6|Чужое племя будет жить в Азоте, и Я уничтожу высокомерие Филистимлян.
ZECH|9|7|Исторгну кровь из уст его и мерзости его из зубов его, и он достанется Богу нашему, и будет как тысяченачальник в Иуде, и Екрон будет, как Иевусей.
ZECH|9|8|И Я расположу стан у дома Моего против войска, против проходящих вперед и назад, и не будет более проходить притеснитель, ибо ныне Моими очами Я буду взирать на это.
ZECH|9|9|Ликуй от радости, дщерь Сиона, торжествуй, дщерь Иерусалима: се Царь твой грядет к тебе, праведный и спасающий, кроткий, сидящий на ослице и на молодом осле, сыне подъяремной.
ZECH|9|10|Тогда истреблю колесницы у Ефрема и коней в Иерусалиме, и сокрушен будет бранный лук; и Он возвестит мир народам, и владычество Его будет от моря до моря и от реки до концов земли.
ZECH|9|11|А что до тебя, ради крови завета твоего Я освобожу узников твоих изо рва, в котором нет воды.
ZECH|9|12|Возвращайтесь на твердыню вы, пленники надеющиеся! Что теперь возвещаю, воздам тебе вдвойне.
ZECH|9|13|Ибо как лук Я натяну Себе Иуду и наполню лук Ефремом, и воздвигну сынов твоих, Сион, против сынов твоих, Иония, и сделаю тебя мечом ратоборца.
ZECH|9|14|И явится над ними Господь, и как молния вылетит стрела Его, и возгремит Господь Бог трубою, и шествовать будет в бурях полуденных.
ZECH|9|15|Господь Саваоф будет защищать их, и они будут истреблять и попирать пращные камни, и будут пить и шуметь как бы от вина, и наполнятся как жертвенные чаши, как углы жертвенника.
ZECH|9|16|И спасет их Господь Бог их в тот день, как овец, народ Свой; ибо, подобно камням в венце, они воссияют на земле Его.
ZECH|9|17|О, как велика благость его и какая красота его! Хлеб одушевит язык у юношей и вино – у отроковиц!
ZECH|10|1|Просите у Господа дождя во время благопотребное; Господь блеснет молниею и даст вам обильный дождь, каждому злак на поле.
ZECH|10|2|Ибо терафимы говорят пустое, и вещуны видят ложное и рассказывают сны лживые; они утешают пустотою; поэтому они бродят как овцы, бедствуют, потому что нет пастыря.
ZECH|10|3|На пастырей воспылал гнев Мой, и козлов Я накажу; ибо посетит Господь Саваоф стадо Свое, дом Иудин, и поставит их, как славного коня Своего на брани.
ZECH|10|4|Из него будет краеугольный камень, из него – гвоздь, из него – лук для брани, из него произойдут все народоправители.
ZECH|10|5|И они будут, как герои, попирающие [врагов] на войне, как уличную грязь, и сражаться, потому что Господь с ними, и посрамят всадников на конях.
ZECH|10|6|И укреплю дом Иудин, и спасу дом Иосифов, и возвращу их, потому что Я умилосердился над ними, и они будут, как бы Я не оставлял их: ибо Я Господь Бог их, и услышу их.
ZECH|10|7|Как герой будет Ефрем; возвеселится сердце их, как от вина; и увидят это сыны их в возрадуются; в восторге будет сердце их о Господе.
ZECH|10|8|Я дам им знак и соберу их, потому что Я искупил их; они будут так же многочисленны, как прежде;
ZECH|10|9|и расселю их между народами, и в отдаленных странах они будут воспоминать обо Мне и будут жить с детьми своими, и возвратятся;
ZECH|10|10|и возвращу их из земли Египетской, и из Ассирии соберу их, и приведу их в землю Галаадскую и на Ливан, и недостанет [места] для них.
ZECH|10|11|И пройдет бедствие по морю, и поразит волны морские, и иссякнут все глубины реки, и смирится гордость Ассура, и скипетр отнимется у Египта.
ZECH|10|12|Укреплю их в Господе, и они будут ходить во имя Его, говорит Господь.
ZECH|11|1|Отворяй, Ливан, ворота твои, и да пожрет огонь кедры твои.
ZECH|11|2|Рыдай, кипарис, ибо упал кедр, ибо и величавые опустошены; рыдайте, дубы Васанские, ибо повалился непроходимый лес.
ZECH|11|3|Слышен голос рыдания пастухов, потому что опустошено приволье их; слышно рыкание молодых львов, потому что опустошена краса Иордана.
ZECH|11|4|Так говорит Господь Бог мой: паси овец, обреченных на заклание,
ZECH|11|5|которых купившие убивают ненаказанно, а продавшие говорят: "благословен Господь; я разбогател!" и пастухи их не жалеют о них.
ZECH|11|6|Ибо Я не буду более миловать жителей земли сей, говорит Господь; и вот, Я предам людей, каждого в руки ближнего его и в руки царя его, и они будут поражать землю, и Я не избавлю от рук их.
ZECH|11|7|И буду пасти овец, обреченных на заклание, овец поистине бедных. И возьму Себе два жезла, и назову один – благоволением, другой – узами, и ими буду пасти овец.
ZECH|11|8|И истреблю трех из пастырей в один месяц; и отвратится душа Моя от них, как и их душа отвращается от Меня.
ZECH|11|9|Тогда скажу: не буду пасти вас: умирающая – пусть умирает, и гибнущая – пусть гибнет, а остающиеся пусть едят плоть одна другой.
ZECH|11|10|И возьму жезл Мой – благоволения и переломлю его, чтобы уничтожить завет, который заключил Я со всеми народами.
ZECH|11|11|И он уничтожен будет в тот день, и тогда узнают бедные из овец, ожидающие Меня, что это слово Господа.
ZECH|11|12|И скажу им: если угодно вам, то дайте Мне плату Мою; если же нет, – не давайте; и они отвесят в уплату Мне тридцать сребренников.
ZECH|11|13|И сказал мне Господь: брось их в церковное хранилище, – высокая цена, в какую они оценили Меня! И взял Я тридцать сребренников и бросил их в дом Господень для горшечника.
ZECH|11|14|И переломил Я другой жезл Мой – "узы", чтобы расторгнуть братство между Иудою и Израилем.
ZECH|11|15|И Господь сказал мне: еще возьми себе снаряд одного из глупых пастухов.
ZECH|11|16|Ибо вот, Я поставлю на этой земле пастуха, который о погибающих не позаботится, потерявшихся не будет искать и больных не будет лечить, здоровых не будет кормить, а мясо тучных будет есть и копыта их оторвет.
ZECH|11|17|Горе негодному пастуху, оставляющему стадо! меч на руку его и на правый глаз его! рука его совершенно иссохнет, и правый глаз его совершенно потускнет.
ZECH|12|1|Пророческое слово Господа об Израиле. Господь, распростерший небо, основавший землю и образовавший дух человека внутри него, говорит:
ZECH|12|2|вот, Я сделаю Иерусалим чашею исступления для всех окрестных народов, и также для Иуды во время осады Иерусалима.
ZECH|12|3|И будет в тот день, сделаю Иерусалим тяжелым камнем для всех племен; все, которые будут поднимать его, надорвут себя, а соберутся против него все народы земли.
ZECH|12|4|В тот день, говорит Господь, Я поражу всякого коня бешенством и всадника его безумием, а на дом Иудин отверзу очи Мои; всякого же коня у народов поражу слепотою.
ZECH|12|5|И скажут князья Иудины в сердцах своих: сила моя – жители Иерусалима в Господе Саваофе, Боге их.
ZECH|12|6|В тот день Я сделаю князей Иудиных, как жаровню с огнем между дровами и как горящий светильник среди снопов, и они истребят все окрестные народы, справа и слева, и снова населен будет Иерусалим на своем месте, в Иерусалиме.
ZECH|12|7|И спасет Господь сначала шатры Иуды, чтобы величие дома Давидова и величие жителей Иерусалима не возносилось над Иудою.
ZECH|12|8|В тот день защищать будет Господь жителей Иерусалима, и самый слабый между ними в тот день будет как Давид, а дом Давида будет как Бог, как Ангел Господень перед ними.
ZECH|12|9|И будет в тот день, Я истреблю все народы, нападающие на Иерусалим.
ZECH|12|10|А на дом Давида и на жителей Иерусалима изолью дух благодати и умиления, и они воззрят на Него, Которого пронзили, и будут рыдать о Нем, как рыдают об единородном сыне, и скорбеть, как скорбят о первенце.
ZECH|12|11|В тот день поднимется большой плач в Иерусалиме, как плач Гададриммона в долине Мегиддонской.
ZECH|12|12|И будет рыдать земля, каждое племя особо: племя дома Давидова особо, и жены их особо; племя дома Нафанова особо, и жены их особо;
ZECH|12|13|племя дома Левиина особо, и жены их особо; племя Симеоново особо, и жены их особо.
ZECH|12|14|Все остальные племена – каждое племя особо, и жены их особо.
ZECH|13|1|В тот день откроется источник дому Давидову и жителям Иерусалима для омытия греха и нечистоты.
ZECH|13|2|И будет в тот день, говорит Господь Саваоф, Я истреблю имена идолов с этой земли, и они не будут более упоминаемы, равно как лжепророков и нечистого духа удалю с земли.
ZECH|13|3|Тогда, если кто будет прорицать, то отец его и мать его, родившие его, скажут ему: тебе не должно жить, потому что ты ложь говоришь во имя Господа; и поразят его отец его и мать его, родившие его, когда он будет прорицать.
ZECH|13|4|И будет в тот день, устыдятся такие прорицатели, каждый видения своего, когда будут прорицать, и не будут надевать на себя власяницы, чтобы обманывать.
ZECH|13|5|И каждый скажет: я не пророк, я земледелец, потому что некто сделал меня рабом от детства моего.
ZECH|13|6|Ему скажут: отчего же на руках у тебя рубцы? И он ответит: от того, что меня били в доме любящих меня.
ZECH|13|7|О, меч! поднимись на пастыря Моего и на ближнего Моего, говорит Господь Саваоф: порази пастыря, и рассеются овцы! И Я обращу руку Мою на малых.
ZECH|13|8|И будет на всей земле, говорит Господь, две части на ней будут истреблены, вымрут, а третья останется на ней.
ZECH|13|9|И введу эту третью часть в огонь, и расплавлю их, как плавят серебро, и очищу их, как очищают золото: они будут призывать имя Мое, и Я услышу их и скажу: "это Мой народ", и они скажут: "Господь – Бог мой!"
ZECH|14|1|Вот наступает день Господень, и разделят награбленное у тебя среди тебя.
ZECH|14|2|И соберу все народы на войну против Иерусалима, и взят будет город, и разграблены будут домы, и обесчещены будут жены, и половина города пойдет в плен; но остальной народ не будет истреблен из города.
ZECH|14|3|Тогда выступит Господь и ополчится против этих народов, как ополчился в день брани.
ZECH|14|4|И станут ноги Его в тот день на горе Елеонской, которая перед лицем Иерусалима к востоку; и раздвоится гора Елеонская от востока к западу весьма большою долиною, и половина горы отойдет к северу, а половина ее – к югу.
ZECH|14|5|И вы побежите в долину гор Моих, ибо долина гор будет простираться до Асила; и вы побежите, как бежали от землетрясения во дни Озии, царя Иудейского; и придет Господь Бог мой и все святые с Ним.
ZECH|14|6|И будет в тот день: не станет света, светила удалятся.
ZECH|14|7|День этот будет единственный, ведомый только Господу: ни день, ни ночь; лишь в вечернее время явится свет.
ZECH|14|8|И будет в тот день, живые воды потекут из Иерусалима, половина их к морю восточному и половина их к морю западному: летом и зимой так будет.
ZECH|14|9|И Господь будет Царем над всею землею; в тот день будет Господь един, и имя Его едино.
ZECH|14|10|Вся эта земля будет, как равнина, от Гаваона до Реммона, на юг от Иерусалима, который высоко будет стоять на своем месте и населится от ворот Вениаминовых до места первых ворот, до угловых ворот, и от башни Анамеила до царских точил.
ZECH|14|11|И будут жить в нем, и проклятия не будет более, но будет стоять Иерусалим безопасно.
ZECH|14|12|И вот какое будет поражение, которым поразит Господь все народы, которые воевали против Иерусалима: у каждого исчахнет тело его, когда он еще стоит на своих ногах, и глаза у него истают в яминах своих, и язык его иссохнет во рту у него.
ZECH|14|13|И будет в тот день: произойдет между ними великое смятение от Господа, так что один схватит руку другого, и поднимется рука его на руку ближнего его.
ZECH|14|14|Но и сам Иуда будет воевать против Иерусалима, и собрано будет богатство всех окрестных народов: золото, серебро и одежды в великом множестве.
ZECH|14|15|Будет такое же поражение и коней, и лошаков, и верблюдов, и ослов, и всякого скота, какой будет в станах у них.
ZECH|14|16|Затем все остальные из всех народов, приходивших против Иерусалима, будут приходить из года в год для поклонения Царю, Господу Саваофу, и для празднования праздника кущей.
ZECH|14|17|И будет: если какое из племен земных не пойдет в Иерусалим для поклонения Царю, Господу Саваофу, то не будет дождя у них.
ZECH|14|18|И если племя Египетское не поднимется в путь и не придет, то и у него не будет [дождя] и постигнет его поражение, каким поразит Господь народы, не приходящие праздновать праздника кущей.
ZECH|14|19|Вот что будет за грех Египта и за грех всех народов, которые не придут праздновать праздника кущей!
ZECH|14|20|В то время даже на конских уборах будет [начертано]: "Святыня Господу", и котлы в доме Господнем будут, как жертвенные чаши перед алтарем.
ZECH|14|21|И все котлы в Иерусалиме и Иудее будут святынею Господа Саваофа, и будут приходить все приносящие жертву и брать их и варить в них, и не будет более ни одного Хананея в доме Господа Саваофа в тот день.
