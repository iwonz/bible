LAM|1|1|Как одиноко сидит город, некогда многолюдный! он стал, как вдова; великий между народами, князь над областями сделался данником.
LAM|1|2|Горько плачет он ночью, и слезы его на ланитах его. Нет у него утешителя из всех, любивших его; все друзья его изменили ему, сделались врагами ему.
LAM|1|3|Иуда переселился по причине бедствия и тяжкого рабства, поселился среди язычников, и не нашел покоя; все, преследовавшие его, настигли его в тесных местах.
LAM|1|4|Пути Сиона сетуют, потому что нет идущих на праздник; все ворота его опустели; священники его вздыхают, девицы его печальны, горько и ему самому.
LAM|1|5|Враги его стали во главе, неприятели его благоденствуют, потому что Господь наслал на него горе за множество беззаконий его; дети его пошли в плен впереди врага.
LAM|1|6|И отошло от дщери Сиона все ее великолепие; князья ее – как олени, не находящие пажити; обессиленные они пошли вперед погонщика.
LAM|1|7|Вспомнил Иерусалим, во дни бедствия своего и страданий своих, о всех драгоценностях своих, какие были у него в прежние дни, тогда как народ его пал от руки врага, и никто не помогает ему; неприятели смотрят на него и смеются над его субботами.
LAM|1|8|Тяжко согрешил Иерусалим, за то и сделался отвратительным; все, прославлявшие его, смотрят на него с презрением, потому что увидели наготу его; и сам он вздыхает и отворачивается назад.
LAM|1|9|На подоле у него была нечистота, но он не помышлял о будущности своей, и поэтому необыкновенно унизился, и нет у него утешителя. "Воззри, Господи, на бедствие мое, ибо враг возвеличился!"
LAM|1|10|Враг простер руку свою на все самое драгоценное его; он видит, как язычники входят во святилище его, о котором Ты заповедал, чтобы они не вступали в собрание Твое.
LAM|1|11|Весь народ его вздыхает, ища хлеба, отдает драгоценности свои за пищу, чтобы подкрепить душу. "Воззри, Господи, и посмотри, как я унижен!"
LAM|1|12|Да не будет этого с вами, все проходящие путем! взгляните и посмотрите, есть ли болезнь, как моя болезнь, какая постигла меня, какую наслал на меня Господь в день пламенного гнева Своего?
LAM|1|13|Свыше послал Он огонь в кости мои, и он овладел ими; раскинул сеть для ног моих, опрокинул меня, сделал меня бедным и томящимся всякий день.
LAM|1|14|Ярмо беззаконий моих связано в руке Его; они сплетены и поднялись на шею мою; Он ослабил силы мои. Господь отдал меня в руки, из которых не могу подняться.
LAM|1|15|Всех сильных моих Господь низложил среди меня, созвал против меня собрание, чтобы истребить юношей моих; как в точиле, истоптал Господь деву, дочь Иуды.
LAM|1|16|Об этом плачу я; око мое, око мое изливает воды, ибо далеко от меня утешитель, который оживил бы душу мою; дети мои разорены, потому что враг превозмог.
LAM|1|17|Сион простирает руки свои, но утешителя нет ему. Господь дал повеление о Иакове врагам его окружить его; Иерусалим сделался мерзостью среди них.
LAM|1|18|Праведен Господь, ибо я непокорен был слову Его. Послушайте, все народы, и взгляните на болезнь мою: девы мои и юноши мои пошли в плен.
LAM|1|19|Зову друзей моих, но они обманули меня; священники мои и старцы мои издыхают в городе, ища пищи себе, чтобы подкрепить душу свою.
LAM|1|20|Воззри, Господи, ибо мне тесно, волнуется во мне внутренность, сердце мое перевернулось во мне за то, что я упорно противился Тебе; отвне обесчадил меня меч, а дома – как смерть.
LAM|1|21|Услышали, что я стенаю, а утешителя у меня нет; услышали все враги мои о бедствии моем и обрадовались, что Ты соделал это: о, если бы Ты повелел наступить дню, предреченному Тобою, и они стали бы подобными мне!
LAM|1|22|Да предстанет пред лице Твое вся злоба их; и поступи с ними так же, как Ты поступил со мною за все грехи мои, ибо тяжки стоны мои, и сердце мое изнемогает.
LAM|2|1|Как помрачил Господь во гневе Своем дщерь Сиона! с небес поверг на землю красу Израиля и не вспомнил о подножии ног Своих в день гнева Своего.
LAM|2|2|Погубил Господь все жилища Иакова, не пощадил, разрушил в ярости Своей укрепления дщери Иудиной, поверг на землю, отверг царство и князей его, как нечистых:
LAM|2|3|в пылу гнева сломил все роги Израилевы, отвел десницу Свою от неприятеля и воспылал в Иакове, как палящий огонь, пожиравший все вокруг;
LAM|2|4|натянул лук Свой, как неприятель, направил десницу Свою, как враг, и убил все, вожделенное для глаз; на скинию дщери Сиона излил ярость Свою, как огонь.
LAM|2|5|Господь стал как неприятель, истребил Израиля, разорил все чертоги его, разрушил укрепления его и распространил у дщери Иудиной сетование и плач.
LAM|2|6|И отнял ограду Свою, как у сада; разорил Свое место собраний, заставил Господь забыть на Сионе празднества и субботы; и в негодовании гнева Своего отверг царя и священника.
LAM|2|7|Отверг Господь жертвенник Свой, отвратил сердце Свое от святилища Своего, предал в руки врагов стены чертогов его; в доме Господнем они шумели, как в праздничный день.
LAM|2|8|Господь определил разрушить стену дщери Сиона, протянул вервь, не отклонил руки Своей от разорения; истребил внешние укрепления, и стены вместе разрушены.
LAM|2|9|Ворота ее вдались в землю; Он разрушил и сокрушил запоры их; царь ее и князья ее – среди язычников; не стало закона, и пророки ее не сподобляются видений от Господа.
LAM|2|10|Сидят на земле безмолвно старцы дщери Сионовой, посыпали пеплом свои головы, препоясались вретищем; опустили к земле головы свои девы Иерусалимские.
LAM|2|11|Истощились от слез глаза мои, волнуется во мне внутренность моя, изливается на землю печень моя от гибели дщери народа моего, когда дети и грудные младенцы умирают от голода среди городских улиц.
LAM|2|12|Матерям своим говорят они: "где хлеб и вино?", умирая, подобно раненым, на улицах городских, изливая души свои в лоно матерей своих.
LAM|2|13|Что мне сказать тебе, с чем сравнить тебя, дщерь Иерусалима? чему уподобить тебя, чтобы утешить тебя, дева, дщерь Сиона? ибо рана твоя велика, как море; кто может исцелить тебя?
LAM|2|14|Пророки твои провещали тебе пустое и ложное и не раскрывали твоего беззакония, чтобы отвратить твое пленение, и изрекали тебе откровения ложные и приведшие тебя к изгнанию.
LAM|2|15|Руками всплескивают о тебе все проходящие путем, свищут и качают головою своею о дщери Иерусалима, говоря: "это ли город, который называли совершенством красоты, радостью всей земли?"
LAM|2|16|Разинули на тебя пасть свою все враги твои, свищут и скрежещут зубами, говорят: "поглотили мы его, только этого дня и ждали мы, дождались, увидели!"
LAM|2|17|Совершил Господь, что определил, исполнил слово Свое, изреченное в древние дни, разорил без пощады и дал врагу порадоваться над тобою, вознес рог неприятелей твоих.
LAM|2|18|Сердце их вопиет к Господу: стена дщери Сиона! лей ручьем слезы день и ночь, не давай себе покоя, не спускай зениц очей твоих.
LAM|2|19|Вставай, взывай ночью, при начале каждой стражи; изливай, как воду, сердце твое пред лицем Господа; простирай к Нему руки твои о душе детей твоих, издыхающих от голода на углах всех улиц.
LAM|2|20|"Воззри, Господи, и посмотри: кому Ты сделал так, чтобы женщины ели плод свой, младенцев, вскормленных ими? чтобы убиваемы были в святилище Господнем священник и пророк?
LAM|2|21|Дети и старцы лежат на земле по улицам; девы мои и юноши мои пали от меча; Ты убивал их в день гнева Твоего, заколал без пощады.
LAM|2|22|Ты созвал отовсюду, как на праздник, ужасы мои, и в день гнева Господня никто не спасся, никто не уцелел; тех, которые были мною вскормлены и вырощены, враг мой истребил".
LAM|3|1|Я человек, испытавший горе от жезла гнева Его.
LAM|3|2|Он повел меня и ввел во тьму, а не во свет.
LAM|3|3|Так, Он обратился на меня и весь день обращает руку Свою;
LAM|3|4|измождил плоть мою и кожу мою, сокрушил кости мои;
LAM|3|5|огородил меня и обложил горечью и тяготою;
LAM|3|6|посадил меня в темное место, как давно умерших;
LAM|3|7|окружил меня стеною, чтобы я не вышел, отяготил оковы мои,
LAM|3|8|и когда я взывал и вопиял, задерживал молитву мою;
LAM|3|9|каменьями преградил дороги мои, извратил стези мои.
LAM|3|10|Он стал для меня как бы медведь в засаде, [как бы] лев в скрытном месте;
LAM|3|11|извратил пути мои и растерзал меня, привел меня в ничто;
LAM|3|12|натянул лук Свой и поставил меня как бы целью для стрел;
LAM|3|13|послал в почки мои стрелы из колчана Своего.
LAM|3|14|Я стал посмешищем для всего народа моего, вседневною песнью их.
LAM|3|15|Он пресытил меня горечью, напоил меня полынью.
LAM|3|16|Сокрушил камнями зубы мои, покрыл меня пеплом.
LAM|3|17|И удалился мир от души моей; я забыл о благоденствии,
LAM|3|18|и сказал я: погибла сила моя и надежда моя на Господа.
LAM|3|19|Помысли о моем страдании и бедствии моем, о полыни и желчи.
LAM|3|20|Твердо помнит это душа моя и падает во мне.
LAM|3|21|Вот что я отвечаю сердцу моему и потому уповаю:
LAM|3|22|по милости Господа мы не исчезли, ибо милосердие Его не истощилось.
LAM|3|23|Оно обновляется каждое утро; велика верность Твоя!
LAM|3|24|Господь часть моя, говорит душа моя, итак буду надеяться на Него.
LAM|3|25|Благ Господь к надеющимся на Него, к душе, ищущей Его.
LAM|3|26|Благо тому, кто терпеливо ожидает спасения от Господа.
LAM|3|27|Благо человеку, когда он несет иго в юности своей;
LAM|3|28|сидит уединенно и молчит, ибо Он наложил его на него;
LAM|3|29|полагает уста свои в прах, [помышляя]: "может быть, еще есть надежда";
LAM|3|30|подставляет ланиту свою биющему его, пресыщается поношением,
LAM|3|31|ибо не навек оставляет Господь.
LAM|3|32|Но послал горе, и помилует по великой благости Своей.
LAM|3|33|Ибо Он не по изволению сердца Своего наказывает и огорчает сынов человеческих.
LAM|3|34|Но, когда попирают ногами своими всех узников земли,
LAM|3|35|когда неправедно судят человека пред лицем Всевышнего,
LAM|3|36|когда притесняют человека в деле его: разве не видит Господь?
LAM|3|37|Кто это говорит: "и то бывает, чему Господь не повелел быть"?
LAM|3|38|Не от уст ли Всевышнего происходит бедствие и благополучие?
LAM|3|39|Зачем сетует человек живущий? всякий сетуй на грехи свои.
LAM|3|40|Испытаем и исследуем пути свои, и обратимся к Господу.
LAM|3|41|Вознесем сердце наше и руки к Богу, [сущему] на небесах:
LAM|3|42|мы отпали и упорствовали; Ты не пощадил.
LAM|3|43|Ты покрыл Себя гневом и преследовал нас, умерщвлял, не щадил;
LAM|3|44|Ты закрыл Себя облаком, чтобы не доходила молитва наша;
LAM|3|45|сором и мерзостью Ты сделал нас среди народов.
LAM|3|46|Разинули на нас пасть свою все враги наши.
LAM|3|47|Ужас и яма, опустошение и разорение – доля наша.
LAM|3|48|Потоки вод изливает око мое о гибели дщери народа моего.
LAM|3|49|Око мое изливается и не перестает, ибо нет облегчения,
LAM|3|50|доколе не призрит и не увидит Господь с небес.
LAM|3|51|Око мое опечаливает душу мою ради всех дщерей моего города.
LAM|3|52|Всячески усиливались уловить меня, как птичку, враги мои, без всякой причины;
LAM|3|53|повергли жизнь мою в яму и закидали меня камнями.
LAM|3|54|Воды поднялись до головы моей; я сказал: "погиб я".
LAM|3|55|Я призывал имя Твое, Господи, из ямы глубокой.
LAM|3|56|Ты слышал голос мой; не закрой уха Твоего от воздыхания моего, от вопля моего.
LAM|3|57|Ты приближался, когда я взывал к Тебе, и говорил: "не бойся".
LAM|3|58|Ты защищал, Господи, дело души моей; искуплял жизнь мою.
LAM|3|59|Ты видишь, Господи, обиду мою; рассуди дело мое.
LAM|3|60|Ты видишь всю мстительность их, все замыслы их против меня.
LAM|3|61|Ты слышишь, Господи, ругательство их, все замыслы их против меня,
LAM|3|62|речи восстающих на меня и их ухищрения против меня всякий день.
LAM|3|63|Воззри, сидят ли они, встают ли, я для них – песнь.
LAM|3|64|Воздай им, Господи, по делам рук их;
LAM|3|65|пошли им помрачение сердца и проклятие Твое на них;
LAM|3|66|преследуй их, Господи, гневом, и истреби их из поднебесной.
LAM|4|1|Как потускло золото, изменилось золото наилучшее! камни святилища раскиданы по всем перекресткам.
LAM|4|2|Сыны Сиона драгоценные, равноценные чистейшему золоту, как они сравнены с глиняною посудою, изделием рук горшечника!
LAM|4|3|И чудовища подают сосцы и кормят своих детенышей, а дщерь народа моего стала жестока подобно страусам в пустыне.
LAM|4|4|Язык грудного младенца прилипает к гортани его от жажды; дети просят хлеба, и никто не подает им.
LAM|4|5|Евшие сладкое истаевают на улицах; воспитанные на багрянице жмутся к навозу.
LAM|4|6|Наказание нечестия дщери народа моего превышает казнь за грехи Содома: тот низринут мгновенно, и руки человеческие не касались его.
LAM|4|7|Князья ее [были] в ней чище снега, белее молока; они были телом краше коралла, вид их был, как сапфир;
LAM|4|8|а теперь темнее всего черного лице их; не узнают их на улицах; кожа их прилипла к костям их, стала суха, как дерево.
LAM|4|9|Умерщвляемые мечом счастливее умерщвляемых голодом, потому что сии истаевают, поражаемые недостатком плодов полевых.
LAM|4|10|Руки мягкосердых женщин варили детей своих, чтобы они были для них пищею во время гибели дщери народа моего.
LAM|4|11|Совершил Господь гнев Свой, излил ярость гнева Своего и зажег на Сионе огонь, который пожрал основания его.
LAM|4|12|Не верили цари земли и все живущие во вселенной, чтобы враг и неприятель вошел во врата Иерусалима.
LAM|4|13|[Все это] – за грехи лжепророков его, за беззакония священников его, которые среди него проливали кровь праведников;
LAM|4|14|бродили как слепые по улицам, осквернялись кровью, так что невозможно было прикоснуться к одеждам их.
LAM|4|15|"Сторонитесь! нечистый!" кричали им; "сторонитесь, сторонитесь, не прикасайтесь"; и они уходили в смущении; а между народом говорили: "их более не будет!
LAM|4|16|лице Господне рассеет их; Он уже не призрит на них", потому что они лица священников не уважают, старцев не милуют.
LAM|4|17|Наши глаза истомлены в напрасном ожидании помощи; со сторожевой башни нашей мы ожидали народ, который не мог спасти нас.
LAM|4|18|А они подстерегали шаги наши, чтобы мы не могли ходить по улицам нашим; приблизился конец наш, дни наши исполнились; пришел конец наш.
LAM|4|19|Преследовавшие нас были быстрее орлов небесных; гонялись за нами по горам, ставили засаду для нас в пустыне.
LAM|4|20|Дыхание жизни нашей, помазанник Господень пойман в ямы их, тот, о котором мы говорили: "под тенью его будем жить среди народов".
LAM|4|21|Радуйся и веселись, дочь Едома, обитательница земли Уц! И до тебя дойдет чаша; напьешься допьяна и обнажишься.
LAM|4|22|Дщерь Сиона! наказание за беззаконие твое кончилось; Он не будет более изгонять тебя; но твое беззаконие, дочь Едома, Он посетит и обнаружит грехи твои.
LAM|5|1|Вспомни, Господи, что над нами совершилось; призри и посмотри на поругание наше.
LAM|5|2|Наследие наше перешло к чужим, домы наши – к иноплеменным;
LAM|5|3|мы сделались сиротами, без отца; матери наши – как вдовы.
LAM|5|4|Воду свою пьем за серебро, дрова наши достаются нам за деньги.
LAM|5|5|Нас погоняют в шею, мы работаем, [и] не имеем отдыха.
LAM|5|6|Протягиваем руку к Египтянам, к Ассириянам, чтобы насытиться хлебом.
LAM|5|7|Отцы наши грешили: их уже нет, а мы несем наказание за беззакония их.
LAM|5|8|Рабы господствуют над нами, и некому избавить от руки их.
LAM|5|9|С опасностью жизни от меча, в пустыне достаем хлеб себе.
LAM|5|10|Кожа наша почернела, как печь, от жгучего голода.
LAM|5|11|Жен бесчестят на Сионе, девиц – в городах Иудейских.
LAM|5|12|Князья повешены руками их, лица старцев не уважены.
LAM|5|13|Юношей берут к жерновам, и отроки падают под ношами дров.
LAM|5|14|Старцы уже не сидят у ворот; юноши не поют.
LAM|5|15|Прекратилась радость сердца нашего; хороводы наши обратились в сетование.
LAM|5|16|Упал венец с головы нашей; горе нам, что мы согрешили!
LAM|5|17|От сего–то изнывает сердце наше; от сего померкли глаза наши.
LAM|5|18|От того, что опустела гора Сион, лисицы ходят по ней.
LAM|5|19|Ты, Господи, пребываешь во веки; престол Твой – в род и род.
LAM|5|20|Для чего совсем забываешь нас, оставляешь нас на долгое время?
LAM|5|21|Обрати нас к Тебе, Господи, и мы обратимся; обнови дни наши, как древле.
LAM|5|22|Неужели Ты совсем отверг нас, прогневался на нас безмерно?
