LAM|1|1|ALEPH quomodo sedit sola civitas plena populo facta est quasi vidua domina gentium princeps provinciarum facta est sub tributo
LAM|1|2|BETH plorans ploravit in nocte et lacrimae eius in maxillis eius non est qui consoletur eam ex omnibus caris eius omnes amici eius spreverunt eam et facti sunt ei inimici
LAM|1|3|GIMEL migravit Iuda propter adflictionem et multitudinem servitutis habitavit inter gentes nec invenit requiem omnes persecutores eius adprehenderunt eam inter angustias
LAM|1|4|DELETH viae Sion lugent eo quod non sint qui veniant ad sollemnitatem omnes portae eius destructae sacerdotes eius gementes virgines eius squalidae et ipsa oppressa amaritudine
LAM|1|5|HE facti sunt hostes eius in capite inimici illius locupletati sunt quia Dominus locutus est super eam propter multitudinem iniquitatum eius parvuli eius ducti sunt captivi ante faciem tribulantis
LAM|1|6|VAV et egressus est a filia Sion omnis decor eius facti sunt principes eius velut arietes non invenientes pascuam et abierunt absque fortitudine ante faciem subsequentis
LAM|1|7|ZAI recordata est Hierusalem dierum adflictionis suae et praevaricationis omnium desiderabilium suorum quae habuerat a diebus antiquis cum caderet populus eius in manu hostili et non esset auxiliator viderunt eam hostes et deriserunt sabbata eius
LAM|1|8|HETH peccatum peccavit Hierusalem propterea instabilis facta est omnes qui glorificabant eam spreverunt illam quia viderunt ignominiam eius ipsa autem gemens et conversa retrorsum
LAM|1|9|TETH sordes eius in pedibus eius nec recordata est finis sui deposita est vehementer non habens consolatorem vide Domine adflictionem meam quoniam erectus est inimicus
LAM|1|10|IOTH manum suam misit hostis ad omnia desiderabilia eius quia vidit gentes ingressas sanctuarium suum de quibus praeceperas ne intrarent in ecclesiam tuam
LAM|1|11|CAPH omnis populus eius gemens et quaerens panem dederunt pretiosa quaeque pro cibo ad refocilandam animam vide Domine considera quoniam facta sum vilis
LAM|1|12|LAMED o vos omnes qui transitis per viam adtendite et videte si est dolor sicut dolor meus quoniam vindemiavit me ut locutus est Dominus in die irae furoris sui
LAM|1|13|MEM de excelso misit ignem in ossibus meis et erudivit me expandit rete pedibus meis convertit me retrorsum posuit me desolatam tota die maerore confectam
LAM|1|14|NUN vigilavit iugum iniquitatum mearum in manu eius convolutae sunt et inpositae collo meo infirmata est virtus mea dedit me Dominus in manu de qua non potero surgere
LAM|1|15|SAMECH abstulit omnes magnificos meos Dominus de medio mei vocavit adversum me tempus ut contereret electos meos torcular calcavit Dominus virgini filiae Iuda
LAM|1|16|AIN idcirco ego plorans et oculus meus deducens aquam quia longe factus est a me consolator convertens animam meam facti sunt filii mei perditi quoniam invaluit inimicus
LAM|1|17|FE expandit Sion manus suas non est qui consoletur eam mandavit Dominus adversum Iacob in circuitu eius hostes eius facta est Hierusalem quasi polluta menstruis inter eos
LAM|1|18|SADE iustus est Dominus quia os eius ad iracundiam provocavi audite obsecro universi populi et videte dolorem meum virgines meae et iuvenes mei abierunt in captivitatem
LAM|1|19|COPH vocavi amicos meos et ipsi deceperunt me sacerdotes mei et senes mei in urbe consumpti sunt quia quaesierunt cibum sibi ut refocilarent animam suam
LAM|1|20|RES vide Domine quoniam tribulor venter meus conturbatus est subversum est cor meum in memet ipsa quoniam amaritudine plena sum foris interfecit gladius et domi mors similis est
LAM|1|21|SEN audierunt quia ingemesco ego et non est qui consoletur me omnes inimici mei audierunt malum meum laetati sunt quoniam tu fecisti adduxisti diem consolationis et fient similes mei
LAM|1|22|THAU ingrediatur omne malum eorum coram te et devindemia eos sicut vindemiasti me propter omnes iniquitates meas multi enim gemitus mei et cor meum maerens
LAM|2|1|ALEPH quomodo obtexit caligine in furore suo Dominus filiam Sion proiecit de caelo terram inclitam Israhel et non recordatus est scabilli pedum suorum in die furoris sui
LAM|2|2|BETH praecipitavit Dominus nec pepercit omnia speciosa Iacob destruxit in furore suo munitiones virginis Iuda deiecit in terram polluit regnum et principes eius
LAM|2|3|GIMEL confregit in ira furoris omne cornu Israhel avertit retrorsum dexteram suam a facie inimici et succendit in Iacob quasi ignem flammae devorantis in gyro
LAM|2|4|DELETH tetendit arcum suum quasi inimicus firmavit dexteram suam quasi hostis et occidit omne quod pulchrum erat visu in tabernaculo filiae Sion effudit quasi ignem indignationem suam
LAM|2|5|HE factus est Dominus velut inimicus praecipitavit Israhel praecipitavit omnia moenia eius dissipavit munitiones eius et replevit in filia Iuda humiliatum et humiliatam
LAM|2|6|VAV et dissipavit quasi hortum tentorium suum demolitus est tabernaculum suum oblivioni tradidit Dominus in Sion festivitatem et sabbatum et obprobrio in indignatione furoris sui regem et sacerdotem
LAM|2|7|ZAI reppulit Dominus altare suum maledixit sanctificationi suae tradidit in manu inimici muros turrium eius vocem dederunt in domo Domini sicut in die sollemni
LAM|2|8|HETH cogitavit Dominus dissipare murum filiae Sion tetendit funiculum suum et non avertit manum suam a perditione luxitque antemurale et murus pariter dissipatus est
LAM|2|9|TETH defixae sunt in terra portae eius perdidit et contrivit vectes eius regem eius et principes eius in gentibus non est lex et prophetae eius non invenerunt visionem a Domino
LAM|2|10|IOTH sederunt in terra conticuerunt senes filiae Sion consperserunt cinere capita sua accincti sunt ciliciis abiecerunt in terra capita sua virgines Hierusalem
LAM|2|11|CAPH defecerunt prae lacrimis oculi mei conturbata sunt viscera mea effusum est in terra iecur meum super contritione filiae populi mei cum deficeret parvulus et lactans in plateis oppidi
LAM|2|12|LAMED matribus suis dixerunt ubi est triticum et vinum cum deficerent quasi vulnerati in plateis civitatis cum exhalarent animas suas in sinu matrum suarum
LAM|2|13|MEM cui conparabo te vel cui adsimilabo te filia Hierusalem cui exaequabo te et consolabor te virgo filia Sion magna enim velut mare contritio tua quis medebitur tui
LAM|2|14|NUN prophetae tui viderunt tibi falsa et stulta nec aperiebant iniquitatem tuam ut te ad paenitentiam provocarent viderunt autem tibi adsumptiones falsas et eiectiones
LAM|2|15|SAMECH plauserunt super te manibus omnes transeuntes per viam sibilaverunt et moverunt caput suum super filiam Hierusalem haecine est urbs dicentes perfecti decoris gaudium universae terrae
LAM|2|16|FE aperuerunt super te os suum omnes inimici tui sibilaverunt et fremuerunt dentibus dixerunt devoravimus en ista est dies quam expectabamus invenimus vidimus
LAM|2|17|AIN fecit Dominus quae cogitavit conplevit sermonem suum quem praeceperat a diebus antiquis destruxit et non pepercit et laetificavit super te inimicum et exaltavit cornu hostium tuorum
LAM|2|18|SADE clamavit cor eorum ad Dominum super muros filiae Sion deduc quasi torrentem lacrimas per diem et per noctem non des requiem tibi neque taceat pupilla oculi tui
LAM|2|19|COPH consurge lauda in nocte in principio vigiliarum effunde sicut aqua cor tuum ante conspectum Domini leva ad eum manus tuas pro anima parvulorum tuorum qui defecerunt in fame in capite omnium conpetorum
LAM|2|20|RES vide Domine et considera quem vindemiaveris ita ergone comedent mulieres fructum suum parvulos ad mensuram palmae si occidetur in sanctuario Domini sacerdos et propheta
LAM|2|21|SEN iacuerunt in terra foris puer et senex virgines meae et iuvenes mei ceciderunt in gladio interfecisti in die furoris tui percussisti nec misertus es
LAM|2|22|THAU vocasti quasi ad diem sollemnem qui terrerent me de circuitu et non fuit in die furoris Domini qui effugeret et relinqueretur quos educavi et enutrivi inimicus meus consumpsit eos
LAM|3|1|ALEPH ego vir videns paupertatem meam in virga indignationis eius
LAM|3|2|ALEPH me minavit et adduxit in tenebris et non in lucem
LAM|3|3|ALEPH tantum in me vertit et convertit manum suam tota die
LAM|3|4|BETH vetustam fecit pellem meam et carnem meam contrivit ossa mea
LAM|3|5|BETH aedificavit in gyro meo et circumdedit me felle et labore
LAM|3|6|BETH in tenebrosis conlocavit me quasi mortuos sempiternos
LAM|3|7|GIMEL circumaedificavit adversum me ut non egrediar adgravavit conpedem meam
LAM|3|8|GIMEL sed et cum clamavero et rogavero exclusit orationem meam
LAM|3|9|GIMEL conclusit vias meas lapidibus quadris semitas meas subvertit
LAM|3|10|DELETH ursus insidians factus est mihi leo in absconditis
LAM|3|11|DELETH semitas meas subvertit et confregit me posuit me desolatam
LAM|3|12|DELETH tetendit arcum suum et posuit me quasi signum ad sagittam
LAM|3|13|HE misit in renibus meis filias faretrae suae
LAM|3|14|HE factus sum in derisu omni populo meo canticum eorum tota die
LAM|3|15|HE replevit me amaritudinibus inebriavit me absinthio
LAM|3|16|VAV et fregit ad numerum dentes meos cibavit me cinere
LAM|3|17|VAV et repulsa est anima mea oblitus sum bonorum
LAM|3|18|VAV et dixi periit finis meus et spes mea a Domino
LAM|3|19|ZAI recordare paupertatis et transgressionis meae absinthii et fellis
LAM|3|20|ZAI memoria memor ero et tabescet in me anima mea
LAM|3|21|ZAI hoc recolens in corde meo ideo sperabo
LAM|3|22|HETH misericordiae Domini quia non sumus consumpti quia non defecerunt miserationes eius
LAM|3|23|HETH novae diluculo multa est fides tua
LAM|3|24|HETH pars mea Dominus dixit anima mea propterea expectabo eum
LAM|3|25|TETH bonus est Dominus sperantibus in eum animae quaerenti illum
LAM|3|26|TETH bonum est praestolari cum silentio salutare Domini
LAM|3|27|TETH bonum est viro cum portaverit iugum ab adulescentia sua
LAM|3|28|IOTH sedebit solitarius et tacebit quia levavit super se
LAM|3|29|IOTH ponet in pulvere os suum si forte sit spes
LAM|3|30|IOTH dabit percutienti se maxillam saturabitur obprobriis
LAM|3|31|CAPH quia non repellet in sempiternum Dominus
LAM|3|32|CAPH quia si abiecit et miserebitur secundum multitudinem misericordiarum suarum
LAM|3|33|CAPH non enim humiliavit ex corde suo et abiecit filios hominis
LAM|3|34|LAMED ut contereret sub pedibus suis omnes vinctos terrae
LAM|3|35|LAMED ut declinaret iudicium viri in conspectu vultus Altissimi
LAM|3|36|LAMED ut perverteret hominem in iudicio suo Dominus ignoravit
LAM|3|37|MEM quis est iste qui dixit ut fieret Domino non iubente
LAM|3|38|MEM ex ore Altissimi non egredientur nec mala nec bona
LAM|3|39|MEM quid murmuravit homo vivens vir pro peccatis suis
LAM|3|40|NUN scrutemur vias nostras et quaeramus et revertamur ad Dominum
LAM|3|41|NUN levemus corda nostra cum manibus ad Dominum in caelos
LAM|3|42|NUN nos inique egimus et ad iracundiam provocavimus idcirco tu inexorabilis es
LAM|3|43|SAMECH operuisti in furore et percussisti nos occidisti nec pepercisti
LAM|3|44|SAMECH opposuisti nubem tibi ne transeat oratio
LAM|3|45|SAMECH eradicationem et abiectionem posuisti me in medio populorum
LAM|3|46|FE aperuerunt super nos os suum omnes inimici
LAM|3|47|FE formido et laqueus facta est nobis vaticinatio et contritio
LAM|3|48|FE divisiones aquarum deduxit oculus meus in contritione filiae populi mei
LAM|3|49|AIN oculus meus adflictus est nec tacuit eo quod non esset requies
LAM|3|50|AIN donec respiceret et videret Dominus de caelis
LAM|3|51|AIN oculus meus depraedatus est animam meam in cunctis filiabus urbis meae
LAM|3|52|SADE venatione ceperunt me quasi avem inimici mei gratis
LAM|3|53|SADE lapsa est in lacu vita mea et posuerunt lapidem super me
LAM|3|54|SADE inundaverunt aquae super caput meum dixi perii
LAM|3|55|COPH invocavi nomen tuum Domine de lacis novissimis
LAM|3|56|COPH vocem meam audisti ne avertas aurem tuam a singultu meo et clamoribus
LAM|3|57|COPH adpropinquasti in die quando invocavi te dixisti ne timeas
LAM|3|58|RES iudicasti Domine causam animae meae redemptor vitae meae
LAM|3|59|RES vidisti Domine iniquitatem adversum me iudica iudicium meum
LAM|3|60|RES vidisti omnem furorem universas cogitationes eorum adversum me
LAM|3|61|SEN audisti obprobria eorum Domine omnes cogitationes eorum adversum me
LAM|3|62|SEN labia insurgentium mihi et meditationes eorum adversum me tota die
LAM|3|63|SEN sessionem eorum et resurrectionem eorum vide ego sum psalmus eorum
LAM|3|64|THAU reddes eis vicem Domine iuxta opera manuum suarum
LAM|3|65|THAU dabis eis scutum cordis laborem tuum
LAM|3|66|THAU persequeris in furore et conteres eos sub caelis Domine
LAM|4|1|ALEPH quomodo obscuratum est aurum mutatus est color optimus dispersi sunt lapides sanctuarii in capite omnium platearum
LAM|4|2|BETH filii Sion incliti et amicti auro primo quomodo reputati sunt in vasa testea opus manuum figuli
LAM|4|3|GIMEL sed et lamiae nudaverunt mammam lactaverunt catulos suos filia populi mei crudelis quasi strutio in deserto
LAM|4|4|DELETH adhesit lingua lactantis ad palatum eius in siti parvuli petierunt panem et non erat qui frangeret eis
LAM|4|5|HE qui vescebantur voluptuose interierunt in viis qui nutriebantur in croceis amplexati sunt stercora
LAM|4|6|VAV et maior effecta est iniquitas filiae populi mei peccato Sodomorum quae subversa est in momento et non ceperunt in ea manus
LAM|4|7|ZAI candidiores nazarei eius nive nitidiores lacte rubicundiores ebore antiquo sapphyro pulchriores
LAM|4|8|HETH denigrata est super carbones facies eorum et non sunt cogniti in plateis adhesit cutis eorum ossibus aruit et facta est quasi lignum
LAM|4|9|TETH melius fuit occisis gladio quam interfectis fame quoniam isti extabuerunt consumpti ab sterilitate terrae
LAM|4|10|IOTH manus mulierum misericordium coxerunt filios suos facti sunt cibus earum in contritione filiae populi mei
LAM|4|11|CAPH conplevit Dominus furorem suum effudit iram indignationis suae et succendit ignem in Sion et devoravit fundamenta eius
LAM|4|12|LAMED non crediderunt reges terrae et universi habitatores orbis quoniam ingrederetur hostis et inimicus per portas Hierusalem
LAM|4|13|MEM propter peccata prophetarum eius iniquitates sacerdotum eius qui effuderunt in medio eius sanguinem iustorum
LAM|4|14|NUN erraverunt caeci in plateis polluti sunt sanguine cumque non possent tenuerunt lacinias suas
LAM|4|15|SAMECH recedite polluti clamaverunt eis recedite abite nolite tangere iurgati quippe sunt et commoti dixerunt inter gentes non addet ultra ut habitet in eis
LAM|4|16|FE facies Domini divisit eos non addet ut respiciat eos facies sacerdotum non erubuerunt neque senum miserti sunt
LAM|4|17|AIN cum adhuc subsisteremus defecerunt oculi nostri ad auxilium nostrum vanum cum respiceremus adtenti ad gentem quae salvare non poterat
LAM|4|18|SADE lubricaverunt vestigia nostra in itinere platearum nostrarum adpropinquavit finis noster conpleti sunt dies nostri quia venit finis noster
LAM|4|19|COPH velociores fuerunt persecutores nostri aquilis caeli super montes persecuti sunt nos in deserto insidiati sunt nobis
LAM|4|20|RES spiritus oris nostri christus dominus captus est in peccatis nostris cui diximus in umbra tua vivemus in gentibus
LAM|4|21|SEN gaude et laetare filia Edom quae habitas in terra Hus ad te quoque perveniet calix inebriaberis atque nudaberis
LAM|4|22|THAU conpleta est iniquitas tua filia Sion non addet ultra ut transmigret te visitavit iniquitatem tuam filia Edom discoperuit peccata tua
LAM|5|1|recordare Domine quid acciderit nobis intuere et respice obprobrium nostrum
LAM|5|2|hereditas nostra versa est ad alienos domus nostrae ad extraneos
LAM|5|3|pupilli facti sumus absque patre matres nostrae quasi viduae
LAM|5|4|aquam nostram pecunia bibimus ligna nostra pretio conparavimus
LAM|5|5|cervicibus minabamur lassis non dabatur requies
LAM|5|6|Aegypto dedimus manum et Assyriis ut saturaremur pane
LAM|5|7|patres nostri peccaverunt et non sunt et nos iniquitates eorum portavimus
LAM|5|8|servi dominati sunt nostri non fuit qui redimeret de manu eorum
LAM|5|9|in animabus nostris adferebamus panem nobis a facie gladii in deserto
LAM|5|10|pellis nostra quasi clibanus exusta est a facie tempestatum famis
LAM|5|11|mulieres in Sion humiliaverunt virgines in civitatibus Iuda
LAM|5|12|principes manu suspensi sunt facies senum non erubuerunt
LAM|5|13|adulescentibus inpudice abusi sunt et pueri in ligno corruerunt
LAM|5|14|senes de portis defecerunt iuvenes de choro psallentium
LAM|5|15|defecit gaudium cordis nostri versus est in luctu chorus noster
LAM|5|16|cecidit corona capitis nostri vae nobis quia peccavimus
LAM|5|17|propterea maestum factum est cor nostrum ideo contenebrati sunt oculi nostri
LAM|5|18|propter montem Sion quia disperiit vulpes ambulaverunt in eo
LAM|5|19|tu autem Domine in aeternum permanebis solium tuum in generatione et generatione
LAM|5|20|quare in perpetuum oblivisceris nostri derelinques nos in longitudinem dierum
LAM|5|21|converte nos Domine ad te et convertemur innova dies nostros sicut a principio
LAM|5|22|sed proiciens reppulisti nos iratus es contra nos vehementer
