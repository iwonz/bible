PS|1|1|不從惡人的計謀， 不站罪人的道路， 不坐傲慢人的座位， 惟喜愛耶和華的律法， 晝夜思想 他的律法； 這人便為有福！
PS|1|2|
PS|1|3|他要像一棵樹栽在溪水旁， 按時候結果子， 葉子也不枯乾。 凡他所做的盡都順利。
PS|1|4|惡人並不是這樣， 卻像糠秕被風吹散。
PS|1|5|因此，當審判的時候惡人必站立不住， 罪人在義人的會眾中也是如此。
PS|1|6|因為耶和華知道義人的道路， 惡人的道路卻必滅亡。
PS|2|1|列國為甚麼爭鬧？ 萬民為甚麼圖謀虛妄？
PS|2|2|世上的君王都站穩， 臣宰一同算計， 要對抗耶和華， 對抗他的受膏者：
PS|2|3|「我們要掙脫他們的捆綁， 脫去他們的繩索。」
PS|2|4|那坐在天上的必譏笑， 主必嗤笑他們。
PS|2|5|那時，他要在怒中責備他們， 在烈怒中驚嚇他們：
PS|2|6|「我已經在 錫安 －我的聖山 膏立了我的君王。」
PS|2|7|我要傳耶和華的聖旨， 他對我說：「你是我的兒子， 我今日生了你。
PS|2|8|你求我，我就將列國賜你為基業， 將地極賜你為田產。
PS|2|9|你必用鐵杖打破他們， 把他們如同陶匠的瓦器摔碎。」
PS|2|10|現在，君王啊，應當謹慎！ 世上的審判官哪，要聽勸戒！
PS|2|11|當存敬畏的心事奉耶和華， 又當戰兢而快樂。
PS|2|12|當親吻兒子，免得他發怒， 你們就在半途中滅亡， 因為他的怒氣快要發作。 凡投靠他的，都是有福的。
PS|3|1|耶和華啊，我的敵人何其增多！ 許多人起來攻擊我。
PS|3|2|許多人議論我： 「他得不到上帝的幫助。」（細拉）
PS|3|3|但你－耶和華是我四圍的盾牌， 是我的榮耀，又是令我抬起頭來的。
PS|3|4|我用我的聲音求告耶和華， 他就從他的聖山上應允我。（細拉）
PS|3|5|我躺下，我睡覺，我醒來， 耶和華都保佑我。
PS|3|6|雖有成萬的百姓周圍攻擊我， 我也不懼怕。
PS|3|7|耶和華啊，求你興起！ 我的上帝啊，求你救我！ 因為你打斷我所有仇敵的腮骨， 敲碎了惡人的牙齒。
PS|3|8|救恩屬於耶和華； 願你賜福給你的百姓。（細拉）
PS|4|1|顯我為義的上帝啊， 我呼求的時候，求你應允我！ 我在困境中，你曾使我寬暢； 求你憐憫我，聽我的禱告！
PS|4|2|你們這些人哪，你們把我的尊榮變為羞辱，要到幾時呢？ 你們喜愛虛妄，尋找虛假，要到幾時呢？ （細拉）
PS|4|3|你們要知道，耶和華已將虔誠人分別出來歸他自己； 我求告耶和華，他必垂聽。
PS|4|4|應當畏懼，不可犯罪； 在床上的時候，要心裏思想，並要安靜。（細拉）
PS|4|5|當獻上公義的祭， 又當倚靠耶和華。
PS|4|6|有許多人說：「誰能指示我們甚麼好處？ 耶和華啊，求你用你臉上的光照耀我們。」
PS|4|7|你使我心裏喜樂， 勝過那豐收五穀新酒的人。
PS|4|8|我必平安地躺下睡覺， 因為獨有你－耶和華使我安然居住。
PS|5|1|耶和華啊，求你側耳聽我的言語， 顧念我的心思！
PS|5|2|我的王，我的上帝啊，求你留心聽我呼求的聲音！ 因為我向你祈禱。
PS|5|3|耶和華啊，早晨你必聽我的聲音； 早晨我要向你陳明我的心思，並要警醒。
PS|5|4|因為你不是喜愛邪惡的上帝， 惡人不能與你同住。
PS|5|5|狂傲的人不能站在你眼前； 凡作惡的，都是你所恨惡的。
PS|5|6|說謊言的，你必滅絕； 好流人血、玩弄詭詐的，都為耶和華所憎惡。
PS|5|7|至於我，我必憑你豐盛的慈愛進入你的居所， 我要存敬畏你的心向你的聖殿下拜。
PS|5|8|耶和華啊，求你因我仇敵的緣故，憑你的公義引領我， 使你的道路在我面前正直。
PS|5|9|因為他們口中沒有誠實， 心裏充滿邪惡， 他們的喉嚨是敞開的墳墓； 他們用舌頭諂媚人。
PS|5|10|上帝啊，求你定他們的罪！ 願他們因自己的計謀跌倒； 求你因他們過犯眾多趕逐他們， 因為他們背叛了你。
PS|5|11|凡投靠你的，願他們喜樂，時常歡呼， 因為你庇護他們； 又願那愛你名的人都靠你歡欣。
PS|5|12|耶和華啊，因為你必賜福給義人， 你必用恩惠如同盾牌四面護衛他。
PS|6|1|耶和華啊，求你不要在怒中責備我， 不要在烈怒中懲罰我！
PS|6|2|耶和華啊，求你憐憫我，因為我軟弱。 耶和華啊，求你醫治我，因為我的骨頭戰抖。
PS|6|3|我的心也大大驚惶。 耶和華啊，你要等到幾時呢？
PS|6|4|耶和華啊，求你轉回搭救我， 因你的慈愛拯救我。
PS|6|5|因為死了的人不會記念你， 在陰間有誰稱謝你？
PS|6|6|我因呻吟而困乏； 我每夜流淚，使床鋪漂起， 把褥子濕透。
PS|6|7|我的眼睛因憂愁而昏花， 因敵人的緣故，我的眼目模糊不清。
PS|6|8|你們所有作惡的人，離開我吧！ 因為耶和華聽了我哀哭的聲音。
PS|6|9|耶和華聽了我的懇求， 耶和華必接納我的禱告。
PS|6|10|我所有的仇敵都必羞愧，大大驚惶； 轉眼之間，他們要羞愧撤退。
PS|7|1|耶和華－我的上帝啊，我投靠你！ 求你救我脫離所有追趕我的人，搭救我出來！
PS|7|2|免得他們像獅子撕裂我， 甚至撕碎，無人搭救。
PS|7|3|耶和華－我的上帝啊，我若行了這事， 若有罪孽在我手裏，
PS|7|4|我若以惡回報我的朋友， 連那無故與我為敵的，我也救了他 ，
PS|7|5|就任憑仇敵追趕我，直到追上， 把我的性命踏在地上， 使我的榮耀歸於灰塵。（細拉）
PS|7|6|耶和華啊，求你在怒中起來， 挺身而立，抵擋我敵人的烈怒！ 求你為我興起！你已經發令施行審判。
PS|7|7|願萬民聚集環繞你！ 願你居高位統治他們！
PS|7|8|耶和華向萬民施行審判； 耶和華啊，求你按我的公義 和我心中的純正判斷我。
PS|7|9|願惡人的惡斷絕！ 願你堅立義人！ 因為公義的上帝察驗人的心腸肺腑。
PS|7|10|上帝是我的盾牌， 他拯救心裏正直的人。
PS|7|11|上帝是公義的審判者， 又是天天向惡人發怒的上帝。
PS|7|12|若有人不回頭，他的刀必磨快， 弓必上弦，預備妥當。
PS|7|13|他也預備了致死的兵器， 他所射的是火箭。
PS|7|14|看哪，惡人懷邪惡， 養毒害，生虛假。
PS|7|15|他掘了坑，挖得太深， 竟掉在自己所挖的陷阱裏。
PS|7|16|他的毒害必回到自己頭上， 他的殘暴必落到自己的腦袋上。
PS|7|17|我要照著耶和華的公義稱謝他， 要歌頌耶和華至高者的名。
PS|8|1|耶和華－我們的主啊， 你的名在全地何其美！ 你將你的榮耀彰顯於天 。
PS|8|2|你因敵人的緣故， 從孩童和吃奶的口中建立了能力， 使仇敵和報仇的閉口無言。
PS|8|3|我觀看你手指所造的天， 並你所陳設的月亮星宿。
PS|8|4|人算甚麼，你竟顧念他！ 世人算甚麼，你竟眷顧他！
PS|8|5|你使他比上帝 微小一點， 賜他榮耀尊貴為冠冕。
PS|8|6|你派他管理你手所造的， 使萬物，就是一切的牛羊、 田野的牲畜、空中的鳥、海裏的魚， 凡游在水裏的，都服在他的腳下。
PS|8|7|
PS|8|8|
PS|8|9|耶和華－我們的主啊， 你的名在全地何其美！
PS|9|1|我要一心稱謝耶和華， 傳揚你一切奇妙的作為。
PS|9|2|我要因你歡喜快樂； 至高者啊，我要歌頌你的名！
PS|9|3|我的仇敵回轉撤退的時候， 他們在你面前跌倒滅亡。
PS|9|4|因你已經為我伸冤，為我辯護； 你坐在寶座上，按公義審判。
PS|9|5|你曾斥責列國，滅絕惡人； 你曾塗去他們的名，直到永永遠遠。
PS|9|6|仇敵到了盡頭； 他們遭毀壞，直到永遠。 你拆毀他們的城鎮， 連他們的名字 也都消滅！
PS|9|7|惟耶和華坐在王位上，直到永遠； 他已經為審判擺設寶座。
PS|9|8|他要按公義審判世界， 按正直判斷萬民。
PS|9|9|耶和華要作受欺壓者的庇護所， 在患難時的庇護所。
PS|9|10|耶和華啊，認識你名的人要倚靠你， 因你沒有離棄尋求你的人。
PS|9|11|應當歌頌居於 錫安 的耶和華， 將他所做的傳揚在萬民中。
PS|9|12|那位追討流人血的， 他記念受屈的人， 不忘記困苦人的哀求。
PS|9|13|耶和華啊，求你憐憫我！ 你是從死門把我提升起來的， 求你看那恨我的人所加給我的苦難，
PS|9|14|好讓我述說你一切的美德。 我要在 錫安 的城門因你的救恩歡樂。
PS|9|15|外邦人陷在自己所掘的坑中， 他們的腳被自己暗設的網羅纏住了。
PS|9|16|耶和華已將自己顯明，他已施行審判； 惡人被自己手所做的纏住了 。（細拉）
PS|9|17|惡人，就是忘記上帝的外邦人， 都必歸到陰間。
PS|9|18|貧窮人必不永久被忘， 困苦人的指望必不永遠落空。
PS|9|19|耶和華啊，求你興起，不容世人得勝！ 願外邦人在你面前受審判！
PS|9|20|耶和華啊，求你使他們恐懼， 願外邦人知道自己不過是人。（細拉）
PS|10|1|耶和華啊，你為甚麼站在遠處？ 在患難的時候為甚麼隱藏？
PS|10|2|惡人驕橫地追逼困苦人； 願他們陷在自己所設的計謀裏。
PS|10|3|因為惡人以自己的心願自誇， 貪財的背棄耶和華，並且輕慢他 。
PS|10|4|惡人面帶驕傲，不尋找耶和華； 他的思想中全無上帝。
PS|10|5|他的路時常亨通， 你的審判不在他眼裏。 至於他所有的敵人，他都向他們發怒氣。
PS|10|6|他心裏說：「我必不動搖， 世世代代不遭災難。」
PS|10|7|他滿口咒罵、詭詐、欺壓， 舌底盡是毒害、奸惡。
PS|10|8|他在村莊埋伏等候， 在隱密處殺害無辜的人， 他的眼睛窺探無倚無靠的人。
PS|10|9|他埋伏在暗地，如獅子蹲在洞中。 他埋伏，要俘擄困苦人； 他拉網，就把困苦人擄去。
PS|10|10|他屈身蹲伏， 無倚無靠的人就倒在他的暴力之下。
PS|10|11|他心裏說：「上帝竟忘記了， 上帝轉臉永不觀看。」
PS|10|12|耶和華啊，求你興起！ 上帝啊，求你舉手！ 不要忘記困苦人！
PS|10|13|惡人為何輕慢上帝， 心裏說「你必不追究」？
PS|10|14|你已經察看， 顧念人的憂患和愁苦， 放在你的手中。 無倚無靠的人把自己交託給你， 你向來是幫助孤兒的。
PS|10|15|求你打斷惡人的膀臂， 至於壞人，求你追究他的惡，直到淨盡。
PS|10|16|耶和華永永遠遠為王， 外邦人從他的地已經滅絕了。
PS|10|17|耶和華啊，困苦人的心願你早已聽見； 你必堅固他們的心，也必側耳聽他們的祈求，
PS|10|18|為要給孤兒和受欺壓的人伸冤， 使世上的人不再威嚇他們。
PS|11|1|我投靠耶和華； 你們怎麼對我說：「你當像鳥逃到你們的山去；
PS|11|2|看哪，惡人彎弓，把箭搭在弦上， 要在暗中射那心裏正直的人。
PS|11|3|根基若毀壞， 義人還能做甚麼呢？」
PS|11|4|耶和華在他的聖殿裏， 耶和華在天上的寶座上； 他的眼睛察看， 他的眼目 察驗世人。
PS|11|5|耶和華考驗義人； 惟有惡人和喜愛暴力的人，他心裏恨惡。
PS|11|6|他要向惡人密佈羅網， 烈火、硫磺、熱風作他們杯中的份。
PS|11|7|因為耶和華是公義的，他喜愛義行， 正直人必得見他的面。
PS|12|1|耶和華啊，求你幫助，因虔誠人斷絕了， 世人中間忠信的人消失了。
PS|12|2|人人向鄰舍說謊； 他們說話嘴唇油滑，心口不一。
PS|12|3|願耶和華剪除一切油滑的嘴唇， 誇大的舌頭。
PS|12|4|他們說：「我們必能以舌頭取勝， 我們的嘴唇是自己的， 誰能作我們的主呢？」
PS|12|5|耶和華說：「因為困苦人的冤屈 和貧窮人的嘆息， 我現在要起來， 把他安置在他所切慕的穩妥之地。」
PS|12|6|耶和華的言語是純淨的言語， 如同銀子在泥做的爐中煉過七次。
PS|12|7|耶和華啊，你必保護他們， 你必保佑他們永遠脫離這世代的人。
PS|12|8|卑鄙的人在世人中高升時， 就有惡人四處橫行。
PS|13|1|耶和華啊，你忘記我要到幾時呢？要到永遠嗎？ 你轉臉不顧我要到幾時呢？
PS|13|2|我心裏籌算，終日愁苦，要到幾時呢？ 我的仇敵升高壓制我，要到幾時呢？
PS|13|3|耶和華－我的上帝啊，求你看顧我，應允我！ 求你使我眼目明亮，免得我沉睡至死；
PS|13|4|免得我的仇敵說「我勝了他」； 免得我的敵人在我動搖的時候喜樂。
PS|13|5|但我倚靠你的慈愛， 我的心因你的救恩快樂。
PS|13|6|我要向耶和華歌唱， 因他厚厚地恩待我。
PS|14|1|愚頑人心裏說：「沒有上帝。」 他們都敗壞，行了可憎惡的事， 沒有一個人行善。
PS|14|2|耶和華從天上垂看世人， 要看有明白的沒有， 有尋求上帝的沒有。
PS|14|3|他們都偏離正路，一同變為污穢， 沒有行善的， 連一個也沒有。
PS|14|4|作惡的都沒有知識嗎？ 他們吞吃我的百姓如同吃飯一樣， 並不求告耶和華。
PS|14|5|他們在那裏大大害怕， 因為上帝在義人的族類中。
PS|14|6|你們叫困苦人的籌算變為羞辱， 然而耶和華是他的避難所。
PS|14|7|但願 以色列 的救恩出自 錫安 。 當耶和華救回他被擄子民的時候， 雅各 要快樂， 以色列 要歡喜。
PS|15|1|耶和華啊，誰能寄居你的帳幕？ 誰能居住你的聖山？
PS|15|2|就是行為正直、做事公義、 心裏說實話的人。
PS|15|3|他不以舌頭讒害人， 不惡待朋友， 也不隨夥毀謗鄰舍。
PS|15|4|他眼中藐視匪類， 卻尊重那敬畏耶和華的人。 他發了誓，雖然自己吃虧也不更改。
PS|15|5|他不放債取利， 不受賄賂以害無辜。 做這些事的人必永不動搖。
PS|16|1|上帝啊，求你保佑我， 因為我投靠你。
PS|16|2|我 曾對耶和華說：「你是我的主， 我的福氣惟獨從你而來。」
PS|16|3|論到世上的聖民，他們是尊貴的人， 是我最喜悅的。
PS|16|4|追逐 別神的， 他們的愁苦必增加； 他們所澆奠的血我不獻上， 我嘴唇也不提別神的名號。
PS|16|5|耶和華是我的產業，是我杯中的福分； 我所得的，你為我持守。
PS|16|6|用繩量給我的地界，坐落在佳美之處； 我的產業實在美好。
PS|16|7|我要稱頌那指引我的耶和華， 在夜間我的心腸也指教我。
PS|16|8|我讓耶和華常在我面前， 因他在我右邊，我就不致動搖。
PS|16|9|因此，我的心歡喜，我的靈 快樂； 我的肉身也要安然居住。
PS|16|10|因為你必不將我的靈魂 撇在陰間， 也不讓你的聖者見地府 。
PS|16|11|你必將生命的道路指示我。 在你面前有滿足的喜樂， 在你右手中有永遠的福樂。
PS|17|1|耶和華啊，求你垂聽公義的呼聲， 留心聽我的呼求！ 求你側耳聽我這沒有詭詐的嘴唇的祈禱！
PS|17|2|願判我公正的話從你面前發出， 願你的眼睛察看正直。
PS|17|3|你已經考驗我的心， 你在夜間鑒察我。 你熬煉我，卻找不到錯失， 我立志叫我口中沒有過失。
PS|17|4|論到人的行為，我謹守你嘴唇的言語， 不走殘暴人的道路。
PS|17|5|我的腳緊緊跟隨你的腳蹤， 我的兩腳未曾滑跌。
PS|17|6|上帝啊，我求告你，因為你必應允我； 求你向我側耳，聽我的言語。
PS|17|7|求你顯出你奇妙的慈愛， 你用右手拯救投靠你的人，脫離那起來攻擊他們的人。
PS|17|8|求你保護我，如同保護眼中的瞳人， 把我隱藏在你翅膀的蔭下，
PS|17|9|使我脫離欺壓我的惡人， 脫離那圍困我要害我命的仇敵。
PS|17|10|他們的心被油脂包裹， 用口說驕傲的話。
PS|17|11|他們追逼我 ，現在他們圍困了我們， 瞪著眼，要把我們推倒在地。
PS|17|12|他像獅子要貪吃獵物， 又像少壯獅子蹲伏在暗處。
PS|17|13|耶和華啊，求你興起，前去迎敵，把他打倒！ 求你用你的刀救我的命脫離惡人。
PS|17|14|耶和華啊，求你用手救我脫離世人， 脫離那只在今生有福分的世人！ 你以財寶充滿他們的肚腹， 他們因有兒女就滿足， 將其餘的財物留給他們的孩子。
PS|17|15|至於我，我必因公正得見你的面； 我醒了的時候，你的形像使我滿足。
PS|18|1|耶和華我的力量啊，我愛你！
PS|18|2|耶和華是我的巖石、我的山寨、我的救主、 我的上帝、我的磐石、我所投靠的。 他是我的盾牌， 是拯救我的角，是我的碉堡。
PS|18|3|我要求告當讚美的耶和華， 我必從仇敵手中被救出來。
PS|18|4|死亡的繩索勒住我， 毀滅的急流驚嚇我，
PS|18|5|陰間的繩索纏繞我， 死亡的圈套臨到我。
PS|18|6|我在急難中求告耶和華， 向我的上帝呼求。 他從殿中聽了我的聲音， 我在他面前的呼求必進入他耳中。
PS|18|7|那時，因他發怒地就震動戰抖， 山的根基也震動挪移。
PS|18|8|他的鼻孔冒煙上騰， 他的口發火焚燒，連煤炭也燒著了。
PS|18|9|他使天垂下，親自降臨， 黑雲在他腳下。
PS|18|10|他乘坐基路伯飛行， 藉著風的翅膀快飛，
PS|18|11|以黑暗為藏身之處， 以水的黑暗、天空的密雲作四圍的行宮。
PS|18|12|因他發出光輝， 冰雹和火炭穿透密雲。
PS|18|13|耶和華在天上打雷， 至高者發出聲音，就有冰雹和火炭 。
PS|18|14|他射出箭來，使仇敵四散； 發出連串的閃電，擊潰他們。
PS|18|15|耶和華啊，你的斥責一發， 你鼻孔的氣一出， 海底就顯現， 大地的根基也暴露。
PS|18|16|他從高天伸手抓住我， 把我從大水中拉上來。
PS|18|17|他救我脫離強敵和那些恨我的人， 因為他們比我強盛。
PS|18|18|我遭遇災難的日子，他們來攻擊我； 但耶和華是我的倚靠。
PS|18|19|他領我到寬闊之處， 他救拔我，因他喜愛我。
PS|18|20|耶和華必按我的公義報答我， 按我手中的清潔賞賜我。
PS|18|21|因為我遵守耶和華的道， 未曾作惡離開我的上帝。
PS|18|22|他的一切典章常在我面前， 他的律例我也未曾丟棄。
PS|18|23|我在他面前作了完全人， 我也保護自己遠離罪孽。
PS|18|24|所以耶和華按我的公義， 在他眼前按我手中的清潔賞賜我。
PS|18|25|慈愛的人，你以慈愛待他； 完全的人，你以完善待他。
PS|18|26|清潔的人，你以清潔待他； 歪曲的人，你以彎曲待他。
PS|18|27|困苦的百姓，你必拯救； 高傲的眼目，你使他降卑。
PS|18|28|你必點亮我的燈； 耶和華－我的上帝必照明我的黑暗。
PS|18|29|我藉著你衝入敵軍， 藉著我的上帝跳過城牆。
PS|18|30|至於上帝，他的道是完全的； 耶和華的話是純淨的。 凡投靠他的，他就作他們的盾牌。
PS|18|31|除了耶和華，誰是上帝呢？ 除了我們的上帝，誰是磐石呢？
PS|18|32|惟有那以力量束我的腰、 使我行為完全的，他是上帝。
PS|18|33|他使我的腳快如母鹿， 使我站穩在高處。
PS|18|34|他教導我的手能爭戰， 我的膀臂能開銅造的弓。
PS|18|35|你賜救恩給我作盾牌， 你的右手扶持我， 你的庇護 使我為大。
PS|18|36|你使我腳步寬闊， 我的腳踝未曾滑跌。
PS|18|37|我要追趕我的仇敵，且要追上他們； 若不將他們滅絕，我總不歸回。
PS|18|38|我要打傷他們，使他們站不起來； 他們必倒在我的腳下。
PS|18|39|你曾以力量束我的腰，使我能爭戰； 也曾使那起來攻擊我的，都服在我以下。
PS|18|40|你又使我的仇敵在我面前轉身逃跑， 使我剪除那恨我的人。
PS|18|41|他們呼求，卻無人拯救； 就是呼求耶和華，他也不應允。
PS|18|42|我搗碎他們，如同風前的灰塵； 傾倒 他們，如同街上的泥土。
PS|18|43|你救我脫離百姓的紛爭， 立我作列國的元首； 我素不認識的百姓必事奉我。
PS|18|44|他們一聽見我的名聲就必順從我， 外邦人要投降我。
PS|18|45|外邦人要喪膽， 戰戰兢兢地出營寨。
PS|18|46|耶和華永遠活著。 願我的磐石被稱頌， 願救我的上帝受尊崇。
PS|18|47|這位上帝為我伸冤， 使萬民服在我以下。
PS|18|48|他拯救我脫離仇敵， 又把我舉起，高過那些起來攻擊我的人， 救我脫離殘暴的人。
PS|18|49|耶和華啊，因此我要在外邦中稱謝你， 歌頌你的名。
PS|18|50|耶和華賜極大的救恩給他所立的王， 施慈愛給他的受膏者， 就是給 大衛 和他的後裔，直到永遠。
PS|19|1|諸天述說上帝的榮耀， 穹蒼傳揚他手的作為。
PS|19|2|這日到那日發出言語， 這夜到那夜傳出知識。
PS|19|3|無言無語， 也無聲音可聽。
PS|19|4|它們的聲浪 傳遍天下， 它們的言語傳到地極。 上帝在其中為太陽安設帳幕，
PS|19|5|太陽如同新郎步出洞房， 又如勇士歡然奔路。
PS|19|6|它從天這邊出來，繞到天那邊， 沒有一物可隱藏得不到它的熱氣。
PS|19|7|耶和華的律法全備，使人甦醒； 耶和華的法度確定，使愚蒙人有智慧。
PS|19|8|耶和華的訓詞正直，使人心快活； 耶和華的命令清潔，使人眼目明亮。
PS|19|9|耶和華的典章真實，全然公義， 敬畏耶和華是純潔的，存到永遠，
PS|19|10|比金子可羨慕，比極多的純金可羨慕； 比蜜甘甜，比蜂房下滴的蜜甘甜。
PS|19|11|因此你的僕人受警戒， 遵守這些有極大的賞賜。
PS|19|12|誰能察覺自己的錯失呢？ 求你赦免我隱藏的過犯。
PS|19|13|求你攔阻僕人不犯任意妄為的罪， 不容這罪轄制我， 我就完全，免犯大罪。
PS|19|14|耶和華－我的磐石，我的救贖主啊， 願我口中的言語，心裏的意念在你面前蒙悅納。
PS|20|1|願耶和華在你患難的日子應允你， 願 雅各 的上帝的名保護你。
PS|20|2|願他從聖所救助你， 從 錫安 堅固你，
PS|20|3|記念你的一切祭物， 悅納你的燔祭，（細拉）
PS|20|4|將你心所願的賜給你， 成就你的一切籌算。
PS|20|5|我們要因你的救恩誇勝， 要奉我們上帝的名豎立旌旗。 願耶和華成就你一切所求的！
PS|20|6|現在我知道耶和華必救護他的受膏者， 從他神聖的天上應允他， 用右手的能力救護他。
PS|20|7|有人靠車，有人靠馬， 但我們要提耶和華－我們上帝的名。
PS|20|8|他們都屈身仆倒， 我們卻起來，堅立不移。
PS|20|9|耶和華啊，求你拯救； 我們呼求的時候，願王應允我們！
PS|21|1|耶和華啊，王必因你的能力歡喜； 因你的救恩，他的快樂何其大！
PS|21|2|他心裏所願的，你已經賜給他； 他嘴唇所求的，你未嘗不應允。（細拉）
PS|21|3|你以美善的福氣迎接他， 把純金的冠冕戴在他頭上。
PS|21|4|他向你祈求長壽，你就賜給他， 就是日子長久，直到永遠。
PS|21|5|他因你的救恩大有榮耀， 你將尊榮威嚴加在他身上。
PS|21|6|你使他有洪福，直到永遠， 又使他在你面前歡喜快樂。
PS|21|7|王倚靠耶和華， 因至高者的慈愛，王必不動搖。
PS|21|8|你的手要搜出所有的仇敵， 你的右手要搜出那些恨你的人。
PS|21|9|你的臉出現的時候，要使他們如在炎熱的火爐中。 耶和華要在他的震怒中吞滅他們， 那火要把他們燒盡。
PS|21|10|你必從世上滅絕他們的幼苗， 從人間滅絕他們的後裔。
PS|21|11|因為他們有意加害於你； 他們想出計謀，卻不能做成。
PS|21|12|你必使他們轉身逃跑， 向著他們的臉搭箭在弦。
PS|21|13|耶和華啊，願你因自己的能力顯為至高！ 這樣，我們就唱詩，歌頌你的大能。
PS|22|1|我的上帝，我的上帝，為甚麼離棄我？ 為甚麼遠離不救我，不聽我的呻吟？
PS|22|2|我的上帝啊，我白日呼求，你不應允； 夜間呼求，也不得安寧。
PS|22|3|但你是神聖的， 用 以色列 的讚美為寶座。
PS|22|4|我們的祖宗倚靠你； 他們倚靠你，你解救他們。
PS|22|5|他們哀求你，就蒙解救； 他們倚靠你，就不羞愧。
PS|22|6|但我是蟲，不是人， 被眾人羞辱，被百姓藐視。
PS|22|7|凡看見我的都嗤笑我； 他們撇嘴搖頭：
PS|22|8|「他把自己交託給耶和華，讓耶和華救他吧！ 耶和華既喜愛他，可以搭救他吧！」
PS|22|9|但你是叫我出母腹的， 我在母懷裏，你就使我有倚靠的心。
PS|22|10|我自出母胎就交在你手裏， 自我出母腹，你就是我的上帝。
PS|22|11|求你不要遠離我！ 因為災難臨頭，無人幫助。
PS|22|12|許多公牛環繞我， 巴珊 大力的公牛四面圍困我。
PS|22|13|牠們向我張口， 好像獵食吼叫的獅子。
PS|22|14|我如水被倒出， 我的骨頭都脫了節， 我的心如蠟，在我裏面熔化。
PS|22|15|我的精力枯乾，如同瓦片， 我的舌頭緊貼上顎。 你將我安置在死灰中。
PS|22|16|犬類圍著我，惡黨環繞我； 他們扎了我的手、我的腳。
PS|22|17|我數遍我的骨頭； 他們瞪著眼看我。
PS|22|18|他們分我的外衣， 為我的內衣抽籤。
PS|22|19|耶和華啊，求你不要遠離我！ 我的救主啊，求你快來幫助我！
PS|22|20|求你救我的性命脫離刀劍， 使我僅有的 脫離犬類，
PS|22|21|求你救我脫離獅子的口； 你已經應允我，使我脫離野牛的角。
PS|22|22|我要將你的名傳給我的弟兄， 在會眾中我要讚美你。
PS|22|23|敬畏耶和華的人哪，要讚美他！ 雅各 的後裔啊，要榮耀他！ 以色列 的後裔啊，要懼怕他！
PS|22|24|因為他沒有藐視、憎惡受苦的人， 也沒有轉臉不顧他們； 那受苦之人呼求的時候，他就垂聽。
PS|22|25|我在大會中讚美你的話是從你而來， 我要在敬畏耶和華的人面前還我的願。
PS|22|26|願困苦的人吃得飽足， 願尋求耶和華的人讚美他。 願你們的心永遠活著！
PS|22|27|地的四極都要想念耶和華，並且歸順他， 列國的萬族都要在你面前敬拜。
PS|22|28|因為國度屬於耶和華， 他是管理列國的。
PS|22|29|地上富足的人都必吃喝而敬拜， 凡下到塵土中不能存活自己性命的人， 都要在他面前下拜 ；
PS|22|30|必有後裔事奉他， 主所做的事必傳給後代。
PS|22|31|他們必來傳他的公義給尚未出生的子民， 這是他的作為。
PS|23|1|耶和華是我的牧者， 我必不致缺乏。
PS|23|2|他使我躺臥在青草地上， 領我在可安歇的水邊。
PS|23|3|他使我的靈魂甦醒 ， 為自己的名引導我走義路。
PS|23|4|我雖然行過死蔭的幽谷， 也不怕遭害， 因為你與我同在； 你的杖、你的竿，都安慰我。
PS|23|5|在我敵人面前，你為我擺設筵席； 你用油膏了我的頭，使我的福杯滿溢。
PS|23|6|我一生一世必有恩惠慈愛隨著我； 我且要住在 耶和華的殿中，直到永遠。
PS|24|1|地和其中所充滿的， 世界和住在其中的，都屬耶和華。
PS|24|2|他把地建立在海上， 安定在江河之上。
PS|24|3|誰能登耶和華的山？ 誰能站在他的聖所？
PS|24|4|就是手潔心清，意念不向虛妄， 起誓不懷詭詐的人。
PS|24|5|他必蒙耶和華賜福， 又蒙救他的上帝使他成義。
PS|24|6|這是尋求耶和華的族類， 是尋求你面的 雅各 。（細拉）
PS|24|7|眾城門哪，要抬起頭來！ 永久的門戶啊，你們要被舉起！ 榮耀的王將要進來！
PS|24|8|這榮耀的王是誰呢？ 就是有力有能的耶和華， 在戰場上大有能力的耶和華！
PS|24|9|眾城門哪，要抬起頭來！ 永久的門戶啊，你們要高舉！ 榮耀的王將要進來！
PS|24|10|這榮耀的王是誰呢？ 萬軍之耶和華是榮耀的王！（細拉）
PS|25|1|耶和華啊，我的心仰望你。
PS|25|2|我的上帝啊，我素來倚靠你； 求你不要叫我羞愧， 不要叫我的仇敵向我誇勝。
PS|25|3|凡等候你的必不羞愧， 惟有那無故行奸詐的必要羞愧。
PS|25|4|耶和華啊，求你將你的道指示我， 將你的路指教我！
PS|25|5|求你指教我，引導我進入你的真理， 因為你是救我的上帝。 我整日等候你。
PS|25|6|耶和華啊，求你記念你的憐憫和慈愛， 因為這是亙古以來所常有的。
PS|25|7|求你不要記得我幼年的罪愆和我的過犯； 耶和華啊，求你因你的良善，按你的慈愛記念我。
PS|25|8|耶和華是良善正直的， 因此，他必教導罪人走正路。
PS|25|9|他要按公平引領謙卑人， 將他的道指教他們。
PS|25|10|凡遵守他的約和他法度的人， 耶和華都以慈愛信實待他。
PS|25|11|耶和華啊，求你因你名的緣故赦免我的罪， 因我的罪重大。
PS|25|12|誰敬畏耶和華， 耶和華必教導他當選擇的道路。
PS|25|13|他要安然居住， 他的後裔必承受土地。
PS|25|14|耶和華與敬畏他的人親密， 他要將自己的約指示他們。
PS|25|15|我的眼目時常仰望耶和華， 因他必將我的腳從網裏拉出來。
PS|25|16|求你轉向我，憐憫我， 因我孤獨困苦。
PS|25|17|我心裏愁苦甚多， 求你救我脫離我的禍患。
PS|25|18|求你看顧我的困苦、我的艱難， 赦免我一切的罪。
PS|25|19|求你察看我的仇敵， 因為他們人數眾多，並且痛恨我。
PS|25|20|求你保護我的性命，搭救我， 使我不致羞愧，因為我投靠你。
PS|25|21|願純全、正直保護我， 因為我等候你。
PS|25|22|上帝啊，求你救贖 以色列 脫離他一切的愁苦。
PS|26|1|耶和華啊，求你為我伸冤， 因我向來行事純正； 我倚靠耶和華，必不動搖。
PS|26|2|耶和華啊，求你察看我，考驗我， 熬煉我的肺腑心腸。
PS|26|3|因為你的慈愛常在我眼前， 我也按你的真理而行。
PS|26|4|我未曾與虛妄的人同坐， 也不與偽善的人來往。
PS|26|5|我痛恨惡人的集會， 必不與惡人同坐。
PS|26|6|耶和華啊，我要洗手表明無辜， 才環繞你的祭壇；
PS|26|7|我好發出稱謝的聲音， 述說你一切奇妙的作為。
PS|26|8|耶和華啊，我喜愛你所住的殿 和你顯榮耀的居所。
PS|26|9|不要把我的性命和罪人一同除掉， 不要把我的生命和好流人血的一同除掉。
PS|26|10|他們的手中有奸惡， 他們的右手滿有賄賂。
PS|26|11|至於我，卻要行事純正； 求你救贖我，憐憫我！
PS|26|12|我的腳站在平坦的地方， 在聚會中我要稱頌耶和華！
PS|27|1|耶和華是我的亮光，是我的拯救， 我還怕誰呢？ 耶和華是我生命的保障， 我還懼誰呢？
PS|27|2|那作惡的就是我的仇敵， 前來吃我肉的時候就絆跌仆倒。
PS|27|3|雖有軍隊安營攻擊我，我的心也不害怕； 雖然興起戰爭攻擊我，我仍舊安穩。
PS|27|4|有一件事，我曾求耶和華，我仍要尋求， 就是一生一世住在耶和華的殿中， 瞻仰他的榮美，在他的殿宇裏求問。
PS|27|5|因為我遭遇患難，他必將我隱藏在他的帳棚裏， 把我藏在他帳幕的隱密處， 將我高舉在磐石上。
PS|27|6|現在我得以昂首，高過四面的仇敵。 我要在他的帳幕裏歡然獻祭， 我要唱詩歌頌耶和華。
PS|27|7|耶和華啊，我呼求的時候，求你垂聽我的聲音； 求你憐憫我，應允我。
PS|27|8|你說：「你們當尋求我的面。」 那時我的心向你說： 「耶和華啊，你的面我正要尋求。」
PS|27|9|求你不要轉臉不顧我， 不要發怒趕逐你的僕人， 你向來是幫助我的。 救我的上帝啊，不要離開我， 也不要撇棄我。
PS|27|10|即使我的父母撇棄我， 耶和華終必收留我。
PS|27|11|耶和華啊，求你將你的道指教我， 因我仇敵的緣故引導我走平坦的路。
PS|27|12|求你不要把我交給敵人，遂其所願； 因為妄作見證的和口吐凶言的都起來攻擊我。
PS|27|13|我深信在活人之地 必得見耶和華的恩惠。
PS|27|14|要等候耶和華， 當壯膽，堅固你的心， 要等候耶和華！
PS|28|1|耶和華啊，我要求告你！ 我的磐石啊，求你不要向我緘默！ 倘若你向我閉口， 我就如下入地府的人一樣。
PS|28|2|我呼求你，向你至聖所舉手的時候， 求你垂聽我懇求的聲音！
PS|28|3|不要把我和壞人並作惡的一同除掉； 他們跟鄰舍說平安，心裏卻是奸惡。
PS|28|4|求你按著他們所做的， 按他們的惡行對待他們； 求你照著他們手所做的對待他們， 將他們應得的報應加給他們。
PS|28|5|他們既然不尊重耶和華的作為， 也不尊重他手所做的， 耶和華就必毀壞他們，不建立他們。
PS|28|6|耶和華是應當稱頌的， 因為他聽了我懇求的聲音。
PS|28|7|耶和華是我的力量，是我的盾牌， 我心裏倚靠他就得幫助。 我心中歡樂， 我要用詩歌稱謝他。
PS|28|8|耶和華是他百姓的力量， 又是他受膏者得救的保障。
PS|28|9|求你拯救你的百姓，賜福給你的產業； 求你牧養他們，扶持他們，直到永遠。
PS|29|1|上帝的子民 哪，你們要將榮耀、能力歸給耶和華， 都歸給耶和華！
PS|29|2|要將耶和華的名的榮耀歸給他， 要敬拜神聖榮耀的耶和華 。
PS|29|3|耶和華的聲音在眾水上， 榮耀的上帝打雷； 耶和華打雷在大水之上。
PS|29|4|耶和華的聲音大有能力， 耶和華的聲音滿有威嚴。
PS|29|5|耶和華的聲音震碎香柏樹， 耶和華震碎 黎巴嫩 的香柏樹。
PS|29|6|他使 黎巴嫩 跳躍如牛犢， 使 西連 跳躍如野牛犢。
PS|29|7|耶和華的聲音使火焰分岔。
PS|29|8|耶和華的聲音震動曠野， 耶和華震動 加低斯 的曠野。
PS|29|9|耶和華的聲音驚動母鹿落胎， 樹林也脫落淨光。 凡在他殿中的，都述說他的榮耀。
PS|29|10|耶和華坐在洪水之上為王； 耶和華坐著為王，直到永遠。
PS|29|11|耶和華必賜力量給他的百姓， 耶和華必賜平安的福給他的百姓。
PS|30|1|耶和華啊，我要尊崇你， 因為你救了我，不讓仇敵向我誇耀。
PS|30|2|耶和華－我的上帝啊， 我呼求你，你醫治了我。
PS|30|3|耶和華啊，你救我的性命脫離陰間， 使我存活，不至於下入地府。
PS|30|4|耶和華的聖民哪，你們要歌頌他， 要頌揚他神聖的名字 。
PS|30|5|因為，他的怒氣不過是轉眼之間； 他的恩典乃是一生之久。 一宿雖然有哭泣， 早晨便必歡呼。
PS|30|6|至於我，我凡事順利，就說： 「我永不動搖。」
PS|30|7|耶和華啊，你曾施恩，使我穩固如山； 你轉臉不顧，我就驚惶。
PS|30|8|耶和華啊，我曾求告你； 我向耶和華懇求：
PS|30|9|「我被害流血，下到地府，有何益處呢？ 塵土豈能稱謝你、傳揚你的信實嗎？
PS|30|10|耶和華啊，求你應允我，憐憫我！ 耶和華啊，求你幫助我！」
PS|30|11|你將我的哀哭變為跳舞， 脫去我的麻衣，為我披上喜樂，
PS|30|12|使我的靈 歌頌你，不致緘默。 耶和華－我的上帝啊，我要稱謝你，直到永遠！
PS|31|1|耶和華啊，我投靠你， 求你使我永不羞愧， 憑你的公義搭救我！
PS|31|2|求你側耳聽我， 快快救我！ 求你作我堅固的磐石， 拯救我的保障！
PS|31|3|你真是我的巖石、我的山寨， 求你為你名的緣故引導我，指教我。
PS|31|4|求你救我脫離人為我暗設的網羅， 因為你是我的保障。
PS|31|5|我將我的靈交在你手裏； 耶和華─信實的上帝啊，你救贖了我。
PS|31|6|我 恨惡那信奉虛無神明 的人； 我卻倚靠耶和華。
PS|31|7|我要因你的慈愛歡喜快樂， 因為你見過我的困苦， 知道我心中的艱難。
PS|31|8|你未曾把我交在仇敵手裏， 你使我的腳站在寬闊的地方。
PS|31|9|耶和華啊，求你憐憫我， 因為我在急難之中； 我的眼睛因憂愁而昏花， 我的身心也已耗盡。
PS|31|10|我的生命為愁苦所消耗， 我的年歲為嘆息所荒廢； 我的力量因我的罪孽 衰敗， 我的骨頭也枯乾。
PS|31|11|我因所有的敵人成了羞辱， 在我鄰舍跟前更加羞辱； 那認識我的都懼怕我， 在街上看見我的都躲避我。
PS|31|12|我被遺忘，如同死人，無人記念； 我好像破碎的器皿。
PS|31|13|我聽見許多人的毀謗， 四圍盡是驚嚇； 他們一同商議攻擊我， 圖謀害我的性命。
PS|31|14|耶和華啊，我仍要倚靠你； 我說：「你是我的上帝。」
PS|31|15|我終生的事在你手中， 求你救我脫離仇敵的手和那些迫害我的人。
PS|31|16|求你使你的臉向僕人發光， 憑你的慈愛拯救我。
PS|31|17|耶和華啊，求你叫我不致羞愧， 因為我曾呼求你； 求你使惡人羞愧， 使他們在陰間緘默無聲。
PS|31|18|那撒謊的人逞驕傲輕慢， 出狂妄的話攻擊義人， 願他的嘴啞而無言。
PS|31|19|在世人眼前， 你為敬畏你的人所積存的， 為投靠你的人所施行的， 是何等大的恩惠啊！
PS|31|20|你必將他們藏在你面前的隱密處， 免得遭人暗算； 你要隱藏他們在棚子裏， 免受口舌的爭鬧。
PS|31|21|耶和華是應當稱頌的， 因為我在圍城裏，他向我施展奇妙的慈愛。
PS|31|22|至於我，我曾驚惶地說： 「我從你眼前被隔絕。」 然而，我呼求你的時候， 你仍聽我懇求的聲音。
PS|31|23|耶和華的聖民哪，你們都要愛他！ 耶和華保護誠實可靠的人， 卻加倍報應行事驕傲的人。
PS|31|24|凡仰望耶和華的人， 你們都要壯膽，堅固你們的心！
PS|32|1|過犯得赦免， 罪惡蒙遮蓋的人有福了！
PS|32|2|耶和華不算為有罪， 內心沒有詭詐的人有福了！
PS|32|3|我閉口不認罪的時候， 因終日呻吟而骨頭枯乾。
PS|32|4|黑夜白日，你的手壓在我身上沉重； 我的精力耗盡 ，如同夏天的乾旱。（細拉）
PS|32|5|我向你陳明我的罪， 不隱瞞我的惡。 我說：「我要向耶和華承認我的過犯」； 你就赦免我的罪惡。（細拉）
PS|32|6|為此，凡虔誠人都當趁你可尋找 的時候向你禱告； 大水氾濫的時候，必不臨到他。
PS|32|7|你是我藏身之處， 你必保佑我脫離苦難， 以得救的歡呼 四面環繞我。（細拉）
PS|32|8|我要教導你，指示你當行的路， 我要定睛在你身上勸戒你。
PS|32|9|你不可像那無知的騾馬， 須用嚼環韁繩勒住， 不然，牠就不會靠近你。
PS|32|10|惡人必多受苦楚； 惟獨倚靠耶和華的，必有慈愛四面環繞他。
PS|32|11|義人哪，你們應當靠耶和華歡喜快樂， 心裏正直的人哪，你們都當歡呼。
PS|33|1|義人哪，你們當因耶和華歡呼， 正直人理當讚美耶和華。
PS|33|2|你們要彈琴稱謝耶和華， 用十弦瑟歌頌他。
PS|33|3|應當向他唱新歌， 彈得巧妙，聲音洪亮。
PS|33|4|因為耶和華的言語正直， 他的作為盡都信實。
PS|33|5|他喜愛公義和公平， 遍地滿了耶和華的慈愛。
PS|33|6|諸天藉耶和華的話而造， 萬象藉他口中的氣而成。
PS|33|7|他聚集海水如壘， 收藏深洋在倉庫。
PS|33|8|願全地都敬畏耶和華！ 願世上的居民都懼怕他！
PS|33|9|因為他說有，就有， 命立，就立。
PS|33|10|耶和華使列國的籌算歸於無有， 使萬民的計謀全無功效。
PS|33|11|耶和華的籌算永遠立定， 他心中的計劃萬代長存。
PS|33|12|以耶和華為上帝的，那國有福了！ 耶和華揀選為自己產業的，那民有福了！
PS|33|13|耶和華從天上觀看， 看見所有的人，
PS|33|14|從他的居所察看地上每一個居民，
PS|33|15|他塑造他們的心， 洞察他們一切的作為。
PS|33|16|君王不能因兵多得勝， 勇士不能因力大得救。
PS|33|17|靠馬得救是枉然的， 馬也不能因力大救人。
PS|33|18|看哪，耶和華的眼目看顧敬畏他的人 和仰望他慈愛的人，
PS|33|19|要救他們的性命脫離死亡， 使他們在饑荒中存活。
PS|33|20|我們的心向來等候耶和華； 他是我們的幫助，是我們的盾牌。
PS|33|21|我們的心必靠他歡喜， 因為我們向來倚靠他的聖名。
PS|33|22|耶和華啊，求你照著我們所仰望你的， 向我們施行慈愛！
PS|34|1|我要時時稱頌耶和華， 讚美他的話常在我口中。
PS|34|2|我的心必因耶和華誇耀， 謙卑的人聽見就喜樂。
PS|34|3|你們要和我一同尊耶和華為大， 讓我們一同高舉他的名。
PS|34|4|我曾尋求耶和華，他就應允我， 救我脫離一切的恐懼。
PS|34|5|仰望他的人，就有光榮； 他們 的臉必不蒙羞。
PS|34|6|這困苦人呼求，耶和華就垂聽， 救他脫離一切的患難。
PS|34|7|耶和華的使者在敬畏他的人四圍安營， 要搭救他們。
PS|34|8|你們要嘗嘗主恩的滋味，便知道他是美善； 投靠他的人有福了！
PS|34|9|耶和華的聖民哪，你們當敬畏他， 因敬畏他的一無所缺。
PS|34|10|少壯獅子尚且缺食忍餓， 但尋求耶和華的甚麼好處都不缺。
PS|34|11|孩子們哪，來聽我！ 我要將敬畏耶和華的道教導你們。
PS|34|12|有誰喜愛生命， 愛慕長壽，得享美福？
PS|34|13|你要禁止舌頭不出惡言， 嘴唇不說詭詐的話。
PS|34|14|要棄惡行善， 尋求和睦，一心追求。
PS|34|15|耶和華的眼目看顧義人， 他的耳朵聽他們的呼求。
PS|34|16|耶和華向行惡的人變臉， 要從地上除滅他們的名字 。
PS|34|17|義人呼求，耶和華聽見了， 就拯救他們脫離一切患難。
PS|34|18|耶和華靠近傷心的人， 拯救心靈痛悔的人。
PS|34|19|義人多有苦難， 但耶和華救他脫離這一切，
PS|34|20|又保護他全身的骨頭， 連一根也不折斷。
PS|34|21|惡必害死惡人， 恨惡義人的，必被定罪。
PS|34|22|耶和華救贖他僕人的性命， 凡投靠他的，必不致定罪。
PS|35|1|耶和華啊，與我相爭的，求你與他們相爭！ 與我爭戰的，求你與他們爭戰！
PS|35|2|求你拿著大小盾牌， 起來幫助我；
PS|35|3|舉起槍來，抵擋那追趕我的。 求你對我說：「我是拯救你的。」
PS|35|4|願那尋索我命的，蒙羞受辱！ 願那謀害我的，退後羞愧！
PS|35|5|願他們像風前的糠秕， 有耶和華的使者趕逐他們。
PS|35|6|願他們的道路又暗又滑， 有耶和華的使者追趕他們。
PS|35|7|因他們無故為我暗設網羅， 無故挖坑，要害我的命。
PS|35|8|願災禍忽然臨到他身上！ 願他暗設的網羅纏住自己！ 願他落在其中遭災禍！
PS|35|9|我的心必靠耶和華快樂， 靠他的救恩歡喜。
PS|35|10|我全身的骨頭要說： 「耶和華啊，誰能像你 救護困苦人脫離那比他強壯的， 救護困苦貧窮人脫離那搶奪他的？」
PS|35|11|兇惡的見證人起來， 盤問我所不知道的事。
PS|35|12|他們向我以惡報善， 使我喪失兒子。
PS|35|13|至於我，他們有病的時候， 我穿麻衣，禁食，刻苦己心； 我所求的都歸到自己身上。
PS|35|14|我如此行，好像他是我的朋友，我的兄弟； 我屈身悲哀，如同哀悼自己的母親。
PS|35|15|我在患難中，他們卻歡喜，大家聚集， 我所不認識的卑賤人 聚集攻擊我， 他們不住地撕裂我。
PS|35|16|他們試探我，不斷嘲笑我 ， 向我咬牙切齒。
PS|35|17|主啊，你看著不理要到幾時呢？ 求你救我的性命脫離他們的殘害， 救我僅有的 脫離少壯獅子！
PS|35|18|我在大會中要稱謝你， 在許多百姓中要讚美你。
PS|35|19|求你不容那無理與我為仇的向我誇耀！ 不容那無故恨我的向我瞪眼！
PS|35|20|因為他們不說平安， 倒想出詭詐的言語擾害地上安靜的人。
PS|35|21|他們大大張口攻擊我，說： 「啊哈，啊哈，我們已經親眼看見了！」
PS|35|22|耶和華啊，你已經看見了，求你不要沉默！ 主啊，求你不要遠離我！
PS|35|23|我的上帝─我的主啊，求你醒來，求你奮起， 還我公正，伸明我冤！
PS|35|24|耶和華－我的上帝啊，求你按你的公義判斷我， 不容他們向我誇耀！
PS|35|25|不容他們心裏說：「啊哈，遂我們的心願了！」 不容他們說：「我們已經把他吞了！」
PS|35|26|願那喜歡我遭難的一同抱愧蒙羞！ 願那向我妄自尊大的披戴慚愧，蒙受羞辱！
PS|35|27|願那喜悅我被判為義 的歡呼快樂； 願他們常說：「當尊耶和華為大！ 耶和華喜悅他的僕人平安。」
PS|35|28|我的舌頭要論說你的公義， 要常常讚美你。
PS|36|1|過犯在惡人的心底向他說話 ， 他的眼中不怕上帝。
PS|36|2|他自誇自媚， 以致罪孽無法察覺，不被恨惡。
PS|36|3|他口中的言語盡是罪孽詭詐， 他不再有智慧，也不再行善。
PS|36|4|他在床上圖謀罪孽， 定意行不善的道，不憎惡惡事。
PS|36|5|耶和華啊，你的慈愛上及諸天， 你的信實達到穹蒼，
PS|36|6|你的公義好像高山， 你的判斷如同深淵； 耶和華啊，人民、牲畜，你都救護。
PS|36|7|上帝啊，你的慈愛何其寶貴！ 世人投靠在你翅膀的蔭下。
PS|36|8|他們必因你殿裏的豐盛得以飽足， 你也必叫他們喝你那喜樂的泉水。
PS|36|9|因為在你那裏有生命的泉源， 在你的光中，我們必得見光。
PS|36|10|願你常施慈愛給認識你的人， 常以公義待心裏正直的人。
PS|36|11|不容驕傲人的腳踐踏我， 不容兇惡人的手趕逐我。
PS|36|12|在那裏，作惡的人已經仆倒； 他們被推倒，不能再起來。
PS|37|1|不要為作惡的心懷不平， 也不要嫉妒那行不義的人。
PS|37|2|因為他們如草快被割下， 又如綠色的嫩草快要枯乾。
PS|37|3|你當倚靠耶和華而行善， 安居地上，以他的信實為糧；
PS|37|4|又當以耶和華為樂， 他就將你心裏所求的賜給你。
PS|37|5|當將你的道路交託耶和華， 並倚靠他，他就必成全。
PS|37|6|他要使你的公義如光發出， 使你的公平明如正午。
PS|37|7|你當安心倚靠耶和華，耐性等候他， 不要因那道路通達的和那惡謀成就的心懷不平。
PS|37|8|當止住怒氣，離棄憤怒； 不要心懷不平，以致作惡。
PS|37|9|因為作惡的必被剪除； 惟有等候耶和華的必承受土地。
PS|37|10|還有片時，惡人要歸於無有； 你就是細察他的住處，也不存在。
PS|37|11|但謙卑的人必承受土地， 以豐盛的平安為樂。
PS|37|12|惡人設謀要害義人， 向他咬牙。
PS|37|13|但主必笑他， 因見他受罰的日子將要來到。
PS|37|14|惡人刀已出鞘，弓已上弦， 要砍倒困苦貧窮的人， 要殺害行為正直的人。
PS|37|15|他們的刀必刺入自己的心， 他們的弓必折斷。
PS|37|16|一個義人所有的雖少， 強過許多惡人的富餘。
PS|37|17|因為惡人的膀臂必折斷； 但耶和華扶持義人。
PS|37|18|耶和華知道完全人的日子， 他們的產業要存到永遠。
PS|37|19|他們在患難的時候必不致羞愧， 在饑荒的日子必得飽足。
PS|37|20|惡人卻要滅亡。 耶和華的仇敵要像草地的華美 ； 他們要毀滅，在煙中消失 。
PS|37|21|惡人借貸卻不償還； 義人恩待人，並且施捨。
PS|37|22|蒙耶和華賜福的必承受土地； 他所詛咒的必被剪除。
PS|37|23|義人的腳步為耶和華所穩定； 他的道路，耶和華也喜愛。
PS|37|24|他雖失腳也不致全身仆倒， 因為耶和華攙扶他的手。
PS|37|25|我從前年幼，現在年老， 卻未見過義人被棄， 也未見過他的後裔求乞。
PS|37|26|他常常恩待人，借貸給人， 他的後裔也必蒙福。
PS|37|27|你當離惡行善， 就可永遠安居。
PS|37|28|因為耶和華喜愛公平， 不撇棄他的聖民， 他們永蒙保佑； 但惡人的後裔必被剪除。
PS|37|29|義人必承受土地， 永居其上。
PS|37|30|義人的口發出智慧， 他的舌頭講說公平。
PS|37|31|上帝的律法在他心裏， 他的步伐總不搖動。
PS|37|32|惡人窺探義人， 想要殺他。
PS|37|33|耶和華必不把他交在惡人手中， 當審判的時候，也不定他的罪。
PS|37|34|你當等候耶和華，遵守他的道， 他就抬舉你，使你承受土地； 你必看到惡人被剪除。
PS|37|35|我見過惡人大有勢力， 高聳如本地青翠的樹木。
PS|37|36|有人 從那裏經過，看哪，他已不存在， 我尋找他，卻尋不著了。
PS|37|37|你要細察那完全人，觀看那正直人， 因為和平的人有好結局。
PS|37|38|至於罪人，必一同滅絕， 惡人的結局必被剪除。
PS|37|39|義人得救是出於耶和華， 在患難時耶和華作他們的避難所。
PS|37|40|耶和華幫助他們，解救他們； 他解救他們脫離惡人，把他們救出來， 因為他們投靠他。
PS|38|1|耶和華啊，求你不要在怒中責備我， 不要在烈怒中懲罰我！
PS|38|2|因為你的箭射入我身， 你的手壓住我。
PS|38|3|因你的惱怒，我的肉無一完全； 因我的罪過，我的骨頭也不安寧。
PS|38|4|我的罪孽高過我的頭， 如同重擔叫我擔當不起。
PS|38|5|因我的愚昧， 我的傷發臭流膿。
PS|38|6|我疼痛，大大蜷曲， 整日哀痛。
PS|38|7|我滿腰灼熱， 我的肉無一完全。
PS|38|8|我被壓碎，身心虛弱； 因心裏痛苦，我就呻吟。
PS|38|9|主啊，我的心願都在你面前， 我的嘆息不向你隱瞞。
PS|38|10|我心顫慄，體力衰微， 眼中無光。
PS|38|11|我遭遇災病，良朋密友都袖手旁觀， 我的親戚本家也遠遠站立。
PS|38|12|那尋索我命的設下羅網， 那想要害我的口出惡言， 整日思想詭計。
PS|38|13|但我如聾子聽不見， 像啞巴不能開口。
PS|38|14|我如聽不見的人， 無法用口答辯。
PS|38|15|耶和華啊，我仰望你！ 主－我的上帝啊，你必應允我！
PS|38|16|我曾說：「恐怕他們向我誇耀， 我失腳的時候，他們向我誇口。」
PS|38|17|我就要跌倒， 我的痛苦常在我面前。
PS|38|18|我要承認我的罪孽， 要因我的罪憂愁。
PS|38|19|但我的仇敵又活潑又強壯， 無理恨我的增多了。
PS|38|20|以惡報善的與我作對， 但我追求良善。
PS|38|21|耶和華啊，求你不要撇棄我！ 我的上帝啊，求你不要遠離我！
PS|38|22|拯救我的主啊， 求你快快幫助我！
PS|39|1|我曾說：「我要謹慎我的言行， 免得我的舌頭犯罪； 惡人在我面前的時候， 我要用嚼環勒住我的口。」
PS|39|2|我默然無聲，連好話也不出口， 我的愁苦就更加深。
PS|39|3|我的心在我裏面發熱； 我默想的時候，火就燒起， 我用舌頭說話：
PS|39|4|「耶和華啊，求你讓我曉得我的結局， 我的壽數幾何， 使我知道我的生命何等短暫！
PS|39|5|看哪，你使我的年日窄如手掌， 我一生的年數，在你面前如同無有； 各人最穩妥的時候，真是全然虛幻。（細拉）
PS|39|6|世人行動實係幻影， 他們忙亂，真是枉然， 積蓄財寶，不知將來有誰收取。
PS|39|7|「主啊，如今我等甚麼呢？ 我的指望在乎你！
PS|39|8|求你救我脫離一切的過犯， 不要使我受愚頑人的羞辱。
PS|39|9|我保持沉默，閉口不言， 因為這一切都是你所做的。
PS|39|10|求你從我身上免去你的責罰； 因你手的責打，我就消滅。
PS|39|11|因人的罪惡你懲罰管教他的時候， 如蛀蟲一般，吃掉他所喜愛的。 世人真是虛幻！（細拉）
PS|39|12|「耶和華啊，求你聽我的禱告， 側耳聽我的呼求！ 我流淚，求你不要靜默無聲！ 因為在你面前我是客旅， 是寄居的，像我列祖一般。
PS|39|13|求你寬容我， 使我在去而不返之先可以喜樂。」
PS|40|1|我曾耐性等候耶和華， 他垂聽我的呼求。
PS|40|2|他從泥坑裏， 從淤泥中，把我拉上來， 使我的腳立在磐石上， 使我腳步穩健。
PS|40|3|他使我口唱新歌， 就是讚美我們上帝的話。 許多人必看見而懼怕， 並要倚靠耶和華。
PS|40|4|那倚靠耶和華、 不理會狂傲和偏向虛假的， 這人有福了！
PS|40|5|耶和華－我的上帝啊，你所行的奇事 和你為我們設想的計劃，多到無法盡述； 若要述說陳明，不可勝數。
PS|40|6|祭物和禮物，你不喜愛， 你已經開通我的耳朵； 燔祭和贖罪祭非你所要。
PS|40|7|那時我說：「看哪，我來了！ 我的事在經卷上已經記載了。
PS|40|8|我的上帝啊，我樂意照你的旨意行， 你的律法在我心裏。」
PS|40|9|我在大會中傳講公義的佳音， 看哪，必不制止我的嘴唇； 耶和華啊，這一切你都知道。
PS|40|10|我未曾把你的公義藏在心裏， 我已陳明你的信實和你的救恩； 在大會中我未曾隱瞞你的慈愛和信實。
PS|40|11|耶和華啊，求你不要向我止住你的憐憫！ 願你的慈愛和信實常常保佑我！
PS|40|12|因有無數的禍患圍困我， 我的罪孽追上了我，使我不能看見， 這罪孽比我的頭髮還多， 我的膽量喪失了。
PS|40|13|耶和華啊，求你開恩搭救我！ 耶和華啊，求你速速幫助我！
PS|40|14|願那些尋找我、要滅我命的，一同抱愧蒙羞！ 願那些喜悅我遭害的，退後受辱！
PS|40|15|願那些對我說「啊哈、啊哈」的， 因羞愧而敗亡！
PS|40|16|願一切尋求你的，因你歡喜快樂！ 願那些喜愛你救恩的，常說：「當尊耶和華為大！」
PS|40|17|我本是困苦貧窮的，主卻顧念我。 你是幫助我的，搭救我的； 我的上帝啊，求你不要耽延！
PS|41|1|眷顧貧寒人的有福了 ！ 在患難的日子，耶和華必搭救他。
PS|41|2|耶和華必保全他，使他存活， 他要在地上享福。 求你不要把他交給仇敵，遂其所願。
PS|41|3|他病重在榻，耶和華必扶持他； 他在病中，你必使他離開病床。
PS|41|4|我曾說：「耶和華啊，求你憐憫我， 醫治我，因為我得罪了你。」
PS|41|5|我的仇敵用惡言議論我： 「他幾時才會死，他的名幾時才會消滅呢？」
PS|41|6|當他來看我的時候，說的是假話； 他心存奸惡，走到外邊才說出來。
PS|41|7|所有恨我的，都一同交頭接耳議論我， 他們設計要害我。
PS|41|8|他們說：「他有怪病纏身， 他已躺下，必不能再起來。」
PS|41|9|連我知己的朋友， 我所信賴、吃我飯的人也用腳踢我。
PS|41|10|耶和華啊，求你憐憫我， 使我起來，好報復他們！
PS|41|11|我因此就知道你喜愛我， 我的仇敵不得向我誇勝。
PS|41|12|你因我純正就扶持我， 使我永遠站立在你面前。
PS|41|13|耶和華－ 以色列 的上帝是應當稱頌的， 從亙古直到永遠。阿們！阿們！ 可拉後裔的詩。交給聖詠團長。
PS|42|1|上帝啊，我的心切慕你， 如鹿切慕溪水。
PS|42|2|我的心渴想上帝，就是永生上帝， 我幾時得朝見上帝呢？
PS|42|3|我晝夜以眼淚當食物， 人不住地對我說：「你的上帝在哪裏呢？」
PS|42|4|我從前與眾人同往， 領他們到上帝的殿裏， 大家用歡呼稱頌的聲音守節； 我追想這些事， 我的心極其悲傷。
PS|42|5|我的心哪，你為何憂悶？ 為何在我裏面煩躁？ 應當仰望上帝， 因我還要稱謝他，我當面的拯救，
PS|42|6|我的上帝。我的心在我裏面憂悶， 所以我從 約旦 地， 從 黑門嶺 ，從 米薩山 記念你。
PS|42|7|你的瀑布發聲，深淵就與深淵響應， 你的波浪洪濤漫過我身。
PS|42|8|白晝，耶和華必施慈愛； 黑夜，我要歌頌祈禱賜我生命的上帝。
PS|42|9|我要對上帝－我的磐石說： 「你為何忘記我呢？ 我為何因仇敵的欺壓時常哀痛呢？」
PS|42|10|我的敵人辱罵我， 好像敲碎我的骨頭， 他們不住地對我說： 「你的上帝在哪裏呢？」
PS|42|11|我的心哪，你為何憂悶？ 為何在我裏面煩躁？ 應當仰望上帝， 因我還要稱謝他，我當面的拯救，我的上帝。
PS|43|1|上帝啊，求你為我伸冤， 向不虔誠的國為我辯護； 求你救我脫離詭詐不義的人。
PS|43|2|你是作我保障 的上帝，為何丟棄我呢？ 我為何因仇敵的欺壓時常哀痛呢？
PS|43|3|求你發出你的亮光和信實，好引導我， 帶我到你的聖山，到你的居所！
PS|43|4|我就走到上帝的祭壇， 到賜我喜樂的上帝那裏。 上帝，我的上帝啊， 我要彈琴稱謝你！
PS|43|5|我的心哪，你為何憂悶？ 為何在我裏面煩躁？ 應當仰望上帝， 我還要稱謝他，我當面的拯救，我的上帝。
PS|44|1|上帝啊，你在古時， 我們列祖的日子所做的事， 我們親耳聽見了， 我們的列祖曾為我們述說。
PS|44|2|你曾用手趕出外邦人， 卻栽培了我們的列祖； 你苦待萬民， 卻叫我們的列祖發達。
PS|44|3|因為他們不是靠自己的刀劍承受土地， 也不是靠自己的膀臂得勝， 而是靠你的右手、你的膀臂， 和你臉上的亮光， 因為你喜愛他們。
PS|44|4|上帝啊，你是我的君王， 求你發命令使 雅各 得勝。
PS|44|5|靠你，我們要推倒我們的敵人； 靠你的名，我們要踐踏那興起攻擊我們的人。
PS|44|6|因為我必不倚靠我的弓， 我的刀也不能使我得勝。
PS|44|7|惟有你拯救我們脫離敵人， 使恨我們的人羞愧。
PS|44|8|我們要常常因上帝誇耀， 要永遠頌揚你的名。（細拉）
PS|44|9|但如今你丟棄了我們，使我們受辱， 不和我們的軍隊同去。
PS|44|10|你使我們在敵人前轉身撤退， 使那恨我們的人任意搶奪。
PS|44|11|你使我們如羊當作食物， 把我們分散在列國中。
PS|44|12|你賣了你的子民也不獲利， 所得的並未加添你的資財。
PS|44|13|你使我們受鄰國的羞辱， 被四圍的人嗤笑譏諷。
PS|44|14|你使我們在列國中成了笑柄， 在萬民中使人搖頭。
PS|44|15|因辱罵者和毀謗者的聲音， 因仇敵和報仇者的緣故， 我的凌辱常常在我面前， 我臉上的羞愧將我遮蔽，
PS|44|16|
PS|44|17|這些事都臨到我們身上， 我們卻沒有忘記你， 也沒有違背你的約；
PS|44|18|我們的心並未退縮， 我們的腳也沒有偏離你的路。
PS|44|19|你在野狗出沒之處壓傷我們， 以死蔭籠罩我們。
PS|44|20|倘若我們忘記上帝的名， 或向外邦神明舉手，
PS|44|21|上帝豈不鑒察這事嗎？ 因為他曉得人心裏的隱祕。
PS|44|22|我們為你的緣故終日被殺， 人看我們如將宰的羊。
PS|44|23|主啊，求你睡醒，為何儘睡呢？ 求你醒來，不要永遠丟棄我們！
PS|44|24|你為何轉臉， 不顧我們所遭的苦難和所受的欺壓呢？
PS|44|25|我們俯伏在塵土上， 我們的肚腹緊貼地面。
PS|44|26|求你興起幫助我們！ 因你的慈愛救贖我們！
PS|45|1|我心裏湧出美辭， 我為王朗誦我的詩章， 我的舌頭是敏捷文士的手筆。
PS|45|2|你比世人更美， 你嘴裏滿有恩惠； 所以上帝賜福給你，直到永遠。
PS|45|3|勇士啊，願你腰間佩刀， 大展榮耀和威嚴，
PS|45|4|為真理、謙卑、公義威嚴地駕車前進，無不得勝； 願你的右手顯明可畏的事。
PS|45|5|你的箭鋒快，射中王的仇敵的心， 萬民仆倒在你之下。
PS|45|6|上帝啊，你的寶座是永永遠遠的， 你國度的權杖是正直的權杖。
PS|45|7|你喜愛公義，恨惡罪惡， 所以上帝，就是你的上帝，用喜樂油膏你， 勝過膏你的同伴。
PS|45|8|你的衣服散發沒藥、沉香、肉桂的香氣， 象牙宮中絲弦樂器的聲音使你歡喜。
PS|45|9|你的妃嬪之中有列王的女兒， 王后佩戴 俄斐 金飾站立在你右邊。
PS|45|10|女子啊，要傾聽，要思想，要側耳而聽！ 不要記念你本族和你父家，
PS|45|11|王就羨慕你的美貌； 因為他是你的主，你當向他下拜。
PS|45|12|推羅 必來送禮， 百姓中富足的人也必向你求恩。
PS|45|13|君王的女兒在宮裏極其榮華， 她的衣服是金線繡的；
PS|45|14|她穿錦繡的衣服，引到王面前， 陪伴她的童女隨從她，也被帶到你面前。
PS|45|15|她們要歡喜快樂， 被引導進入王宮。
PS|45|16|你的子孫要接續你列祖， 你要立他們在各地作王。
PS|45|17|我必使萬代記念你的名， 萬民要永永遠遠稱謝你。
PS|46|1|上帝是我們的避難所，是我們的力量， 是我們在患難中隨時的幫助。
PS|46|2|所以，地雖改變， 山雖搖動到海心，
PS|46|3|其中的水雖澎湃翻騰， 山雖因海漲而戰抖， 我們也不害怕。（細拉）
PS|46|4|有一道河，這河的分汊使上帝的城歡喜， 這城就是至高者居住的聖所。
PS|46|5|上帝在其中，城必不動搖； 到天一亮，上帝必幫助這城。
PS|46|6|萬邦喧嚷，國度動搖； 上帝出聲，地就熔化。
PS|46|7|萬軍之耶和華與我們同在， 雅各 的上帝是我們的避難所！（細拉）
PS|46|8|你們來看耶和華的作為， 看他使地怎樣荒涼。
PS|46|9|他止息戰爭，直到地極； 他折弓、斷槍，把戰車焚燒在火中。
PS|46|10|你們要休息，要知道我是上帝！ 我必在列國中受尊崇，在全地也受尊崇。
PS|46|11|萬軍之耶和華與我們同在， 雅各 的上帝是我們的避難所！
PS|47|1|萬民哪，你們都要鼓掌！ 用歡呼的聲音向上帝呼喊！
PS|47|2|因為耶和華至高者是可畏的， 他是治理全地的大君王。
PS|47|3|他使萬民服在我們以下， 又使萬族服在我們腳下。
PS|47|4|他為我們選擇產業， 就是他所愛之 雅各 的榮耀。（細拉）
PS|47|5|上帝上升，有喊聲相送； 耶和華上升，有角聲相送。
PS|47|6|你們要向上帝歌頌，歌頌！ 向我們的王歌頌，歌頌！
PS|47|7|因為上帝是全地的王， 你們要用聖詩歌頌！
PS|47|8|上帝作王治理列國， 上帝坐在他的聖寶座上。
PS|47|9|萬民的君王聚集， 要作 亞伯拉罕 的上帝的子民， 因為地上的盾牌是屬上帝的， 他為至高！
PS|48|1|耶和華本為大！ 在我們上帝的城中， 在他的聖山上， 當受大讚美。
PS|48|2|錫安山 －大君王的城， 在北面居高華美， 為全地所喜悅。
PS|48|3|上帝在城的宮殿中， 自顯為避難所。
PS|48|4|看哪，諸王會合， 一同經過。
PS|48|5|他們見了這城就驚奇喪膽， 急忙逃跑。
PS|48|6|戰兢在那裏抓住他們， 他們好像臨產的婦人一樣陣痛。
PS|48|7|上帝啊，你用東風擊破 他施 的船隻。
PS|48|8|我們在萬軍之耶和華的城裏， 就是我們上帝的城裏， 所看見的正如我們所聽見的。 上帝必堅立這城，直到永遠。（細拉）
PS|48|9|上帝啊，我們在你的殿中 想念你的慈愛。
PS|48|10|上帝啊，你受的讚美正與你的名相稱，直到地極！ 你的右手滿了公義。
PS|48|11|因你的判斷， 錫安山 應當歡喜， 猶大 的城鎮 應當快樂。
PS|48|12|你們當周遊 錫安 ， 四圍環繞，數點城樓，
PS|48|13|細看它的城郭， 察看它的宮殿， 為要傳揚給後代。
PS|48|14|因為這上帝永永遠遠為我們的上帝， 他必作我們引路的，直到死時 。
PS|49|1|萬民哪，你們都當聽這話！ 世上所有的居民， 無論貴賤貧富， 都當側耳而聽！
PS|49|2|
PS|49|3|我口要說智慧的言語， 我心思想通達的道理。
PS|49|4|我要側耳聽比喻， 用琴解謎語。
PS|49|5|在患難的日子，追逼我的人的奸惡 環繞我， 我何必懼怕？
PS|49|6|他們那些倚靠財貨， 自誇錢財多的人，
PS|49|7|沒有一個能贖自己的弟兄 ， 能將贖價給上帝，
PS|49|8|讓他長遠活著，不見地府 ； 因為贖生命的價值極貴， 只可永遠罷休。
PS|49|9|
PS|49|10|他要見智慧人死， 愚昧人和畜牲一般的人一同滅亡， 把他們的財貨留給別人。
PS|49|11|他們雖以自己的名叫自己的地， 墳墓卻作他們永遠的家， 作他們世世代代的居所。
PS|49|12|人居尊貴中不能長久， 如同死亡的畜類一樣。
PS|49|13|他們所行之道本為自己的愚昧， 後來的人卻還佩服他們的話語。（細拉）
PS|49|14|他們如同羊群註定要下陰間， 死亡必作他們的牧者； 到了早晨，正直人必管轄他們。 他們的形像必被陰間所滅，無處可容身。
PS|49|15|然而上帝必救贖我的命脫離陰間的掌控， 因他必收納我。（細拉）
PS|49|16|見人發財、家室日益顯赫的時候， 你不要懼怕；
PS|49|17|因為他死的時候甚麼也不能帶去， 他的榮耀不能隨他下去。
PS|49|18|他活著的時候，雖然自誇為有福 ─你若自己行得好，人必誇獎你─
PS|49|19|他仍必與歷代的祖宗一樣同歸死亡， 永不見光。
PS|49|20|人在尊貴中而不醒悟， 就如死亡的畜類一樣。
PS|50|1|大能者上帝－耶和華已經發言呼召天下， 從日出之地到日落之處。
PS|50|2|從全然美麗的 錫安 中， 上帝已經發光了。
PS|50|3|我們的上帝要來，絕不閉口； 有烈火在他面前吞滅， 有暴風在他四圍颳起。
PS|50|4|他呼召上天下地， 為要審判他的子民：
PS|50|5|「召集我的聖民， 就是那些用祭物與我立約的人，到我這裏來。」
PS|50|6|諸天必表明他的公義， 因為上帝是施行審判的。（細拉）
PS|50|7|「聽啊，我的子民，我要說話！ 以色列 啊，我要審問你； 我是上帝，是你的上帝！
PS|50|8|我並不因你的祭物責備你； 你的燔祭常在我面前。
PS|50|9|我不從你家中取公牛， 也不從你圈內取公山羊；
PS|50|10|因為，林中的百獸是我的， 千山的牲畜也是我的。
PS|50|11|山中 的飛鳥，我都知道， 田野的走獸也都屬我。
PS|50|12|「我若是飢餓，不用告訴你， 因為世界和其中所充滿的都是我的。
PS|50|13|我豈吃公牛的肉呢？ 我豈喝公山羊的血呢？
PS|50|14|你們要以感謝為祭獻給上帝， 又要向至高者還你的願，
PS|50|15|並要在患難之日求告我， 我必搭救你，你也要榮耀我。」
PS|50|16|但上帝對惡人說：「你怎敢傳講我的律例， 口中提到我的約呢？
PS|50|17|其實你恨惡管教， 將我的言語拋在腦後。
PS|50|18|你見了盜賊就樂意與他同夥， 又和行姦淫的人同流合污。
PS|50|19|「你的口出惡言， 你的舌編造詭詐。
PS|50|20|你坐著，毀謗你的兄弟， 讒害你親母的兒子。
PS|50|21|你做了這些事，我閉口不言， 你想我正如你一樣； 其實我要責備你，將這些事擺在你眼前。
PS|50|22|「你們忘記上帝的，要思想這事， 免得我把你們撕碎，無人搭救。
PS|50|23|凡以感謝獻祭的就是榮耀我； 那按正路而行的，我必使他得著上帝的救恩。」
PS|51|1|上帝啊，求你按你的慈愛恩待我！ 按你豐盛的憐憫塗去我的過犯！
PS|51|2|求你將我的罪孽洗滌淨盡， 潔除我的罪！
PS|51|3|因為我知道我的過犯； 我的罪常在我面前。
PS|51|4|我向你犯罪，惟獨得罪了你， 在你眼前行了這惡， 以致你責備的時候顯為公義， 判斷的時候顯為清白。
PS|51|5|看哪，我是在罪孽裏生的， 在我母親懷胎的時候就有了罪。
PS|51|6|你所喜愛的是內心的誠實； 求你在我隱密處使我得智慧。
PS|51|7|求你用牛膝草潔淨我，我就乾淨； 求你洗滌我，我就比雪更白。
PS|51|8|求你使我得聽歡喜快樂的聲音， 使你所壓傷的骨頭可以踴躍。
PS|51|9|求你轉臉不看我的罪， 塗去我一切的罪孽。
PS|51|10|上帝啊，求你為我造清潔的心， 使我裏面重新有正直 的靈。
PS|51|11|不要丟棄我，使我離開你的面； 不要從我收回你的聖靈。
PS|51|12|求你使我重得救恩之樂， 以樂意的靈來扶持我，
PS|51|13|我就把你的道指教有過犯的人， 罪人必歸順你。
PS|51|14|上帝啊，你是拯救我的上帝； 求你救我脫離流人血的罪！ 我的舌頭就高唱你的公義。
PS|51|15|主啊，求你使我嘴唇張開， 我的口就傳揚讚美你的話！
PS|51|16|你本不喜愛祭物，若喜愛，我就獻上； 燔祭你也不喜悅。
PS|51|17|上帝所要的祭就是憂傷的靈； 上帝啊，憂傷痛悔的心，你必不輕看。
PS|51|18|求你隨你的美意善待 錫安 ， 建造 耶路撒冷 的城牆。
PS|51|19|那時，你必喜愛公義的祭 和燔祭，全牲的燔祭； 那時，人必將公牛獻在你壇上。
PS|52|1|勇士啊，你為何作惡自誇？ 上帝的慈愛是常存的。
PS|52|2|你這行詭詐的人哪， 你的舌頭像快利的剃刀，圖謀毀滅。
PS|52|3|你愛惡勝似愛善， 又愛說謊，勝於愛說公義。（細拉）
PS|52|4|詭詐的舌頭啊， 你愛說一切毀滅的話！
PS|52|5|上帝也要毀滅你，直到永遠。 他要抓住你，從帳棚中拉你出來， 從活人之地將你拔除。（細拉）
PS|52|6|義人要看見而懼怕， 並要笑他。
PS|52|7|看哪，這就是那不以上帝為保障的人， 他只倚靠豐富的財物，在邪惡上堅立自己。
PS|52|8|至於我，就像上帝殿中的青橄欖樹， 我永永遠遠倚靠上帝的慈愛。
PS|52|9|我要稱謝你，直到永遠， 因為你做了這事。 我也要在你聖民面前仰望你的名， 這名本為美好。
PS|53|1|愚頑人心裏說：「沒有上帝。」 他們都敗壞，行了可憎惡的罪孽， 沒有一個人行善。
PS|53|2|上帝從天上垂看世人， 要看有明白的沒有， 有尋求上帝的沒有。
PS|53|3|他們全都退後，一同變為污穢， 沒有行善的， 連一個也沒有。
PS|53|4|作惡的都沒有知識嗎？ 他們吞吃我的百姓如同吃飯一樣， 並不求告上帝。
PS|53|5|他們在無可懼怕之處就大大害怕， 因為上帝使那安營攻擊你之人的骨頭散開了。 你使他們蒙羞，因為上帝棄絕了他們。
PS|53|6|但願 以色列 的救恩出自 錫安 。 當上帝救回他被擄子民的時候， 雅各 要快樂， 以色列 要歡喜。
PS|54|1|上帝啊，求你因你的名拯救我， 憑你的大能為我伸冤。
PS|54|2|上帝啊，求你聽我的禱告， 側耳聽我口中的言語。
PS|54|3|因為陌生人興起攻擊我， 強橫的人尋索我的性命； 他們眼中沒有上帝。（細拉）
PS|54|4|看哪，上帝是幫助我的， 主是扶持我性命的，
PS|54|5|他要報應我仇敵所作的惡； 求你憑你的信實滅絕他們。
PS|54|6|我要把甘心祭獻給你； 耶和華啊，我要頌揚你的名，這名本為美好。
PS|54|7|他從一切的急難中把我救出來， 我的眼睛也看見了我的仇敵遭報。
PS|55|1|上帝啊，求你側耳聽我的禱告， 不要隱藏不聽我的懇求！
PS|55|2|求你留心聽我，應允我。 我哀嘆不安，發出呻吟，
PS|55|3|都因仇敵的聲音，惡人的欺壓； 他們將罪孽加在我身上，發怒氣加害我。
PS|55|4|我的心在我裏面陣痛， 死亡的恐怖落在我身。
PS|55|5|恐懼戰兢臨到了我， 驚恐籠罩我。
PS|55|6|我說：「但願我有翅膀像鴿子， 我就飛去，得享安息。
PS|55|7|看哪，我要遠走高飛， 宿在曠野。（細拉）
PS|55|8|我要速速逃到避難之所， 脫離狂風暴雨。」
PS|55|9|主啊，求你吞滅他們，變亂他們的言語！ 因為我在城中見了兇暴爭吵的事。
PS|55|10|他們晝夜在城牆上繞行， 城內也有罪孽和奸惡。
PS|55|11|邪惡在其中， 欺壓和詭詐不離街市。
PS|55|12|原來，不是仇敵辱罵我， 若是仇敵，還可忍受； 也不是恨我的人向我狂妄自大， 若是恨我的人，我必躲避他。
PS|55|13|不料是你；你原與我同等， 是我的朋友，是我的知己！
PS|55|14|我們素常彼此交談，以為甘甜； 我們結伴在上帝的殿中同行。
PS|55|15|願死亡忽然臨到他們！ 願他們活生生地下入陰間！ 因為他們的住處都是邪惡， 他們的內心充滿奸惡。
PS|55|16|至於我，我要求告上帝， 耶和華必拯救我。
PS|55|17|晚上、早晨、中午我要哀聲悲嘆， 他就垂聽我的聲音。
PS|55|18|他救贖我的命脫離攻擊我的人， 使我得享平安， 因為與我相爭的人很多。
PS|55|19|那不願改變、不敬畏上帝的人， 從太古常存的上帝必聽見而使他受苦。（細拉）
PS|55|20|他背了約， 伸手攻擊與他和好的人。
PS|55|21|他的口如奶油光滑， 他的心卻懷著敵意； 他的話比油柔和， 其實是拔出的刀。
PS|55|22|你要把你的重擔卸給耶和華， 他必扶持你， 他永不叫義人動搖。
PS|55|23|上帝啊，你必使惡人墜入滅亡的坑； 那好流人血、行詭詐的人必活不過半生， 但我要倚靠你。
PS|56|1|上帝啊，求你憐憫我，因為有人踐踏我， 終日攻擊欺壓我。
PS|56|2|我的仇敵終日踐踏我， 逞驕傲攻擊我的人很多。
PS|56|3|我懼怕的時候要倚靠你。
PS|56|4|我倚靠上帝，我要讚美他的話語； 我倚靠上帝，必不懼怕。 血肉之軀能把我怎麼樣呢？
PS|56|5|他們終日扭曲我的話， 千方百計加害於我。
PS|56|6|他們聚集，埋伏，窺探我的腳蹤， 等候要害我的命。
PS|56|7|他們豈能脫罪呢 ？ 上帝啊，求你在怒中使萬民敗落！
PS|56|8|我幾次流離，你都數算； 求你把我的眼淚裝在你的皮袋裏。 這一切不都記在你的冊子上嗎？
PS|56|9|我呼求的日子，仇敵都要轉身撤退。 上帝幫助我，這是我所知道的。
PS|56|10|我倚靠上帝，我要讚美他的話語； 我倚靠耶和華，我要讚美他的話語。
PS|56|11|我倚靠上帝，必不懼怕。 人能把我怎麼樣呢？
PS|56|12|上帝啊，我要向你還所許的願， 我要以感謝祭回報你；
PS|56|13|因為你救我的命脫離死亡。 你保護我的腳不跌倒， 使我在生命的光中行在上帝面前。
PS|57|1|上帝啊，求你憐憫我，憐憫我， 因為我的心投靠你。 我要投靠在你翅膀蔭下， 直等到災害過去。
PS|57|2|我要求告至高的上帝， 就是為我成全萬事的上帝。
PS|57|3|那踐踏我的人辱罵我的時候， 上帝必從天上施恩救我，(細拉) 他必向我施行慈愛和信實。
PS|57|4|至於我的性命， 我好像躺臥在吞噬人的獅子當中； 他們的牙齒是槍、箭， 他們的舌頭是快刀。
PS|57|5|上帝啊，願你崇高過於諸天！ 願你的榮耀高過全地！
PS|57|6|他們為我的腳設下網羅，壓迫我； 他們在我面前掘了坑，自己反掉在其中。（細拉）
PS|57|7|上帝啊，我心堅定，我心堅定； 我要唱詩，我要歌頌！
PS|57|8|我的靈 啊，你當醒起！ 琴瑟啊，當醒起！ 我自己要極早醒起！
PS|57|9|主啊，我要在萬民中稱謝你， 在萬族中歌頌你！
PS|57|10|因為你的慈愛高及諸天， 你的信實達到穹蒼。
PS|57|11|上帝啊，願你崇高過於諸天！ 願你的榮耀高過全地！
PS|58|1|你們緘默不語，真合公義嗎？ 你們審判世人，豈按正直嗎？
PS|58|2|不然！你們心中作惡， 量出你們在地上手中的殘暴。
PS|58|3|惡人一出母胎就與上帝疏遠， 一離母腹就走錯路，說謊話。
PS|58|4|他們的毒氣好像蛇的毒氣， 他們好像聾的毒蛇塞住耳朵，
PS|58|5|聽不見弄蛇者的聲音， 也聽不見魔術師的咒語。
PS|58|6|上帝啊，求你敲碎他們口中的牙！ 耶和華啊，求你敲掉少壯獅子的大牙！
PS|58|7|願他們消滅，如急流的水一般； 他們瞄準射箭的時候，箭頭彷彿折斷。
PS|58|8|願他們像蝸牛腐爛消失， 又像婦人流掉的胎兒，未見天日。
PS|58|9|你們用荊棘燒火，鍋還未熱， 上帝就用旋風把未燒著的和已燒著的一齊颳去。
PS|58|10|義人見仇敵遭報就歡喜， 他要在惡人的血中洗腳。
PS|58|11|因此，人必說：「義人誠然有善報， 在地上果然有施行審判的上帝！」
PS|59|1|我的上帝啊，求你救我脫離仇敵， 把我安置在高處，脫離那些起來攻擊我的人。
PS|59|2|求你救我脫離作惡的人， 救我脫離好流人血的人！
PS|59|3|因為他們埋伏要害我命， 強悍的人聚集攻擊我， 耶和華啊，不是為我的過犯， 也不是為我的罪愆。
PS|59|4|我雖然無過，他們急忙擺陣攻擊我。 求你興起，來幫助我，來鑒察！
PS|59|5|萬軍之耶和華上帝－ 以色列 的上帝啊， 求你醒起，懲治萬國！ 不要憐憫行詭詐的惡人！（細拉）
PS|59|6|他們晚上轉回， 叫號如狗，圍城繞行。
PS|59|7|看哪，他們口中噴吐惡言， 嘴裏有刀： 「有誰聽見呢？」
PS|59|8|但你－耶和華必譏笑他們， 你要嗤笑萬國。
PS|59|9|我 的力量啊，我要等候你， 因為上帝是我的庇護所。
PS|59|10|我的上帝要以慈愛 迎接我， 上帝要叫我看見我的仇敵遭報。
PS|59|11|主，我們的盾牌啊， 不要殺他們，免得我的子民遺忘； 求你用你的能力使他們四散， 使他們降為卑。
PS|59|12|願他們因口中的罪和嘴唇的言語， 被自己的驕傲抓住， 他們所說的盡是咒罵和謊話。
PS|59|13|求你發怒，使他們消滅， 求你使他們消滅，歸於無有， 使他們知道上帝在 雅各 中間掌權， 直到地極。（細拉）
PS|59|14|他們晚上轉回， 叫號如狗，圍城繞行。
PS|59|15|他們到處走動覓食， 若不飽足就咆哮不已。
PS|59|16|但我要歌頌你的能力， 早晨要高唱你的慈愛； 因為你是我的庇護所， 在急難的日子作過我的避難所。
PS|59|17|我的力量啊，我要歌頌你； 因為上帝是我的庇護所， 是賜恩給我的上帝。
PS|60|1|上帝啊，你丟棄了我們，破壞了我們； 你曾發怒，求你使我們復興！
PS|60|2|你使地震動，崩裂； 求你將裂口補好，因為地在搖動。
PS|60|3|你讓你的子民遇見艱難， 使我們喝那令人東倒西歪的酒。
PS|60|4|你把旌旗賜給敬畏你的人， 可以躲避弓箭 。（細拉）
PS|60|5|求你應允我們 ，用右手施行拯救， 好讓你所親愛的人得救。
PS|60|6|上帝在他的聖所 說： 「我要歡樂； 要劃分 示劍 ， 丈量 疏割谷 。
PS|60|7|基列 是我的， 瑪拿西 是我的。 以法蓮 是護衛我頭的， 猶大 是我的權杖。
PS|60|8|摩押 是我的沐浴盆， 我要向 以東 扔鞋。 非利士 啊，你還能因我歡呼嗎？」
PS|60|9|誰能領我進堅固城？ 誰能引我到 以東 地？
PS|60|10|上帝啊，你真的丟棄了我們嗎？ 上帝啊，你不和我們的軍隊同去嗎？
PS|60|11|求你幫助我們攻擊敵人， 因為人的幫助是枉然的。
PS|60|12|我們倚靠上帝才得施展大能， 因為踐踏我們敵人的就是他。
PS|61|1|上帝啊，求你聽我的呼求， 留心聽我的禱告！
PS|61|2|我心裏發昏的時候， 要從地極求告你。 求你領我到那比我更高的磐石，
PS|61|3|因為你是我的避難所， 是我的堅固臺，使我脫離仇敵。
PS|61|4|我要永遠住在你的帳幕裏！ 我要投靠在你翅膀下的隱密處！（細拉）
PS|61|5|上帝啊，你聽了我所許的願； 你將產業賜給敬畏你名的人。
PS|61|6|求你加添王的壽數， 使他的年歲存到世世代代。
PS|61|7|願他在上帝面前永遠坐在王位上， 求你預備慈愛和信實保佑他！
PS|61|8|這樣，我要歌頌你的名，直到永遠， 天天還我所許的願。
PS|62|1|我的心默默無聲，專等候上帝， 我的救恩從他而來。
PS|62|2|惟獨他是我的磐石，我的拯救； 他是我的庇護所，我必不大大動搖。
PS|62|3|你們大家攻擊一人，使他被殺， 如歪斜的牆、將倒的壁，要到幾時呢？
PS|62|4|他們彼此商議，要把他從高位上拉下來； 他們喜愛謊話，口雖祝福，心卻詛咒。（細拉）
PS|62|5|我的心哪，你當默默無聲，專等候上帝， 因為我的盼望是從他而來。
PS|62|6|惟獨他是我的磐石，我的拯救； 他是我的庇護所，我必不動搖。
PS|62|7|我的拯救、我的榮耀都在於上帝； 我力量的磐石、我的避難所都在於上帝。
PS|62|8|百姓啊，要時時倚靠他， 在他面前傾心吐意； 上帝是我們的避難所。（細拉）
PS|62|9|人真是虛空， 人真是虛假； 放在天平裏就必浮起， 他們一共比空氣還輕。
PS|62|10|不要仗勢欺人， 也不要因搶奪而驕傲； 若財寶加增，不要放在心上。
PS|62|11|上帝說了一次、兩次，我都聽見了， 就是能力屬乎上帝。
PS|62|12|主啊，慈愛也是屬乎你， 因為你照著各人所做的報應他。
PS|63|1|上帝啊，你是我的上帝， 我要切切尋求你； 在乾旱疲乏無水之地， 我的心靈渴想你，我的肉身切慕你。
PS|63|2|我在聖所中曾如此瞻仰你， 為要見你的能力和你的榮耀。
PS|63|3|因你的慈愛比生命更好， 我的嘴唇要頌讚你。
PS|63|4|我還活著的時候要這樣稱頌你， 我要奉你的名舉手。
PS|63|5|我在床上記念你， 在夜更的時候思念你； 我的心像吃飽了骨髓肥油， 我也要以歡樂的嘴唇讚美你。
PS|63|6|
PS|63|7|因為你曾幫助了我， 我要在你翅膀的蔭下歡呼。
PS|63|8|我的心緊緊跟隨你； 你的右手扶持了我。
PS|63|9|但那些尋索要滅我命的人 必往地底下去；
PS|63|10|他們必被刀劍所殺， 成為野狗的食物。
PS|63|11|但是王必因上帝歡喜， 凡指著他發誓的都要誇耀， 因為說謊之人的口必被塞住。
PS|64|1|上帝啊，我哀嘆的時候，求你聽我的聲音！ 求你保護我的性命，不受仇敵的驚嚇！
PS|64|2|求你把我隱藏， 使我脫離作惡之人的暗謀， 脫離作孽之人的擾亂。
PS|64|3|他們磨舌如刀， 發出苦毒的言語，好像瞄準了的箭，
PS|64|4|要在暗地裏射完全人； 他們忽然射他，並不懼怕。
PS|64|5|他們彼此勉勵，設下惡計； 他們商量，暗設圈套， 說：「誰能看見呢？」
PS|64|6|他們圖謀奸惡： 「我們完成了精密的策劃。」 各人的意念心思是深沉的。
PS|64|7|但上帝要用箭射他們， 他們忽然受了傷。
PS|64|8|他們必然絆跌，被自己的舌頭所害； 凡看見他們的都必搖頭。
PS|64|9|眾人都要害怕， 要傳揚上帝的工作， 並且明白他的作為。
PS|64|10|義人必因耶和華歡喜，並要投靠他； 凡心裏正直的人都必誇耀。
PS|65|1|上帝啊，在 錫安 ，人都等候讚美你， 也要向你還所許的願。
PS|65|2|聽禱告的主啊， 凡有血肉之軀的都要來就你。
PS|65|3|罪孽勝了我； 至於我們的過犯，你都要赦免。
PS|65|4|你所揀選、使他親近你、住在你院中的， 這人有福了！ 我們要因你居所、你聖殿的美福知足。
PS|65|5|拯救我們的上帝啊，你必以威嚴秉公義應允我們； 地極和海角遠方的人都倚靠你。
PS|65|6|你既以大能束腰， 就用力量安定諸山，
PS|65|7|使諸海的響聲和其中波浪的響聲， 並萬民的喧嘩，都平靜了。
PS|65|8|住在地極的人因你的神蹟懼怕， 你使日出日落之地都歡呼。
PS|65|9|你眷顧地， 降雨使地大大肥沃。 上帝的河滿了水； 你這樣澆灌了地， 好為人預備五穀。
PS|65|10|你澆透地的犁溝，潤澤犁脊， 降甘霖，使地鬆軟； 其中生長的，蒙你賜福。
PS|65|11|你以恩惠為年歲的冠冕， 你的路徑都滴下油脂，
PS|65|12|滴在曠野的草場上。 小山以歡樂束腰，
PS|65|13|草場以羊群為衣， 谷中也長滿了五穀； 這一切都歡呼歌唱。
PS|66|1|全地都當向上帝歡呼！
PS|66|2|當歌頌他名的榮耀， 使讚美他的話大有榮耀！
PS|66|3|當對上帝說：「你的作為何等可畏！ 因你的大能，仇敵要向你投降。
PS|66|4|全地要敬拜你，歌頌你， 要歌頌你的名。」（細拉）
PS|66|5|你們來看上帝所做的， 他向世人所做之事是可畏的。
PS|66|6|他將海變成乾地，使百姓步行過河； 我們在那裏要因他歡喜。
PS|66|7|他用權能治理，直到永遠。 他的眼睛鑒察萬民； 悖逆的人不可自高。（細拉）
PS|66|8|萬民哪，你們當稱頌我們的上帝， 使人得聽讚美他的聲音。
PS|66|9|他使我們的性命存活， 不叫我們的腳搖動。
PS|66|10|上帝啊，你曾考驗我們， 你熬煉我們，如煉銀子一樣。
PS|66|11|你使我們進入羅網， 把重擔放在我們身上。
PS|66|12|你使人坐車軋我們的頭； 我們經過水火， 你卻使我們到豐富之地。
PS|66|13|我要帶著燔祭進你的殿， 向你還我的願，
PS|66|14|就是在急難時我嘴唇所發的、 口中所許的。
PS|66|15|我要將肥牛的燔祭 和公羊的香祭獻給你， 又要把公牛和公山羊獻上。（細拉）
PS|66|16|敬畏上帝的人哪，你們都來聽！ 我要述說他為我所做的事。
PS|66|17|我曾用口求告他， 我的舌頭也稱他為高。
PS|66|18|我若心裏注重罪孽， 主必不聽。
PS|66|19|但上帝實在聽見了， 他留心聽了我禱告的聲音。
PS|66|20|上帝是應當稱頌的！ 他沒有推卻我的禱告， 也沒有使他的慈愛離開我。
PS|67|1|願上帝憐憫我們，賜福給我們， 使他的臉向我們發光，（細拉）
PS|67|2|好讓全地得知你的道路， 萬國得知你的救恩。
PS|67|3|上帝啊，願萬民稱謝你！ 願萬民都稱謝你！
PS|67|4|願萬族都快樂歡呼； 因為你必按公正審判萬民， 引導地上的萬族。（細拉）
PS|67|5|上帝啊，願萬民稱謝你！ 願萬民都稱謝你！
PS|67|6|地已經出了土產， 上帝，我們的上帝，要賜福給我們。
PS|67|7|上帝要賜福給我們， 地的四極都要敬畏他！
PS|68|1|願上帝興起，使他的仇敵四散， 使那恨他的人從他面前逃跑。
PS|68|2|你驅逐他們 ，如煙被吹散； 惡人見上帝的面就消滅，如蠟被火熔化。
PS|68|3|惟有義人必然歡喜， 在上帝面前快樂， 他們要在喜樂中歡欣。
PS|68|4|你們當向上帝唱詩，歌頌他的名； 為那駕車經過曠野的修平道路 。 他的名是耶和華， 你們要在他面前歡樂！
PS|68|5|上帝在他的聖所作孤兒的父， 作寡婦的伸冤者。
PS|68|6|上帝使孤獨的有家， 使被囚的出來享福； 惟有悖逆的要住在乾旱之地。
PS|68|7|上帝啊，當你走在百姓前頭， 在曠野行進，（細拉）
PS|68|8|地見上帝的面就震動，天也降雨； 西奈山 見 以色列 上帝的面也震動。
PS|68|9|上帝啊，你降下大雨； 你的產業 以色列 疲乏的時候，你使他堅固。
PS|68|10|你的會眾住在境內； 上帝啊，你在恩惠中為困苦人預備所需的。
PS|68|11|主發命令， 傳好信息的婦女成了大群：
PS|68|12|「統領大軍的君王逃跑了，逃跑了！」 在家等候的婦女也分得了掠物。
PS|68|13|你們躺臥在羊圈， 好像鴿子的翅膀鍍銀，翎毛鍍金一般。
PS|68|14|全能者在境內趕散列王的時候， 勢如飄雪在 撒們 。
PS|68|15|巴珊山 是極其宏偉 的山， 巴珊山 是多峰多嶺的山。
PS|68|16|你們多峰多嶺的山哪， 為何以妒忌的眼光看上帝所願居住的山？ 耶和華必住這山，直到永遠！
PS|68|17|上帝的車輦累萬盈千； 主在其中，好像在 西奈 聖山一樣。
PS|68|18|你已經升上高天，擄掠了俘虜； 你在人間，就是在悖逆的人中，受了供獻， 使耶和華上帝可以與他們同住。
PS|68|19|天天背負我們重擔的主， 就是拯救我們的上帝， 是應當稱頌的！（細拉）
PS|68|20|上帝是為我們施行拯救的上帝； 人能脫離死亡是在乎主─耶和華。
PS|68|21|但上帝要打破他仇敵的頭， 就是那常犯罪之人的頭顱。
PS|68|22|主說：「我要使百姓從 巴珊 歸來， 使他們從深海轉回，
PS|68|23|好叫你打碎仇敵，使你的腳踹在血中， 使你狗的舌頭也有份。」
PS|68|24|上帝啊，你是我的上帝，我的王； 人已經看見你行走，進入聖所。
PS|68|25|歌唱的行在前，作樂的隨在後， 都在擊鼓的童女中間：
PS|68|26|「從 以色列 源頭而來的啊， 你們當在各會中稱頌上帝─耶和華！」
PS|68|27|在那裏，有統管他們的小 便雅憫 ， 有 猶大 的領袖和他們的一群人， 有 西布倫 的領袖， 有 拿弗他利 的領袖。
PS|68|28|你的上帝已賜給你力量 ； 上帝啊，求你堅固你為我們所成全的事！
PS|68|29|因你 耶路撒冷 的殿， 列王必帶貢物獻給你。
PS|68|30|求你斥責蘆葦中的野獸和公牛群， 並萬民中的牛犢。 直到他們帶著銀塊來朝貢 ； 上帝已經趕散好戰的萬民 。
PS|68|31|埃及 的使臣要出來， 古實 人要急忙向上帝伸出手來。
PS|68|32|地上的國度啊， 你們要向上帝歌唱， 要歌頌主，（細拉）
PS|68|33|就是那駕行在亙古的諸天之上的主！ 聽啊，他發出聲音，是極大的聲音。
PS|68|34|你們要將能力歸給上帝； 他的威榮在 以色列 之上， 他的能力顯在天上。
PS|68|35|上帝啊，你從聖所顯為可畏， 以色列 的上帝是那將力量權能賜給他百姓的。 上帝是應當稱頌的！
PS|69|1|上帝啊，求你救我！ 因為眾水就要淹沒我。
PS|69|2|我深陷在淤泥中，沒有立腳之地； 我到了深水之中，波濤漫過我身。
PS|69|3|我因呼求困乏，喉嚨發乾； 我因等候上帝，眼睛失明。
PS|69|4|無故恨我的，比我的頭髮還多； 無理與我為仇、要把我剪除的，甚為強盛。 我沒有搶奪，他們竟然要我償還！
PS|69|5|上帝啊，我的愚昧，你原知道， 我的罪愆不能向你隱瞞。
PS|69|6|萬軍之主耶和華啊， 求你不要讓那等候你的因我蒙羞！ 以色列 的上帝啊， 求你不要讓那尋求你的因我受辱！
PS|69|7|因我為你的緣故受了辱罵， 滿面羞愧。
PS|69|8|我的兄弟把我當陌生人， 我母親的兒子把我當外邦人。
PS|69|9|因我為你的殿心裏焦急，如同火燒， 並且辱罵你的人的辱罵都落在我身上。
PS|69|10|我哭泣，以禁食刻苦我心； 這倒成了我的羞辱。
PS|69|11|我拿麻布當衣裳， 卻成了他們的笑柄。
PS|69|12|坐在城門口的談論我， 酒徒也以我為歌曲。
PS|69|13|至於我，耶和華啊，在悅納的時候我向你祈禱。 上帝啊，求你按你豐盛的慈愛， 憑你拯救的信實應允我！
PS|69|14|求你搭救我脫離淤泥， 不叫我陷在其中； 求你使我脫離那些恨我的人， 使我脫離深水。
PS|69|15|求你不容波濤漫過我， 不容深淵吞滅我， 不容深坑在我以上合口。
PS|69|16|耶和華啊，求你應允我！ 因為你的慈愛本為美好； 求你按你豐盛的憐憫轉回眷顧我！
PS|69|17|不要轉臉不顧你的僕人； 我在急難之中，求你速速應允我！
PS|69|18|求你親近我，救贖我！ 求你因我仇敵的緣故將我贖回！
PS|69|19|你知道我所受的辱罵、欺凌、羞辱； 我的敵人都在你面前。
PS|69|20|辱罵刺傷我的心， 使我憂愁。 我指望有人體恤，卻沒有一個； 指望有人安慰，卻找不著一個。
PS|69|21|他們拿苦膽給我當食物； 我渴了，他們拿醋給我喝。
PS|69|22|願他們的筵席在他們面前變為羅網， 在他們平安的時候 變為圈套。
PS|69|23|願他們的眼睛昏花，看不見； 求你使他們的腰常常戰抖。
PS|69|24|求你將你的惱恨倒在他們身上， 使你的烈怒追上他們。
PS|69|25|願他們的住處變為廢墟， 他們的帳棚無人居住。
PS|69|26|因為你所擊打的，他們就迫害； 你所擊傷的，他們述說 他的愁苦。
PS|69|27|求你使他們罪上加罪， 不容他們在你面前稱義。
PS|69|28|願他們從生命冊上被塗去， 不得名列在義人之中。
PS|69|29|但我困苦憂傷； 上帝啊，願你的救恩將我安置在高處。
PS|69|30|我要以詩歌讚美上帝的名， 以感謝尊他為大！
PS|69|31|這就讓耶和華喜悅，勝似獻牛， 獻有角有蹄的公牛。
PS|69|32|謙卑的人看見了就喜樂； 尋求上帝的人，願你們的心甦醒。
PS|69|33|因為耶和華聽了窮乏的人， 不藐視被囚的人。
PS|69|34|願天和地、 海洋和其中一切的動物都讚美他！
PS|69|35|因為上帝要拯救 錫安 ，建造 猶大 的城鎮； 他的子民要在那裏居住，得地為業。
PS|69|36|他僕人的後裔要承受這地， 愛他名的人要住在其中。
PS|70|1|上帝啊，求你快快搭救我！ 耶和華啊，求你速速幫助我！
PS|70|2|願那些尋索我命的，抱愧蒙羞； 願那些喜悅我遭害的，退後受辱。
PS|70|3|願那些對我說「啊哈、啊哈」的， 因羞愧退後。
PS|70|4|願所有尋求你的，因你歡喜快樂； 願那些喜愛你救恩的，常說：「當尊上帝為大！」
PS|70|5|但我是困苦貧窮的； 上帝啊，求你速速到我這裏來！ 你是幫助我的，搭救我的； 耶和華啊，求你不要耽延！
PS|71|1|耶和華啊，我投靠你， 求你叫我永不羞愧！
PS|71|2|求你憑你的公義搭救我，救拔我； 側耳聽我，拯救我！
PS|71|3|求你作我常來棲身 的磐石， 你已經吩咐要救我， 因為你是我的巖石、我的山寨。
PS|71|4|我的上帝啊，求你救我脫離惡人的手， 脫離不義和殘暴之人的手。
PS|71|5|主耶和華啊，你是我所盼望的； 自我年幼，你是我所倚靠的。
PS|71|6|我自出母胎被你扶持， 使我出母腹的是你。 我要常常讚美你！
PS|71|7|許多人看我為異類， 但你是我堅固的避難所。
PS|71|8|我要滿口述說讚美你的話 終日榮耀你。
PS|71|9|我年老的時候，求你不要丟棄我！ 我體力衰弱時，求你不要離棄我！
PS|71|10|我的仇敵議論我， 那些窺探要害我命的一同商議，
PS|71|11|說：「上帝已經離棄他； 你們去追趕他，捉拿他吧！ 因為沒有人搭救。」
PS|71|12|上帝啊，求你不要遠離我！ 我的上帝啊，求你速速幫助我！
PS|71|13|願那與我為敵的，羞愧滅亡； 願那謀害我的，受辱蒙羞。
PS|71|14|我卻要常常仰望， 並要越發讚美你。
PS|71|15|我的口要終日述說你的公義和你的救恩， 因我無從計算其數。
PS|71|16|我要述說主耶和華的大能， 我單要提說你的公義。
PS|71|17|上帝啊，自我年幼，你就教導我； 直到如今，我傳揚你奇妙的作為。
PS|71|18|上帝啊，我年老髮白的時候， 求你不要離棄我！ 等我宣揚你的能力給下一代， 宣揚你的大能給後世的人。
PS|71|19|上帝啊，你的公義極高； 行過大事的上帝啊，誰能像你？
PS|71|20|你是叫我多經歷重大急難的， 必使我再活過來， 從地的深處救我上來。
PS|71|21|你必使我越發昌大， 又轉來安慰我。
PS|71|22|我的上帝啊，我要鼓瑟稱謝你， 稱謝你的信實！ 以色列 的聖者啊，我要彈琴歌頌你！
PS|71|23|我歌頌你的時候，我的嘴唇要歡呼； 我的性命，就是你所救贖的，也要歡呼。
PS|71|24|我的舌頭也必終日講論你的公義， 因為那些謀害我的人已經蒙羞受辱了。
PS|72|1|上帝啊，求你將你的公平賜給王， 將你的公義賜給王的兒子。
PS|72|2|使他按公義審判你的子民， 按公平審判你的困苦人。
PS|72|3|大山小山都要因公義 使百姓得享平安。
PS|72|4|他必為百姓中困苦的人伸冤， 拯救貧窮之輩， 壓碎那欺壓人的人。
PS|72|5|太陽還存，月亮猶在， 人要敬畏你 ，直到萬代！
PS|72|6|他必降臨，像雨降在已割的草地上， 如甘霖滋潤田地。
PS|72|7|在他的日子，公義 要興旺， 大有平安，除非月亮不在。
PS|72|8|他要執掌權柄，從這海直到那海， 從 大河 直到地極。
PS|72|9|住在曠野的必在他面前下拜， 他的仇敵必要舔土。
PS|72|10|他施 和海島的王要進貢， 示巴 和 西巴 的王要獻禮物。
PS|72|11|眾王都要叩拜他， 萬國都要事奉他。
PS|72|12|貧窮人呼求，他要搭救， 無人幫助的困苦人，他也搭救。
PS|72|13|他要憐憫貧寒和貧窮的人， 拯救貧窮人的性命。
PS|72|14|他要救贖他們脫離欺壓和殘暴， 他們的血在他眼中看為寶貴。
PS|72|15|願他永遠活著， 示巴 的金子要獻給他； 願人常常為他禱告，終日祝福他。
PS|72|16|在地的山頂上，願五穀茂盛， 所結的穀實響動，如 黎巴嫩 的樹林； 願城裏的人興旺，如地上的草。
PS|72|17|願他的名存到永遠， 他的名如太陽之長久 ； 願人因他蒙福， 萬國稱他為有福。
PS|72|18|惟獨耶和華－ 以色列 的上帝能行奇事， 他是應當稱頌的！
PS|72|19|他榮耀的名也當稱頌，直到永遠。 願他的榮耀充滿全地！ 阿們！阿們！
PS|72|20|耶西 的兒子－ 大衛 的祈禱完畢。 亞薩的詩。
PS|73|1|上帝實在恩待 以色列 那些清心的人！
PS|73|2|至於我，我的腳幾乎失閃， 我的步伐險些走偏；
PS|73|3|因為我嫉妒狂傲的人， 我看見惡人享平安。
PS|73|4|他們的力氣強壯， 他們死的時候也沒有疼痛。
PS|73|5|他們不像別人受苦， 也不像別人遭災。
PS|73|6|所以，驕傲如鏈子戴在他們項上， 殘暴像衣裳覆蓋在他們身上。
PS|73|7|他們的眼睛 因體胖而凸出， 他們的內心放任不羈 。
PS|73|8|他們譏笑人，憑惡意說欺壓人的話。 他們說話自高；
PS|73|9|他們的口褻瀆上天， 他們的舌毀謗全地。
PS|73|10|所以他的百姓歸到這裏， 享受滿杯的水 。
PS|73|11|他們說：「上帝怎能曉得？ 至高者哪會知道呢？」
PS|73|12|看哪，這就是惡人， 他們常享安逸，財寶增多。
PS|73|13|我實在徒然潔淨了我的心， 徒然洗手表明我的無辜，
PS|73|14|因為我終日遭災難， 每日早晨受懲治。
PS|73|15|我若說「我要這樣講」， 就是愧對這世代的眾兒女了。
PS|73|16|我思索要明白這事， 眼看實係為難，
PS|73|17|直到我進了上帝的聖所， 思想他們的結局。
PS|73|18|你實在把他們安放在滑地， 使他們跌倒滅亡；
PS|73|19|他們轉眼之間成了何等荒涼！ 他們被驚恐滅盡了。
PS|73|20|人睡醒了，怎樣看夢， 主啊，你醒了也必照樣輕看他們的影像。
PS|73|21|因此，我心裏苦惱， 肺腑被刺。
PS|73|22|我這樣愚昧無知， 在你面前如同畜牲。
PS|73|23|然而，我常與你同在； 你攙扶我的右手。
PS|73|24|你要以你的訓言引導我， 以後你必接我到榮耀裏。
PS|73|25|除你以外，在天上我有誰呢？ 除你以外，在地上我也沒有所愛慕的。
PS|73|26|我的肉體和我的心腸衰殘； 但上帝是我心裏的力量， 又是我的福分，直到永遠。
PS|73|27|看哪，遠離你的，必要死亡； 凡離棄你行淫的，你都滅絕了。
PS|73|28|但我親近上帝是於我有益； 我以主耶和華為我的避難所， 好叫我述說你一切的作為。
PS|74|1|上帝啊，你為何永遠丟棄我們呢？ 為何向你草場的羊發怒，如煙冒出呢？
PS|74|2|求你記念你古時得來的會眾， 就是你所贖、作你產業支派的， 並記念你向來居住的 錫安山 。
PS|74|3|求你舉步去看那日久荒涼之地， 看仇敵在聖所中所做的一切惡事。
PS|74|4|你的敵人在你會中吼叫， 他們豎起自己的標幟為記號，
PS|74|5|好像人揚起斧子 對著林中的樹，
PS|74|6|現在將聖所中的雕刻 ， 全都用斧子錘子打壞。
PS|74|7|他們用火焚燒你的聖所， 褻瀆你名的居所於地。
PS|74|8|他們心裏說「我們要盡行毀滅」； 就在遍地燒燬敬拜上帝聚會的所在。
PS|74|9|我們看不見自己的標幟，不再有先知， 我們當中也無人知道這災禍要到幾時。
PS|74|10|上帝啊，敵人辱罵要到幾時呢？ 仇敵藐視你的名要到永遠嗎？
PS|74|11|你為甚麼縮回你的右手？ 求你從懷中伸出手來，毀滅他們。
PS|74|12|上帝自古以來是我的王， 在這地上施行拯救。
PS|74|13|你曾用能力將海分開， 你打破水裏大魚的頭。
PS|74|14|你曾壓碎 力威亞探 的頭， 把牠給曠野的禽獸作食物。
PS|74|15|你曾分裂泉源和溪流； 使長流的江河枯乾。
PS|74|16|白晝屬你，黑夜也屬你； 亮光和太陽是你預備的。
PS|74|17|地的一切疆界是你立的， 夏天和冬天是你定的。
PS|74|18|耶和華啊，仇敵辱罵，愚頑之輩藐視你的名； 求你記念這事。
PS|74|19|不要將屬你的斑鳩 交給野獸， 不要永遠忘記你困苦人的性命。
PS|74|20|求你顧念所立的約， 因為地上黑暗之處遍滿了兇暴。
PS|74|21|不要讓受欺壓的人蒙羞回去； 要使困苦貧窮的人讚美你的名。
PS|74|22|上帝啊，求你起來為自己辯護！ 求你記念愚頑人怎樣終日辱罵你。
PS|74|23|不要忘記你敵人的喧鬧， 就是那時常上升、起來對抗你之人的喧嘩。
PS|75|1|上帝啊，我們稱謝你，我們稱謝你！ 你的名臨近，人 都述說你奇妙的作為。
PS|75|2|我選定了日期， 必按正直施行審判。
PS|75|3|地和其上的居民都熔化了； 我親自堅立地的柱子。（細拉）
PS|75|4|我對狂傲的人說：「不要狂傲！」 對兇惡的人說：「不要舉角！」
PS|75|5|不要把你們的角高舉， 不要挺著頸項 說話。
PS|75|6|因為高舉非從東，非從西， 也非從南而來。
PS|75|7|惟有上帝斷定， 他使這人降卑，使那人升高。
PS|75|8|耶和華的手裏有杯， 杯內滿了調和起沫的酒； 他倒出來， 地上的惡人都必喝，直到喝盡它的渣滓。
PS|75|9|但我要宣揚，直到永遠！ 我要歌頌 雅各 的上帝！
PS|75|10|惡人一切的角，我要砍斷； 惟有義人的角必被高舉。
PS|76|1|在 猶大 ，上帝為人所認識； 在 以色列 ，他的名為大。
PS|76|2|在 撒冷 有他的住處， 在 錫安 有他的居所。
PS|76|3|他在那裏折斷弓上的火箭、 盾牌、刀劍和戰爭的兵器。（細拉）
PS|76|4|你是光榮的， 比獵物 之山更威嚴。
PS|76|5|心中勇敢的人都被掠奪； 他們睡了長覺，沒有一個英雄能措手。
PS|76|6|雅各 的上帝啊，你的斥責一發， 戰車和戰馬都沉睡了。
PS|76|7|你，惟獨你是可畏的！ 你的怒氣一發，誰能在你面前站得住呢？
PS|76|8|你從天上使人聽判斷。 上帝起來施行審判， 要救地上所有困苦的人； 那時地就懼怕而靜默。（細拉）
PS|76|9|
PS|76|10|人的憤怒終必稱謝你， 你要以人的餘怒束腰。
PS|76|11|你們當向耶和華－你們的上帝許願，還願； 在他四圍的人都當拿貢物獻給那可畏的主。
PS|76|12|他要挫折王子的驕氣， 向地上的君王顯為可畏。
PS|77|1|我要向上帝發聲呼求； 我向上帝發聲，他必側耳聽我。
PS|77|2|我在患難之日尋求主， 在夜間不住地舉手禱告 ， 我的心不肯受安慰。
PS|77|3|我想念上帝，就煩躁不安； 我沉思默想，心靈發昏。（細拉）
PS|77|4|你使我不能閉眼； 我心煩亂，甚至不能說話。
PS|77|5|我追想古時之日， 上古之年。
PS|77|6|夜間我想起我的歌曲 ， 我的心默想，我的靈仔細省察：
PS|77|7|「難道主要永遠丟棄我， 不再施恩嗎？
PS|77|8|難道他的慈愛永遠窮盡， 他的應許世世廢棄嗎？
PS|77|9|難道上帝忘記施恩， 因發怒就止住他的憐憫嗎？」（細拉）
PS|77|10|我說，至高者右手的能力已改變， 這是我的悲哀。
PS|77|11|我要記念耶和華所做的， 要記念你古時的奇事；
PS|77|12|我要思想你所做的， 默念你的作為。
PS|77|13|上帝啊，你的道是神聖的； 有何神明大如上帝呢？
PS|77|14|你是行奇事的上帝， 你曾在萬民中彰顯能力。
PS|77|15|你曾用膀臂贖了你的子民， 就是 雅各 和 約瑟 的子孫。（細拉）
PS|77|16|上帝啊，眾水見你， 眾水一見你就都驚惶， 深淵也都戰抖。
PS|77|17|密雲倒出水來， 天空發出響聲， 你的箭也飛行四方。
PS|77|18|你的雷聲在旋風之中， 閃電照亮世界， 大地戰抖震動。
PS|77|19|你的道在海中， 你的路在大水之中， 你的腳蹤無人知道。
PS|77|20|你曾藉 摩西 和 亞倫 的手引導你的百姓， 好像領羊群一般。
PS|78|1|我的子民哪，要側耳聽我的訓誨， 豎起耳朵聽我口中的言語。
PS|78|2|我要開口說比喻， 我要解開古時的謎語，
PS|78|3|是我們所聽見、所知道， 我們的祖宗告訴我們的。
PS|78|4|我們不要向子孫隱瞞這些事， 而要將耶和華的美德和他的能力， 並他所行的奇事，述說給後代聽。
PS|78|5|他在 雅各 中立法度， 在 以色列 中設律法； 他吩咐我們的祖宗要傳給子孫，
PS|78|6|使將要生的後代子孫可以曉得。 他們也要起來告訴他們的子孫，
PS|78|7|好讓他們仰望上帝， 不忘記上帝的作為， 惟遵守他的命令；
PS|78|8|不要像他們的祖宗， 是頑梗悖逆、心不堅定， 向上帝心不忠實之輩。
PS|78|9|以法蓮 人帶著兵器，拿著弓， 臨陣之日轉身退後。
PS|78|10|他們不遵守上帝的約， 不肯照他的律法行；
PS|78|11|又忘記他的作為 和他所彰顯的奇事。
PS|78|12|他在 埃及 地，在 瑣安 田， 在他們祖宗眼前施行奇事。
PS|78|13|他把海分開，使他們過去， 又叫水立起如壘。
PS|78|14|他白日用雲彩， 終夜用火光引導他們。
PS|78|15|他在曠野使磐石裂開， 多多地給他們水喝，如從深淵而出。
PS|78|16|他使水從磐石湧出， 叫水如江河下流。
PS|78|17|他們卻仍舊得罪他， 在乾旱之地悖逆至高者。
PS|78|18|他們心中試探上帝， 隨自己所欲的求食物，
PS|78|19|並且妄論上帝說： 「上帝豈能在曠野擺設筵席嗎？
PS|78|20|他雖曾擊打磐石，使水湧出，如江河氾濫； 他還能賜糧食嗎？ 還能為他的百姓預備吃的肉嗎？」
PS|78|21|所以，耶和華聽見就發怒， 有烈火向 雅各 點燃， 有怒氣向 以色列 上騰；
PS|78|22|因為他們不信服上帝， 不倚賴他的拯救。
PS|78|23|然而他卻吩咐天空， 又敞開天上的門，
PS|78|24|降嗎哪像雨，給他們吃， 將天上的糧食賜給他們。
PS|78|25|各人就吃大能者的食物； 他賜下糧食，使他們飽足。
PS|78|26|他令東風吹在天空， 用能力引來南風。
PS|78|27|他降肉像雨，多如塵土， 降飛鳥，多如海沙，
PS|78|28|落在他自己的營中， 在他帳幕的四周圍。
PS|78|29|他們吃了，而且飽足； 這樣就隨了他們所欲的。
PS|78|30|但在他們滿足食慾以前， 食物還在他們口中的時候，
PS|78|31|上帝的怒氣就向他們上騰， 殺了他們當中肥壯的人， 打倒 以色列 的青年。
PS|78|32|雖是這樣，他們仍舊犯罪， 不信他奇妙的作為。
PS|78|33|因此，他使他們的日子全歸虛空， 叫他們的年歲盡屬驚恐。
PS|78|34|他殺他們的時候，他們才求問他， 回心轉意，切切尋求上帝。
PS|78|35|他們追念上帝是他們的磐石， 至高的上帝是他們的救贖主。
PS|78|36|他們卻用口諂媚他， 用舌向他說謊。
PS|78|37|他們的心向他不堅定， 不忠於他的約。
PS|78|38|但他有憐憫， 赦免他們的罪孽， 沒有滅絕他們， 而且屢次撤銷他的怒氣， 不發盡他的憤怒。
PS|78|39|他想念他們不過是血肉之軀， 是一陣去而不返的風。
PS|78|40|他們在曠野悖逆他， 在荒地令他擔憂，何其多呢！
PS|78|41|他們再三試探上帝， 惹動 以色列 的聖者。
PS|78|42|他們不追念他手的能力， 和他救贖他們脫離敵人的日子；
PS|78|43|他怎樣在 埃及 顯神蹟， 在 瑣安 田顯奇事，
PS|78|44|把江河並河汊的水都變為血， 使他們不能喝。
PS|78|45|他使蒼蠅成群落在他們當中，吃盡他們， 又叫青蛙滅了他們，
PS|78|46|將他們的果實交給螞蚱， 把他們勞碌得來的交給蝗蟲。
PS|78|47|他降冰雹打壞他們的葡萄樹， 下寒霜打壞他們的桑樹，
PS|78|48|將他們的牲畜交給冰雹， 把他們的群畜交給閃電。
PS|78|49|他使猛烈的怒氣和憤怒、惱恨、苦難， 成了一群降災的使者，臨到他們。
PS|78|50|他為自己的怒氣修平了路， 將他們的性命交給瘟疫， 使他們死亡，
PS|78|51|在 埃及 擊殺所有的長子， 在 含 的帳棚中擊殺他們壯年時頭生的。
PS|78|52|他卻領出自己的子民如羊， 在曠野引導他們如羊群。
PS|78|53|他領他們穩穩妥妥地，使他們不致害怕； 海卻淹沒他們的仇敵。
PS|78|54|他帶他們到自己聖地的邊界， 到他右手所得的這山地。
PS|78|55|他在他們面前趕出外邦人， 用繩子抽籤量地給他們為業， 讓 以色列 支派的人住在自己的帳棚裏。
PS|78|56|他們仍舊試探，悖逆至高的上帝， 不遵守他的法度，
PS|78|57|反倒退後，行詭詐，像他們的祖宗一樣， 他們翻轉，如同鬆弛的弓，
PS|78|58|以丘壇惹他發怒， 以雕刻的偶像使他忌恨。
PS|78|59|上帝聽見就發怒， 全然棄絕了 以色列 ，
PS|78|60|甚至離棄 示羅 的帳幕， 就是他在人間所搭的帳棚；
PS|78|61|又將他有能力的約櫃 交給人擄去， 將他的榮耀交在敵人手中；
PS|78|62|並將他的百姓交給刀劍， 向他的產業發怒。
PS|78|63|壯丁被火燒滅， 童女也無婚禮頌歌。
PS|78|64|祭司倒在刀下， 寡婦卻不哀哭。
PS|78|65|那時，主像睡覺的人醒來， 如勇士飲酒呼喊。
PS|78|66|他擊退敵人， 叫他們永蒙羞辱。
PS|78|67|他撇棄 約瑟 的帳棚， 不揀選 以法蓮 支派，
PS|78|68|卻揀選 猶大 支派， 揀選他所喜愛的 錫安山 ；
PS|78|69|建造他的聖所如同高峰， 又像他所建立的永存之地。
PS|78|70|他揀選他的僕人 大衛 ， 從羊圈中將他召來，
PS|78|71|叫他不再牧放那些母羊， 為要牧養自己的百姓 雅各 和自己的產業 以色列 。
PS|78|72|於是，他以純正的心牧養他們， 用巧妙的手引導他們。
PS|79|1|上帝啊，外邦人侵犯你的產業， 玷污你的聖殿，使 耶路撒冷 變成廢墟，
PS|79|2|將你僕人的屍首交給天空的飛鳥為食， 把你聖民的肉交給地上的走獸，
PS|79|3|耶路撒冷 的周圍流出他們的血如水， 無人埋葬。
PS|79|4|我們成為鄰國羞辱的對象， 被四圍的人嗤笑譏刺。
PS|79|5|耶和華啊，你發怒要到幾時呢？ 要到永遠嗎？ 你的忌恨要如火焚燒嗎？
PS|79|6|求你將你的憤怒傾倒在那不認識你的萬邦 和那不求告你名的國度。
PS|79|7|因為他們吞了 雅各 ， 將他的住處變為廢墟。
PS|79|8|求你不要記得我們先前世代的罪孽； 願你的憐憫速速臨到我們， 因為我們落到極卑微的地步。
PS|79|9|拯救我們的上帝啊，求你因你名的榮耀幫助我們！ 為你名的緣故搭救我們，赦免我們的罪。
PS|79|10|為何讓列國說「他們的上帝在哪裏」呢？ 求你讓列國知道， 你在我們眼前伸你僕人流血的冤。
PS|79|11|願被囚之人的嘆息達到你面前， 求你以強大的膀臂存留那些將死的人。
PS|79|12|主啊，求你將我們鄰邦所加給你的羞辱 七倍歸到他們身上。
PS|79|13|這樣，你的子民，你草場的羊， 要稱謝你，直到永遠； 要述說讚美你的話，直到萬代。
PS|80|1|領 約瑟 如領羊群的 以色列 牧者啊，求你側耳而聽！ 在基路伯之上坐寶座的啊，求你發出光來！
PS|80|2|在 以法蓮 、 便雅憫 、 瑪拿西 面前 求你施展你的大能，拯救我們。
PS|80|3|上帝啊，求你使我們回轉 ， 使你的臉發光，我們就會得救！
PS|80|4|耶和華─萬軍之上帝啊， 你因你百姓的禱告發怒，要到幾時呢？
PS|80|5|你以眼淚當食物給他們吃， 量出滿碗的眼淚給他們喝。
PS|80|6|你使鄰邦因我們紛爭， 我們的仇敵彼此戲笑。
PS|80|7|萬軍之上帝啊，求你使我們回轉， 使你的臉發光，我們就會得救！
PS|80|8|你從 埃及 拔出一棵葡萄樹， 趕出外邦人，把這樹栽上。
PS|80|9|你在它面前清除雜物， 它就深深扎根，蔓延滿地。
PS|80|10|它的影子遮蔽群山， 枝子好像高大的香柏樹。
PS|80|11|它長出枝子，直到大海， 伸展嫩枝，延到 大河 。
PS|80|12|你為何拆毀這樹的籬笆， 任憑路人摘取？
PS|80|13|林中的野豬踐踏它， 田裏的走獸吞吃它。
PS|80|14|萬軍之上帝啊，求你轉回， 從天上垂看觀察，眷顧這葡萄樹；
PS|80|15|保護你右手所栽的根， 你為自己所堅固的幼苗。
PS|80|16|這樹已經被火焚燒，被刀砍伐， 因你臉上的怒容就滅亡了。
PS|80|17|願你的手扶持你右邊的人， 你為自己所堅固的人子。
PS|80|18|這樣，我們就不背離你； 求你救活我們，讓我們得以求告你的名。
PS|80|19|耶和華─萬軍之上帝啊，求你使我們回轉， 使你的臉發光，我們就會得救！
PS|81|1|你們當向上帝－我們的力量大聲歌唱， 向 雅各 的上帝歡呼！
PS|81|2|高唱詩歌，擊打手鼓， 彈奏悅耳的琴瑟。
PS|81|3|當在新月和滿月－ 我們過節的日期吹角，
PS|81|4|因這是為 以色列 所定的律例， 是 雅各 上帝的典章。
PS|81|5|他攻擊 埃及 地的時候， 曾立此為 約瑟 的法度。 我聽見我所不明白的語言：
PS|81|6|「我使你 的肩頭得脫重擔， 使你的手放下筐子。
PS|81|7|你在急難中呼求，我就搭救你， 在雷的隱密處應允你， 在 米利巴 水那裏考驗你。（細拉）
PS|81|8|聽啊，我的子民，我要勸戒你； 以色列 啊，我真願你肯聽從我。
PS|81|9|在你當中，不可有外族的神明； 外邦的神明，你也不可下拜。
PS|81|10|我是耶和華－你的上帝， 曾將你從 埃及 地領上來； 你要大大張口，我就使你滿足。
PS|81|11|「無奈，我的子民不聽我的聲音， 以色列 不肯聽從我。
PS|81|12|我就任憑他們心裏頑梗， 隨自己的計謀而行。
PS|81|13|我的子民若肯聽從我， 以色列 肯行我的道，
PS|81|14|我就速速制伏他們的仇敵， 反手攻擊他們的敵人。
PS|81|15|恨耶和華的人必來投降， 願他們的厄運直到永遠。
PS|81|16|他必拿上好的麥子給 以色列 吃， 又拿磐石出的蜂蜜使你飽足。 」
PS|82|1|上帝站立在神聖的會中， 在諸神中施行審判。
PS|82|2|你們審判不秉公義， 抬舉惡人的臉面，要到幾時呢？（細拉）
PS|82|3|當為貧寒的人和孤兒伸冤， 為困苦和窮乏的人施行公義。
PS|82|4|當保護貧寒和貧窮的人， 救他們脫離惡人的手。
PS|82|5|他們愚昧，他們無知， 在黑暗中走來走去； 地的根基都搖動了。
PS|82|6|我曾說：「你們是諸神， 都是至高者的兒子。
PS|82|7|然而，你們要死去，與世人一樣， 要仆倒，像任何一位王子一般。」
PS|82|8|上帝啊，求你起來審判全地， 因為你必得萬國為業。
PS|83|1|上帝啊，求你不要靜默！ 上帝啊，求你不要閉口，不要不作聲！
PS|83|2|因為你的仇敵喧嚷， 恨你的抬起頭來。
PS|83|3|他們同謀奸詐要害你的百姓， 彼此商議要害你所保護的人。
PS|83|4|他們說：「來吧，我們將他們除滅， 使他們不再成國！ 使 以色列 的名不再被人記念！」
PS|83|5|他們同心商議， 彼此結盟，要抵擋你；
PS|83|6|他們就是住帳棚的 以東 和 以實瑪利 人， 摩押 和 夏甲 人，
PS|83|7|迦巴勒 、 亞捫 、 亞瑪力 、 非利士 和 推羅 的居民。
PS|83|8|亞述 也與他們聯合， 作 羅得 子孫的幫手。（細拉）
PS|83|9|求你待他們，如待 米甸 ， 如在 基順河 待 西西拉 和 耶賓 一樣。
PS|83|10|他們在 隱‧多珥 滅亡， 成了地上的糞土。
PS|83|11|求你使他們的貴族像 俄立 和 西伊伯 ， 使他們的王子都像 西巴 和 撒慕拿 。
PS|83|12|因為他們說：「我們要得上帝的住處， 作自己的產業。」
PS|83|13|我的上帝啊，求你使他們像旋風中的塵土， 如風前的碎秸。
PS|83|14|火怎樣焚燒樹林， 火焰怎樣燒著山嶺，
PS|83|15|求你也照樣用狂風追趕他們， 用暴雨恐嚇他們。
PS|83|16|耶和華啊，求你使他們滿面羞恥， 好叫他們尋求你的名！
PS|83|17|願他們永遠羞愧驚惶！ 願他們慚愧滅亡！
PS|83|18|願他們認識你的名是耶和華， 惟獨你是掌管全地的至高者！
PS|84|1|萬軍之耶和華啊， 你的居所何等可愛！
PS|84|2|我羨慕渴想耶和華的院宇， 我的內心，我的肉體向永生上帝歡呼。
PS|84|3|萬軍之耶和華－我的王，我的上帝啊， 在你祭壇那裏，麻雀為自己找到了家， 燕子為自己找著菢雛之窩。
PS|84|4|如此住在你殿中的有福了！ 他們不斷地讚美你。（細拉）
PS|84|5|靠你有力量、心中嚮往 錫安 大道的， 這人有福了！
PS|84|6|他們經過「流淚谷」 ，叫這谷變為泉源之地； 且有秋雨之福蓋滿了全谷。
PS|84|7|他們行走，力上加力， 各人到 錫安 朝見上帝。
PS|84|8|萬軍之耶和華上帝啊，求你聽我的禱告！ 雅各 的上帝啊，求你側耳而聽！（細拉）
PS|84|9|上帝啊，我們的盾牌，求你觀看， 求你垂顧你受膏者的面！
PS|84|10|在你的院宇一日， 勝似千日； 寧可在我上帝的殿中看門， 不願住在惡人的帳棚裏。
PS|84|11|因為耶和華上帝是太陽，是盾牌， 耶和華要賜下恩惠和榮耀。 他未嘗留下福氣不給那些行動正直的人。
PS|84|12|萬軍之耶和華啊， 倚靠你的人有福了！
PS|85|1|耶和華啊，你已經向你的地施恩， 救回被擄的 雅各 。
PS|85|2|你赦免了你百姓的罪孽， 遮蓋了他們一切的過犯。（細拉）
PS|85|3|你收回所發的憤怒， 撤銷你猛烈的怒氣。
PS|85|4|拯救我們的上帝啊，求你使我們回轉， 使你向我們所發的憤怒止息。
PS|85|5|你要向我們發怒到永遠嗎？ 要將你的怒氣延留到萬代嗎？
PS|85|6|你不再將我們救活， 使你的百姓因你歡喜嗎？
PS|85|7|耶和華啊，求你使我們得見你的慈愛， 又將你的救恩賜給我們。
PS|85|8|我要聽上帝－耶和華所說的話， 因為他必應許賜平安給他的百姓，就是他的聖民； 他們卻不可再轉向愚昧 。
PS|85|9|他的救恩誠然與敬畏他的人相近， 使榮耀住在我們的地上。
PS|85|10|慈愛和誠實彼此相遇， 公義與和平彼此相親。
PS|85|11|誠實從地而生， 公義從天而現。
PS|85|12|耶和華必賜福氣給我們； 我們的地也要出土產。
PS|85|13|公義要行在他面前， 使他的腳蹤有可走之路。
PS|86|1|耶和華啊，求你側耳應允我， 因我是困苦貧窮的。
PS|86|2|求你保住我的性命，因我是虔誠的人。 我的上帝啊，求你拯救我這倚靠你的僕人！
PS|86|3|主啊，求你憐憫我， 因我終日求告你。
PS|86|4|主啊，求你使你的僕人心裏歡喜， 因為我的心仰望你。
PS|86|5|主啊，你本為良善，樂於饒恕人， 以豐盛的慈愛對待凡求告你的人。
PS|86|6|耶和華啊，求你側耳聽我的禱告， 留心聽我懇求的聲音。
PS|86|7|我在患難之日要求告你， 因為你必應允我。
PS|86|8|主啊，諸神之中沒有可與你相比的， 你的作為也無以為比。
PS|86|9|主啊，你所造的萬民都要來敬拜你， 他們要榮耀你的名。
PS|86|10|因你本為大，且行奇妙的事， 惟獨你是上帝。
PS|86|11|耶和華啊，求你將你的道指教我， 我要照你的真理而行； 求你使我專心敬畏你的名！
PS|86|12|主－我的上帝啊，我要一心稱謝你； 我要榮耀你的名，直到永遠。
PS|86|13|因為你的慈愛在我身上浩大， 你救了我的性命免入陰間的深處。
PS|86|14|上帝啊，驕傲的人起來攻擊我， 又有一群強橫的人尋索我的命； 他們沒有將你放在眼裏。
PS|86|15|主啊，你是有憐憫，有恩惠的上帝， 不輕易發怒，並有豐盛的慈愛和信實。
PS|86|16|求你轉向我，憐憫我， 將你的力量賜給僕人，拯救你使女的兒子。
PS|86|17|求你向我顯出恩待我的憑據， 使恨我的人看見就羞愧， 因為你－耶和華幫助我，安慰了我。
PS|87|1|耶和華所立的根基在聖山上。
PS|87|2|耶和華愛 錫安 的門， 勝於愛 雅各 一切的住處。
PS|87|3|上帝的城啊， 有榮耀的事是指著你說的。（細拉）
PS|87|4|我要提起 拉哈伯 和 巴比倫 人， 是在認識我之中的； 看哪， 非利士 、 推羅 和 古實 人， 個個生在那裏。
PS|87|5|論到 錫安 ，必有話說： 「這一個、那一個都生在其中」； 而且至高者必親自堅立這城。
PS|87|6|當耶和華記錄萬民的時候， 他要寫出人的出生地。（細拉）
PS|87|7|歌唱的、跳舞的，都要說： 「我的泉源都在你裏面。」
PS|88|1|耶和華－拯救我的上帝啊， 我晝夜在你面前呼求；
PS|88|2|願我的禱告達到你面前， 求你側耳聽我的懇求！
PS|88|3|因為我心裏滿了患難， 我的性命臨近陰間；
PS|88|4|我與下到地府的人同列， 如同無人幫助的人一樣。
PS|88|5|我被丟在死人中， 好像被殺的人躺在墳墓裏， 不再被你記得， 與你的手隔絕了。
PS|88|6|你把我放在極深的地府裏， 在黑暗地，在深處。
PS|88|7|你的憤怒重壓我身， 你用一切的波浪困住我。（細拉）
PS|88|8|你把我所認識的人隔在遠處， 使我為他們所憎惡； 我被拘禁，不能出來。
PS|88|9|我的眼睛因困苦而昏花； 耶和華啊，我天天求告你，向你舉手。
PS|88|10|你豈要行奇事給死人看嗎？ 陰魂還能起來稱謝你嗎？（細拉）
PS|88|11|你的慈愛豈能在墳墓裏被人述說嗎？ 你的信實豈能在冥府 被人傳揚嗎？
PS|88|12|你的奇事豈能在幽暗裏為人所知嗎？ 你的公義豈能在遺忘之地為人所識嗎？
PS|88|13|耶和華啊，至於我，我要呼求你； 每早晨，我的禱告要達到你面前。
PS|88|14|耶和華啊，你為何丟棄我？ 為何轉臉不顧我？
PS|88|15|我自幼受苦，幾乎死亡； 你使我驚恐，煩亂不安。
PS|88|16|你的烈怒漫過我身， 你用驚嚇把我除滅。
PS|88|17|這些如水終日環繞我， 一起圍困我。
PS|88|18|你把我的良朋密友隔在遠處， 使我所認識的人都在黑暗裏 。
PS|89|1|我要歌唱耶和華的慈愛，直到永遠， 我要用口將你的信實傳到萬代。
PS|89|2|因我曾說：「你的慈愛必建立到永遠， 你的信實必堅立在天上。」
PS|89|3|「我與我所揀選的人立了約， 向我的僕人 大衛 起了誓：
PS|89|4|『我要堅立你的後裔，直到永遠， 要建立你的寶座，直到萬代。』」（細拉）
PS|89|5|耶和華啊，諸天要稱謝你的奇事； 在聖者的會中，要稱謝你的信實。
PS|89|6|因在天空誰能比耶和華呢？ 諸神之中，誰能像耶和華呢？
PS|89|7|在聖者的會中，他是大有威嚴的上帝， 比在他四圍所有的更可畏懼。
PS|89|8|耶和華－萬軍之上帝啊， 哪一個大能者像耶和華？ 你的信實在你四圍。
PS|89|9|你管轄海的狂傲； 波浪翻騰，你使它平靜了。
PS|89|10|你打碎了 拉哈伯 ，使牠如遭刺殺的人； 你用大能的膀臂打散了你的仇敵。
PS|89|11|天屬你，地也屬你； 世界和其中所充滿的都為你所建立。
PS|89|12|南北為你所創造； 他泊 和 黑門 都因你的名歡呼。
PS|89|13|你有大能的膀臂， 你的手有力，你的右手也高舉。
PS|89|14|公義和公平是你寶座的根基， 慈愛和信實行在你前面。
PS|89|15|知道向你歡呼的，那民有福了！ 耶和華啊，他們要行走在你臉的光中。
PS|89|16|他們因你的名終日歡樂， 因你的公義得以高舉。
PS|89|17|你是他們力量的榮耀。 我們的角必被高舉，因為你喜愛我們。
PS|89|18|我們的盾牌是耶和華， 我們的王是 以色列 的聖者。
PS|89|19|當時，你在異象中吩咐你的聖民，說： 「我已把救助之力加在壯士身上， 高舉了那從百姓中所揀選的人。
PS|89|20|我尋得我的僕人 大衛 ， 用我的聖膏膏他。
PS|89|21|我的手必使他堅立， 我的膀臂也必堅固他。
PS|89|22|仇敵必不勒索他， 兇惡之子也不苦害他。
PS|89|23|我要在他面前打碎他的敵人， 擊殺那些恨他的人。
PS|89|24|我的信實和我的慈愛要與他同在； 因我的名，他的角必被高舉。
PS|89|25|我要使他的手伸到海上， 右手伸到河上。
PS|89|26|他要稱呼我說：『你是我的父， 是我的上帝，是拯救我的磐石。』
PS|89|27|我也要立他為長子， 為世上最高的君王。
PS|89|28|我要為他存留我的慈愛，直到永遠， 我與他所立的約必堅定不移。
PS|89|29|我也要使他的後裔存到永遠， 使他的寶座如天之久。
PS|89|30|「倘若他的子孫離棄我的律法， 不照我的典章行，
PS|89|31|背棄我的律例， 不遵守我的誡命，
PS|89|32|我就要用杖責罰他們的過犯， 用鞭責罰他們的罪孽。
PS|89|33|只是我不將我的慈愛全然收回， 也不叫我的信實廢除。
PS|89|34|我必不毀損我的約， 也不改變我口中所出的話。
PS|89|35|我僅此一次指著自己的神聖起誓， 我絕不向 大衛 說謊！
PS|89|36|他的後裔要存到永遠， 他的寶座在我面前如太陽，
PS|89|37|又如月亮永遠堅立； 天上的見證是確實的。」（細拉）
PS|89|38|但你惱怒你的受膏者， 拒絕他，離棄了他。
PS|89|39|你厭惡與你僕人所立的約， 將他的冠冕踐踏於地。
PS|89|40|你拆毀了他一切的圍牆， 使他的堡壘變為廢墟。
PS|89|41|過路的人都搶奪他， 他成了鄰邦羞辱的對象。
PS|89|42|你高舉了他敵人的右手， 使他所有的仇敵歡喜。
PS|89|43|你叫他的刀劍捲刃， 使他在戰爭中站立不住。
PS|89|44|你使他的光輝止息， 將他的寶座推倒於地。
PS|89|45|你減少他年輕的日子， 又使他蒙羞。（細拉）
PS|89|46|耶和華啊，這要到幾時呢？ 你要隱藏自己到永遠嗎？ 你的憤怒如火焚燒要到幾時呢？
PS|89|47|求你想念我的生命是何等短暫。 你創造世人，要使他們歸於何等的虛空呢？
PS|89|48|誰能常活不見死亡、 救自己脫離陰間的掌控呢？（細拉）
PS|89|49|主啊，你從前憑你的信實 向 大衛 起誓要施行的慈愛在哪裏呢？
PS|89|50|主啊，求你記念僕人們所受的羞辱， 記念我怎樣將萬族所加的羞辱都放在我的胸懷。
PS|89|51|耶和華啊，這是你仇敵所加的羞辱， 羞辱了你受膏者的腳蹤。
PS|89|52|耶和華是應當稱頌的，直到永遠。 阿們！阿們！ 神人摩西的祈禱。
PS|90|1|主啊，你世世代代作我們的居所。
PS|90|2|諸山未曾生出， 地與世界你未曾造成， 從亙古到永遠，你是上帝。
PS|90|3|你使人歸於塵土，說： 「世人哪，你們要歸回。」
PS|90|4|在你看來，千年如已過的昨日， 又如夜間的一更。
PS|90|5|你叫他們如水沖去， 他們如睡一覺。 早晨，他們如生長的草；
PS|90|6|早晨發芽生長， 晚上割下枯乾。
PS|90|7|我們因你的怒氣而消滅， 因你的憤怒而驚惶。
PS|90|8|你將我們的罪孽擺在你面前， 將我們的隱惡擺在你面光之中。
PS|90|9|我們經過的日子，都在你震怒之下， 我們度盡的年歲，好像一聲嘆息。
PS|90|10|我們一生的年日是七十歲， 若是強壯可到八十歲； 但其中所矜誇的不過是勞苦愁煩， 轉眼即逝，我們便如飛而去。
PS|90|11|誰曉得你怒氣的權勢？ 誰因著敬畏你而曉得你的憤怒呢？
PS|90|12|求你指教我們怎樣數算自己的日子， 好叫我們得著智慧的心。
PS|90|13|耶和華啊，我們要等到幾時呢？ 求你轉回，憐憫你的僕人們。
PS|90|14|求你使我們早早飽得你的慈愛， 好叫我們一生一世歡呼喜樂。
PS|90|15|求你照著你使我們受苦的日子， 和我們遭難的年歲，使我們喜樂。
PS|90|16|願你的作為向你僕人們顯現， 願你的榮耀向他們子孫顯明。
PS|90|17|願主－我們上帝的恩寵歸於我們身上。 願你堅立我們手所做的工， 我們手所做的工，願你堅立。
PS|91|1|住在至高者隱密處的， 必住在全能者的蔭下。
PS|91|2|我要向耶和華說： 「我的避難所、我的山寨、 我的上帝，你是我所倚靠的。」
PS|91|3|他必救你脫離捕鳥者的羅網 和毀滅人的瘟疫。
PS|91|4|他必用自己的翎毛遮蔽你； 你要投靠在他翅膀底下， 他的信實是大小的盾牌。
PS|91|5|你必不怕黑夜的驚駭， 或是白日飛的箭，
PS|91|6|也不怕黑夜流行的瘟疫， 或是午間滅人的災害。
PS|91|7|雖有千人仆倒在你旁邊， 萬人仆倒在你右邊， 這災卻不得臨近你。
PS|91|8|你惟親眼觀看， 見惡人遭報。
PS|91|9|因為耶和華是我的避難所， 你以至高者為居所，
PS|91|10|禍患必不臨到你， 災害也不挨近你的帳棚。
PS|91|11|因他要為你命令他的使者， 在你所行的一切道路上保護你。
PS|91|12|他們要用手托住你， 免得你的腳碰在石頭上。
PS|91|13|你要踹踏獅子和毒蛇， 踐踏少壯獅子和大蛇。
PS|91|14|「因為他專心愛我，我要搭救他； 因為他認識我的名，我要把他安置在高處。
PS|91|15|他若求告我，我就應允他； 他在急難中，我與他同在； 我要搭救他，使他尊貴。
PS|91|16|我要使他享足長壽， 將我的救恩顯明給他。」
PS|92|1|這是多麼好啊！ 稱謝耶和華， 歌頌你至高者的名，
PS|92|2|早晨傳揚你的慈愛， 每夜傳揚你的信實。
PS|92|3|用十弦的樂器和瑟， 用琴優雅的聲音；
PS|92|4|因你－耶和華藉著你的作為使我高興， 我要因你手的工作歡呼。
PS|92|5|耶和華啊，你的工作何其大！ 你的心思極其深！
PS|92|6|畜牲一般的人不曉得， 愚昧人也不明白。
PS|92|7|惡人雖茂盛如草， 作惡的人雖全都興旺， 他們卻要滅亡， 直到永遠。
PS|92|8|耶和華啊，惟有你是至高， 直到永遠。
PS|92|9|耶和華啊，看哪，你的仇敵， 看哪，你的仇敵都要滅亡； 作惡的全都要離散。
PS|92|10|你卻高舉了我的角，如野牛的角； 我是被新油膏抹的。
PS|92|11|我的眼睛看見我的仇敵遭報， 我的耳朵聽見那些起來攻擊我的惡人受罰。
PS|92|12|義人要興旺如棕樹， 生長如 黎巴嫩 的香柏樹。
PS|92|13|他們栽於耶和華的殿中， 發旺在我們上帝的院裏。
PS|92|14|他們髮白的時候仍結果子， 而且鮮美多汁，
PS|92|15|好顯明耶和華是正直的； 他是我的磐石，在他毫無不義。
PS|93|1|耶和華作王！ 他以威嚴為衣穿上； 耶和華以能力為衣，以能力束腰， 世界就堅定，不得動搖。
PS|93|2|你的寶座從太初立定， 你從亙古就有。
PS|93|3|耶和華啊，大水揚起， 大水發聲，大水澎湃。
PS|93|4|耶和華在高處大有威力， 勝過諸水的響聲，洋海的大浪。
PS|93|5|耶和華啊，你的法度最為確定； 你的殿宜稱為聖，直到永遠。
PS|94|1|耶和華啊，你是伸冤的上帝； 伸冤的上帝啊，求你發出光來！
PS|94|2|審判世界的主啊，求你挺身而立， 使驕傲的人受應得的報應！
PS|94|3|耶和華啊，惡人誇勝要到幾時呢？ 要到幾時呢？
PS|94|4|他們咆哮，說狂妄的話， 作惡的人全都誇耀自己。
PS|94|5|耶和華啊，他們強壓你的百姓， 苦害你的產業。
PS|94|6|他們殺死寡婦和寄居的人， 又殺害孤兒。
PS|94|7|他們說：「耶和華必不看見， 雅各 的上帝必不留意。」
PS|94|8|百姓中像畜牲一般的人當思想， 你們愚昧人要到幾時才有智慧呢？
PS|94|9|造耳朵的，難道自己聽不見嗎？ 造眼睛的，難道自己看不見嗎？
PS|94|10|管教列國的，就是叫人得知識的， 難道自己不懲治人嗎？
PS|94|11|耶和華知道人的意念是虛妄的。
PS|94|12|耶和華啊，你所管教、 用律法教導的人有福了！
PS|94|13|你使他在遭難的日子仍得平安， 直到為惡人挖好了坑。
PS|94|14|因為耶和華必不丟棄他的百姓， 也不離棄他的產業。
PS|94|15|審判要回復公義， 心裏正直的，都必跟隨它。
PS|94|16|誰肯為我起來攻擊邪惡的？ 誰肯為我站起抵擋作惡的？
PS|94|17|若不是耶和華幫助我， 我早就住在寂靜 之中了。
PS|94|18|我若說：「我失了腳！」 耶和華啊，你的慈愛必扶持我。
PS|94|19|我心裏多憂多疑， 你的安慰使我歡樂。
PS|94|20|那藉著律例玩弄奸惡、 以權位肆行殘害的，豈能與你交往呢？
PS|94|21|他們大家聚集攻擊義人， 將無辜的人定了死罪。
PS|94|22|但耶和華向來作我的碉堡， 我的上帝作了我投靠的磐石。
PS|94|23|他叫他們的罪孽歸到自己身上， 要因他們的邪惡剪除他們； 耶和華－我們的上帝要把他們剪除。
PS|95|1|來啊，我們要向耶和華歌唱， 向拯救我們的磐石歡呼！
PS|95|2|我們要以感謝來到他面前， 用詩歌向他歡呼！
PS|95|3|因耶和華是偉大的上帝， 是超越萬神的大君王。
PS|95|4|地的深處在他手中； 山的高峰也屬他。
PS|95|5|海洋屬他，是他造的； 旱地也是他手造成的。
PS|95|6|來啊，我們要俯伏敬拜， 在造我們的耶和華面前跪拜。
PS|95|7|因為他是我們的上帝； 我們是他草場的百姓，是他手中的羊。 惟願你們今天聽他的話！
PS|95|8|你們不可硬著心，像在 米利巴 ， 就是在曠野 瑪撒 的日子。
PS|95|9|那時，你們的祖宗試我，探我， 並且觀看我的作為。
PS|95|10|四十年之久，我厭煩那世代，說： 「這是心裏迷糊的百姓， 竟不知道我的道路！」
PS|95|11|所以，我在怒中起誓： 「他們斷不可進入我的安息！」
PS|96|1|你們要向耶和華唱新歌！ 全地都要向耶和華歌唱！
PS|96|2|要向耶和華歌唱，稱頌他的名！ 天天傳揚他的救恩！
PS|96|3|在列國中述說他的榮耀！ 在萬民中述說他的奇事！
PS|96|4|因耶和華本為大，當受極大的讚美； 他在萬神之上，當受敬畏。
PS|96|5|因萬民的神明都屬虛無； 惟獨耶和華創造諸天。
PS|96|6|有尊榮和威嚴在他面前， 有能力與華美在他聖所。
PS|96|7|民中的萬族啊，要將榮耀、能力歸給耶和華， 都歸給耶和華！
PS|96|8|要將耶和華的名所當得的榮耀歸給他， 拿供物來進入他的院宇。
PS|96|9|當敬拜神聖榮耀的耶和華 ， 全地都要在他面前戰抖！
PS|96|10|要在列國中說：「耶和華作王了！ 世界堅定，不得動搖； 他要按公正審判萬民。」
PS|96|11|願天歡喜，願地快樂！ 願海和其中所充滿的澎湃！
PS|96|12|願田和其中所有的都歡樂！ 那時，林中的樹木都要在耶和華面前歡呼。
PS|96|13|因為他來了，他來要審判全地。 他要按公義審判世界， 按信實審判萬民。
PS|97|1|耶和華作王！願地快樂！ 願眾海島歡喜！
PS|97|2|密雲和幽暗在他四圍， 公義和公平是他寶座的根基。
PS|97|3|烈火在他前頭行， 燒滅他四圍的敵人。
PS|97|4|他的閃電光照世界， 大地看見就震動。
PS|97|5|諸山見耶和華的面， 就是全地之主的面，就如蠟熔化。
PS|97|6|諸天表明他的公義， 萬民看見他的榮耀。
PS|97|7|願所有事奉雕刻偶像、 靠虛無神明自誇的，都蒙羞愧。 萬神哪，你們都當拜他。
PS|97|8|耶和華啊，因你的判斷， 錫安 聽見就歡喜； 猶大 的城鎮 也都快樂。
PS|97|9|因為你－耶和華至高，超乎全地； 受尊崇，遠超萬神之上。
PS|97|10|你們愛耶和華的，都當恨惡罪惡； 他保護聖民的性命， 搭救他們脫離惡人的手。
PS|97|11|散播亮光是為義人 ， 喜樂歸於心裏正直的人。
PS|97|12|義人哪，你們當靠耶和華歡喜， 當頌揚他神聖的名字 。
PS|98|1|你們要向耶和華唱新歌！ 因為他行過奇妙的事， 他的右手和聖臂施行救恩。
PS|98|2|耶和華顯明了他的救恩， 在列國眼前顯出公義；
PS|98|3|記念他對 以色列 家的慈愛和信實。 地的四極都看見我們上帝的救恩。
PS|98|4|全地都要向耶和華歡呼， 要揚聲，歡唱，歌頌！
PS|98|5|用琴歌頌耶和華， 用琴和詩歌的聲音歌頌他！
PS|98|6|用號筒和角聲， 在大君王耶和華面前歡呼！
PS|98|7|願海和其中所充滿的澎湃， 願世界和住在其間的發聲。
PS|98|8|願大水拍掌， 願諸山在耶和華面前一同歡呼；
PS|98|9|因為他來要審判全地。 他要按公義審判世界， 按公正審判萬民。
PS|99|1|耶和華作王，萬民當戰抖！ 他坐在基路伯的寶座上，地當動搖。
PS|99|2|耶和華在 錫安 為大， 他超越萬民之上。
PS|99|3|願他們頌揚他大而可畏的名， 他本為聖！
PS|99|4|喜愛公平、大能的王啊，你堅立公正， 在 雅各 中施行公平和公義。
PS|99|5|當尊崇耶和華－我們的上帝， 在他腳凳前下拜。 他本為聖！
PS|99|6|在他的祭司中有 摩西 和 亞倫 ， 在求告他名的人中有 撒母耳 。 他們求告耶和華，他就應允他們。
PS|99|7|他在雲柱中向他們說話， 他們遵守他的法度和他所賜給他們的律例。
PS|99|8|耶和華－我們的上帝啊，你應允了他們； 你是赦免他們的上帝， 卻按他們所做的報應他們。
PS|99|9|當尊崇耶和華－我們的上帝， 在他的聖山下拜， 因為耶和華－我們的上帝本為聖！
PS|100|1|普天下當向耶和華歡呼！
PS|100|2|當樂意事奉耶和華， 當歡唱來到他面前！
PS|100|3|當認識耶和華是上帝！ 我們是他造的，也是屬他的； 我們是他的民，是他草場的羊。
PS|100|4|當稱謝進入他的門， 當讚美進入他的院。 當感謝他，稱頌他的名！
PS|100|5|因為耶和華本為善； 他的慈愛存到永遠， 他的信實直到萬代。
PS|101|1|我要歌唱慈愛和公平， 耶和華啊，我要向你歌頌！
PS|101|2|我要用智慧行完全的道。 你幾時到我這裏來呢？ 我要以純正的心行在我家中。
PS|101|3|邪僻的事，我都不擺在我眼前； 悖逆的人所做的事，我甚恨惡， 不容沾在我身上。
PS|101|4|歪曲的心思，我必遠離； 邪惡的事情，我不知道。
PS|101|5|暗中讒害他鄰居的，我必將他滅絕； 眼目高傲、心裏驕縱的，我必不容忍。
PS|101|6|我眼要看顧地上誠實可靠的人，使他們與我同住； 行正直路的，他要侍候我。
PS|101|7|行詭詐的，必不得住在我家裏； 說謊言的，必不得立在我眼前。
PS|101|8|我每日早晨要滅絕地上所有的惡人， 把作惡的從耶和華的城裏全都剪除。
PS|102|1|耶和華啊，求你聽我的禱告， 願我的呼求達到你面前！
PS|102|2|我急難的日子，求你不要轉臉不顧我！ 我呼求的日子，求你向我側耳，快快應允我！
PS|102|3|因為我的年日在煙中消失 ， 我的骨頭如火把燒著。
PS|102|4|我的心如草被踩碎而枯乾， 甚至我忘記吃飯。
PS|102|5|因我嘆息的聲音， 我的肉緊貼骨頭。
PS|102|6|我如同曠野的鵜鶘， 好像荒地的貓頭鷹。
PS|102|7|我清醒難以入眠， 如同房頂上孤單的麻雀。
PS|102|8|我的仇敵整日辱罵我， 向我叫號的人指著我賭咒。
PS|102|9|我吃灰燼如同吃飯， 我喝的有眼淚攙雜。
PS|102|10|這都因你的惱恨和憤怒， 你把我舉起，又把我摔下。
PS|102|11|我的年日如夕陽， 我也如草枯乾。
PS|102|12|惟你－耶和華必永遠坐在寶座上， 你的名 存到萬代。
PS|102|13|你必起來憐憫 錫安 ； 因現在是可憐它的時候， 因所定的日期已經到了。
PS|102|14|你的僕人們喜愛 錫安 的石頭， 憐憫它的塵土。
PS|102|15|列國要敬畏耶和華的名， 地上眾王都要敬畏你的榮耀。
PS|102|16|因為耶和華建造了 錫安 ， 在他的榮耀裏顯現。
PS|102|17|他垂聽窮乏人的禱告， 不藐視他們的祈求。
PS|102|18|這必為後代的人記下， 將來受造的百姓要讚美耶和華。
PS|102|19|因為他從至高的聖所垂看； 耶和華從天向地觀看，
PS|102|20|要垂聽被囚之人的嘆息， 要釋放將死的人，
PS|102|21|使人在 錫安 傳揚耶和華的名， 在 耶路撒冷 傳揚讚美他的話，
PS|102|22|就是在萬民和列國 聚集事奉耶和華的時候。
PS|102|23|他使我的力量半途衰弱， 使我的年日短少。
PS|102|24|我說：「我的上帝啊， 不要使我中年去世。 你的年數世世無窮！」
PS|102|25|你起初立了地的根基， 天也是你手所造的。
PS|102|26|天地都會消滅，你卻長存； 天地都會像外衣漸漸舊了。 你要將天地如內衣更換， 天地就都改變了。
PS|102|27|惟有你永不改變， 你的年數沒有窮盡。
PS|102|28|你僕人的子孫要安然居住， 他們的後裔要堅立在你面前。
PS|103|1|我的心哪，你要稱頌耶和華！ 凡在我裏面的，都要稱頌他的聖名！
PS|103|2|我的心哪，你要稱頌耶和華！ 不可忘記他一切的恩惠！
PS|103|3|他赦免你一切的罪孽， 醫治你一切的疾病。
PS|103|4|他救贖你的命脫離地府， 以仁愛和憐憫為你的冠冕。
PS|103|5|他用美物使你的生命 得以滿足， 以致你如鷹返老還童。
PS|103|6|耶和華施行公義， 為所有受欺壓的人伸冤。
PS|103|7|他使 摩西 知道他的法則， 使 以色列 人曉得他的作為。
PS|103|8|耶和華有憐憫，有恩惠， 不輕易發怒，且有豐盛的慈愛。
PS|103|9|他不長久責備， 也不永遠懷怒。
PS|103|10|他沒有按我們的罪待我們， 也沒有照我們的罪孽報應我們。
PS|103|11|天離地何等的高， 他的慈愛向敬畏他的人也是何等的大！
PS|103|12|東離西有多遠， 他叫我們的過犯離我們也有多遠！
PS|103|13|父親怎樣憐憫他的兒女， 耶和華也怎樣憐憫敬畏他的人！
PS|103|14|因為他知道我們的本體， 思念我們不過是塵土。
PS|103|15|至於世人，他的年日如草一樣。 他興旺如野地的花，
PS|103|16|經風一吹，就歸無有， 它的原處也不再認識它。
PS|103|17|但耶和華的慈愛歸於敬畏他的人， 從亙古到永遠； 他的公義也歸於子子孫孫，
PS|103|18|就是那些遵守他的約、 記念他的訓詞而遵行的人。
PS|103|19|耶和華在天上立定寶座， 他的國統管萬有。
PS|103|20|聽從他命令、成全他旨意、 有大能的天使啊，你們都要稱頌耶和華！
PS|103|21|你們行他所喜悅的， 作他諸軍，作他僕役的啊，都要稱頌耶和華！
PS|103|22|你們一切被他造的， 在他所治理的各處， 都要稱頌耶和華！ 我的心哪，你要稱頌耶和華！
PS|104|1|我的心哪，你要稱頌耶和華！ 耶和華－我的上帝啊，你為至大！ 你以尊榮威嚴為衣，
PS|104|2|披上亮光，如披外袍， 鋪張穹蒼，如鋪幔子，
PS|104|3|在水中立樓閣的棟梁， 用雲彩為車輦， 藉著風的翅膀而行，
PS|104|4|以風為使者， 以火焰為僕役，
PS|104|5|將地立在根基上， 使地永不動搖。
PS|104|6|你用深水遮蓋地面，猶如衣裳； 諸水高過山嶺。
PS|104|7|你的斥責一發，水就奔逃； 你的雷聲一發，水就奔流。
PS|104|8|諸山上升，諸谷下沉， 歸你為它所立定之地。
PS|104|9|你定了界限，使水不能超越， 不再轉回淹沒大地。
PS|104|10|耶和華使泉源湧在山谷， 流在山間，
PS|104|11|使野地的走獸有水喝， 野驢得解其渴。
PS|104|12|天上的飛鳥在水旁住宿， 在枝幹間啼叫。
PS|104|13|他從樓閣中澆灌山嶺； 因他作為的功效，地就豐足。
PS|104|14|他使草生長，給牲畜吃， 使菜蔬生長，供給人用 ， 使人從地裏得食物，
PS|104|15|得酒能悅人心， 得油能潤人面， 得糧能養人心。
PS|104|16|佳美的樹木， 就是耶和華所栽種的 黎巴嫩 的香柏樹， 都滿了汁漿。
PS|104|17|雀鳥在其上搭窩， 鸛以松樹 為家。
PS|104|18|高山為野山羊的居所， 巖石為石獾的藏身處。
PS|104|19|你安置月亮以定季節， 太陽自知沉落。
PS|104|20|你造黑暗為夜， 林中的百獸就都爬出來。
PS|104|21|少壯獅子吼叫覓食， 向上帝尋求食物。
PS|104|22|太陽一出，獸就躲避， 躺臥在洞裏。
PS|104|23|人出去做工， 勞碌直到晚上。
PS|104|24|耶和華啊，你所造的何其多！ 都是你用智慧造成的， 全地遍滿了你所造之物。
PS|104|25|那裏有海，又大又廣， 其中有無數的動物， 大小活物都有。
PS|104|26|那裏有船行走， 有你所造的 力威亞探 悠游在其中。
PS|104|27|這些都仰望你按時給牠們食物。
PS|104|28|你給牠們，牠們就拾起來； 你張手，牠們就飽得美食。
PS|104|29|你轉臉，牠們就驚惶； 你收回牠們的氣，牠們就死亡，歸於塵土。
PS|104|30|你差遣你的靈，牠們就受造； 你使地面更換為新。
PS|104|31|願耶和華的榮耀存到永遠！ 願耶和華喜愛自己所造的！
PS|104|32|他看地，地便震動； 他摸山，山就冒煙。
PS|104|33|我一生要向耶和華唱詩！ 我還活的時候，要向我的上帝歌頌！
PS|104|34|願他悅納我的默念！ 我要因耶和華歡喜！
PS|104|35|願罪人從世上消滅！ 願惡人歸於無有！ 我的心哪，你要稱頌耶和華！ 哈利路亞 ！
PS|105|1|你們要稱謝耶和華，求告他的名， 在萬民中傳揚他的作為！
PS|105|2|要向他唱詩，向他歌頌， 述說他一切奇妙的作為！
PS|105|3|要誇耀他的聖名！ 願尋求耶和華的人心中歡喜！
PS|105|4|要尋求耶和華與他的能力， 時常尋求他的面。
PS|105|5|他僕人 亞伯拉罕 的後裔， 他所揀選 雅各 的子孫哪， 要記念他奇妙的作為和他的奇事， 並他口中的判語。
PS|105|6|
PS|105|7|他是耶和華－我們的上帝， 全地都有他的判斷。
PS|105|8|他記念他的約，直到永遠； 記念他吩咐的話，直到千代，
PS|105|9|就是與 亞伯拉罕 所立的約， 向 以撒 所起的誓。
PS|105|10|他將這約向 雅各 定為律例， 向 以色列 定為永遠的約，
PS|105|11|說：「我必將 迦南 地賜給你， 作你們應得的產業。」
PS|105|12|當時，他們人丁有限， 數目稀少，在那地寄居。
PS|105|13|他們從這邦遊到那邦， 從這國去到另一民族。
PS|105|14|他不容人欺負他們， 為他們的緣故責備君王：
PS|105|15|「不可傷害我的受膏者， 也不可惡待我的先知。」
PS|105|16|他命饑荒降在那地， 斷絕日用的糧食 ，
PS|105|17|在他們以先差遣一個人前往， 約瑟 被賣為奴。
PS|105|18|人用腳鐐傷他的腳， 他被鐵的項鏈捆鎖。
PS|105|19|耶和華的話試煉他， 直等所說的應驗了。
PS|105|20|王差人將他解開， 治理萬民的把他釋放，
PS|105|21|立他為王家之主， 掌管他一切所有的，
PS|105|22|使他隨意捆綁他的臣宰， 將智慧教導他的長老。
PS|105|23|以色列 也到了 埃及 ， 雅各 在 含 地寄居。
PS|105|24|耶和華使他的百姓生養眾多， 使他們比敵人強盛，
PS|105|25|他使敵人的心轉去恨他的百姓， 用詭計待他的僕人。
PS|105|26|他差遣他的僕人 摩西 和他所揀選的 亞倫 ，
PS|105|27|在敵人中間顯他的神蹟， 在 含 地顯他的奇事。
PS|105|28|他差遣黑暗，就有黑暗； 他們沒有違背他的話。
PS|105|29|他使 埃及 的水變為血， 令他們的魚死了。
PS|105|30|在他們的地上，青蛙多多滋生， 王宮的內室也是如此。
PS|105|31|他一吩咐，蒼蠅就成群飛來， 並有蚊子進入他們四境。
PS|105|32|他給他們降下冰雹為雨， 在他們的地上降下火焰。
PS|105|33|他擊打他們的葡萄樹和無花果樹， 毀壞他們境內的樹木。
PS|105|34|他一吩咐，就有蝗蟲蝻子上來， 不計其數，
PS|105|35|吃光他們地上各樣的菜蔬， 吞盡他們田地的出產。
PS|105|36|他又擊殺他們國內 所有的長子， 就是他們強壯時頭生的。
PS|105|37|他卻帶領自己的百姓帶著金子銀子出來， 他支派中沒有一個走不動的。
PS|105|38|他們出來的時候， 埃及 人就歡喜； 因為 埃及 人懼怕他們。
PS|105|39|他鋪張雲彩當遮蔽， 夜間使火光照。
PS|105|40|他們祈求，他就使鵪鶉飛來， 並用天上的糧食使他們飽足。
PS|105|41|他敲開磐石，水就湧出； 在乾旱之處，水流成河。
PS|105|42|這都因他記念他的聖言 和他的僕人 亞伯拉罕 。
PS|105|43|他帶領自己的百姓歡樂而出， 帶領自己的選民歡呼前往。
PS|105|44|他把列國的地賜給他們， 他們就承受萬民勞碌得來的，
PS|105|45|好讓他們遵他的律例， 守他的律法。 哈利路亞！
PS|106|1|哈利路亞！ 你們要稱謝耶和華，因他本為善， 他的慈愛永遠長存！
PS|106|2|誰能傳揚耶和華的大能？ 誰能表明他一切的美德？
PS|106|3|凡遵守公平、常行公義的， 這人有福了！
PS|106|4|耶和華啊，你恩待你百姓的時候，求你記念我； 你拯救他們的時候，求你眷顧我，
PS|106|5|好使我經歷你選民的福分， 享受你國民的喜樂， 與你的產業一同誇耀。
PS|106|6|我們與我們的祖宗一同犯罪， 偏邪行惡。
PS|106|7|我們的祖宗在 埃及 不明白你的奇事， 不記念你豐盛的慈愛， 反倒在 紅海 行了悖逆。
PS|106|8|然而，他因自己的名拯救他們， 為要彰顯他的大能。
PS|106|9|他斥責 紅海 ，海就乾了， 帶領他們走過深海，如走曠野。
PS|106|10|他拯救他們脫離恨他們之人的手， 從仇敵手中救贖他們。
PS|106|11|水淹沒他們的敵人， 沒有一個存留。
PS|106|12|那時，他們才信他的話， 歌唱讚美他。
PS|106|13|很快地，他們就忘了他的作為， 不仰望他的指引，
PS|106|14|反倒在曠野起了貪婪之心， 在荒地試探上帝。
PS|106|15|他將他們所求的賜給他們， 卻使他們心靈軟弱。
PS|106|16|他們在營中嫉妒 摩西 和耶和華的聖者 亞倫 。
PS|106|17|地就裂開，吞下 大坍 ， 掩蓋 亞比蘭 一夥的人。
PS|106|18|有火在他們黨中點燃， 有火焰燒燬了惡人。
PS|106|19|他們在 何烈山 造了牛犢， 叩拜鑄成的像，
PS|106|20|將他們榮耀的主 換為吃草之牛的像，
PS|106|21|忘了上帝－他們的救主， 就是曾在 埃及 行大事，
PS|106|22|在 含 地行奇事， 在 紅海 行可畏之事的那位。
PS|106|23|因此，他說要滅絕他們； 若非他所揀選的 摩西 在他面前站在破裂之處， 使他的憤怒轉消， 恐怕他就滅絕他們了。
PS|106|24|他們又藐視那美地， 不信他的話，
PS|106|25|在自己帳棚內發怨言， 不聽耶和華的聲音。
PS|106|26|所以他向他們起誓， 必叫他們倒在曠野，
PS|106|27|叫他們的後裔倒在列國之中， 分散在各地。
PS|106|28|他們又與 巴力‧毗珥 連合， 吃了祭死人的物。
PS|106|29|他們這樣行，惹耶和華發怒， 就有瘟疫流行在他們中間。
PS|106|30|那時， 非尼哈 起而干預， 瘟疫這才止息。
PS|106|31|那就算他為義， 世世代代，直到永遠。
PS|106|32|他們在 米利巴 水又惹耶和華發怒， 甚至 摩西 也因他們的緣故受虧損，
PS|106|33|是因他們觸怒了他的靈， 摩西就用嘴說了急躁的話。
PS|106|34|他們不照耶和華所吩咐的 滅絕外邦人，
PS|106|35|反倒與列國相交， 學習他們的行為，
PS|106|36|事奉他們的偶像， 這就成了自己的圈套。
PS|106|37|他們把自己的兒女祭祀鬼魔，
PS|106|38|流無辜人的血， 就是自己兒女的血， 用他們祭祀 迦南 的偶像， 那地就被血玷污了。
PS|106|39|這樣，他們被自己所做的玷污了， 在行為上犯了淫亂。
PS|106|40|耶和華的怒氣向他的百姓發作， 他憎惡自己的產業，
PS|106|41|將他們交在外邦人手裏， 恨他們的人就轄制他們。
PS|106|42|他們的仇敵欺壓他們， 他們伏在敵人手下。
PS|106|43|他屢次搭救他們， 他們卻圖謀悖逆， 就因自己的罪孽降為卑下。
PS|106|44|然而，他聽見他們哀告的時候， 就眷顧他們的急難，
PS|106|45|為了他們，他記念自己的約， 照他豐盛的慈愛改變心意，
PS|106|46|使他們在凡擄掠他們的人面前蒙憐憫。
PS|106|47|耶和華－我們的上帝啊，求你拯救我們， 從列國中召集我們， 我們好頌揚你的聖名， 以讚美你為誇勝。
PS|106|48|耶和華－ 以色列 的上帝是應當稱頌的， 從亙古直到永遠。 願全體百姓都說：「阿們！」 哈利路亞！
PS|107|1|你們要稱謝耶和華，因他本為善， 他的慈愛永遠長存！
PS|107|2|願耶和華救贖的百姓說這話， 就是他從敵人手中所救贖，
PS|107|3|從各地，從東從西， 從北從海那邊召集來的。
PS|107|4|他們在曠野、在荒地飄流， 找不到可居住的城，
PS|107|5|又飢又渴， 心裏發昏。
PS|107|6|於是他們在急難中哀求耶和華， 他就搭救他們脫離禍患，
PS|107|7|又領他們行走直路， 前往可居住的城。
PS|107|8|但願人因耶和華的慈愛 和他向人所做的奇事都稱謝他；
PS|107|9|因他使心裏渴慕的人得以滿足， 使飢餓的人得飽美食。
PS|107|10|那些坐在黑暗中、死蔭裏的人， 被困苦和鐵鏈捆鎖，
PS|107|11|是因他們違背上帝的言語， 藐視至高者的旨意。
PS|107|12|所以，他用勞苦制伏他們的心； 他們仆倒，無人扶助。
PS|107|13|於是他們在急難中哀求耶和華， 他就拯救他們脫離禍患。
PS|107|14|他從黑暗中、從死蔭裏領他們出來， 扯斷他們的捆綁。
PS|107|15|但願人因耶和華的慈愛 和他向人所做的奇事都稱謝他；
PS|107|16|因為他打破了銅門， 砍斷了鐵閂。
PS|107|17|愚妄人因自己叛逆的行徑 和自己的罪孽受苦楚。
PS|107|18|他們心裏厭惡各樣的食物， 就臨近死亡之門。
PS|107|19|於是他們在急難中哀求耶和華， 他就拯救他們脫離禍患。
PS|107|20|他發出自己的話語醫治他們， 救他們脫離陰府。
PS|107|21|但願人因耶和華的慈愛 和他向人所做的奇事都稱謝他。
PS|107|22|願他們以感謝為祭獻給他， 歡呼述說他的作為！
PS|107|23|那些搭船出海， 在大水中做生意的，
PS|107|24|他們看見耶和華的作為， 並他在深海中的奇事。
PS|107|25|他一出令，狂風捲起， 波浪翻騰。
PS|107|26|他們上到天空，下到海底， 他們的心因患難而消沉。
PS|107|27|他們搖搖晃晃，東倒西歪，好像醉酒的人， 他們的智慧無法可施。
PS|107|28|於是他們在急難中哀求耶和華， 他就領他們脫離禍患。
PS|107|29|他使狂風止息， 波浪平靜，
PS|107|30|既平靜了，他們就歡喜， 他就領他們到想要去的海港。
PS|107|31|但願人因耶和華的慈愛 和他向人所做的奇事都稱謝他。
PS|107|32|願他們在百姓的會中尊崇他， 在長老的座位上讚美他！
PS|107|33|他使江河變為曠野， 叫水泉變為乾涸之地，
PS|107|34|使肥沃之地變為荒蕪的鹽地， 都因當地居民的邪惡。
PS|107|35|他使曠野變為水潭， 叫旱地變為水泉，
PS|107|36|使飢餓的人住在那裏， 建造可居住的城，
PS|107|37|又種田地，栽葡萄園， 得享所出產的果實。
PS|107|38|他賜福給他們，使他們生養眾多， 也不叫他們的牲畜減少。
PS|107|39|但他們因欺壓、患難、愁苦， 人口減少而且卑微。
PS|107|40|他使貴族蒙羞受辱， 使他們迷失在荒涼無路之地；
PS|107|41|卻將窮乏人安置在高處，脫離苦難， 使他的家屬多如羊群。
PS|107|42|正直的人看見就歡喜， 罪孽之輩卻要啞口無言。
PS|107|43|凡有智慧的必在這些事上留心， 他必思想耶和華的慈愛。
PS|108|1|上帝啊，我心堅定； 我口 要唱詩歌頌！
PS|108|2|琴瑟啊，當醒起！ 我要喚起曙光！
PS|108|3|耶和華啊，我要在萬民中稱謝你， 在萬族中歌頌你！
PS|108|4|因為你的慈愛大過諸天， 你的信實達到穹蒼。
PS|108|5|上帝啊，願你崇高過於諸天！ 願你的榮耀高過全地！
PS|108|6|求你應允我，用右手施行拯救， 好讓你所親愛的人得救。
PS|108|7|上帝在他的聖所 說： 「我要歡樂； 要劃分 示劍 ， 丈量 疏割谷 。
PS|108|8|基列 是我的， 瑪拿西 是我的， 以法蓮 是護衛我頭的， 猶大 是我的權杖。
PS|108|9|摩押 是我的沐浴盆， 我要向 以東 扔鞋， 我必因勝 非利士 而歡呼。」
PS|108|10|誰能領我進堅固城？ 誰能引我到 以東 地？
PS|108|11|上帝啊，你真的丟棄了我們嗎？ 上帝啊，你不和我們的軍隊同去嗎？
PS|108|12|求你幫助我們攻擊敵人， 因為人的幫助是枉然的。
PS|108|13|我們倚靠上帝才得施展大能， 因為踐踏我們敵人的就是他。
PS|109|1|我所讚美的上帝啊， 求你不要閉口不言。
PS|109|2|因為惡人的嘴和詭詐人的口張開攻擊我， 他們用撒謊的舌頭對我說話。
PS|109|3|他們圍繞我，說怨恨的話， 又無故地攻打我。
PS|109|4|他們與我作對回報我的愛， 但我專心祈禱。
PS|109|5|他們向我以惡報善， 以恨報愛。
PS|109|6|求你派惡人轄制他， 派對頭站在他右邊！
PS|109|7|他受審判的時候， 願他背負罪名而出！ 願他的祈禱反成為罪！
PS|109|8|願他的年歲短少！ 願別人得他的職分！
PS|109|9|願他的兒女成為孤兒， 他的妻子成為寡婦！
PS|109|10|願他的兒女飄流討飯， 從荒涼之處出來求乞 ！
PS|109|11|願債主牢籠他一切所有的！ 願陌生人搶走他勞碌得來的！
PS|109|12|願無人向他佈施恩惠， 無人恩待他的孤兒！
PS|109|13|願他的後人斷絕， 名字被塗去，不傳於下代！
PS|109|14|願耶和華記得他祖宗的罪孽， 不塗去他母親的罪過！
PS|109|15|願這些罪常在耶和華面前！ 願他們的名字 從地上除滅！
PS|109|16|因為他從未想過要施恩， 卻迫害困苦貧窮的和傷心的人， 把他們處死。
PS|109|17|他愛咒罵，咒罵就臨到他； 他不喜愛祝福，祝福就遠離他！
PS|109|18|他拿咒罵當衣服穿上； 這咒罵就如水進到他裏面， 如油進入他骨頭。
PS|109|19|願這咒罵當他遮身的衣服， 作他經常束腰的帶子！
PS|109|20|這就是那些與我作對、用惡言議論我的人 從耶和華所受的報應。
PS|109|21|但是你，主－耶和華啊， 求你因你的名採取行動； 因你的慈愛美好，求你搭救我！
PS|109|22|因為我困苦貧窮， 內心受傷。
PS|109|23|我如日影偏斜而去， 如蝗蟲被抖出來。
PS|109|24|我因禁食，膝蓋軟弱； 我身體消瘦，不再豐潤。
PS|109|25|我受他們的羞辱， 他們看見我就搖頭。
PS|109|26|耶和華－我的上帝啊，求你幫助我， 照你的慈愛拯救我，
PS|109|27|好讓他們知道這是你的手， 是你－耶和華所做的事。
PS|109|28|任憑他們咒罵，你卻要賜福； 他們幾時起來就必蒙羞， 你的僕人卻要歡喜。
PS|109|29|願與我作對的人披戴羞辱！ 願他們以自己的羞愧作外袍遮身！
PS|109|30|我要用口極力稱謝耶和華， 我要在眾人中間讚美他；
PS|109|31|因為他必站在貧窮人的右邊， 救他脫離定他死罪的人。
PS|110|1|耶和華對我主說： 「你坐在我的右邊， 等我使你仇敵作你的腳凳。」
PS|110|2|耶和華必使你從 錫安 伸出你能力的權杖； 你務要在仇敵中掌權。
PS|110|3|你在聖山上 掌權的日子， 你的子民必甘心跟隨 ； 從晨曦初現， 你就有清晨 的甘露。
PS|110|4|耶和華起了誓，絕不改變： 「你是照著 麥基洗德 的體系永遠為祭司。」
PS|110|5|在你右邊的主， 當他發怒的日子，必打傷列王。
PS|110|6|他要審判列國， 屍首就佈滿各處； 他要痛擊遍地的領袖。
PS|110|7|他要喝路旁的河水， 因此必抬起頭來。
PS|111|1|哈利路亞！ 我要在正直人的大會和會眾中 一心稱謝耶和華。
PS|111|2|耶和華的作為本為大， 被所有喜愛的人所探尋。
PS|111|3|他所做的是尊榮和威嚴， 他的公義存到永遠。
PS|111|4|他行了奇事，使人記念； 耶和華有恩惠，有憐憫。
PS|111|5|他賜糧食給敬畏他的人， 他必永遠記念他的約。
PS|111|6|他向百姓顯出大能的作為， 將列國賜給他們為業。
PS|111|7|他手所做的信實公平， 他的訓詞全然可靠，
PS|111|8|是永永遠遠堅定的， 是按信實正直設立的。
PS|111|9|他向百姓施行救贖， 頒佈他的約，直到永遠； 他的名聖而可畏。
PS|111|10|敬畏耶和華是智慧的開端， 凡遵行他命令的有美好的見識。 耶和華是永遠當讚美的！
PS|112|1|哈利路亞！ 敬畏耶和華，甚喜愛他命令的， 這人有福了！
PS|112|2|他的後裔在世必強盛， 正直人的後代必蒙福。
PS|112|3|他的家中有金銀財寶， 他的義行存到永遠。
PS|112|4|正直人在黑暗中有光向他照耀， 他有恩惠，有憐憫，有公義。
PS|112|5|施恩與人、借貸與人、秉公處事的人 必享美福，
PS|112|6|他永不動搖。 義人被記念，直到永遠。
PS|112|7|他不懼怕兇惡的信息， 他的心堅定，倚靠耶和華。
PS|112|8|他的心確定，總不懼怕， 直到他看見敵人遭報。
PS|112|9|他施捨，賙濟貧窮， 他的義行存到永遠， 他的角必被高舉，大有榮耀。
PS|112|10|惡人看見就憤怒，必咬牙而消亡， 惡人的心願要歸於幻滅。
PS|113|1|哈利路亞！ 耶和華的僕人哪，你們要讚美， 讚美耶和華的名！
PS|113|2|耶和華的名是應當稱頌的， 從今時直到永遠！
PS|113|3|從日出之地到日落之處， 耶和華的名是應當讚美的！
PS|113|4|耶和華超乎萬國之上， 他的榮耀高過諸天。
PS|113|5|誰像耶和華－我們的上帝呢？ 他坐在至高之處，
PS|113|6|自己謙卑， 觀看天上地下的事。
PS|113|7|他從灰塵裏抬舉貧寒的人， 從糞堆中提拔貧窮的人，
PS|113|8|使他們與貴族同坐， 與本國的貴族同坐。
PS|113|9|他使不孕的婦女安居家中， 成為快樂的母親，兒女成群。 哈利路亞！
PS|114|1|以色列 出 埃及 ， 雅各 家離開說陌生語言之民時，
PS|114|2|猶大 作主的聖所， 以色列 為他所治理的國。
PS|114|3|滄海看見就奔逃， 約旦河 也倒流。
PS|114|4|大山踴躍如公羊， 小山跳舞如羔羊。
PS|114|5|滄海啊，你為何奔逃？ 約旦 哪，你為何倒流？
PS|114|6|大山哪，你為何踴躍如公羊？ 小山哪，你為何跳舞如羔羊？
PS|114|7|大地啊，在主的面前， 在 雅各 的上帝的面前，震動吧！
PS|114|8|他叫磐石變為水池， 使堅石變為泉源。
PS|115|1|耶和華啊，榮耀不要歸與我們， 不要歸與我們； 要因你的慈愛和信實歸在你的名下！
PS|115|2|為何讓列國說 「他們的上帝在哪裏」呢？
PS|115|3|但是，我們的上帝在天上， 萬事都隨自己的旨意而行。
PS|115|4|他們的偶像是金的，是銀的， 是人手所造的，
PS|115|5|有口卻不能言， 有眼卻不能看，
PS|115|6|有耳卻不能聽， 有鼻卻不能聞，
PS|115|7|有手卻不能摸， 有腳卻不能走， 有喉卻不能說話。
PS|115|8|造它們的要像它們一樣， 凡靠它們的也必如此。
PS|115|9|以色列 啊，要倚靠耶和華！ 他是人的幫助和盾牌。
PS|115|10|亞倫 家啊，要倚靠耶和華！ 他是人的幫助和盾牌。
PS|115|11|敬畏耶和華的人哪，要倚靠耶和華！ 他是人的幫助和盾牌。
PS|115|12|耶和華向來眷念我們， 他還要賜福， 賜福給 以色列 家， 賜福給 亞倫 家。
PS|115|13|凡敬畏耶和華的，無論大小， 主必賜福給他。
PS|115|14|願耶和華使你們 和你們的子孫日見增加。
PS|115|15|你們蒙了耶和華的福， 他是創造天地的主宰。
PS|115|16|天，是耶和華的天； 地，他卻給了世人。
PS|115|17|死人不能讚美耶和華， 下到寂靜 中的也都不能。
PS|115|18|但我們要稱頌耶和華， 從今時直到永遠。 哈利路亞！
PS|116|1|我愛耶和華， 因為他聽了我的聲音和我的懇求。
PS|116|2|他既向我側耳， 我一生要求告他。
PS|116|3|死亡的繩索勒住我， 陰間的痛苦抓住我， 我遭遇患難愁苦。
PS|116|4|那時，我求告耶和華的名： 「耶和華啊，求你救我！」
PS|116|5|耶和華有恩惠，有公義， 我們的上帝有憐憫。
PS|116|6|耶和華保護愚蒙的人； 我落到卑微的地步，他救了我。
PS|116|7|我的心哪！你要復歸安寧， 因為耶和華用厚恩待你。
PS|116|8|主啊，你救我的命脫離死亡， 使我的眼不再流淚， 使我的腳不致跌倒。
PS|116|9|我行在耶和華面前， 走在活人之地。
PS|116|10|我信，儘管我說： 「我受了極大的困苦。」
PS|116|11|我曾驚惶地說： 「人都是說謊的！」
PS|116|12|耶和華向我賞賜一切厚恩， 我拿甚麼來報答他呢？
PS|116|13|我要舉起救恩的杯， 稱揚耶和華的名。
PS|116|14|我要在他的全體百姓面前 向耶和華還我所許的願。
PS|116|15|在耶和華眼中， 聖民之死極為寶貴。
PS|116|16|耶和華啊，哦，我是你的僕人； 我是你的僕人，是你使女的兒子。 你已經解開我的捆索。
PS|116|17|我要以感謝為祭獻給你， 又要求告耶和華的名。
PS|116|18|我要在 耶路撒冷 當中， 在耶和華殿的院內， 在他的全體百姓面前， 向耶和華還我所許的願。 哈利路亞！
PS|116|19|
PS|117|1|萬國啊，你們要讚美耶和華！ 萬族啊，你們都要頌讚他！
PS|117|2|因為他向我們大施慈愛， 耶和華的信實存到永遠。 哈利路亞！
PS|118|1|你們要稱謝耶和華，因他本為善； 他的慈愛永遠長存！
PS|118|2|願 以色列 說： 「他的慈愛永遠長存！」
PS|118|3|願 亞倫 家說： 「他的慈愛永遠長存！」
PS|118|4|願敬畏耶和華的人說： 「他的慈愛永遠長存！」
PS|118|5|我在急難中求告耶和華， 耶和華就應允我，把我安置在寬闊之地。
PS|118|6|耶和華在我這邊 ，我必不懼怕， 人能把我怎麼樣呢？
PS|118|7|在那幫助我的人中，有耶和華幫助我， 所以我要看見那些恨我的人遭報。
PS|118|8|投靠耶和華， 強似倚賴人；
PS|118|9|投靠耶和華， 強似倚賴權貴。
PS|118|10|列邦圍繞我， 我靠耶和華的名必剿滅他們。
PS|118|11|他們圍繞我，圍困我， 我靠耶和華的名必剿滅他們。
PS|118|12|他們如同蜜蜂一般地圍繞我， 他們熄滅，好像燒荊棘的火； 我靠耶和華的名，必剿滅他們。
PS|118|13|你用力推我，要叫我跌倒， 但耶和華幫助了我。
PS|118|14|耶和華是我的力量，是我的詩歌， 他也成了我的拯救。
PS|118|15|在義人的帳棚裏，有歡呼拯救的聲音， 耶和華的右手施展大能。
PS|118|16|耶和華的右手高舉， 耶和華的右手施展大能。
PS|118|17|我不至於死，仍要存活， 並要傳揚耶和華的作為。
PS|118|18|耶和華雖嚴嚴地懲治我， 卻未曾將我交於死亡。
PS|118|19|給我敞開義門， 我要進去稱謝耶和華！
PS|118|20|這是耶和華的門， 義人要進去！
PS|118|21|我要稱謝你，因為你已經應允我， 又成了我的拯救！
PS|118|22|匠人所丟棄的石頭 已成了房角的頭塊石頭。
PS|118|23|這是耶和華所做的， 在我們眼中看為奇妙。
PS|118|24|這是耶和華所定的日子， 我們在其中要高興歡喜！
PS|118|25|耶和華啊，求你拯救 ！ 耶和華啊，求你使我們順利！
PS|118|26|奉耶和華的名來的是應當稱頌的！ 我們從耶和華的殿中為你們祝福！
PS|118|27|耶和華是上帝， 他光照了我們。 你們要用繩索把祭牲拴住， 直牽到壇角。
PS|118|28|你是我的上帝，我要稱謝你！ 我的上帝啊，我要尊崇你 ！
PS|118|29|你們要稱謝耶和華，因他本為善； 他的慈愛永遠長存！
PS|119|1|行為正直、遵行耶和華律法的， 這人有福了！
PS|119|2|遵守他的法度、一心尋求他的， 這人有福了！
PS|119|3|他們不做不義的事， 但遵行他的道。
PS|119|4|耶和華啊，你曾將你的訓詞吩咐我們， 為要我們切實遵守。
PS|119|5|但願我行事堅定， 得以遵守你的律例。
PS|119|6|我看重你的一切命令， 就不致羞愧。
PS|119|7|我學習你公義的典章， 要以正直的心稱謝你。
PS|119|8|我必遵守你的律例， 求你不要把我全然棄絕！
PS|119|9|青年要如何保持純潔呢？ 是要遵行你的話！
PS|119|10|我曾一心尋求你， 求你不要使我偏離你的命令。
PS|119|11|我將你的話藏在心裏， 免得我得罪你。
PS|119|12|耶和華啊，你是應當稱頌的！ 求你將你的律例教導我！
PS|119|13|我用嘴唇傳揚 你口中一切的典章。
PS|119|14|我喜愛你的法度， 如同喜愛一切的財物。
PS|119|15|我要默想你的訓詞， 看重你的道路。
PS|119|16|我要以你的律例為樂， 我不忘記你的話。
PS|119|17|求你用厚恩待你的僕人，使我存活， 我就遵守你的話。
PS|119|18|求你開我的眼睛， 使我看出你律法中的奇妙。
PS|119|19|我在地上是寄居的人， 求你不要向我隱藏你的命令！
PS|119|20|我時常切慕你的典章， 耗盡心力。
PS|119|21|受詛咒、偏離你命令的驕傲人， 你已經責備他們。
PS|119|22|求你除掉我所受的羞辱和藐視， 因我遵守你的法度。
PS|119|23|雖有掌權者坐著妄論我， 你僕人卻思想你的律例。
PS|119|24|你的法度也是我的喜樂， 我的導師 。
PS|119|25|我的性命幾乎歸於塵土， 求你照你的話將我救活！
PS|119|26|我述說我所做的，你應允了我； 求你將你的律例教導我！
PS|119|27|求你使我明白你的訓詞， 我要默想你的奇事。
PS|119|28|我因愁苦身心耗盡， 求你照你的話使我堅立！
PS|119|29|求你使我離開奸詐的道路， 開恩將你的律法賜給我！
PS|119|30|我選擇了忠信的道路， 將你的典章擺在我面前。
PS|119|31|我持守你的法度； 耶和華啊，求你不要叫我羞愧！
PS|119|32|你使我心胸開闊的時候， 我就往你命令的道路直奔。
PS|119|33|耶和華啊，求你將你的律例指教我， 我必遵守到底！
PS|119|34|求你賜我悟性，我就遵守你的律法， 且要一心遵守。
PS|119|35|求你叫我遵行你的命令， 因為這是我所喜愛的。
PS|119|36|求你使我的心趨向你的法度， 不趨向不義之財。
PS|119|37|求你叫我轉眼不看虛假， 使我活在你的道路 中。
PS|119|38|求你向敬畏你的僕人 堅守你的話！
PS|119|39|求你使我所懼怕的羞辱遠離我， 因你的典章本為美。
PS|119|40|看哪，我切慕你的訓詞， 求你因你的公義賜我生命 ！
PS|119|41|耶和華啊，求你使你的慈愛臨到我， 照你的話使你的救恩臨到我，
PS|119|42|我就有話回答那羞辱我的， 因我倚靠你的話。
PS|119|43|求你叫真理的話總不離開我的口， 因我仰望你的典章。
PS|119|44|我要常守你的律法， 直到永永遠遠。
PS|119|45|我要自由而行 ， 因我尋求了你的訓詞。
PS|119|46|我要在列王面前宣講你的法度， 也不致羞愧。
PS|119|47|我以你的命令為樂， 這命令是我所喜愛的。
PS|119|48|我向我所愛的，就是你的命令高舉雙手 ， 我也要默想你的律例。
PS|119|49|求你記念你向僕人所說的話， 這話使我有盼望。
PS|119|50|你的話將我救活了； 這是我在患難中的安慰。
PS|119|51|驕傲的人極度地侮慢我， 我卻未曾偏離你的律法。
PS|119|52|耶和華啊，我記念你從古以來的典章， 就得了安慰。
PS|119|53|我因惡人離棄你的律法， 怒火中燒。
PS|119|54|我在世寄居， 以你的律例為詩歌。
PS|119|55|耶和華啊，我夜間記念你的名， 我也要遵守你的律法。
PS|119|56|這臨到我， 是因我謹守你的訓詞。
PS|119|57|耶和華是我的福分； 我曾說，我要遵守你的話。
PS|119|58|我一心懇求你的面， 求你照你的話憐憫我！
PS|119|59|我思想自己所行的道路， 我的腳步就轉向你的法度。
PS|119|60|我速速遵守你的命令， 並不遲延。
PS|119|61|惡人的繩索纏繞我， 我卻沒有忘記你的律法。
PS|119|62|我因你公義的典章， 夜半起來稱謝你。
PS|119|63|凡敬畏你、守你訓詞的人， 我都與他作伴。
PS|119|64|耶和華啊，遍地滿了你的慈愛； 求你將你的律例教導我！
PS|119|65|耶和華啊，你照你的話， 善待你的僕人。
PS|119|66|求你教我明辨和知識， 因我信靠你的命令。
PS|119|67|我未受苦以先曾經迷失， 現在卻遵守你的話。
PS|119|68|你本為善，所行的也善； 求你將你的律例教導我！
PS|119|69|驕傲的人編造謊言攻擊我， 我卻要一心遵守你的訓詞。
PS|119|70|他們的心蒙昧如蒙油脂， 我卻喜愛你的律法。
PS|119|71|我受苦是與我有益， 為要使我學習你的律例。
PS|119|72|你口中的律法與我有益， 勝於千萬金銀。
PS|119|73|你的手造了我，塑造我； 求你賜我悟性學習你的命令！
PS|119|74|敬畏你的人看見我就歡喜， 因我仰望你的話。
PS|119|75|耶和華啊，我知道你的典章是公義的； 你使我受苦是以信實待我。
PS|119|76|求你照著你向僕人所說的話， 以慈愛安慰我。
PS|119|77|求你的憐憫臨到我，使我存活， 因你的律法是我的喜樂。
PS|119|78|願驕傲的人蒙羞，因為他們無理傾覆我； 但我要默想你的訓詞。
PS|119|79|願敬畏你的人和知道你法度的人 都歸向我。
PS|119|80|願我的心在你的律例上完全， 使我不致蒙羞。
PS|119|81|我渴想你的救恩身心耗盡， 我仰望你的話。
PS|119|82|我因渴望你的話眼睛失明，說： 「你何時安慰我呢？」
PS|119|83|我雖像煙薰的皮囊， 卻不忘記你的律例。
PS|119|84|你僕人的年日有多少呢？ 你幾時向迫害我的人施行審判呢？
PS|119|85|不順從你律法的驕傲人 為我掘了坑。
PS|119|86|你的命令盡都信實； 他們無理迫害我，求你幫助我！
PS|119|87|他們幾乎把我從世上除滅； 但我沒有離棄你的訓詞。
PS|119|88|求你照你的慈愛將我救活， 我就遵守你口中的法度。
PS|119|89|耶和華啊，你的話安定在天， 直到永遠。
PS|119|90|你的信實存到萬代； 你堅立了地，地就長存。
PS|119|91|天地照你的典章存到今日； 萬物都是你的僕役。
PS|119|92|我若不以你的律法為樂， 早就在苦難中滅絕了！
PS|119|93|我永不忘記你的訓詞， 因你用這訓詞將我救活。
PS|119|94|我是屬你的，求你救我， 因我尋求了你的訓詞。
PS|119|95|惡人等著要滅絕我， 我卻要揣摩你的法度。
PS|119|96|我看萬事盡都有限， 惟有你的命令極其寬廣。
PS|119|97|我何等愛慕你的律法， 終日不住地思想。
PS|119|98|你的命令常存在我心裏， 使我比仇敵有智慧。
PS|119|99|我比我的教師更通達， 因我思想你的法度。
PS|119|100|我比年老的更明白， 因我謹守你的訓詞。
PS|119|101|我阻止我的腳走一切邪路， 為要遵守你的話。
PS|119|102|我沒有偏離你的典章， 因為你教導了我。
PS|119|103|你的言語在我上膛何等甘美， 在我口中比蜜更甜！
PS|119|104|我藉著你的訓詞得以明白， 因此，我恨惡一切虛假的行徑。
PS|119|105|你的話是我腳前的燈， 是我路上的光。
PS|119|106|你公義的典章，我曾起誓遵守， 我必按著誓言而行。
PS|119|107|我極其痛苦； 耶和華啊，求你照你的話將我救活！
PS|119|108|耶和華啊，求你悅納我口中的讚美為甘心祭， 又將你的典章教導我！
PS|119|109|我的性命常在我手掌中 ， 我卻不忘記你的律法。
PS|119|110|惡人為我設下羅網， 我卻沒有偏離你的訓詞。
PS|119|111|我以你的法度為永遠的產業， 因這是我心中所喜愛的。
PS|119|112|我的心傾向你的律例， 謹守到底，直到永遠。
PS|119|113|心懷二意的人為我所恨； 但你的律法為我所愛。
PS|119|114|你是我藏身之處，是我的盾牌； 我仰望你的話。
PS|119|115|作惡的人哪，你們離開我吧！ 我要遵守我上帝的命令。
PS|119|116|求你照你的話扶持我，使我存活， 不要叫我因失望而蒙羞。
PS|119|117|求你扶持我，使我得救， 時常看重你的律例。
PS|119|118|凡偏離你律例的人，你都輕看他們， 因為他們的詭詐必歸虛空。
PS|119|119|你除掉地上所有的惡人，好像除掉渣滓 ； 因此我喜愛你的法度。
PS|119|120|我因懼怕你，肉體戰慄； 我害怕你的典章。
PS|119|121|我行公平和公義， 求你不要撇下我，交給欺壓我的人！
PS|119|122|求你保證你的僕人得福， 不容驕傲的人欺壓我！
PS|119|123|我因盼望你的救恩 和你公義的言語眼睛失明。
PS|119|124|求你照你的慈愛待僕人， 將你的律例教導我。
PS|119|125|我是你的僕人，求你賜我悟性， 得以認識你的法度。
PS|119|126|這是耶和華採取行動的時候， 因人廢棄了你的律法。
PS|119|127|所以，我喜愛你的命令勝於金子， 更勝於純金。
PS|119|128|你的一切訓詞，在萬事上我都以為正直； 我恨惡一切虛假的行徑。
PS|119|129|你的法度奇妙， 所以我一心謹守。
PS|119|130|你的話一開啟就發出亮光， 使愚蒙人通達。
PS|119|131|我大大張口，呼吸急促， 因我切慕你的命令。
PS|119|132|求你轉向我，憐憫我， 就像你待那些喜愛你名的人。
PS|119|133|求你用你的言語使我腳步穩健， 不容罪孽轄制我。
PS|119|134|求你救我脫離人的欺壓， 我要遵守你的訓詞。
PS|119|135|求你使你的臉向僕人發光， 又將你的律例教導我。
PS|119|136|我的眼睛流淚成河， 因為他們不守你的律法。
PS|119|137|耶和華啊，你是公義的； 你的典章正直！
PS|119|138|你所頒佈的法度是公義的， 極其可靠。
PS|119|139|我的狂熱把我燒滅， 因我敵人忘記你的話。
PS|119|140|你的言語極其精煉， 令你僕人喜愛。
PS|119|141|我渺小，被人藐視， 卻不忘記你的訓詞。
PS|119|142|你的公義永遠公義， 你的律法是確實的。
PS|119|143|我遭遇患難愁苦， 你的命令是我的喜樂。
PS|119|144|你的法度永遠公義； 求你賜我悟性，使我存活。
PS|119|145|耶和華啊，我一心呼求你，求你應允我！ 我必謹守你的律例。
PS|119|146|我向你呼求，求你救我！ 我要遵守你的法度。
PS|119|147|天尚未亮我呼喊求救， 我仰望你的話。
PS|119|148|我終夜雙眼睜開， 為要思想你的言語。
PS|119|149|求你按你的慈愛聽我的聲音， 耶和華啊，求你照你的典章將我救活！
PS|119|150|追逐奸惡的人 迫近了， 他們遠離你的律法。
PS|119|151|耶和華啊，你就在我身邊， 你一切的命令是確實的！
PS|119|152|我從你的法度早已知道， 這法度是你永遠立定的。
PS|119|153|求你看顧我的苦難，搭救我， 因我不忘記你的律法。
PS|119|154|求你為我的冤屈辯護，救贖我， 照你的言語將我救活。
PS|119|155|救恩遠離惡人， 因為他們不尋求你的律例。
PS|119|156|耶和華啊，你的憐憫本為大； 求你照你的典章將我救活。
PS|119|157|迫害我的、抵擋我的甚多， 我卻沒有偏離你的法度。
PS|119|158|我看見奸惡的人就憎惡， 因為他們不遵守你的言語。
PS|119|159|你看我何等喜愛你的訓詞！ 耶和華啊，求你按你的慈愛將我救活！
PS|119|160|你話語的精髓是真實的， 你一切公義的典章永遠長存。
PS|119|161|掌權者無故迫害我， 然而我的心畏懼你的話。
PS|119|162|我喜愛你的言語， 好像人得到許多戰利品。
PS|119|163|我恨惡，憎惡虛假； 惟喜愛你的律法。
PS|119|164|我因你公義的典章 一天七次讚美你。
PS|119|165|喜愛你律法的人大有平安， 任何事都不能使他們跌倒。
PS|119|166|耶和華啊，我仰望你的救恩， 遵行你的命令。
PS|119|167|我心謹守你的法度， 這法度我極其喜愛。
PS|119|168|我遵守你的訓詞和法度， 因我所行的道路都在你的面前。
PS|119|169|耶和華啊，願我的呼求達到你面前， 求你照你的話賜我悟性。
PS|119|170|願我的懇求達到你面前， 求你照你的言語搭救我。
PS|119|171|願我的嘴唇發出讚美， 因為你將律例教導我。
PS|119|172|願我的舌頭歌唱你的言語， 因你一切的命令盡都公義。
PS|119|173|求你用你的手幫助我， 因我選擇你的訓詞。
PS|119|174|耶和華啊，我切慕你的救恩！ 你的律法是我的喜樂。
PS|119|175|願我的性命存活，得以讚美你！ 願你的典章幫助我！
PS|119|176|我走迷了路如同失喪的羊，求你尋找你的僕人， 因我不忘記你的命令。
PS|120|1|我在急難中求告耶和華， 他就應允我。
PS|120|2|耶和華啊，求你救我脫離 說謊的嘴唇和詭詐的舌頭！
PS|120|3|詭詐的舌頭啊，他會給你甚麼呢？ 會加給你甚麼呢？
PS|120|4|就是勇士的利箭、 羅騰木 的炭火。
PS|120|5|禍哉！我寄居在 米設 ， 住在 基達 帳棚之中。
PS|120|6|我與那恨惡和平的人 許久同住。
PS|120|7|我願和平， 當我發言，他們卻要戰爭。
PS|121|1|我要向山舉目， 我的幫助從何而來？
PS|121|2|我的幫助 從造天地的耶和華而來。
PS|121|3|他不叫你的腳搖動， 保護你的必不打盹！
PS|121|4|保護 以色列 的 必不打盹，也不睡覺。
PS|121|5|保護你的是耶和華， 耶和華在你右邊蔭庇你。
PS|121|6|白日，太陽必不傷你； 夜間，月亮也不害你。
PS|121|7|耶和華要保護你，免受一切的災害， 他要保護你的性命。
PS|121|8|你出你入，耶和華要保護你， 從今時直到永遠。
PS|122|1|我喜樂， 因人對我說：「我們到耶和華的殿去。」
PS|122|2|耶路撒冷 啊， 我們的腳站在你門內。
PS|122|3|耶路撒冷 被建造， 如同連結整齊的一座城。
PS|122|4|眾支派就是耶和華的支派，上那裏去， 按 以色列 的法度頌揚耶和華的名。
PS|122|5|他們在那裏設立審判的寶座， 就是 大衛 家的寶座。
PS|122|6|你們要為 耶路撒冷 求平安： 「願愛你的人興旺！
PS|122|7|願你城中有平安！ 願你宮內得平靜！」
PS|122|8|為我弟兄和同伴的緣故，我要說： 「願你平安！」
PS|122|9|為耶和華－我們上帝殿的緣故， 我要為你求福！
PS|123|1|坐在天上的主啊， 我向你舉目。
PS|123|2|看哪，僕人的眼睛怎樣仰望主人的手， 婢女的眼睛怎樣仰望女主人的手， 我們的眼睛也照樣仰望耶和華－我們的上帝， 直到他憐憫我們。
PS|123|3|耶和華啊，求你憐憫我們，憐憫我們！ 因為我們受盡了藐視。
PS|123|4|我們受盡了安逸人的譏誚 和驕傲人的藐視。
PS|124|1|說吧， 以色列 ： 「若不是耶和華幫助我們，
PS|124|2|若不是耶和華幫助我們， 當人起來攻擊我們，
PS|124|3|那時，人向我們發怒， 就把我們活活吞了；
PS|124|4|那時，波濤必漫過我們， 河水必淹沒我們；
PS|124|5|那時，狂傲的水 必淹沒我們。」
PS|124|6|耶和華是應當稱頌的！ 他沒有把我們交給他們，作牙齒的獵物。
PS|124|7|我們好像雀鳥，從捕鳥人的羅網裏逃脫， 羅網破裂，我們就逃脫了。
PS|124|8|我們得幫助， 是因造天地之耶和華的名。
PS|125|1|倚靠耶和華的人好像 錫安山 ， 安穩坐鎮，永不動搖。
PS|125|2|眾山怎樣圍繞 耶路撒冷 ， 耶和華也照樣圍繞他的百姓，從今時直到永遠。
PS|125|3|惡人的杖必不在義人的土地上停留， 免得義人伸手作惡。
PS|125|4|耶和華啊，求你善待 行善和心裏正直的人。
PS|125|5|至於那偏行彎曲道路的人， 耶和華必將他們和作惡的人一同驅逐出去。 願平安歸於 以色列 ！
PS|126|1|當耶和華使 錫安 被擄的人歸回的時候， 我們好像做夢的人。
PS|126|2|那時，我們滿口喜笑、 滿舌歡呼； 那時，列國中就有人說： 「耶和華為他們行了大事！」
PS|126|3|耶和華果然為我們行了大事， 我們就歡喜。
PS|126|4|耶和華啊，求你使我們這些被擄的人歸回， 好像 尼革夫 的河水復流。
PS|126|5|流淚撒種的， 必歡呼收割！
PS|126|6|那帶種流淚出去的， 必歡呼地帶禾捆回來！
PS|127|1|若不是耶和華建造房屋， 建造的人就枉然勞力； 若不是耶和華看守城池， 看守的人就枉然警醒。
PS|127|2|你們清晨早起，夜晚安歇， 吃勞碌得來的飯，本是枉然； 惟有耶和華所親愛的， 必叫他安然睡覺。
PS|127|3|看哪，兒女是耶和華所賜的產業， 所懷的胎是他所給的賞賜。
PS|127|4|人在年輕時生的兒女 好像勇士手中的箭。
PS|127|5|箭袋充滿的人有福了！ 他們在城門口和仇敵爭論時必不蒙羞。
PS|128|1|凡敬畏耶和華、 遵行他道的人有福了！
PS|128|2|你要吃勞碌得來的； 你要享福，凡事順利。
PS|128|3|你妻子在你內室，好像多結果子的葡萄樹； 你兒女圍繞你的桌子，如同橄欖樹苗。
PS|128|4|看哪，敬畏耶和華的人 必要這樣蒙福！
PS|128|5|願耶和華從 錫安 賜福給你！ 願你一生一世看見 耶路撒冷 興旺！
PS|128|6|願你看見 你的子子孫孫！ 願平安歸於 以色列 ！
PS|129|1|說吧， 以色列 ： 「從我幼年以來，人屢次苦害我；
PS|129|2|從我幼年以來，人屢次苦害我， 卻沒有勝過我。
PS|129|3|扶犁的人在我背上扶犁而耕， 耕的犁溝很長。」
PS|129|4|耶和華是公義的， 他砍斷了惡人的繩索。
PS|129|5|願恨惡 錫安 的 都蒙羞退後！
PS|129|6|願他們像房頂上的草， 一發芽就枯乾，
PS|129|7|收割的不夠用手抓一把， 捆禾的也不夠抱滿懷。
PS|129|8|過路的也不說：「願耶和華所賜的福歸與你們！ 我們奉耶和華的名給你們祝福！」
PS|130|1|耶和華啊， 我從深處求告你！
PS|130|2|主啊，求你聽我的聲音！ 求你側耳聽我懇求的聲音！
PS|130|3|耶和華啊，你若究察罪孽， 主啊，誰能站得住呢？
PS|130|4|但在你有赦免之恩， 要叫人敬畏你。
PS|130|5|我等候耶和華，我的心等候； 我也仰望他的話。
PS|130|6|我的心等候主，勝於守夜的等候天亮， 勝於守夜的等候天亮。
PS|130|7|以色列 啊，你當仰望耶和華， 因耶和華有慈愛，有豐盛的救恩。
PS|130|8|他必救贖 以色列 脫離一切的罪孽。
PS|131|1|耶和華啊，我的心不狂妄， 我的眼不高傲； 重大和測不透的事， 我也不敢行。
PS|131|2|我使我心安穩平靜，好像母親懷中斷奶的孩子； 我的心在我裏面如同斷過奶的孩子。
PS|131|3|以色列 啊，你當仰望耶和華， 從今時直到永遠！
PS|132|1|耶和華啊，求你記念 大衛 ， 記念他所受的一切苦難！
PS|132|2|他怎樣向耶和華起誓， 向 雅各 的大能者許願：
PS|132|3|「我必不進我的帳幕， 也不上我的床鋪；
PS|132|4|我不容我的眼睛睡覺， 也不容我的眼皮打盹；
PS|132|5|直等到我為耶和華尋得所在， 為 雅各 的大能者尋得居所。」
PS|132|6|我們聽說約櫃在 以法他 ， 我們在 雅珥 的田野尋見它。
PS|132|7|「我們要進他的居所， 在他腳凳前下拜。」
PS|132|8|耶和華啊，求你興起， 與你有能力的約櫃同入安歇之所！
PS|132|9|願你的祭司披上公義！ 願你的聖民歡呼！
PS|132|10|求你因你僕人 大衛 的緣故， 不要厭棄你的受膏者！
PS|132|11|耶和華憑信實向 大衛 起了誓，絕不改變： 「我要立你身所生的 坐在你的寶座上。
PS|132|12|你的眾子若謹守我的約和我所教導他們的法度， 他們的子孫必永遠坐在你的寶座上。」
PS|132|13|因為耶和華揀選了 錫安 ， 願意當作自己的居所：
PS|132|14|「這是我永遠安歇之所； 我要住在這地方，因為我願意在這裏。
PS|132|15|我要賜福使糧食豐足， 使其中的貧窮人飽享食物。
PS|132|16|我要使祭司披上救恩， 聖民就要大聲歡呼！
PS|132|17|在那裏我要使 大衛 的角茁壯， 為我的受膏者預備明燈。
PS|132|18|我要使他的仇敵披上羞恥； 但他的冠冕要在他頭上發光。」
PS|133|1|看哪，弟兄和睦同住 是何等的善，何等的美！
PS|133|2|這好比那貴重的油澆在 亞倫 的頭上， 流到鬍鬚，又流到他的衣襟；
PS|133|3|又好比 黑門 的甘露降在 錫安山 ； 因為在那裏有耶和華所命定的福，就是永遠的生命。
PS|134|1|來，稱頌耶和華！ 夜間侍立在耶和華殿中，耶和華的僕人，
PS|134|2|當向聖所舉手， 稱頌耶和華！
PS|134|3|願造天地的耶和華 從 錫安 賜福給你們！
PS|135|1|哈利路亞！ 你們要讚美耶和華的名！ 侍立在耶和華殿中，耶和華的僕人， 侍立在我們上帝殿院中的，要讚美他！
PS|135|2|
PS|135|3|你們要讚美耶和華， 因耶和華本為善； 要歌頌他的名， 因為這是美好的。
PS|135|4|耶和華揀選 雅各 歸自己， 揀選 以色列 作他寶貴的產業。
PS|135|5|我知道耶和華本為大， 也知道我們的主超乎萬神之上。
PS|135|6|在天，在地，在海洋，在各深淵， 耶和華都隨自己的旨意而行。
PS|135|7|他使雲霧從地極上騰， 造電隨雨而閃， 從倉庫中吹出風來。
PS|135|8|他將 埃及 頭生的， 連人帶牲畜都擊殺了。
PS|135|9|埃及 啊，他施行神蹟奇事， 在你們中間，在法老和他所有臣僕身上。
PS|135|10|他擊打許多國家， 殺戮大能的君王，
PS|135|11|就是 亞摩利 王 西宏 、 巴珊 王 噩 ， 和 迦南 一切的國度，
PS|135|12|他賞賜他們的地為業， 作為自己百姓 以色列 的產業。
PS|135|13|耶和華啊，你的名字存到永遠！ 耶和華啊，你的稱號 存到萬代！
PS|135|14|耶和華要為自己的百姓伸冤， 為自己的僕人發憐憫。
PS|135|15|外邦的偶像是金的，是銀的， 是人手所造的，
PS|135|16|有口卻不能言， 有眼卻不能看，
PS|135|17|有耳卻不能聽， 口中也沒有氣息。
PS|135|18|造它們的要像它們一樣， 凡靠它們的也必如此。
PS|135|19|以色列 家啊，要稱頌耶和華！ 亞倫 家啊，要稱頌耶和華！
PS|135|20|利未 家啊，要稱頌耶和華！ 你們敬畏耶和華的，要稱頌耶和華！
PS|135|21|住在 耶路撒冷 的、 錫安 的耶和華， 是應當稱頌的。 哈利路亞！
PS|136|1|你們要稱謝耶和華，因他本為善； 他的慈愛永遠長存。
PS|136|2|你們要稱謝萬神之神， 因他的慈愛永遠長存。
PS|136|3|你們要稱謝萬主之主， 因他的慈愛永遠長存。
PS|136|4|稱謝那惟一能行大 奇事的， 因他的慈愛永遠長存。
PS|136|5|稱謝那用智慧造天的， 因他的慈愛永遠長存。
PS|136|6|稱謝那鋪地在水以上的， 因他的慈愛永遠長存。
PS|136|7|稱謝那造成大光的， 因他的慈愛永遠長存。
PS|136|8|他造太陽管白晝， 因他的慈愛永遠長存。
PS|136|9|他造月亮星宿管黑夜， 因他的慈愛永遠長存。
PS|136|10|稱謝那擊殺 埃及 凡是頭生的， 因他的慈愛永遠長存。
PS|136|11|他以大能的手和伸出來的膀臂， 因他的慈愛永遠長存。 領 以色列 人從 埃及 人中出來， 因他的慈愛永遠長存。
PS|136|12|
PS|136|13|稱謝那分裂 紅海 的， 因他的慈愛永遠長存。
PS|136|14|他領 以色列 從其中經過， 因他的慈愛永遠長存；
PS|136|15|卻把法老和他的軍隊推落 紅海 裏， 因他的慈愛永遠長存。
PS|136|16|稱謝那引導自己子民行走曠野的， 因他的慈愛永遠長存。
PS|136|17|稱謝那擊殺大君王的， 因他的慈愛永遠長存。
PS|136|18|他殺戮威武的君王， 因他的慈愛永遠長存；
PS|136|19|殺戮 亞摩利 王 西宏 ， 因他的慈愛永遠長存；
PS|136|20|殺戮 巴珊 王 噩 ， 因他的慈愛永遠長存。
PS|136|21|他賞賜他們的地為業， 因他的慈愛永遠長存；
PS|136|22|作為他僕人 以色列 的產業， 因他的慈愛永遠長存。
PS|136|23|我們身處卑微，他顧念我們， 因他的慈愛永遠長存。
PS|136|24|他搭救我們脫離敵人， 因他的慈愛永遠長存。
PS|136|25|凡有血有肉的，他賜糧食， 因他的慈愛永遠長存。
PS|136|26|你們要稱謝天上的上帝， 因他的慈愛永遠長存。
PS|137|1|我們在 巴比倫 河邊， 坐在那裏，追想 錫安 ，就哭了。
PS|137|2|在一排柳樹中， 我們掛上我們的豎琴。
PS|137|3|擄掠我們的在那裏 要我們唱歌； 搶奪我們的要我們為他們作樂： 「給我們唱一首 錫安 的歌吧！」
PS|137|4|我們怎能在外邦之土 唱耶和華的歌呢？
PS|137|5|耶路撒冷 啊，我若忘記你， 寧願我的右手枯萎；
PS|137|6|我若不記得你，不看你過於我最喜樂的， 寧願我的舌頭貼於上膛！
PS|137|7|耶路撒冷 攻破的日子， 以東 人說：「拆毀！拆毀！ 直拆到根基！」 耶和華啊，求你記得！
PS|137|8|將要被滅的 巴比倫 哪， 用你待我們的惡行報復你的，那人有福了。
PS|137|9|抓起你的嬰孩摔在磐石上的， 那人有福了。
PS|138|1|我要一心稱謝你 ， 在諸神面前歌頌你。
PS|138|2|我要向你的聖殿下拜， 我要因你的慈愛和信實頌揚你的名； 因你使你的名和你的言語顯為大， 超乎一切 。
PS|138|3|我呼求的日子，你應允我， 使我壯膽，心裏有能力。
PS|138|4|耶和華啊，地上的君王都要稱謝你， 因他們聽見了你口中的言語。
PS|138|5|他們要歌頌耶和華的作為， 因耶和華大有榮耀。
PS|138|6|耶和華雖崇高，卻看顧卑微的人； 驕傲的人，他從遠處即能認出。
PS|138|7|我雖困在患難中，你必將我救活； 我的仇敵發怒，你必伸手抵擋他們， 你的右手也必拯救我。
PS|138|8|耶和華必成全他在我身上的旨意； 耶和華啊，你的慈愛永遠長存！ 求你不要離棄你手所造的。
PS|139|1|耶和華啊，你已經鑒察我， 認識我。
PS|139|2|我坐下，我起來，你都曉得； 你從遠處知道我的意念。
PS|139|3|我行路，我躺臥，你都細察； 你也深知我一切所行的。
PS|139|4|耶和華啊，我舌頭上的話， 你沒有一句不知道的。
PS|139|5|你前後環繞我， 按手在我身上。
PS|139|6|這樣的知識奇妙，是我不能測的； 至高，是我不能及的。
PS|139|7|我往哪裏去，躲避你的靈？ 我往哪裏逃，躲避你的面？
PS|139|8|我若升到天上，你在那裏； 我若躺在陰間，你也在那裏。
PS|139|9|我若展開清晨的翅膀， 飛到海極居住，
PS|139|10|就是在那裏，你的手必引導我， 你的右手也必扶持我。
PS|139|11|我若說「黑暗必定壓碎我， 我周圍的亮光必成為黑夜」，
PS|139|12|黑暗對你不再是黑暗， 黑夜卻如白晝發亮。 黑暗和光明， 在你看來都是一樣。
PS|139|13|我的肺腑是你所造的， 我在母腹中，你已編織 我。
PS|139|14|我要稱謝你，因我受造奇妙可畏， 你的作為奇妙，這是我心深知道的。
PS|139|15|我在暗中受造，在地的深處被塑造； 那時，我的形體並不向你隱藏。
PS|139|16|我未成形的體質， 你的眼早已看見了； 你所定的日子，我尚未度一日， 都在你的冊子寫上了。
PS|139|17|上帝啊，你的意念向我何等寶貴！ 其數何等眾多！
PS|139|18|我若數點，比海沙更多； 我睡醒的時候，仍和你同在。
PS|139|19|上帝啊，惟願你殺戮惡人； 你們好流人血的，離開我去吧！
PS|139|20|他們說惡言頂撞你， 你的仇敵妄稱你的名 。
PS|139|21|耶和華啊，恨惡你的，我豈不恨惡他們嗎？ 攻擊你的，我豈不憎惡他們嗎？
PS|139|22|我恨惡他們到極點， 以他們為我的仇敵。
PS|139|23|上帝啊，求你鑒察我，知道我的心思， 試煉我，知道我的意念；
PS|139|24|看在我裏面有甚麼惡行沒有， 引導我走永生的道路。
PS|140|1|耶和華啊，求你救我脫離邪惡的人， 保護我脫離殘暴的人！
PS|140|2|他們心中圖謀奸惡， 日日不停挑起戰爭。
PS|140|3|他們的舌頭銳利如蛇， 嘴唇裏有毒蛇的毒液。（細拉）
PS|140|4|耶和華啊，求你庇護我脫離惡人的手， 保護我脫離殘暴的人，他們想要推倒我。
PS|140|5|驕傲的人為我暗設羅網和繩索； 他們在路旁張開網，為我設下圈套。（細拉）
PS|140|6|我曾對耶和華說：「你是我的上帝。」 耶和華啊，求你側耳聽我懇求的聲音！
PS|140|7|主－耶和華、我救恩的力量啊， 在戰爭的日子，你遮蔽了我的頭。
PS|140|8|耶和華啊，求你不要遂惡人的心願； 不要成就他們的計謀，免得他們自高。（細拉）
PS|140|9|至於那些昂首圍困我的人， 願他們嘴唇的奸惡陷害 自己！
PS|140|10|願他們被丟在火中，火炭落在他們身上； 願他們被拋在深坑裏，不能再起來！
PS|140|11|願說惡言的人在地上站立不住； 願禍患獵取殘暴的人，把他打倒。
PS|140|12|我知道耶和華必為困苦人伸冤， 為貧窮人辯護。
PS|140|13|義人必頌揚你的名， 正直人要在你面前居住。
PS|141|1|耶和華啊，我曾求告你， 求你快快臨到我這裏！ 我求告你的時候， 求你側耳聽我的聲音！
PS|141|2|願我的禱告如香呈到你面前！ 願我的手舉起 ，如獻晚祭！
PS|141|3|耶和華啊，求你看守我的口， 把守我的嘴唇！
PS|141|4|不要使我的心偏向邪惡的事， 以致我和作惡的人一同行惡； 也不叫我吃他們的美食。
PS|141|5|任憑義人擊打我，這算為仁慈； 任憑他責備我，這算為頭上的膏油； 我的頭不躲閃。 人正行惡的時候，我仍要祈禱。
PS|141|6|他們的審判官被扔在巖下， 他們就要聽我的話，因為這話甘甜。
PS|141|7|我們的 骨頭散落在陰間的口， 就像人耕田刨地 一樣。
PS|141|8|主－耶和華啊，我的眼目仰望你； 我投靠你，求你不要使我的性命陷入危險！
PS|141|9|求你保護我脫離惡人為我設的羅網 和作惡之人的圈套！
PS|141|10|願惡人落在自己的網中， 我卻得以逃脫。
PS|142|1|我出聲哀告耶和華， 出聲懇求耶和華。
PS|142|2|我在他面前傾訴我的苦情， 在他面前陳說我的患難。
PS|142|3|我的靈在我裏面發昏的時候， 你知道我的道路。 在我所行的路上， 人為我暗設羅網。
PS|142|4|求你留意向我右邊觀看， 無人認識我； 我無避難之處， 也無人眷顧我。
PS|142|5|耶和華啊，我曾向你哀求。 我說：「你是我的避難所， 在活人之地，你是我的福分。」
PS|142|6|求你留心聽我的呼求， 因我落到極卑微之地； 求你救我脫離迫害我的人， 因為他們比我強盛。
PS|142|7|求你從被囚之地領我出來， 我好頌揚你的名。 義人必環繞我， 因為你用厚恩待我。
PS|143|1|耶和華啊，求你聽我的禱告， 側耳聽我的懇求，憑你的信實和公義應允我。
PS|143|2|求你不要審問僕人， 因為在你面前，凡活著的人沒有一個是義的。
PS|143|3|因為仇敵迫害我， 將我打倒在地， 使我住在幽暗之處， 像死了許久的人一樣。
PS|143|4|我的靈在我裏面發昏， 我的心在我裏面顫慄。
PS|143|5|我追想古時之日，思想你的一切作為， 默念你手的工作。
PS|143|6|我向你舉手， 我的心渴想你，如乾旱之地盼雨一樣。（細拉）
PS|143|7|耶和華啊，求你速速應允我！ 我的心神耗盡！ 求你不要轉臉不顧我， 免得我像那些下入地府的人一樣。
PS|143|8|求你使我清晨得聽你慈愛的聲音， 因我倚靠你； 求你使我知道當走的路， 因我的心仰望你。
PS|143|9|耶和華啊，求你救我脫離我的仇敵！ 我往你那裏藏身。
PS|143|10|求你指教我遵行你的旨意， 因你是我的上帝； 願你至善的靈 引我到平坦之地。
PS|143|11|耶和華啊，求你為你名的緣故將我救活， 憑你的公義，將我從患難中領出來，
PS|143|12|憑你的慈愛剪除我的仇敵， 滅絕所有苦待我的人，因我是你的僕人。
PS|144|1|耶和華─我的磐石是應當稱頌的！ 他教導我的手爭戰， 教導我的指頭打仗。
PS|144|2|他是我慈愛的主、我的山寨、 我的碉堡、我的救主、 我的盾牌，是我所投靠的。 他使我的百姓 服在我以下。
PS|144|3|耶和華啊，人算甚麼，你竟認識他！ 世人算甚麼，你竟顧念他！
PS|144|4|人不過像一口氣， 他的年日如影消逝。
PS|144|5|耶和華啊，求你使天下垂，親自降臨； 求你摸山，使山冒煙。
PS|144|6|求你發出閃電，使仇敵四散， 射出你的箭，使他們混亂。
PS|144|7|求你從高處伸手救拔我， 救我脫離大水，脫離外邦人的手。
PS|144|8|他們的口說謊話， 他們的右手起假誓。
PS|144|9|上帝啊，我要向你唱新歌， 用十弦瑟向你歌頌。
PS|144|10|你是那拯救君王的， 你是那救僕人 大衛 脫離害命之刀的。
PS|144|11|求你救拔我， 救我脫離外邦人的手。 他們的口說謊話， 他們的右手起假誓。
PS|144|12|我們的兒子從幼年好像樹苗長大， 我們的女兒如同房角石，按照建宮殿的樣式鑿成。
PS|144|13|我們的倉盈滿，能供應各種糧食； 我們的羊在田野孳生千萬。
PS|144|14|我們的牲口馱滿貨物， 沒有人闖進來搶奪， 也沒有人出去爭戰； 我們的街市上也沒有哭號的聲音。
PS|144|15|這樣情況的百姓有福了！ 以耶和華為他們上帝的百姓有福了！
PS|145|1|我的上帝、我的王啊、我要尊崇你！ 我要永永遠遠稱頌你的名！
PS|145|2|我要天天稱頌你， 也要永永遠遠讚美你的名！
PS|145|3|耶和華本為大，該受大讚美， 其大無法測度。
PS|145|4|這一代要對那一代頌讚你的作為， 他們要傳揚你的大能。
PS|145|5|他們要述說你威嚴榮耀的尊榮， 我要默念你奇妙的作為 。
PS|145|6|人要傳講你可畏的能力， 我也要傳揚你的偉大。
PS|145|7|他們要將你可記念的大恩傳開， 並要高唱你的公義。
PS|145|8|耶和華有恩惠，有憐憫， 不輕易發怒，大有慈愛。
PS|145|9|耶和華善待萬有， 他的憐憫覆庇他一切所造的。
PS|145|10|耶和華啊，你一切所造的都要稱謝你， 你的聖民也要稱頌你。
PS|145|11|他們要傳講你國度的榮耀， 談論你的大能，
PS|145|12|好讓世人知道你大能的作為 和你國度威嚴的榮耀。
PS|145|13|你的國是永遠的國！ 你執掌的權柄存到萬代！ 耶和華一切的話信實可靠， 他一切的作為都有慈愛 。
PS|145|14|耶和華扶起所有跌倒的， 扶起所有被壓下的。
PS|145|15|萬有的眼目都仰望你， 你按時給他們食物。
PS|145|16|你張手， 使一切有生命的都隨願飽足。
PS|145|17|耶和華一切所行的，無不公義， 一切所做的，都有慈愛。
PS|145|18|耶和華臨近凡求告他的， 臨近所有誠心求告他的人。
PS|145|19|敬畏他的，他必成就他們的心願， 也必聽他們的呼求，拯救他們。
PS|145|20|耶和華保護凡愛他的人， 卻要滅絕所有的惡人。
PS|145|21|我的口要述說讚美耶和華的話； 惟願有血肉之軀的都永永遠遠稱頌他的聖名。
PS|146|1|哈利路亞！ 我的心哪，你要讚美耶和華！
PS|146|2|我一生要讚美耶和華！ 我還活著的時候要歌頌我的上帝！
PS|146|3|你們不要倚靠君王，不要倚靠世人， 他一點也不能幫助。
PS|146|4|他的氣一斷，就歸回塵土， 他所打算的，當日就消滅了。
PS|146|5|以 雅各 的上帝為幫助、 仰望耶和華－他上帝的，這人有福了！
PS|146|6|耶和華造天、地、海和其中的萬物， 他守信實，直到永遠。
PS|146|7|他為受欺壓的伸冤， 賜食物給飢餓的人。 耶和華釋放被囚的，
PS|146|8|耶和華開了盲人的眼睛， 耶和華扶起被壓下的人， 耶和華喜愛義人。
PS|146|9|耶和華保護寄居的，扶持孤兒和寡婦， 卻使惡人的道路彎曲。
PS|146|10|耶和華要作王，直到永遠！ 錫安 哪，你的上帝要作王，直到萬代！ 哈利路亞！
PS|147|1|哈利路亞！ 歌頌我們的上帝是美善的， 因為他是美好的，讚美他是合宜的。
PS|147|2|耶和華建造 耶路撒冷 ， 聚集 以色列 中被趕散的人。
PS|147|3|他醫好傷心的人， 包紮他們的傷處。
PS|147|4|他數點星宿的數目， 一一稱它們的名。
PS|147|5|我們的主本為大，大有能力， 他的智慧無法測度。
PS|147|6|耶和華扶持謙卑的人， 將惡人傾覆於地。
PS|147|7|你們要以感謝向耶和華歌唱， 用琴向我們的上帝歌頌。
PS|147|8|他用密雲遮天，為地預備雨水， 使草生長在山上。
PS|147|9|他賜食物給走獸 和啼叫的小烏鴉。
PS|147|10|他不喜悅馬的力大， 不喜愛人的腿快。
PS|147|11|耶和華喜愛敬畏他 和盼望他慈愛的人。
PS|147|12|耶路撒冷 啊，要頌讚耶和華！ 錫安 哪，要讚美你的上帝！
PS|147|13|因為他堅固了你的門閂， 賜福給你中間的兒女。
PS|147|14|他使你境內平安， 用上好的麥子使你滿足。
PS|147|15|他向大地發出命令， 他的話速速頒行。
PS|147|16|他降雪如羊毛， 撒霜如灰燼。
PS|147|17|他擲下冰雹如碎渣， 他發出寒冷，誰能當得起呢？
PS|147|18|他一出令，這些就都融化， 他使風颳起，水便流動。
PS|147|19|他將他的道指示 雅各 ， 將他的律例典章指示 以色列 。
PS|147|20|他未曾這樣對待別國， 至於他的典章，他們向來都不知道 。 哈利路亞！
PS|148|1|哈利路亞！ 你們要從天上讚美耶和華， 在高處讚美他！
PS|148|2|他的眾使者啊，要讚美他！ 他的諸軍啊，都要讚美他！
PS|148|3|太陽月亮啊，要讚美他！ 放光的星宿啊，都要讚美他！
PS|148|4|天上的天和天上的水啊， 你們都要讚美他！
PS|148|5|願這些都讚美耶和華的名！ 因他一吩咐就都造成。
PS|148|6|他將這些設定，直到永永遠遠； 他訂了律例，不能廢去。
PS|148|7|你們哪，都當讚美耶和華： 地上一切所有的，大魚和深洋，
PS|148|8|火和冰雹，雪和霧氣， 成就他命令的狂風，
PS|148|9|大山和小山， 結果子的樹木和一切香柏樹，
PS|148|10|野獸和一切牲畜， 昆蟲和飛鳥，
PS|148|11|世上的君王和萬民， 領袖和世上所有的審判官，
PS|148|12|少年和少女， 老人和孩童，
PS|148|13|願這些都讚美耶和華的名！ 因為獨有他的名被尊崇，他的榮耀在天地之上。
PS|148|14|他高舉自己百姓的角， 使他的聖民 以色列 人，就是與他相近的百姓得榮耀 。 哈利路亞！
PS|149|1|哈利路亞！ 你們要向耶和華唱新歌， 在聖民的會中讚美他！
PS|149|2|願 以色列 因造他的主歡喜！ 願 錫安 的民因他們的王快樂！
PS|149|3|願他們跳舞讚美他的名， 擊鼓彈琴歌頌他！
PS|149|4|因為耶和華喜愛自己的百姓， 他要用救恩當作謙卑人的妝飾。
PS|149|5|願聖民因所得的榮耀歡樂！ 願他們在床上也歡呼！
PS|149|6|願他們口中稱頌上帝為至高， 手裏有兩刃的劍，
PS|149|7|為要報復列國， 懲罰萬民。
PS|149|8|要用鏈子捆他們的君王， 用鐵鐐鎖他們的貴族，
PS|149|9|要在他們身上施行所記錄的審判。 他的聖民都享榮耀。 哈利路亞！
PS|150|1|哈利路亞！ 你們要在上帝的聖所讚美他！ 在他顯能力的穹蒼讚美他！
PS|150|2|要因他大能的作為讚美他， 因他極其偉大讚美他！
PS|150|3|要用角聲讚美他， 鼓瑟彈琴讚美他！
PS|150|4|擊鼓跳舞讚美他！ 用絲弦的樂器和簫的聲音讚美他！
PS|150|5|用大響的鈸讚美他！ 用高聲的鈸讚美他！
PS|150|6|凡有生命的都要讚美耶和華！ 哈利路亞！
