JAS|1|1|Яків, раб Бога й Господа Ісуса Христа, дванадцятьом племенам, які в Розпорошенні, вітаю я вас!
JAS|1|2|Майте, брати мої, повну радість, коли впадаєте в усілякі випробовування,
JAS|1|3|знаючи, що досвідчення вашої віри дає терпеливість.
JAS|1|4|А терпеливість нехай має чин досконалий, щоб ви досконалі та бездоганні були, і недостачі ні в чому не мали.
JAS|1|5|А якщо кому з вас не стачає мудрости, нехай просить від Бога, що всім дає просто, та не докоряє, і буде вона йому дана.
JAS|1|6|Але нехай просить із вірою, без жадного сумніву. Бо хто має сумнів, той подібний до морської хвилі, яку жене й кидає вітер.
JAS|1|7|Нехай бо така людина не гадає, що дістане що від Господа.
JAS|1|8|Двоєдушна людина непостійна на всіх дорогах своїх.
JAS|1|9|А понижений брат нехай хвалиться високістю своєю,
JAS|1|10|а багатий пониженням своїм, бо він промине, як той цвіт трав'яний,
JAS|1|11|бо сонце зійшло зо спекотою, і траву посушило, і відпав цвіт її, і зникла краса її виду... Так само зів'яне й багатий у дорогах своїх!
JAS|1|12|Блаженна людина, що витерпить пробу, бо, бувши випробувана, дістане вінця життя, якого Господь обіцяв тим, хто любить Його.
JAS|1|13|Випробовуваний, хай не каже ніхто: Я від Бога спокушуваний. Бо Бог злом не спокушується, і нікого Він Сам не спокушує.
JAS|1|14|Але кожен спокушується, як надиться й зводиться пожадливістю власною.
JAS|1|15|Пожадливість потому, зачавши, народжує гріх, а зроблений гріх народжує смерть.
JAS|1|16|Не обманюйтесь, брати мої любі!
JAS|1|17|Усяке добре давання та дар досконалий походить згори від Отця світил, що в Нього нема переміни чи тіні відміни.
JAS|1|18|Захотівши, Він нас породив словом правди, щоб ми стали якимсь первопочином творів Його.
JAS|1|19|Отож, мої брати любі, нехай буде кожна людина швидка послухати, забарна говорити, повільна на гнів.
JAS|1|20|Бо гнів людський не чинить правди Божої.
JAS|1|21|Тому то відкиньте всіляку нечисть та залишок злоби, і прийміть із лагідністю всіяне слово, що може спасти ваші душі.
JAS|1|22|Будьте ж виконавцями слова, а не слухачами самими, що себе самих обманюють.
JAS|1|23|Бо хто слухач слова, а не виконавець, той подібний людині, що риси обличчя свого розглядає у дзеркалі,
JAS|1|24|бо розгляне себе та й відійде, і зараз забуде, яка вона є.
JAS|1|25|А хто заглядає в закон досконалий, закон волі, і в нім пробуває, той не буде забудько слухач, але виконавець діла, і він буде блаженний у діянні своїм!
JAS|1|26|Коли ж хто гадає, що він побожний, і свого язика не вгамовує, та своє серце обманює, марна побожність того!
JAS|1|27|Чиста й непорочна побожність перед Богом і Отцем оця: зглянутися над сиротами та вдовицями в утисках їхніх, себе берегти чистим від світу.
JAS|2|1|Брати мої, не зважаючи на обличчя, майте віру в нашого Господа слави, Ісуса Христа.
JAS|2|2|Бо коли до вашого зібрання ввійде чоловік із золотим перснем, у шаті блискучій, увійде й бідар у вбогім вбранні,
JAS|2|3|і ви поглянете на того, хто в шаті блискучій, і скажете йому: Ти сідай вигідно отут, а бідареві прокажете: Ти стань там, чи сідай собі тут на підніжку моїм,
JAS|2|4|то чи не стало між вами поділення, і не стали ви злодумними суддями?
JAS|2|5|Послухайте, мої брати любі, чи ж не вибрав Бог бідарів цього світу за багатих вірою й за спадкоємців Царства, яке обіцяв Він тим, хто любить Його?
JAS|2|6|А ви бідаря зневажили! Хіба не багачі переслідують вас, хіба не вони тягнуть вас на суди?
JAS|2|7|Хіба не вони зневажають те добре ім'я, що ви ним називаєтесь?
JAS|2|8|Коли ви Закона Царського виконуєте, за Писанням: Люби свого ближнього, як самого себе, то ви робите добре.
JAS|2|9|Коли ж дивитеся на обличчя, то чините гріх, бо Закон удоводнює, що ви винуватці.
JAS|2|10|Бо хто всього Закона виконує, а згрішить в одному, той винним у всьому стає.
JAS|2|11|Бо Той, Хто сказав: Не чини перелюбства, також наказав: Не вбивай. А хоч ти перелюбства не чиниш, а вб'єш, то ти переступник Закону.
JAS|2|12|Отак говоріть і отак чиніть, як такі, що будете суджені законом волі.
JAS|2|13|Бо суд немилосердний на того, хто не вчинив милосердя. Милосердя бо ставиться вище за суд.
JAS|2|14|Яка користь, брати мої, коли хто говорить, що має віру, але діл не має? Чи може спасти його віра?
JAS|2|15|Коли ж брат чи сестра будуть нагі, і позбавлені денного покорму,
JAS|2|16|а хтонебудь із вас до них скаже: Ідіть з миром, грійтесь та їжте, та не дасть їм потрібного тілу, що ж то поможе?
JAS|2|17|Так само й віра, коли діл не має, мертва в собі!
JAS|2|18|Але скаже хтонебудь: Маєш ти віру, а я маю діла; покажи мені віру свою без діл твоїх, а я покажу тобі віру свою від діл моїх.
JAS|2|19|Чи віруєш ти, що Бог один? Добре робиш! Та й демони вірують, і тремтять.
JAS|2|20|Чи хочеш ти знати, о марна людино, що віра без діл мертва?
JAS|2|21|Авраам, отець наш, чи він не з діл виправданий був, як поклав був на жертівника свого сина Ісака?
JAS|2|22|Чи ти бачиш, що віра помогла його ділам, і вдосконалилась віра із діл?
JAS|2|23|І здійснилося Писання, що каже: Авраам же ввірував Богові, і це йому зараховане в праведність, і був названий він другом Божим.
JAS|2|24|Отож, чи ви бачите, що людина виправдується від діл, а не тільки від віри?
JAS|2|25|Чи так само і блудниця Рахав не з діл виправдалась, коли прийняла посланців, і дорогою іншою випустила?
JAS|2|26|Бо як тіло без духа мертве, так і віра без діл мертва!
JAS|3|1|Не багато-хто ставайте, брати мої, учителями, знавши, що більший осуд приймемо.
JAS|3|2|Бо багато ми всі помиляємось. Коли хто не помиляється в слові, то це муж досконалий, спроможний приборкувати й усе тіло.
JAS|3|3|От і коням вкладаєм уздечки до рота, щоб корилися нам, і ми всім їхнім тілом керуємо.
JAS|3|4|От і кораблі, хоч які величезні та гнані вітрами жорстокими, проте найменшим стерном скеровуються, куди хоче стерничий.
JAS|3|5|Так само й язик, малий член, але хвалиться вельми! Ось маленький огонь, а запалює величезного ліса!
JAS|3|6|І язик то огонь. Як світ неправости, поставлений так поміж нашими членами, язик сквернить усе тіло, запалює круг життя, і сам запалюється від геєнни.
JAS|3|7|Бо всяка природа звірів і пташок, гадів і морських потвор приборкується, і приборкана буде природою людською,
JAS|3|8|та не може ніхто із людей язика вгамувати, він зло безупинне, він повний отрути смертельної!
JAS|3|9|Ним ми благословляємо Бога й Отця, і ним проклинаєм людей, що створені на Божу подобу.
JAS|3|10|Із тих самих уст виходить благословення й прокляття. Не повинно, брати мої, щоб так це було!
JAS|3|11|Хіба з одного отвору виходить вода солодка й гірка?
JAS|3|12|Хіба може, брати мої, фіґове дерево родити оливки, або виноград фіґи? Солодка вода не тече з солонця.
JAS|3|13|Хто мудрий і розумний між вами? Нехай він покаже діла свої в лагідній мудрості добрим поводженням!
JAS|3|14|Коли ж гірку заздрість та сварку ви маєте в серці своєму, то не величайтесь та не говоріть неправди на правду,
JAS|3|15|це не мудрість, що ніби зверху походить вона, але земна, тілесна та демонська.
JAS|3|16|Бо де заздрість та сварка, там безлад та всяка зла річ!
JAS|3|17|А мудрість, що зверху вона, насамперед чиста, а потім спокійна, лагідна, покірлива, повна милосердя та добрих плодів, безстороння та нелукава.
JAS|3|18|А плід правди сіється творцями миру.
JAS|4|1|Звідки війни та свари між вами? Чи не звідси, від ваших пожадливостей, які в ваших членах воюють?
JAS|4|2|Бажаєте ви та й не маєте, убиваєте й заздрите та досягнути не можете, сваритеся та воюєте та не маєте, бо не прохаєте,
JAS|4|3|прохаєте та не одержуєте, бо прохаєте на зле, щоб ужити на розкоші свої.
JAS|4|4|Перелюбники та перелюбниці, чи ж ви не знаєте, що дружба зо світом то ворожнеча супроти Бога? Бо хто хоче бути світові приятелем, той ворогом Божим стається.
JAS|4|5|Чи ви думаєте, що даремно Писання говорить: Жадає аж до заздрости дух, що в нас пробуває?
JAS|4|6|Та ще більшу благодать дає, через що й промовляє: Бог противиться гордим, а смиренним дає благодать.
JAS|4|7|Тож підкоріться Богові та спротивляйтесь дияволові, то й утече він від вас.
JAS|4|8|Наблизьтесь до Бога, то й Бог наблизиться до вас. Очистьте руки, грішні, та серця освятіть, двоєдушні!
JAS|4|9|Журіться, сумуйте та плачте! Хай обернеться сміх ваш у плач, а радість у сум!
JAS|4|10|Упокоріться перед Господнім лицем, і Він вас підійме!
JAS|4|11|Не обмовляйте, брати, один одного! Бо хто брата свого обмовляє або судить брата, той Закона обмовляє та судить Закона. А коли ти Закона осуджуєш, то ти не виконавець Закона, але суддя.
JAS|4|12|Один Законодавець і Суддя, що може спасти й погубити. А ти хто такий, що осуджуєш ближнього?
JAS|4|13|А ну тепер ви, що говорите: Сьогодні чи взавтра ми підем у те чи те місто, і там рік проживемо, та будемо торгувати й заробляти,
JAS|4|14|ви, що не відаєте, що трапиться взавтра, яке ваше життя? Бо це пара, що на хвильку з'являється, а потім зникає!...
JAS|4|15|Замість того, щоб вам говорити: Як схоче Господь та будемо живі, то зробимо це або те.
JAS|4|16|А тепер ви хвалитеся в своїх гордощах, лиха всяка подібна хвальба!
JAS|4|17|Отож, хто знає, як чинити добро, та не чинить, той має гріх!
JAS|5|1|А ну ж тепер ви, багачі, плачте й ридайте над лихом своїм, що вас має спіткати:
JAS|5|2|ваше багатство згнило, а ваші вбрання міль поїла!
JAS|5|3|Золото ваше та срібло поіржавіло, а їхня іржа буде свідчити проти вас, і поїсть ваше тіло, немов той огонь! Ви скарби зібрали собі на останні дні!
JAS|5|4|Ось голосить заплата, що ви затримали в робітників, які жали на ваших полях, і голосіння женців досягли вух Господа Саваота!
JAS|5|5|Ви розкошували на землі й насолоджувались, серця свої вигодували, немов би на день заколення.
JAS|5|6|Ви Праведного засудили й убили, Він вам не противився!
JAS|5|7|Отож, браття, довготерпіть аж до приходу Господа! Ось чекає рільник дорогоцінного плоду землі, довготерпить за нього, аж поки одержить дощ ранній та пізній.
JAS|5|8|Довготерпіть же й ви, зміцніть серця ваші, бо наблизився прихід Господній!
JAS|5|9|Не нарікайте один на одного, браття, щоб вас не засуджено, он Суддя стоїть перед дверима!
JAS|5|10|Візьміть, браття, пророків за приклад страждання та довготерпіння, вони промовляли Господнім Ім'ям!
JAS|5|11|Отож, за блаженних ми маємо тих, хто витерпів. Ви чули про Йовове терпіння та бачили Господній кінець його, що вельми Господь милостивий та щедрий.
JAS|5|12|А найперше, браття мої, не кляніться ні небом, ані землею, і ніякою іншою клятвою! Слово ж ваше хай буде: Так, так та Ні, ні, щоб не впасти вам в осуд.
JAS|5|13|Чи страждає хто з вас? Нехай молиться! Чи тішиться хтось? Хай співає псалми!
JAS|5|14|Чи хворіє хто з вас? Хай покличе пресвітерів Церкви, і над ним хай помоляться, намастивши його оливою в Господнє Ім'я,
JAS|5|15|і молитва віри вздоровить недужого, і Господь його підійме, а коли він гріхи був учинив, то вони йому простяться.
JAS|5|16|Отже, признавайтесь один перед одним у своїх прогріхах, і моліться один за одного, щоб вам уздоровитись. Бо дуже могутня ревна молитва праведного!
JAS|5|17|Ілля був людина, подібна до нас пристрастями, і він помолився молитвою, щоб дощу не було, і дощу не було на землі аж три роки й шість місяців...
JAS|5|18|І він знов помолився, і дощу дало небо, а земля вродила свій плід!
JAS|5|19|Браття мої, коли хто з-поміж вас заблудить від правди, і його хто наверне,
JAS|5|20|хай знає, що той, хто грішника навернув від його блудної дороги, той душу його спасає від смерти та безліч гріхів покриває!
