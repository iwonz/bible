PHIL|1|1|基督耶穌的僕人 保羅 和 提摩太 寫信給住 腓立比 、在基督耶穌裏的眾聖徒，以及諸位監督和執事。
PHIL|1|2|願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
PHIL|1|3|我每逢想念你們，就感謝我的上帝，
PHIL|1|4|每逢為你們眾人祈求的時候，總是歡歡喜喜地祈求，
PHIL|1|5|因為從第一天直到如今，你們都同心合意興旺福音。
PHIL|1|6|我深信，那在你們心裏動了美好工作的，到了耶穌基督的日子必完成這工作。
PHIL|1|7|我為你們眾人有這樣的想法原是應當的，因為你們常在我心裏；無論我是在捆鎖中，在辯明並證實福音的時候，你們都與我一同蒙恩。
PHIL|1|8|我以基督耶穌的心腸切切想念你們眾人，這是上帝可以為我作證的。
PHIL|1|9|我所禱告的就是：要你們的愛心，在知識和各樣見識上，不斷增長，
PHIL|1|10|使你們能分辨是非，在基督的日子作真誠無可指責的人，
PHIL|1|11|更靠著耶穌基督結滿仁義的果子，歸榮耀稱讚給上帝。
PHIL|1|12|弟兄們，我要你們知道，我所遭遇的事反而使福音更興旺，
PHIL|1|13|以致御營全軍和其餘的人都知道我是為基督的緣故受捆鎖的；
PHIL|1|14|而且那在主裏的弟兄，多半都因我受的捆鎖而篤信不疑，越發放膽無所懼怕地傳道。
PHIL|1|15|有些人傳基督是出於嫉妒紛爭；有些人是出於好意。
PHIL|1|16|後者是出於愛心，知道我奉差遣是為福音辯護的。
PHIL|1|17|前者傳基督是出於自私，動機不純，企圖要加增我捆鎖的苦楚。
PHIL|1|18|這又何妨呢？或是假意或是真心，無論如何，只要基督被傳開了，為此我就歡喜。 我還要歡喜，
PHIL|1|19|因為我知道，這事藉著你們的祈禱和耶穌基督的靈的幫助，終必使我得到釋放。
PHIL|1|20|這就是我所切慕、所盼望的：沒有一事能使我羞愧；反倒凡事坦然無懼，無論是生是死，總要讓基督在我身上照常顯大。
PHIL|1|21|因為我活著就是基督，死了就有益處。
PHIL|1|22|但是，我在肉身活著，若能有工作的成果，我就不知道該挑選甚麼。
PHIL|1|23|我處在兩難之間：我情願離世與基督同在，因為這是好得無比的；
PHIL|1|24|然而，我為你們肉身活著更加要緊。
PHIL|1|25|既然我這樣深信，就知道仍要留在世間，且與你們眾人一起存留，使你們在所信的道上又長進又喜樂，
PHIL|1|26|為了我再到你們那裏時，你們在基督耶穌裏的誇耀越發加增。
PHIL|1|27|最重要的是：你們行事為人要與基督的福音相稱，這樣，無論我來見你們，或不在你們那裏，都可以聽到你們的景況，知道你們同有一個心志，站立得穩，為福音的信仰齊心努力，
PHIL|1|28|絲毫不怕敵人的威脅；以此證明他們會沉淪，你們會得救，這是出於上帝。
PHIL|1|29|因為你們蒙恩，不但得以信服基督，而且要為他受苦。
PHIL|1|30|你們的爭戰，就與你們曾在我身上見過、現在所聽到的是一樣的。
PHIL|2|1|所以，在基督裏若有任何勸勉，若有任何愛心的安慰，若有任何聖靈的團契，若有任何慈悲憐憫，
PHIL|2|2|你們就要意志相同，愛心相同，有一致的心思，一致的想法，使我的喜樂得以滿足。
PHIL|2|3|凡事不可自私自利，不可貪圖虛榮；只要心存謙卑，各人看別人比自己強。
PHIL|2|4|各人不要單顧自己的事，也要顧別人的事。
PHIL|2|5|你們當以基督耶穌的心為心：
PHIL|2|6|他本有上帝的形像， 卻不堅持自己與上帝同等 ；
PHIL|2|7|反倒虛己， 取了奴僕的形像， 成為人的樣式； 既有人的樣子，
PHIL|2|8|就謙卑自己， 存心順服，以至於死， 且死在十字架上。
PHIL|2|9|所以上帝把他升為至高， 又賜給他超乎萬名之上的名，
PHIL|2|10|使一切在天上的、地上的和地底下的， 因耶穌的名， 眾膝都要跪下，
PHIL|2|11|眾口都要宣認： 耶穌基督是主， 歸榮耀給父上帝。
PHIL|2|12|我親愛的，這樣看來，你們向來是順服的，不但我在你們那裏，就是我現在不在你們那裏的時候更是順服的，就當恐懼戰兢完成你們自己得救的事；
PHIL|2|13|因為是上帝在你們心裏運行，使你們又立志又實行，為要成就他的美意。
PHIL|2|14|你們無論做甚麼事，都不要發怨言起爭論，
PHIL|2|15|好使你們無可指責，誠實無偽，在這彎曲悖謬的世代作上帝無瑕疵的兒女。你們在這世代中要像明光照耀，
PHIL|2|16|將生命的道顯明出來，使我在基督的日子得以誇耀我沒有白跑，也沒有徒勞。
PHIL|2|17|我以你們的信心為供獻的祭物，我若被澆獻在其上也是喜樂，並且與你們眾人一同喜樂。
PHIL|2|18|你們也要照樣喜樂，並且與我一同喜樂。
PHIL|2|19|我靠主耶穌希望很快能差 提摩太 去見你們，好讓我知道你們的事而心裏得著安慰。
PHIL|2|20|因為我沒有別人與我同心，真正關懷你們的事。
PHIL|2|21|其他的人都求自己的事，並不求耶穌基督的事。
PHIL|2|22|但你們知道 提摩太 是經得起考驗的，他與我為了福音一同服侍，待我像兒子待父親一樣。
PHIL|2|23|所以，我一看出我的事怎樣了結，我希望立刻差他去，
PHIL|2|24|但我靠著主自信我不久也會去。
PHIL|2|25|然而，我想必須差 以巴弗提 到你們那裏去。他是我的弟兄、同工和戰友，是你們差遣來供應我需要的。
PHIL|2|26|他很想念 你們眾人，並且極其難過，因為你們聽見他病了。
PHIL|2|27|他真的生病了，幾乎要死。然而上帝憐憫他，不但憐憫他，也憐憫我，免得我憂上加憂。
PHIL|2|28|所以，我更要盡快送他回去，好讓你們再見到他而喜樂，我也可以減少憂愁。
PHIL|2|29|故此，你們要在主裏歡歡喜喜地接待他，而且要尊重這樣的人，
PHIL|2|30|因他為做基督的工作不顧性命，幾乎至死，為要補足你們供應我不夠的地方。
PHIL|3|1|末了，我的弟兄們，你們要靠主喜樂。我把這些話再寫給你們，對我並不困難，對你們卻是妥當的。
PHIL|3|2|應當防備犬類，防備作惡的，防備妄自行割的。
PHIL|3|3|因為真受割禮的，就是我們這藉著上帝的靈敬拜、以基督耶穌為誇耀、不依靠肉體的。
PHIL|3|4|其實，我也可以靠肉體；若是別人以為他可以依靠肉體，我更可以。
PHIL|3|5|我出生後第八天受割禮；我是 以色列 族、 便雅憫 支派的人，是 希伯來 人所生的 希伯來 人。就律法說，我是法利賽人；
PHIL|3|6|就熱心說，我是迫害教會的；就律法上的義說，我是無可指責的。
PHIL|3|7|只是我先前以為對我是有益的，我現在因基督的緣故而當作是有損的。
PHIL|3|8|不但如此，我已把萬事當作是有損的，因我以認識我主基督耶穌為至寶。我為他已經丟棄萬事，看作糞土，為要贏得基督，
PHIL|3|9|並且得以在他裏面，不是有自己因律法而得的義，而是有信基督的義 ，就是基於信，從上帝而來的義，
PHIL|3|10|使我認識基督，知道他復活的大能，並且知道和他一同受苦，效法他的死，
PHIL|3|11|或許我也得以從死人中復活。
PHIL|3|12|這不是說我已經得著了，已經完全了；而是竭力追求，或許可以得著基督耶穌 所要我得著的 。
PHIL|3|13|弟兄們，我不是以為自己已經得著了；我只有一件事，就是忘記背後，努力面前的，
PHIL|3|14|向著標竿直跑，要得上帝在基督耶穌裏從上面召我來得的獎賞。
PHIL|3|15|所以，我們中間凡是成熟的人，總要存這樣的心；若在甚麼事上存別樣的心，上帝也會把這些事指示你們。
PHIL|3|16|然而，我們達到甚麼地步，就當照這個地步行。
PHIL|3|17|弟兄們，你們要一同效法我，也當留意看那些效法我們榜樣的人。
PHIL|3|18|因為，我屢次告訴你們，現在又流淚告訴你們：許多人行事是基督十字架的仇敵。
PHIL|3|19|他們的結局就是滅亡。他們的神明是自己的肚腹；他們以自己的羞辱為光榮，專以地上的事為念。
PHIL|3|20|我們卻是天上的國民，並且等候救主，就是主耶穌基督從天上降臨。
PHIL|3|21|他要按著那能使萬有歸服自己的大能，把我們這卑賤的身體改變形狀，和他自己榮耀的身體相似。
PHIL|4|1|我所親愛、所想念的弟兄們，你們就是我的喜樂，我的冠冕。我親愛的，你們應當靠主站立得穩。
PHIL|4|2|我勸 友阿蝶 和 循都基 要在主裏同心。
PHIL|4|3|我也求你這真實同負一軛的，要幫助這兩個女人，因為她們在福音上曾與我、 革利免 和我其餘的同工一同勞苦，他們的名字都在生命冊上。
PHIL|4|4|你們要靠主常常喜樂。我再說，你們要喜樂。
PHIL|4|5|要讓眾人知道你們謙讓的心。主已經近了。
PHIL|4|6|應當一無掛慮，只要凡事藉著禱告、祈求和感謝，將你們所要的告訴上帝。
PHIL|4|7|上帝所賜那超越人所能了解的平安 ，必在基督耶穌裏，保守你們的心懷意念。
PHIL|4|8|末了，弟兄們，凡是真實的、凡是可敬的、凡是公義的、凡是清潔的、凡是可愛的、凡是有美名的，若有甚麼德行，若有甚麼稱讚，你們都要留意。
PHIL|4|9|你們從我所學習的，所領受的，所聽見的，所看見的事，你們都要繼續去做，賜平安的上帝就必與你們同在。
PHIL|4|10|我靠主大大喜樂，因為你們關懷我的心如今又表現了出來；其實你們一直都關懷我，只是沒有機會罷了。
PHIL|4|11|我並不是因缺乏而說這話，因為我已經學會無論在甚麼景況都可以知足。
PHIL|4|12|我知道怎樣處卑賤，也知道怎樣處豐富；或飽足或飢餓，或有餘或缺乏，任何事情，任何景況，我都得了祕訣。
PHIL|4|13|我靠著那加給我力量的，凡事都能做。
PHIL|4|14|然而，你們能和我分擔憂患是一件好事。
PHIL|4|15|腓立比 人哪，你們也知道我開始傳福音、離開 馬其頓 的時候，在收支的事上，除了你們以外，並沒有別的教會和我分擔。
PHIL|4|16|就是我在 帖撒羅尼迦 ，你們也一再差人來供給我的需用。
PHIL|4|17|我並不求甚麼饋贈，只求你們的果子不斷增多，歸在你們的賬上。
PHIL|4|18|但我已經如數收到，並且有餘；我已經充足，因我從 以巴弗提 受了你們的饋贈，當作極美的香氣，為上帝所接納、所喜悅的祭物。
PHIL|4|19|我的上帝必照他榮耀的豐富，在基督耶穌裏，使你們一切所需用的都充足。
PHIL|4|20|願榮耀歸給我們的父上帝，直到永永遠遠。阿們！
PHIL|4|21|請問候在基督耶穌裏的各位聖徒。跟我一起的眾弟兄都問候你們。
PHIL|4|22|眾聖徒都問候你們，特別在凱撒家裏的人問候你們。
PHIL|4|23|願主耶穌基督的恩與你們的靈同在！
