SONG|1|1|osculetur me osculo oris sui quia meliora sunt ubera tua vino
SONG|1|2|fraglantia unguentis optimis oleum effusum nomen tuum ideo adulescentulae dilexerunt te
SONG|1|3|trahe me post te curremus introduxit me rex in cellaria sua exultabimus et laetabimur in te memores uberum tuorum super vinum recti diligunt te
SONG|1|4|nigra sum sed formonsa filiae Hierusalem sicut tabernacula Cedar sicut pelles Salomonis
SONG|1|5|nolite me considerare quod fusca sim quia decoloravit me sol filii matris meae pugnaverunt contra me posuerunt me custodem in vineis vineam meam non custodivi
SONG|1|6|indica mihi quem diligit anima mea ubi pascas ubi cubes in meridie ne vagari incipiam per greges sodalium tuorum
SONG|1|7|si ignoras te o pulchra inter mulieres egredere et abi post vestigia gregum et pasce hedos tuos iuxta tabernacula pastorum
SONG|1|8|equitatui meo in curribus Pharaonis adsimilavi te amica mea
SONG|1|9|pulchrae sunt genae tuae sicut turturis collum tuum sicut monilia
SONG|1|10|murenulas aureas faciemus tibi vermiculatas argento
SONG|1|11|dum esset rex in accubitu suo nardus mea dedit odorem suum
SONG|1|12|fasciculus murrae dilectus meus mihi inter ubera mea commorabitur
SONG|1|13|botrus cypri dilectus meus mihi in vineis Engaddi
SONG|1|14|ecce tu pulchra es amica mea ecce tu pulchra oculi tui columbarum
SONG|1|15|ecce tu pulcher es dilecte mi et decorus lectulus noster floridus
SONG|1|16|tigna domorum nostrarum cedrina laquearia nostra cypressina
SONG|2|1|ego flos campi et lilium convallium
SONG|2|2|sicut lilium inter spinas sic amica mea inter filias
SONG|2|3|sicut malum inter ligna silvarum sic dilectus meus inter filios sub umbra illius quam desideraveram sedi et fructus eius dulcis gutturi meo
SONG|2|4|introduxit me in cellam vinariam ordinavit in me caritatem
SONG|2|5|fulcite me floribus stipate me malis quia amore langueo
SONG|2|6|leva eius sub capite meo et dextera illius amplexabitur me
SONG|2|7|adiuro vos filiae Hierusalem per capreas cervosque camporum ne suscitetis neque evigilare faciatis dilectam quoadusque ipsa velit
SONG|2|8|vox dilecti mei ecce iste venit saliens in montibus transiliens colles
SONG|2|9|similis est dilectus meus capreae hinuloque cervorum en ipse stat post parietem nostrum despiciens per fenestras prospiciens per cancellos
SONG|2|10|et dilectus meus loquitur mihi surge propera amica mea formonsa mea et veni
SONG|2|11|iam enim hiemps transiit imber abiit et recessit
SONG|2|12|flores apparuerunt in terra tempus putationis advenit vox turturis audita est in terra nostra
SONG|2|13|ficus protulit grossos suos vineae florent dederunt odorem surge amica mea speciosa mea et veni
SONG|2|14|columba mea in foraminibus petrae in caverna maceriae ostende mihi faciem tuam sonet vox tua in auribus meis vox enim tua dulcis et facies tua decora
SONG|2|15|capite nobis vulpes vulpes parvulas quae demoliuntur vineas nam vinea nostra floruit
SONG|2|16|dilectus meus mihi et ego illi qui pascitur inter lilia
SONG|2|17|donec adspiret dies et inclinentur umbrae revertere similis esto dilecte mi capreae aut hinulo cervorum super montes Bether
SONG|3|1|in lectulo meo per noctes quaesivi quem diligit anima mea quaesivi illum et non inveni
SONG|3|2|surgam et circuibo civitatem per vicos et plateas quaeram quem diligit anima mea quaesivi illum et non inveni
SONG|3|3|invenerunt me vigiles qui custodiunt civitatem num quem dilexit anima mea vidistis
SONG|3|4|paululum cum pertransissem eos inveni quem diligit anima mea tenui eum nec dimittam donec introducam illum in domum matris meae et in cubiculum genetricis meae
SONG|3|5|adiuro vos filiae Hierusalem per capreas cervosque camporum ne suscitetis neque evigilare faciatis dilectam donec ipsa velit
SONG|3|6|quae est ista quae ascendit per desertum sicut virgula fumi ex aromatibus murrae et turis et universi pulveris pigmentarii
SONG|3|7|en lectulum Salomonis sexaginta fortes ambiunt ex fortissimis Israhel
SONG|3|8|omnes tenentes gladios et ad bella doctissimi uniuscuiusque ensis super femur suum propter timores nocturnos
SONG|3|9|ferculum fecit sibi rex Salomon de lignis Libani
SONG|3|10|columnas eius fecit argenteas reclinatorium aureum ascensum purpureum media caritate constravit propter filias Hierusalem
SONG|3|11|egredimini et videte filiae Sion regem Salomonem in diademate quo coronavit eum mater sua in die disponsionis illius et in die laetitiae cordis eius
SONG|4|1|quam pulchra es amica mea quam pulchra es oculi tui columbarum absque eo quod intrinsecus latet capilli tui sicut greges caprarum quae ascenderunt de monte Galaad
SONG|4|2|dentes tui sicut greges tonsarum quae ascenderunt de lavacro omnes gemellis fetibus et sterilis non est inter eas
SONG|4|3|sicut vitta coccinea labia tua et eloquium tuum dulce sicut fragmen mali punici ita genae tuae absque eo quod intrinsecus latet
SONG|4|4|sicut turris David collum tuum quae aedificata est cum propugnaculis mille clypei pendent ex ea omnis armatura fortium
SONG|4|5|duo ubera tua sicut duo hinuli capreae gemelli qui pascuntur in liliis
SONG|4|6|donec adspiret dies et inclinentur umbrae vadam ad montem murrae et ad collem turis
SONG|4|7|tota pulchra es amica mea et macula non est in te
SONG|4|8|veni de Libano sponsa veni de Libano veni coronaberis de capite Amana de vertice Sanir et Hermon de cubilibus leonum de montibus pardorum
SONG|4|9|vulnerasti cor meum soror mea sponsa vulnerasti cor meum in uno oculorum tuorum et in uno crine colli tui
SONG|4|10|quam pulchrae sunt mammae tuae soror mea sponsa pulchriora ubera tua vino et odor unguentorum tuorum super omnia aromata
SONG|4|11|favus distillans labia tua sponsa mel et lac sub lingua tua et odor vestimentorum tuorum sicut odor turis
SONG|4|12|hortus conclusus soror mea sponsa hortus conclusus fons signatus
SONG|4|13|emissiones tuae paradisus malorum punicorum cum pomorum fructibus cypri cum nardo
SONG|4|14|nardus et crocus fistula et cinnamomum cum universis lignis Libani murra et aloe cum omnibus primis unguentis
SONG|4|15|fons hortorum puteus aquarum viventium quae fluunt impetu de Libano
SONG|4|16|surge aquilo et veni auster perfla hortum meum et fluant aromata illius
SONG|5|1|veniat dilectus meus in hortum suum et comedat fructum pomorum suorum veni in hortum meum soror mea sponsa messui murram meam cum aromatibus meis comedi favum cum melle meo bibi vinum meum cum lacte meo comedite amici bibite et inebriamini carissimi
SONG|5|2|ego dormio et cor meum vigilat vox dilecti mei pulsantis aperi mihi soror mea amica mea columba mea inmaculata mea quia caput meum plenum est rore et cincinni mei guttis noctium
SONG|5|3|expoliavi me tunica mea quomodo induar illa lavi pedes meos quomodo inquinabo illos
SONG|5|4|dilectus meus misit manum suam per foramen et venter meus intremuit ad tactum eius
SONG|5|5|surrexi ut aperirem dilecto meo manus meae stillaverunt murra digiti mei pleni murra probatissima
SONG|5|6|pessulum ostii aperui dilecto meo at ille declinaverat atque transierat anima mea liquefacta est ut locutus est quaesivi et non inveni illum vocavi et non respondit mihi
SONG|5|7|invenerunt me custodes qui circumeunt civitatem percusserunt me vulneraverunt me tulerunt pallium meum mihi custodes murorum
SONG|5|8|adiuro vos filiae Hierusalem si inveneritis dilectum meum ut nuntietis ei quia amore langueo
SONG|5|9|qualis est dilectus tuus ex dilecto o pulcherrima mulierum qualis est dilectus tuus ex dilecto quia sic adiurasti nos
SONG|5|10|dilectus meus candidus et rubicundus electus ex milibus
SONG|5|11|caput eius aurum optimum comae eius sicut elatae palmarum nigrae quasi corvus
SONG|5|12|oculi eius sicut columbae super rivulos aquarum quae lacte sunt lotae et resident iuxta fluenta plenissima
SONG|5|13|genae illius sicut areolae aromatum consitae a pigmentariis labia eius lilia distillantia murram primam
SONG|5|14|manus illius tornatiles aureae plenae hyacinthis venter eius eburneus distinctus sapphyris
SONG|5|15|crura illius columnae marmoreae quae fundatae sunt super bases aureas species eius ut Libani electus ut cedri
SONG|5|16|guttur illius suavissimum et totus desiderabilis talis est dilectus meus et iste est amicus meus filiae Hierusalem
SONG|5|17|quo abiit dilectus tuus o pulcherrima mulierum quo declinavit dilectus tuus et quaeremus eum tecum
SONG|6|1|dilectus meus descendit in hortum suum ad areolam aromatis ut pascatur in hortis et lilia colligat
SONG|6|2|ego dilecto meo et dilectus meus mihi qui pascitur inter lilia
SONG|6|3|pulchra es amica mea suavis et decora sicut Hierusalem terribilis ut castrorum acies ordinata
SONG|6|4|averte oculos tuos a me quia ipsi me avolare fecerunt capilli tui sicut grex caprarum quae apparuerunt de Galaad
SONG|6|5|dentes tui sicut grex ovium quae ascenderunt de lavacro omnes gemellis fetibus et sterilis non est in eis
SONG|6|6|sicut cortex mali punici genae tuae absque occultis tuis
SONG|6|7|sexaginta sunt reginae et octoginta concubinae et adulescentularum non est numerus
SONG|6|8|una est columba mea perfecta mea una est matris suae electa genetrici suae viderunt illam filiae et beatissimam praedicaverunt reginae et concubinae et laudaverunt eam
SONG|6|9|quae est ista quae progreditur quasi aurora consurgens pulchra ut luna electa ut sol terribilis ut acies ordinata
SONG|6|10|descendi ad hortum nucum ut viderem poma convallis ut inspicerem si floruisset vinea et germinassent mala punica
SONG|6|11|nescivi anima mea conturbavit me propter quadrigas Aminadab
SONG|6|12|revertere revertere Sulamitis revertere revertere ut intueamur te
SONG|7|1|quid videbis in Sulamiten nisi choros castrorum quam pulchri sunt gressus tui in calciamentis filia principis iunctura feminum tuorum sicut monilia quae fabricata sunt manu artificis
SONG|7|2|umbilicus tuus crater tornatilis numquam indigens poculis venter tuus sicut acervus tritici vallatus liliis
SONG|7|3|duo ubera tua sicut duo hinuli gemelli capreae
SONG|7|4|collum tuum sicut turris eburnea oculi tui sicut piscinae in Esebon quae sunt in porta filiae multitudinis nasus tuus sicut turris Libani quae respicit contra Damascum
SONG|7|5|caput tuum ut Carmelus et comae capitis tui sicut purpura regis vincta canalibus
SONG|7|6|quam pulchra es et quam decora carissima in deliciis
SONG|7|7|statura tua adsimilata est palmae et ubera tua botris
SONG|7|8|dixi ascendam in palmam adprehendam fructus eius et erunt ubera tua sicut botri vineae et odor oris tui sicut malorum
SONG|7|9|guttur tuum sicut vinum optimum dignum dilecto meo ad potandum labiisque et dentibus illius ruminandum
SONG|7|10|ego dilecto meo et ad me conversio eius
SONG|7|11|veni dilecte mi egrediamur in agrum commoremur in villis
SONG|7|12|mane surgamus ad vineas videamus si floruit vinea si flores fructus parturiunt si floruerunt mala punica ibi dabo tibi ubera mea
SONG|7|13|mandragorae dederunt odorem in portis nostris omnia poma nova et vetera dilecte mi servavi tibi
SONG|8|1|quis mihi det te fratrem meum sugentem ubera matris meae ut inveniam te foris et deosculer et iam me nemo despiciat
SONG|8|2|adprehendam te et ducam in domum matris meae ibi me docebis et dabo tibi poculum ex vino condito et mustum malorum granatorum meorum
SONG|8|3|leva eius sub capite meo et dextera illius amplexabitur me
SONG|8|4|adiuro vos filiae Hierusalem ne suscitetis et evigilare faciatis dilectam donec ipsa velit
SONG|8|5|quae est ista quae ascendit de deserto deliciis affluens et nixa super dilectum suum sub arbore malo suscitavi te ibi corrupta est mater tua ibi violata est genetrix tua
SONG|8|6|pone me ut signaculum super cor tuum ut signaculum super brachium tuum quia fortis est ut mors dilectio dura sicut inferus aemulatio lampades eius lampades ignis atque flammarum
SONG|8|7|aquae multae non poterunt extinguere caritatem nec flumina obruent illam si dederit homo omnem substantiam domus suae pro dilectione quasi nihil despicient eum
SONG|8|8|soror nostra parva et ubera non habet quid faciemus sorori nostrae in die quando adloquenda est
SONG|8|9|si murus est aedificemus super eum propugnacula argentea si ostium est conpingamus illud tabulis cedrinis
SONG|8|10|ego murus et ubera mea sicut turris ex quo facta sum coram eo quasi pacem repperiens
SONG|8|11|vinea fuit Pacifico in ea quae habet populos tradidit eam custodibus vir adfert pro fructu eius mille argenteos
SONG|8|12|vinea mea coram me est mille tui Pacifice et ducenti his qui custodiunt fructus eius
SONG|8|13|quae habitas in hortis amici auscultant fac me audire vocem tuam
SONG|8|14|fuge dilecte mi et adsimilare capreae hinuloque cervorum super montes aromatum
