REV|1|1|The revelation of Jesus Christ, which God gave him to show his servants what must soon take place. He made it known by sending his angel to his servant John,
REV|1|2|who testifies to everything he saw--that is, the word of God and the testimony of Jesus Christ.
REV|1|3|Blessed is the one who reads the words of this prophecy, and blessed are those who hear it and take to heart what is written in it, because the time is near.
REV|1|4|John, To the seven churches in the province of Asia: Grace and peace to you from him who is, and who was, and who is to come, and from the seven spirits
REV|1|5|before his throne, and from Jesus Christ, who is the faithful witness, the firstborn from the dead, and the ruler of the kings of the earth.
REV|1|6|To him who loves us and has freed us from our sins by his blood, and has made us to be a kingdom and priests to serve his God and Father--to him be glory and power for ever and ever! Amen.
REV|1|7|Look, he is coming with the clouds, and every eye will see him, even those who pierced him; and all the peoples of the earth will mourn because of him. So shall it be! Amen.
REV|1|8|"I am the Alpha and the Omega," says the Lord God, "who is, and who was, and who is to come, the Almighty."
REV|1|9|I, John, your brother and companion in the suffering and kingdom and patient endurance that are ours in Jesus, was on the island of Patmos because of the word of God and the testimony of Jesus.
REV|1|10|On the Lord's Day I was in the Spirit, and I heard behind me a loud voice like a trumpet,
REV|1|11|which said: "Write on a scroll what you see and send it to the seven churches: to Ephesus, Smyrna, Pergamum, Thyatira, Sardis, Philadelphia and Laodicea."
REV|1|12|I turned around to see the voice that was speaking to me. And when I turned I saw seven golden lampstands,
REV|1|13|and among the lampstands was someone "like a son of man," dressed in a robe reaching down to his feet and with a golden sash around his chest.
REV|1|14|His head and hair were white like wool, as white as snow, and his eyes were like blazing fire.
REV|1|15|His feet were like bronze glowing in a furnace, and his voice was like the sound of rushing waters.
REV|1|16|In his right hand he held seven stars, and out of his mouth came a sharp double-edged sword. His face was like the sun shining in all its brilliance.
REV|1|17|When I saw him, I fell at his feet as though dead. Then he placed his right hand on me and said: "Do not be afraid. I am the First and the Last.
REV|1|18|I am the Living One; I was dead, and behold I am alive for ever and ever! And I hold the keys of death and Hades.
REV|1|19|"Write, therefore, what you have seen, what is now and what will take place later.
REV|1|20|The mystery of the seven stars that you saw in my right hand and of the seven golden lampstands is this: The seven stars are the angels of the seven churches, and the seven lampstands are the seven churches.
REV|2|1|"To the angel of the church in Ephesus write: These are the words of him who holds the seven stars in his right hand and walks among the seven golden lampstands:
REV|2|2|I know your deeds, your hard work and your perseverance. I know that you cannot tolerate wicked men, that you have tested those who claim to be apostles but are not, and have found them false.
REV|2|3|You have persevered and have endured hardships for my name, and have not grown weary.
REV|2|4|Yet I hold this against you: You have forsaken your first love.
REV|2|5|Remember the height from which you have fallen! Repent and do the things you did at first. If you do not repent, I will come to you and remove your lampstand from its place.
REV|2|6|But you have this in your favor: You hate the practices of the Nicolaitans, which I also hate.
REV|2|7|He who has an ear, let him hear what the Spirit says to the churches. To him who overcomes, I will give the right to eat from the tree of life, which is in the paradise of God.
REV|2|8|"To the angel of the church in Smyrna write: These are the words of him who is the First and the Last, who died and came to life again.
REV|2|9|I know your afflictions and your poverty-yet you are rich! I know the slander of those who say they are Jews and are not, but are a synagogue of Satan.
REV|2|10|Do not be afraid of what you are about to suffer. I tell you, the devil will put some of you in prison to test you, and you will suffer persecution for ten days. Be faithful, even to the point of death, and I will give you the crown of life.
REV|2|11|He who has an ear, let him hear what the Spirit says to the churches. He who overcomes will not be hurt at all by the second death.
REV|2|12|"To the angel of the church in Pergamum write: These are the words of him who has the sharp, doubleedged sword.
REV|2|13|I know where you live-where Satan has his throne. Yet you remain true to my name. You did not renounce your faith in me, even in the days of Antipas, my faithful witness, who was put to death in your city-where Satan lives.
REV|2|14|Nevertheless, I have a few things against you: You have people there who hold to the teaching of Balaam, who taught Balak to entice the Israelites to sin by eating food sacrificed to idols and by committing sexual immorality.
REV|2|15|Likewise you also have those who hold to the teaching of the Nicolaitans.
REV|2|16|Repent therefore! Otherwise, I will soon come to you and will fight against them with the sword of my mouth.
REV|2|17|He who has an ear, let him hear what the Spirit says to the churches. To him who overcomes, I will give some of the hidden manna. I will also give him a white stone with a new name written on it, known only to him who receives it.
REV|2|18|"To the angel of the church in Thyatira write: These are the words of the Son of God, whose eyes are like blazing fire and whose feet are like burnished bronze.
REV|2|19|I know your deeds, your love and faith, your service and perseverance, and that you are now doing more than you did at first.
REV|2|20|Nevertheless, I have this against you: You tolerate that woman Jezebel, who calls herself a prophetess. By her teaching she misleads my servants into sexual immorality and the eating of food sacrificed to idols.
REV|2|21|I have given her time to repent of her immorality, but she is unwilling.
REV|2|22|So I will cast her on a bed of suffering, and I will make those who commit adultery with her suffer intensely, unless they repent of her ways.
REV|2|23|I will strike her children dead. Then all the churches will know that I am he who searches hearts and minds, and I will repay each of you according to your deeds.
REV|2|24|Now I say to the rest of you in Thyatira, to you who do not hold to her teaching and have not learned Satan's so-called deep secrets (I will not impose any other burden on you):
REV|2|25|Only hold on to what you have until I come.
REV|2|26|To him who overcomes and does my will to the end, I will give authority over the nations--
REV|2|27|'He will rule them with an iron scepter; he will dash them to pieces like pottery'--
REV|2|28|just as I have received authority from my Father. I will also give him the morning star.
REV|2|29|He who has an ear, let him hear what the Spirit says to the churches.
REV|3|1|"To the angel of the church in Sardis write: These are the words of him who holds the seven spirits of God and the seven stars. I know your deeds; you have a reputation of being alive, but you are dead.
REV|3|2|Wake up! Strengthen what remains and is about to die, for I have not found your deeds complete in the sight of my God.
REV|3|3|Remember, therefore, what you have received and heard; obey it, and repent. But if you do not wake up, I will come like a thief, and you will not know at what time I will come to you.
REV|3|4|Yet you have a few people in Sardis who have not soiled their clothes. They will walk with me, dressed in white, for they are worthy.
REV|3|5|He who overcomes will, like them, be dressed in white. I will never blot out his name from the book of life, but will acknowledge his name before my Father and his angels.
REV|3|6|He who has an ear, let him hear what the Spirit says to the churches.
REV|3|7|"To the angel of the church in Philadelphia write: These are the words of him who is holy and true, who holds the key of David. What he opens no one can shut, and what he shuts no one can open.
REV|3|8|I know your deeds. See, I have placed before you an open door that no one can shut. I know that you have little strength, yet you have kept my word and have not denied my name.
REV|3|9|I will make those who are of the synagogue of Satan, who claim to be Jews though they are not, but are liars--I will make them come and fall down at your feet and acknowledge that I have loved you.
REV|3|10|Since you have kept my command to endure patiently, I will also keep you from the hour of trial that is going to come upon the whole world to test those who live on the earth.
REV|3|11|I am coming soon. Hold on to what you have, so that no one will take your crown.
REV|3|12|Him who overcomes I will make a pillar in the temple of my God. Never again will he leave it. I will write on him the name of my God and the name of the city of my God, the new Jerusalem, which is coming down out of heaven from my God; and I will also write on him my new name.
REV|3|13|He who has an ear, let him hear what the Spirit says to the churches.
REV|3|14|"To the angel of the church in Laodicea write: These are the words of the Amen, the faithful and true witness, the ruler of God's creation.
REV|3|15|I know your deeds, that you are neither cold nor hot. I wish you were either one or the other!
REV|3|16|So, because you are lukewarm--neither hot nor cold--I am about to spit you out of my mouth.
REV|3|17|You say, 'I am rich; I have acquired wealth and do not need a thing.' But you do not realize that you are wretched, pitiful, poor, blind and naked.
REV|3|18|I counsel you to buy from me gold refined in the fire, so you can become rich; and white clothes to wear, so you can cover your shameful nakedness; and salve to put on your eyes, so you can see.
REV|3|19|Those whom I love I rebuke and discipline. So be earnest, and repent.
REV|3|20|Here I am! I stand at the door and knock. If anyone hears my voice and opens the door, I will come in and eat with him, and he with me.
REV|3|21|To him who overcomes, I will give the right to sit with me on my throne, just as I overcame and sat down with my Father on his throne.
REV|3|22|He who has an ear, let him hear what the Spirit says to the churches."
REV|4|1|After this I looked, and there before me was a door standing open in heaven. And the voice I had first heard speaking to me like a trumpet said, "Come up here, and I will show you what must take place after this."
REV|4|2|At once I was in the Spirit, and there before me was a throne in heaven with someone sitting on it.
REV|4|3|And the one who sat there had the appearance of jasper and carnelian. A rainbow, resembling an emerald, encircled the throne.
REV|4|4|Surrounding the throne were twenty-four other thrones, and seated on them were twenty-four elders. They were dressed in white and had crowns of gold on their heads.
REV|4|5|From the throne came flashes of lightning, rumblings and peals of thunder. Before the throne, seven lamps were blazing. These are the seven spirits of God.
REV|4|6|Also before the throne there was what looked like a sea of glass, clear as crystal.
REV|4|7|In the center, around the throne, were four living creatures, and they were covered with eyes, in front and in back. The first living creature was like a lion, the second was like an ox, the third had a face like a man, the fourth was like a flying eagle.
REV|4|8|Each of the four living creatures had six wings and was covered with eyes all around, even under his wings. Day and night they never stop saying: "Holy, holy, holy is the Lord God Almighty, who was, and is, and is to come."
REV|4|9|Whenever the living creatures give glory, honor and thanks to him who sits on the throne and who lives for ever and ever,
REV|4|10|the twenty-four elders fall down before him who sits on the throne, and worship him who lives for ever and ever. They lay their crowns before the throne and say:
REV|4|11|"You are worthy, our Lord and God, to receive glory and honor and power, for you created all things, and by your will they were created and have their being."
REV|5|1|Then I saw in the right hand of him who sat on the throne a scroll with writing on both sides and sealed with seven seals.
REV|5|2|And I saw a mighty angel proclaiming in a loud voice, "Who is worthy to break the seals and open the scroll?"
REV|5|3|But no one in heaven or on earth or under the earth could open the scroll or even look inside it.
REV|5|4|I wept and wept because no one was found who was worthy to open the scroll or look inside.
REV|5|5|Then one of the elders said to me, "Do not weep! See, the Lion of the tribe of Judah, the Root of David, has triumphed. He is able to open the scroll and its seven seals."
REV|5|6|Then I saw a Lamb, looking as if it had been slain, standing in the center of the throne, encircled by the four living creatures and the elders. He had seven horns and seven eyes, which are the seven spirits of God sent out into all the earth.
REV|5|7|He came and took the scroll from the right hand of him who sat on the throne.
REV|5|8|And when he had taken it, the four living creatures and the twenty-four elders fell down before the Lamb. Each one had a harp and they were holding golden bowls full of incense, which are the prayers of the saints.
REV|5|9|And they sang a new song: "You are worthy to take the scroll and to open its seals, because you were slain, and with your blood you purchased men for God from every tribe and language and people and nation.
REV|5|10|You have made them to be a kingdom and priests to serve our God, and they will reign on the earth."
REV|5|11|Then I looked and heard the voice of many angels, numbering thousands upon thousands, and ten thousand times ten thousand. They encircled the throne and the living creatures and the elders.
REV|5|12|In a loud voice they sang: "Worthy is the Lamb, who was slain, to receive power and wealth and wisdom and strength and honor and glory and praise!"
REV|5|13|Then I heard every creature in heaven and on earth and under the earth and on the sea, and all that is in them, singing: "To him who sits on the throne and to the Lamb be praise and honor and glory and power, for ever and ever!"
REV|5|14|The four living creatures said, "Amen," and the elders fell down and worshiped.
REV|6|1|I watched as the Lamb opened the first of the seven seals. Then I heard one of the four living creatures say in a voice like thunder, "Come!"
REV|6|2|I looked, and there before me was a white horse! Its rider held a bow, and he was given a crown, and he rode out as a conqueror bent on conquest.
REV|6|3|When the Lamb opened the second seal, I heard the second living creature say, "Come!"
REV|6|4|Then another horse came out, a fiery red one. Its rider was given power to take peace from the earth and to make men slay each other. To him was given a large sword.
REV|6|5|When the Lamb opened the third seal, I heard the third living creature say, "Come!" I looked, and there before me was a black horse! Its rider was holding a pair of scales in his hand.
REV|6|6|Then I heard what sounded like a voice among the four living creatures, saying, "A quart of wheat for a day's wages, and three quarts of barley for a day's wages, and do not damage the oil and the wine!"
REV|6|7|When the Lamb opened the fourth seal, I heard the voice of the fourth living creature say, "Come!"
REV|6|8|I looked, and there before me was a pale horse! Its rider was named Death, and Hades was following close behind him. They were given power over a fourth of the earth to kill by sword, famine and plague, and by the wild beasts of the earth.
REV|6|9|When he opened the fifth seal, I saw under the altar the souls of those who had been slain because of the word of God and the testimony they had maintained.
REV|6|10|They called out in a loud voice, "How long, Sovereign Lord, holy and true, until you judge the inhabitants of the earth and avenge our blood?"
REV|6|11|Then each of them was given a white robe, and they were told to wait a little longer, until the number of their fellow servants and brothers who were to be killed as they had been was completed.
REV|6|12|I watched as he opened the sixth seal. There was a great earthquake. The sun turned black like sackcloth made of goat hair, the whole moon turned blood red,
REV|6|13|and the stars in the sky fell to earth, as late figs drop from a fig tree when shaken by a strong wind.
REV|6|14|The sky receded like a scroll, rolling up, and every mountain and island was removed from its place.
REV|6|15|Then the kings of the earth, the princes, the generals, the rich, the mighty, and every slave and every free man hid in caves and among the rocks of the mountains.
REV|6|16|They called to the mountains and the rocks, "Fall on us and hide us from the face of him who sits on the throne and from the wrath of the Lamb!
REV|6|17|For the great day of their wrath has come, and who can stand?"
REV|7|1|After this I saw four angels standing at the four corners of the earth, holding back the four winds of the earth to prevent any wind from blowing on the land or on the sea or on any tree.
REV|7|2|Then I saw another angel coming up from the east, having the seal of the living God. He called out in a loud voice to the four angels who had been given power to harm the land and the sea:
REV|7|3|"Do not harm the land or the sea or the trees until we put a seal on the foreheads of the servants of our God."
REV|7|4|Then I heard the number of those who were sealed: 144,000 from all the tribes of Israel.
REV|7|5|From the tribe of Judah 12,000 were sealed, from the tribe of Reuben 12,000, from the tribe of Gad 12,000,
REV|7|6|from the tribe of Asher 12,000, from the tribe of Naphtali 12,000, from the tribe of Manasseh 12,000,
REV|7|7|from the tribe of Simeon 12,000, from the tribe of Levi 12,000, from the tribe of Issachar 12,000,
REV|7|8|from the tribe of Zebulun 12,000, from the tribe of Joseph 12,000, from the tribe of Benjamin 12,000.
REV|7|9|After this I looked and there before me was a great multitude that no one could count, from every nation, tribe, people and language, standing before the throne and in front of the Lamb. They were wearing white robes and were holding palm branches in their hands.
REV|7|10|And they cried out in a loud voice: "Salvation belongs to our God, who sits on the throne, and to the Lamb."
REV|7|11|All the angels were standing around the throne and around the elders and the four living creatures. They fell down on their faces before the throne and worshiped God,
REV|7|12|saying: "Amen! Praise and glory and wisdom and thanks and honor and power and strength be to our God for ever and ever. Amen!"
REV|7|13|Then one of the elders asked me, "These in white robes--who are they, and where did they come from?"
REV|7|14|I answered, "Sir, you know."
REV|7|15|And he said, "These are they who have come out of the great tribulation; they have washed their robes and made them white in the blood of the Lamb. Therefore, "they are before the throne of God and serve him day and night in his temple; and he who sits on the throne will spread his tent over them.
REV|7|16|Never again will they hunger; never again will they thirst. The sun will not beat upon them, nor any scorching heat.
REV|7|17|For the Lamb at the center of the throne will be their shepherd; he will lead them to springs of living water. And God will wipe away every tear from their eyes."
REV|8|1|When he opened the seventh seal, there was silence in heaven for about half an hour.
REV|8|2|And I saw the seven angels who stand before God, and to them were given seven trumpets.
REV|8|3|Another angel, who had a golden censer, came and stood at the altar. He was given much incense to offer, with the prayers of all the saints, on the golden altar before the throne.
REV|8|4|The smoke of the incense, together with the prayers of the saints, went up before God from the angel's hand.
REV|8|5|Then the angel took the censer, filled it with fire from the altar, and hurled it on the earth; and there came peals of thunder, rumblings, flashes of lightning and an earthquake.
REV|8|6|Then the seven angels who had the seven trumpets prepared to sound them.
REV|8|7|The first angel sounded his trumpet, and there came hail and fire mixed with blood, and it was hurled down upon the earth. A third of the earth was burned up, a third of the trees were burned up, and all the green grass was burned up.
REV|8|8|The second angel sounded his trumpet, and something like a huge mountain, all ablaze, was thrown into the sea. A third of the sea turned into blood,
REV|8|9|a third of the living creatures in the sea died, and a third of the ships were destroyed.
REV|8|10|The third angel sounded his trumpet, and a great star, blazing like a torch, fell from the sky on a third of the rivers and on the springs of water--
REV|8|11|the name of the star is Wormwood. A third of the waters turned bitter, and many people died from the waters that had become bitter.
REV|8|12|The fourth angel sounded his trumpet, and a third of the sun was struck, a third of the moon, and a third of the stars, so that a third of them turned dark. A third of the day was without light, and also a third of the night.
REV|8|13|As I watched, I heard an eagle that was flying in midair call out in a loud voice: "Woe! Woe! Woe to the inhabitants of the earth, because of the trumpet blasts about to be sounded by the other three angels!"
REV|9|1|The fifth angel sounded his trumpet, and I saw a star that had fallen from the sky to the earth. The star was given the key to the shaft of the Abyss.
REV|9|2|When he opened the Abyss, smoke rose from it like the smoke from a gigantic furnace. The sun and sky were darkened by the smoke from the Abyss.
REV|9|3|And out of the smoke locusts came down upon the earth and were given power like that of scorpions of the earth.
REV|9|4|They were told not to harm the grass of the earth or any plant or tree, but only those people who did not have the seal of God on their foreheads.
REV|9|5|They were not given power to kill them, but only to torture them for five months. And the agony they suffered was like that of the sting of a scorpion when it strikes a man.
REV|9|6|During those days men will seek death, but will not find it; they will long to die, but death will elude them.
REV|9|7|The locusts looked like horses prepared for battle. On their heads they wore something like crowns of gold, and their faces resembled human faces.
REV|9|8|Their hair was like women's hair, and their teeth were like lions' teeth.
REV|9|9|They had breastplates like breastplates of iron, and the sound of their wings was like the thundering of many horses and chariots rushing into battle.
REV|9|10|They had tails and stings like scorpions, and in their tails they had power to torment people for five months.
REV|9|11|They had as king over them the angel of the Abyss, whose name in Hebrew is Abaddon, and in Greek, Apollyon.
REV|9|12|The first woe is past; two other woes are yet to come.
REV|9|13|The sixth angel sounded his trumpet, and I heard a voice coming from the horns of the golden altar that is before God.
REV|9|14|It said to the sixth angel who had the trumpet, "Release the four angels who are bound at the great river Euphrates."
REV|9|15|And the four angels who had been kept ready for this very hour and day and month and year were released to kill a third of mankind.
REV|9|16|The number of the mounted troops was two hundred million. I heard their number.
REV|9|17|The horses and riders I saw in my vision looked like this: Their breastplates were fiery red, dark blue, and yellow as sulfur. The heads of the horses resembled the heads of lions, and out of their mouths came fire, smoke and sulfur.
REV|9|18|A third of mankind was killed by the three plagues of fire, smoke and sulfur that came out of their mouths.
REV|9|19|The power of the horses was in their mouths and in their tails; for their tails were like snakes, having heads with which they inflict injury.
REV|9|20|The rest of mankind that were not killed by these plagues still did not repent of the work of their hands; they did not stop worshiping demons, and idols of gold, silver, bronze, stone and wood--idols that cannot see or hear or walk.
REV|9|21|Nor did they repent of their murders, their magic arts, their sexual immorality or their thefts.
REV|10|1|Then I saw another mighty angel coming down from heaven. He was robed in a cloud, with a rainbow above his head; his face was like the sun, and his legs were like fiery pillars.
REV|10|2|He was holding a little scroll, which lay open in his hand. He planted his right foot on the sea and his left foot on the land,
REV|10|3|and he gave a loud shout like the roar of a lion. When he shouted, the voices of the seven thunders spoke.
REV|10|4|And when the seven thunders spoke, I was about to write; but I heard a voice from heaven say, "Seal up what the seven thunders have said and do not write it down."
REV|10|5|Then the angel I had seen standing on the sea and on the land raised his right hand to heaven.
REV|10|6|And he swore by him who lives for ever and ever, who created the heavens and all that is in them, the earth and all that is in it, and the sea and all that is in it, and said, "There will be no more delay!
REV|10|7|But in the days when the seventh angel is about to sound his trumpet, the mystery of God will be accomplished, just as he announced to his servants the prophets."
REV|10|8|Then the voice that I had heard from heaven spoke to me once more: "Go, take the scroll that lies open in the hand of the angel who is standing on the sea and on the land."
REV|10|9|So I went to the angel and asked him to give me the little scroll. He said to me, "Take it and eat it. It will turn your stomach sour, but in your mouth it will be as sweet as honey."
REV|10|10|I took the little scroll from the angel's hand and ate it. It tasted as sweet as honey in my mouth, but when I had eaten it, my stomach turned sour.
REV|10|11|Then I was told, "You must prophesy again about many peoples, nations, languages and kings."
REV|11|1|I was given a reed like a measuring rod and was told, "Go and measure the temple of God and the altar, and count the worshipers there.
REV|11|2|But exclude the outer court; do not measure it, because it has been given to the Gentiles. They will trample on the holy city for 42 months.
REV|11|3|And I will give power to my two witnesses, and they will prophesy for 1,260 days, clothed in sackcloth."
REV|11|4|These are the two olive trees and the two lampstands that stand before the Lord of the earth.
REV|11|5|If anyone tries to harm them, fire comes from their mouths and devours their enemies. This is how anyone who wants to harm them must die.
REV|11|6|These men have power to shut up the sky so that it will not rain during the time they are prophesying; and they have power to turn the waters into blood and to strike the earth with every kind of plague as often as they want.
REV|11|7|Now when they have finished their testimony, the beast that comes up from the Abyss will attack them, and overpower and kill them.
REV|11|8|Their bodies will lie in the street of the great city, which is figuratively called Sodom and Egypt, where also their Lord was crucified.
REV|11|9|For three and a half days men from every people, tribe, language and nation will gaze on their bodies and refuse them burial.
REV|11|10|The inhabitants of the earth will gloat over them and will celebrate by sending each other gifts, because these two prophets had tormented those who live on the earth.
REV|11|11|But after the three and a half days a breath of life from God entered them, and they stood on their feet, and terror struck those who saw them.
REV|11|12|Then they heard a loud voice from heaven saying to them, "Come up here." And they went up to heaven in a cloud, while their enemies looked on.
REV|11|13|At that very hour there was a severe earthquake and a tenth of the city collapsed. Seven thousand people were killed in the earthquake, and the survivors were terrified and gave glory to the God of heaven.
REV|11|14|The second woe has passed; the third woe is coming soon.
REV|11|15|The seventh angel sounded his trumpet, and there were loud voices in heaven, which said: "The kingdom of the world has become the kingdom of our Lord and of his Christ, and he will reign for ever and ever."
REV|11|16|And the twenty-four elders, who were seated on their thrones before God, fell on their faces and worshiped God,
REV|11|17|saying: "We give thanks to you, Lord God Almighty, the One who is and who was, because you have taken your great power and have begun to reign.
REV|11|18|The nations were angry; and your wrath has come. The time has come for judging the dead, and for rewarding your servants the prophets and your saints and those who reverence your name, both small and great--and for destroying those who destroy the earth."
REV|11|19|Then God's temple in heaven was opened, and within his temple was seen the ark of his covenant. And there came flashes of lightning, rumblings, peals of thunder, an earthquake and a great hailstorm.
REV|12|1|A great and wondrous sign appeared in heaven: a woman clothed with the sun, with the moon under her feet and a crown of twelve stars on her head.
REV|12|2|She was pregnant and cried out in pain as she was about to give birth.
REV|12|3|Then another sign appeared in heaven: an enormous red dragon with seven heads and ten horns and seven crowns on his heads.
REV|12|4|His tail swept a third of the stars out of the sky and flung them to the earth. The dragon stood in front of the woman who was about to give birth, so that he might devour her child the moment it was born.
REV|12|5|She gave birth to a son, a male child, who will rule all the nations with an iron scepter. And her child was snatched up to God and to his throne.
REV|12|6|The woman fled into the desert to a place prepared for her by God, where she might be taken care of for 1,260 days.
REV|12|7|And there was war in heaven. Michael and his angels fought against the dragon, and the dragon and his angels fought back.
REV|12|8|But he was not strong enough, and they lost their place in heaven.
REV|12|9|The great dragon was hurled down--that ancient serpent called the devil, or Satan, who leads the whole world astray. He was hurled to the earth, and his angels with him.
REV|12|10|Then I heard a loud voice in heaven say: "Now have come the salvation and the power and the kingdom of our God, and the authority of his Christ. For the accuser of our brothers, who accuses them before our God day and night, has been hurled down.
REV|12|11|They overcame him by the blood of the Lamb and by the word of their testimony; they did not love their lives so much as to shrink from death.
REV|12|12|Therefore rejoice, you heavens and you who dwell in them! But woe to the earth and the sea, because the devil has gone down to you! He is filled with fury, because he knows that his time is short."
REV|12|13|When the dragon saw that he had been hurled to the earth, he pursued the woman who had given birth to the male child.
REV|12|14|The woman was given the two wings of a great eagle, so that she might fly to the place prepared for her in the desert, where she would be taken care of for a time, times and half a time, out of the serpent's reach.
REV|12|15|Then from his mouth the serpent spewed water like a river, to overtake the woman and sweep her away with the torrent.
REV|12|16|But the earth helped the woman by opening its mouth and swallowing the river that the dragon had spewed out of his mouth.
REV|12|17|Then the dragon was enraged at the woman and went off to make war against the rest of her offspring--those who obey God's commandments and hold to the testimony of Jesus.
REV|13|1|And the dragon stood on the shore of the sea.
REV|13|2|And I saw a beast coming out of the sea. He had ten horns and seven heads, with ten crowns on his horns, and on each head a blasphemous name. The beast I saw resembled a leopard, but had feet like those of a bear and a mouth like that of a lion. The dragon gave the beast his power and his throne and great authority.
REV|13|3|One of the heads of the beast seemed to have had a fatal wound, but the fatal wound had been healed. The whole world was astonished and followed the beast.
REV|13|4|Men worshiped the dragon because he had given authority to the beast, and they also worshiped the beast and asked, "Who is like the beast? Who can make war against him?"
REV|13|5|The beast was given a mouth to utter proud words and blasphemies and to exercise his authority for forty-two months.
REV|13|6|He opened his mouth to blaspheme God, and to slander his name and his dwelling place and those who live in heaven.
REV|13|7|He was given power to make war against the saints and to conquer them. And he was given authority over every tribe, people, language and nation.
REV|13|8|All inhabitants of the earth will worship the beast--all whose names have not been written in the book of life belonging to the Lamb that was slain from the creation of the world.
REV|13|9|He who has an ear, let him hear.
REV|13|10|If anyone is to go into captivity, into captivity he will go. If anyone is to be killed with the sword, with the sword he will be killed. This calls for patient endurance and faithfulness on the part of the saints.
REV|13|11|Then I saw another beast, coming out of the earth. He had two horns like a lamb, but he spoke like a dragon.
REV|13|12|He exercised all the authority of the first beast on his behalf, and made the earth and its inhabitants worship the first beast, whose fatal wound had been healed.
REV|13|13|And he performed great and miraculous signs, even causing fire to come down from heaven to earth in full view of men.
REV|13|14|Because of the signs he was given power to do on behalf of the first beast, he deceived the inhabitants of the earth. He ordered them to set up an image in honor of the beast who was wounded by the sword and yet lived.
REV|13|15|He was given power to give breath to the image of the first beast, so that it could speak and cause all who refused to worship the image to be killed.
REV|13|16|He also forced everyone, small and great, rich and poor, free and slave, to receive a mark on his right hand or on his forehead,
REV|13|17|so that no one could buy or sell unless he had the mark, which is the name of the beast or the number of his name.
REV|13|18|This calls for wisdom. If anyone has insight, let him calculate the number of the beast, for it is man's number. His number is 666.
REV|14|1|Then I looked, and there before me was the Lamb, standing on Mount Zion, and with him 144,000 who had his name and his Father's name written on their foreheads.
REV|14|2|And I heard a sound from heaven like the roar of rushing waters and like a loud peal of thunder. The sound I heard was like that of harpists playing their harps.
REV|14|3|And they sang a new song before the throne and before the four living creatures and the elders. No one could learn the song except the 144,000 who had been redeemed from the earth.
REV|14|4|These are those who did not defile themselves with women, for they kept themselves pure. They follow the Lamb wherever he goes. They were purchased from among men and offered as firstfruits to God and the Lamb.
REV|14|5|No lie was found in their mouths; they are blameless.
REV|14|6|Then I saw another angel flying in midair, and he had the eternal gospel to proclaim to those who live on the earth--to every nation, tribe, language and people.
REV|14|7|He said in a loud voice, "Fear God and give him glory, because the hour of his judgment has come. Worship him who made the heavens, the earth, the sea and the springs of water."
REV|14|8|A second angel followed and said, "Fallen! Fallen is Babylon the Great, which made all the nations drink the maddening wine of her adulteries."
REV|14|9|A third angel followed them and said in a loud voice: "If anyone worships the beast and his image and receives his mark on the forehead or on the hand,
REV|14|10|he, too, will drink of the wine of God's fury, which has been poured full strength into the cup of his wrath. He will be tormented with burning sulfur in the presence of the holy angels and of the Lamb.
REV|14|11|And the smoke of their torment rises for ever and ever. There is no rest day or night for those who worship the beast and his image, or for anyone who receives the mark of his name."
REV|14|12|This calls for patient endurance on the part of the saints who obey God's commandments and remain faithful to Jesus.
REV|14|13|Then I heard a voice from heaven say, "Write: Blessed are the dead who die in the Lord from now on.Yes," says the Spirit, "they will rest from their labor, for their deeds will follow them."
REV|14|14|I looked, and there before me was a white cloud, and seated on the cloud was one "like a son of man" with a crown of gold on his head and a sharp sickle in his hand.
REV|14|15|Then another angel came out of the temple and called in a loud voice to him who was sitting on the cloud, "Take your sickle and reap, because the time to reap has come, for the harvest of the earth is ripe."
REV|14|16|So he who was seated on the cloud swung his sickle over the earth, and the earth was harvested.
REV|14|17|Another angel came out of the temple in heaven, and he too had a sharp sickle.
REV|14|18|Still another angel, who had charge of the fire, came from the altar and called in a loud voice to him who had the sharp sickle, "Take your sharp sickle and gather the clusters of grapes from the earth's vine, because its grapes are ripe."
REV|14|19|The angel swung his sickle on the earth, gathered its grapes and threw them into the great winepress of God's wrath.
REV|14|20|They were trampled in the winepress outside the city, and blood flowed out of the press, rising as high as the horses' bridles for a distance of 1,600 stadia.
REV|15|1|I saw in heaven another great and marvelous sign: seven angels with the seven last plagues--last, because with them God's wrath is completed.
REV|15|2|And I saw what looked like a sea of glass mixed with fire and, standing beside the sea, those who had been victorious over the beast and his image and over the number of his name. They held harps given them by God
REV|15|3|and sang the song of Moses the servant of God and the song of the Lamb: "Great and marvelous are your deeds, Lord God Almighty. Just and true are your ways, King of the ages.
REV|15|4|Who will not fear you, O Lord, and bring glory to your name? For you alone are holy. All nations will come and worship before you, for your righteous acts have been revealed."
REV|15|5|After this I looked and in heaven the temple, that is, the tabernacle of the Testimony, was opened.
REV|15|6|Out of the temple came the seven angels with the seven plagues. They were dressed in clean, shining linen and wore golden sashes around their chests.
REV|15|7|Then one of the four living creatures gave to the seven angels seven golden bowls filled with the wrath of God, who lives for ever and ever.
REV|15|8|And the temple was filled with smoke from the glory of God and from his power, and no one could enter the temple until the seven plagues of the seven angels were completed.
REV|16|1|Then I heard a loud voice from the temple saying to the seven angels, "Go, pour out the seven bowls of God's wrath on the earth."
REV|16|2|The first angel went and poured out his bowl on the land, and ugly and painful sores broke out on the people who had the mark of the beast and worshiped his image.
REV|16|3|The second angel poured out his bowl on the sea, and it turned into blood like that of a dead man, and every living thing in the sea died.
REV|16|4|The third angel poured out his bowl on the rivers and springs of water, and they became blood.
REV|16|5|Then I heard the angel in charge of the waters say: "You are just in these judgments, you who are and who were, the Holy One, because you have so judged;
REV|16|6|for they have shed the blood of your saints and prophets, and you have given them blood to drink as they deserve."
REV|16|7|And I heard the altar respond: "Yes, Lord God Almighty, true and just are your judgments."
REV|16|8|The fourth angel poured out his bowl on the sun, and the sun was given power to scorch people with fire.
REV|16|9|They were seared by the intense heat and they cursed the name of God, who had control over these plagues, but they refused to repent and glorify him.
REV|16|10|The fifth angel poured out his bowl on the throne of the beast, and his kingdom was plunged into darkness. Men gnawed their tongues in agony
REV|16|11|and cursed the God of heaven because of their pains and their sores, but they refused to repent of what they had done.
REV|16|12|The sixth angel poured out his bowl on the great river Euphrates, and its water was dried up to prepare the way for the kings from the East.
REV|16|13|Then I saw three evil spirits that looked like frogs; they came out of the mouth of the dragon, out of the mouth of the beast and out of the mouth of the false prophet.
REV|16|14|They are spirits of demons performing miraculous signs, and they go out to the kings of the whole world, to gather them for the battle on the great day of God Almighty.
REV|16|15|"Behold, I come like a thief! Blessed is he who stays awake and keeps his clothes with him, so that he may not go naked and be shamefully exposed."
REV|16|16|Then they gathered the kings together to the place that in Hebrew is called Armageddon.
REV|16|17|The seventh angel poured out his bowl into the air, and out of the temple came a loud voice from the throne, saying, "It is done!"
REV|16|18|Then there came flashes of lightning, rumblings, peals of thunder and a severe earthquake. No earthquake like it has ever occurred since man has been on earth, so tremendous was the quake.
REV|16|19|The great city split into three parts, and the cities of the nations collapsed. God remembered Babylon the Great and gave her the cup filled with the wine of the fury of his wrath.
REV|16|20|Every island fled away and the mountains could not be found.
REV|16|21|From the sky huge hailstones of about a hundred pounds each fell upon men. And they cursed God on account of the plague of hail, because the plague was so terrible.
REV|17|1|One of the seven angels who had the seven bowls came and said to me, "Come, I will show you the punishment of the great prostitute, who sits on many waters.
REV|17|2|With her the kings of the earth committed adultery and the inhabitants of the earth were intoxicated with the wine of her adulteries."
REV|17|3|Then the angel carried me away in the Spirit into a desert. There I saw a woman sitting on a scarlet beast that was covered with blasphemous names and had seven heads and ten horns.
REV|17|4|The woman was dressed in purple and scarlet, and was glittering with gold, precious stones and pearls. She held a golden cup in her hand, filled with abominable things and the filth of her adulteries.
REV|17|5|This title was written on her forehead: MYSTERY BABYLON THE GREAT THE MOTHER OF PROSTITUTES AND OF THE ABOMINATIONS OF THE EARTH.
REV|17|6|I saw that the woman was drunk with the blood of the saints, the blood of those who bore testimony to Jesus.
REV|17|7|When I saw her, I was greatly astonished. Then the angel said to me: "Why are you astonished? I will explain to you the mystery of the woman and of the beast she rides, which has the seven heads and ten horns.
REV|17|8|The beast, which you saw, once was, now is not, and will come up out of the Abyss and go to his destruction. The inhabitants of the earth whose names have not been written in the book of life from the creation of the world will be astonished when they see the beast, because he once was, now is not, and yet will come.
REV|17|9|"This calls for a mind with wisdom. The seven heads are seven hills on which the woman sits.
REV|17|10|They are also seven kings. Five have fallen, one is, the other has not yet come; but when he does come, he must remain for a little while.
REV|17|11|The beast who once was, and now is not, is an eighth king. He belongs to the seven and is going to his destruction.
REV|17|12|"The ten horns you saw are ten kings who have not yet received a kingdom, but who for one hour will receive authority as kings along with the beast.
REV|17|13|They have one purpose and will give their power and authority to the beast.
REV|17|14|They will make war against the Lamb, but the Lamb will overcome them because he is Lord of lords and King of kings--and with him will be his called, chosen and faithful followers."
REV|17|15|Then the angel said to me, "The waters you saw, where the prostitute sits, are peoples, multitudes, nations and languages.
REV|17|16|The beast and the ten horns you saw will hate the prostitute. They will bring her to ruin and leave her naked; they will eat her flesh and burn her with fire.
REV|17|17|For God has put it into their hearts to accomplish his purpose by agreeing to give the beast their power to rule, until God's words are fulfilled.
REV|17|18|The woman you saw is the great city that rules over the kings of the earth."
REV|18|1|After this I saw another angel coming down from heaven. He had great authority, and the earth was illuminated by his splendor.
REV|18|2|With a mighty voice he shouted: "Fallen! Fallen is Babylon the Great! She has become a home for demons and a haunt for every evil spirit, a haunt for every unclean and detestable bird.
REV|18|3|For all the nations have drunk the maddening wine of her adulteries. The kings of the earth committed adultery with her, and the merchants of the earth grew rich from her excessive luxuries."
REV|18|4|Then I heard another voice from heaven say: "Come out of her, my people, so that you will not share in her sins, so that you will not receive any of her plagues;
REV|18|5|for her sins are piled up to heaven, and God has remembered her crimes.
REV|18|6|Give back to her as she has given; pay her back double for what she has done. Mix her a double portion from her own cup.
REV|18|7|Give her as much torture and grief as the glory and luxury she gave herself. In her heart she boasts, 'I sit as queen; I am not a widow, and I will never mourn.'
REV|18|8|Therefore in one day her plagues will overtake her: death, mourning and famine. She will be consumed by fire, for mighty is the Lord God who judges her.
REV|18|9|"When the kings of the earth who committed adultery with her and shared her luxury see the smoke of her burning, they will weep and mourn over her.
REV|18|10|Terrified at her torment, they will stand far off and cry: "'Woe! Woe, O great city, O Babylon, city of power! In one hour your doom has come!'
REV|18|11|"The merchants of the earth will weep and mourn over her because no one buys their cargoes any more--
REV|18|12|cargoes of gold, silver, precious stones and pearls; fine linen, purple, silk and scarlet cloth; every sort of citron wood, and articles of every kind made of ivory, costly wood, bronze, iron and marble;
REV|18|13|cargoes of cinnamon and spice, of incense, myrrh and frankincense, of wine and olive oil, of fine flour and wheat; cattle and sheep; horses and carriages; and bodies and souls of men.
REV|18|14|"They will say, 'The fruit you longed for is gone from you. All your riches and splendor have vanished, never to be recovered.'
REV|18|15|The merchants who sold these things and gained their wealth from her will stand far off, terrified at her torment. They will weep and mourn
REV|18|16|and cry out: "'Woe! Woe, O great city, dressed in fine linen, purple and scarlet, and glittering with gold, precious stones and pearls!
REV|18|17|In one hour such great wealth has been brought to ruin!'
REV|18|18|"Every sea captain, and all who travel by ship, the sailors, and all who earn their living from the sea, will stand far off. When they see the smoke of her burning, they will exclaim, 'Was there ever a city like this great city?'
REV|18|19|They will throw dust on their heads, and with weeping and mourning cry out: "'Woe! Woe, O great city, where all who had ships on the sea became rich through her wealth! In one hour she has been brought to ruin!
REV|18|20|Rejoice over her, O heaven! Rejoice, saints and apostles and prophets! God has judged her for the way she treated you.'"
REV|18|21|Then a mighty angel picked up a boulder the size of a large millstone and threw it into the sea, and said: "With such violence the great city of Babylon will be thrown down, never to be found again.
REV|18|22|The music of harpists and musicians, flute players and trumpeters, will never be heard in you again. No workman of any trade will ever be found in you again. The sound of a millstone will never be heard in you again.
REV|18|23|The light of a lamp will never shine in you again. The voice of bridegroom and bride will never be heard in you again. Your merchants were the world's great men. By your magic spell all the nations were led astray.
REV|18|24|In her was found the blood of prophets and of the saints, and of all who have been killed on the earth."
REV|19|1|After this I heard what sounded like the roar of a great multitude in heaven shouting: "Hallelujah! Salvation and glory and power belong to our God,
REV|19|2|for true and just are his judgments. He has condemned the great prostitute who corrupted the earth by her adulteries. He has avenged on her the blood of his servants."
REV|19|3|And again they shouted: "Hallelujah! The smoke from her goes up for ever and ever."
REV|19|4|The twenty-four elders and the four living creatures fell down and worshiped God, who was seated on the throne. And they cried: "Amen, Hallelujah!"
REV|19|5|Then a voice came from the throne, saying: "Praise our God, all you his servants, you who fear him, both small and great!"
REV|19|6|Then I heard what sounded like a great multitude, like the roar of rushing waters and like loud peals of thunder, shouting: "Hallelujah! For our Lord God Almighty reigns.
REV|19|7|Let us rejoice and be glad and give him glory! For the wedding of the Lamb has come, and his bride has made herself ready.
REV|19|8|Fine linen, bright and clean, was given her to wear." (Fine linen stands for the righteous acts of the saints.)
REV|19|9|Then the angel said to me, "Write: 'Blessed are those who are invited to the wedding supper of the Lamb!'" And he added, "These are the true words of God."
REV|19|10|At this I fell at his feet to worship him. But he said to me, "Do not do it! I am a fellow servant with you and with your brothers who hold to the testimony of Jesus. Worship God! For the testimony of Jesus is the spirit of prophecy."
REV|19|11|I saw heaven standing open and there before me was a white horse, whose rider is called Faithful and True. With justice he judges and makes war.
REV|19|12|His eyes are like blazing fire, and on his head are many crowns. He has a name written on him that no one knows but he himself.
REV|19|13|He is dressed in a robe dipped in blood, and his name is the Word of God.
REV|19|14|The armies of heaven were following him, riding on white horses and dressed in fine linen, white and clean.
REV|19|15|Out of his mouth comes a sharp sword with which to strike down the nations. "He will rule them with an iron scepter." He treads the winepress of the fury of the wrath of God Almighty.
REV|19|16|On his robe and on his thigh he has this name written: KING OF KINGS AND LORD OF LORDS.
REV|19|17|And I saw an angel standing in the sun, who cried in a loud voice to all the birds flying in midair, "Come, gather together for the great supper of God,
REV|19|18|so that you may eat the flesh of kings, generals, and mighty men, of horses and their riders, and the flesh of all people, free and slave, small and great."
REV|19|19|Then I saw the beast and the kings of the earth and their armies gathered together to make war against the rider on the horse and his army.
REV|19|20|But the beast was captured, and with him the false prophet who had performed the miraculous signs on his behalf. With these signs he had deluded those who had received the mark of the beast and worshiped his image. The two of them were thrown alive into the fiery lake of burning sulfur.
REV|19|21|The rest of them were killed with the sword that came out of the mouth of the rider on the horse, and all the birds gorged themselves on their flesh.
REV|20|1|And I saw an angel coming down out of heaven, having the key to the Abyss and holding in his hand a great chain.
REV|20|2|He seized the dragon, that ancient serpent, who is the devil, or Satan, and bound him for a thousand years.
REV|20|3|He threw him into the Abyss, and locked and sealed it over him, to keep him from deceiving the nations anymore until the thousand years were ended. After that, he must be set free for a short time.
REV|20|4|I saw thrones on which were seated those who had been given authority to judge. And I saw the souls of those who had been beheaded because of their testimony for Jesus and because of the word of God. They had not worshiped the beast or his image and had not received his mark on their foreheads or their hands. They came to life and reigned with Christ a thousand years.
REV|20|5|(The rest of the dead did not come to life until the thousand years were ended.) This is the first resurrection.
REV|20|6|Blessed and holy are those who have part in the first resurrection. The second death has no power over them, but they will be priests of God and of Christ and will reign with him for a thousand years.
REV|20|7|When the thousand years are over, Satan will be released from his prison
REV|20|8|and will go out to deceive the nations in the four corners of the earth--Gog and Magog--to gather them for battle. In number they are like the sand on the seashore.
REV|20|9|They marched across the breadth of the earth and surrounded the camp of God's people, the city he loves. But fire came down from heaven and devoured them.
REV|20|10|And the devil, who deceived them, was thrown into the lake of burning sulfur, where the beast and the false prophet had been thrown. They will be tormented day and night for ever and ever.
REV|20|11|Then I saw a great white throne and him who was seated on it. Earth and sky fled from his presence, and there was no place for them.
REV|20|12|And I saw the dead, great and small, standing before the throne, and books were opened. Another book was opened, which is the book of life. The dead were judged according to what they had done as recorded in the books.
REV|20|13|The sea gave up the dead that were in it, and death and Hades gave up the dead that were in them, and each person was judged according to what he had done.
REV|20|14|Then death and Hades were thrown into the lake of fire. The lake of fire is the second death.
REV|20|15|If anyone's name was not found written in the book of life, he was thrown into the lake of fire.
REV|21|1|Then I saw a new heaven and a new earth, for the first heaven and the first earth had passed away, and there was no longer any sea.
REV|21|2|I saw the Holy City, the new Jerusalem, coming down out of heaven from God, prepared as a bride beautifully dressed for her husband.
REV|21|3|And I heard a loud voice from the throne saying, "Now the dwelling of God is with men, and he will live with them. They will be his people, and God himself will be with them and be their God.
REV|21|4|He will wipe every tear from their eyes. There will be no more death or mourning or crying or pain, for the old order of things has passed away."
REV|21|5|He who was seated on the throne said, "I am making everything new!" Then he said, "Write this down, for these words are trustworthy and true."
REV|21|6|He said to me: "It is done. I am the Alpha and the Omega, the Beginning and the End. To him who is thirsty I will give to drink without cost from the spring of the water of life.
REV|21|7|He who overcomes will inherit all this, and I will be his God and he will be my son.
REV|21|8|But the cowardly, the unbelieving, the vile, the murderers, the sexually immoral, those who practice magic arts, the idolaters and all liars--their place will be in the fiery lake of burning sulfur. This is the second death."
REV|21|9|One of the seven angels who had the seven bowls full of the seven last plagues came and said to me, "Come, I will show you the bride, the wife of the Lamb."
REV|21|10|And he carried me away in the Spirit to a mountain great and high, and showed me the Holy City, Jerusalem, coming down out of heaven from God.
REV|21|11|It shone with the glory of God, and its brilliance was like that of a very precious jewel, like a jasper, clear as crystal.
REV|21|12|It had a great, high wall with twelve gates, and with twelve angels at the gates. On the gates were written the names of the twelve tribes of Israel.
REV|21|13|There were three gates on the east, three on the north, three on the south and three on the west.
REV|21|14|The wall of the city had twelve foundations, and on them were the names of the twelve apostles of the Lamb.
REV|21|15|The angel who talked with me had a measuring rod of gold to measure the city, its gates and its walls.
REV|21|16|The city was laid out like a square, as long as it was wide. He measured the city with the rod and found it to be 12,000 stadia in length, and as wide and high as it is long.
REV|21|17|He measured its wall and it was 144 cubits thick, by man's measurement, which the angel was using.
REV|21|18|The wall was made of jasper, and the city of pure gold, as pure as glass.
REV|21|19|The foundations of the city walls were decorated with every kind of precious stone. The first foundation was jasper, the second sapphire, the third chalcedony, the fourth emerald,
REV|21|20|the fifth sardonyx, the sixth carnelian, the seventh chrysolite, the eighth beryl, the ninth topaz, the tenth chrysoprase, the eleventh jacinth, and the twelfth amethyst.
REV|21|21|The twelve gates were twelve pearls, each gate made of a single pearl. The great street of the city was of pure gold, like transparent glass.
REV|21|22|I did not see a temple in the city, because the Lord God Almighty and the Lamb are its temple.
REV|21|23|The city does not need the sun or the moon to shine on it, for the glory of God gives it light, and the Lamb is its lamp.
REV|21|24|The nations will walk by its light, and the kings of the earth will bring their splendor into it.
REV|21|25|On no day will its gates ever be shut, for there will be no night there.
REV|21|26|The glory and honor of the nations will be brought into it.
REV|21|27|Nothing impure will ever enter it, nor will anyone who does what is shameful or deceitful, but only those whose names are written in the Lamb's book of life.
REV|22|1|Then the angel showed me the river of the water of life, as clear as crystal, flowing from the throne of God and of the Lamb
REV|22|2|down the middle of the great street of the city. On each side of the river stood the tree of life, bearing twelve crops of fruit, yielding its fruit every month. And the leaves of the tree are for the healing of the nations.
REV|22|3|No longer will there be any curse. The throne of God and of the Lamb will be in the city, and his servants will serve him.
REV|22|4|They will see his face, and his name will be on their foreheads.
REV|22|5|There will be no more night. They will not need the light of a lamp or the light of the sun, for the Lord God will give them light. And they will reign for ever and ever.
REV|22|6|The angel said to me, "These words are trustworthy and true. The Lord, the God of the spirits of the prophets, sent his angel to show his servants the things that must soon take place."
REV|22|7|"Behold, I am coming soon! Blessed is he who keeps the words of the prophecy in this book."
REV|22|8|I, John, am the one who heard and saw these things. And when I had heard and seen them, I fell down to worship at the feet of the angel who had been showing them to me.
REV|22|9|But he said to me, "Do not do it! I am a fellow servant with you and with your brothers the prophets and of all who keep the words of this book. Worship God!"
REV|22|10|Then he told me, "Do not seal up the words of the prophecy of this book, because the time is near.
REV|22|11|Let him who does wrong continue to do wrong; let him who is vile continue to be vile; let him who does right continue to do right; and let him who is holy continue to be holy."
REV|22|12|"Behold, I am coming soon! My reward is with me, and I will give to everyone according to what he has done.
REV|22|13|I am the Alpha and the Omega, the First and the Last, the Beginning and the End.
REV|22|14|"Blessed are those who wash their robes, that they may have the right to the tree of life and may go through the gates into the city.
REV|22|15|Outside are the dogs, those who practice magic arts, the sexually immoral, the murderers, the idolaters and everyone who loves and practices falsehood.
REV|22|16|"I, Jesus, have sent my angel to give you this testimony for the churches. I am the Root and the Offspring of David, and the bright Morning Star."
REV|22|17|The Spirit and the bride say, "Come!" And let him who hears say, "Come!" Whoever is thirsty, let him come; and whoever wishes, let him take the free gift of the water of life.
REV|22|18|I warn everyone who hears the words of the prophecy of this book: If anyone adds anything to them, God will add to him the plagues described in this book.
REV|22|19|And if anyone takes words away from this book of prophecy, God will take away from him his share in the tree of life and in the holy city, which are described in this book.
REV|22|20|He who testifies to these things says, "Yes, I am coming soon." Amen. Come, Lord Jesus.
REV|22|21|The grace of the Lord Jesus be with God's people. Amen.
