MIC|1|1|Слово Господне, которое было к Михею Морасфитину во дни Иоафама, Ахаза и Езекии, царей Иудейских, и которое открыто ему о Самарии и Иерусалиме.
MIC|1|2|Слушайте, все народы, внимай, земля и все, что наполняет ее! Да будет Господь Бог свидетелем против вас, Господь из святаго храма Своего!
MIC|1|3|Ибо вот, Господь исходит от места Своего, низойдет и наступит на высоты земли, –
MIC|1|4|и горы растают под Ним, долины распадутся, как воск от огня, как воды, льющиеся с крутизны.
MIC|1|5|Все это – за нечестие Иакова, за грех дома Израилева. От кого нечестие Иакова? не от Самарии ли? Кто [устроил] высоты в Иудее? не Иерусалим ли?
MIC|1|6|За то сделаю Самарию грудою развалин в поле, местом для разведения винограда; низрину в долину камни ее и обнажу основания ее.
MIC|1|7|Все истуканы ее будут разбиты и все любодейные дары ее сожжены будут огнем, и всех идолов ее предам разрушению, ибо из любодейных даров она устраивала их, на любодейные дары они и будут обращены.
MIC|1|8|Об этом буду я плакать и рыдать, буду ходить, как ограбленный и обнаженный, выть, как шакалы, и плакать, как страусы,
MIC|1|9|потому что болезненно поражение ее, дошло до Иуды, достигло даже до ворот народа моего, до Иерусалима.
MIC|1|10|Не объявляйте об этом в Гефе, не плачьте там громко; но в селении Офра покрой себя пеплом.
MIC|1|11|Переселяйтесь, жительницы Шафира, срамно обнаженные; не убежит и живущая в Цаане; плач в селении Ецель не даст вам остановиться в нем.
MIC|1|12|Горюет о своем добре жительница Марофы, ибо сошло бедствие от Господа к воротам Иерусалима.
MIC|1|13|Запрягай в колесницу быстрых, жительница Лахиса; ты – начало греха дщери Сионовой, ибо у тебя появились преступления Израиля.
MIC|1|14|Посему ты посылать будешь дары в Морешеф–Геф; но селения Ахзива будут обманом для царей Израилевых.
MIC|1|15|Еще наследника приведу к тебе, жительница Мореша; он пройдет до Одоллама, славы Израиля.
MIC|1|16|Сними с себя волосы, остригись, скорбя о нежно любимых сынах твоих; расширь из–за них лысину, как у линяющего орла, ибо они переселены будут от тебя.
MIC|2|1|Горе замышляющим беззаконие и на ложах своих придумывающим злодеяния, которые совершают утром на рассвете, потому что есть в руке их сила!
MIC|2|2|Пожелают полей и берут их силою, домов, – и отнимают их; обирают человека и его дом, мужа и его наследие.
MIC|2|3|Посему так говорит Господь: вот, Я помышляю навести на этот род такое бедствие, которого вы не свергнете с шеи вашей, и не будете ходить выпрямившись; ибо это время злое.
MIC|2|4|В тот день произнесут о вас притчу и будут плакать горьким плачем и говорить: "мы совершенно разорены! удел народа моего отдан другим; как возвратится ко мне! поля наши уже разделены иноплеменникам".
MIC|2|5|Посему не будет у тебя никого, кто бросил бы жребий для измерения в собрании пред Господом.
MIC|2|6|Не пророчествуйте, пророки; не пророчествуйте им, чтобы не постигло вас бесчестие.
MIC|2|7|О, называющийся домом Иакова! разве умалился Дух Господень? таковы ли действия Его? не благотворны ли слова Мои для того, кто поступает справедливо?
MIC|2|8|Народ же, который был прежде Моим, восстал как враг, и вы отнимаете как верхнюю, так и нижнюю одежду у проходящих мирно, отвращающихся войны.
MIC|2|9|Жен народа Моего вы изгоняете из приятных домов их; у детей их вы навсегда отнимаете украшение Мое.
MIC|2|10|Встаньте и уходите, ибо [страна] сия не есть место покоя; за нечистоту она будет разорена и притом жестоким разорением.
MIC|2|11|Если бы какой–либо ветреник выдумал ложь и сказал: "я буду проповедывать тебе о вине и сикере", то он и был бы угодным проповедником для этого народа.
MIC|2|12|Непременно соберу всего тебя, Иаков, непременно соединю остатки Израиля, совокуплю их воедино, как овец в Восоре, как стадо в овечьем загоне; зашумят они от многолюдства.
MIC|2|13|Перед ними пойдет стенорушитель; они сокрушат преграды, войдут сквозь ворота и выйдут ими; и царь их пойдет перед ними, а во главе их Господь.
MIC|3|1|И сказал я: слушайте, главы Иакова и князья дома Израилева: не вам ли должно знать правду?
MIC|3|2|А вы ненавидите доброе и любите злое; сдираете с них кожу их и плоть с костей их,
MIC|3|3|едите плоть народа Моего и сдираете с них кожу их, а кости их ломаете и дробите как бы в горшок, и плоть – как бы в котел.
MIC|3|4|И будут они взывать к Господу, но Он не услышит их и сокроет лице Свое от них на то время, как они злодействуют.
MIC|3|5|Так говорит Господь на пророков, вводящих в заблуждение народ Мой, которые грызут зубами своими – и проповедуют мир, а кто ничего не кладет им в рот, против того объявляют войну.
MIC|3|6|Посему ночь будет вам вместо видения, и тьма – вместо предвещаний; зайдет солнце над пророками и потемнеет день над ними.
MIC|3|7|И устыдятся прозорливцы, и посрамлены будут гадатели, и закроют уста свои все они, потому что не будет ответа от Бога.
MIC|3|8|А я исполнен силы Духа Господня, правоты и твердости, чтобы высказать Иакову преступление его и Израилю грех его.
MIC|3|9|Слушайте же это, главы дома Иаковлева и князья дома Израилева, гнушающиеся правосудием и искривляющие все прямое,
MIC|3|10|созидающие Сион кровью и Иерусалим – неправдою!
MIC|3|11|Главы его судят за подарки и священники его учат за плату, и пророки его предвещают за деньги, а между тем опираются на Господа, говоря: "не среди ли нас Господь? не постигнет нас беда!"
MIC|3|12|Посему за вас Сион распахан будет как поле, и Иерусалим сделается грудою развалин, и гора дома сего будет лесистым холмом.
MIC|4|1|И будет в последние дни: гора дома Господня поставлена будет во главу гор и возвысится над холмами, и потекут к ней народы.
MIC|4|2|И пойдут многие народы и скажут: придите, и взойдем на гору Господню и в дом Бога Иаковлева, и Он научит нас путям Своим, и будем ходить по стезям Его, ибо от Сиона выйдет закон и слово Господне – из Иерусалима.
MIC|4|3|И будет Он судить многие народы, и обличит многие племена в отдаленных странах; и перекуют они мечи свои на орала и копья свои – на серпы; не поднимет народ на народ меча, и не будут более учиться воевать.
MIC|4|4|Но каждый будет сидеть под своею виноградною лозою и под своею смоковницею, и никто не будет устрашать их, ибо уста Господа Саваофа изрекли это.
MIC|4|5|Ибо все народы ходят, каждый во имя своего бога; а мы будем ходить во имя Господа Бога нашего во веки веков.
MIC|4|6|В тот день, говорит Господь, соберу хромлющее и совокуплю разогнанное и тех, на кого Я навел бедствие.
MIC|4|7|И сделаю хромлющее остатком и далеко рассеянное сильным народом, и Господь будет царствовать над ними на горе Сионе отныне и до века.
MIC|4|8|А ты, башня стада, холм дщери Сиона! к тебе придет и возвратится прежнее владычество, царство – к дщерям Иерусалима.
MIC|4|9|Для чего же ты ныне так громко вопиешь? Разве нет у тебя царя? Или не стало у тебя советника, что тебя схватили муки, как рождающую?
MIC|4|10|Страдай и мучься болями, дщерь Сиона, как рождающая, ибо ныне ты выйдешь из города и будешь жить в поле, и дойдешь до Вавилона: там будешь спасена, там искупит тебя Господь от руки врагов твоих.
MIC|4|11|А теперь собрались против тебя многие народы и говорят: "да будет она осквернена, и да наглядится око наше на Сион!"
MIC|4|12|Но они не знают мыслей Господних и не разумеют совета Его, что Он собрал их как снопы на гумно.
MIC|4|13|Встань и молоти, дщерь Сиона, ибо Я сделаю рог твой железным и копыта твои сделаю медными, и сокрушишь многие народы, и посвятишь Господу стяжания их и богатства их Владыке всей земли.
MIC|5|1|Теперь ополчись, дщерь полчищ; обложили нас осадою, тростью будут бить по ланите судью Израилева.
MIC|5|2|И ты, Вифлеем–Ефрафа, мал ли ты между тысячами Иудиными? из тебя произойдет Мне Тот, Который должен быть Владыкою в Израиле и Которого происхождение из начала, от дней вечных.
MIC|5|3|Посему Он оставит их до времени, доколе не родит имеющая родить; тогда возвратятся к сынам Израиля и оставшиеся братья их.
MIC|5|4|И станет Он, и будет пасти в силе Господней, в величии имени Господа Бога Своего, и они будут жить безопасно, ибо тогда Он будет великим до краев земли.
MIC|5|5|И будет Он мир. Когда Ассур придет в нашу землю и вступит в наши чертоги, мы выставим против него семь пастырей и восемь князей.
MIC|5|6|И будут они пасти землю Ассура мечом и землю Немврода в самых воротах ее, и Он–то избавит от Ассура, когда тот придет в землю нашу и когда вступит в пределы наши.
MIC|5|7|И будет остаток Иакова среди многих народов как роса от Господа, как ливень на траве, и он не будет зависеть от человека и полагаться на сынов Адамовых.
MIC|5|8|И будет остаток Иакова между народами, среди многих племен, как лев среди зверей лесных, как скимен среди стада овец, который, когда выступит, то попирает и терзает, и никто не спасет от него.
MIC|5|9|Поднимется рука твоя над врагами твоими, и все неприятели твои будут истреблены.
MIC|5|10|И будет в тот день, говорит Господь: истреблю коней твоих из среды твоей и уничтожу колесницы твои,
MIC|5|11|истреблю города в земле твоей и разрушу все укрепления твои,
MIC|5|12|исторгну чародеяния из руки твоей, и гадающих по облакам не будет у тебя;
MIC|5|13|истреблю истуканов твоих и кумиров из среды твоей, и не будешь более поклоняться изделиям рук твоих.
MIC|5|14|Искореню из среды твоей священные рощи твои и разорю города твои.
MIC|5|15|И совершу в гневе и негодовании мщение над народами, которые будут непослушны.
MIC|6|1|Слушайте, что говорит Господь: встань, судись перед горами, и холмы да слышат голос твой!
MIC|6|2|Слушайте, горы, суд Господень, и вы, твердые основы земли: ибо у Господа суд с народом Своим, и с Израилем Он состязуется.
MIC|6|3|Народ Мой! что сделал Я тебе и чем отягощал тебя? отвечай Мне.
MIC|6|4|Я вывел тебя из земли Египетской и искупил тебя из дома рабства, и послал перед тобою Моисея, Аарона и Мариам.
MIC|6|5|Народ Мой! вспомни, что замышлял Валак, царь Моавитский, и что отвечал ему Валаам, сын Веоров, и что [происходило] от Ситтима до Галгал, чтобы познать тебе праведные действия Господни.
MIC|6|6|"С чем предстать мне пред Господом, преклониться пред Богом небесным? Предстать ли пред Ним со всесожжениями, с тельцами однолетними?
MIC|6|7|Но можно ли угодить Господу тысячами овнов или неисчетными потоками елея? Разве дам Ему первенца моего за преступление мое и плод чрева моего – за грех души моей?"
MIC|6|8|О, человек! сказано тебе, что – добро и чего требует от тебя Господь: действовать справедливо, любить дела милосердия и смиренномудренно ходить пред Богом твоим.
MIC|6|9|Глас Господа взывает к городу, и мудрость благоговеет пред именем Твоим: слушайте жезл и Того, Кто поставил его.
MIC|6|10|Не находятся ли и теперь в доме нечестивого сокровища нечестия и уменьшенная мера, отвратительная?
MIC|6|11|Могу ли я быть чистым с весами неверными и с обманчивыми гирями в суме?
MIC|6|12|Так как богачи его исполнены неправды, и жители его говорят ложь, и язык их есть обман в устах их,
MIC|6|13|то и Я неисцельно поражу тебя опустошением за грехи твои.
MIC|6|14|Ты будешь есть, и не будешь сыт; пустота будет внутри тебя; будешь хранить, но не убережешь, а что сбережешь, то предам мечу.
MIC|6|15|Будешь сеять, а жать не будешь; будешь давить оливки, и не будешь умащаться елеем; выжмешь виноградный сок, а вина пить не будешь.
MIC|6|16|Сохранились у вас обычаи Амврия и все дела дома Ахавова, и вы поступаете по советам их; и предам Я тебя опустошению и жителей твоих посмеянию, и вы понесете поругание народа Моего.
MIC|7|1|Горе мне! ибо со мною теперь – как по собрании летних плодов, как по уборке винограда: ни одной ягоды для еды, ни спелого плода, которого желает душа моя.
MIC|7|2|Не стало милосердых на земле, нет правдивых между людьми; все строят ковы, чтобы проливать кровь; каждый ставит брату своему сеть.
MIC|7|3|Руки их обращены к тому, чтобы уметь делать зло; начальник требует подарков, и судья судит за взятки, а вельможи высказывают злые хотения души своей и извращают дело.
MIC|7|4|Лучший из них – как терн, и справедливый – хуже колючей изгороди, день провозвестников Твоих, посещение Твое наступает; ныне постигнет их смятение.
MIC|7|5|Не верьте другу, не полагайтесь на приятеля; от лежащей на лоне твоем стереги двери уст твоих.
MIC|7|6|Ибо сын позорит отца, дочь восстает против матери, невестка – против свекрови своей; враги человеку – домашние его.
MIC|7|7|А я буду взирать на Господа, уповать на Бога спасения моего: Бог мой услышит меня.
MIC|7|8|Не радуйся ради меня, неприятельница моя! хотя я упал, но встану; хотя я во мраке, но Господь свет для меня.
MIC|7|9|Гнев Господень я буду нести, потому что согрешил пред Ним, доколе Он не решит дела моего и не совершит суда надо мною; тогда Он выведет меня на свет, и я увижу правду Его.
MIC|7|10|И увидит это неприятельница моя и стыд покроет ее, говорившую мне: "где Господь Бог твой?" Насмотрятся на нее глаза мои, как она будет попираема подобно грязи на улицах.
MIC|7|11|В день сооружения стен твоих, в этот день отдалится определение.
MIC|7|12|В тот день придут к тебе из Ассирии и городов Египетских, и от Египта до реки [Евфрата], и от моря до моря, и от горы до горы.
MIC|7|13|А земля та будет пустынею за [вину] жителей ее, за плоды деяний их.
MIC|7|14|Паси народ Твой жезлом Твоим, овец наследия Твоего, обитающих уединенно в лесу среди Кармила; да пасутся они на Васане и Галааде, как во дни древние!
MIC|7|15|Как во дни исхода твоего из земли Египетской, явлю ему дивные дела.
MIC|7|16|Увидят это народы и устыдятся при всем могуществе своем; положат руку на уста, уши их сделаются глухими;
MIC|7|17|будут лизать прах как змея, как черви земные выползут они из укреплений своих; устрашатся Господа Бога нашего и убоятся Тебя.
MIC|7|18|Кто Бог, как Ты, прощающий беззаконие и не вменяющий преступления остатку наследия Твоего? не вечно гневается Он, потому что любит миловать.
MIC|7|19|Он опять умилосердится над нами, изгладит беззакония наши. Ты ввергнешь в пучину морскую все грехи наши.
MIC|7|20|Ты явишь верность Иакову, милость Аврааму, которую с клятвою обещал отцам нашим от дней первых.
