AMOS|1|1|這是 猶大 王 烏西雅 在位與 約阿施 的兒子 以色列 王 耶羅波安 在位的時候，大地震前二年，從 提哥亞 來的牧人 阿摩司 所見的─他的話論到 以色列 。
AMOS|1|2|他說：「耶和華必從 錫安 吼叫， 從 耶路撒冷 出聲； 牧人的草場哀傷， 迦密 的山頂枯乾。」
AMOS|1|3|耶和華如此說： 「 大馬士革 三番四次犯罪， 以鐵的打穀機擊打 基列 ， 我必不撤銷對它的懲罰。
AMOS|1|4|我要降火在 哈薛 的王宮， 吞滅 便‧哈達 的宮殿；
AMOS|1|5|我要折斷 大馬士革 的門閂， 剪除 亞文 平原的居民 和 伯‧伊甸 的掌權者， 亞蘭 人必被擄到 吉珥 。」 這是耶和華說的。
AMOS|1|6|耶和華如此說： 「 迦薩 三番四次犯罪， 擄掠全體百姓交給 以東 ， 我必不撤銷對它的懲罰。
AMOS|1|7|我要降火在 迦薩 城內， 吞滅它的宮殿；
AMOS|1|8|我要剪除 亞實突 的居民 和 亞實基倫 的掌權者， 反手攻擊 以革倫 ， 剩餘的 非利士 人都必滅亡。」 這是主耶和華說的。
AMOS|1|9|耶和華如此說： 「 推羅 三番四次犯罪， 將全體百姓交給 以東 ， 不顧念弟兄的盟約， 我必不撤銷對它的懲罰，
AMOS|1|10|我要降火在 推羅 城內， 吞滅它的宮殿。」
AMOS|1|11|耶和華如此說： 「 以東 三番四次犯罪， 怒氣不停發作，永遠懷著憤怒， 拿刀追趕兄弟，絲毫不存憐憫， 我必不撤銷對它的懲罰。
AMOS|1|12|我要降火在 提幔 ， 吞滅 波斯拉 的宮殿。」
AMOS|1|13|耶和華如此說： 「 亞捫 人三番四次犯罪， 剖開 基列 的孕婦， 擴張自己的疆界， 我必不撤銷對它的懲罰。
AMOS|1|14|我要在戰爭吶喊的日子， 在旋風狂吹時， 在 拉巴 城內放火， 吞滅它的宮殿；
AMOS|1|15|他們的君王和官長必一同被擄。」 這是耶和華說的。
AMOS|2|1|耶和華如此說： 「 摩押 三番四次犯罪， 把 以東 王的骸骨焚燒成灰， 我必不撤銷對它的懲罰。
AMOS|2|2|我要降火在 摩押 ， 吞滅 加略 的宮殿， 摩押 必在鬧鬨、吶喊、吹角聲中滅亡；
AMOS|2|3|我要剪除 摩押 的領袖， 把所有的官長和他一同殺戮。」 這是耶和華說的。
AMOS|2|4|耶和華如此說： 「 猶大 三番四次犯罪， 厭棄耶和華的訓誨， 不遵守他的律例； 他們祖先所隨從虛假的偶像 使他們走迷了， 我必不撤銷對它的懲罰。
AMOS|2|5|我要降火在 猶大 ， 吞滅 耶路撒冷 的宮殿。」
AMOS|2|6|耶和華如此說： 「 以色列 三番四次犯罪， 為銀子賣了義人， 為一雙鞋賣了窮人， 我必不撤銷對它的懲罰。
AMOS|2|7|他們把貧寒人的頭踐踏在地的塵土上 ， 又阻礙困苦人的道路。 父子與同一個女子行淫， 以致褻瀆我的聖名。
AMOS|2|8|他們在各祭壇旁邊， 躺臥在人所典當的衣服上， 又在他們上帝的殿裏 喝受罰之人的酒。
AMOS|2|9|「我從他們面前除滅 亞摩利 人； 他雖高大如香柏樹，強壯如橡樹， 我卻上滅其果，下絕其根。
AMOS|2|10|我曾將你們從 埃及 地領上來， 在曠野裏引導你們四十年， 使你們得 亞摩利 人之地為業；
AMOS|2|11|我從你們子孫中興起先知， 又從你們少年中興起拿細耳人。 以色列 人哪，不是這樣嗎？」 這是耶和華說的。
AMOS|2|12|「你們卻把酒給拿細耳人喝， 囑咐先知說：『不要說預言。』
AMOS|2|13|「看哪，我要把你們壓下去， 如同裝滿禾捆的車壓過一樣。
AMOS|2|14|快跑的無從避難， 壯士無法使力， 勇士也不能自救；
AMOS|2|15|拿弓的站立不住， 腿快的不能逃脫， 騎馬的也不能自救。
AMOS|2|16|到那日，勇士中最有膽量的， 必赤身逃跑。」 這是耶和華說的。
AMOS|3|1|以色列 人哪，當聽耶和華責備你們的話，責備我從 埃及 地領上來的全家，說：
AMOS|3|2|「在地上萬族中，我只認識你們； 因此，我必懲罰你們一切的罪孽。」
AMOS|3|3|二人若不同心， 豈能同行呢？
AMOS|3|4|獅子若無獵物， 豈會在林中咆哮呢？ 少壯獅子若無所得， 豈會從洞裏吼叫呢？
AMOS|3|5|若未設圈套， 雀鳥豈能陷入地上的羅網呢？ 羅網若無所得， 豈會從地上翻起呢？
AMOS|3|6|城中若吹角， 百姓豈不戰兢嗎？ 災禍若臨到一城， 豈非耶和華所降的嗎？
AMOS|3|7|主耶和華不會做任何事情， 除非先將奧祕指示他的僕人眾先知。
AMOS|3|8|獅子吼叫，誰不懼怕呢？ 主耶和華既已說了，誰能不說預言呢？
AMOS|3|9|你們要在 亞實突 的宮殿 和 埃及 地的宮殿傳揚，說： 「要聚集在 撒瑪利亞 的山上， 看城裏有何等大的擾亂與欺壓。」
AMOS|3|10|「他們以暴力搶奪， 堆積在自己的宮殿裏， 卻不懂得行正直的事。」 這是耶和華說的。
AMOS|3|11|所以主耶和華如此說： 「敵人必來圍攻這地， 削弱你的勢力， 搶掠你的宮殿。」
AMOS|3|12|耶和華如此說：「牧人怎樣從獅子口中搶回兩條腿或耳朵的一小片，住 撒瑪利亞 的 以色列 人得救也是如此，不過搶回床的一角和床榻的靠枕 而已。」
AMOS|3|13|主耶和華－萬軍之上帝說： 「當聽這話，警戒 雅各 家。
AMOS|3|14|我懲罰 以色列 罪孽的日子， 也要懲罰 伯特利 的祭壇； 祭壇的角必被砍下，墜落於地。
AMOS|3|15|我要拆毀過冬和避暑的房屋， 象牙的房屋必毀滅， 廣廈豪宅都歸無有。」 這是耶和華說的。
AMOS|4|1|「你們這些 撒瑪利亞山 上的 巴珊 母牛啊， 當聽這話！ 你們欺負貧寒人，壓碎貧窮人， 對主人說：『拿酒來，我們喝吧！』
AMOS|4|2|主耶和華指著自己的神聖起誓說： 『看哪，日子將到，人必用鉤子將你們鉤去， 用魚鉤把你們中最後一個鉤去。
AMOS|4|3|你們必從城牆的缺口 出去， 各人直往前行， 投向 哈門 。』」 這是耶和華說的。
AMOS|4|4|「 以色列 人哪，任你們往 伯特利 去犯罪， 到 吉甲 增加罪過， 每早晨獻上你們的祭物， 每三日納你們的十一奉獻；
AMOS|4|5|任你們獻上有酵的感謝祭， 宣揚你們的甘心祭，使人聽見， 因為這是你們所喜愛的。」 這是主耶和華說的。
AMOS|4|6|「我使你們在每一座城裏牙齒乾淨， 使你們各處的糧食缺乏， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|7|「在收割的前三個月， 我不降雨在你們那裏， 我降雨在這城， 不降雨在那城； 這塊地有雨， 那塊無雨的地就必枯乾。
AMOS|4|8|兩三城的人擠到一個城去找水喝， 卻喝不足， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|9|「我以焚風 和霉爛攻擊你們， 你們許多的菜園、葡萄園、 無花果樹、橄欖樹屢屢被剪蟲 所吃， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|10|「我降瘟疫在你們中間， 如在 埃及 的樣子； 用刀殺戮你們的年輕人 和你們遭擄掠的馬匹， 營中臭氣撲鼻， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|11|「我傾覆你們， 如同上帝從前傾覆 所多瑪 、 蛾摩拉 一樣； 你們好像從火中搶救出來的一根柴， 你們仍不歸向我。」 這是耶和華說的。
AMOS|4|12|「因此， 以色列 啊，我要如此對待你； 因為我要這樣對待你， 以色列 啊， 你當預備迎見你的上帝。」
AMOS|4|13|看哪，那創山，造風，將其心意指示人， 使晨光變幽暗，踩行在地之高處的， 他的名是耶和華－萬軍之上帝。
AMOS|5|1|以色列 家啊，聽我為你們所作的哀歌：
AMOS|5|2|「 以色列 民 跌倒，不得再起； 躺在地上，無人扶起。」
AMOS|5|3|主耶和華如此說： 「 以色列 家的城派出一千，只剩一百； 派出一百，只剩十個。」
AMOS|5|4|耶和華向 以色列 家如此說： 「你們要尋求我，就必存活。
AMOS|5|5|不要往 伯特利 尋求， 不要進入 吉甲 ， 也不要過到 別是巴 ； 因為 吉甲 必被擄走， 伯特利 必歸無有。」
AMOS|5|6|要尋求耶和華，就必存活， 免得他在 約瑟 家如火發出， 焚燒 伯特利 ，無人撲滅。
AMOS|5|7|你們這使公平變為茵蔯， 將公義丟棄於地的人哪！
AMOS|5|8|那造昴星和參星， 使死蔭變為晨光， 使白晝變為黑夜， 召喚海水、 使其傾倒在地面上的， 耶和華是他的名。
AMOS|5|9|他快速摧毀強壯的人， 毀滅就臨到堡壘。
AMOS|5|10|你們怨恨那在城門口斷是非的， 憎惡那說正直話的。
AMOS|5|11|所以，因你們踐踏貧寒人， 向他們勒索糧稅； 你們雖建造石鑿的房屋， 卻不得住在其內； 雖栽植美好的葡萄園， 卻不得喝其中所出的酒。
AMOS|5|12|我知道你們的罪過何其多， 你們的罪惡何其大； 你們迫害義人，收受賄賂， 在城門口屈枉貧窮人。
AMOS|5|13|所以智慧人在這樣的時候必靜默不言， 因為這是險惡的時候。
AMOS|5|14|你們要尋求良善， 不要尋求邪惡，就必存活。 這樣，耶和華－萬軍之上帝 必照你們所說的與你們同在。
AMOS|5|15|要恨惡邪惡，喜愛良善， 在城門口秉公行義； 或者耶和華－萬軍之上帝 會施恩給 約瑟 的餘民。
AMOS|5|16|因此，主耶和華－萬軍之上帝如此說： 「在一切的廣場上必有哀號的聲音； 在各街市上必有人說： 『哀哉！哀哉！』 他們叫農夫來哭號， 叫善唱哀歌的來舉哀；
AMOS|5|17|各葡萄園都有哀號的聲音， 因為我必從你中間經過。」 這是耶和華說的。
AMOS|5|18|想望耶和華日子的人有禍了！ 為甚麼你們要耶和華的日子呢？ 那是黑暗沒有光明的日子，
AMOS|5|19|好像人躲避獅子卻遇見熊； 進房屋以手靠牆，卻被蛇咬。
AMOS|5|20|耶和華的日子豈不是黑暗沒有光明， 幽暗毫無光輝嗎？
AMOS|5|21|「我厭惡你們的節期， 也不喜悅你們的嚴肅會。
AMOS|5|22|你們雖然向我獻燔祭和素祭， 我卻不悅納， 也不看你們用肥畜獻的平安祭。
AMOS|5|23|要使你們歌唱的聲音遠離我， 因為我不聽你們琴瑟的樂曲。
AMOS|5|24|惟願公平如大水滾滾， 公義如江河滔滔。
AMOS|5|25|「 以色列 家啊，你們在曠野四十年，何嘗將祭物和供物獻給我呢？
AMOS|5|26|你們抬著你們的 撒古特 君王 ，和你們為自己所造之偶像 迦溫 ，你們的神明之星。
AMOS|5|27|所以我要把你們擄到 大馬士革 以外。」這是耶和華說的，他的名為萬軍之上帝。
AMOS|6|1|「那在 錫安 安逸， 在 撒瑪利亞山 安穩， 為列國之首，具有名望， 且為 以色列 家所歸向的，有禍了！
AMOS|6|2|你們要過到 甲尼 察看， 從那裏往 哈馬 大城去， 又下到 非利士 人的 迦特 ， 你們比這些國更好嗎？ 或是他們的疆界比你們的疆界廣大呢？
AMOS|6|3|你們以為降禍的日子尚遠， 卻使殘暴的統治 臨近。
AMOS|6|4|「那些躺臥在象牙床上，舒身在榻上的， 吃群中的羔羊和棚裏的牛犢。
AMOS|6|5|他們以琴瑟逍遙歌唱， 為自己作曲 ，像 大衛 一樣；
AMOS|6|6|以大碗喝酒，用上等油抹身， 卻不為 約瑟 所受的苦難憂傷；
AMOS|6|7|所以，現在這些人必首先被擄， 逍遙的歡宴必消失。」
AMOS|6|8|主耶和華指著自己起誓說： 「我憎惡 雅各 的驕傲，厭棄他的宮殿； 我必將城和其中一切所有的都交給敵人。」 這是耶和華－萬軍之上帝說的 。
AMOS|6|9|那時，若一房之內剩下十個人，也都必死。
AMOS|6|10|死人的叔伯要把屍首抬到屋外焚燒，就問房屋內間的人說：「你那裏還有別人嗎？」他說：「沒有。」又說：「不要作聲，不可提耶和華的名。」
AMOS|6|11|看哪，耶和華發命令， 把大房子拆成碎片， 小屋子裂為小塊。
AMOS|6|12|馬豈能在巖石上奔跑？ 人豈能在那裏 用牛耕種呢？ 你們卻使公平變為苦膽， 使公義的果子變為茵蔯。
AMOS|6|13|你們這些喜愛 羅‧底巴 的，自誇說： 「我們不是憑自己的力量攻佔了 加寧 嗎？」
AMOS|6|14|耶和華─萬軍之上帝說： 「 以色列 家，看哪，我必興起一國攻擊你們； 他們必欺壓你們， 從 哈馬口 直到 亞拉巴 的河。」
AMOS|7|1|主耶和華指示我一件事，在春天作物剛長出時，看哪，主 造了蝗蟲；看哪，這是王收割後長出的春天作物。
AMOS|7|2|蝗蟲吃盡那地青草的時候，我說： 「主耶和華啊，求你赦免； 因為 雅各 弱小， 他怎能站立得住呢？」
AMOS|7|3|耶和華對這事改變心意， 耶和華說：「這災可以免了。」
AMOS|7|4|主耶和華又指示我一件事，看哪，主耶和華命火施行審判，火就吞滅深淵，燒盡產業。
AMOS|7|5|我就說： 「主耶和華啊，求你止息； 因為 雅各 弱小， 他怎能站立得住呢？」
AMOS|7|6|耶和華對這事改變心意， 主耶和華說：「這災也可免了。」
AMOS|7|7|他又指示我一件事，看哪，主手拿鉛垂線，站立在依鉛垂線建好的牆邊。
AMOS|7|8|耶和華對我說：「 阿摩司 ，你看見甚麼？」我說：「鉛垂線。」主說： 「看哪，我要在我子民 以色列 中 吊起鉛垂線， 不再寬恕他們。
AMOS|7|9|以撒 的丘壇必荒涼， 以色列 的聖所必荒廢； 我要起來用刀攻擊 耶羅波安 的家。」
AMOS|7|10|伯特利 的祭司 亞瑪謝 派人到 以色列 王 耶羅波安 那裏，說：「 阿摩司 在 以色列 家中圖謀背叛你，他所說的一切話，這地不能承擔；
AMOS|7|11|因為 阿摩司 這樣說： 『 耶羅波安 必被刀殺， 以色列 百姓必被擄， 離開本地。』」
AMOS|7|12|於是 亞瑪謝 對 阿摩司 說：「你這先見哪，要逃到 猶大 地，在那裏過活 ，在那裏說預言；
AMOS|7|13|卻不要在 伯特利 再說預言，因為這裏有王的聖所，有王的宮殿。」
AMOS|7|14|阿摩司 對 亞瑪謝 說：「我原不是先知，也不是先知的門徒；我是牧人，是修剪桑樹的。
AMOS|7|15|耶和華帶領我，叫我不再牧放羊群，對我說：『你去向我子民 以色列 說預言。』
AMOS|7|16|「現在你要聽耶和華的話。 你說：『不要向 以色列 說預言， 也不要向 以撒 家傳講 。』
AMOS|7|17|所以耶和華如此說： 『你的妻子要在城中作妓女， 你的兒女要倒在刀下； 你的地必有人用繩子量了瓜分， 你自己必死在不潔淨之地； 以色列 百姓必被擄， 離開本地。』」
AMOS|8|1|主耶和華又指示我一件事，看哪，有一筐夏天的果子。
AMOS|8|2|他說：「 阿摩司 ，你看見甚麼？」我說：「一筐夏天的果子。」耶和華對我說： 「我子民 以色列 的結局 到了， 我必不再寬恕他們。
AMOS|8|3|那日，宮殿裏的詩歌要變為哀號 ； 必有許多屍首拋在各處， 安靜無聲。」 這是主耶和華說的。
AMOS|8|4|你們這些踐踏貧窮人、 使這地困苦人衰敗的， 當聽這話！
AMOS|8|5|你們說：「初一幾時過去， 我們好賣糧； 安息日幾時過去， 我們好擺開穀物； 我們要把伊法變小， 把舍客勒變大， 以詭詐的天平欺哄人，
AMOS|8|6|用銀子買貧寒人， 以一雙鞋換貧窮人， 把壞的穀物賣給人。」
AMOS|8|7|耶和華指著 雅各 的驕傲起誓說： 「他們這一切的行為，我必永遠不忘。
AMOS|8|8|地豈不因這事震動？ 其中的居民豈不悲哀嗎？ 全地必如 尼羅河 漲起， 如 埃及 的 尼羅河 湧起退落。
AMOS|8|9|「到那日， 我要使太陽在正午落下， 使這地在白晝黑暗。」 這是主耶和華說的。
AMOS|8|10|「我要使你們的節期變為悲哀， 你們一切的歌曲變為哀歌； 我要使眾人腰束麻布， 頭上光禿； 我要使這悲哀如喪獨子， 其結局如悲痛的日子。
AMOS|8|11|「看哪，日子將到， 我必命饑荒降在地上； 人飢餓非因無餅，乾渴非因無水， 而是因不聽耶和華的話。」 這是主耶和華說的。
AMOS|8|12|他們必飄流，從這海到那海， 從北邊到東邊，往來奔跑， 尋求耶和華的話， 卻尋不著。
AMOS|8|13|「當那日，少年和美貌的少女 必因乾渴而發昏。
AMOS|8|14|那些指著 撒瑪利亞 的罪孽 起誓的，說： 『 但 哪，我們指著你那裏的神明起誓』， 又說：『我們指著通往 別是巴 的路起誓』， 這些人都必仆倒，永不再起。」
AMOS|9|1|我看見主站在祭壇旁，說： 「你要擊打柱頂，使門檻震動， 要剪除眾人當中為首的， 他們中最後的 ，我必用刀殺戮； 無一人能逃避，無一人能逃脫。
AMOS|9|2|「雖然他們挖透陰間， 我的手必從那裏拉出他們； 雖然他們爬到天上， 我必從那裏拿下他們；
AMOS|9|3|雖然藏在 迦密山 頂， 我必在那裏搜尋，擒拿他們； 雖然離開我眼前藏在海底， 我必在那裏命令蛇咬他們；
AMOS|9|4|雖然被仇敵擄去， 我也必在那裏命令刀劍殺戮他們； 我必定睛在他們身上， 降禍不降福。」
AMOS|9|5|萬軍的主耶和華觸摸地，地就融化， 凡住在地上的都必悲哀； 全地必如 尼羅河 漲起， 如同 埃及 的 尼羅河 落下。
AMOS|9|6|那在天上建造樓閣、 在地上奠定穹蒼、 召喚海水、 使其傾倒在地面上的， 耶和華是他的名。
AMOS|9|7|耶和華說：「 以色列 人哪， 我豈不是看你們如 古實 人嗎？ 我豈不是領 以色列 人出 埃及 地， 也領 非利士 人出 迦斐託 ， 領 亞蘭 人出 吉珥 嗎？
AMOS|9|8|看哪，主耶和華的眼目 察看這有罪的國度， 要把它從地面上滅絕， 卻不將 雅各 家滅絕淨盡。」 這是耶和華說的。
AMOS|9|9|「看哪，我發命令， 使 以色列 家在萬國中飄流， 好像人用篩子篩穀， 連一粒也不落在地上。
AMOS|9|10|我子民中所有的罪人， 就是那些說 『災禍必不靠近，必不追上我們』的， 都必死在刀下。」
AMOS|9|11|「在那日，我必重建 大衛 倒塌的帳幕， 修補其中的缺口； 我必建立那遭破壞的， 重新修造，如古時一般，
AMOS|9|12|使 以色列 人接管 以東 所剩餘的 和所有稱為我名下的國。 這是耶和華說的，他要行這事。
AMOS|9|13|「看哪，日子將到， 耕種的必接續收割的， 踹葡萄的必接續撒種的； 大山要滴下甜酒， 小山也被漫過。」 這是耶和華說的。
AMOS|9|14|「我要使 以色列 被擄的子民歸回； 他們要重修荒廢的城鎮， 居住在其中； 栽植葡萄園，喝其中所出的酒， 修造果園，吃其中的果子。
AMOS|9|15|我要將他們栽植於本地， 他們必不再從我所賜給他們的地上被拔出。」 這是耶和華－你的上帝說的。
