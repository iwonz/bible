COL|1|1|Paul, an apostle of Christ Jesus by the will of God, and Timothy our brother,
COL|1|2|To the holy and faithful brothers in Christ at Colosse: Grace and peace to you from God our Father.
COL|1|3|We always thank God, the Father of our Lord Jesus Christ, when we pray for you,
COL|1|4|because we have heard of your faith in Christ Jesus and of the love you have for all the saints--
COL|1|5|the faith and love that spring from the hope that is stored up for you in heaven and that you have already heard about in the word of truth, the gospel
COL|1|6|that has come to you. All over the world this gospel is bearing fruit and growing, just as it has been doing among you since the day you heard it and understood God's grace in all its truth.
COL|1|7|You learned it from Epaphras, our dear fellow servant, who is a faithful minister of Christ on our behalf,
COL|1|8|and who also told us of your love in the Spirit.
COL|1|9|For this reason, since the day we heard about you, we have not stopped praying for you and asking God to fill you with the knowledge of his will through all spiritual wisdom and understanding.
COL|1|10|And we pray this in order that you may live a life worthy of the Lord and may please him in every way: bearing fruit in every good work, growing in the knowledge of God,
COL|1|11|being strengthened with all power according to his glorious might so that you may have great endurance and patience, and joyfully
COL|1|12|giving thanks to the Father, who has qualified you to share in the inheritance of the saints in the kingdom of light.
COL|1|13|For he has rescued us from the dominion of darkness and brought us into the kingdom of the Son he loves,
COL|1|14|in whom we have redemption, the forgiveness of sins.
COL|1|15|He is the image of the invisible God, the firstborn over all creation.
COL|1|16|For by him all things were created: things in heaven and on earth, visible and invisible, whether thrones or powers or rulers or authorities; all things were created by him and for him.
COL|1|17|He is before all things, and in him all things hold together.
COL|1|18|And he is the head of the body, the church; he is the beginning and the firstborn from among the dead, so that in everything he might have the supremacy.
COL|1|19|For God was pleased to have all his fullness dwell in him,
COL|1|20|and through him to reconcile to himself all things, whether things on earth or things in heaven, by making peace through his blood, shed on the cross.
COL|1|21|Once you were alienated from God and were enemies in your minds because of your evil behavior.
COL|1|22|But now he has reconciled you by Christ's physical body through death to present you holy in his sight, without blemish and free from accusation--
COL|1|23|if you continue in your faith, established and firm, not moved from the hope held out in the gospel. This is the gospel that you heard and that has been proclaimed to every creature under heaven, and of which I, Paul, have become a servant.
COL|1|24|Now I rejoice in what was suffered for you, and I fill up in my flesh what is still lacking in regard to Christ's afflictions, for the sake of his body, which is the church.
COL|1|25|I have become its servant by the commission God gave me to present to you the word of God in its fullness--
COL|1|26|the mystery that has been kept hidden for ages and generations, but is now disclosed to the saints.
COL|1|27|To them God has chosen to make known among the Gentiles the glorious riches of this mystery, which is Christ in you, the hope of glory.
COL|1|28|We proclaim him, admonishing and teaching everyone with all wisdom, so that we may present everyone perfect in Christ.
COL|1|29|To this end I labor, struggling with all his energy, which so powerfully works in me.
COL|2|1|I want you to know how much I am struggling for you and for those at Laodicea, and for all who have not met me personally.
COL|2|2|My purpose is that they may be encouraged in heart and united in love, so that they may have the full riches of complete understanding, in order that they may know the mystery of God, namely, Christ,
COL|2|3|in whom are hidden all the treasures of wisdom and knowledge.
COL|2|4|I tell you this so that no one may deceive you by fine-sounding arguments.
COL|2|5|For though I am absent from you in body, I am present with you in spirit and delight to see how orderly you are and how firm your faith in Christ is.
COL|2|6|So then, just as you received Christ Jesus as Lord, continue to live in him,
COL|2|7|rooted and built up in him, strengthened in the faith as you were taught, and overflowing with thankfulness.
COL|2|8|See to it that no one takes you captive through hollow and deceptive philosophy, which depends on human tradition and the basic principles of this world rather than on Christ.
COL|2|9|For in Christ all the fullness of the Deity lives in bodily form,
COL|2|10|and you have been given fullness in Christ, who is the head over every power and authority.
COL|2|11|In him you were also circumcised, in the putting off of the sinful nature, not with a circumcision done by the hands of men but with the circumcision done by Christ,
COL|2|12|having been buried with him in baptism and raised with him through your faith in the power of God, who raised him from the dead.
COL|2|13|When you were dead in your sins and in the uncircumcision of your sinful nature, God made you alive with Christ. He forgave us all our sins,
COL|2|14|having canceled the written code, with its regulations, that was against us and that stood opposed to us; he took it away, nailing it to the cross.
COL|2|15|And having disarmed the powers and authorities, he made a public spectacle of them, triumphing over them by the cross.
COL|2|16|Therefore do not let anyone judge you by what you eat or drink, or with regard to a religious festival, a New Moon celebration or a Sabbath day.
COL|2|17|These are a shadow of the things that were to come; the reality, however, is found in Christ.
COL|2|18|Do not let anyone who delights in false humility and the worship of angels disqualify you for the prize. Such a person goes into great detail about what he has seen, and his unspiritual mind puffs him up with idle notions.
COL|2|19|He has lost connection with the Head, from whom the whole body, supported and held together by its ligaments and sinews, grows as God causes it to grow.
COL|2|20|Since you died with Christ to the basic principles of this world, why, as though you still belonged to it, do you submit to its rules:
COL|2|21|"Do not handle! Do not taste! Do not touch!"?
COL|2|22|These are all destined to perish with use, because they are based on human commands and teachings.
COL|2|23|Such regulations indeed have an appearance of wisdom, with their self-imposed worship, their false humility and their harsh treatment of the body, but they lack any value in restraining sensual indulgence.
COL|3|1|Since, then, you have been raised with Christ, set your hearts on things above, where Christ is seated at the right hand of God.
COL|3|2|Set your minds on things above, not on earthly things.
COL|3|3|For you died, and your life is now hidden with Christ in God.
COL|3|4|When Christ, who is your life, appears, then you also will appear with him in glory.
COL|3|5|Put to death, therefore, whatever belongs to your earthly nature: sexual immorality, impurity, lust, evil desires and greed, which is idolatry.
COL|3|6|Because of these, the wrath of God is coming.
COL|3|7|You used to walk in these ways, in the life you once lived.
COL|3|8|But now you must rid yourselves of all such things as these: anger, rage, malice, slander, and filthy language from your lips.
COL|3|9|Do not lie to each other, since you have taken off your old self with its practices
COL|3|10|and have put on the new self, which is being renewed in knowledge in the image of its Creator.
COL|3|11|Here there is no Greek or Jew, circumcised or uncircumcised, barbarian, Scythian, slave or free, but Christ is all, and is in all.
COL|3|12|Therefore, as God's chosen people, holy and dearly loved, clothe yourselves with compassion, kindness, humility, gentleness and patience.
COL|3|13|Bear with each other and forgive whatever grievances you may have against one another. Forgive as the Lord forgave you.
COL|3|14|And over all these virtues put on love, which binds them all together in perfect unity.
COL|3|15|Let the peace of Christ rule in your hearts, since as members of one body you were called to peace. And be thankful.
COL|3|16|Let the word of Christ dwell in you richly as you teach and admonish one another with all wisdom, and as you sing psalms, hymns and spiritual songs with gratitude in your hearts to God.
COL|3|17|And whatever you do, whether in word or deed, do it all in the name of the Lord Jesus, giving thanks to God the Father through him.
COL|3|18|Wives, submit to your husbands, as is fitting in the Lord.
COL|3|19|Husbands, love your wives and do not be harsh with them.
COL|3|20|Children, obey your parents in everything, for this pleases the Lord.
COL|3|21|Fathers, do not embitter your children, or they will become discouraged.
COL|3|22|Slaves, obey your earthly masters in everything; and do it, not only when their eye is on you and to win their favor, but with sincerity of heart and reverence for the Lord.
COL|3|23|Whatever you do, work at it with all your heart, as working for the Lord, not for men,
COL|3|24|since you know that you will receive an inheritance from the Lord as a reward. It is the Lord Christ you are serving.
COL|3|25|Anyone who does wrong will be repaid for his wrong, and there is no favoritism.
COL|4|1|Masters, provide your slaves with what is right and fair, because you know that you also have a Master in heaven.
COL|4|2|Devote yourselves to prayer, being watchful and thankful.
COL|4|3|And pray for us, too, that God may open a door for our message, so that we may proclaim the mystery of Christ, for which I am in chains.
COL|4|4|Pray that I may proclaim it clearly, as I should.
COL|4|5|Be wise in the way you act toward outsiders; make the most of every opportunity.
COL|4|6|Let your conversation be always full of grace, seasoned with salt, so that you may know how to answer everyone.
COL|4|7|Tychicus will tell you all the news about me. He is a dear brother, a faithful minister and fellow servant in the Lord.
COL|4|8|I am sending him to you for the express purpose that you may know about our circumstances and that he may encourage your hearts.
COL|4|9|He is coming with Onesimus, our faithful and dear brother, who is one of you. They will tell you everything that is happening here.
COL|4|10|My fellow prisoner Aristarchus sends you his greetings, as does Mark, the cousin of Barnabas. (You have received instructions about him; if he comes to you, welcome him.)
COL|4|11|Jesus, who is called Justus, also sends greetings. These are the only Jews among my fellow workers for the kingdom of God, and they have proved a comfort to me.
COL|4|12|Epaphras, who is one of you and a servant of Christ Jesus, sends greetings. He is always wrestling in prayer for you, that you may stand firm in all the will of God, mature and fully assured.
COL|4|13|I vouch for him that he is working hard for you and for those at Laodicea and Hierapolis.
COL|4|14|Our dear friend Luke, the doctor, and Demas send greetings.
COL|4|15|Give my greetings to the brothers at Laodicea, and to Nympha and the church in her house.
COL|4|16|After this letter has been read to you, see that it is also read in the church of the Laodiceans and that you in turn read the letter from Laodicea.
COL|4|17|Tell Archippus: "See to it that you complete the work you have received in the Lord."
COL|4|18|I, Paul, write this greeting in my own hand. Remember my chains. Grace be with you.
