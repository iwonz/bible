1COR|1|1|奉上帝旨意，蒙召作基督耶稣使徒的 保罗 ，同弟兄 所提尼 ，
1COR|1|2|写信给在 哥林多 上帝的教会—就是在基督耶稣里成圣、蒙召作圣徒的—以及所有在各处求告我主耶稣基督之名的人。基督是他们的主，也是我们的主。
1COR|1|3|愿恩惠、平安 从我们的父上帝并主耶稣基督归给你们！
1COR|1|4|我常为你们感谢我的上帝，因上帝在基督耶稣里所赐给你们的恩惠。
1COR|1|5|因为你们在他里面凡事富足，具有各种口才、各样知识，
1COR|1|6|正如我为基督作的见证在你们心里得以坚固，
1COR|1|7|以致你们在恩赐上一无欠缺，切切等候我们主耶稣基督的显现。
1COR|1|8|他也必坚固你们到底，使你们在我们主耶稣基督 的日子无可指责。
1COR|1|9|上帝是信实的，他呼召你们好与他儿子—我们的主耶稣基督—共享团契。
1COR|1|10|弟兄们，我藉我们主耶稣基督的名劝你们说话要一致。你们中间不可分裂，只要一心一意彼此团结。
1COR|1|11|我的弟兄们， 革来 氏家里的人曾对我提起你们，说你们中间有纷争。
1COR|1|12|我的意思是，你们各人说：“我是属 保罗 的”；“我是属 亚波罗 的”；“我是属 矶法 的”；“我是属基督的。”
1COR|1|13|基督是分裂的吗？ 保罗 为你们钉了十字架吗？你们是奉 保罗 的名受了洗吗？
1COR|1|14|我感谢上帝 ，除了 基利司布 和 该犹 以外，我没有给你们中的任何一个人施洗，
1COR|1|15|免得有人说你们是奉我的名受洗的。
1COR|1|16|我曾为 司提法那 家施过洗；此外我已记不清有没有给别人施过洗。
1COR|1|17|因为基督差遣我不是为施洗，而是为传福音；并不是用智慧的言论，免得基督的十字架落了空。
1COR|1|18|因为十字架的道理，在那灭亡的人是愚拙，在我们得救的人却是上帝的大能。
1COR|1|19|就如经上所记： “我要摧毁智慧人的智慧， 废弃聪明人的聪明。”
1COR|1|20|智慧人在哪里？文士在哪里？这世上的辩士在哪里？上帝岂不是已使这世上的智慧变成愚拙了吗？
1COR|1|21|既然世人凭自己的智慧不认识上帝，上帝就本着自己的智慧乐意藉着人所传愚拙的话拯救那些信的人。
1COR|1|22|犹太 人要的是神迹， 希腊 人求的是智慧，
1COR|1|23|我们却是传被钉十字架的基督，这对 犹太 人是绊脚石，对外邦人是愚拙；
1COR|1|24|但对那蒙召的，无论是 犹太 人、 希腊 人，基督总是上帝的大能，上帝的智慧。
1COR|1|25|因为，上帝的愚拙总比人智慧；上帝的软弱总比人强壮。
1COR|1|26|弟兄们哪，想一想你们的蒙召，按着人的观点，有智慧的不多，有能力的不多，有尊贵地位的也不多。
1COR|1|27|但是，上帝拣选了世上愚拙的，为了使有智慧的羞愧；又拣选了世上软弱的，为了使强壮的羞愧。
1COR|1|28|上帝也拣选了世上卑贱的，被人厌恶的，以及那一无所有的，为要废掉那样样都有的，
1COR|1|29|使凡血肉之躯的，在上帝面前，一个也不能自夸。
1COR|1|30|但你们得以在基督耶稣里是本乎上帝，他使基督成为我们的智慧，成为公义、圣洁、救赎。
1COR|1|31|如经上所记：“要夸耀的，该夸耀主。”
1COR|2|1|弟兄们，从前我到你们那里去，并没有用高言大智对你们宣讲上帝的奥秘。
1COR|2|2|因为我曾定了主意，在你们中间不知道别的，只知道耶稣基督并他钉十字架。
1COR|2|3|我在你们那里时，又软弱，又惧怕，又战战兢兢。
1COR|2|4|我说的话、讲的道不是用委婉智慧的言语 ，而是以圣灵的大能来证明，
1COR|2|5|为要使你们的信不靠着人的智慧，而是靠着上帝的大能。
1COR|2|6|然而，在成熟的人中，我们也讲智慧，但不是今世的智慧，也不是今世有权有位、将要灭亡的人的智慧。
1COR|2|7|我们讲的是从前隐藏的、上帝奥秘的智慧，就是上帝在万世以前预定使我们得荣耀的智慧；
1COR|2|8|这智慧，今世有权有位的人没有一个知道，若知道，他们就不会把荣耀的主钉在十字架上了。
1COR|2|9|如经上所记： “上帝为爱他的人所预备的 是眼睛未曾看见，耳朵未曾听见， 人心也未曾想到的。”
1COR|2|10|只有上帝藉着圣灵把这事向我们显明了；因为圣灵参透万事，就是上帝深奥的事也参透了。
1COR|2|11|除了在人里头的灵，谁知道人的事？照样，除了上帝的灵，也没有人知道上帝的事。
1COR|2|12|我们所领受的并不是世上的灵，而是从上帝来的灵，为使我们知道上帝把恩赐赏给我们的事。
1COR|2|13|我们也讲说这些事，不是用人的智慧所教的言语，而是用圣灵所教的言语，用属灵的话解释属灵的事 。
1COR|2|14|然而，属血气的人不接受上帝的灵的事，他反倒以这为愚拙，并且他不能了解，因为这些事惟有属灵的人才能领悟。
1COR|2|15|属灵的人能看透万事，却没有一人能看透他。
1COR|2|16|“谁曾知道主的心？ 谁会教导他？” 至于我们，我们有基督的心。
1COR|3|1|弟兄们，我从前对你们说话，还不能把你们当作属灵的，只能把你们当作属肉体的，你们在基督里仅是婴孩。
1COR|3|2|我用奶喂你们，没有用饭喂你们，因为那时你们不能吃。就是如今还是不能，
1COR|3|3|因为你们仍是属肉体的。你们中间有嫉妒、纷争，这岂不是属乎肉体，照着世人的样子生活吗？
1COR|3|4|有人说：“我是属 保罗 的”；有人说：“我是属 亚波罗 的”；这样你们岂不是和世人一样吗？
1COR|3|5|亚波罗 算什么？ 保罗 算什么？我们都是上帝的执事，藉着我们，你们信了；这不过是照着主给各人的恩赐去做罢了。
1COR|3|6|我栽种了， 亚波罗 浇灌了，惟有上帝使它生长。
1COR|3|7|可见，栽种的算不了什么，浇灌的也算不了什么；惟有上帝能使它生长。
1COR|3|8|栽种的和浇灌的都是一样，但将来各人要照自己的劳苦得到自己的报酬。
1COR|3|9|因为我们是上帝的同工，而你们是上帝的田地，上帝的房屋。
1COR|3|10|我照上帝所给我的恩典，好像一个聪明的工头，立好了根基，别人在上面建造；只是各人要谨慎怎样在上面建造。
1COR|3|11|因为，那已经立好的根基就是耶稣基督，此外没有人能立别的根基。
1COR|3|12|若有人用金银、宝石，草木、禾秸，在这根基上建造，
1COR|3|13|各人的工程必将显露，因为那日子要将它显明，有火把它暴露出来，这火要试炼各人的工程怎样。
1COR|3|14|人在那根基上所建造的工程若能保得住，他将要得赏赐。
1COR|3|15|人的工程若被烧了，他将损失，虽然他自己将得救，却要像从火里经过一样。
1COR|3|16|难道不知你们是上帝的殿，上帝的灵住在你们里面吗？
1COR|3|17|若有人毁坏上帝的殿，上帝一定要毁灭那人；因为上帝的殿是神圣的，这殿就是你们。
1COR|3|18|谁都不可自欺。你们中间若有人自以为在今世有智慧，倒不如变为愚拙，好成为有智慧的。
1COR|3|19|因为这世界的智慧在上帝看来是愚拙的。如经上记着： “主使有智慧的人中了自己的诡计；”
1COR|3|20|又说： “主知道智慧人的意念， 因为它们是虚妄的。”
1COR|3|21|所以，无论谁都不可夸耀人；因为万有都是你们的，
1COR|3|22|或 保罗 ，或 亚波罗 ，或 矶法 ，或世界，或生，或死，或现今的事，或将来的事，全是你们的，
1COR|3|23|而你们是属基督的，基督是属上帝的。
1COR|4|1|人应该把我们看为基督的执事，为上帝的奥秘的管家。
1COR|4|2|所求于管家的，是要他忠心。
1COR|4|3|我被你们评断，或被别人评断，我都以为是极小的事；连我自己也不评断自己。
1COR|4|4|虽然我不觉得自己有错，却也不能因此判为无罪；审断我的是主。
1COR|4|5|所以，时候未到，在主来以前什么都不要评断，他要照出暗中的隐情，揭发人的动机。那时，各人要从上帝那里得著称赞。
1COR|4|6|弟兄们，为你们的缘故，我拿这些事应用到我自己和 亚波罗 身上，让你们从我们学到“不可过于圣经所记”这话的意思，免得你们自高自大，看重这个，看轻那个。
1COR|4|7|使你与人不同的是谁呢？你所有的有哪一个不是领受的呢？若是领受的，为何自夸，仿佛不是领受的呢？
1COR|4|8|你们已经饱足了，已经富足了，用不着我们，自己就作王了。我愿意你们果真作王，让我们也可以与你们一同作王！
1COR|4|9|我想，上帝把我们作使徒的明显地列在末后，好像定死罪的囚犯，因为我们成了一台戏，给世界、天使和众人观看。
1COR|4|10|我们为基督的缘故成为愚拙的；你们在基督里倒是聪明的。我们软弱，你们倒强壮；你们有荣耀，我们倒被藐视。
1COR|4|11|直到如今，我们还是又饥又渴，又赤身露体，又挨打，又到处漂泊，
1COR|4|12|并且劳碌，亲手做工；被人咒骂，我们就祝福；被人迫害，我们就忍受；
1COR|4|13|被人毁谤，我们就劝导。直到如今，人还把我们看作世上的污秽，万物中的渣滓。
1COR|4|14|我写这些话，不是要使你们羞愧，而是要警戒你们，好像我所爱的儿女一样。
1COR|4|15|虽然你们在基督里有无数的导师，却没有许多父亲，因我是在基督耶稣里用福音生了你们。
1COR|4|16|所以，我求你们要效法我。
1COR|4|17|因此，我已差 提摩太 到你们那里去。他在主里面是我亲爱和忠心的儿子；他要提醒你们，我在基督耶稣 里怎样行事为人，在各处各教会中怎样教导人。
1COR|4|18|有些人以为我不到你们那里去而自高自大。
1COR|4|19|但是，主若准许，我会很快到你们那里去；我所要知道的，不是那些自高自大者的言语，而是他们的权能。
1COR|4|20|因为上帝的国不在乎言语，而在乎权能。
1COR|4|21|你们愿意怎么样呢？要我带着棍子到你们那里去呢，还是带着慈爱温柔的心呢？
1COR|5|1|我确实听说在你们中间有淫乱的事；这种淫乱连外邦人中也没有，就是有人和他的继母同居。
1COR|5|2|你们还自高自大！你们不是该觉得痛心，把做这事的人从你们中间赶出去吗？
1COR|5|3|我人虽然不在你们那里，心却在你们那里，好像亲自与你们同在。我奉我们主耶稣 的名，已经判断了做这事的人。你们聚会的时候，我的心和你们同在。你们藉着我们主耶稣的权能，
1COR|5|4|
1COR|5|5|要把这样的人交给撒但，使他的肉体败坏，好让他的灵魂在主的日子可以得救。
1COR|5|6|你们这样自夸是不好的。你们不知道一点面酵能使全团发起来吗？
1COR|5|7|既然你们是无酵的面，要把旧酵除净，好使你们成为新团；因为我们逾越节的羔羊—基督已经被杀献为祭牲了。
1COR|5|8|所以，我们来守这节，不可用旧酵，就是不可用恶毒、邪恶的酵，只用纯洁真实的无酵饼。
1COR|5|9|我先前写信告诉过你们，不可与淫乱的人交往。
1COR|5|10|此话不是泛指这世上所有行淫乱的，或贪婪的，勒索的，或拜偶像的；若是这样，你们非离开这世界不可。
1COR|5|11|但现在，我写信告诉你们，若有称为弟兄的人却仍犯淫乱，或贪婪，或拜偶像，或辱骂，或醉酒，或勒索，这样的人不可跟他交往，就是跟他吃饭都不可以。
1COR|5|12|因为审判教外的人与我何干？教内的人岂不是你们要审判吗？
1COR|5|13|至于外人有上帝审判他们。如经上说：“要从你们中间把那邪恶的人赶出去。”
1COR|6|1|你们中间有彼此争吵的事，怎敢告到不义的人面前，而不告到圣徒面前呢？
1COR|6|2|你们岂不知圣徒要审判世界吗？若世界要受你们的审判，难道你们不配审判这最小的事吗？
1COR|6|3|你们岂不知我们要审判天使吗？何况今生的事呢！
1COR|6|4|既是这样，你们若有今生当审判的事，会让教会所轻看的人来审判吗？
1COR|6|5|我说这话是要使你们惭愧。难道你们中间没有一个有智慧的人能审断弟兄中的事吗？
1COR|6|6|你们竟然有弟兄去告弟兄，而且告到不信主的人面前。
1COR|6|7|你们彼此告状，这已经是你们的大错了。为什么不情愿受冤屈呢？为什么不情愿吃亏呢？
1COR|6|8|你们反倒去冤枉人，亏负人，况且所冤枉所亏负的就是弟兄。
1COR|6|9|你们岂不知不义的人不能承受上帝的国吗？不要自欺！无论是淫乱的、拜偶像的、奸淫的、作娼妓 的，亲男色的、
1COR|6|10|偷窃的、贪婪的、醉酒的、辱骂的、勒索的，都不能承受上帝的国。
1COR|6|11|从前你们中间也有人是这样；但现在你们奉主耶稣基督 的名，并藉着我们上帝的灵，已经洗净，已经成圣，已经称义了。
1COR|6|12|“凡事我都可行”，但不是凡事都有益处。“凡事我都可行”，但无论哪一件，我都不受它的辖制。
1COR|6|13|“食物是为肚腹，肚腹是为食物”；但上帝要使这两样都毁坏。身体不是为淫乱，而是为主；主也是为身体。
1COR|6|14|上帝已经使主复活，也要用他自己的能力使我们复活。
1COR|6|15|你们岂不知道你们的身体是基督的肢体吗？我可以把基督的肢体作为娼妓的肢体吗？绝对不可！
1COR|6|16|你们岂不知道与娼妓苟合的，就是与她成为一体吗？因为主说：“二人要成为一体。”
1COR|6|17|但与主联合的，就是与主成为一灵。
1COR|6|18|你们要远避淫行。人所犯的，无论什么罪，都在身体以外；惟有行淫的，是得罪自己的身体。
1COR|6|19|你们岂不知道你们的身体是圣灵的殿吗？这圣灵是从上帝而来，住在你们里面的。而且你们不是属自己的人，
1COR|6|20|因为你们是重价买来的。所以，要在你们的身体上荣耀上帝。
1COR|7|1|关于你们信上所提的事，男人不亲近女人倒好。
1COR|7|2|但为了避免淫乱的事，男人当各有自己的妻子，女人也当各有自己的丈夫。
1COR|7|3|丈夫对妻子要尽本分；妻子对丈夫也要如此。
1COR|7|4|妻子对自己的身体没有主张的权柄，权柄在丈夫；丈夫对自己的身体也没有主张的权柄，权柄在妻子。
1COR|7|5|夫妻不可忽略对方的需求，除非为了要专心祷告，在两相情愿下暂时分房；以后仍要同房，免得撒但趁着你们情不自禁而引诱你们。
1COR|7|6|我说这话是出于容忍，不是命令。
1COR|7|7|我愿众人像我一样；但是各人都有来自上帝的恩赐，一个是这样，一个是那样。
1COR|7|8|我对没有嫁娶的和寡妇说，他们若能维持独身像我一样就好。
1COR|7|9|但他们若不能自制，就应该嫁娶，与其欲火攻心，倒不如结婚为妙。
1COR|7|10|至于那已经嫁娶的，我吩咐他们—其实不是我，而是主吩咐的：妻子不可离开丈夫，
1COR|7|11|若是离开了，不可再嫁，不然要跟丈夫复和；丈夫也不可离弃妻子。
1COR|7|12|我对其余的人说—是我，不是主说—倘若某弟兄有不信的妻子，妻子也情愿和他一起生活，他就不可离弃妻子。
1COR|7|13|妻子有不信的丈夫，丈夫也情愿和她一起生活，她就不可离弃丈夫。
1COR|7|14|因为不信的丈夫会因着妻子成了圣洁；不信的妻子也会因着丈夫 成了圣洁。不然，你们的儿女就不洁净了，但现在他们是圣洁的。
1COR|7|15|倘若那不信的人要离开，就由他离开吧！无论是弟兄是姊妹，遇着这样的事都不必拘束。上帝召你们原是要你们和睦。
1COR|7|16|你这作妻子的怎么知道不能救你的丈夫呢？你这作丈夫的怎么知道不能救你的妻子呢？
1COR|7|17|无论如何，要照主所分给各人的恩赐和上帝所召各人的情况生活。我在各教会里都是这样规定的。
1COR|7|18|有人受割礼后才蒙召，他就不必除去割礼的记号。有人未受割礼前蒙召，他就不必受割礼。
1COR|7|19|受割礼算不了什么，不受割礼也算不了什么，只要谨守上帝的诫命就是了。
1COR|7|20|各人蒙召的时候是什么身份，要守住这身份。
1COR|7|21|你是作奴隶时蒙召的吗？不要介意；若能获得自由，就争取自由更好。
1COR|7|22|因为，蒙主呼召的奴仆是主所释放的人；蒙主呼召的自由之人是基督的奴仆。
1COR|7|23|你们是重价买来的；不要作人的奴仆。
1COR|7|24|弟兄们，你们各人蒙召的时候是什么身份，要在上帝面前守住这身份。
1COR|7|25|关于未婚女子，我没有主的命令，但我既蒙主怜悯、作为一个可信靠的人，把自己的意见告诉你们。
1COR|7|26|因现今的艰难，据我看来，人不如安于现状。
1COR|7|27|你已经有了妻子，就不要求摆脱；你还没有妻子，就不要想娶妻。
1COR|7|28|你若娶妻，并不是犯罪；未婚女子若出嫁，也不是犯罪。然而，这等人会遭受肉身上的苦难，我宁愿你们免受这苦难。
1COR|7|29|弟兄们，我是说：时候不多了。从此以后，那有妻子的，要像没有一样；
1COR|7|30|哀哭的，不像在哀哭；快乐的，不像在快乐；购买的，像一无所得；
1COR|7|31|享受这世界的，不像在享受这世界；因为这世界的局面将要过去了。
1COR|7|32|我愿你们一无挂虑。没有结婚的是为主的事挂虑，想怎样令主喜悦；
1COR|7|33|结了婚的是为世上的事挂虑，想怎样让妻子喜悦，
1COR|7|34|于是，他就分心了。没有结婚的和未婚的女子是为主的事挂虑，为要身体和心灵都圣洁；已经出嫁的是为世上的事挂虑，想怎样让丈夫喜悦。
1COR|7|35|我说这话是为你们的益处，不是要限制你们，而是要你们做合宜的事，得以不分心地对主忠诚。
1COR|7|36|若有人认为自己待他的女儿 不合宜，女儿也过了适婚年龄 ，他可以随意处理，不算有罪，让两人结婚就是了。
1COR|7|37|倘若有人心里坚定，没有不得已的事，并且由得自己作主，心里又决定了不让女儿结婚 ，这样做也好。
1COR|7|38|这样看来，让自己的女儿结婚 固然是好，不让她结婚更好。
1COR|7|39|丈夫活着的时候，妻子是受约束的；丈夫若长眠了，妻子就自由了，可以随意再嫁，只是要嫁给主里面的人。
1COR|7|40|然而，按我的意见，她若能守节就更有福气。我想我自己也有上帝的灵的感动。
1COR|8|1|关于祭过偶像的食物，我们晓得“我们都有知识”，但知识使人自高自大，惟有爱心能造就人。
1COR|8|2|若有人自以为知道什么，他其实仍不知道他所应当知道的。
1COR|8|3|若有人爱上帝，他就是上帝所认识的人了。
1COR|8|4|关于吃祭过偶像的食物，我们知道“偶像在世上算不得什么”；也知道“上帝只有一位，没有别的”。
1COR|8|5|虽然在天上或地上有许多所谓的神明，就如他们中间有许多的神明，许多的主，
1COR|8|6|但是我们只有一位上帝，就是父，万物都出于他，我们也归于他；并只有一位主，就是耶稣基督，万物都是藉着他而有，我们也是藉着他而有。
1COR|8|7|可是，不是人人都有这知识。有人到现在因拜惯了偶像，仍以为所吃的是祭过偶像的食物；既然他们的良心软弱，也就污秽了。
1COR|8|8|其实，食物不能使我们更接近上帝，因为我们不吃也无损，吃也无益。
1COR|8|9|可是，你们要谨慎，免得你们这自由竟成了软弱人的绊脚石。
1COR|8|10|若有人见你这有知识的在偶像的庙里坐席，而这人的良心是软弱的，他岂不放胆去吃那祭过偶像的食物吗？
1COR|8|11|因此，基督为他死的那软弱弟兄，也就因你的知识沉沦了。
1COR|8|12|你们这样得罪弟兄，伤了他们软弱的良心，就是得罪基督。
1COR|8|13|所以，食物若使我的弟兄跌倒，我就永远不吃肉，免得使我的弟兄跌倒了。
1COR|9|1|我不是自由的吗？我不是使徒吗？我不是见过我们的主耶稣吗？你们不是我在主里面工作的成果吗？
1COR|9|2|假若对别人来说，我不是使徒，对你们来说，我总是使徒；因为你们在主里正是我作使徒的印证。
1COR|9|3|对那些质问我的人，这就是我的答辩。
1COR|9|4|难道我们没有权利靠着传福音吃喝吗？
1COR|9|5|难道我们没有权利带着信主的妻子一起出入，如同其余的使徒，和主的兄弟们，和 矶法 一样吗？
1COR|9|6|只有我和 巴拿巴 没有权利不做工吗？
1COR|9|7|有谁当兵而自备粮饷呢？有谁栽葡萄园而不吃园里的果子呢？有谁牧养牛羊而不喝牛羊的奶呢？
1COR|9|8|我说这些话岂是照一般人的看法？律法不也是这样说吗？
1COR|9|9|就如 摩西 的律法记着：“牛在踹谷的时候，不可笼住它的嘴。”难道上帝所挂念的是牛吗？
1COR|9|10|他不全是为我们说的吗？的确是为我们说的！因为耕种的要存着指望去耕种；收割的也要存着分享谷物的指望去收割。
1COR|9|11|我们既然把属灵的种子撒在你们中间，若从你们收取养生之物，这还算大事吗？
1COR|9|12|假如别人在你们身上享有这权利，何况我们呢？ 然而，我们并没有用过这权利，倒是凡事忍受，免得基督的福音受到阻碍。
1COR|9|13|你们岂不知在圣殿供职的人吃圣殿中的食物吗？在祭坛伺候的人分享坛上的供物吗？
1COR|9|14|主也是这样命令，要传福音的人靠着福音养生。
1COR|9|15|但这权利我全然没有用过。我写这些话，并非要你们这样待我，因为我宁可死也不让人使我所夸的落了空。
1COR|9|16|我传福音原没有可夸耀的，因为我是不得已的，若不传福音，我就有祸了。
1COR|9|17|我若甘心做这事，就有赏赐；若不甘心，责任却已经托付给我了。
1COR|9|18|这样，我的赏赐是什么呢？就是我传福音的时候，使人不花钱得福音，免得我用尽了传福音的权利。
1COR|9|19|我虽然是自由的，不受人管辖，但我甘心作了众人的仆人，为赢得更多的人。
1COR|9|20|对 犹太 人，我就作 犹太 人，为要赢得 犹太 人；对律法以下的人，我虽不在律法以下，还是作律法以下的人，为要赢得律法以下的人。
1COR|9|21|对没有律法的人，我就作没有律法的人，为要赢得没有律法的人；其实我在上帝面前，不是没有律法，而是在基督的律法之下。
1COR|9|22|对软弱的人，我就作软弱的人，为要赢得软弱的人。对什么样的人，我就作什么样的人。无论如何我总要救一些人。
1COR|9|23|凡我所做的，都是为福音的缘故，为要与人共享这福音的好处。
1COR|9|24|你们不知道在运动场上赛跑的，大家都跑，但得奖赏的只有一人？你们也要这样跑，好使你们得着奖赏。
1COR|9|25|凡参加竞赛的，在各方面都要有节制，他们不过是要得会朽坏的冠冕；我们却是要得不会朽坏的冠冕。
1COR|9|26|所以，我奔跑，不像无目标的；我斗拳，不像打空气的。
1COR|9|27|我克制己身，使它完全顺服，免得我传福音给别人，自己反而被淘汰了。
1COR|10|1|弟兄们，我不愿意你们不知道，我们的祖宗从前都在云下，都从海中经过，
1COR|10|2|都在云里、海里受洗 归了 摩西 ，
1COR|10|3|并且都吃了一样的灵粮，
1COR|10|4|也都喝了一样的灵水，所喝的是出于跟随着他们的灵磐石；那磐石就是基督。
1COR|10|5|但他们中间多半是上帝不喜欢的人，所以倒毙在旷野里了。
1COR|10|6|这些事都是我们的鉴戒，使我们不要贪恋恶事，像他们贪恋过的一样。
1COR|10|7|也不要拜偶像，像他们中有些人曾经拜过。如经上所记：“百姓坐下吃喝，起来玩乐。”
1COR|10|8|我们也不可犯奸淫，像他们中有些人曾经犯过，一天就倒毙了二万三千人。
1COR|10|9|也不可试探主 ，像他们中有些人曾试探主就被蛇咬死。
1COR|10|10|你们也不可发怨言，像他们中有些人曾经发过，就被毁灭者所灭。
1COR|10|11|这些事发生在他们身上，要作为鉴戒，而且写下来正是要警戒我们这末世的人。
1COR|10|12|所以，自以为站得稳的人必须谨慎，免得跌倒。
1COR|10|13|你们所受的考验无非是人所承受得了的。上帝是信实的，他不会让你们遭受无法承受的考验，在受考验的时候，总会给你们开一条出路，让你们能忍受得了。
1COR|10|14|所以，我亲爱的，你们要远避拜偶像的事。
1COR|10|15|我好像对精明人说的；你们要辨别我的话。
1COR|10|16|我们所祝谢的杯，岂不是同领基督的血吗？我们所擘开的饼，岂不是同领基督的身体吗？
1COR|10|17|因为饼只是一个，我们虽然人多，仍是一体，我们同享一个饼。
1COR|10|18|你们看那按肉体是 以色列 人的，那些吃祭物的人岂不是与祭坛有份吗？
1COR|10|19|那么，我怎么说呢？是说祭偶像之物算得了什么吗？或说偶像算得了什么吗？
1COR|10|20|不，我是说，他们 所献的祭是祭鬼，不是祭上帝；我不愿意你们与鬼来往。
1COR|10|21|你们不能喝主的杯，又喝鬼的杯；不能吃主的筵席，又吃鬼的筵席。
1COR|10|22|我们要惹主的嫉恨吗？我们比他更强吗？
1COR|10|23|“凡事都可行”，但不都有益处。“凡事都可行”，但不都造就人。
1COR|10|24|无论什么人，不要求自己的益处，而要求别人的益处。
1COR|10|25|凡市场上所卖的，你们只管吃，不要为良心的缘故问什么，
1COR|10|26|“因为地和其中所充满的都属于主”。
1COR|10|27|倘若有一个不信的人请你们吃饭，而你们也愿意去，凡摆在你们面前的，只管吃，不要为良心的缘故问什么。
1COR|10|28|若有人对你们说：“这是献过祭的物”，那么为了那告诉你们的人，并为了良心的缘故就不吃。
1COR|10|29|我说的良心不是你自己的，而是他的。我的自由为什么被别人的良心评断呢？
1COR|10|30|我若谢恩而吃，为什么因我谢恩的物被人毁谤呢？
1COR|10|31|所以，你们或吃或喝，无论做什么，都要为荣耀上帝而做。
1COR|10|32|你们不要使 犹太 人、 希腊 人，或上帝教会中的人跌倒；
1COR|10|33|但要像我一样，凡事都使众人喜欢，不求自己的益处，只求众人的益处，使他们得救。
1COR|11|1|你们该效法我，像我效法基督一样。
1COR|11|2|我称赞你们，因为你们凡事记得我，又坚守我所传授给你们的。
1COR|11|3|但是我要你们知道：基督是男人的头；男人是女人的头 ；上帝是基督的头。
1COR|11|4|凡男人祷告或讲道 ，若蒙着头，就是羞辱自己的头。
1COR|11|5|凡女人祷告或讲道，若不蒙着头，就是羞辱自己的头，因为这就如同剃了头发一样。
1COR|11|6|女人若不蒙着头，就该剪了头发；女人若以剪发剃发为羞愧，就该蒙着头。
1COR|11|7|男人本不该蒙着头，因为他是上帝的形像和荣耀；但女人是男人的荣耀。
1COR|11|8|起初，男人不是由女人而出，女人却是由男人而出。
1COR|11|9|而且男人不是为女人造的，女人却是为男人造的。
1COR|11|10|因此，女人为天使的缘故应当在头上有服权柄的记号。
1COR|11|11|然而，照主的安排，女人不可没有男人，男人也不可没有女人。
1COR|11|12|因为女人原是由男人而出，男人是藉着女人而生；但万有都是出于上帝。
1COR|11|13|你们自己要判断，女人祷告上帝，不蒙着头合宜吗？
1COR|11|14|你们的本性不也教导你们，男人若留长头发是他的羞辱吗？
1COR|11|15|但女人留长头发是她的荣耀，因为这头发是给她盖头的 。
1COR|11|16|若有人想要辩驳，我们却没有这样的规矩，上帝的众教会也没有。
1COR|11|17|我现在吩咐你们这话不是在称赞你们，因为你们聚会是有损无益的。
1COR|11|18|首先，我听说你们教会聚会的时候有分裂的事，我也有些相信这话。
1COR|11|19|在你们中间必然有分门结党的事，好使那些经得起考验的人显明出来。
1COR|11|20|你们聚会的时候，不是在吃主的晚餐，
1COR|11|21|因为吃的时候，各人先吃自己的饭，甚至有人饥饿，有人酒醉。
1COR|11|22|难道你们没有家可以吃喝吗？还是你们藐视上帝的教会，使那没有的羞愧呢？我该对你们说什么呢？我要称赞你们吗？在这事上我绝不称赞你们！
1COR|11|23|我当日传给你们的是从主所领受的。主耶稣被出卖的那一夜，拿起饼来，
1COR|11|24|祝谢了，就擘开，说：“这是我的身体，为你们舍 的；你们要如此行，为的是记念我。”
1COR|11|25|饭后，他也照样拿起杯来，说：“这杯是用我的血所立的新约；你们每逢喝的时候，要如此行，来记念我。”
1COR|11|26|你们每逢吃这饼，喝这杯，是宣告主的死，直到他来。
1COR|11|27|所以，任何不按规矩吃了主的饼，喝了主的杯，就是干犯主的身体和主的血了。
1COR|11|28|人应该省察自己，然后吃这饼，喝这杯。
1COR|11|29|因为人吃喝，若不分辨是主的身体，他的吃喝就是定自己的罪了。
1COR|11|30|因此，在你们中间有好些软弱的与患病的，长眠了的也不少。
1COR|11|31|我们若是先省察自己，就不至于受审判。
1COR|11|32|我们受审判的时候，就是被主管教，这样就免得和世人一同被定罪。
1COR|11|33|所以，我的弟兄们，你们聚会吃晚餐的时候，要彼此等待。
1COR|11|34|若有人饿了，要在家里先吃，免得你们聚会，反被定罪。其余的事等我来的时候再安排。
1COR|12|1|弟兄们，关于属灵的恩赐 ，我不愿意你们不明白。
1COR|12|2|你们知道，你们作外邦人的时候，随事被引诱，受了迷惑去拜不会出声的偶像。
1COR|12|3|所以，我要你们知道，被上帝的灵感动的，没有人会说“耶稣该受诅咒”；若不是被圣灵感动的，也没有人能说“耶稣是主”。
1COR|12|4|恩赐有许多种，却是同一位圣灵所赐。
1COR|12|5|事奉有许多种，却是事奉同一位主。
1COR|12|6|工作有许多种，却是同一位上帝在万人中运行万事。
1COR|12|7|圣灵彰显在各人身上，是要使人得益处。
1COR|12|8|有人藉着圣灵领受智慧的言语；有人也靠着同一位圣灵领受知识的言语；
1COR|12|9|又有人由同一位圣灵领受信心；还有人由同一位圣灵领受医病的恩赐；
1COR|12|10|又有人能行异能，又有人能作先知，又有人能辨别诸灵，又有人能说方言 ，又有人能翻方言。
1COR|12|11|这一切都是由惟一的、同一位圣灵所运行，随着自己的旨意分给各人的。
1COR|12|12|就如身体是一个，却有许多肢体，身体的肢体虽多，仍是一个身体；基督也是这样。
1COR|12|13|我们无论是 犹太 人是 希腊 人，是为奴的是自主的，都从一位圣灵受洗成了一个身体，并且共享这位圣灵。
1COR|12|14|身体原不只是一个肢体，而是许多肢体。
1COR|12|15|假如脚说：“我不是手，所以不属于身体”，它不能因此就不属于身体。
1COR|12|16|假如耳朵说：“我不是眼睛，所以不属于身体”，它也不能因此就不属于身体。
1COR|12|17|假如全身是眼睛，听觉在哪里呢？假如全身是耳朵，嗅觉在哪里呢？
1COR|12|18|但现在上帝随自己的意思把肢体一一安置在身体上了。
1COR|12|19|假如全都是一个肢体，身体在哪里呢？
1COR|12|20|但现在肢体虽多，身体还是一个。
1COR|12|21|眼睛不能对手说：“我用不着你。”头也不能对脚说：“我用不着你。”
1COR|12|22|不但如此，身上的肢体，人以为软弱的，更是不可缺少的；
1COR|12|23|身上的肢体，我们认为不体面的，越发给它加上体面；我们不雅观的，越发装饰得雅观。
1COR|12|24|我们雅观的肢体自然用不着装饰；但上帝配搭这身子，把加倍的体面给那有缺欠的肢体，
1COR|12|25|免得身体不协调，总要肢体彼此照顾。
1COR|12|26|假如一个肢体受苦，所有的肢体就一同受苦；假如一个肢体得光荣，所有的肢体就一同快乐。
1COR|12|27|你们是基督的身体，并且各自都是肢体。
1COR|12|28|上帝在教会所设立的：第一是使徒；第二是先知；第三是教师；其次是行异能的；再次是医病的恩赐，帮助人的，治理事的，说方言的。
1COR|12|29|难道个个都是使徒吗？难道个个都是先知吗？难道个个都是教师吗？难道个个都是行异能的吗？
1COR|12|30|难道个个都是有医病的恩赐吗？难道个个都是说方言的吗？难道个个都是翻方言的吗？
1COR|12|31|你们要追求那更大的恩赐。 我现今把最妙的道指示你们。
1COR|13|1|我若能说人间的方言，甚至天使的语言，却没有爱，我就成为鸣的锣、响的钹一般。
1COR|13|2|我若有先知讲道的能力，也明白各样的奥秘，各样的知识，而且有齐备的信心，使我能够移山，却没有爱，我就算不了什么。
1COR|13|3|我若将所有的财产救济穷人，又牺牲自己的身体让人夸赞 ，却没有爱，仍然对我无益。
1COR|13|4|爱是恒久忍耐；又有恩慈；爱是不嫉妒；爱是不自夸，不张狂，
1COR|13|5|不做害羞的事，不求自己的益处，不轻易发怒，不计算人的恶，
1COR|13|6|不喜欢不义，只喜欢真理；
1COR|13|7|凡事包容，凡事相信，凡事盼望，凡事忍耐。
1COR|13|8|爱是永不止息。先知讲道之能终必归于无有；说方言 之能终必停止；知识也终必归于无有。
1COR|13|9|我们现在所知道的有限，先知所讲的也有限，
1COR|13|10|等那完全的来到，这有限的必消逝。
1COR|13|11|我作孩子的时候，说话像孩子，心思像孩子，意念像孩子；既长大成人，就把孩子的事丢弃了。
1COR|13|12|我们现在是对着镜子观看，模糊不清 ；到那时，就要面对面了。我如今所认识的有限，到那时就全认识，如同主认识我一样。
1COR|13|13|如今常存的有信，有望，有爱这三样，其中最大的是爱。
1COR|14|1|你们要追求爱，也要切慕属灵的恩赐，尤其是作先知讲道 。
1COR|14|2|那说方言 的，不是对人说，而是对上帝说，因为没有人听得懂；他是藉着圣灵说各样的奥秘。
1COR|14|3|但作先知讲道的，是对人说，要造就、安慰、劝勉人。
1COR|14|4|说方言的，是造就自己；作先知讲道的，是造就教会。
1COR|14|5|我希望你们都说方言，更希望你们作先知讲道；因为说方言的，若不解释出来，使教会得造就，那作先知讲道的就比他强了。
1COR|14|6|弟兄们，我到你们那里去，若只说方言，不用启示，或知识，或预言，或教导，给你们讲解，我对你们有什么益处呢？
1COR|14|7|就连那有声而没有生命的东西，如箫，如琴，发出来的音若没有分别，怎能知道所吹所弹的是什么呢？
1COR|14|8|号角吹出来的音若不清楚，谁会预备打仗呢？
1COR|14|9|你们也是如此；若用舌头说听不懂的信息，怎能知道所说的是什么呢？你们就是向空气说话了。
1COR|14|10|世上有许多种语言，却没有一样是无意思的。
1COR|14|11|我若不明白那语言的意思，说话的人必以我为未开化的人，我也以他为未开化的人。
1COR|14|12|你们也是如此，既然你们切慕属灵的恩赐，就当追求多得造就教会的恩赐。
1COR|14|13|所以，那说方言的，就当祈求有翻方言的恩赐。
1COR|14|14|我若用方言祷告，是我的灵在祷告；但我的理智没有效果。
1COR|14|15|我应该怎么做呢？我要用灵祷告，也要用理智祷告；我要用灵歌唱，也要用理智歌唱。
1COR|14|16|不然，你用灵祝谢，那在座不通方言的人，既然不明白你的话，怎能在你感谢的时候说“阿们”呢？
1COR|14|17|你的感谢固然是好，不过不能造就别人。
1COR|14|18|我感谢上帝，我说方言比你们众人还多；
1COR|14|19|但在教会中，我宁可用理智说五句教导人的话，强过说万句方言。
1COR|14|20|弟兄们，在心志上不要作小孩子。但是，在恶事上要作婴孩，而在心志上总要作大人。
1COR|14|21|律法上记着：“主说： 我要用外邦人的舌头 和外邦人的嘴唇 向这百姓说话； 虽然如此，他们还是不听从我。”
1COR|14|22|这样看来，说方言不是为信的人作标记，而是为不信的人；作先知讲道不是为不信的人作标记，而是为信的人。
1COR|14|23|所以，全教会聚在一处的时候，若都说方言，偶然有不通方言的或是不信的人进来，岂不会说你们疯了吗？
1COR|14|24|若个个都作先知讲道，偶然有不信的或是不懂方言的人进来，就被众人劝戒，被众人审问，
1COR|14|25|他心里的隐情被显露出来，就必将脸伏地，敬拜上帝，宣告说：“上帝真的是在你们中间了。”
1COR|14|26|弟兄们，那么，你们该怎么做呢？你们聚会的时候，各人或有诗歌，或有教导，或有启示，或有方言，或有翻出来，凡事都应当造就人。
1COR|14|27|若有说方言的，只可有两个人，至多三个人，且要轮流着说，也要有一个人翻出来。
1COR|14|28|若没有人翻，就当在会中闭口，只对自己和上帝说就是了。
1COR|14|29|至于作先知讲道的，只可有两个人或是三个人，其余的人当慎思明辨。
1COR|14|30|假如旁边坐着的得了启示，那先说话的就当闭口不言。
1COR|14|31|因为你们都可以一个一个地作先知讲道，使众人都可以学习，使众人都得劝勉。
1COR|14|32|先知的灵是顺服先知的，
1COR|14|33|因为上帝不是叫人混乱，而是叫人和谐的上帝。 在圣徒的众教会中，
1COR|14|34|妇女应该闭口不言；因为，不准她们说话，总要顺服，正如律法所说的。
1COR|14|35|她们若要学什么，应该在家里问自己的丈夫，因为妇女在会中说话是可耻的。
1COR|14|36|难道上帝的话是从你们出来的吗？难道是单临到你们的吗？
1COR|14|37|若有人自以为是先知，或是属灵的，就应该知道，我所写给你们的是主的命令。
1COR|14|38|若有不理会的，你们也不必理会他。
1COR|14|39|所以，我的弟兄们，你们要切慕作先知讲道的恩赐，不要禁止说方言。
1COR|14|40|凡事都要规规矩矩地按着次序行。
1COR|15|1|弟兄们，我要你们认清我先前传给你们的福音；这福音你们领受了，又靠着它站立得住，
1COR|15|2|你们若能够持守我传给你们的信息，就必因这福音得救，否则你们是徒然相信。
1COR|15|3|我当日所领受又传给你们的，最重要的就是：照圣经所说，基督为我们的罪死了，
1COR|15|4|而且埋葬了；又照圣经所说，第三天复活了，
1COR|15|5|还显给 矶法 看，又显给十二使徒看，
1COR|15|6|后来一次显给五百多弟兄看，其中一大半到现在还在，却也有已经睡了的。
1COR|15|7|以后他显给 雅各 看，再显给众使徒看，
1COR|15|8|最后也显给我看；我如同未到产期而生的人一般。
1COR|15|9|我原是使徒中最小的，不配称为使徒，因为我曾迫害过上帝的教会。
1COR|15|10|然而，由于上帝的恩典，我才成了今日的我，并且他所赐给我的恩典不是徒然的。我比众使徒格外劳苦；其实不是我，而是上帝的恩典与我同在。
1COR|15|11|无论是我或是其他使徒，我们都如此传，你们也都如此信了。
1COR|15|12|既然我们传基督是从死人中复活了，怎么在你们中间有人说没有死人复活的事呢？
1COR|15|13|若没有死人复活的事，基督就没有复活了。
1COR|15|14|基督若没有复活，我们所传的就是枉然，你们所信的也是枉然。
1COR|15|15|这样，我们甚至被当作是为上帝妄作见证的，因为我们见证上帝是使基督复活了。如果死人真的没有复活，上帝就没有使基督复活了。
1COR|15|16|因为死人若不复活，基督也就没有复活了。
1COR|15|17|基督若没有复活，你们的信就是徒然，你们仍活在罪里。
1COR|15|18|就是在基督里睡了的人也灭亡了。
1COR|15|19|我们若靠基督只在今生有指望，就比所有的人更可怜了。
1COR|15|20|其实，基督已经从死人中复活，成为睡了之人初熟的果子。
1COR|15|21|既然死是因一人而来，死人复活也因一人而来。
1COR|15|22|在 亚当 里众人都死了；同样，在基督里众人也都要复活。
1COR|15|23|但各人是按着自己的次序复活：初熟的果子是基督；然后在他来的时候，是那些属于基督的。
1COR|15|24|再后，终结到了，那时基督既将一切执政的、掌权的、有权能的都毁灭了，就把国交给父上帝。
1COR|15|25|因为基督必须掌权，等上帝把一切仇敌都放在他的脚下。
1COR|15|26|他要毁灭的最后仇敌就是死亡。
1COR|15|27|因为经上说：“上帝使万物都服在他的脚下。”既然说万物都服了他，那使万物屈服的，很明显地是不在其内了。
1COR|15|28|既然万物服了他，那时，子也要自己顺服那叫万物服他的，好使上帝在万物之中，在万物之上。
1COR|15|29|不然，那些为死人受洗的，能做什么呢？如果死人不会复活，为什么替他们受洗呢？
1COR|15|30|我们为什么要时刻冒险呢？
1COR|15|31|弟兄们 ，我在我们的主基督耶稣里，指着你们—我所夸的极力地说，我天天冒死。
1COR|15|32|从人的观点看来，我当日在 以弗所 同野兽搏斗，对我有什么益处呢？如果死人没有复活， “让我们吃吃喝喝吧！ 因为明天要死了。”
1COR|15|33|不要被欺骗了； “滥交朋友败坏品德。”
1COR|15|34|你们要醒悟为善，不再犯罪；因为有人不认识上帝。我说这话是要使你们羞愧。
1COR|15|35|但是有人会问：“死人怎样复活呢？他们带着什么身体来呢？”
1COR|15|36|无知的人哪，你所种的若不死就不能生。
1COR|15|37|并且你所种的不是那将来要有的形体，无论是麦子或别样谷物，都不过是子粒。
1COR|15|38|但上帝随自己的意思给它一个形体，并叫各样子粒各有自己的形体。
1COR|15|39|不是所有的肉体都是同样的：人是一个样子，兽又是一个样子，鸟又是一个样子，鱼又是一个样子。
1COR|15|40|有天上的形体，也有地上的形体；但天上形体的荣光是一个样子，地上形体的荣光又是一个样子。
1COR|15|41|日有日的光辉，月有月的光辉，星有星的光辉；这星和那星的光辉也有区别。
1COR|15|42|死人复活也是这样。所种的是会朽坏的，复活的是不朽坏的；
1COR|15|43|所种的是羞辱的，复活的是荣耀的；所种的是软弱的，复活的是强壮的；
1COR|15|44|所种的是血肉的身体，复活的是灵性的身体。既有血肉的身体，也就有灵性的身体。
1COR|15|45|经上也是这样记着说：“首先的人 亚当 成了有生命的人”；末后的 亚当 成了赐生命的灵。
1COR|15|46|但是，不是属灵的在先，而是属血肉的在先，然后才是属灵的。
1COR|15|47|第一个人是出于地，是属于尘土；第二个人是出于天。
1COR|15|48|那属尘土的怎样，凡属尘土的也都怎样；属天的怎样，凡属天的也都怎样。
1COR|15|49|就如我们既有属尘土的形像，将来也必有属天的形像。
1COR|15|50|弟兄们，我要告诉你们的是：血肉之躯不能承受上帝的国，必朽坏的也不能承受不朽坏的。
1COR|15|51|我如今把一件奥秘的事告诉你们：我们不是都要睡觉，而是都要改变，
1COR|15|52|就在一刹那，眨眼之间，号筒末次吹响的时候。因号筒要吹响，死人要复活成为不朽坏的，我们也要改变。
1COR|15|53|这会朽坏的必须变成 不朽坏的；这会死的总要变成不会死的。
1COR|15|54|当这会朽坏的变成不朽坏的，这会死的变成不会死的，那时经上所记“死亡已被胜利吞灭了”的话就应验了。
1COR|15|55|“死亡啊！你得胜的权势在哪里？ 死亡啊！你的毒刺在哪里？”
1COR|15|56|死亡的毒刺就是罪，罪的权势就是律法。
1COR|15|57|感谢上帝，他使我们藉着我们的主耶稣基督得胜。
1COR|15|58|所以，我亲爱的弟兄们，你们务要坚固，不可动摇，常常竭力多做主工，因为你们知道，你们在主里的劳苦不是徒然的。
1COR|16|1|关于为圣徒捐款的事，我从前怎样吩咐 加拉太 的众教会，你们也该怎样做。
1COR|16|2|每逢七日的第一日，每人要照自己的收入抽出若干，保留起来，免得我来的时候现凑。
1COR|16|3|等到我来了，你们写信举荐谁，我就差遣他们，把你们的款项送到 耶路撒冷 去。
1COR|16|4|如果我也该去，他们可以和我同去。
1COR|16|5|我想穿越 马其顿 ；我经过了 马其顿 后，就到你们那里去，
1COR|16|6|可能会和你们同住一些时候，甚至和你们一起过冬。这样无论我往哪里去，你们可以给我送行。
1COR|16|7|我现在不愿意在路过的时候见你们；主若允许，我就指望和你们同住一些时候。
1COR|16|8|不过我要仍旧住在 以弗所 ，直到五旬节，
1COR|16|9|因为有又宽大又有效的门为我开了，虽然反对的人也多。
1COR|16|10|若是 提摩太 来到，你们要留心照顾他，使他在你们那里无所惧怕，因为他做主的工作像我一样。
1COR|16|11|所以，无论谁都不可藐视他。只要送他平安前行，让他到我这里来，因为我等着他和弟兄们同来。
1COR|16|12|至于 亚波罗 弟兄，我再三劝他同弟兄们到你们那里去；但现在他绝不愿意去，等有机会他就会去。
1COR|16|13|你们要警醒，在信仰上要站稳，要勇敢，要刚强。
1COR|16|14|你们所做的一切都要凭爱心而做。
1COR|16|15|弟兄们，你们知道 司提法那 一家，是 亚该亚 初结的果子；他们专以服事圣徒为念。
1COR|16|16|我劝你们顺服这样的人，和一切与他同工同劳的人。
1COR|16|17|司提法那 、 福徒拿都 和 亚该古 到这里来，我很高兴，因为他们补上了你们不在我身边的遗憾。
1COR|16|18|他们使我和你们心里都快慰；这样的人，你们务要敬重。
1COR|16|19|亚细亚 的众教会向你们问安。 亚居拉 、 百基拉 ，和在他们家里的教会，在主里热切地向你们问安。
1COR|16|20|众弟兄都向你们问安。要用圣洁的吻彼此问安。
1COR|16|21|我— 保罗 亲笔问安。
1COR|16|22|若有人不爱主，这人该受诅咒。主啊，愿你来！
1COR|16|23|愿主耶稣基督的恩常与你们众人同在。
1COR|16|24|我在基督耶稣里的爱与你们同在！
