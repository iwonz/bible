1JOHN|1|1|Що було від початку, що ми чули, що бачили власними очима, що розглядали, і чого руки наші торкалися, про Слово життя,
1JOHN|1|2|а життя з'явилось, і ми бачили, і свідчимо, і звіщаємо вам життя вічне, що в Отця перебувало й з'явилося нам,
1JOHN|1|3|що ми бачили й чули про те ми звіщаємо вам, щоб і ви мали спільність із нами. Спільність же наша з Отцем і Сином Його Ісусом Христом.
1JOHN|1|4|А це пишемо вам, щоб повна була ваша радість!
1JOHN|1|5|А це звістка, що ми її чули від Нього і звіщаємо вам: Бог є світло, і немає в Нім жадної темряви!
1JOHN|1|6|Коли ж кажемо, що маємо спільність із Ним, а ходимо в темряві, то неправду говоримо й правди не чинимо!
1JOHN|1|7|Коли ж ходимо в світлі, як Сам Він у світлі, то маємо спільність один із одним, і кров Ісуса Христа, Його Сина, очищує нас від усякого гріха.
1JOHN|1|8|Коли ж кажемо, що не маєм гріха, то себе обманюємо, і немає в нас правди!
1JOHN|1|9|Коли ми свої гріхи визнаємо, то Він вірний та праведний, щоб гріхи нам простити, та очистити нас від неправди всілякої.
1JOHN|1|10|А як кажемо, що ми не згрішили, то чинимо з Нього неправдомовця, і слова Його нема в нас!
1JOHN|2|1|Діточки мої, це пишу я до вас, щоб ви не грішили! А коли хто згрішить, то маємо Заступника перед Отцем, Ісуса Христа, Праведного.
1JOHN|2|2|Він ублагання за наші гріхи, і не тільки за наші, але й за гріхи всього світу.
1JOHN|2|3|А що ми пізнали Його, пізнаємо це з того, коли заповіді Його додержуємо.
1JOHN|2|4|Хто говорить: Пізнав я Його, але не додержує Його заповідів, той неправдомовець, і немає в нім правди!
1JOHN|2|5|А хто додержує Його слово, у тому Божа любов справді вдосконалилась. Із того ми пізнаємо, що в Нім пробуваємо.
1JOHN|2|6|А хто каже, що в Нім пробуває, той повинен поводитись так, як поводився Він.
1JOHN|2|7|Улюблені, не пишу я для вас нову заповідь, але заповідь давню, яку мали від початку: заповідь давня, то слово, що чули його від початку.
1JOHN|2|8|Але нову заповідь я вам пишу, що справді вона в Нім та в вас, що минається темрява, і світло правдиве вже світить.
1JOHN|2|9|Хто говорить, що він пробуває у світлі, та ненавидить брата свого, той у темряві досі.
1JOHN|2|10|А хто любить брата свого, той пробуває у світлі, і в ньому спотикання немає.
1JOHN|2|11|Хто ж ненавидить брата свого, пробуває той у темряві й ходить у темряві, і не знає, куди він іде, бо темрява очі йому осліпила.
1JOHN|2|12|Пишу я вам, дітоньки, що гріхи вам прощаються ради Ймення Його.
1JOHN|2|13|Пишу вам, батьки, бо ви пізнали Того, Хто від початку. Пишу вам, юнаки, бо перемогли ви лукавого.
1JOHN|2|14|Пишу, діти, вам, бо ви пізнали Отця. Я писав вам, батьки, бо ви пізнали Того, Хто від початку. Писав я до вас, юнаки, бо міцні ви, і Слово Боже в вас пробуває, і лукавого перемогли ви.
1JOHN|2|15|Не любіть світу, ані того, що в світі. Коли любить хто світ, у тім немає любови Отцівської,
1JOHN|2|16|бо все, що в світі: пожадливість тілесна, і пожадливість очам, і пиха життєва, це не від Отця, а від світу.
1JOHN|2|17|Минається і світ, і його пожадливість, а хто Божу волю виконує, той повік пробуває!
1JOHN|2|18|Діти остання година! А що чули були, що антихрист іде, а тепер з'явилось багато антихристів, з цього ми пізнаємо, що остання година настала!
1JOHN|2|19|Із нас вони вийшли, та до нас не належали. Коли б були належали до нас, то залишилися б з нами; але вийшли, щоб відкрилось, що не всі вони наші.
1JOHN|2|20|А ви маєте помазання від Святого, і знаєте все.
1JOHN|2|21|Я не писав вам, немов ви не знаєте правди, але що знаєте її, і що всяка лжа не від правди.
1JOHN|2|22|Хто неправдомовець, як не той, хто відкидає, що Ісус є Христос? Це антихрист, що відрікається Отця й Сина!
1JOHN|2|23|Кожен, хто відрікається Сина, не має Отця; хто визнає Сина, той має Отця.
1JOHN|2|24|Тож, що ви чули з початку, нехай в вас пробуває воно; якщо в вас пробуватиме те, що ви чули з початку, то й ви пробуватимете в Сині й Отці.
1JOHN|2|25|А оце та обітниця, яку Він Сам обіцяв нам: вічне життя.
1JOHN|2|26|Це я написав вам про тих, хто обманює вас.
1JOHN|2|27|А помазання, яке прийняли ви від Нього, воно в вас залишається, і ви не потребуєте, щоб вас хто навчав. А що те помазання само вас навчає про все, воно бо правдиве й нехибне, то як вас навчило воно, у тім пробувайте.
1JOHN|2|28|А тепер, діточки, залишайтеся в Нім, щоб, як з'явиться Він, то щоб ми мали відвагу та не були засоромлені Ним під час Його приходу.
1JOHN|2|29|Коли знаєте, що Він праведний, то знайте, що всякий, хто чинить справедливість, народився від Нього.
1JOHN|3|1|Подивіться, яку любов дав нам Отець, щоб ми були дітьми Божими, і ними ми є. Світ нас не знає тому, що Його не пізнав.
1JOHN|3|2|Улюблені, ми тепер Божі діти, але ще не виявилось, що ми будемо. Та знаємо, що, коли з'явиться, то будем подібні до Нього, бо будемо бачити Його, як Він є.
1JOHN|3|3|І кожен, хто має на Нього надію оцю, очищає себе так же само, як чистий і Він.
1JOHN|3|4|Кожен, хто чинить гріх, чинить і беззаконня. Бо гріх то беззаконня.
1JOHN|3|5|І ви знаєте, що Він був з'явився, щоб гріхи наші взяти, а гріха в Нім нема.
1JOHN|3|6|Кожен, хто в Нім пробуває, не грішить; усякий, хто грішить, не бачив Його, і не пізнав Його.
1JOHN|3|7|Діточки, хай ніхто вас не зводить! Хто чинить правду, той праведний, як праведний Він!
1JOHN|3|8|Хто чинить гріх, той від диявола, бо диявол грішить від початку. Тому то з'явився Син Божий, щоб знищити справи диявола.
1JOHN|3|9|Кожен, хто родився від Бога, не чинить гріха, бо в нім пробуває насіння Його. І не може грішити, бо від Бога народжений він.
1JOHN|3|10|Цим пізнаються діти Божі та діти дияволові: Кожен, хто праведности не чинить, той не від Бога, як і той, хто брата свого не любить!
1JOHN|3|11|Бо це та звістка, яку від початку ви чули, щоб любили один одного,
1JOHN|3|12|не так, як той Каїн, що був від лукавого, і брата свого забив. А за що він забив його? Бо лукаві були його вчинки, а брата його праведні.
1JOHN|3|13|Не дивуйтеся, браття мої, коли світ вас ненавидить!
1JOHN|3|14|Ми знаємо, що ми перейшли від смерти в життя, бо любимо братів. А хто брата не любить, пробуває той в смерті.
1JOHN|3|15|Кожен, хто ненавидить брата свого, той душогуб. А ви знаєте, що жаден душогуб не має вічного життя, що в нім перебувало б.
1JOHN|3|16|Ми з того пізнали любов, що душу Свою Він поклав був за нас. І ми мусимо класти душі за братів!
1JOHN|3|17|А хто має достаток на світі, і бачить брата свого в недостачі, та серце своє зачиняє від нього, то як Божа любов пробуває в такому?
1JOHN|3|18|Діточки, любімо не словом, ані язиком, але ділом та правдою!
1JOHN|3|19|Із цього довідуємось, що ми з правди, і впокорюєм наші серця перед Ним,
1JOHN|3|20|бо коли винуватить нас серце, то Бог більший від нашого серця та відає все!
1JOHN|3|21|Улюблені, коли не винуватить нас серце, то маємо відвагу до Бога,
1JOHN|3|22|і чого тільки попросимо, одержимо від Нього, бо виконуємо Його заповіді та чинимо любе для Нього.
1JOHN|3|23|І оце Його заповідь, щоб ми вірували в Ім'я Сина Його Ісуса Христа, і щоб любили один одного, як Він нам заповідь дав!
1JOHN|3|24|А хто Його заповіді береже, той у Нім пробуває, а Він у ньому. А що в нас пробуває, пізнаємо це з того Духа, що Він нам Його дав.
1JOHN|4|1|Улюблені, не кожному духові вірте, але випробовуйте духів, чи від Бога вони, бо неправдивих пророків багато з'явилося в світ.
1JOHN|4|2|Духа Божого цим пізнавайте: кожен дух, який визнає, що Ісус Христос прийшов був у тілі, той від Бога.
1JOHN|4|3|А кожен дух, який не визнає Ісуса, той не від Бога, але він антихристів, про якого ви чули, що йде, а тепер уже він у світі.
1JOHN|4|4|Ви від Бога, дітки, і ви перемогли їх, більший бо Той, Хто в вас, аніж той, хто в світі.
1JOHN|4|5|Вони від світу, тому то говорять від світу, а світ слухає їх.
1JOHN|4|6|Ми від Бога, хто знає Бога, той слухає нас, хто не від Бога, той не слухає нас. Цим пізнаємо Духа правди та духа обмани.
1JOHN|4|7|Улюблені, любім один одного, бо від Бога любов, і кожен, хто любить, родився від Бога та відає Бога!
1JOHN|4|8|Хто не любить, той Бога не пізнав, бо Бог є любов!
1JOHN|4|9|Любов Божа до нас з'явилася тим, що Бог Сина Свого Однородженого послав у світ, щоб ми через Нього жили.
1JOHN|4|10|Не в тому любов, що ми полюбили Бога, а що Він полюбив нас, і послав Свого Сина вблаганням за наші гріхи.
1JOHN|4|11|Улюблені, коли Бог полюбив нас отак, то повинні любити і ми один одного!
1JOHN|4|12|Бога не бачив ніколи ніхто. Коли один одного любимо, то Бог в нас пробуває, а любов Його в нас удосконалилась.
1JOHN|4|13|Що ми пробуваємо в Ньому, а Він у нас, пізнаємо це тим, що Він дав нам від Духа Свого.
1JOHN|4|14|І ми бачили й свідчимо, що Отець послав Сина Спасителем світу.
1JOHN|4|15|Коли хто визнає, що Ісус то Син Божий, то в нім Бог пробуває, а він у Бозі.
1JOHN|4|16|Ми познали й увірували в ту любов, що Бог її має до нас. Бог є любов, і хто пробуває в любові, пробуває той в Бозі, і в нім Бог пробуває!
1JOHN|4|17|Любов удосконалюється з нами так, що ми маємо відвагу на день судний, бо який Він, такі й ми на цім світі.
1JOHN|4|18|Страху немає в любові, але досконала любов проганяє страх геть, бо страх має муку. Хто ж боїться, той не досконалий в любові.
1JOHN|4|19|Ми любимо Його, бо Він перше нас полюбив.
1JOHN|4|20|Як хто скаже: Я Бога люблю, та ненавидить брата свого, той неправдомовець. Бо хто не любить брата свого, якого бачить, як може він Бога любити, Якого не бачить?
1JOHN|4|21|І ми оцю заповідь маємо від Нього, щоб, хто любить Бога, той і брата свого любив!
1JOHN|5|1|Кожен, хто вірує, що Ісус то Христос, той родився від Бога. І кожен, хто любить Того, Хто породив, любить і Того, Хто народився від Нього.
1JOHN|5|2|Що ми любимо Божих дітей, дізнаємося з того, коли любимо Бога і Його заповіді додержуємо.
1JOHN|5|3|Бо то любов Божа, щоб ми додержували Його заповіді, Його ж заповіді не тяжкі.
1JOHN|5|4|Бо кожен, хто родився від Бога, перемагає світ. А оце перемога, що світ перемогла, віра наша.
1JOHN|5|5|А хто світ перемагає, як не той, хто вірує, що Ісус то Син Божий?
1JOHN|5|6|То Той, що прийшов був водою та кров'ю, Ісус Христос. І не тільки водою, а водою та кров'ю. І Дух свідчить, бо Дух то правда.
1JOHN|5|7|Бо троє свідкують на небі: Отець, Слово й Святий Дух, і ці Троє Одно.
1JOHN|5|8|І троє свідкують на землі: дух, і вода, і кров, і троє в одно.
1JOHN|5|9|Коли ми приймаємо свідчення людське, то свідчення Боже вартніше, бо це свідчення Бога, яким свідчив про Сина Свого.
1JOHN|5|10|Хто вірує в Божого Сина, той свідчення має в собі. Хто не вірує Богові, той учинив Його неправдомовцем, бо не вірив у свідчення, яким Бог свідчив про Сина Свого.
1JOHN|5|11|А це свідчення, що Бог життя вічне нам дав, а життя це у Сині Його.
1JOHN|5|12|Хто має Сина, той має життя; хто не має Сина Божого, той не має життя.
1JOHN|5|13|Оце написав я до вас, що віруєте в Ім'я Божого Сина, щоб ви знали, що ви віруючи в Ім'я Божого Сина, маєте вічне життя.
1JOHN|5|14|І оце та відвага, що ми маємо до Нього, що коли чого просимо згідно волі Його, то Він слухає нас.
1JOHN|5|15|А як знаємо, що Він слухає нас, чого тільки ми просимо, то знаємо, що одержуємо те, чого просимо від Нього.
1JOHN|5|16|Коли хто бачить брата свого, що грішить гріхом не на смерть, нехай молиться за нього, і Він життя йому дасть, тим, хто грішить не на смерть. Є й гріх на смерть, не про нього кажу, щоб молився.
1JOHN|5|17|Усяка неправда то гріх. Та є гріх не на смерть.
1JOHN|5|18|Ми знаємо, що кожен, хто народився від Бога, не грішить, бо хто народився від Бога, той себе береже, і лукавий його не торкається.
1JOHN|5|19|Ми знаємо, що ми від Бога, і що ввесь світ лежить у злі.
1JOHN|5|20|Ми знаємо, що Син Божий прийшов, і розум нам дав, щоб пізнати Правдивого, і щоб бути в правдивому Сині Його, Ісусі Христі. Він Бог правдивий і вічне життя!
1JOHN|5|21|Дітоньки, бережіться від ідолів! Амінь.
