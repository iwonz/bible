JOB|1|1|乌斯 地有一个人名叫 约伯 。这人完全、正直、敬畏上帝、远离恶事。
JOB|1|2|他生了七个儿子，三个女儿。
JOB|1|3|他的家产有七千只羊，三千匹骆驼，五百对牛，五百匹母驴，并有许多仆婢。这人在东方人中为至大。
JOB|1|4|他的儿子按着日子各在自己家里摆设宴席，派人去请他们的三个姊妹来，与他们一同吃喝。
JOB|1|5|宴席的日子过了， 约伯 派人去叫他们自洁。他清早起来，按着他们众人的数目献燔祭，因为他说：“恐怕我的儿子犯了罪，心中背弃 上帝。” 约伯 常常这样行。
JOB|1|6|有一天，上帝的众使者 来侍立在耶和华面前，撒但也来在其中。
JOB|1|7|耶和华对撒但说：“你从哪里来？”撒但回答耶和华说：“我从地上走来走去，在那里往返。”
JOB|1|8|耶和华对撒但说：“你曾用心察看我的仆人 约伯 没有？地上再没有人像他那样完全、正直、敬畏上帝、远离恶事。”
JOB|1|9|撒但回答耶和华说：“ 约伯 敬畏上帝，岂是无故呢？
JOB|1|10|你岂不是四面圈上篱笆围护他和他的家，以及他一切所有的吗？他手所做的都蒙你赐福，他的家产也在地上增多。
JOB|1|11|但你若伸手毁他一切所有的，他必当面背弃你。”
JOB|1|12|耶和华对撒但说：“看哪，凡他所有的都在你手中；只是不可伸手加害于他。”于是撒但从耶和华面前退出去。
JOB|1|13|有一天， 约伯 的儿女正在他们长兄的家里吃饭喝酒，
JOB|1|14|有报信的来见 约伯 ，说：“牛正耕地，母驴在旁边吃草，
JOB|1|15|示巴 人忽然闯来，把牲畜掳去，并用刀杀了仆人；惟有我一人逃脱，来报信给你。”
JOB|1|16|他还说话的时候，又有人来说：“上帝从天上降下火来，把羊群和仆人都吞灭了；惟有我一人逃脱，来报信给你。”
JOB|1|17|他还说话的时候，又有人来说：“ 迦勒底 人分成三队忽然闯来，把骆驼掳去，并用刀杀了仆人；惟有我一人逃脱，来报信给你。”
JOB|1|18|他还说话的时候，又有人来说：“你的儿女正在他们长兄的家里吃饭喝酒，
JOB|1|19|看哪，有狂风从旷野刮来，袭击房屋的四角，房屋倒塌在年轻人身上，他们就都死了；惟有我一人逃脱，来报信给你。”
JOB|1|20|约伯 就起来，撕裂外袍，剃了头，俯伏在地敬拜，
JOB|1|21|说：“我赤身出于母胎，也必赤身归回；赏赐的是耶和华，收取的也是耶和华。耶和华的名是应当称颂的。”
JOB|1|22|在这一切的事上， 约伯 并没有犯罪，也不以上帝为狂妄。
JOB|2|1|又有一天，上帝的众使者 来侍立在耶和华面前，撒但也来在其中。
JOB|2|2|耶和华问撒但说：“你从哪里来？”撒但回答说：“我从地上走来走去，在那里往返。”
JOB|2|3|耶和华对撒但说：“你曾用心察看我的仆人 约伯 没有？地上再没有人像他那样完全、正直、敬畏上帝、远离恶事。你虽激起我攻击他，无故吞灭他，他仍然持守他的纯正。”
JOB|2|4|撒但回答耶和华说：“人以皮代皮，情愿舍去一切所有的，来保全性命。
JOB|2|5|但你若伸手伤他的骨头和他的肉，他必当面背弃 你。”
JOB|2|6|耶和华对撒但说：“看哪，他在你手中，只要留下他的性命。”
JOB|2|7|于是撒但从耶和华面前退出去，击打 约伯 ，使他从脚掌到头顶长毒疮。
JOB|2|8|约伯 就坐在灰烬中，拿瓦片刮身体。
JOB|2|9|他的妻子对他说：“你仍然持守你的纯正吗？你背弃上帝，死了吧！”
JOB|2|10|约伯 却对她说：“你说话，正如愚顽的妇人。唉！难道我们从上帝手里得福，不也受祸吗？”在这一切的事上， 约伯 并没有以口犯罪。
JOB|2|11|约伯 的三个朋友， 提幔 人 以利法 、 书亚 人 比勒达 、 拿玛 人 琐法 ，听说这一切的灾祸临到他身上，各人就从自己的地方相约同来，为他悲伤，安慰他。
JOB|2|12|他们远远地举目观看，认不出他来，就放声大哭。各人撕裂外袍，向空中撒尘土，落在自己的头上。
JOB|2|13|他们同他七天七夜坐在地上，一句话也不对他说，因为他们见到了极大的痛苦。
JOB|3|1|此后， 约伯 开口诅咒自己的生日 。
JOB|3|2|约伯 说：
JOB|3|3|“愿我生的那日灭没， 说‘怀了男胎’的那夜也灭没。
JOB|3|4|愿那日变为黑暗， 愿上帝不从上面寻找它， 愿亮光不照于其上。
JOB|3|5|愿黑暗和死荫索取那日， 愿密云停在其上， 愿白天的昏暗 恐吓它。
JOB|3|6|愿那夜被幽暗夺取， 不在一年的日子中喜乐， 也不列入月中的数目。
JOB|3|7|看哪，愿那夜没有生育， 其间也没有欢乐的声音。
JOB|3|8|愿那些诅咒日子且能惹动 力威亚探 的， 诅咒那夜。
JOB|3|9|愿那夜黎明的星宿变为黑暗， 盼亮却不亮， 也不见晨曦破晓 ；
JOB|3|10|因它没有把怀我胎的门关闭， 也没有从我的眼中隐藏患难。
JOB|3|11|“我为何不出母胎而死？ 为何不出母腹就气绝呢？
JOB|3|12|为何有膝盖接收我？ 为何有奶哺养我呢？
JOB|3|13|不然，我现在已躺卧安睡， 而且，早已长眠安息；
JOB|3|14|与那些为自己重建荒凉之处， 地上的君王和谋士在一起；
JOB|3|15|或与把银子装满房屋， 拥有金子的王子在一起；
JOB|3|16|我为何不像流产的胎儿被埋藏， 如同未见光的婴孩？
JOB|3|17|在那里恶人止息搅扰， 在那里困乏人得享安息，
JOB|3|18|被囚的人同得安逸， 不再听见监工的声音。
JOB|3|19|大的小的都在那里， 奴仆脱离主人得自由。
JOB|3|20|“遭受患难的人为何有光赐给他呢？ 心中愁苦的人为何有生命赐给他呢？
JOB|3|21|他们等死，却不得死； 求死，胜于求隐藏的珍宝。
JOB|3|22|他们寻见坟墓， 就欢喜快乐，极其高兴。
JOB|3|23|这人的道路遮隐， 上帝又四面围困他。
JOB|3|24|我吃饭前就发出叹息， 我的唉哼涌出如水。
JOB|3|25|因我所恐惧的临到我， 我所惧怕的迎向我；
JOB|3|26|我不得安逸，不得平静， 也不得安息，却有患难来到。”
JOB|4|1|提幔 人 以利法 回答说：
JOB|4|2|“人想与你说话，你就厌烦吗？ 但谁能忍住不发言呢？
JOB|4|3|看哪，你素来教导许多人， 又坚固软弱的手。
JOB|4|4|你的言语曾扶助跌倒的人； 你使软弱的膝盖稳固。
JOB|4|5|但现在祸患临到 你，你就烦躁了； 它挨近你，你就惊惶。
JOB|4|6|你的倚靠不是在于你敬畏上帝吗？ 你的盼望不是在于你行事纯正吗？
JOB|4|7|“请你追想：无辜的人有谁灭亡？ 正直的人何处被剪除？
JOB|4|8|按我所见，耕罪孽的， 种毒害的，照样收割。
JOB|4|9|上帝一嘘气，他们就灭亡； 上帝一发怒，他们就消失。
JOB|4|10|狮子吼叫，猛狮咆哮， 少壮狮子的牙齿被敲断。
JOB|4|11|公狮因缺猎物而死， 母狮的幼狮都离散。
JOB|4|12|“有话暗中传递给我， 耳朵听其微小的声音。
JOB|4|13|世人沉睡的时候， 从夜间异象的杂念中，
JOB|4|14|恐惧战兢临到我身， 使我百骨战抖。
JOB|4|15|有灵从我面前经过， 我身上的毫毛竖立。
JOB|4|16|那灵停住， 我却不能辨其形状； 有形像在我眼前。 我在静默中听见有声音：
JOB|4|17|‘必死的人能比上帝公义吗？ 壮士能比造他的主纯洁吗？
JOB|4|18|看哪，主不信靠他的仆人， 尚且指他的使者为愚昧，
JOB|4|19|何况那些住在泥屋、 根基在尘土里、 被蛀虫所毁坏的人呢？
JOB|4|20|早晚之间，他们就被毁灭， 永归无有，无人理会。
JOB|4|21|他们帐棚的绳索岂不从中拔出来呢？ 他们死，且是无智慧而死。’”
JOB|5|1|“你呼求吧，有谁回答你呢？ 圣者之中，你转向哪一位呢？
JOB|5|2|愤怒害死愚妄人， 嫉妒杀死愚蠢的人。
JOB|5|3|我曾见愚妄人扎下根， 但我忽然诅咒他的住处。
JOB|5|4|他的儿女远离稳妥之地， 在城门口被欺压，无人搭救。
JOB|5|5|他的庄稼被饥饿的人吃尽了， 就是在荆棘里的也抢去了； 他的财宝被陷阱 张口吞没了。
JOB|5|6|因为祸患不是从尘土中出来， 患难也不是从土地里长出。
JOB|5|7|人生出来必遭遇患难， 如同火花 飞腾。
JOB|5|8|“至于我，我必寻求上帝， 把我的事情交托给他。
JOB|5|9|他行大事不可测度， 行奇事不可胜数。
JOB|5|10|他降雨在地面， 赐水于田野。
JOB|5|11|他将卑微的人安置在高处， 将哀痛的人举到稳妥之地。
JOB|5|12|他破坏通达人的计谋， 使他们手所做的不得成就。
JOB|5|13|他使有智慧的人中了自己的诡计， 叫狡诈人的计谋速速落空。
JOB|5|14|他们白昼遇见黑暗， 午间摸索如在夜间。
JOB|5|15|上帝拯救贫穷人脱离残暴人的手， 脱离他们口中的刀。
JOB|5|16|这样，贫寒人有指望， 不义的人闭口无言。
JOB|5|17|“看哪，上帝所惩治的人是有福的！ 所以你不可轻看全能者的管教。
JOB|5|18|因为他打伤，又包扎； 他击伤，又亲手医治。
JOB|5|19|你六次遭难，他必救你； 就是七次，灾祸也无法害你。
JOB|5|20|在饥荒中，他必救你脱离死亡； 在战争中，他必救你脱离刀剑的权势。
JOB|5|21|你必被隐藏，不受口舌之害； 灾害临到，你也不惧怕。
JOB|5|22|对于灾害饥馑，你必讥笑； 至于地上的野兽，你也不惧怕。
JOB|5|23|因为你必与田间的石头立约， 田里的野兽也必与你和好。
JOB|5|24|你必知道你的帐棚平安， 你查看你的羊圈，一无所失。
JOB|5|25|你也必知道你的后裔众多， 你的子孙像地上的青草。
JOB|5|26|你必寿高年迈才归坟墓， 好像禾捆按时收藏。
JOB|5|27|看哪，这道理我们已经考察，本是如此。 你须要听，要亲自明白。”
JOB|6|1|约伯 回答说：
JOB|6|2|“惟愿我的烦恼被秤一秤， 我一切的灾害放在天平里，
JOB|6|3|现今都比海沙更重， 所以我说话急躁。
JOB|6|4|因全能者的箭射中了我， 我的灵喝尽其毒； 上帝的惊吓摆阵攻击我。
JOB|6|5|野驴有草岂会叫唤？ 牛有饲料岂会吼叫？
JOB|6|6|食物淡而无盐岂可吃呢？ 蛋白有什么滋味呢？
JOB|6|7|那些可厌的食物， 我心不肯挨近。
JOB|6|8|“惟愿我得着所求的， 上帝赏赐我所切望的，
JOB|6|9|愿上帝把我压碎， 伸手将我剪除。
JOB|6|10|我因没有违弃那圣者的言语， 就仍以此为安慰， 在不止息的痛苦中还可欢跃。
JOB|6|11|我有什么气力使我等候？ 我有什么结局使我忍耐？
JOB|6|12|我的气力岂是石头的气力？ 我的肉身岂是铜呢？
JOB|6|13|在我里面岂不是无助吗？ 智慧岂不是从我心中被赶逐吗？
JOB|6|14|“灰心的人，他的朋友当以慈爱待他， 因为他将离弃敬畏全能者的心。
JOB|6|15|我的弟兄诡诈，好像河道， 像溪水流过的河床，
JOB|6|16|因结冰而混浊， 有雪藏在其中，
JOB|6|17|暖和的时候就溶化， 炎热时便从原处干涸。
JOB|6|18|商队偏离道路， 上到荒凉之地而死亡。
JOB|6|19|提玛 的商队瞻望， 示巴 的旅客等候。
JOB|6|20|他们因希望落空就抱愧， 来到那里便蒙羞。
JOB|6|21|现在你们正是这样 ， 看见惊吓的事就惧怕。
JOB|6|22|我岂说：‘请你们供给我， 从你们的财物中送礼给我’？
JOB|6|23|或说：‘请你们拯救我脱离敌人的手， 救赎我脱离残暴人的手’吗？
JOB|6|24|“请你们指教我，我就不作声； 我在何事上有错，请使我明白。
JOB|6|25|正直言语的力量何其大！ 但你们责备是责备什么呢？
JOB|6|26|绝望人的讲论既然如风， 你们还计划批驳言语吗？
JOB|6|27|你们甚至为孤儿抽签， 把朋友当货物。
JOB|6|28|“现在，请你们看着我， 我绝不当面说谎。
JOB|6|29|请你们转意，不要不公义； 请再转意，正义在我这里。
JOB|6|30|我的舌头岂有不公义吗？ 我的上膛岂不辨奸恶吗？”
JOB|7|1|“人在世上岂无劳役呢？ 他的日子不像雇工的日子吗？
JOB|7|2|像奴仆切慕阴凉， 像雇工等待工钱，
JOB|7|3|我也照样度过虚空的岁月， 愁烦的夜晚指定给我。
JOB|7|4|我躺卧的时候就说： ‘我何时可以起来呢？’漫漫长夜， 我总是翻来覆去，直到天亮。
JOB|7|5|我的肉体以虫子和尘土为衣， 我的皮肤才收了口又流脓。
JOB|7|6|我的日子比织布的梭更快， 都消耗在没有指望之中。
JOB|7|7|“你要记得，我的生命不过是一口气， 我的眼睛必不再看见福乐。
JOB|7|8|观看我的人，他的眼必不看见我； 你的眼目投向我，我却不在了。
JOB|7|9|云彩消散而去； 照样，人下阴间也不再上来。
JOB|7|10|他不再回自己的家， 他自己的地方也不再认得他。
JOB|7|11|“我甚至不封我的口； 我灵愁苦，要发出言语； 我心苦恼，要吐露哀情。
JOB|7|12|我岂是海洋，岂是大鱼， 你竟防守着我呢？
JOB|7|13|我若说：‘我的床必安慰我， 我的榻必分担我的苦情’，
JOB|7|14|你就用梦惊扰我， 用异象恐吓我。
JOB|7|15|甚至我宁可窒息死亡， 胜似留我这副骨头。
JOB|7|16|我厌弃生命，不愿永远活着。 你任凭我吧，因我的日子都是虚空。
JOB|7|17|人算什么，你竟看他为大， 将他放在心上，
JOB|7|18|每早晨鉴察他， 每时刻考验他？
JOB|7|19|你到何时才转眼不看我， 任凭我咽下唾沫呢？
JOB|7|20|鉴察人的主啊，我若有罪，于你何妨？ 为何以我当你的箭靶， 使我成为你的重担呢？
JOB|7|21|为何不赦免我的过犯， 除掉我的罪孽呢？ 我现今要躺卧在尘土中； 你要切切寻找我，我却不在了。”
JOB|8|1|书亚 人 比勒达 回答说：
JOB|8|2|“这些话你要说到几时？ 你口中的言语如狂风要到几时呢？
JOB|8|3|上帝岂能偏离公平？ 全能者岂能偏离公义？
JOB|8|4|或者你的儿女得罪了他， 他就把他们交在过犯的掌控中。
JOB|8|5|你若切切寻求上帝， 向全能者恳求；
JOB|8|6|你若纯洁正直， 他必定为你兴起， 使你公义的居所兴旺。
JOB|8|7|你起初虽然微小， 日后必非常强盛。
JOB|8|8|“请你询问上代， 思念他们祖先所查究的。
JOB|8|9|我们不过从昨日才有，一无所知， 因我们在世的日子好像影子。
JOB|8|10|他们岂不指教你，告诉你， 说出发自内心的言语呢？
JOB|8|11|“蒲草没有泥岂能生长？ 芦荻没有水岂能长大？
JOB|8|12|它还青翠，没有割下的时候， 比百样的草先枯槁。
JOB|8|13|凡忘记上帝的人，路途也是这样； 不虔敬人的指望要灭没。
JOB|8|14|他所仰赖的必折断， 他所倚靠的是蜘蛛网。
JOB|8|15|他要倚靠房屋，房屋却站立不住； 他要抓住房屋，房屋却不能存留。
JOB|8|16|他在日光之下茂盛， 嫩枝在园中蔓延；
JOB|8|17|他的根盘绕石堆， 钻入石缝 。
JOB|8|18|他若从本地被拔出， 那地就不认识他，说：‘我没有见过你。’
JOB|8|19|看哪，这就是他道路中的喜乐， 以后必另有人从尘土而生。
JOB|8|20|看哪，上帝必不丢弃完全人， 也不扶助邪恶人的手。
JOB|8|21|他还要以喜笑充满你的口， 以欢呼充满你的嘴唇。
JOB|8|22|恨恶你的要披戴羞愧， 恶人的帐棚必归于无有。”
JOB|9|1|约伯 回答说：
JOB|9|2|“我真的知道是这样， 但人在上帝前怎能成为义呢？
JOB|9|3|人若想要与他争辩， 千次中也不能回答一次。
JOB|9|4|他心里有智慧，且大有能力。 谁向上帝刚硬而得平安呢？
JOB|9|5|他把山挪移，山却不知， 他在怒气中，把山翻倒。
JOB|9|6|他使地震动，离其本位， 地的柱子就摇撼。
JOB|9|7|他吩咐太阳，太阳就不出来， 又封住众星。
JOB|9|8|他独自铺张诸天， 步行在海浪之上。
JOB|9|9|他造北斗、参星、昴星， 以及南方的星宿 ；
JOB|9|10|他行大事不可测度， 行奇事不可胜数。
JOB|9|11|看哪，他从我旁边经过，我看不见； 他走过，我没有察觉他。
JOB|9|12|看哪，他夺去，谁能阻挡他？ 谁敢对他说：‘你做什么呢？’
JOB|9|13|“上帝必不收回他的怒气， 扶助 拉哈伯 的，屈身在上帝以下。
JOB|9|14|既是这样，我怎敢回答他， 怎敢在他之前选择辩词呢？
JOB|9|15|我虽有义，也不能回答， 我要向那审判我的恳求。
JOB|9|16|我若呼求，纵然他应允我， 我仍不信他会侧耳听我的声音。
JOB|9|17|他用暴风 摧折我， 无故加增我的损伤。
JOB|9|18|他不容我喘一口气， 倒使我饱受苦恼。
JOB|9|19|若论力量，看哪，他真有能力！ 若论审判，‘谁能传我呢？’
JOB|9|20|我虽有义，我的口要定我有罪； 我虽完全，他必证明我为弯曲。
JOB|9|21|我虽完全，不顾自己； 我厌弃我的性命。
JOB|9|22|所以我说，都是一样； 完全人和恶人，他都灭绝。
JOB|9|23|若灾祸忽然带来死亡， 他必戏笑无辜人的苦难。
JOB|9|24|世界交在恶人手中； 他蒙蔽世界审判官的脸， 若不是他，那么是谁呢？
JOB|9|25|“我的日子比奔跑者更快， 急速过去，不见福乐。
JOB|9|26|我的日子如蒲草船掠过， 如鹰俯冲抓食。
JOB|9|27|我若说：‘我要忘记我的苦情， 强颜欢笑’，
JOB|9|28|我就因一切的愁苦而惧怕； 我知道你必不以我为无辜。
JOB|9|29|我必被定罪， 我何必徒然劳苦呢？
JOB|9|30|我若用雪水洗身， 用碱洁净我的手掌，
JOB|9|31|你还要把我扔在坑里， 我的衣服都憎恶我。
JOB|9|32|他不像我是个人，使我可以回答他， 使我们可以一同受审判。
JOB|9|33|我们中间没有仲裁者， 可以按手在我们两造之间。
JOB|9|34|愿他使他的杖离开我， 不使他的威严恐吓我，
JOB|9|35|我就说话，不惧怕他； 但对我来说，我却不是这样。”
JOB|10|1|“我厌恶自己的性命， 任由我述说自己的苦情； 因心里苦恼，我要说话。
JOB|10|2|我对上帝说，不要定我有罪， 要指示我，你为何与我争辩？
JOB|10|3|你手所造的，你又欺压，又藐视， 却光照恶人的计谋。 这事你以为美吗？
JOB|10|4|你的眼岂是肉眼？ 你察看岂像人察看吗？
JOB|10|5|你的日子岂像人的日子， 你的年岁岂像壮士的年岁，
JOB|10|6|你就追问我的罪孽， 寻察我的罪过吗？
JOB|10|7|其实，你知道我没有行恶， 也无人能施行拯救，脱离你的手。
JOB|10|8|你的手塑造我，造了我， 但我整个人却要一起被你吞灭。
JOB|10|9|求你记得，你制造我如泥土， 你还要使我归回尘土吗？
JOB|10|10|你不是倒出我来好像奶， 使我凝结如同奶酪吗？
JOB|10|11|你以皮和肉给我穿上， 用骨与筋把我联结起来。
JOB|10|12|你将生命和慈爱赐给我， 你也眷顾保全我的灵。
JOB|10|13|然而，你把这些事藏在你心里， 我知道这是你的旨意。
JOB|10|14|我若犯罪，你就察看我， 并不赦免我的罪。
JOB|10|15|我若行恶，我就有祸了； 我若行义，也不敢抬头， 而是饱受羞辱， 看见我的痛苦。
JOB|10|16|你如狮子昂首追捕我 ， 又在我身上显出奇事。
JOB|10|17|你更新你的见证对付我， 向我加增恼怒， 调遣军队攻击我。
JOB|10|18|“你为何使我出母胎呢？ 甚愿我当时气绝，没有眼睛看见我。
JOB|10|19|这样，就如从未有过我， 我一出母胎就被送入坟墓。
JOB|10|20|我的日子不是短少吗？求你停止， 求你放过我 ，使我可以稍得喜乐，
JOB|10|21|就是在我去而不返， 往黑暗和死荫之地以先。
JOB|10|22|那是乌黑之地， 犹如幽暗的死荫， 毫无秩序； 发出的光辉也像幽暗。”
JOB|11|1|拿玛 人 琐法 回答说：
JOB|11|2|“这许多的话岂不该回答吗？ 多嘴多舌的人岂可成为义呢？
JOB|11|3|你夸大的话岂能使人不作声吗？ 你戏笑的时候岂没有人使你受辱吗？
JOB|11|4|你说：‘我的教导纯全， 我在你眼前是清洁的。’
JOB|11|5|但是，惟愿上帝说话， 愿他张开嘴唇攻击你。
JOB|11|6|愿他将智慧的奥秘指示你， 因为健全的知识是两面的。 你当知道，上帝使你忘记你的一些罪孽。
JOB|11|7|你能寻见上帝的奥秘吗？ 你能寻见全能者的极限吗？
JOB|11|8|高如诸天，你能做什么？ 比阴间深，你能知道什么？
JOB|11|9|其量度比地长， 比海更宽。
JOB|11|10|他若经过，把人拘禁， 召集会众，谁能阻挡他呢？
JOB|11|11|因为他知道虚妄的人； 当他看见罪恶，岂不留意吗？
JOB|11|12|空虚的人若获得知识， 野驴生下的驹子也成了人。
JOB|11|13|“至于你，若坚固己心， 又向主举手；
JOB|11|14|你若远远脱离你手中的罪孽， 不容许不义住在你帐棚之中；
JOB|11|15|这样，你必仰起脸来，毫无瑕疵； 你也必安稳，无所惧怕。
JOB|11|16|你必忘记你的苦楚， 就是想起来，也如流过的水。
JOB|11|17|你在世要升高，比正午更明， 虽有黑暗，仍像早晨。
JOB|11|18|你因有指望就必稳固， 也必四围察看 ，安然躺下。
JOB|11|19|你躺卧，无人惊吓， 并有许多人向你求恩。
JOB|11|20|但恶人的眼睛要失明； 他们无路可逃， 他们的指望就是气绝身亡。”
JOB|12|1|约伯 回答说：
JOB|12|2|“你们果真是人物啊！ 智慧要与你们一同去死。
JOB|12|3|但我也有聪明，跟你们一样， 并非不及你们。 这些事，谁不知道呢？
JOB|12|4|我这求告上帝、蒙他应允的人 竟成了朋友所讥笑的； 又公义又完全的人竟遭受讥笑。
JOB|12|5|安逸的人心里藐视灾祸， 这灾祸在等待失足滑跌的人。
JOB|12|6|强盗的帐棚安宁， 惹上帝发怒的人稳固， 他们把上帝 握在自己手中 。
JOB|12|7|“你问走兽，走兽必指教你； 你问空中的飞鸟，飞鸟必告诉你；
JOB|12|8|或者你与地说话，地必指教你 ； 海中的鱼也必向你说明。
JOB|12|9|在这一切当中， 有谁不知道这是耶和华的手做成的呢？
JOB|12|10|凡动物的生命 和人类的气息都在他手中。
JOB|12|11|耳朵岂不辨别言语， 正如上膛品尝食物吗？
JOB|12|12|年老的有智慧， 寿高的有知识。
JOB|12|13|“在上帝有智慧和能力， 他有谋略和知识。
JOB|12|14|看哪，他拆毁，就不能重建； 他拘禁人，人就不得释放。
JOB|12|15|看哪，他使水止住，水就干了； 他把水放出，水就淹没大地。
JOB|12|16|在他有能力和智慧， 走迷的和使人迷路的都属他。
JOB|12|17|他把谋士剥衣掳去， 使审判官变为愚妄。
JOB|12|18|他解除君王的权势 ， 用带子捆住他们的腰。
JOB|12|19|他把祭司剥衣掳去， 使有权能的人倾覆。
JOB|12|20|他废去忠信者的言论， 夺去长者的见识。
JOB|12|21|他使贵族蒙羞受辱， 放松勇士的腰带。
JOB|12|22|他从黑暗中彰显深奥的事， 使死荫显出光明。
JOB|12|23|他使邦国兴旺而又毁灭， 使邦国扩展又被掠夺。
JOB|12|24|他将地上百姓中领袖的聪明夺去， 使他们迷失在荒凉无路之地。
JOB|12|25|他们在无光的黑暗中摸索； 他使他们摇晃像醉酒的人一样。”
JOB|13|1|“看哪，这一切，我眼都见过； 我耳都听过，而且明白。
JOB|13|2|你们所知道的，我也知道， 并非不及你们。
JOB|13|3|然而我要对全能者说话， 我愿与上帝理论。
JOB|13|4|但你们是编造谎言的， 全都是无用的医生。
JOB|13|5|惟愿你们全然不作声， 这就是你们的智慧！
JOB|13|6|请你们听我的答辩， 留心听我嘴唇的诉求。
JOB|13|7|你们要为上帝说不义的话吗？ 要为他说诡诈的言语吗？
JOB|13|8|你们要看上帝的情面吗？ 要为他争辩吗？
JOB|13|9|他查究你们，这岂是好事吗？ 人欺骗人，你们也要照样欺骗他吗？
JOB|13|10|你们若暗中看人的情面， 他必定要责备你们。
JOB|13|11|他的尊荣岂不叫你们惧怕吗？ 他岂不使惊吓临到你们吗？
JOB|13|12|你们可记念的谚语是灰烬的箴言； 你们的后盾是泥土的后盾。
JOB|13|13|“你们不要向我作声， 让我说话，无论如何我都承当。
JOB|13|14|我为何把我的肉挂在我的牙上， 将我的命放在我的手掌中呢？
JOB|13|15|看哪，他要杀我，我毫无指望 ， 然而我还要在他面前辩明我所行的。
JOB|13|16|这要成为我的拯救， 因为不虔诚的人不可到他面前。
JOB|13|17|你们要细听我的言语， 让我的申辩入你们耳中。
JOB|13|18|看哪，我已陈明我的案， 知道自己有义。
JOB|13|19|还有谁要和我争辩， 我现在就缄默不言，气绝而死。
JOB|13|20|惟有两件事不要向我施行， 我就不躲开你的面：
JOB|13|21|就是把你的手缩回，远离我身； 又不使你的威严恐吓我。
JOB|13|22|这样，你呼叫，我就回答； 或是让我说话，你回答我。
JOB|13|23|我的罪孽和我的罪有多少呢？ 求你叫我知道我的过犯与我的罪。
JOB|13|24|你为何转脸， 拿我当仇敌呢？
JOB|13|25|你要惊动被风吹的叶子吗？ 要追赶枯干的碎秸吗？
JOB|13|26|你写下苦楚对付我， 又使我担当幼年的罪孽。
JOB|13|27|你把我的脚锁上木枷， 察看我一切的道路， 为我的脚掌划定界限。
JOB|13|28|人像灭绝的烂物， 像虫蛀的衣裳。”
JOB|14|1|“人为妇人所生， 日子短少，多有患难。
JOB|14|2|他出来如花，凋谢而去； 他飞逝如影，不能存留。
JOB|14|3|这样的人你岂会睁眼看他， 又叫我 来，在你那里受审吗？
JOB|14|4|谁能使洁净出于污秽呢？ 谁也不能！
JOB|14|5|既然人的日子限定， 他的月数在于你， 你划定他的界限，他不能越过；
JOB|14|6|求你转眼不看他，使他得歇息， 直到他像雇工享受他的一天。
JOB|14|7|“因树有指望， 若被砍下，还可发芽， 嫩枝生长不息。
JOB|14|8|树根若衰老在地里， 树干也死在土中，
JOB|14|9|及至得了水气，还会发芽， 长出枝条，像新栽的树一样。
JOB|14|10|但壮士一死就消逝了； 人一气绝，他在何处呢？
JOB|14|11|海中的水枯竭， 江河消散干涸。
JOB|14|12|人一躺下就不再起来， 等到诸天没有了 ，仍不复醒， 也不能从睡中唤醒。
JOB|14|13|惟愿你把我藏在阴间， 把我隐藏，直到你的愤怒过去； 愿你为我定下期限，并记得我。
JOB|14|14|壮士若死了能再活吗？ 我在一切服役的日子中等待， 直到我退伍的时候来到。
JOB|14|15|你呼叫，我就回答你； 你手所做的，你必期待。
JOB|14|16|但如今你数点我的脚步， 不察看我的罪。
JOB|14|17|我的过犯被你密封在囊中， 你遮掩了我的罪孽。
JOB|14|18|“然而，山崩变为无有， 磐石从原处挪移。
JOB|14|19|流水冲蚀石头， 急流洗去地上的尘土； 你也照样灭绝人的指望。
JOB|14|20|你终必胜过人，使他消逝； 你改变他的容貌，把他送走。
JOB|14|21|他的儿子得尊荣，他不知道； 他们降为卑，他也不晓得。
JOB|14|22|他只觉得身上疼痛， 心中为自己悲哀。”
JOB|15|1|提幔 人 以利法 回答说：
JOB|15|2|“智慧人岂可用虚空的知识回答， 用东风充满自己的肚腹呢？
JOB|15|3|他岂可用无益的话， 用无济于事的言语理论呢？
JOB|15|4|你诚然废弃敬畏， 不在上帝面前默想。
JOB|15|5|你的罪孽指教你的口； 你选用诡诈人的舌头。
JOB|15|6|你自己的口定你有罪，并非是我； 你自己的嘴唇见证你的不是。
JOB|15|7|“你是头一个生下来的人吗？ 你受造在诸山之先吗？
JOB|15|8|你曾听见上帝的密旨吗？ 你要独自得尽智慧吗？
JOB|15|9|什么是你知道，我们不知道的呢？ 什么是你明白，我们不明白的呢？
JOB|15|10|我们这里有白发的和年老的， 比你父亲还年长。
JOB|15|11|上帝的安慰和对你温和的话， 你以为太小吗？
JOB|15|12|你的心为何失控， 你的眼为何冒火，
JOB|15|13|以致你的灵反对上帝， 你的口说出这样的言语呢？
JOB|15|14|人是什么，竟算为洁净呢？ 妇人所生的是什么，竟算为义呢？
JOB|15|15|看哪，上帝不信任他的众圣者； 在他眼前，天也不洁净，
JOB|15|16|何况那污秽可憎， 喝罪孽如水的世人呢！
JOB|15|17|“我指示你，你要听我； 我要陈述我所看见的，
JOB|15|18|就是智慧人从列祖所受， 传讲而不隐瞒的事。
JOB|15|19|这地惟独赐给他们， 并没有外人从他们中间经过。
JOB|15|20|恶人一生的日子绞痛难熬， 残暴人存留的年数也是如此。
JOB|15|21|惊吓的声音常在他耳中； 在平安时，毁灭者必临到他。
JOB|15|22|他不信自己能从黑暗中转回； 他被刀剑看守。
JOB|15|23|他飘流在外求食：‘哪里有食物呢？’ 他知道黑暗的日子在他手边预备好了。
JOB|15|24|急难困苦叫他害怕， 而且胜过他，好像君王预备上阵。
JOB|15|25|因他伸手攻击上帝， 逞强对抗全能者，
JOB|15|26|挺着颈项， 用盾牌坚厚的凸面向全能者直闯；
JOB|15|27|又因他的脸蒙上油脂， 腰上积满肥肉。
JOB|15|28|他住在荒凉的城镇， 房屋无人居住， 将成为废墟。
JOB|15|29|他不得富足， 财物不得常存， 产业在地上也不加增。
JOB|15|30|他不得脱离黑暗， 火焰要把他的嫩枝烧干； 因上帝口中的气，他要离去。
JOB|15|31|不要让他倚靠虚假，欺骗自己， 因虚假必成为他的报应。
JOB|15|32|他的日期未到之先，这事必实现； 他的枝子不得青绿。
JOB|15|33|他必像葡萄树，葡萄未熟就掉落； 又像橄榄树，一开花就凋谢。
JOB|15|34|因不敬虔之辈必不能生育， 受贿赂之人的帐棚必被火吞灭。
JOB|15|35|他们所怀的是毒害，所生的是罪孽， 肚腹里所预备的是诡诈。”
JOB|16|1|约伯 回答说：
JOB|16|2|“这样的话我听了许多； 你们全都是使人愁烦的安慰者。
JOB|16|3|如风的言语有穷尽吗？ 或者什么惹动你回答呢？
JOB|16|4|我也能说你们那样的话， 你们若处在我的景况， 我也可以堆砌言词攻击你们， 又可以向你们摇头。
JOB|16|5|但我必用口坚固你们， 颤动的嘴唇带来舒解。
JOB|16|6|“我若说话，痛苦仍不得缓解； 我若停止，痛苦就离开我吗？
JOB|16|7|但现在上帝使我困倦， 你使所有的亲友远离我，
JOB|16|8|你抓住我 ，成为见证起来攻击我； 我的枯瘦也当着我的面作证。
JOB|16|9|上帝发怒撕裂我，逼迫我， 向我咬牙切齿； 我的敌人怒目瞪我。
JOB|16|10|他们向我大大张口， 打我的耳光羞辱我， 聚在一起攻击我。
JOB|16|11|上帝把我交给不敬虔的人， 把我扔到恶人的手中。
JOB|16|12|我本是安逸，他折断我， 掐住我的颈项，把我摔碎， 又立我作他的箭靶。
JOB|16|13|他的弓箭手围绕我。 他刺破我的肾脏，并不留情， 把我的胆汁倾倒在地上。
JOB|16|14|他使我破裂，破裂又破裂， 如同勇士向我直闯。
JOB|16|15|“我把麻布缝在我的皮肤上， 把我的角放在尘土中。
JOB|16|16|我的脸因哭泣变红， 我的眼皮上有死荫。
JOB|16|17|我的手中却没有暴力， 我的祈祷也是纯洁的。
JOB|16|18|“地啊，不要遮盖我的血！ 不要让我的哀求有藏匿之处！
JOB|16|19|现今，看哪，在天有我的见证， 在上有我的保人。
JOB|16|20|我的朋友讥诮我， 我却向上帝眼泪汪汪。
JOB|16|21|愿人可与上帝理论， 如同人与朋友一样；
JOB|16|22|因为再过几年， 我必走那往而不返之路。”
JOB|17|1|“我的灵耗尽，我的日子消逝； 坟墓为我预备好了。
JOB|17|2|戏笑的人果真陪伴着我， 我的眼睛盯住他们的悖逆。
JOB|17|3|“愿你亲自为我付押担保。 谁还会与我击掌呢？
JOB|17|4|因你蒙蔽他们的心，使不明理， 所以你必不高举他们。
JOB|17|5|控告 朋友为了分享产业的， 他儿女的眼睛要失明。
JOB|17|6|“上帝使我成为人群中的笑谈， 他们吐唾沫在我脸上。
JOB|17|7|我的眼睛因忧愁昏花， 我的肢体全像影儿。
JOB|17|8|正直人因此必惊奇； 无辜的人要兴起攻击不敬虔之辈。
JOB|17|9|然而，义人要持守所行的道， 手洁的人要力上加力。
JOB|17|10|至于你们众人，再回来吧！ 你们中间，我找不到一个智慧人。
JOB|17|11|我的日子已经过去了， 我的谋算、我心的愿望已经断绝了。
JOB|17|12|他们以黑夜为白昼， 即使面临黑暗，以为亮光已近。
JOB|17|13|我若盼望阴间为我的家， 若下榻在黑暗中，
JOB|17|14|若对地府呼叫：‘你是我的父亲’， 若对虫呼叫：‘你是我的母亲、姊妹’，
JOB|17|15|这样，我的盼望在哪里呢？ 我所盼望的，谁能看见呢？
JOB|17|16|这盼望要下到阴间的门闩吗 ？ 要一起在尘土中安息吗 ？”
JOB|18|1|书亚 人 比勒达 回答说：
JOB|18|2|“你们寻索言语要到几时呢 ？ 你们要明白，然后我们才说话。
JOB|18|3|我们为何被视为畜生， 在你们眼中看为愚笨 呢？
JOB|18|4|在怒气中将自己撕裂的人哪， 难道大地要因你见弃、 磐石要挪开原处吗？
JOB|18|5|“恶人的亮光必要熄灭， 他的火焰必不照耀。
JOB|18|6|他帐棚中的亮光要变黑暗， 他上面的灯也必熄灭。
JOB|18|7|他强横的脚步必遭阻碍， 他的计谋必将自己绊倒。
JOB|18|8|他因自己的脚陷入网中， 走在缠人的网子上。
JOB|18|9|罗网必抓住他的脚跟， 陷阱必擒获他。
JOB|18|10|绳索为他藏在土里， 羁绊为他藏在路上。
JOB|18|11|四面的惊吓使他害怕， 在他脚跟后面追赶他。
JOB|18|12|他的力量必因饥饿衰败， 祸患要在他的旁边等候，
JOB|18|13|侵蚀他肢体的皮肤； 死亡的长子吞吃他的肢体。
JOB|18|14|他要从所倚靠的帐棚被拔出来， 带到使人惊恐的王那里。
JOB|18|15|不属他的必住在他的帐棚里， 硫磺必撒在他所住之处。
JOB|18|16|下边，他的根要枯干； 上边，他的枝子要剪除。
JOB|18|17|他的称号 从地上消失， 他的名字不在街上存留。
JOB|18|18|他必从光明中被驱逐到黑暗里， 他必被赶出世界。
JOB|18|19|他在自己百姓中必无子无孙， 在寄居之地也没有幸存者。
JOB|18|20|以后的人 要因他的日子惊讶， 以前的人 也被惊骇抓住。
JOB|18|21|不义之人的住处总是这样， 这就是不认识上帝之人的下场。”
JOB|19|1|约伯 回答说：
JOB|19|2|“你们搅扰我的心， 用言语压碎我要到几时呢？
JOB|19|3|你们这十次羞辱我， 苦待我也不以为耻。
JOB|19|4|果真我有错， 这错是在于我。
JOB|19|5|若你们真要向我夸大， 以我的羞辱来责备我，
JOB|19|6|就该知道是上帝倾覆我， 用罗网围绕我。
JOB|19|7|看哪，我喊冤叫屈，却不蒙应允； 我呼求，却没有公正。
JOB|19|8|上帝拦住我的道路，使我不得经过； 他使黑暗笼罩我的路径。
JOB|19|9|他剥去我的荣光， 摘去我头上的冠冕。
JOB|19|10|他在四围攻击我，我就走了； 他将我的指望如树拔出。
JOB|19|11|他向我发烈怒， 以我为他的敌人。
JOB|19|12|他的军队一齐上来， 修筑道路攻击我， 在我帐棚的四围安营。
JOB|19|13|“他把我的兄弟隔在远处， 使我认识的人全然与我生疏。
JOB|19|14|我的亲戚都离开了我； 我的密友都忘记了我。
JOB|19|15|在我家寄居的和我的使女， 都当我是陌生人； 我在他们眼中被视为外邦人。
JOB|19|16|我呼唤仆人，他却不回答； 我必须亲口求他。
JOB|19|17|我口的气味令我妻子厌恶， 我的同胞都憎恶我。
JOB|19|18|连小男孩也藐视我； 我起来，他们都嘲笑我。
JOB|19|19|我的知心朋友都憎恶我； 我平日所爱的人向我翻脸。
JOB|19|20|我的皮和肉紧贴骨头， 我得以逃脱，仅剩牙齿 。
JOB|19|21|我的朋友啊，可怜我！可怜我！ 因为上帝的手攻击我。
JOB|19|22|你们为什么仿佛上帝逼迫我， 吃我的肉还不满足呢？
JOB|19|23|“惟愿我的言语现在就写上， 都记录在书上；
JOB|19|24|用铁笔和铅， 刻在磐石上，存到永远。
JOB|19|25|我知道我的救赎主 活着， 末后他必站在尘土上。
JOB|19|26|我这皮肉灭绝之后 ， 我必在肉体之外 得见上帝。
JOB|19|27|我自己要见他， 亲眼要看他，并不像陌生人。 我的心肠在我里面耗尽了！
JOB|19|28|你们若说：‘我们怎么逼迫他呢？ 事情的根源是在于他 ’，
JOB|19|29|你们就当惧怕刀剑， 因为愤怒带来刀剑的刑罚。 这样，你们就知道有审判。”
JOB|20|1|拿玛 人 琐法 回答说：
JOB|20|2|“这样，我的思念叫我回答， 因为我心中急躁。
JOB|20|3|我听见那羞辱我的责备； 我悟性的灵回答我。
JOB|20|4|你岂不知道吗？亘古以来， 自从人被安置在地，
JOB|20|5|恶人欢乐的声音是暂时的， 不敬虔人的喜乐不过是转眼之间。
JOB|20|6|他的尊荣虽达到天上， 头虽顶到云中，
JOB|20|7|他必永远灭亡，像自己的粪一样。 看见他的人要说：‘他在哪里呢？’
JOB|20|8|他必如梦飞去，不再寻见； 他被赶走，如夜间的异象。
JOB|20|9|亲眼见过他的，必不再见他； 他自己的地方也不再见到他。
JOB|20|10|他的儿女要向穷人求恩； 他的手要赔还钱财。
JOB|20|11|他的骨头虽然满有年轻的活力， 却要和他一同躺卧在尘土之中。
JOB|20|12|“他口中以恶为甘甜， 把恶藏在舌头底下，
JOB|20|13|爱恋不舍， 含在口中。
JOB|20|14|他的食物在肚里却要翻转， 在他里面成为虺蛇的毒液。
JOB|20|15|他吞了财宝，还要吐出； 上帝要从他腹中掏出来。
JOB|20|16|他必吸饮虺蛇的毒汁， 毒蛇的舌头必杀他。
JOB|20|17|他不再看见溪流， 流奶与蜜之河。
JOB|20|18|他劳碌得来的要赔还，不得吞下； 赚取了财货，也不得欢乐。
JOB|20|19|他欺压穷人，弃之不顾， 强取非自己所盖的房屋 。
JOB|20|20|“他的肚腹不知安逸， 所贪恋的连一样也不放过，
JOB|20|21|剩余的没有一样他不吞吃， 所以他的福乐不能长久。
JOB|20|22|他在满足有余的时候，必有困苦临到； 凡受苦楚之人的手必加在他身上。
JOB|20|23|他的肚腹正要满足的时候， 上帝必将猛烈的愤怒降在他身上； 他正在吃饭的时候， 上帝要将这愤怒如雨降在他身上。
JOB|20|24|他要躲避铁的武器， 铜弓要将他射透。
JOB|20|25|箭一抽，就从他背上出来， 发亮的箭头从他胆中出来； 有惊惶临到他身上。
JOB|20|26|他的财宝隐藏在深沉的黑暗里； 有非人吹起的火要把他吞灭， 把他帐棚中所剩下的烧毁。
JOB|20|27|天要显明他的罪孽， 地要兴起去攻击他。
JOB|20|28|他家里出产的必消失， 在上帝愤怒的日子被冲走。
JOB|20|29|这是恶人从上帝所得的份， 是上帝为他所定的产业。”
JOB|21|1|约伯 回答说：
JOB|21|2|“你们要细心听我的言语， 这就算是你们的安慰。
JOB|21|3|请宽容我，我又要说话； 说了以后，任凭你嗤笑吧！
JOB|21|4|我岂是向人诉苦？ 我为何不是没有耐心呢？
JOB|21|5|你们要转向我而惊奇， 要用手捂口。
JOB|21|6|我每逢思想，心就惊惶， 战兢抓住我身。
JOB|21|7|恶人为何存活， 得享高寿，势力强盛呢？
JOB|21|8|他们的后裔与他们一起 ，坚立在他们面前， 他们得以眼见自己的子孙。
JOB|21|9|他们的家宅平安无惧， 上帝的杖不加在他们身上。
JOB|21|10|他们的公牛传种而不断绝， 母牛生牛犊而不掉胎。
JOB|21|11|他们打发小男孩出去，多如羊群， 他们的孩子踊跃跳舞。
JOB|21|12|他们随着琴鼓歌唱， 因箫声欢喜。
JOB|21|13|他们度日诸事亨通， 在平安中下到阴间。
JOB|21|14|他们对上帝说：‘离开我们吧！ 我们不想知道你的道路。
JOB|21|15|全能者是谁，我们何必事奉他呢？ 求告他有什么益处呢？’
JOB|21|16|看哪，他们亨通不是靠自己的手； 恶人的计谋离我好远。
JOB|21|17|“恶人的灯何尝熄灭？ 患难何尝临到他们呢？ 上帝何尝发怒，把灾祸分给他们呢？
JOB|21|18|他们何尝像风前的碎秸， 如暴风刮去的糠秕呢？
JOB|21|19|上帝为恶人的儿女积蓄罪孽， 不如本人遭报，好使他亲自知道。
JOB|21|20|愿他亲眼看见自己败亡， 亲自饮全能者的愤怒。
JOB|21|21|他的岁月既尽， 他身后还顾他的家吗？
JOB|21|22|谁能将知识教导上帝呢？ 是他审判那些居高位的。
JOB|21|23|有人至死身体强壮， 尽得平顺安逸；
JOB|21|24|他的肚腹充满奶汁 ， 他的骨髓滋润。
JOB|21|25|有人至死心中痛苦， 从未尝过福乐的滋味；
JOB|21|26|他们同样躺卧于尘土， 虫子覆盖他们。
JOB|21|27|“看哪，我知道你们的意念， 并残害我的计谋。
JOB|21|28|你们说：‘权贵的房屋在哪里？ 恶人住过的帐棚在哪里？’
JOB|21|29|你们没有询问那些过路的人吗？ 你们不承认他们的证据吗？
JOB|21|30|就是恶人在患难的日子得存留， 在愤怒的日子得逃脱。
JOB|21|31|他所行的，有谁当面给他说明？ 他所做的，有谁报应他呢？
JOB|21|32|然而他要被抬到坟地， 并有人看守墓穴。
JOB|21|33|他要以谷中的土块为甘甜； 人人要跟在他后面， 在他前面去的无数。
JOB|21|34|你们怎能以空话安慰我呢？ 你们的对答全都错谬！”
JOB|22|1|提幔 人 以利法 回答说：
JOB|22|2|“人能使上帝有益吗？ 智慧人能使他有益吗？
JOB|22|3|你为人公义，岂能叫全能者喜悦呢？ 你行为完全，岂能使他得利呢？
JOB|22|4|他岂是因你敬畏的心就责备你， 审判你吗？
JOB|22|5|你的罪恶岂不是大吗？ 你的罪孽不是没有穷尽吗？
JOB|22|6|因你无故强取弟兄的抵押， 剥去赤身者的衣服。
JOB|22|7|疲乏的人，你没有给他水喝； 饥饿的人，你没有给他食物。
JOB|22|8|有能力的人得土地； 尊贵的人住在其中。
JOB|22|9|你打发寡妇空手回去， 你折断孤儿的膀臂。
JOB|22|10|因此，有罗网环绕你， 有恐惧忽然使你惊惶；
JOB|22|11|或有黑暗使你看不见 ， 有洪水淹没你。
JOB|22|12|“上帝岂不是在高天吗？ 你看星宿的顶点何其高呢！
JOB|22|13|你说：‘上帝知道什么？ 他岂能透过幽暗施行审判呢？
JOB|22|14|密云将他遮盖，使他不能看见； 他周游穹苍。’
JOB|22|15|你要依从上古的道吗？ 这道是恶人行过的。
JOB|22|16|他们未到时候就被抓去 ； 他们的根基被江河冲去。
JOB|22|17|他们向上帝说：‘离开我们吧！’ 全能者能把他们怎么样呢？
JOB|22|18|然而，是上帝以美物充满他们的房屋； 恶人的计谋离我好远！
JOB|22|19|义人看见他们的结局 就欢喜； 无辜的人嗤笑他们：
JOB|22|20|‘攻击我们的果然被剪除， 剩余的都被火吞灭。’
JOB|22|21|“你要与上帝和好，要和平， 这样，福气必临到你。
JOB|22|22|你当领受他口中的教导， 将他的言语存在心里。
JOB|22|23|你若归向全能者，就必得建立。 你要从你帐棚中远离不义，
JOB|22|24|你要将黄金丢到尘土里， 将 俄斐 的金子丢在溪河石头之间；
JOB|22|25|全能者就必作你的黄金， 作你成堆的银子。
JOB|22|26|那时，你要以全能者为喜乐， 向上帝仰脸。
JOB|22|27|你要向他祷告，他就听你； 你也要还你的愿。
JOB|22|28|你定意要做何事，必然为你成就； 亮光也必照耀你的路。
JOB|22|29|当人降卑，你说：是因骄傲； 眼目谦卑的人，上帝必然拯救。
JOB|22|30|不是无辜的人，上帝尚且要搭救他 ； 他必因你手中的清洁得蒙拯救。”
JOB|23|1|约伯 回答说：
JOB|23|2|“如今我的哀告还算为悖逆； 我虽唉哼，他的手仍然重重责罚我 。
JOB|23|3|惟愿我知道哪里可以寻见上帝， 能到他的台前，
JOB|23|4|我就在他面前陈明我的案件， 满口辩诉。
JOB|23|5|我必知道他回答我的言语， 明白他向我所要说的。
JOB|23|6|他岂用大能与我争辩呢？ 不！他必理会我。
JOB|23|7|在那里正直人可以与他辩论， 我就必永远脱离那审判我的。
JOB|23|8|“看哪，我往前走，他不在那里； 往后退，也没有察觉他。
JOB|23|9|他在左边行事，我却看不见他； 他转向右边 ，我也见不到他。
JOB|23|10|然而他知道我所走的路； 他试炼我，我就如纯金。
JOB|23|11|我的脚紧跟他的步伐； 我谨守他的道，并不偏离。
JOB|23|12|他嘴唇的命令，我未曾背弃； 我看重他口中的言语，过于我需用的饮食 。
JOB|23|13|只是他心志已定，谁能使他转意呢？ 他心里所愿的，就行出来。
JOB|23|14|因此，为我所定的，他必做成， 这类的事他还有许多。
JOB|23|15|所以我在他面前惊惶； 我思想就惧怕他。
JOB|23|16|上帝使我丧胆， 全能者使我惊惶。
JOB|23|17|但我并非被黑暗剪除， 只是幽暗遮盖了我的脸。
JOB|24|1|“为何全能者不定下期限？ 为何认识他的人看不到那些日子呢？
JOB|24|2|有人挪移地界， 抢夺群畜去放牧。
JOB|24|3|他们拉走孤儿的驴， 强取寡妇的牛作抵押。
JOB|24|4|他们使贫穷人离开正道； 世上的困苦人尽都隐藏。
JOB|24|5|看哪，他们如同野驴出到旷野，殷勤寻找食物， 在野地给孩童糊口。
JOB|24|6|他们收割别人田间的庄稼， 摘取恶人剩余的葡萄。
JOB|24|7|他们终夜赤身无衣， 在寒冷中毫无遮盖。
JOB|24|8|他们在山上被大雨淋湿， 因没有避身之处就拥抱磐石。
JOB|24|9|又有人从母怀中抢走孤儿， 在困苦人身上强取抵押品 。
JOB|24|10|困苦人赤身无衣，到处流浪， 饿着肚子扛抬禾捆，
JOB|24|11|他们在围墙内榨油， 踹压酒池，自己却口渴。
JOB|24|12|在城内垂死的人呻吟， 受伤的人哀号； 上帝却不理会狂妄的事。
JOB|24|13|“又有人背弃光明， 不认识光明的道， 不留在光明的路上。
JOB|24|14|杀人者黎明起来， 杀害困苦人和贫穷人， 夜间又作盗贼。
JOB|24|15|奸夫的眼等候黄昏， 说：‘没有眼睛能见我’， 就把脸蒙住。
JOB|24|16|盗贼黑夜挖洞； 他们白日躲藏， 并不认识光明。
JOB|24|17|他们全都看早晨如死荫， 因为他们熟悉死荫的惊骇。
JOB|24|18|“恶人在水面上快速飘荡， 他们在地上所得的产业被诅咒； 无人再回到他们的葡萄园。
JOB|24|19|干旱炎热融化雪水； 阴间也如此吞没犯罪的人。
JOB|24|20|怀他的母胎忘记他； 虫子要吃他，觉得甘甜； 他不再被人记念； 不义的人必如树折断。
JOB|24|21|“他与不怀孕不生育的妇人交往 ， 却不善待寡妇。
JOB|24|22|然而上帝用能力保全有势力的人； 那性命难保的人仍然兴起。
JOB|24|23|上帝使他安稳，他就有所倚靠； 上帝的眼目看顾他们的道路。
JOB|24|24|他们高升，不过片刻就没有了； 他们降为卑，被除灭，与众人一样 ， 又如谷的穗子被割下。
JOB|24|25|若不是这样，谁能指证我是说谎的， 以我的言语为毫无根据呢？”
JOB|25|1|书亚 人 比勒达 回答说：
JOB|25|2|“上帝有统治之权，威严可畏； 他在高处施行和平。
JOB|25|3|他的军队岂能数算？ 他的光向谁不会升起呢 ？
JOB|25|4|这样，在上帝面前人怎能称义？ 妇人所生的怎能洁净？
JOB|25|5|看哪，在上帝眼前，月亮无光， 星宿也不皎洁，
JOB|25|6|更何况是如虫的人， 如蛆的世人呢！
JOB|26|1|约伯 回答说：
JOB|26|2|“无能的人蒙你何等的帮助！ 膀臂无力的人蒙你何等的拯救！
JOB|26|3|无智慧的人蒙你何等的指教！ 你向他显出丰富的知识。
JOB|26|4|你向谁发出言语？ 谁的灵从你而出？
JOB|26|5|在大水和水族以下， 阴魂战兢。
JOB|26|6|在上帝面前，阴间显露； 冥府 也不得遮掩。
JOB|26|7|上帝将北极铺在空中， 将大地悬在虚空。
JOB|26|8|他将水包在密云中， 盛水的云却不破裂。
JOB|26|9|他遮蔽宝座的正面， 把他的云彩铺在其上。
JOB|26|10|他在水面上划一圆圈， 直到光明与黑暗的交界。
JOB|26|11|天的柱子震动， 因他的斥责惊奇。
JOB|26|12|他以能力搅动 大海 ， 藉知识打伤 拉哈伯 。
JOB|26|13|他藉自己的灵使天空晴朗； 他的手刺杀爬得快的蛇。
JOB|26|14|看哪，这不过是上帝工作的些微； 我们听见他的话，是何等细微的声音！ 他大能的雷声谁能明白呢？”
JOB|27|1|约伯 继续发表他的言论说：
JOB|27|2|“我指着夺去我公道的永生上帝， 并使我心中愁苦的全能者起誓：
JOB|27|3|只要我的生命尚在我里面， 上帝所赐的气息仍在我鼻孔内，
JOB|27|4|我的唇绝不说不义， 我的舌也不说诡诈。
JOB|27|5|我断不以你们为义； 我至死不放弃自己的纯正！
JOB|27|6|我持定我的义，并不放松； 在世的日子，我的心不责备我。
JOB|27|7|“愿我的仇敌如恶人一样； 愿那起来攻击我的，如不义之人一般。
JOB|27|8|不敬虔的人有什么指望呢？ 上帝要剪除他，取他的性命。
JOB|27|9|患难临到他， 上帝岂听他的呼求？
JOB|27|10|他岂以全能者为乐， 随时求告上帝呢？
JOB|27|11|上帝手所做的，我要指教你们； 全能者所行的，我也不会隐瞒。
JOB|27|12|看哪，你们自己也都见过， 为何全变为这样虚妄呢？
JOB|27|13|“这是上帝为恶人所定的份， 残暴人从全能者所得的产业：
JOB|27|14|倘若他的儿女增多，仍被刀所杀； 他的子孙必不得饱食。
JOB|27|15|他遗留的人必死而埋葬， 他的寡妇也不哀哭。
JOB|27|16|他虽积蓄银子如尘沙， 堆积衣服如泥土，
JOB|27|17|他尽管堆积，义人却要穿上， 无辜的人却要分取银子。
JOB|27|18|他建造房屋如虫做窝， 又如守望者所搭的棚。
JOB|27|19|他虽富足躺卧，却不得收殓 ， 他张开眼睛，就不在了。
JOB|27|20|惊恐如洪水将他追上， 暴风在夜间将他刮去。
JOB|27|21|东风把他吹去，他就走了； 风将他刮离原地。
JOB|27|22|风 无情地击打他， 他试图逃脱风的手。
JOB|27|23|风要因他拍掌， 并要发叱声，使他离开原地。”
JOB|28|1|“银子有矿； 炼金有场。
JOB|28|2|铁从土里开采， 铜从矿石镕出。
JOB|28|3|人探索黑暗的尽头， 查究矿石直到极处， 那是幽暗和死荫；
JOB|28|4|他在无人居住之处开凿矿穴， 在无足迹之地被遗忘 ， 与人远离，悬空摇摆。
JOB|28|5|地出产粮食， 地底翻腾如火。
JOB|28|6|地的石头是蓝宝石之处， 那里还有金沙。
JOB|28|7|鸷鸟不知那条路， 鹰眼也未曾见过。
JOB|28|8|狂傲的野兽未曾踩踏， 猛烈的狮子也未曾经过。
JOB|28|9|“人动手凿开坚石， 翻倒山的根基，
JOB|28|10|在磐石中凿出水道， 亲眼看见各样宝物。
JOB|28|11|他封闭河川不得涓滴 ， 使隐藏之物显露出来。
JOB|28|12|“然而，智慧何处可寻？ 聪明之地在哪里？
JOB|28|13|智慧的价值 无人能知， 活人之地也无处可寻。
JOB|28|14|深渊说：‘不在我里面。’ 沧海说：‘不在我这里。’
JOB|28|15|智慧不可用黄金换取， 也不能用白银秤她的价值。
JOB|28|16|俄斐 的金子和贵重的红玛瑙， 以及蓝宝石，不足与她比拟；
JOB|28|17|黄金和玻璃不足与她比较； 纯金的器皿不足兑换她。
JOB|28|18|珊瑚、水晶都不值得提； 智慧的价值胜过宝石 。
JOB|28|19|古实 的红璧玺不足与她比较； 纯金也不足与她比拟。
JOB|28|20|“智慧从何处来呢？ 聪明之地在哪里？
JOB|28|21|她隐藏，远离众生的眼目， 她掩蔽，远离空中的飞鸟。
JOB|28|22|毁灭和死亡说： ‘我们风闻其名。’
JOB|28|23|“上帝明白智慧的道路， 知道智慧的所在。
JOB|28|24|因为他鉴察直到地极， 遍观普天之下，
JOB|28|25|要为风定轻重， 又度量诸水，
JOB|28|26|为雨定律例， 为雷电定道路。
JOB|28|27|那时他看见智慧，就谈论她， 坚定她，并且查究她。
JOB|28|28|他对人说：‘看哪，敬畏主就是智慧； 远离恶事就是聪明。’”
JOB|29|1|约伯 继续发表他的言论说：
JOB|29|2|“惟愿我如从前的岁月， 如上帝保护我的日子。
JOB|29|3|那时他的灯照在我头上， 我藉他的光行过黑暗。
JOB|29|4|在我壮年的时候， 上帝亲密的情谊临到我的帐棚中。
JOB|29|5|全能者仍与我同在， 我的儿女都环绕我。
JOB|29|6|我的脚洗在乳酪当中； 磐石为我流出油河。
JOB|29|7|我出到城门， 在广场安排座位，
JOB|29|8|年轻人见我而回避， 老年人起身站立。
JOB|29|9|王子都停止说话， 用手捂口；
JOB|29|10|领袖静默无声， 舌头贴住上膛。
JOB|29|11|耳朵听见了，称我有福； 眼睛看见了，就称赞我。
JOB|29|12|因我拯救了哀求的困苦人 和无人帮助的孤儿。
JOB|29|13|将要灭亡的为我祝福， 我使寡妇心中欢呼。
JOB|29|14|我穿上公义，它遮蔽我； 我的公平如外袍和冠冕。
JOB|29|15|我作瞎子的眼， 瘸子的脚。
JOB|29|16|我作贫穷人的父； 我不认识之人的案件，我也去查明。
JOB|29|17|我打破不义之人的大牙， 从他牙齿中夺走他所抢的。
JOB|29|18|我说：‘我要增添我的日子如尘沙， 我必死在自己家中 。
JOB|29|19|我的根伸展到水边， 露水夜宿我的枝上。
JOB|29|20|我的荣耀在我身上更新， 我的弓在我手中日新。’
JOB|29|21|“人听我说话而等候， 为我的教导而静默。
JOB|29|22|我说话之后，他们就不再说； 我的言语滴在他们身上。
JOB|29|23|他们等候我如等雨水， 又张口如切慕春雨。
JOB|29|24|我向他们微笑，他们不敢相信； 他们不使我脸上的光失色。
JOB|29|25|我为他们选择道路，又坐首位； 我如君王在军队中居住， 又如人安慰哀伤的人。”
JOB|30|1|“但如今，比我年轻的人讥笑我； 我曾藐视他们的父亲， 不放在我的牧羊犬中。
JOB|30|2|他们的精力既已衰败， 手中的气力于我何益？
JOB|30|3|他们因穷乏饥饿，没有生气， 在荒废凄凉的幽暗中啃干燥之地。
JOB|30|4|他们在草丛之中采咸草， 罗腾 树的根成为他们的食物。
JOB|30|5|他们从人群中被赶出， 人追喊他们如贼一般，
JOB|30|6|以致他们住在荒谷， 住在地洞和岩穴中。
JOB|30|7|他们在草丛中叫唤， 在荆棘下挤成一团。
JOB|30|8|这都是愚顽卑微人的儿女； 他们被鞭打，赶出境外。
JOB|30|9|“现在这些人以我为歌曲， 以我为笑谈。
JOB|30|10|他们厌恶我，躲避我， 不住地吐唾沫在我脸上。
JOB|30|11|上帝松开我的弓弦 使我受苦， 他们就在我面前脱去辔头。
JOB|30|12|这伙人在我右边起来， 他们推开我的脚， 筑灾难之路攻击我。
JOB|30|13|他们毁坏我的道， 加增我的灾害； 他们毋须人帮助。
JOB|30|14|他们来，如同闯进大缺口， 在暴风间滚动。
JOB|30|15|惊恐倾倒在我身上， 我的尊荣被逐如风； 我的福禄如云飘去。
JOB|30|16|“现在我的心极其悲伤， 困苦的日子将我抓住。
JOB|30|17|夜间，我里面的骨头刺痛， 啃着我的没有止息。
JOB|30|18|我的外衣因大力扭皱 ， 内衣的领子把我勒住。
JOB|30|19|上帝把我扔在淤泥之中， 我就像尘土和灰烬一样。
JOB|30|20|我呼求你，你不应允我； 我站起来，你只是望着我。
JOB|30|21|你对我变得残忍， 大能的手追逼我。
JOB|30|22|你把我提到风中，使我乘风而去， 使我消失在烈风之中。
JOB|30|23|我知道你要使我归于死亡， 到那为众生所定的阴宅。
JOB|30|24|“然而，人在废墟岂不伸手？ 遇灾难时一定呼救。
JOB|30|25|人遭难的日子，我岂不为他哭泣呢？ 人贫穷的时候，我岂不为他忧愁呢？
JOB|30|26|我仰望福气，灾祸就来到； 我等待光明，黑暗便来临。
JOB|30|27|我内心烦扰不安， 困苦的日子临到我身。
JOB|30|28|我在阴暗中行走，没有日光 ， 我在会众中站立求救。
JOB|30|29|我与野狗为弟兄， 我跟鸵鸟为同伴。
JOB|30|30|我的皮肤变黑脱落， 我的骨头因热烧焦。
JOB|30|31|我的琴音变为哀泣； 我的箫声变为哭声。”
JOB|31|1|“我与眼睛立约， 怎能凝望少女呢？
JOB|31|2|从至上的上帝所得之分， 从至高全能者所得之业是什么呢？
JOB|31|3|岂不是祸患临到不义的， 灾害临到作恶的吗？
JOB|31|4|上帝岂不察看我的道路， 数点我所有的脚步吗？
JOB|31|5|“我若与虚谎同行， 我脚若紧跟诡诈，
JOB|31|6|愿上帝用公道的天平秤我， 愿他知道我的纯正。
JOB|31|7|我的脚步若偏离正路， 我的心若随从我眼目， 我的手掌若粘有污秽；
JOB|31|8|愿我栽种，别人来吃， 我的农作物连根拔出。
JOB|31|9|“我心若因妇人受迷惑， 在邻舍的门外等候，
JOB|31|10|就愿我妻子给别人推磨， 别人与她同寝。
JOB|31|11|因为这是邪恶的事， 审判官裁定的罪孽。
JOB|31|12|这是一场火，直烧到毁灭 ， 必拔除我一切的家产。
JOB|31|13|“我的仆婢与我争辩， 我若藐视不听他们的冤情，
JOB|31|14|上帝兴起的时候，我怎样行呢？ 他察问的时候，我怎样回答他呢？
JOB|31|15|造我在母腹中的，不也是造了他吗？ 在母胎中使我们成形的，岂不是同一位吗？
JOB|31|16|“我若不让贫寒人遂其所愿， 或是叫寡妇眼中失望，
JOB|31|17|或独自吃自己的食物， 孤儿没有吃其中些许；
JOB|31|18|从我年轻时，孤儿就与我一同长大，我好像他的父亲， 我从出母腹就扶助寡妇 ；
JOB|31|19|我若见人因无衣死亡， 或见贫穷人毫无遮盖；
JOB|31|20|我若不使他真心为我祝福， 不使他因我羊的毛得暖；
JOB|31|21|我若举手攻击孤儿， 因为在城门口见有帮助我的；
JOB|31|22|情愿我的肩膀从肩胛骨脱落， 我的膀臂从肱骨折断。
JOB|31|23|因上帝降的灾祸使我恐惧 ， 因他的威严，我什么都不能。
JOB|31|24|“我若以黄金为我的指望， 对纯金说：你是我的倚靠；
JOB|31|25|我若因财物丰裕， 因手多得资财而欢喜；
JOB|31|26|我若见太阳发光， 明月运行，
JOB|31|27|心就暗暗被引诱， 口亲吻自己的手；
JOB|31|28|这也是审判官裁定的罪孽， 因为我背弃了至上的上帝。
JOB|31|29|“我若见恨我的遇难就欢喜， 见他遭灾就高兴；
JOB|31|30|其实我没有容许口犯罪， 以诅咒要他的性命；
JOB|31|31|若我帐棚中的人未曾说： ‘谁不以他的肉食吃饱呢？’
JOB|31|32|我未曾让旅客在街上过夜， 却开门迎接行路的人；
JOB|31|33|我若像 亚当 遮掩自己的过犯， 将罪孽藏在怀中；
JOB|31|34|我若因大大惧怕众人， 又因宗族的藐视而恐惧， 以致我缄默不言，闭门不出；
JOB|31|35|惟愿有一位肯听我！ 看哪，我的记号，愿全能者回答我！ 愿那与我争讼的写下状词！
JOB|31|36|我必把它带在肩上， 绑在头上为冠冕。
JOB|31|37|我必向上帝述说我脚步的数目， 如同王子进到他面前。
JOB|31|38|“若我的田地喊冤告我， 犁沟也一同哭泣；
JOB|31|39|我若吃地的出产不给银钱， 或叫地的原主丧命；
JOB|31|40|愿蒺藜生长代替麦子， 恶臭的草代替大麦。” 约伯 的话说完了。
JOB|32|1|于是这三个人因 约伯 看自己为义就停止，不再回答他。
JOB|32|2|那时 布西 人， 兰 族 巴拉迦 的儿子 以利户 发怒了。他向 约伯 发怒，因 约伯 自以为义，不以上帝为义。
JOB|32|3|他又向 约伯 的三个朋友发怒，因为他们想不出回答的话来，仍以 约伯 为有罪。
JOB|32|4|以利户 因为他们比自己年老，就等候要与 约伯 说话。
JOB|32|5|以利户 见这三个人口中无话回答，就发怒。
JOB|32|6|布西 人 巴拉迦 的儿子 以利户 回答说： “我年轻，你们年长， 因此我退让，不敢向你们陈述我的意见。
JOB|32|7|我说：‘年长的当先说话； 寿高的当以智慧教导人。’
JOB|32|8|其实，是人里面的灵， 全能者的气使人有聪明。
JOB|32|9|寿高的不都有智慧， 年老的不都明白公平。
JOB|32|10|因此我说：‘你们要听我， 我也要陈述我的意见。’
JOB|32|11|“看哪，我等候你们的话， 侧耳听你们的高见； 直到你们找到要说的言语。
JOB|32|12|我留心听你们， 看哪，你们中间无一人能折服 约伯 ， 回答他的话。
JOB|32|13|你们切不可说：‘我们寻得智慧； 上帝能胜他 ，人却不能。’
JOB|32|14|约伯 没有用言语与我争辩； 我也不用你们的话回答他。
JOB|32|15|“他们惊惶不再回答， 一言不发。
JOB|32|16|我岂因他们不说话， 因他们站住不再回答，仍旧等候呢？
JOB|32|17|我也要以我的一番话回答， 我也要陈述我的意见。
JOB|32|18|因为我满怀言语， 我里面的灵激动我。
JOB|32|19|看哪，我的肚腹如酒囊没有气孔， 又如新皮袋 快要破裂。
JOB|32|20|我要说话，使我舒畅； 我要张开嘴唇回答。
JOB|32|21|我必不看人的情面， 也不奉承人。
JOB|32|22|我不懂得奉承； 不然，造我的主必快快除灭我。”
JOB|33|1|“但是， 约伯 啊，请听我的言语， 侧耳听我一切的话。
JOB|33|2|看哪，我开口， 我的舌在上膛发言。
JOB|33|3|我的言语要表明心中的正直， 我嘴唇所知道的就诚实地说。
JOB|33|4|上帝的灵造了我， 全能者的气使我得生。
JOB|33|5|你若能够，就请回答我； 请你站起来，在我面前陈明。
JOB|33|6|看哪，我在上帝面前与你一样， 也是用泥土造成的。
JOB|33|7|看哪，我不用威严恐吓你， 也不用势力重压你。
JOB|33|8|“其实，你向我耳朵说话， 我听见你言语的声音：
JOB|33|9|‘我是纯洁无过的， 我是无辜的，在我里面没有罪孽。
JOB|33|10|看哪，上帝找机会攻击我， 以我为他的仇敌，
JOB|33|11|把我的脚锁上木枷， 察看我一切的道路。’
JOB|33|12|“看哪，你这话无理，我要回答你， 因上帝比世人更大。
JOB|33|13|你为何与他争论： ‘他任何事都不向人解答’？
JOB|33|14|上帝说一次、两次， 人却不理会。
JOB|33|15|世人在床上沉睡安眠时， 在梦中和夜间的异象里，
JOB|33|16|上帝就开通世人的耳朵， 把警告印在他们心上 ，
JOB|33|17|好叫人转离自己的行为， 叫壮士远离骄傲，
JOB|33|18|拦阻人不陷入地府， 不让他命丧刀下 。
JOB|33|19|“人在床上被疼痛惩治， 骨头不住地挣扎，
JOB|33|20|以致生命厌弃食物， 心中厌恶美味。
JOB|33|21|他的肉消瘦，难以看见； 先前看不见的骨头都凸出来。
JOB|33|22|他的性命临近地府， 他的生命挨近灭命者。
JOB|33|23|一千天使中， 若有一个作传话的临到他， 指示人所当行的事，
JOB|33|24|上帝就施恩给他，说： ‘要救赎他 免得下入地府， 我已经得了赎价。
JOB|33|25|他的肉要比孩童的肉更嫩； 他就返老还童。’
JOB|33|26|他向上帝祷告，上帝就悦纳他； 他必欢呼朝见上帝的面， 因上帝恢复他的义。
JOB|33|27|他在人前歌唱说： ‘我犯了罪，颠倒是非， 却没有受该得的报应。
JOB|33|28|上帝救赎我的性命免入地府， 我的生命也必见光。’
JOB|33|29|“看哪，上帝两次、三次 向人行这一切的事，
JOB|33|30|为要从地府救回人的性命， 使他被生命之光照耀。
JOB|33|31|约伯 啊，你当留心听我； 不要作声，我要说话。
JOB|33|32|你若有话说，可以回答我； 你只管说，因我愿以你为义。
JOB|33|33|若不然，你当听我； 不要作声，我要把智慧教导你。”
JOB|34|1|以利户 继续说：
JOB|34|2|“你们智慧人要听我的言语， 有知识的人要侧耳听我。
JOB|34|3|因为耳朵辨别言语， 好像上膛品尝食物。
JOB|34|4|我们当选择公理， 彼此知道何为善。
JOB|34|5|约伯 曾说：‘我是公义的， 上帝夺去我的公理。
JOB|34|6|我有理，岂能说谎呢？ 我无过，受的箭伤却不能医治。’
JOB|34|7|哪一个人像 约伯 ， 喝讥诮如同喝水呢？
JOB|34|8|他与作恶的结伴， 和恶人同行。
JOB|34|9|他说：‘人以上帝为乐， 总是无益。’
JOB|34|10|“所以，你们明理的人要听我， 上帝断不致行恶， 全能者断不致不义。
JOB|34|11|他必按人所做的报应人， 使各人照所行的得报。
JOB|34|12|确实地，上帝必不作恶， 全能者必不偏离公平。
JOB|34|13|谁派他治理大地？ 谁安定全世界呢？
JOB|34|14|他若专心为己， 将灵和气收归自己，
JOB|34|15|凡血肉之躯必一同死亡； 世人必归于尘土。
JOB|34|16|“你若明理，当听这话， 侧耳听我言语的声音。
JOB|34|17|难道恨恶公平的可以掌权吗？ 那有公义、有大能的，你岂可定他有罪呢？
JOB|34|18|你会对君王说：‘你是卑鄙的’； 对贵族说：‘你们是邪恶的’吗？
JOB|34|19|他待王子不徇情面， 也不看重富足的过于贫寒的， 因为他们都是他手所造的。
JOB|34|20|一瞬间他们就死亡。 百姓在半夜中被震动而去世； 有权力的被夺去，非藉人手。
JOB|34|21|“上帝的眼目观看人的道路， 察看他每一脚步。
JOB|34|22|没有黑暗，没有死荫， 能给作恶者在那里藏身。
JOB|34|23|上帝不必再三传人 到他面前受审判。
JOB|34|24|他毋须调查就粉碎有大能的人， 指定别人代替他们。
JOB|34|25|所以他知道他们的行为， 使他们在夜间倾倒压碎。
JOB|34|26|他在众目睽睽下击打他们， 如同击打恶人。
JOB|34|27|因为他们转离不跟从他， 不留心他一切的道，
JOB|34|28|甚至使贫寒人的哀声达到他那里； 他也听了困苦人的哀声。
JOB|34|29|他安静，谁能定罪呢？ 他转脸，谁能见他呢？ 无论一国或一人都是如此。
JOB|34|30|不虔敬的人不得作王， 免得百姓陷入圈套。
JOB|34|31|“有谁对上帝说： ‘我受了责罚，必不再犯罪；
JOB|34|32|我所看不明的，求你指教我； 我若行了不义，必不再行’？
JOB|34|33|他因你拒绝不接受， 就随你的心愿施行报应吗？ 选择的是你，不是我。 你所知道的，只管说吧！
JOB|34|34|明理的人必对我说， 听我的智慧人也说：
JOB|34|35|‘ 约伯 说话没有知识， 他的言语毫无智慧。’
JOB|34|36|愿 约伯 被考验到底， 因他回答像恶人一样。
JOB|34|37|他在罪上又加悖逆； 在我们中间引起疑惑 ， 用许多言语轻慢上帝。”
JOB|35|1|以利户 继续说：
JOB|35|2|“你以为这话有理， 说：‘我在上帝面前是公义的。’
JOB|35|3|你说：‘这对你有什么益处？ 我不犯罪有什么好处呢？’
JOB|35|4|至于我，我要用言语回答你 和跟你一起的朋友。
JOB|35|5|你要向天观看， 瞻望那高于你的穹苍。
JOB|35|6|你若犯罪，能使上帝受何害呢？ 你的过犯加增，能使上帝受何损呢？
JOB|35|7|你若是公义，能加增他什么呢？ 他从你手里还接受什么呢？
JOB|35|8|你的罪恶只影响像你这类的人； 你的公义也只影响世人。
JOB|35|9|“人因多受欺压就哀求， 因强权者的膀臂而求救。
JOB|35|10|但无人说：‘造我的上帝在哪里？ 他使人夜间歌唱，
JOB|35|11|教导我们多过地上的走兽， 使我们比空中的飞鸟更聪明。’
JOB|35|12|因为恶人骄傲， 他们在那里呼求，他却不回答。
JOB|35|13|虚妄的呼求，上帝必不垂听； 全能者必不留意。
JOB|35|14|何况你说，你不得见他。 案件就在他面前，你等候他吧。
JOB|35|15|但如今因他未曾发怒降罚， 也一点都不理会狂傲，
JOB|35|16|所以 约伯 开口说虚妄的话， 多多发表无知识的言语。”
JOB|36|1|以利户 继续说：
JOB|36|2|“你再给我片时，我就指示你， 因我还有话要为上帝说。
JOB|36|3|我要把我的知识从远处引来， 我要将公义归给造我的主。
JOB|36|4|我的言语绝不虚假， 有全备知识的与你同在。
JOB|36|5|“看哪，上帝有大能，并不藐视人； 他的心智能力广大。
JOB|36|6|他不让恶人活着， 却为困苦人伸冤。
JOB|36|7|他的眼目不远离义人， 却使他们和君王同坐宝座， 永远被高举 。
JOB|36|8|他们若被锁链捆住， 被苦难的绳索缠住，
JOB|36|9|他就向他们指示他们的作为和过犯， 以及他们的狂妄自大。
JOB|36|10|他也开通他们的耳朵来领受教导， 吩咐他们回转离开罪孽。
JOB|36|11|他们若听从事奉他， 就必度日亨通， 历年享福。
JOB|36|12|他们若不听从，就要被刀杀灭， 无知无识而死。
JOB|36|13|“那心中不敬虔的人积蓄怒气； 上帝捆绑他们，他们竟不求救。
JOB|36|14|他们必在青年时死亡， 与神庙娼妓一样丧命。
JOB|36|15|上帝藉着困苦救拔困苦人， 藉所受的欺压开通他们的耳朵。
JOB|36|16|上帝也必引你脱离患难， 进入宽阔不狭窄之地； 摆在你席上的必满有肥甘。
JOB|36|17|“但你充满着恶人的辩辞， 辩辞和审判抓住你。
JOB|36|18|不可让愤怒触动你，使你破口谩骂 ； 也不可因赎价大而偏行。
JOB|36|19|你的呼求 和一切的势力， 果真有用，使你不遭患难吗？
JOB|36|20|不要切慕黑夜， 就是众民在本处被除灭的时候。
JOB|36|21|你要谨慎，不可偏向罪孽， 因你选择罪孽过于苦难。
JOB|36|22|看哪，上帝因他的能力而崇高； 有谁像他那样作教师呢？
JOB|36|23|谁派定他的道路呢？ 谁能说：‘你行了不义’？
JOB|36|24|“你要记得颂赞他的作为， 就是人所歌颂的。
JOB|36|25|他的作为，万人都看见； 世人也从远处观看。
JOB|36|26|看哪，上帝崇高，我们不能知道； 他的年数，不能测度。
JOB|36|27|因他吸取水点， 水点就从云雾中变成雨；
JOB|36|28|云彩将雨落下， 沛然降于世人。
JOB|36|29|又有谁能明白密云如何铺张， 和上帝行宫的雷声呢？
JOB|36|30|看哪，他的亮光普照自己的四围； 他覆盖海的深处。
JOB|36|31|因他用这些审判 众民， 又赐丰富的粮食。
JOB|36|32|他以闪电遮手掌， 命令它击中靶子。
JOB|36|33|所发的雷声将他显明， 牲畜也指明要起暴风 。”
JOB|37|1|“因此我心战兢， 从原处移动。
JOB|37|2|听啊，听他轰轰的声音， 是上帝口中所发的响声。
JOB|37|3|他发响声震遍天下， 他的闪电直到地极。
JOB|37|4|随后，人听见他的声音， 是那轰轰的声音； 他发出威严的雷声， 而不加以遏止。
JOB|37|5|上帝发出奇妙的雷声； 他行大事，我们不能测透。
JOB|37|6|他对雪说：‘要降在地上’； 对大雨和暴雨也是这样说。
JOB|37|7|他封住各人的手， 叫所造的万人都知道他的作为。
JOB|37|8|野兽进入穴中， 卧在自己洞内。
JOB|37|9|暴风来自内宫， 寒冷出于狂风。
JOB|37|10|上帝嘘气成冰， 凝结宽阔之水，
JOB|37|11|使密云盛满水气， 乌云散布闪电。
JOB|37|12|云藉着他的指引游行旋转， 在世界的地面上行他一切所吩咐的，
JOB|37|13|或为责罚，或为他的地， 或为慈爱，都是他所行的。
JOB|37|14|“ 约伯 啊，侧耳听这话， 要站立，思想上帝奇妙的作为。
JOB|37|15|你知道上帝如何安排这些， 如何使云中的闪电照耀吗？
JOB|37|16|你知道云彩如何浮于空中， 知识全备者奇妙的作为吗？
JOB|37|17|你知道南风使地寂静， 你的衣服就变为热吗？
JOB|37|18|你岂能与上帝同铺穹苍， 坚固如同铸成的镜子吗？
JOB|37|19|我们因在黑暗中，不会陈说， 请你指教我们该对他说什么。
JOB|37|20|有人告诉他我要说话吗？ 岂有人说他愿被吞灭吗？
JOB|37|21|“现在，人不得见穹苍的亮光； 风一吹过，天色晴朗。
JOB|37|22|金色的光辉来自北方， 在上帝那里有可畏的威严。
JOB|37|23|全能者，我们不能测度； 他大有能力，又有公平， 满有公义，必不苦待人。
JOB|37|24|所以，世人敬畏他； 凡自以为 有智慧的，他都不看顾。”
JOB|38|1|那时，耶和华从旋风中回答 约伯 说：
JOB|38|2|“谁用无知的言语使我的旨意暗昧不明？
JOB|38|3|你要如勇士束腰； 我问你，你可以让我知道。
JOB|38|4|“我立大地根基的时候，你在哪里？ 你若明白事理，只管说吧！
JOB|38|5|你知道是谁定地的尺度， 是谁把准绳拉在其上吗？
JOB|38|6|地的根基安置在何处？ 地的角石是谁安放的？
JOB|38|7|那时，晨星一同歌唱； 上帝的众使者也都欢呼。
JOB|38|8|“当海水冲出，如出母胎， 谁用门将它关闭呢？
JOB|38|9|是我用云彩当海的衣服， 用幽暗当包裹它的布，
JOB|38|10|为它定界限， 又安门和闩，
JOB|38|11|说：‘你只可到这里，不可越过； 你狂傲的浪要到此止住。’
JOB|38|12|“你有生以来，曾命定晨光， 曾使黎明知道自己的地位，
JOB|38|13|抓住地的四极， 把恶人从其中驱逐出来吗？
JOB|38|14|地改变如泥上盖印， 万物出现如衣服一样。
JOB|38|15|亮光不照恶人， 高举的膀臂也必折断。
JOB|38|16|“你曾进到海之源， 或在深渊的隐密处行走吗？
JOB|38|17|死亡的门曾向你显露吗？ 死荫的门你曾见过吗？
JOB|38|18|地的广大，你能测透吗？ 你若全知道，只管说吧！
JOB|38|19|“往光明居所的路在哪里？ 黑暗的地方在何处？
JOB|38|20|你能将它带到其领域， 能辨明其居所之路吗？
JOB|38|21|你知道的，因为那时你已出生， 你活的日子数目也多。
JOB|38|22|“你曾进入雪之库， 或见过雹的仓吗？
JOB|38|23|雪雹是我为灾难的时候， 为打仗和战争的日子所预备。
JOB|38|24|光亮从何路分开？ 东风从何路分散遍地？
JOB|38|25|“谁为大雨分道， 谁为雷电开路，
JOB|38|26|使雨降在无人之地， 在无人居住的旷野，
JOB|38|27|使荒废凄凉之地得以丰足， 青草得以生长？
JOB|38|28|“雨有父亲吗？ 露珠是谁生的呢？
JOB|38|29|冰出于谁的胎？ 天上的霜是谁生的呢？
JOB|38|30|诸水坚硬如石头， 深渊之面凝结成冰。
JOB|38|31|“你能为昴星系结吗？ 你能为参星解带吗？
JOB|38|32|你能按时领出星宿吗？ 能引导北斗与其众星吗？
JOB|38|33|你知道天的定律吗？ 你能使地归其权下吗？
JOB|38|34|“你能向密云扬起声来， 使倾盆的雨遮盖你吗？
JOB|38|35|你能发出闪电，使它们 行走， 并对你说：‘我们在这里’吗？
JOB|38|36|谁将智慧放在朱鹭 中？ 谁将聪明赐给雄鸡 ？
JOB|38|37|谁能用智慧数算云彩？ 谁能倾倒天上的瓶呢？
JOB|38|38|那时，尘土聚集成团， 土块紧紧结连。
JOB|38|39|“你能为母狮抓取猎物， 使少壮的狮子饱足吗？
JOB|38|40|那时，它们在洞中蹲伏， 在隐密处埋伏。
JOB|38|41|谁能为乌鸦预备食物呢？ 那时，乌鸦之雏哀求上帝， 因无食物飞来飞去。”
JOB|39|1|“你知道岩石间的野山羊几时生产吗？ 你能观察母鹿下小鹿吗？
JOB|39|2|你能数算它们怀胎的月数吗？ 你知道它们几时生产吗？
JOB|39|3|它们屈身，生下幼儿， 就解除了阵痛。
JOB|39|4|其子渐渐肥壮，在荒野长大； 它们出去，不再归回。
JOB|39|5|“谁放野驴自由？ 谁解开快驴的绳索？
JOB|39|6|我使旷野作它的住处， 使盐地当它的居所。
JOB|39|7|它嘲笑城内的喧嚷， 不听赶牲口的喝声。
JOB|39|8|诸山是它漫游的草场， 它寻找各样青绿之物。
JOB|39|9|“野牛岂肯服事你？ 岂肯在你的槽旁过夜？
JOB|39|10|你岂能用套绳将野牛系于犁沟？ 它岂肯随你耙松山谷之地？
JOB|39|11|你岂可因它力大就倚靠它？ 岂可把你的工交给它做呢？
JOB|39|12|你岂能靠它把你的谷物运回， 又收聚在你的禾场上吗？
JOB|39|13|“鸵鸟的翅膀欢然拍动， 但岂是鹳的翎毛和羽毛吗 ？
JOB|39|14|因它把蛋留在地上， 使蛋在尘土中得温暖，
JOB|39|15|却忘记脚会把蛋踹碎， 野兽会践踏它。
JOB|39|16|它粗暴待雏，似乎不是自己生的； 虽徒然劳苦 ，也不惧怕。
JOB|39|17|因为上帝使它忘记智慧， 也未将悟性分给它。
JOB|39|18|它几时挺身展开翅膀， 就嘲笑马和骑马的人。
JOB|39|19|“马的力量是你所赐的吗？ 它颈项上的鬃是你披上的吗？
JOB|39|20|是你叫它跳跃像蝗虫吗？ 它喷气之威严使人惊惶。
JOB|39|21|它用蹄在谷中挖地 ，以能力欢跃； 它出去迎击仇敌 。
JOB|39|22|它嘲笑惧怕，并不惊惶， 也不因刀剑退却。
JOB|39|23|箭袋在它身上铮铮有声， 枪和短枪闪闪发亮。
JOB|39|24|它震颤激动，将地吞下 ； 一听角声就站不住。
JOB|39|25|每逢角声一响，它说：‘啊哈！’ 它从远处闻到战争的气息， 听见军官如雷的吼声和呐喊。
JOB|39|26|“鹰展开翅膀向南飞翔， 岂是藉着你的智慧吗？
JOB|39|27|大鹰上腾在高处搭窝， 岂是听你的指示吗？
JOB|39|28|它住在山岩， 以山峰和坚固之所为家，
JOB|39|29|从那里窥察食物， 眼睛自远方了望。
JOB|39|30|它的雏吸血； 被杀的人在哪里，它也在哪里。”
JOB|40|1|耶和华继续对 约伯 说：
JOB|40|2|“强辩的岂可与全能者争论？ 与上帝辩驳的可以回答吧！”
JOB|40|3|于是， 约伯 回答耶和华说：
JOB|40|4|“看哪，我是卑贱的！我用什么回答你呢？ 我只好用手捂住我的口。
JOB|40|5|我说了一次，就不回答； 说了两次，不再说了。”
JOB|40|6|于是，耶和华从旋风中回答 约伯 说：
JOB|40|7|“你要如勇士束腰； 我问你，你可以让我知道。
JOB|40|8|你岂可废弃我的判断？ 岂可定我有罪，好显自己为义吗？
JOB|40|9|你有上帝那样的膀臂吗？ 你能像他那样发雷声吗？
JOB|40|10|“你要以荣耀庄严为妆饰， 以尊荣威严为衣服。
JOB|40|11|你要发出你满溢的怒气， 见一切骄傲的人，使他降卑；
JOB|40|12|你见一切骄傲的人，将他制伏， 把恶人践踏在原来地方。
JOB|40|13|你将他们一同埋藏在尘土中， 把他们的脸遮蔽在隐密处 。
JOB|40|14|这样，我也向你承认， 你的右手能救你自己。
JOB|40|15|“看哪，我造河马， 也造了你； 它吃草像牛一样。
JOB|40|16|看哪，它的力气在腰间， 能力在肚腹的肌肉上。
JOB|40|17|它挺直 尾巴如香柏树， 它大腿的筋紧密结合。
JOB|40|18|它的骨头好像铜管； 它的肢体仿佛铁棍。
JOB|40|19|“它在上帝所造之物中为首， 只有创造它的能携刀临近它。
JOB|40|20|诸山为它产出食物， 百兽也在那里游玩。
JOB|40|21|它伏在莲叶之下， 在芦苇和沼泽的隐密处。
JOB|40|22|莲叶的阴影遮蔽它， 溪旁的柳树环绕它。
JOB|40|23|看哪，河水泛滥，它不慌张； 连 约旦河 涨到它口边，它也安然自若。
JOB|40|24|谁能在它眼前捉拿它呢？ 谁能以圈套穿它鼻子呢？”
JOB|41|1|“你能用鱼钩钓上 力威亚探 吗？ 能用绳子压下它的舌头吗？
JOB|41|2|你能用绳索穿它的鼻子吗？ 能用钩子穿它的腮骨吗？
JOB|41|3|它岂向你连连恳求， 向你说温柔的话吗？
JOB|41|4|它岂肯与你立约， 让你拿它永远作奴仆吗？
JOB|41|5|你岂可拿它当雀鸟玩耍？ 岂可将它系来给你幼女？
JOB|41|6|合伙的鱼贩岂可拿它当货物？ 他们岂可把它分给商人呢？
JOB|41|7|你能用倒钩扎满它的皮， 能用鱼叉叉满它的头吗？
JOB|41|8|把你的手掌按在它身上吧！ 想一想与它搏斗，你就不再这样做了！
JOB|41|9|看哪，对它有指望是徒然的； 一见它，岂不也丧胆吗？
JOB|41|10|没有那么凶猛的人敢惹它。 这样，谁能在我面前站立得住呢？
JOB|41|11|谁能与我对质，使我偿还呢？ 天下万物都是我的。
JOB|41|12|“我不能缄默不提 它的肢体和力量，以及健美的骨骼。
JOB|41|13|谁能剥它的外皮？ 谁能进它的铠甲之间 呢？
JOB|41|14|谁能开它的腮颊？ 它牙齿的四围是可畏的。
JOB|41|15|它的背上有一排排的鳞甲 ， 紧紧闭合，封得严密。
JOB|41|16|这鳞甲一一相连， 气不得透入其间，
JOB|41|17|互相连接， 胶结一起，不能分开。
JOB|41|18|它打喷嚏就发出光来， 它的眼睛好像晨曦 。
JOB|41|19|从它口中发出烧着的火把， 有火星飞迸出来；
JOB|41|20|从它鼻孔冒出烟来， 如烧开的锅在沸腾 。
JOB|41|21|它的气点着煤炭， 有火焰从它口中发出。
JOB|41|22|它颈项中存着劲力， 恐惧在它面前蹦跳。
JOB|41|23|它的肉块紧紧结连， 紧贴其身，不能摇动。
JOB|41|24|它的心结实如石头， 如下面的磨石那样结实。
JOB|41|25|它一起来，神明都恐惧， 因崩溃而惊慌失措。
JOB|41|26|人用刀剑扎它，是无用的， 枪、标枪、尖枪也一样。
JOB|41|27|它以铁为干草， 以铜为烂木。
JOB|41|28|箭不能使它逃走， 它看弹石如碎秸。
JOB|41|29|它当棍棒作碎秸， 它嘲笑短枪的飕飕声。
JOB|41|30|它肚腹下面是尖瓦片； 它如钉耙刮过淤泥。
JOB|41|31|它使深渊滚沸如锅， 使海洋如锅中膏油。
JOB|41|32|它使走过以后的路发光， 令人觉得深渊如同白发。
JOB|41|33|尘世上没有像它那样的受造物， 一无所惧。
JOB|41|34|凡高大的，它盯着看； 它在一切狂傲的野兽中作王。”
JOB|42|1|约伯 回答耶和华说：
JOB|42|2|“我知道，你万事都能做； 你的计划不能拦阻。
JOB|42|3|谁无知使你的旨意隐藏呢？ 因此我说的，我不明白； 这些事太奇妙，是我不知道的。
JOB|42|4|求你听我，我要说话； 我问你，求你让我知道。
JOB|42|5|我从前风闻有你， 现在亲眼看见你。
JOB|42|6|因此我撤回 ， 在尘土和炉灰中懊悔。”
JOB|42|7|耶和华对 约伯 说话以后，耶和华就对 提幔 人 以利法 说：“我的怒气向你和你两个朋友发作，因为你们议论我，不如我的仆人 约伯 说的正确。
JOB|42|8|现在你们要为自己取七头公牛，七只公羊，到我的仆人 约伯 那里去，为自己献上燔祭，我的仆人 约伯 就为你们祈祷。我必悦纳他，不按你们的愚妄处置你们。你们议论我，不如我的仆人 约伯 说的正确。”
JOB|42|9|于是 提幔 人 以利法 、 书亚 人 比勒达 、 拿玛 人 琐法 遵照耶和华所吩咐的去做，耶和华就悦纳 约伯 。
JOB|42|10|约伯 为他的朋友祈祷。耶和华就使 约伯 从苦境 中转回，并且耶和华赐给他的比他从前所有的加倍。
JOB|42|11|约伯 的兄弟、姊妹，和以前所认识的人都来到他那里，在他家里跟他一同吃饭。他们因耶和华所降于他的一切灾祸，都为他悲伤，安慰他。每人送他一块可锡塔 和一个金环。
JOB|42|12|这样，耶和华后来赐福给 约伯 比先前更多。他有一万四千只羊，六千匹骆驼，一千对牛，一千匹母驴。
JOB|42|13|他也有七个儿子，三个女儿。
JOB|42|14|他给长女起名叫 耶米玛 ，次女叫 基洗亚 ，三女叫 基连哈朴 。
JOB|42|15|在全地的妇女中找不着像 约伯 的女儿那样美貌的。她们的父亲使她们在兄弟中得产业。
JOB|42|16|此后， 约伯 又活了一百四十年，得见他的四代儿孙。
JOB|42|17|这样， 约伯 年纪老迈，日子满足而死。
