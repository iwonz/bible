HAG|1|1|大流士 王第二年六月初一，耶和華的話藉 哈該 先知向 撒拉鐵 的兒子 猶大 省長 所羅巴伯 和 約撒答 的兒子 約書亞 大祭司傳講，說：
HAG|1|2|「萬軍之耶和華如此說，這百姓說，建造耶和華殿的時候還沒有到 。」
HAG|1|3|耶和華的話藉 哈該 先知傳講，說：
HAG|1|4|「這殿荒涼，你們自己還住天花板的房屋嗎？
HAG|1|5|現在，萬軍之耶和華如此說，你們要省察自己的行為。
HAG|1|6|你們撒的種多，收的卻少；你們吃，卻不得飽；喝，卻不得足；穿衣服，卻不得暖；領工錢的，領了工錢卻裝入有破洞的袋中。
HAG|1|7|「萬軍之耶和華如此說，你們要省察自己的行為。
HAG|1|8|你們要上山取木料，建造這殿，我就因此喜樂，且得榮耀。這是耶和華說的。
HAG|1|9|你們盼望多得，看哪，所得的卻少；你們收到家中，我就吹去。這是為甚麼呢？因為我的殿荒涼，你們各人卻只為自己的房屋奔走。這是萬軍之耶和華說的。
HAG|1|10|所以，因你們的緣故 ，天不降甘露，地也不出土產。
HAG|1|11|我命令乾旱臨到土地、山岡、五穀、新酒、新油和地上的出產，也臨到人和牲畜，以及一切人手勞碌得來的。」
HAG|1|12|那時， 撒拉鐵 的兒子 所羅巴伯 、 約撒答 的兒子 約書亞 大祭司，和所有倖存的百姓都聽從耶和華－他們上帝的話，就是 哈該 先知奉耶和華－他們上帝差遣所說的話；百姓在耶和華面前存敬畏的心。
HAG|1|13|耶和華的使者 哈該 奉耶和華差遣對百姓說：「我與你們同在。這是耶和華說的。」
HAG|1|14|耶和華激發 撒拉鐵 的兒子 猶大 省長 所羅巴伯 、 約撒答 的兒子 約書亞 大祭司，和所有倖存百姓的心，他們就來為萬軍之耶和華－他們上帝的殿做工。
HAG|1|15|這是在 大流士 王第二年六月二十四日。
HAG|2|1|七月二十一日，耶和華的話藉 哈該 先知傳講，說：
HAG|2|2|「你要曉諭 撒拉鐵 的兒子 猶大 省長 所羅巴伯 、 約撒答 的兒子 約書亞 大祭司，和所有倖存的百姓，說：
HAG|2|3|『你們中間存留的，有誰見過這殿從前的榮耀呢？現在你們看如何？在你們眼中豈不是如同無有嗎？
HAG|2|4|所羅巴伯 啊，現在，你當剛強！這是耶和華說的。 約撒答 的兒子 約書亞 大祭司啊，你當剛強！這是耶和華說的。這地的百姓啊，你們都當剛強做工，因為我與你們同在。這是萬軍之耶和華說的。
HAG|2|5|這是照著你們出 埃及 時我與你們立約的話。我的靈仍要住在你們中間，你們不必懼怕。
HAG|2|6|萬軍之耶和華如此說：過些時候，我必再一次震動天地、滄海與乾地。
HAG|2|7|我必震動萬國，萬國的珍寶都必運來 ，我就使這殿充滿榮耀。這是萬軍之耶和華說的。
HAG|2|8|銀子是我的，金子也是我的。這是萬軍之耶和華說的。
HAG|2|9|這後來的殿的榮耀必大過先前的榮耀。這是萬軍之耶和華說的。在這地方我必賜平安。這是萬軍之耶和華說的。』」
HAG|2|10|大流士 王第二年九月二十四日，耶和華的話臨到 哈該 先知，說：
HAG|2|11|「萬軍之耶和華如此說，你要向祭司請教律法，說：
HAG|2|12|『看哪，若有人用衣服的邊兜聖肉，這衣服的邊接觸了餅，或湯，或酒，或油，或別的食物，這些是否成為聖呢？』」祭司回答說：「不。」
HAG|2|13|哈該 又說：「若有人因摸屍體染了不潔淨，然後接觸任何東西，這東西就變為不潔淨嗎？」祭司回答說：「必不潔淨。」
HAG|2|14|於是 哈該 說：「耶和華說，在我面前這民如此，這國也是如此；他們手裏的各樣工作都是如此；他們在那裏所獻的都不潔淨。」
HAG|2|15|「現在，你們心裏要想一想，從今日起，耶和華的殿還沒有一塊石頭放在石頭上的情況。
HAG|2|16|那時你們怎麼了？ 有人來到二十斗的穀堆那裏，卻只得了十斗；有人來到酒池那裏要取五十桶，卻只得了二十桶。
HAG|2|17|我以焚風 、霉爛、冰雹攻擊你們，和你們手上的各樣工作，你們仍不歸向我。這是耶和華說的。
HAG|2|18|你們心裏要想一想，從今日起，就是從這九月二十四日起，從立耶和華殿根基的日子起，你們心裏想一想：
HAG|2|19|倉裏還有穀種嗎？葡萄樹、無花果樹、石榴樹、橄欖樹雖沒有結果子， 從今日起，我必賜福。」
HAG|2|20|這月二十四日，耶和華的話再次臨到 哈該 ，說：
HAG|2|21|「你要告訴 猶大 省長 所羅巴伯 說，我必震動天地，
HAG|2|22|傾覆列國的寶座，除滅列邦列國的勢力，並傾覆戰車和坐在其上的。馬和騎兵都必跌倒，各人被弟兄的刀所殺。
HAG|2|23|萬軍之耶和華說： 撒拉鐵 的兒子我僕人 所羅巴伯 啊，這是耶和華說的，到那日，我必以你為印，因我揀選了你。這是萬軍之耶和華說的。」
