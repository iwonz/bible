ECCL|1|1|The words of the Preacher, the son of David, king in Jerusalem.
ECCL|1|2|Vanity of vanities, saith the Preacher, vanity of vanities; all is vanity.
ECCL|1|3|What profit hath a man of all his labour which he taketh under the sun?
ECCL|1|4|One generation passeth away, and another generation cometh: but the earth abideth for ever.
ECCL|1|5|The sun also ariseth, and the sun goeth down, and hasteth to his place where he arose.
ECCL|1|6|The wind goeth toward the south, and turneth about unto the north; it whirleth about continually, and the wind returneth again according to his circuits.
ECCL|1|7|All the rivers run into the sea; yet the sea is not full; unto the place from whence the rivers come, thither they return again.
ECCL|1|8|All things are full of labour; man cannot utter it: the eye is not satisfied with seeing, nor the ear filled with hearing.
ECCL|1|9|The thing that hath been, it is that which shall be; and that which is done is that which shall be done: and there is no new thing under the sun.
ECCL|1|10|Is there any thing whereof it may be said, See, this is new? it hath been already of old time, which was before us.
ECCL|1|11|There is no remembrance of former things; neither shall there be any remembrance of things that are to come with those that shall come after.
ECCL|1|12|I the Preacher was king over Israel in Jerusalem.
ECCL|1|13|And I gave my heart to seek and search out by wisdom concerning all things that are done under heaven: this sore travail hath God given to the sons of man to be exercised therewith.
ECCL|1|14|I have seen all the works that are done under the sun; and, behold, all is vanity and vexation of spirit.
ECCL|1|15|That which is crooked cannot be made straight: and that which is wanting cannot be numbered.
ECCL|1|16|I communed with mine own heart, saying, Lo, I am come to great estate, and have gotten more wisdom than all they that have been before me in Jerusalem: yea, my heart had great experience of wisdom and knowledge.
ECCL|1|17|And I gave my heart to know wisdom, and to know madness and folly: I perceived that this also is vexation of spirit.
ECCL|1|18|For in much wisdom is much grief: and he that increaseth knowledge increaseth sorrow.
ECCL|2|1|I said in mine heart, Go to now, I will prove thee with mirth, therefore enjoy pleasure: and, behold, this also is vanity.
ECCL|2|2|I said of laughter, It is mad: and of mirth, What doeth it?
ECCL|2|3|I sought in mine heart to give myself unto wine, yet acquainting mine heart with wisdom; and to lay hold on folly, till I might see what was that good for the sons of men, which they should do under the heaven all the days of their life.
ECCL|2|4|I made me great works; I builded me houses; I planted me vineyards:
ECCL|2|5|I made me gardens and orchards, and I planted trees in them of all kind of fruits:
ECCL|2|6|I made me pools of water, to water therewith the wood that bringeth forth trees:
ECCL|2|7|I got me servants and maidens, and had servants born in my house; also I had great possessions of great and small cattle above all that were in Jerusalem before me:
ECCL|2|8|I gathered me also silver and gold, and the peculiar treasure of kings and of the provinces: I gat me men singers and women singers, and the delights of the sons of men, as musical instruments, and that of all sorts.
ECCL|2|9|So I was great, and increased more than all that were before me in Jerusalem: also my wisdom remained with me.
ECCL|2|10|And whatsoever mine eyes desired I kept not from them, I withheld not my heart from any joy; for my heart rejoiced in all my labour: and this was my portion of all my labour.
ECCL|2|11|Then I looked on all the works that my hands had wrought, and on the labour that I had laboured to do: and, behold, all was vanity and vexation of spirit, and there was no profit under the sun.
ECCL|2|12|And I turned myself to behold wisdom, and madness, and folly: for what can the man do that cometh after the king? even that which hath been already done.
ECCL|2|13|Then I saw that wisdom excelleth folly, as far as light excelleth darkness.
ECCL|2|14|The wise man's eyes are in his head; but the fool walketh in darkness: and I myself perceived also that one event happeneth to them all.
ECCL|2|15|Then said I in my heart, As it happeneth to the fool, so it happeneth even to me; and why was I then more wise? Then I said in my heart, that this also is vanity.
ECCL|2|16|For there is no remembrance of the wise more than of the fool for ever; seeing that which now is in the days to come shall all be forgotten. And how dieth the wise man? as the fool.
ECCL|2|17|Therefore I hated life; because the work that is wrought under the sun is grievous unto me: for all is vanity and vexation of spirit.
ECCL|2|18|Yea, I hated all my labour which I had taken under the sun: because I should leave it unto the man that shall be after me.
ECCL|2|19|And who knoweth whether he shall be a wise man or a fool? yet shall he have rule over all my labour wherein I have laboured, and wherein I have shewed myself wise under the sun. This is also vanity.
ECCL|2|20|Therefore I went about to cause my heart to despair of all the labour which I took under the sun.
ECCL|2|21|For there is a man whose labour is in wisdom, and in knowledge, and in equity; yet to a man that hath not laboured therein shall he leave it for his portion. This also is vanity and a great evil.
ECCL|2|22|For what hath man of all his labour, and of the vexation of his heart, wherein he hath laboured under the sun?
ECCL|2|23|For all his days are sorrows, and his travail grief; yea, his heart taketh not rest in the night. This is also vanity.
ECCL|2|24|There is nothing better for a man, than that he should eat and drink, and that he should make his soul enjoy good in his labour. This also I saw, that it was from the hand of God.
ECCL|2|25|For who can eat, or who else can hasten hereunto, more than I?
ECCL|2|26|For God giveth to a man that is good in his sight wisdom, and knowledge, and joy: but to the sinner he giveth travail, to gather and to heap up, that he may give to him that is good before God. This also is vanity and vexation of spirit.
ECCL|3|1|To every thing there is a season, and a time to every purpose under the heaven:
ECCL|3|2|A time to be born, and a time to die; a time to plant, and a time to pluck up that which is planted;
ECCL|3|3|A time to kill, and a time to heal; a time to break down, and a time to build up;
ECCL|3|4|A time to weep, and a time to laugh; a time to mourn, and a time to dance;
ECCL|3|5|A time to cast away stones, and a time to gather stones together; a time to embrace, and a time to refrain from embracing;
ECCL|3|6|A time to get, and a time to lose; a time to keep, and a time to cast away;
ECCL|3|7|A time to rend, and a time to sew; a time to keep silence, and a time to speak;
ECCL|3|8|A time to love, and a time to hate; a time of war, and a time of peace.
ECCL|3|9|What profit hath he that worketh in that wherein he laboureth?
ECCL|3|10|I have seen the travail, which God hath given to the sons of men to be exercised in it.
ECCL|3|11|He hath made every thing beautiful in his time: also he hath set the world in their heart, so that no man can find out the work that God maketh from the beginning to the end.
ECCL|3|12|I know that there is no good in them, but for a man to rejoice, and to do good in his life.
ECCL|3|13|And also that every man should eat and drink, and enjoy the good of all his labour, it is the gift of God.
ECCL|3|14|I know that, whatsoever God doeth, it shall be for ever: nothing can be put to it, nor any thing taken from it: and God doeth it, that men should fear before him.
ECCL|3|15|That which hath been is now; and that which is to be hath already been; and God requireth that which is past.
ECCL|3|16|And moreover I saw under the sun the place of judgment, that wickedness was there; and the place of righteousness, that iniquity was there.
ECCL|3|17|I said in mine heart, God shall judge the righteous and the wicked: for there is a time there for every purpose and for every work.
ECCL|3|18|I said in mine heart concerning the estate of the sons of men, that God might manifest them, and that they might see that they themselves are beasts.
ECCL|3|19|For that which befalleth the sons of men befalleth beasts; even one thing befalleth them: as the one dieth, so dieth the other; yea, they have all one breath; so that a man hath no preeminence above a beast: for all is vanity.
ECCL|3|20|All go unto one place; all are of the dust, and all turn to dust again.
ECCL|3|21|Who knoweth the spirit of man that goeth upward, and the spirit of the beast that goeth downward to the earth?
ECCL|3|22|Wherefore I perceive that there is nothing better, than that a man should rejoice in his own works; for that is his portion: for who shall bring him to see what shall be after him?
ECCL|4|1|So I returned, and considered all the oppressions that are done under the sun: and behold the tears of such as were oppressed, and they had no comforter; and on the side of their oppressors there was power; but they had no comforter.
ECCL|4|2|Wherefore I praised the dead which are already dead more than the living which are yet alive.
ECCL|4|3|Yea, better is he than both they, which hath not yet been, who hath not seen the evil work that is done under the sun.
ECCL|4|4|Again, I considered all travail, and every right work, that for this a man is envied of his neighbour. This is also vanity and vexation of spirit.
ECCL|4|5|The fool foldeth his hands together, and eateth his own flesh.
ECCL|4|6|Better is an handful with quietness, than both the hands full with travail and vexation of spirit.
ECCL|4|7|Then I returned, and I saw vanity under the sun.
ECCL|4|8|There is one alone, and there is not a second; yea, he hath neither child nor brother: yet is there no end of all his labour; neither is his eye satisfied with riches; neither saith he, For whom do I labour, and bereave my soul of good? This is also vanity, yea, it is a sore travail.
ECCL|4|9|Two are better than one; because they have a good reward for their labour.
ECCL|4|10|For if they fall, the one will lift up his fellow: but woe to him that is alone when he falleth; for he hath not another to help him up.
ECCL|4|11|Again, if two lie together, then they have heat: but how can one be warm alone?
ECCL|4|12|And if one prevail against him, two shall withstand him; and a threefold cord is not quickly broken.
ECCL|4|13|Better is a poor and a wise child than an old and foolish king, who will no more be admonished.
ECCL|4|14|For out of prison he cometh to reign; whereas also he that is born in his kingdom becometh poor.
ECCL|4|15|I considered all the living which walk under the sun, with the second child that shall stand up in his stead.
ECCL|4|16|There is no end of all the people, even of all that have been before them: they also that come after shall not rejoice in him. Surely this also is vanity and vexation of spirit.
ECCL|5|1|Keep thy foot when thou goest to the house of God, and be more ready to hear, than to give the sacrifice of fools: for they consider not that they do evil.
ECCL|5|2|Be not rash with thy mouth, and let not thine heart be hasty to utter any thing before God: for God is in heaven, and thou upon earth: therefore let thy words be few.
ECCL|5|3|For a dream cometh through the multitude of business; and a fool's voice is known by multitude of words.
ECCL|5|4|When thou vowest a vow unto God, defer not to pay it; for he hath no pleasure in fools: pay that which thou hast vowed.
ECCL|5|5|Better is it that thou shouldest not vow, than that thou shouldest vow and not pay.
ECCL|5|6|Suffer not thy mouth to cause thy flesh to sin; neither say thou before the angel, that it was an error: wherefore should God be angry at thy voice, and destroy the work of thine hands?
ECCL|5|7|For in the multitude of dreams and many words there are also divers vanities: but fear thou God.
ECCL|5|8|If thou seest the oppression of the poor, and violent perverting of judgment and justice in a province, marvel not at the matter: for he that is higher than the highest regardeth; and there be higher than they.
ECCL|5|9|Moreover the profit of the earth is for all: the king himself is served by the field.
ECCL|5|10|He that loveth silver shall not be satisfied with silver; nor he that loveth abundance with increase: this is also vanity.
ECCL|5|11|When goods increase, they are increased that eat them: and what good is there to the owners thereof, saving the beholding of them with their eyes?
ECCL|5|12|The sleep of a labouring man is sweet, whether he eat little or much: but the abundance of the rich will not suffer him to sleep.
ECCL|5|13|There is a sore evil which I have seen under the sun, namely, riches kept for the owners thereof to their hurt.
ECCL|5|14|But those riches perish by evil travail: and he begetteth a son, and there is nothing in his hand.
ECCL|5|15|As he came forth of his mother's womb, naked shall he return to go as he came, and shall take nothing of his labour, which he may carry away in his hand.
ECCL|5|16|And this also is a sore evil, that in all points as he came, so shall he go: and what profit hath he that hath laboured for the wind?
ECCL|5|17|All his days also he eateth in darkness, and he hath much sorrow and wrath with his sickness.
ECCL|5|18|Behold that which I have seen: it is good and comely for one to eat and to drink, and to enjoy the good of all his labour that he taketh under the sun all the days of his life, which God giveth him: for it is his portion.
ECCL|5|19|Every man also to whom God hath given riches and wealth, and hath given him power to eat thereof, and to take his portion, and to rejoice in his labour; this is the gift of God.
ECCL|5|20|For he shall not much remember the days of his life; because God answereth him in the joy of his heart.
ECCL|6|1|There is an evil which I have seen under the sun, and it is common among men:
ECCL|6|2|A man to whom God hath given riches, wealth, and honour, so that he wanteth nothing for his soul of all that he desireth, yet God giveth him not power to eat thereof, but a stranger eateth it: this is vanity, and it is an evil disease.
ECCL|6|3|If a man beget an hundred children, and live many years, so that the days of his years be many, and his soul be not filled with good, and also that he have no burial; I say, that an untimely birth is better than he.
ECCL|6|4|For he cometh in with vanity, and departeth in darkness, and his name shall be covered with darkness.
ECCL|6|5|Moreover he hath not seen the sun, nor known any thing: this hath more rest than the other.
ECCL|6|6|Yea, though he live a thousand years twice told, yet hath he seen no good: do not all go to one place?
ECCL|6|7|All the labour of man is for his mouth, and yet the appetite is not filled.
ECCL|6|8|For what hath the wise more than the fool? what hath the poor, that knoweth to walk before the living?
ECCL|6|9|Better is the sight of the eyes than the wandering of the desire: this is also vanity and vexation of spirit.
ECCL|6|10|That which hath been is named already, and it is known that it is man: neither may he contend with him that is mightier than he.
ECCL|6|11|Seeing there be many things that increase vanity, what is man the better?
ECCL|6|12|For who knoweth what is good for man in this life, all the days of his vain life which he spendeth as a shadow? for who can tell a man what shall be after him under the sun?
ECCL|7|1|A good name is better than precious ointment; and the day of death than the day of one's birth.
ECCL|7|2|It is better to go to the house of mourning, than to go to the house of feasting: for that is the end of all men; and the living will lay it to his heart.
ECCL|7|3|Sorrow is better than laughter: for by the sadness of the countenance the heart is made better.
ECCL|7|4|The heart of the wise is in the house of mourning; but the heart of fools is in the house of mirth.
ECCL|7|5|It is better to hear the rebuke of the wise, than for a man to hear the song of fools.
ECCL|7|6|For as the crackling of thorns under a pot, so is the laughter of the fool: this also is vanity.
ECCL|7|7|Surely oppression maketh a wise man mad; and a gift destroyeth the heart.
ECCL|7|8|Better is the end of a thing than the beginning thereof: and the patient in spirit is better than the proud in spirit.
ECCL|7|9|Be not hasty in thy spirit to be angry: for anger resteth in the bosom of fools.
ECCL|7|10|Say not thou, What is the cause that the former days were better than these? for thou dost not enquire wisely concerning this.
ECCL|7|11|Wisdom is good with an inheritance: and by it there is profit to them that see the sun.
ECCL|7|12|For wisdom is a defence, and money is a defence: but the excellency of knowledge is, that wisdom giveth life to them that have it.
ECCL|7|13|Consider the work of God: for who can make that straight, which he hath made crooked?
ECCL|7|14|In the day of prosperity be joyful, but in the day of adversity consider: God also hath set the one over against the other, to the end that man should find nothing after him.
ECCL|7|15|All things have I seen in the days of my vanity: there is a just man that perisheth in his righteousness, and there is a wicked man that prolongeth his life in his wickedness.
ECCL|7|16|Be not righteous over much; neither make thyself over wise: why shouldest thou destroy thyself?
ECCL|7|17|Be not over much wicked, neither be thou foolish: why shouldest thou die before thy time?
ECCL|7|18|It is good that thou shouldest take hold of this; yea, also from this withdraw not thine hand: for he that feareth God shall come forth of them all.
ECCL|7|19|Wisdom strengtheneth the wise more than ten mighty men which are in the city.
ECCL|7|20|For there is not a just man upon earth, that doeth good, and sinneth not.
ECCL|7|21|Also take no heed unto all words that are spoken; lest thou hear thy servant curse thee:
ECCL|7|22|For oftentimes also thine own heart knoweth that thou thyself likewise hast cursed others.
ECCL|7|23|All this have I proved by wisdom: I said, I will be wise; but it was far from me.
ECCL|7|24|That which is far off, and exceeding deep, who can find it out?
ECCL|7|25|I applied mine heart to know, and to search, and to seek out wisdom, and the reason of things, and to know the wickedness of folly, even of foolishness and madness:
ECCL|7|26|And I find more bitter than death the woman, whose heart is snares and nets, and her hands as bands: whoso pleaseth God shall escape from her; but the sinner shall be taken by her.
ECCL|7|27|Behold, this have I found, saith the preacher, counting one by one, to find out the account:
ECCL|7|28|Which yet my soul seeketh, but I find not: one man among a thousand have I found; but a woman among all those have I not found.
ECCL|7|29|Lo, this only have I found, that God hath made man upright; but they have sought out many inventions.
ECCL|8|1|Who is as the wise man? and who knoweth the interpretation of a thing? a man's wisdom maketh his face to shine, and the boldness of his face shall be changed.
ECCL|8|2|I counsel thee to keep the king's commandment, and that in regard of the oath of God.
ECCL|8|3|Be not hasty to go out of his sight: stand not in an evil thing; for he doeth whatsoever pleaseth him.
ECCL|8|4|Where the word of a king is, there is power: and who may say unto him, What doest thou?
ECCL|8|5|Whoso keepeth the commandment shall feel no evil thing: and a wise man's heart discerneth both time and judgment.
ECCL|8|6|Because to every purpose there is time and judgment, therefore the misery of man is great upon him.
ECCL|8|7|For he knoweth not that which shall be: for who can tell him when it shall be?
ECCL|8|8|There is no man that hath power over the spirit to retain the spirit; neither hath he power in the day of death: and there is no discharge in that war; neither shall wickedness deliver those that are given to it.
ECCL|8|9|All this have I seen, and applied my heart unto every work that is done under the sun: there is a time wherein one man ruleth over another to his own hurt.
ECCL|8|10|And so I saw the wicked buried, who had come and gone from the place of the holy, and they were forgotten in the city where they had so done: this is also vanity.
ECCL|8|11|Because sentence against an evil work is not executed speedily, therefore the heart of the sons of men is fully set in them to do evil.
ECCL|8|12|Though a sinner do evil an hundred times, and his days be prolonged, yet surely I know that it shall be well with them that fear God, which fear before him:
ECCL|8|13|But it shall not be well with the wicked, neither shall he prolong his days, which are as a shadow; because he feareth not before God.
ECCL|8|14|There is a vanity which is done upon the earth; that there be just men, unto whom it happeneth according to the work of the wicked; again, there be wicked men, to whom it happeneth according to the work of the righteous: I said that this also is vanity.
ECCL|8|15|Then I commended mirth, because a man hath no better thing under the sun, than to eat, and to drink, and to be merry: for that shall abide with him of his labour the days of his life, which God giveth him under the sun.
ECCL|8|16|When I applied mine heart to know wisdom, and to see the business that is done upon the earth: (for also there is that neither day nor night seeth sleep with his eyes:)
ECCL|8|17|Then I beheld all the work of God, that a man cannot find out the work that is done under the sun: because though a man labour to seek it out, yet he shall not find it; yea farther; though a wise man think to know it, yet shall he not be able to find it.
ECCL|9|1|For all this I considered in my heart even to declare all this, that the righteous, and the wise, and their works, are in the hand of God: no man knoweth either love or hatred by all that is before them.
ECCL|9|2|All things come alike to all: there is one event to the righteous, and to the wicked; to the good and to the clean, and to the unclean; to him that sacrificeth, and to him that sacrificeth not: as is the good, so is the sinner; and he that sweareth, as he that feareth an oath.
ECCL|9|3|This is an evil among all things that are done under the sun, that there is one event unto all: yea, also the heart of the sons of men is full of evil, and madness is in their heart while they live, and after that they go to the dead.
ECCL|9|4|For to him that is joined to all the living there is hope: for a living dog is better than a dead lion.
ECCL|9|5|For the living know that they shall die: but the dead know not any thing, neither have they any more a reward; for the memory of them is forgotten.
ECCL|9|6|Also their love, and their hatred, and their envy, is now perished; neither have they any more a portion for ever in any thing that is done under the sun.
ECCL|9|7|Go thy way, eat thy bread with joy, and drink thy wine with a merry heart; for God now accepteth thy works.
ECCL|9|8|Let thy garments be always white; and let thy head lack no ointment.
ECCL|9|9|Live joyfully with the wife whom thou lovest all the days of the life of thy vanity, which he hath given thee under the sun, all the days of thy vanity: for that is thy portion in this life, and in thy labour which thou takest under the sun.
ECCL|9|10|Whatsoever thy hand findeth to do, do it with thy might; for there is no work, nor device, nor knowledge, nor wisdom, in the grave, whither thou goest.
ECCL|9|11|I returned, and saw under the sun, that the race is not to the swift, nor the battle to the strong, neither yet bread to the wise, nor yet riches to men of understanding, nor yet favour to men of skill; but time and chance happeneth to them all.
ECCL|9|12|For man also knoweth not his time: as the fishes that are taken in an evil net, and as the birds that are caught in the snare; so are the sons of men snared in an evil time, when it falleth suddenly upon them.
ECCL|9|13|This wisdom have I seen also under the sun, and it seemed great unto me:
ECCL|9|14|There was a little city, and few men within it; and there came a great king against it, and besieged it, and built great bulwarks against it:
ECCL|9|15|Now there was found in it a poor wise man, and he by his wisdom delivered the city; yet no man remembered that same poor man.
ECCL|9|16|Then said I, Wisdom is better than strength: nevertheless the poor man's wisdom is despised, and his words are not heard.
ECCL|9|17|The words of wise men are heard in quiet more than the cry of him that ruleth among fools.
ECCL|9|18|Wisdom is better than weapons of war: but one sinner destroyeth much good.
ECCL|10|1|Dead flies cause the ointment of the apothecary to send forth a stinking savour: so doth a little folly him that is in reputation for wisdom and honour.
ECCL|10|2|A wise man's heart is at his right hand; but a fool's heart at his left.
ECCL|10|3|Yea also, when he that is a fool walketh by the way, his wisdom faileth him, and he saith to every one that he is a fool.
ECCL|10|4|If the spirit of the ruler rise up against thee, leave not thy place; for yielding pacifieth great offences.
ECCL|10|5|There is an evil which I have seen under the sun, as an error which proceedeth from the ruler:
ECCL|10|6|Folly is set in great dignity, and the rich sit in low place.
ECCL|10|7|I have seen servants upon horses, and princes walking as servants upon the earth.
ECCL|10|8|He that diggeth a pit shall fall into it; and whoso breaketh an hedge, a serpent shall bite him.
ECCL|10|9|Whoso removeth stones shall be hurt therewith; and he that cleaveth wood shall be endangered thereby.
ECCL|10|10|If the iron be blunt, and he do not whet the edge, then must he put to more strength: but wisdom is profitable to direct.
ECCL|10|11|Surely the serpent will bite without enchantment; and a babbler is no better.
ECCL|10|12|The words of a wise man's mouth are gracious; but the lips of a fool will swallow up himself.
ECCL|10|13|The beginning of the words of his mouth is foolishness: and the end of his talk is mischievous madness.
ECCL|10|14|A fool also is full of words: a man cannot tell what shall be; and what shall be after him, who can tell him?
ECCL|10|15|The labour of the foolish wearieth every one of them, because he knoweth not how to go to the city.
ECCL|10|16|Woe to thee, O land, when thy king is a child, and thy princes eat in the morning!
ECCL|10|17|Blessed art thou, O land, when thy king is the son of nobles, and thy princes eat in due season, for strength, and not for drunkenness!
ECCL|10|18|By much slothfulness the building decayeth; and through idleness of the hands the house droppeth through.
ECCL|10|19|A feast is made for laughter, and wine maketh merry: but money answereth all things.
ECCL|10|20|Curse not the king, no not in thy thought; and curse not the rich in thy bedchamber: for a bird of the air shall carry the voice, and that which hath wings shall tell the matter.
ECCL|11|1|Cast thy bread upon the waters: for thou shalt find it after many days.
ECCL|11|2|Give a portion to seven, and also to eight; for thou knowest not what evil shall be upon the earth.
ECCL|11|3|If the clouds be full of rain, they empty themselves upon the earth: and if the tree fall toward the south, or toward the north, in the place where the tree falleth, there it shall be.
ECCL|11|4|He that observeth the wind shall not sow; and he that regardeth the clouds shall not reap.
ECCL|11|5|As thou knowest not what is the way of the spirit, nor how the bones do grow in the womb of her that is with child: even so thou knowest not the works of God who maketh all.
ECCL|11|6|In the morning sow thy seed, and in the evening withhold not thine hand: for thou knowest not whether shall prosper, either this or that, or whether they both shall be alike good.
ECCL|11|7|Truly the light is sweet, and a pleasant thing it is for the eyes to behold the sun:
ECCL|11|8|But if a man live many years, and rejoice in them all; yet let him remember the days of darkness; for they shall be many. All that cometh is vanity.
ECCL|11|9|Rejoice, O young man, in thy youth; and let thy heart cheer thee in the days of thy youth, and walk in the ways of thine heart, and in the sight of thine eyes: but know thou, that for all these things God will bring thee into judgment.
ECCL|11|10|Therefore remove sorrow from thy heart, and put away evil from thy flesh: for childhood and youth are vanity.
ECCL|12|1|Remember now thy Creator in the days of thy youth, while the evil days come not, nor the years draw nigh, when thou shalt say, I have no pleasure in them;
ECCL|12|2|While the sun, or the light, or the moon, or the stars, be not darkened, nor the clouds return after the rain:
ECCL|12|3|In the day when the keepers of the house shall tremble, and the strong men shall bow themselves, and the grinders cease because they are few, and those that look out of the windows be darkened,
ECCL|12|4|And the doors shall be shut in the streets, when the sound of the grinding is low, and he shall rise up at the voice of the bird, and all the daughters of musick shall be brought low;
ECCL|12|5|Also when they shall be afraid of that which is high, and fears shall be in the way, and the almond tree shall flourish, and the grasshopper shall be a burden, and desire shall fail: because man goeth to his long home, and the mourners go about the streets:
ECCL|12|6|Or ever the silver cord be loosed, or the golden bowl be broken, or the pitcher be broken at the fountain, or the wheel broken at the cistern.
ECCL|12|7|Then shall the dust return to the earth as it was: and the spirit shall return unto God who gave it.
ECCL|12|8|Vanity of vanities, saith the preacher; all is vanity.
ECCL|12|9|And moreover, because the preacher was wise, he still taught the people knowledge; yea, he gave good heed, and sought out, and set in order many proverbs.
ECCL|12|10|The preacher sought to find out acceptable words: and that which was written was upright, even words of truth.
ECCL|12|11|The words of the wise are as goads, and as nails fastened by the masters of assemblies, which are given from one shepherd.
ECCL|12|12|And further, by these, my son, be admonished: of making many books there is no end; and much study is a weariness of the flesh.
ECCL|12|13|Let us hear the conclusion of the whole matter: Fear God, and keep his commandments: for this is the whole duty of man.
ECCL|12|14|For God shall bring every work into judgment, with every secret thing, whether it be good, or whether it be evil.
