2KGS|1|1|praevaricatus est autem Moab in Israhel postquam mortuus est Ahab
2KGS|1|2|ceciditque Ohozias per cancellos cenaculi sui quod habebat in Samaria et aegrotavit misitque nuntios dicens ad eos ite consulite Beelzebub deum Accaron utrum vivere queam de infirmitate mea hac
2KGS|1|3|angelus autem Domini locutus est ad Heliam Thesbiten surge ascende in occursum nuntiorum regis Samariae et dices ad eos numquid non est Deus in Israhel ut eatis ad consulendum Beelzebub deum Accaron
2KGS|1|4|quam ob rem haec dicit Dominus de lectulo super quem ascendisti non descendes sed morte morieris et abiit Helias
2KGS|1|5|reversique sunt nuntii ad Ohoziam qui dixit eis quare reversi estis
2KGS|1|6|at illi responderunt ei vir occurrit nobis et dixit ad nos ite revertimini ad regem qui misit vos et dicetis ei haec dicit Dominus numquid quia non erat Deus in Israhel mittis ut consulatur Beelzebub deus Accaron idcirco de lectulo super quem ascendisti non descendes sed morte morieris
2KGS|1|7|qui dixit eis cuius figurae et habitu est vir qui occurrit vobis et locutus est verba haec
2KGS|1|8|at illi dixerunt vir pilosus et zona pellicia accinctis renibus qui ait Helias Thesbites est
2KGS|1|9|misitque ad eum quinquagenarium principem et quinquaginta qui erant sub eo qui ascendit ad eum sedentique in vertice montis ait homo Dei rex praecepit ut descendas
2KGS|1|10|respondensque Helias dixit quinquagenario si homo Dei sum descendat ignis e caelo et devoret te et quinquaginta tuos descendit itaque ignis e caelo et devoravit eum et quinquaginta qui erant cum eo
2KGS|1|11|rursum misit ad eum principem quinquagenarium alterum et quinquaginta cum eo qui locutus est illi homo Dei haec dicit rex festina descende
2KGS|1|12|respondens Helias ait si homo Dei ego sum descendat ignis e caelo et devoret te et quinquaginta tuos descendit ergo ignis Dei e caelo et devoravit illum et quinquaginta eius
2KGS|1|13|iterum misit principem quinquagenarium tertium et quinquaginta qui erant cum eo qui cum venisset curvavit genua contra Heliam et precatus est eum et ait homo Dei noli despicere animam meam et animam servorum tuorum qui mecum sunt
2KGS|1|14|ecce descendit ignis de caelo et devoravit duos principes quinquagenarios primos et quinquagenos qui cum eis erant sed nunc obsecro ut miserearis animae meae
2KGS|1|15|locutus est autem angelus Domini ad Heliam dicens descende cum eo ne timeas surrexit igitur et descendit cum eo ad regem
2KGS|1|16|et locutus est ei haec dicit Dominus quia misisti nuntios ad consulendum Beelzebub deum Accaron quasi non esset Deus in Israhel a quo possis interrogare sermonem ideo de lectulo super quem ascendisti non descendes sed morte morieris
2KGS|1|17|mortuus est ergo iuxta sermonem Domini quem locutus est Helias et regnavit Ioram frater eius pro eo anno secundo Ioram filii Iosaphat regis Iudae non enim habebat filium
2KGS|1|18|reliqua autem verborum Ohoziae quae operatus est nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|2|1|factum est autem cum levare vellet Dominus Heliam per turbinem in caelum ibant Helias et Heliseus de Galgalis
2KGS|2|2|dixitque Helias ad Heliseum sede hic quia Dominus misit me usque Bethel cui ait Heliseus vivit Dominus et vivit anima tua quia non derelinquam te cumque descendissent Bethel
2KGS|2|3|egressi sunt filii prophetarum qui erant Bethel ad Heliseum et dixerunt ei numquid nosti quia hodie Dominus tollat dominum tuum a te qui respondit et ego novi silete
2KGS|2|4|dixit autem Helias ad Heliseum sede hic quia Dominus misit me in Hiericho et ille ait vivit Dominus et vivit anima tua quia non derelinquam te cumque venissent Hierichum
2KGS|2|5|accesserunt filii prophetarum qui erant in Hiericho ad Heliseum et dixerunt ei numquid nosti quia hodie Dominus tollet dominum tuum a te et ait et ego novi silete
2KGS|2|6|dixit autem ei Helias sede hic quia Dominus misit me ad Iordanem qui ait vivit Dominus et vivit anima tua quia non derelinquam te ierunt igitur ambo pariter
2KGS|2|7|et quinquaginta viri de filiis prophetarum secuti sunt qui et steterunt e contra longe illi autem ambo stabant super Iordanem
2KGS|2|8|tulitque Helias pallium suum et involvit illud et percussit aquas quae divisae sunt in utramque partem et transierunt ambo per siccum
2KGS|2|9|cumque transissent Helias dixit ad Heliseum postula quod vis ut faciam tibi antequam tollar a te dixitque Heliseus obsecro ut fiat duplex spiritus tuus in me
2KGS|2|10|qui respondit rem difficilem postulasti attamen si videris me quando tollor a te erit quod petisti si autem non videris non erit
2KGS|2|11|cumque pergerent et incedentes sermocinarentur ecce currus igneus et equi ignei diviserunt utrumque et ascendit Helias per turbinem in caelum
2KGS|2|12|Heliseus autem videbat et clamabat pater mi pater mi currus Israhel et auriga eius et non vidit eum amplius adprehenditque vestimenta sua et scidit illa in duas partes
2KGS|2|13|et levavit pallium Heliae quod ceciderat ei reversusque stetit super ripam Iordanis
2KGS|2|14|et pallio Heliae quod ceciderat ei percussit aquas et dixit ubi est Deus Heliae etiam nunc percussitque aquas et divisae sunt huc atque illuc et transiit Heliseus
2KGS|2|15|videntes autem filii prophetarum qui erant in Hiericho de contra dixerunt requievit spiritus Heliae super Heliseum et venientes in occursum eius adoraverunt eum proni in terram
2KGS|2|16|dixeruntque illi ecce cum servis tuis sunt quinquaginta viri fortes qui possint ire et quaerere dominum tuum ne forte tulerit eum spiritus Domini et proiecerit in uno montium aut in una vallium qui ait nolite mittere
2KGS|2|17|coegeruntque eum donec adquiesceret et diceret mittite et miserunt quinquaginta viros qui cum quaesissent tribus diebus non invenerunt
2KGS|2|18|et reversi sunt ad eum at ille habitabat in Hiericho dixitque eis numquid non dixi vobis nolite ire
2KGS|2|19|dixerunt quoque viri civitatis ad Heliseum ecce habitatio civitatis huius optima est sicut tu ipse domine perspicis sed aquae pessimae sunt et terra sterilis
2KGS|2|20|at ille ait adferte mihi vas novum et mittite in illud sal qui cum adtulissent
2KGS|2|21|egressus ad fontem aquarum misit in eum sal et ait haec dicit Dominus sanavi aquas has et non erit ultra in eis mors neque sterilitas
2KGS|2|22|sanatae sunt ergo aquae usque ad diem hanc iuxta verbum Helisei quod locutus est
2KGS|2|23|ascendit autem inde Bethel cumque ascenderet per viam pueri parvi egressi sunt de civitate et inludebant ei dicentes ascende calve ascende calve
2KGS|2|24|qui cum se respexisset vidit eos et maledixit eis in nomine Domini egressique sunt duo ursi de saltu et laceraverunt ex eis quadraginta duos pueros
2KGS|2|25|abiit autem inde in montem Carmeli et inde reversus est Samariam
2KGS|3|1|Ioram vero filius Ahab regnavit super Israhel in Samaria anno octavodecimo Iosaphat regis Iudae regnavitque duodecim annis
2KGS|3|2|et fecit malum coram Domino sed non sicut pater suus et mater tulit enim statuas Baal quas fecerat pater eius
2KGS|3|3|verumtamen in peccatis Hieroboam filii Nabath qui peccare fecit Israhel adhesit nec recessit ab eis
2KGS|3|4|porro Mesa rex Moab nutriebat pecora multa et solvebat regi Israhel centum milia agnorum et centum milia arietum cum velleribus suis
2KGS|3|5|cumque mortuus fuisset Ahab praevaricatus est foedus quod habebat cum rege Israhel
2KGS|3|6|egressus est igitur rex Ioram in die illa de Samaria et recensuit universum Israhel
2KGS|3|7|misitque ad Iosaphat regem Iuda dicens rex Moab recessit a me veni mecum contra Moab ad proelium qui respondit ascendam qui meus est tuus est populus meus populus tuus equi mei equi tui
2KGS|3|8|dixitque per quam viam ascendemus at ille respondit per desertum Idumeae
2KGS|3|9|perrexerunt igitur rex Israhel et rex Iuda et rex Edom et circumierunt per viam septem dierum nec erat aqua exercitui et iumentis quae sequebantur eos
2KGS|3|10|dixitque rex Israhel eheu eheu eheu congregavit nos Dominus tres reges ut traderet in manu Moab
2KGS|3|11|et ait Iosaphat estne hic propheta Domini ut deprecemur Dominum per eum et respondit unus de servis regis Israhel est hic Heliseus filius Saphat qui fundebat aquam super manus Heliae
2KGS|3|12|et ait Iosaphat est apud eum sermo Domini descenditque ad eum rex Israhel et Iosaphat et rex Edom
2KGS|3|13|dixit autem Heliseus ad regem Israhel quid mihi et tibi est vade ad prophetas patris tui et matris tuae et ait illi rex Israhel quare congregavit Dominus tres reges hos ut traderet eos in manu Moab
2KGS|3|14|dixit autem Heliseus vivit Dominus exercituum in cuius conspectu sto quod si non vultum Iosaphat regis Iudae erubescerem ne adtendissem quidem te nec respexissem
2KGS|3|15|nunc autem adducite mihi psalten cumque caneret psaltes facta est super eum manus Domini et ait
2KGS|3|16|haec dicit Dominus facite alveum torrentis huius fossas et fossas
2KGS|3|17|haec enim dicit Dominus non videbitis ventum neque pluviam et alveus iste replebitur aquis et bibetis vos et familiae vestrae et iumenta vestra
2KGS|3|18|parumque hoc est in conspectu Domini insuper tradet etiam Moab in manu vestra
2KGS|3|19|et percutietis omnem civitatem munitam et omnem urbem electam et universum lignum fructiferum succidetis cunctosque fontes aquarum obturabitis et omnem agrum egregium operietis lapidibus
2KGS|3|20|factum est igitur mane quando sacrificium offerri solet et ecce aquae veniebant per viam Edom et repleta est terra aquis
2KGS|3|21|universi autem Moabitae audientes quod ascendissent reges ut pugnarent adversum eos convocaverunt omnes qui accincti erant balteo desuper et steterunt in terminis
2KGS|3|22|primoque mane surgentes et orto iam sole ex adverso aquarum viderunt Moabitae contra aquas rubras quasi sanguinem
2KGS|3|23|dixeruntque sanguis est gladii pugnaverunt reges contra se et caesi sunt mutuo nunc perge ad praedam Moab
2KGS|3|24|perrexeruntque in castra Israhel porro consurgens Israhel percussit Moab at illi fugerunt coram eis venerunt igitur qui vicerant et percusserunt Moab
2KGS|3|25|et civitates destruxerunt et omnem agrum optimum mittentes singuli lapides repleverunt et universos fontes aquarum obturaverunt et omnia ligna fructifera succiderunt ita ut muri tantum fictiles remanerent et circumdata est civitas a fundibalariis et magna ex parte percussa
2KGS|3|26|quod cum vidisset rex Moab praevaluisse scilicet hostes tulit secum septingentos viros educentes gladium ut inrumperet ad regem Edom et non potuerunt
2KGS|3|27|arripiensque filium suum primogenitum qui regnaturus erat pro eo obtulit holocaustum super murum et facta est indignatio magna in Israhel statimque recesserunt ab eo et reversi sunt in terram suam
2KGS|4|1|mulier autem quaedam de uxoribus prophetarum clamabat ad Heliseum dicens servus tuus vir meus mortuus est et tu nosti quia servus tuus fuit timens Dominum et ecce creditor venit ut tollat duos filios meos ad serviendum sibi
2KGS|4|2|cui dixit Heliseus quid vis ut faciam tibi dic mihi quid habes in domo tua at illa respondit non habeo ancilla tua quicquam in domo mea nisi parum olei quo unguear
2KGS|4|3|cui ait vade pete mutuo ab omnibus vicinis tuis vasa vacua non pauca
2KGS|4|4|et ingredere et claude ostium cum intrinsecus fueris tu et filii tui et mitte inde in omnia vasa haec et cum plena fuerint tolles
2KGS|4|5|ivit itaque mulier et clusit ostium super se et super filios suos illi offerebant vasa et illa infundebat
2KGS|4|6|cumque plena fuissent vasa dixit ad filium suum adfer mihi adhuc vas et ille respondit non habeo stetitque oleum
2KGS|4|7|venit autem illa et indicavit homini Dei et ille vade inquit vende oleum et redde creditori tuo tu autem et filii tui vivite de reliquo
2KGS|4|8|facta est autem quaedam dies et transiebat Heliseus per Sunam erat autem ibi mulier magna quae tenuit eum ut comederet panem cumque frequenter inde transiret devertebat ad eam ut comederet panem
2KGS|4|9|quae dixit ad virum suum animadverto quod vir Dei sanctus est iste qui transit per nos frequenter
2KGS|4|10|faciamus ergo cenaculum parvum et ponamus ei in eo lectulum et mensam et sellam et candelabrum ut cum venerit ad nos maneat ibi
2KGS|4|11|facta est igitur dies quaedam et veniens devertit in cenaculum et requievit ibi
2KGS|4|12|dixitque ad Giezi puerum suum voca Sunamitin istam qui cum vocasset eam et illa stetisset coram eo
2KGS|4|13|dixit ad puerum loquere ad eam ecce sedule in omnibus ministrasti nobis quid vis ut faciam tibi numquid habes negotium et vis ut loquar regi sive principi militiae quae respondit in medio populi mei habito
2KGS|4|14|et ait quid ergo vult ut faciam ei dixitque Giezi ne quaeras filium enim non habet et vir eius senex est
2KGS|4|15|praecepit itaque ut vocaret eam quae cum vocata fuisset et stetisset ad ostium
2KGS|4|16|dixit ad eam in tempore isto et in hac eadem hora si vita comes fuerit habebis in utero filium at illa respondit noli quaeso domine mi vir Dei noli mentiri ancillae tuae
2KGS|4|17|et concepit mulier et peperit filium in tempore et in hora eadem quam dixerat Heliseus
2KGS|4|18|crevit autem puer et cum esset quaedam dies et egressus isset ad patrem suum ad messores
2KGS|4|19|ait patri suo caput meum caput meum at ille dixit puero tolle et duc eum ad matrem suam
2KGS|4|20|qui cum tulisset et adduxisset eum ad matrem suam posuit eum illa super genua sua usque ad meridiem et mortuus est
2KGS|4|21|ascendit autem et conlocavit eum super lectulum hominis Dei et clusit ostium et egressa
2KGS|4|22|vocavit virum suum et ait mitte mecum obsecro unum de pueris et asinam ut excurram usque ad hominem Dei et revertar
2KGS|4|23|qui ait illi quam ob causam vadis ad eum hodie non sunt kalendae neque sabbatum quae respondit vale
2KGS|4|24|stravitque asinam et praecepit puero mina et propera ne mihi moram facias in eundo et hoc age quod praecipio tibi
2KGS|4|25|profecta est igitur et venit ad virum Dei in montem Carmeli cumque vidisset eam vir Dei de contra ait ad Giezi puerum suum ecce Sunamitis illa
2KGS|4|26|vade ergo in occursum eius et dic ei rectene agitur circa te et circa virum tuum et circa filium tuum quae respondit recte
2KGS|4|27|cumque venisset ad virum Dei in monte adprehendit pedes eius et accessit Giezi ut amoveret eam et ait homo Dei dimitte illam anima enim eius in amaritudine est et Dominus celavit me et non indicavit mihi
2KGS|4|28|quae dixit illi numquid petivi filium a domino meo numquid non dixi tibi ne inludas me
2KGS|4|29|et ille ait ad Giezi accinge lumbos tuos et tolle baculum meum in manu tua et vade si occurrerit tibi homo non salutes eum et si salutaverit te quispiam non respondeas illi et pones baculum meum super faciem pueri
2KGS|4|30|porro mater pueri ait vivit Dominus et vivit anima tua non dimittam te surrexit ergo et secutus est eam
2KGS|4|31|Giezi autem praecesserat eos et posuerat baculum super faciem pueri et non erat vox neque sensus reversusque est in occursum eius et nuntiavit ei dicens non surrexit puer
2KGS|4|32|ingressus est ergo Heliseus domum et ecce puer mortuus iacebat in lectulo eius
2KGS|4|33|ingressusque clusit ostium super se et puerum et oravit ad Dominum
2KGS|4|34|et ascendit et incubuit super puerum posuitque os suum super os eius et oculos suos super oculos eius et manus suas super manus eius et incurvavit se super eum et calefacta est caro pueri
2KGS|4|35|at ille reversus deambulavit in domo semel huc et illuc et ascendit et incubuit super eum et oscitavit puer septies aperuitque oculos
2KGS|4|36|et ille vocavit Giezi et dixit ei voca Sunamitin hanc quae vocata ingressa est ad eum qui ait tolle filium tuum
2KGS|4|37|venit illa et corruit ad pedes eius et adoravit super terram tulitque filium suum et egressa est
2KGS|4|38|et Heliseus reversus est in Galgala erat autem fames in terra et filii prophetarum habitabant coram eo dixitque uni de pueris suis pone ollam grandem et coque pulmentum filiis prophetarum
2KGS|4|39|et egressus est unus in agrum ut colligeret herbas agrestes invenitque quasi vitem silvestrem et collegit ex ea colocyntidas agri et implevit pallium suum et reversus concidit in ollam pulmenti nesciebat enim quid esset
2KGS|4|40|infuderunt ergo sociis ut comederent cumque gustassent de coctione exclamaverunt dicentes mors in olla vir Dei et non potuerunt comedere
2KGS|4|41|at ille adferte inquit farinam et misit in ollam et ait infunde turbae et comedat et non fuit amplius quicquam amaritudinis in olla
2KGS|4|42|vir autem quidam venit de Balsalisa deferens viro Dei panes primitiarum et viginti panes hordiacios et frumentum novum in pera sua at ille dixit da populo ut comedat
2KGS|4|43|responditque ei minister eius quantum est hoc ut adponam coram centum viris rursum ille da ait populo ut comedat haec enim dicit Dominus comedent et supererit
2KGS|4|44|posuit itaque coram eis qui comederunt et superfuit iuxta verbum Domini
2KGS|5|1|Naaman princeps militiae regis Syriae erat vir magnus apud dominum suum et honoratus per illum enim dedit Dominus salutem Syriae erat autem vir fortis et dives sed leprosus
2KGS|5|2|porro de Syria egressi fuerant latrunculi et captivam duxerant de terra Israhel puellam parvulam quae erat in obsequio uxoris Naaman
2KGS|5|3|quae ait ad dominam suam utinam fuisset dominus meus ad prophetam qui est in Samaria profecto curasset eum a lepra quam habet
2KGS|5|4|ingressus est itaque Naaman ad dominum suum et nuntiavit ei dicens sic et sic locuta est puella de terra Israhel
2KGS|5|5|dixitque ei rex Syriae vade et mittam litteras ad regem Israhel qui cum profectus esset et tulisset secum decem talenta argenti et sex milia aureos et decem mutatoria vestimentorum
2KGS|5|6|detulit litteras ad regem Israhel in haec verba cum acceperis epistulam hanc scito quod miserim ad te Naaman servum meum ut cures eum a lepra sua
2KGS|5|7|cumque legisset rex Israhel litteras scidit vestimenta sua et ait numquid Deus sum ut occidere possim et vivificare quia iste misit ad me ut curem hominem a lepra sua animadvertite et videte quod occasiones quaerat adversum me
2KGS|5|8|quod cum audisset Heliseus vir Dei scidisse videlicet regem Israhel vestimenta sua misit ad eum dicens quare scidisti vestimenta tua veniat ad me et sciat esse prophetam in Israhel
2KGS|5|9|venit ergo Naaman cum equis et curribus et stetit ad ostium domus Helisei
2KGS|5|10|misitque ad eum Heliseus nuntium dicens vade et lavare septies in Iordane et recipiet sanitatem caro tua atque mundaberis
2KGS|5|11|iratus Naaman recedebat dicens putabam quod egrederetur ad me et stans invocaret nomen Domini Dei sui et tangeret manu sua locum leprae et curaret me
2KGS|5|12|numquid non meliores sunt Abana et Pharphar fluvii Damasci omnibus aquis Israhel ut laver in eis et munder cum ergo vertisset se et abiret indignans
2KGS|5|13|accesserunt ad eum servi sui et locuti sunt ei pater si rem grandem dixisset tibi propheta certe facere debueras quanto magis quia nunc dixit tibi lavare et mundaberis
2KGS|5|14|descendit et lavit in Iordane septies iuxta sermonem viri Dei et restituta est caro eius sicut caro pueri parvuli et mundatus est
2KGS|5|15|reversusque ad virum Dei cum universo comitatu suo venit et stetit coram eo et ait vere scio quod non sit Deus in universa terra nisi tantum in Israhel obsecro itaque ut accipias benedictionem a servo tuo
2KGS|5|16|at ille respondit vivit Dominus ante quem sto quia non accipiam cumque vim faceret penitus non adquievit
2KGS|5|17|dixitque Naaman ut vis sed obsecro concede mihi servo tuo ut tollam onus duorum burdonum de terra non enim faciet ultra servus tuus holocaustum aut victimam diis alienis nisi Domino
2KGS|5|18|hoc autem solum est de quo depreceris Dominum pro servo tuo quando ingreditur dominus meus templum Remmon ut adoret et illo innitente super manum meam si adoravero in templo Remmon adorante me in eodem loco ut ignoscat mihi Dominus servo tuo pro hac re
2KGS|5|19|qui dixit ei vade in pace abiit ergo ab eo electo terrae tempore
2KGS|5|20|dixitque Giezi puer viri Dei pepercit dominus meus Naaman Syro isti ut non acciperet ab eo quae adtulit vivit Dominus quia curram post eum et accipiam ab eo aliquid
2KGS|5|21|et secutus est Giezi post tergum Naaman quem cum vidisset ille currentem ad se desilivit de curru in occursum eius et ait rectene sunt omnia
2KGS|5|22|et ille ait recte dominus meus misit me dicens modo venerunt ad me duo adulescentes de monte Ephraim ex filiis prophetarum da eis talentum argenti et vestes mutatorias duplices
2KGS|5|23|dixitque Naaman melius est ut accipias duo talenta et coegit eum ligavitque duo talenta argenti in duobus saccis et duplicia vestimenta et inposuit duobus pueris suis qui et portaverunt coram eo
2KGS|5|24|cumque venisset iam vesperi tulit de manu eorum et reposuit in domo dimisitque viros et abierunt
2KGS|5|25|ipse autem ingressus stetit coram domino suo et dixit Heliseus unde venis Giezi qui respondit non ivit servus tuus quoquam
2KGS|5|26|at ille nonne ait cor meum in praesenti erat quando reversus est homo de curru suo in occursum tui nunc igitur accepisti argentum et accepisti vestes ut emas oliveta et vineta et oves et boves et servos et ancillas
2KGS|5|27|sed et lepra Naaman adherebit tibi et semini tuo in sempiternum et egressus est ab eo leprosus quasi nix
2KGS|6|1|dixerunt autem filii prophetarum ad Heliseum ecce locus in quo habitamus coram te angustus est nobis
2KGS|6|2|eamus usque ad Iordanem et tollant singuli de silva materias singulas ut aedificemus nobis ibi locum ad habitandum qui dixit ite
2KGS|6|3|et ait unus ex illis veni ergo et tu cum servis tuis respondit ego veniam
2KGS|6|4|et abiit cum eis cumque venissent ad Iordanem caedebant ligna
2KGS|6|5|accidit autem ut cum unus materiem succidisset caderet ferrum securis in aquam exclamavitque ille et ait eheu eheu eheu domine mi et hoc ipsum mutuo acceperam
2KGS|6|6|dixit autem homo Dei ubi cecidit at ille monstravit ei locum praecidit ergo lignum et misit illuc natavitque ferrum
2KGS|6|7|et ait tolle qui extendit manum et tulit illud
2KGS|6|8|rex autem Syriae pugnabat contra Israhel consiliumque iniit cum servis suis dicens in loco illo et illo ponamus insidias
2KGS|6|9|misit itaque vir Dei ad regem Israhel dicens cave ne transeas in loco illo quia ibi Syri in insidiis sunt
2KGS|6|10|misit rex Israhel ad locum quem dixerat ei vir Dei et praeoccupavit eum et observavit se ibi non semel neque bis
2KGS|6|11|conturbatumque est cor regis Syriae pro hac re et convocatis servis suis ait quare non indicastis mihi quis proditor mei sit apud regem Israhel
2KGS|6|12|dixitque unus servorum eius nequaquam domine mi rex sed Heliseus propheta qui est in Israhel indicat regi Israhel omnia verba quaecumque locutus fueris in conclavi tuo
2KGS|6|13|dixit eis ite et videte ubi sit ut mittam et capiam eum adnuntiaveruntque ei dicentes ecce in Dothan
2KGS|6|14|misit ergo illuc equos et currus et robur exercitus qui cum venissent nocte circumdederunt civitatem
2KGS|6|15|consurgens autem diluculo minister viri Dei egressus est viditque exercitum in circuitu civitatis et equos et currus nuntiavitque ei dicens eheu eheu domine mi quid faciemus
2KGS|6|16|at ille respondit noli timere plures enim nobiscum sunt quam cum illis
2KGS|6|17|cumque orasset Heliseus ait Domine aperi oculos huius ut videat et aperuit Dominus oculos pueri et vidit et ecce mons plenus equorum et curruum igneorum in circuitu Helisei
2KGS|6|18|hostes vero descenderunt ad eum porro Heliseus oravit Dominum dicens percute obsecro gentem hanc caecitate percussitque eos Dominus ne viderent iuxta verbum Helisei
2KGS|6|19|dixit autem ad eos Heliseus non est haec via nec ista est civitas sequimini me et ostendam vobis virum quem quaeritis duxit ergo eos in Samariam
2KGS|6|20|cumque ingressi fuissent in Samaria dixit Heliseus Domine aperi oculos istorum ut videant aperuitque Dominus oculos eorum et viderunt esse se in medio Samariae
2KGS|6|21|dixitque rex Israhel ad Heliseum cum vidisset eos numquid percutiam eos pater mi
2KGS|6|22|at ille ait non percuties neque enim cepisti eos gladio et arcu tuo ut percutias pone panem et aquam coram eis ut comedant et bibant et vadant ad dominum suum
2KGS|6|23|adpositaque est eis ciborum magna praeparatio et comederunt et biberunt et dimisit eos abieruntque ad dominum suum et ultra non venerunt latrones Syriae in terram Israhel
2KGS|6|24|factum est autem post haec congregavit Benadad rex Syriae universum exercitum suum et ascendit et obsidebat Samariam
2KGS|6|25|factaque est fames magna in Samaria et tamdiu obsessa est donec venundaretur caput asini octoginta argenteis et quarta pars cabi stercoris columbarum quinque argenteis
2KGS|6|26|cumque rex Israhel transiret per murum mulier exclamavit ad eum dicens salva me domine mi rex
2KGS|6|27|qui ait non te salvet Dominus unde salvare te possum de area an de torculari dixitque ad eam rex quid tibi vis quae respondit
2KGS|6|28|mulier ista dixit mihi da filium tuum ut comedamus eum hodie et filium meum comedemus cras
2KGS|6|29|coximus ergo filium meum et comedimus dixique ei die altera da filium tuum ut comedamus eum quae abscondit filium suum
2KGS|6|30|quod cum audisset rex scidit vestimenta sua et transiebat super murum viditque omnis populus cilicium quo vestitus erat ad carnem intrinsecus
2KGS|6|31|et ait haec mihi faciat Deus et haec addat si steterit caput Helisei filii Saphat super eum hodie
2KGS|6|32|Heliseus autem sedebat in domo sua et senes sedebant cum eo praemisit itaque virum et antequam veniret nuntius ille dixit ad senes numquid scitis quod miserit filius homicidae hic ut praecidatur caput meum videte ergo cum venerit nuntius cludite ostium et non sinatis eum introire ecce enim sonitus pedum domini eius post eum est
2KGS|6|33|et adhuc illo loquente eis apparuit nuntius qui veniebat ad eum et ait ecce tantum malum a Domino est quid amplius expectabo a Domino
2KGS|7|1|dixit autem Heliseus audite verbum Domini haec dicit Dominus in tempore hoc cras modius similae uno statere erit et duo modii hordei statere uno in porta Samariae
2KGS|7|2|respondens unus de ducibus super cuius manum rex incumbebat homini Dei ait si Dominus fecerit etiam cataractas in caelo numquid poterit esse quod loqueris qui ait videbis oculis tuis et inde non comedes
2KGS|7|3|quattuor ergo viri erant leprosi iuxta introitum portae qui dixerunt ad invicem quid hic esse volumus donec moriamur
2KGS|7|4|sive ingredi voluerimus civitatem fame moriemur sive manserimus hic moriendum nobis est venite igitur et transfugiamus ad castra Syriae si pepercerint nobis vivemus si autem occidere voluerint nihilominus moriemur
2KGS|7|5|surrexerunt igitur vesperi ut venirent ad castra Syriae cumque venissent ad principium castrorum Syriae nullum ibidem reppererunt
2KGS|7|6|siquidem Dominus sonitum audiri fecerat in castris Syriae curruum et equorum et exercitus plurimi dixeruntque ad invicem ecce mercede conduxit adversum nos rex Israhel reges Hettheorum et Aegyptiorum et venerunt super nos
2KGS|7|7|surrexerunt ergo et fugerunt in tenebris et dereliquerunt tentoria sua et equos et asinos in castris fugeruntque animas tantum suas salvare cupientes
2KGS|7|8|igitur cum venissent leprosi illi ad principium castrorum ingressi sunt unum tabernaculum et comederunt et biberunt tuleruntque inde argentum et aurum et vestes et abierunt et absconderunt et rursum reversi sunt ad aliud tabernaculum et inde similiter auferentes absconderunt
2KGS|7|9|dixeruntque ad invicem non recte facimus haec enim dies boni nuntii est si tacuerimus et noluerimus nuntiare usque mane sceleris arguemur venite eamus et nuntiemus in aula regis
2KGS|7|10|cumque venissent ad portam civitatis narraverunt eis dicentes ivimus ad castra Syriae et nullum ibidem repperimus hominum nisi equos et asinos alligatos et fixa tentoria
2KGS|7|11|ierunt ergo portarii et nuntiaverunt in palatio regis intrinsecus
2KGS|7|12|qui surrexit nocte et ait ad servos suos dico vobis quid fecerint nobis Syri sciunt quia fame laboramus et idcirco egressi sunt de castris et latitant in agris dicentes cum egressi fuerint de civitate capiemus eos viventes et tunc civitatem ingredi poterimus
2KGS|7|13|respondit autem unus servorum eius tollamus quinque equos qui remanserunt in urbe quia ipsi tantum sunt in universa multitudine Israhel alii enim consumpti sunt et mittentes explorare poterimus
2KGS|7|14|adduxerunt ergo duos equos misitque rex ad castra Syrorum dicens ite videte
2KGS|7|15|qui abierunt post eos usque ad Iordanem ecce autem omnis via plena erat vestibus et vasis quae proiecerant Syri cum turbarentur reversique nuntii indicaverunt regi
2KGS|7|16|et egressus populus diripuit castra Syriae factusque est modius similae statere uno et duo modii hordei statere uno iuxta verbum Domini
2KGS|7|17|porro rex ducem illum in cuius manu incubuerat constituit ad portam quem conculcavit turba in introitu et mortuus est iuxta quod locutus fuerat vir Dei quando descenderat rex ad eum
2KGS|7|18|factumque est secundum sermonem viri Dei quem dixerat regi quando ait duo modii hordei statere uno erunt et modius similae statere uno hoc eodem tempore cras in porta Samariae
2KGS|7|19|quando responderat dux ille viro Dei et dixerat etiam si Dominus fecerit cataractas in caelo numquid fieri poterit quod loqueris et dixit ei videbis oculis tuis et inde non comedes
2KGS|7|20|evenit ergo ei sicut praedictum erat et conculcavit eum populus in porta et mortuus est
2KGS|8|1|Heliseus autem locutus est ad mulierem cuius vivere fecerat filium dicens surge vade tu et domus tua et peregrinare ubicumque reppereris vocavit enim Dominus famem et veniet super terram septem annis
2KGS|8|2|quae surrexit et fecit iuxta verbum hominis Dei et vadens cum domo sua peregrinata est in terra Philisthim diebus multis
2KGS|8|3|cumque finiti essent anni septem reversa est mulier de terra Philisthim et egressa est ut interpellaret regem pro domo sua et agris suis
2KGS|8|4|rex autem loquebatur cum Giezi puero viri Dei dicens narra mihi omnia magnalia quae fecit Heliseus
2KGS|8|5|cumque ille narraret regi quomodo mortuum suscitasset apparuit mulier cuius vivificaverat filium clamans ad regem pro domo sua et pro agris suis dixitque Giezi domine mi rex haec est mulier et hic filius eius quem suscitavit Heliseus
2KGS|8|6|et interrogavit rex mulierem quae narravit ei deditque ei rex eunuchum unum dicens restitue ei omnia quae sua sunt et universos reditus agrorum a die qua reliquit terram usque ad praesens
2KGS|8|7|venit quoque Heliseus Damascum et Benadad rex Syriae aegrotabat nuntiaveruntque ei dicentes venit vir Dei huc
2KGS|8|8|et ait rex ad Azahel tolle tecum munera et vade in occursum viri Dei et consule Dominum per eum dicens si evadere potero de infirmitate mea hac
2KGS|8|9|ivit igitur Azahel in occursum eius habens secum munera et omnia bona Damasci onera quadraginta camelorum cumque stetisset coram eo ait filius tuus Benadad rex Syriae misit me ad te dicens si sanari potero de infirmitate mea hac
2KGS|8|10|dixitque ei Heliseus vade dic ei sanaberis porro ostendit mihi Dominus quia morte morietur
2KGS|8|11|stetitque cum eo et conturbatus est usque ad suffusionem vultus flevitque vir Dei
2KGS|8|12|cui Azahel ait quare dominus meus flet at ille respondit quia scio quae facturus sis filiis Israhel mala civitates eorum munitas igne succendes et iuvenes eorum interficies gladio et parvulos eorum elides et praegnantes divides
2KGS|8|13|dixitque Azahel quid enim sum servus tuus canis ut faciam rem istam magnam et ait Heliseus ostendit mihi Dominus te regem Syriae fore
2KGS|8|14|qui cum recessisset ab Heliseo venit ad dominum suum qui ait ei quid tibi dixit Heliseus at ille respondit dixit mihi recipiet sanitatem
2KGS|8|15|cumque venisset dies altera tulit sagulum et infudit aqua et expandit super faciem eius quo mortuo regnavit Azahel pro eo
2KGS|8|16|anno quinto Ioram filii Ahab regis Israhel et Iosaphat regis Iuda regnavit Ioram filius Iosaphat rex Iuda
2KGS|8|17|triginta duorum erat annorum cum regnare coepisset et octo annis regnavit in Hierusalem
2KGS|8|18|ambulavitque in viis regum Israhel sicut ambulaverat domus Ahab filia enim Ahab erat uxor eius et fecit quod malum est coram Domino
2KGS|8|19|noluit autem Dominus disperdere Iudam propter David servum suum sicut promiserat ei ut daret illi lucernam et filiis eius cunctis diebus
2KGS|8|20|in diebus eius recessit Edom ne esset sub Iuda et constituit sibi regem
2KGS|8|21|venitque Ioram Seira et omnis currus cum eo et surrexit nocte percussitque Idumeos qui eum circumdederant et principes curruum populus autem fugit in tabernacula sua
2KGS|8|22|recessit ergo Edom ne esset sub Iuda usque ad diem hanc tunc recessit et Lobna in tempore illo
2KGS|8|23|reliqua autem sermonum Ioram et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|8|24|et dormivit Ioram cum patribus suis sepultusque est cum eis in civitate David et regnavit Ahazias filius eius pro eo
2KGS|8|25|anno duodecimo Ioram filii Ahab regis Israhel regnavit Ahazias filius Ioram regis Iudae
2KGS|8|26|viginti duorum annorum erat Ahazias cum regnare coepisset et uno anno regnavit in Hierusalem nomen matris eius Athalia filia Amri regis Israhel
2KGS|8|27|et ambulavit in viis domus Ahab et fecit quod malum est coram Domino sicut domus Ahab gener enim domus Ahab fuit
2KGS|8|28|abiit quoque cum Ioram filio Ahab ad proeliandum contra Azahel regem Syriae in Ramoth Galaad et vulneraverunt Syri Ioram
2KGS|8|29|qui reversus est ut curaretur in Hiezrahel quia vulneraverant eum Syri in Rama proeliantem contra Azahel regem Syriae porro Ahazias filius Ioram rex Iuda descendit invisere Ioram filium Ahab in Hiezrahel quia aegrotabat
2KGS|9|1|Heliseus autem prophetes vocavit unum de filiis prophetarum et ait illi accinge lumbos tuos et tolle lenticulam olei hanc in manu tua et vade in Ramoth Galaad
2KGS|9|2|cumque veneris illuc videbis Hieu filium Iosaphat filii Namsi et ingressus suscitabis eum de medio fratrum suorum et introduces interius cubiculum
2KGS|9|3|tenensque lenticulam olei fundes super caput eius et dices haec dicit Dominus unxi te regem super Israhel aperiesque ostium et fugies et non ibi subsistes
2KGS|9|4|abiit ergo adulescens puer prophetae Ramoth Galaad
2KGS|9|5|et ingressus est ecce autem principes exercitus sedebant et ait verbum mihi ad te princeps dixitque Hieu ad quem ex omnibus nobis at ille dixit ad te o princeps
2KGS|9|6|et surrexit et ingressus est cubiculum at ille fudit oleum super caput eius et ait haec dicit Dominus Deus Israhel unxi te regem super populum Domini Israhel
2KGS|9|7|et percuties domum Ahab domini tui ut ulciscar sanguinem servorum meorum prophetarum et sanguinem omnium servorum Domini de manu Hiezabel
2KGS|9|8|perdamque omnem domum Ahab et interficiam de Ahab mingentem ad parietem et clausum et novissimum in Israhel
2KGS|9|9|et dabo domum Ahab sicut domum Hieroboam filii Nabath et sicut domum Baasa filii Ahia
2KGS|9|10|Hiezabel quoque comedent canes in agro Hiezrahel nec erit qui sepeliat eam aperuitque ostium et fugit
2KGS|9|11|Hieu autem egressus est ad servos domini sui qui dixerunt ei rectene sunt omnia quid venit insanus iste ad te qui ait eis nostis hominem et quid locutus sit
2KGS|9|12|at illi responderunt falsum est sed magis narra nobis qui ait eis haec et haec locutus est mihi et ait haec dicit Dominus unxi te regem super Israhel
2KGS|9|13|festinaverunt itaque et unusquisque tollens pallium suum posuerunt sub pedibus eius in similitudinem tribunalis et cecinerunt tuba atque dixerunt regnavit Hieu
2KGS|9|14|coniuravit ergo Hieu filius Iosaphat filii Namsi contra Ioram porro Ioram obsederat Ramoth Galaad ipse et omnis Israhel contra Azahel regem Syriae
2KGS|9|15|et reversus fuerat ut curaretur in Hiezrahel propter vulnera quia percusserant eum Syri proeliantem contra Azahel regem Syriae dixitque Hieu si placet vobis nemo egrediatur profugus de civitate ne vadat et nuntiet in Hiezrahel
2KGS|9|16|et ascendit et profectus est in Hiezrahel Ioram enim aegrotabat ibi et Ahazia rex Iuda descenderat ad visitandum Ioram
2KGS|9|17|igitur speculator qui stabat super turrem Hiezrahel vidit globum Hieu venientis et ait video ego globum dixitque Ioram tolle currum et mitte in occursum eorum et dicat vadens rectene sunt omnia
2KGS|9|18|abiit igitur qui ascenderat currum in occursum eius et ait haec dicit rex pacata sunt omnia dixitque ei Hieu quid tibi et paci transi et sequere me nuntiavit quoque speculator dicens venit nuntius ad eos et non revertitur
2KGS|9|19|misit etiam currum equorum secundum venitque ad eos et ait haec dicit rex num pax est et ait Hieu quid tibi et paci transi et sequere me
2KGS|9|20|nuntiavit autem speculator dicens venit usque ad eos et non revertitur est autem incessus quasi incessus Hieu filii Namsi praeceps enim graditur
2KGS|9|21|et ait Ioram iunge currum iunxeruntque currum eius et egressus est Ioram rex Israhel et Ahazias rex Iuda singuli in curribus suis egressique sunt in occursum Hieu et invenerunt eum in agro Naboth Hiezrahelitis
2KGS|9|22|cumque vidisset Ioram Hieu dixit pax est Hieu at ille respondit quae pax adhuc fornicationes Hiezabel matris tuae et veneficia eius multa vigent
2KGS|9|23|convertit autem Ioram manum suam et fugiens ait ad Ahaziam insidiae Ahazia
2KGS|9|24|porro Hieu tetendit arcum manu et percussit Ioram inter scapulas et egressa est sagitta per cor eius statimque corruit in curru suo
2KGS|9|25|dixitque Hieu ad Baddacer ducem tolle proice eum in agro Naboth Hiezrahelitae memini enim quando ego et tu sedentes in curru sequebamur Ahab patrem huius quod Dominus onus hoc levaverit super eum dicens
2KGS|9|26|si non pro sanguine Naboth et pro sanguine filiorum eius quem vidi heri ait Dominus reddam tibi in agro isto dicit Dominus nunc igitur tolle proice eum in agro iuxta verbum Domini
2KGS|9|27|Ahazias autem rex Iuda videns hoc fugit per viam domus horti persecutusque est eum Hieu et ait etiam hunc percutite in curru suo in ascensu Gaber qui est iuxta Ieblaam qui fugit in Mageddo et mortuus est ibi
2KGS|9|28|et inposuerunt eum servi eius super currum suum et tulerunt Hierusalem sepelieruntque in sepulchro cum patribus suis in civitate David
2KGS|9|29|anno undecimo Ioram filii Ahab rege Ahazia super Iudam
2KGS|9|30|venit Hieu Hiezrahel porro Hiezabel introitu eius audito depinxit oculos suos stibio et ornavit caput suum et respexit per fenestram
2KGS|9|31|ingredientem Hieu per portam et ait numquid pax esse potest Zamri qui interfecit dominum suum
2KGS|9|32|levavitque Hieu faciem suam ad fenestram et ait quae est ista et inclinaverunt se ad eum duo vel tres eunuchi
2KGS|9|33|at ille dixit eis praecipitate eam deorsum et praecipitaverunt eam aspersusque est sanguine paries et equorum ungulae qui conculcaverunt eam
2KGS|9|34|cumque ingressus esset et comederet bibissetque ait ite videte maledictam illam et sepelite eam quia filia regis est
2KGS|9|35|cumque issent ut sepelirent eam non invenerunt nisi calvariam et pedes et summas manus
2KGS|9|36|reversique nuntiaverunt ei et ait Hieu sermo Domini est quem locutus est per servum suum Heliam Thesbiten dicens in agro Hiezrahel comedent canes carnes Hiezabel
2KGS|9|37|et erunt carnes Hiezabel sicut stercus super faciem terrae in agro Hiezrahel ita ut praetereuntes dicant haecine est illa Hiezabel
2KGS|10|1|erant autem Ahab septuaginta filii in Samaria scripsit ergo Hieu litteras et misit in Samariam ad optimates civitatis et ad maiores natu et ad nutricios Ahab dicens
2KGS|10|2|statim ut acceperitis litteras has qui habetis filios domini vestri et currus et equos et civitates firmas et arma
2KGS|10|3|eligite meliorem et eum qui vobis placuerit de filiis domini vestri et ponite eum super solium patris sui et pugnate pro domo domini vestri
2KGS|10|4|timuerunt illi vehementer et dixerunt ecce duo reges non potuerunt stare coram eo et quomodo nos valebimus resistere
2KGS|10|5|miserunt ergo praepositus domus et praefectus civitatis et maiores natu et nutricii ad Hieu dicentes servi tui sumus quaecumque iusseris faciemus nec constituemus regem quodcumque tibi placet fac
2KGS|10|6|rescripsit autem eis litteras secundo dicens si mei estis et oboeditis mihi tollite capita filiorum domini vestri et venite ad me hac eadem hora cras in Hiezrahel porro filii regis septuaginta viri apud optimates civitatis nutriebantur
2KGS|10|7|cumque venissent litterae ad eos tulerunt filios regis et occiderunt septuaginta viros et posuerunt capita eorum in cofinis et miserunt ad eum in Hiezrahel
2KGS|10|8|venit autem nuntius et indicavit ei dicens adtulerunt capita filiorum regis qui respondit ponite ea duos acervos iuxta introitum portae usque mane
2KGS|10|9|cumque diluxisset egressus est et stans dixit ad omnem populum iusti estis si ego coniuravi contra dominum meum et interfeci eum quis percussit omnes hos
2KGS|10|10|videte ergo nunc quoniam non cecidit de sermonibus Domini in terram quos locutus est Dominus super domum Ahab et Dominus fecit quod locutus est in manu servi sui Heliae
2KGS|10|11|percussit igitur Hieu omnes qui reliqui erant de domo Ahab in Hiezrahel et universos optimates eius et notos et sacerdotes donec non remanerent ex eo reliquiae
2KGS|10|12|et surrexit et venit in Samariam cumque venisset ad Camaram pastorum in via
2KGS|10|13|invenit fratres Ahaziae regis Iuda dixitque ad eos quinam estis vos at illi responderunt fratres Ahaziae sumus et descendimus ad salutandos filios regis et filios reginae
2KGS|10|14|qui ait conprehendite eos vivos quos cum conprehendissent vivos iugulaverunt eos in cisterna iuxta Camaram quadraginta duos viros et non reliquit ex eis quemquam
2KGS|10|15|cumque abisset inde invenit Ionadab filium Rechab in occursum sibi et benedixit ei et ait ad eum numquid est cor tuum rectum sicut cor meum cum corde tuo et ait Ionadab est si est inquit da manum tuam qui dedit manum suam at ille levavit eum ad se in curru
2KGS|10|16|dixitque ad eum veni mecum et vide zelum meum pro Domino et inpositum currui suo
2KGS|10|17|duxit in Samariam et percussit omnes qui reliqui fuerant de Ahab in Samaria usque ad unum iuxta verbum Domini quod locutus est per Heliam
2KGS|10|18|congregavit ergo Hieu omnem populum et dixit ad eos Ahab coluit Baal parum ego autem colam eum amplius
2KGS|10|19|nunc igitur omnes prophetas Baal et universos servos eius et cunctos sacerdotes ipsius vocate ad me nullus sit qui non veniat sacrificium enim grande est mihi Baal quicumque defuerit non vivet porro Hieu faciebat hoc insidiose ut disperderet cultores Baal
2KGS|10|20|dixit sanctificate diem sollemnem Baal vocavitque
2KGS|10|21|et misit in universos terminos Israhel et venerunt cuncti servi Baal non fuit residuus ne unus quidem qui non veniret et ingressi sunt templum Baal et repleta est domus Baal a summo usque ad summum
2KGS|10|22|dixitque his qui erant super vestes proferte vestimenta universis servis Baal et protulerunt eis vestes
2KGS|10|23|ingressusque Hieu et Ionadab filius Rechab templum Baal et ait cultoribus Baal perquirite et videte ne quis forte vobiscum sit de servis Domini sed ut sint soli servi Baal
2KGS|10|24|ingressi sunt igitur ut facerent victimas et holocausta Hieu autem praeparaverat sibi foris octoginta viros et dixerat eis quicumque fugerit de hominibus his quos ego adduxero in manus vestras anima eius erit pro anima illius
2KGS|10|25|factum est ergo cum conpletum esset holocaustum praecepit Hieu militibus et ducibus suis ingredimini et percutite eos nullus evadat percusseruntque eos ore gladii et proiecerunt milites et duces et ierunt in civitatem templi Baal
2KGS|10|26|et protulerunt statuam de fano Baal et conbuserunt
2KGS|10|27|et comminuerunt eam destruxerunt quoque aedem Baal et fecerunt pro ea latrinas usque ad diem hanc
2KGS|10|28|delevit itaque Hieu Baal de Israhel
2KGS|10|29|verumtamen a peccatis Hieroboam filii Nabath qui peccare fecerat Israhel non recessit nec dereliquit vitulos aureos qui erant in Bethel et in Dan
2KGS|10|30|dixit autem Dominus ad Hieu quia studiose fecisti quod rectum erat et placebat in oculis meis et omnia quae erant in corde meo fecisti contra domum Ahab filii tui usque ad quartam generationem sedebunt super thronum Israhel
2KGS|10|31|porro Hieu non custodivit ut ambularet in lege Domini Dei Israhel in toto corde suo non enim recessit a peccatis Hieroboam qui peccare fecerat Israhel
2KGS|10|32|in diebus illis coepit Dominus taedere super Israhel percussitque eos Azahel in universis finibus Israhel
2KGS|10|33|a Iordane contra orientalem plagam omnem terram Galaad et Gad et Ruben et Manasse ab Aroer quae est super torrentem Arnon et Galaad et Basan
2KGS|10|34|reliqua autem verborum Hieu et universa quae fecit et fortitudo eius nonne haec scripta sunt in libro verborum dierum regum Israhel
2KGS|10|35|et dormivit Hieu cum patribus suis sepelieruntque eum in Samaria et regnavit Ioachaz filius eius pro eo
2KGS|10|36|dies autem quos regnavit Hieu super Israhel viginti et octo anni sunt in Samaria
2KGS|11|1|Athalia vero mater Ahaziae videns mortuum filium suum surrexit et interfecit omne semen regium
2KGS|11|2|tollens autem Iosaba filia regis Ioram soror Ahaziae Ioas filium Ahaziae furata est eum de medio filiorum regis qui interficiebantur et nutricem eius de triclinio et abscondit eum a facie Athaliae ut non interficeretur
2KGS|11|3|eratque cum ea in domo Domini clam sex annis porro Athalia regnavit super terram
2KGS|11|4|anno autem septimo misit Ioiada et adsumens centuriones et milites introduxit ad se in templum Domini pepigitque cum eis foedus et adiurans eos in domo Domini ostendit eis filium regis
2KGS|11|5|et praecepit illis dicens iste sermo quem facere debetis
2KGS|11|6|tertia pars vestrum introeat sabbato et observet excubitum domus regis tertia autem pars sit ad portam Sir et tertia pars ad portam quae est post habitaculum scutariorum et custodietis excubitum domus Messa
2KGS|11|7|duae vero partes e vobis omnes egredientes sabbato custodiant excubias domus Domini circum regem
2KGS|11|8|et vallabitis eum habentes arma in manibus vestris si quis autem ingressus fuerit septum templi interficiatur eritisque cum rege introeunte et egrediente
2KGS|11|9|et fecerunt centuriones iuxta omnia quae praeceperat eis Ioiada sacerdos et adsumentes singuli viros suos qui ingrediebantur sabbatum cum his qui egrediebantur e sabbato venerunt ad Ioiada sacerdotem
2KGS|11|10|qui dedit eis hastas et arma regis David quae erant in domo Domini
2KGS|11|11|et steterunt singuli habentes arma in manu sua a parte templi dextra usque ad partem sinistram altaris et aedis circum regem
2KGS|11|12|produxitque filium regis et posuit super eum diadema et testimonium feceruntque eum regem et unxerunt et plaudentes manu dixerunt vivat rex
2KGS|11|13|audivit Athalia vocem currentis populi et ingressa ad turbas in templum Domini
2KGS|11|14|vidit regem stantem super tribunal iuxta morem et cantores et tubas propter eum omnemque populum terrae laetantem et canentem tubis et scidit vestimenta sua clamavitque coniuratio coniuratio
2KGS|11|15|praecepit autem Ioiada centurionibus qui erant super exercitum et ait eis educite eam extra consepta templi et quicumque secutus eam fuerit feriatur gladio dixerat enim sacerdos non occidatur in templo Domini
2KGS|11|16|inposueruntque ei manus et inpegerunt eam per viam introitus equorum iuxta palatium et interfecta est ibi
2KGS|11|17|pepigit igitur Ioiada foedus inter Dominum et inter regem et inter populum ut esset populus Domini et inter regem et populum
2KGS|11|18|ingressusque est omnis populus terrae templum Baal et destruxerunt aras eius et imagines contriverunt valide Matthan quoque sacerdotem Baal occiderunt coram altari et posuit sacerdos custodias in domo Domini
2KGS|11|19|tulitque centuriones et Cherethi et Felethi legiones et omnem populum terrae deduxeruntque regem de domo Domini et venerunt per viam portae scutariorum in palatium et sedit super thronum regum
2KGS|11|20|laetatusque est omnis populus terrae et civitas conquievit Athalia autem occisa est gladio in domo regis
2KGS|11|21|septemque annorum erat Ioas cum regnare coepisset
2KGS|12|1|anno septimo Hieu regnavit Ioas quadraginta annis regnavit in Hierusalem nomen matris eius Sebia de Bersabee
2KGS|12|2|fecitque Ioas rectum coram Domino cunctis diebus quibus docuit eum Ioiada sacerdos
2KGS|12|3|verumtamen excelsa non abstulit adhuc populus immolabat et adolebat in excelsis incensum
2KGS|12|4|dixitque Ioas ad sacerdotes omnem pecuniam sanctorum quae inlata fuerit in templum Domini a praetereuntibus quae offertur pro pretio animae et quam sponte et arbitrio cordis sui inferunt in templum Domini
2KGS|12|5|accipiant illam sacerdotes iuxta ordinem suum et instaurent sarta tecta domus si quid necessarium viderint instauratione
2KGS|12|6|igitur usque ad vicesimum tertium annum regis Ioas non instauraverunt sacerdotes sarta tecta templi
2KGS|12|7|vocavitque rex Ioas Ioiada pontificem et sacerdotes dicens eis quare sarta tecta non instaurastis templi nolite ergo amplius accipere pecuniam iuxta ordinem vestrum sed ad instaurationem templi reddite eam
2KGS|12|8|prohibitique sunt sacerdotes ultra accipere pecuniam a populo et instaurare sarta tecta domus
2KGS|12|9|et tulit Ioiada pontifex gazofilacium unum aperuitque foramen desuper et posuit illud iuxta altare ad dexteram ingredientium domum Domini mittebantque in eo sacerdotes qui custodiebant ostia omnem pecuniam quae deferebatur ad templum Domini
2KGS|12|10|cumque viderent nimiam pecuniam esse in gazofilacio ascendebat scriba regis et pontifex effundebantque et numerabant pecuniam quae inveniebatur in domo Domini
2KGS|12|11|et dabant eam iuxta numerum atque mensuram in manu eorum qui praeerant cementariis domus Domini qui inpendebant eam in fabris lignorum et in cementariis his qui operabantur in domo Domini
2KGS|12|12|et sarta tecta faciebant et in his qui caedebant saxa et ut emerent ligna et lapides qui excidebantur ita ut impleretur instauratio domus Domini in universis quae indigebant expensa ad muniendam domum
2KGS|12|13|verumtamen non fiebant ex eadem pecunia hydriae templi Domini et fuscinulae et turibula et tubae omne vas aureum et argenteum de pecunia quae inferebatur in templum Domini
2KGS|12|14|his enim qui faciebant opus dabatur ut instauraretur templum Domini
2KGS|12|15|et non fiebat ratio his hominibus qui accipiebant pecuniam ut distribuerent eam artificibus sed in fide tractabant eam
2KGS|12|16|pecuniam vero pro delicto et pecuniam pro peccatis non inferebant in templum Domini quia sacerdotum erat
2KGS|12|17|tunc ascendit Azahel rex Syriae et pugnabat contra Geth cepitque eam et direxit faciem suam ut ascenderet in Hierusalem
2KGS|12|18|quam ob rem tulit Ioas rex Iuda omnia sanctificata quae consecraverant Iosaphat et Ioram et Ahazia patres eius reges Iuda et quae ipse obtulerat et universum argentum quod inveniri potuit in thesauris templi Domini et in palatio regis misitque Azaheli regi Syriae et recessit ab Hierusalem
2KGS|12|19|reliqua autem sermonum Ioas et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|12|20|surrexerunt autem servi eius et coniuraverunt inter se percusseruntque Ioas in domo Mello in descensu Sela
2KGS|12|21|Iozachar namque filius Semath et Iozabad filius Somer servi eius percusserunt eum et mortuus est et sepelierunt eum cum patribus suis in civitate David regnavitque Amasias filius eius pro eo
2KGS|13|1|anno vicesimo tertio Ioas filii Ahaziae regis Iudae regnavit Ioachaz filius Hieu super Israhel in Samaria decem et septem annis
2KGS|13|2|et fecit malum coram Domino secutusque est peccata Hieroboam filii Nabath qui peccare fecit Israhel non declinavit ab eis
2KGS|13|3|iratusque est furor Domini contra Israhel et tradidit eos in manu Azahelis regis Syriae et in manu Benadad filii Azahel cunctis diebus
2KGS|13|4|deprecatus est autem Ioachaz faciem Domini et audivit eum Dominus vidit enim angustiam Israhel qua adtriverat eos rex Syriae
2KGS|13|5|et dedit Dominus Israheli salvatorem et liberatus est de manu Syriae habitaveruntque filii Israhel in tabernaculis suis sicut heri et nudius tertius
2KGS|13|6|verumtamen non recesserunt a peccatis domus Hieroboam qui peccare fecit Israhel in ipsis ambulaverunt siquidem et lucus permansit in Samaria
2KGS|13|7|et non sunt derelicti Ioachaz de populo nisi quinquaginta equites et decem currus et decem milia peditum interfecerat enim eos rex Syriae et redegerat quasi pulverem in tritura areae
2KGS|13|8|reliqua autem sermonum Ioachaz et universa quae fecit sed et fortitudo eius nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|13|9|dormivitque Ioachaz cum patribus suis et sepelierunt eum in Samaria regnavitque Ioas filius eius pro eo
2KGS|13|10|anno tricesimo septimo Ioas regis Iuda regnavit Ioas filius Ioachaz super Israhel in Samaria sedecim annis
2KGS|13|11|et fecit quod malum est in conspectu Domini non declinavit ab omnibus peccatis Hieroboam filii Nabath qui peccare fecit Israhel in ipsis ambulavit
2KGS|13|12|reliqua autem sermonum Ioas et universa quae fecit sed et fortitudo eius quomodo pugnaverit contra Amasiam regem Iuda nonne haec scripta sunt in libro sermonum regum Israhel
2KGS|13|13|et dormivit Ioas cum patribus suis Hieroboam autem sedit super solium eius porro Ioas sepultus est in Samaria cum regibus Israhel
2KGS|13|14|Heliseus autem aegrotabat infirmitate qua et mortuus est descenditque ad eum Ioas rex Israhel et flebat coram eo dicebatque pater mi pater mi currus Israhel et auriga eius
2KGS|13|15|et ait illi Heliseus adfer arcum et sagittas cumque adtulisset ad eum arcum et sagittas
2KGS|13|16|dixit ad regem Israhel pone manum tuam super arcum et cum posuisset ille manum suam superposuit Heliseus manus suas manibus regis
2KGS|13|17|et ait aperi fenestram orientalem cumque aperuisset dixit Heliseus iace sagittam et iecit et ait Heliseus sagitta salutis Domini et sagitta salutis contra Syriam percutiesque Syriam in Afec donec consumas eam
2KGS|13|18|et ait tolle sagittas qui cum tulisset rursum dixit ei percute iaculo terram et cum percussisset tribus vicibus et stetisset
2KGS|13|19|iratus est contra eum vir Dei et ait si percussisses quinquies aut sexies sive septies percussisses Syriam usque ad consummationem nunc autem tribus vicibus percuties eam
2KGS|13|20|mortuus est ergo Heliseus et sepelierunt eum latrunculi quoque de Moab venerunt in terra in ipso anno
2KGS|13|21|quidam autem sepelientes hominem viderunt latrunculos et proiecerunt cadaver in sepulchro Helisei quod ambulavit et tetigit ossa Helisei et revixit homo et stetit super pedes suos
2KGS|13|22|igitur Azahel rex Syriae adflixit Israhel cunctis diebus Ioachaz
2KGS|13|23|et misertus est Dominus eorum et reversus est ad eos propter pactum suum quod habebat cum Abraham Isaac et Iacob et noluit disperdere eos neque proicere penitus usque in praesens tempus
2KGS|13|24|mortuus est autem Azahel rex Syriae et regnavit Benadad filius eius pro eo
2KGS|13|25|porro Ioas filius Ioachaz tulit urbes de manu Benadad filii Azahel quas tulerat de manu Ioachaz patris sui iure proelii tribus vicibus percussit eum Ioas et reddidit civitates Israheli
2KGS|14|1|anno secundo Ioas filii Ioachaz regis Israhel regnavit Amasias filius Ioas regis Iuda
2KGS|14|2|viginti quinque annorum erat cum regnare coepisset viginti autem et novem annis regnavit in Hierusalem nomen matris eius Ioaden de Hierusalem
2KGS|14|3|et fecit rectum coram Domino verumtamen non ut David pater eius iuxta omnia quae fecit Ioas pater suus fecit
2KGS|14|4|nisi hoc tantum quod excelsa non abstulit adhuc enim populus immolabat et adolebat in excelsis
2KGS|14|5|cumque obtinuisset regnum percussit servos suos qui interfecerant regem patrem suum
2KGS|14|6|filios autem eorum qui occiderant non occidit iuxta quod scriptum est in libro legis Mosi sicut praecepit Dominus dicens non morientur patres pro filiis neque filii morientur pro patribus sed unusquisque in peccato suo morietur
2KGS|14|7|ipse percussit Edom in valle Salinarum decem milia et adprehendit Petram in proelio vocavitque nomen eius Iecethel usque in praesentem diem
2KGS|14|8|tunc misit Amasias nuntios ad Ioas filium Ioachaz filii Hieu regis Israhel dicens veni et videamus nos
2KGS|14|9|remisitque Ioas rex Israhel ad Amasiam regem Iuda dicens carduus Libani misit ad cedrum quae est in Libano dicens da filiam tuam filio meo uxorem transieruntque bestiae saltus quae sunt in Libano et conculcaverunt carduum
2KGS|14|10|percutiens invaluisti super Edom et sublevavit te cor tuum contentus esto gloria et sede in domo tua quare provocas malum ut cadas tu et Iuda tecum
2KGS|14|11|et non adquievit Amasias ascenditque Ioas rex Israhel et viderunt se ipse et Amasias rex Iuda in Bethsames oppido Iudae
2KGS|14|12|percussusque est Iuda coram Israhel et fugerunt unusquisque in tabernacula sua
2KGS|14|13|Amasiam vero regem Iuda filium Ioas filii Ahaziae cepit Ioas rex Israhel in Bethsames et adduxit eum in Hierusalem et interrupit murum Hierusalem a porta Ephraim usque ad portam Anguli quadringentis cubitis
2KGS|14|14|tulitque omne aurum et argentum et universa vasa quae inventa sunt in domo Domini et in thesauris regis et obsides et reversus est Samariam
2KGS|14|15|reliqua autem verborum Ioas quae fecit et fortitudo eius qua pugnavit contra Amasiam regem Iuda nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|14|16|dormivitque Ioas cum patribus suis et sepultus est in Samaria cum regibus Israhel et regnavit Hieroboam filius eius pro eo
2KGS|14|17|vixit autem Amasias filius Ioas rex Iuda postquam mortuus est Ioas filius Ioachaz regis Israhel viginti quinque annis
2KGS|14|18|reliqua autem sermonum Amasiae nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|14|19|factaque est contra eum coniuratio in Hierusalem at ille fugit in Lachis miseruntque post eum in Lachis et interfecerunt eum ibi
2KGS|14|20|et asportaverunt in equis sepultusque est in Hierusalem cum patribus suis in civitate David
2KGS|14|21|tulit autem universus populus Iudae Azariam annos natum sedecim et constituerunt eum regem pro patre eius Amasia
2KGS|14|22|ipse aedificavit Ahilam et restituit eam Iudae postquam dormivit rex cum patribus suis
2KGS|14|23|anno quintodecimo Amasiae filii Ioas regis Iuda regnavit Hieroboam filius Ioas regis Israhel in Samaria quadraginta et uno anno
2KGS|14|24|et fecit quod malum est coram Domino non recessit ab omnibus peccatis Hieroboam filii Nabath qui peccare fecit Israhel
2KGS|14|25|ipse restituit terminos Israhel ab introitu Emath usque ad mare Solitudinis iuxta sermonem Domini Dei Israhel quem locutus est per servum suum Ionam filium Amathi prophetam qui erat de Geth quae est in Opher
2KGS|14|26|vidit enim Dominus adflictionem Israhel amaram nimis et quod consumpti essent usque ad clausos carcere et extremos et non esset qui auxiliaretur Israhel
2KGS|14|27|nec locutus est Dominus ut deleret nomen Israhel sub caelo sed salvavit eos in manu Hieroboam filii Ioas
2KGS|14|28|reliqua autem sermonum Hieroboam et universa quae fecit et fortitudo eius qua proeliatus est et quomodo restituit Damascum et Emath Iudae in Israhel nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|14|29|dormivitque Hieroboam cum patribus suis regibus Israhel et regnavit Zaccharias filius eius pro eo
2KGS|15|1|anno vicesimo septimo Hieroboam regis Israhel regnavit Azarias filius Amasiae regis Iudae
2KGS|15|2|sedecim annorum erat cum regnare coepisset et quinquaginta duobus annis regnavit in Hierusalem nomen matris eius Iecelia de Hierusalem
2KGS|15|3|fecitque quod erat placitum coram Domino iuxta omnia quae fecit Amasias pater eius
2KGS|15|4|verumtamen excelsa non est demolitus adhuc populus sacrificabat et adolebat incensum in excelsis
2KGS|15|5|percussit autem Dominus regem et fuit leprosus usque in diem mortis suae et habitabat in domo libera seorsum Ioatham vero filius regis gubernabat palatium et iudicabat populum terrae
2KGS|15|6|reliqua autem sermonum Azariae et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|15|7|et dormivit Azarias cum patribus suis sepelieruntque eum cum maioribus suis in civitate David et regnavit Ioatham filius eius pro eo
2KGS|15|8|anno tricesimo octavo Azariae regis Iudae regnavit Zaccharias filius Hieroboam super Israhel in Samaria sex mensibus
2KGS|15|9|et fecit quod malum est coram Domino sicut fecerant patres eius non recessit a peccatis Hieroboam filii Nabath qui peccare fecit Israhel
2KGS|15|10|coniuravit autem contra eum Sellum filius Iabes percussitque eum palam et interfecit regnavitque pro eo
2KGS|15|11|reliqua autem verborum Zacchariae nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|12|ipse est sermo Domini quem locutus est ad Hieu dicens filii usque ad quartam generationem sedebunt de te super thronum Israhel factumque est ita
2KGS|15|13|Sellum filius Iabes regnavit tricesimo nono anno Azariae regis Iudae regnavit autem uno mense in Samaria
2KGS|15|14|et ascendit Manahem filius Gaddi de Thersa venitque Samariam et percussit Sellum filium Iabes in Samaria et interfecit eum regnavitque pro eo
2KGS|15|15|reliqua autem verborum Sellum et coniuratio eius per quam tetendit insidias nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|16|tunc percussit Manahem Thapsam et omnes qui erant in ea et terminos eius de Thersa noluerant enim aperire ei et interfecit omnes praegnantes eius et scidit eas
2KGS|15|17|anno tricesimo nono Azariae regis Iuda regnavit Manahem filius Gaddi super Israhel decem annis in Samaria
2KGS|15|18|fecitque quod erat malum coram Domino non recessit a peccatis Hieroboam filii Nabath qui peccare fecit Israhel cunctis diebus eius
2KGS|15|19|veniebat Phul rex Assyriorum in terram et dabat Manahem Phul mille talenta argenti ut esset ei in auxilio et firmaret regnum eius
2KGS|15|20|indixitque Manahem argentum super Israhel cunctis potentibus et divitibus ut daret regi Assyriorum quinquaginta siclos argenti per singulos reversusque est rex Assyriorum et non est moratus in terra
2KGS|15|21|reliqua autem sermonum Manahem et universa quae fecit nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|22|et dormivit Manahem cum patribus suis regnavitque Phaceia filius eius pro eo
2KGS|15|23|anno quinquagesimo Azariae regis Iudae regnavit Phaceia filius Manahem super Israhel in Samaria biennio
2KGS|15|24|et fecit quod erat malum coram Domino non recessit a peccatis Hieroboam filii Nabath qui peccare fecit Israhel
2KGS|15|25|coniuravit autem adversum eum Phacee filius Romeliae dux eius et percussit eum in Samaria in turre domus regiae iuxta Argob et iuxta Ari et cum eo quinquaginta viros de filiis Galaaditarum et interfecit eum regnavitque pro eo
2KGS|15|26|reliqua autem sermonum Phaceia et universa quae fecit nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|27|anno quinquagesimo secundo Azariae regis Iudae regnavit Phacee filius Romeliae super Israhel in Samaria viginti annis
2KGS|15|28|et fecit quod malum erat coram Domino non recessit a peccatis Hieroboam filii Nabath qui peccare fecit Israhel
2KGS|15|29|in diebus Phacee regis Israhel venit Theglathfalassar rex Assur et cepit Aiom et Abel domum Maacha et Ianoe et Cedes et Asor et Galaad et Galileam universam terram Nepthalim et transtulit eos in Assyrios
2KGS|15|30|coniuravit autem et tetendit insidias Osee filius Hela contra Phacee filium Romeliae et percussit eum et interfecit regnavitque pro eo vicesimo anno Ioatham filii Oziae
2KGS|15|31|reliqua autem sermonum Phacee et universa quae fecit nonne haec scripta sunt in libro sermonum dierum regum Israhel
2KGS|15|32|anno secundo Phacee filii Romeliae regis Israhel regnavit Ioatham filius Oziae regis Iuda
2KGS|15|33|viginti quinque annorum erat cum regnare coepisset et sedecim annis regnavit in Hierusalem nomen matris eius Hierusa filia Sadoc
2KGS|15|34|fecitque quod erat placitum coram Domino iuxta omnia quae fecerat Ozias pater suus operatus est
2KGS|15|35|verumtamen excelsa non abstulit adhuc populus immolabat et adolebat incensum in excelsis ipse aedificavit portam domus Domini sublimissimam
2KGS|15|36|reliqua autem sermonum Ioatham et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|15|37|in diebus illis coepit Dominus mittere in Iudam Rasin regem Syriae et Phacee filium Romeliae
2KGS|15|38|et dormivit Ioatham cum patribus suis sepultusque est cum eis in civitate David patris sui et regnavit Ahaz filius eius pro eo
2KGS|16|1|anno septimodecimo Phacee filii Romeliae regnavit Ahaz filius Ioatham regis Iuda
2KGS|16|2|viginti annorum erat Ahaz cum regnare coepisset et sedecim annis regnavit in Hierusalem non fecit quod erat placitum in conspectu Domini Dei sui sicut David pater eius
2KGS|16|3|sed ambulavit in via regum Israhel insuper et filium suum consecravit transferens per ignem secundum idola gentium quae dissipavit Dominus coram filiis Israhel
2KGS|16|4|immolabat quoque victimas et adolebat incensum in excelsis et in collibus et sub omni ligno frondoso
2KGS|16|5|tunc ascendit Rasin rex Syriae et Phacee filius Romeliae rex Israhel in Hierusalem ad proeliandum cumque obsiderent Ahaz non valuerunt superare eum
2KGS|16|6|in tempore illo restituit Rasin rex Syriae Ahilam Syriae et eiecit Iudaeos de Ahilam et Idumei venerunt in Ahilam et habitaverunt ibi usque in diem hanc
2KGS|16|7|misit autem Ahaz nuntios ad Theglathfalassar regem Assyriorum dicens servus tuus et filius tuus ego sum ascende et salvum me fac de manu regis Syriae et de manu regis Israhel qui consurrexerunt adversum me
2KGS|16|8|et cum collegisset argentum et aurum quod invenire potuit in domo Domini et in thesauris regis misit regi Assyriorum munera
2KGS|16|9|qui et adquievit voluntati eius ascendit enim rex Assyriorum in Damascum et vastavit eam et transtulit habitatores eius Cyrenen Rasin autem interfecit
2KGS|16|10|perrexitque rex Ahaz in occursum Theglathfalassar regis Assyriorum in Damascum cumque vidisset altare Damasci misit rex Ahaz ad Uriam sacerdotem exemplar eius et similitudinem iuxta omne opus eius
2KGS|16|11|extruxitque Urias sacerdos altare iuxta omnia quae praeceperat rex Ahaz de Damasco ita fecit Urias sacerdos donec veniret rex Ahaz de Damasco
2KGS|16|12|cumque venisset rex de Damasco vidit altare et veneratus est illud ascenditque et immolavit holocausta et sacrificium suum
2KGS|16|13|et libavit libamina et fudit sanguinem pacificorum quae obtulerat super altare
2KGS|16|14|porro altare aeneum quod erat coram Domino transtulit de facie templi et de loco altaris et de loco templi Domini posuitque illud ex latere altaris ad aquilonem
2KGS|16|15|praecepit quoque rex Ahaz Uriae sacerdoti dicens super altare maius offer holocaustum matutinum et sacrificium vespertinum et holocaustum regis et sacrificium eius et holocaustum universi populi terrae et sacrificia eorum et libamina eorum et omnem sanguinem holocausti et universum sanguinem victimae super illud effundes altare vero aeneum erit paratum ad voluntatem meam
2KGS|16|16|fecit igitur Urias sacerdos iuxta omnia quae praeceperat rex Ahaz
2KGS|16|17|tulit autem rex Ahaz celatas bases et luterem qui erat desuper et mare deposuit de bubus aeneis qui sustentabant illud et posuit super pavimentum stratum lapide
2KGS|16|18|Musach quoque sabbati quod aedificaverat in templo et ingressum regis exterius convertit in templo Domini propter regem Assyriorum
2KGS|16|19|reliqua autem verborum Ahaz quae fecit nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|16|20|dormivitque Ahaz cum patribus suis et sepultus est cum eis in civitate David et regnavit Ezechias filius eius pro eo
2KGS|17|1|anno duodecimo Ahaz regis Iuda regnavit Osee filius Hela in Samaria super Israhel novem annis
2KGS|17|2|fecitque malum coram Domino sed non sicut reges Israhel qui ante eum fuerant
2KGS|17|3|contra hunc ascendit Salmanassar rex Assyriorum et factus est ei Osee servus reddebatque illi tributa
2KGS|17|4|cumque deprehendisset rex Assyriorum Osee quod rebellare nitens misisset nuntios ad Sua regem Aegypti ne praestaret tributa regi Assyriorum sicut singulis annis solitus erat obsedit eum et vinctum misit in carcerem
2KGS|17|5|pervagatusque est omnem terram et ascendens Samariam obsedit eam tribus annis
2KGS|17|6|anno autem nono Osee cepit rex Assyriorum Samariam et transtulit Israhel in Assyrios posuitque eos in Ala et in Habor iuxta fluvium Gozan in civitatibus Medorum
2KGS|17|7|factum est enim cum peccassent filii Israhel Domino Deo suo qui eduxerat eos de terra Aegypti de manu Pharaonis regis Aegypti coluerunt deos alienos
2KGS|17|8|et ambulaverunt iuxta ritum gentium quas consumpserat Dominus in conspectu filiorum Israhel et regum Israhel quia similiter fecerant
2KGS|17|9|et operuerunt filii Israhel verbis non rectis Dominum Deum suum et aedificaverunt sibi excelsa in cunctis urbibus suis a turre custodum usque ad civitatem munitam
2KGS|17|10|feceruntque sibi statuas et lucos in omni colle sublimi et subter omne lignum nemorosum
2KGS|17|11|et adolebant ibi incensum super aras in more gentium quas transtulerat Dominus a facie eorum feceruntque verba pessima inritantes Dominum
2KGS|17|12|et coluerunt inmunditias de quibus praecepit Dominus eis ne facerent verbum hoc
2KGS|17|13|et testificatus est Dominus in Israhel et in Iuda per manum omnium prophetarum et videntum dicens revertimini a viis vestris pessimis et custodite praecepta mea et caerimonias iuxta omnem legem quam praecepi patribus vestris et sicut misi ad vos in manu servorum meorum prophetarum
2KGS|17|14|qui non audierunt sed induraverunt cervicem suam iuxta cervicem patrum suorum qui noluerunt oboedire Domino Deo suo
2KGS|17|15|et abiecerunt legitima eius et pactum quod pepigit cum patribus eorum et testificationes quibus contestatus est eos secutique sunt vanitates et vane egerunt et secuti sunt gentes quae erant per circuitum eorum super quibus praeceperat Dominus eis ut non facerent sicut et illae faciebant
2KGS|17|16|et dereliquerunt omnia praecepta Domini Dei sui feceruntque sibi conflatiles duos vitulos et lucos et adoraverunt universam militiam caeli servieruntque Baal
2KGS|17|17|et consecrabant ei filios suos et filias suas per ignem et divinationibus inserviebant et auguriis et tradiderunt se ut facerent malum coram Domino et inritarent eum
2KGS|17|18|iratusque est Dominus vehementer Israhel et abstulit eos de conspectu suo et non remansit nisi tribus Iuda tantummodo
2KGS|17|19|sed nec ipse Iuda custodivit mandata Domini Dei sui verum ambulavit in erroribus Israhel quos operatus fuerat
2KGS|17|20|proiecitque Dominus omne semen Israhel et adflixit eos et tradidit in manu diripientium donec proiceret eos a facie sua
2KGS|17|21|ex eo iam tempore quo scissus est Israhel a domo David et constituerunt sibi regem Hieroboam filium Nabath separavit enim Hieroboam Israhel a Domino et peccare eos fecit peccatum magnum
2KGS|17|22|et ambulaverunt filii Israhel in universis peccatis Hieroboam quae fecerat non recesserunt ab eis
2KGS|17|23|usquequo auferret Dominus Israhel a facie sua sicut locutus fuerat in manu omnium servorum suorum prophetarum translatusque est Israhel de terra sua in Assyrios usque in diem hanc
2KGS|17|24|adduxit autem rex Assyriorum de Babylone et de Chutha et de Haiath et de Emath et de Sepharvaim et conlocavit eos in civitatibus Samariae pro filiis Israhel qui possederunt Samariam et habitaverunt in urbibus eius
2KGS|17|25|cumque ibi habitare coepissent non timebant Dominum et inmisit eis Dominus leones qui interficiebant eos
2KGS|17|26|nuntiatumque est regi Assyriorum et dictum gentes quas transtulisti et habitare fecisti in civitatibus Samariae ignorant legitima Dei terrae et inmisit in eos Dominus leones et ecce interficiunt eos eo quod ignorent ritum Dei terrae
2KGS|17|27|praecepit autem rex Assyriorum dicens ducite illuc unum de sacerdotibus quos inde captivos adduxistis et vadat et habitet cum eis et doceat eos legitima Dei terrae
2KGS|17|28|igitur cum venisset unus de sacerdotibus his qui captivi ducti fuerant de Samaria habitavit in Bethel et docebat eos quomodo colerent Dominum
2KGS|17|29|et unaquaeque gens fabricata est deum suum posueruntque eos in fanis excelsis quae fecerant Samaritae gens et gens in urbibus suis in quibus habitabant
2KGS|17|30|viri enim babylonii fecerunt Socchothbenoth viri autem chutheni fecerunt Nergel et viri de Emath fecerunt Asima
2KGS|17|31|porro Evei fecerunt Nebaaz et Tharthac hii autem qui erant de Sepharvaim conburebant filios suos igni Adramelech et Anamelech diis Sepharvaim
2KGS|17|32|et nihilominus colebant Dominum fecerunt autem sibi de novissimis sacerdotes excelsorum et ponebant eos in fanis sublimibus
2KGS|17|33|et cum Dominum colerent diis quoque suis serviebant iuxta consuetudinem gentium de quibus translati fuerant Samariam
2KGS|17|34|usque in praesentem diem morem sequuntur antiquum non timent Dominum neque custodiunt caerimonias eius et iudicia et legem et mandatum quod praeceperat Dominus filiis Iacob quem cognominavit Israhel
2KGS|17|35|et percusserat cum eis pactum et mandaverat eis dicens nolite timere deos alienos et non adoretis eos neque colatis et non immoletis eis
2KGS|17|36|sed Dominum Deum vestrum qui eduxit vos de terra Aegypti in fortitudine magna et in brachio extento ipsum timete illum adorate et ipsi immolate
2KGS|17|37|caerimonias quoque et iudicia et legem et mandatum quod scripsit vobis custodite ut faciatis cunctis diebus et non timeatis deos alienos
2KGS|17|38|et pactum quod percussi vobiscum nolite oblivisci nec colatis deos alienos
2KGS|17|39|sed Dominum Deum vestrum timete et ipse eruet vos de manu omnium inimicorum vestrorum
2KGS|17|40|illi vero non audierunt sed iuxta consuetudinem suam pristinam perpetrabant
2KGS|17|41|fuerunt igitur gentes istae timentes quidem Dominum sed nihilominus et idolis suis servientes nam et filii eorum et nepotes sicut fecerunt parentes sui ita faciunt usque in praesentem diem
2KGS|18|1|anno tertio Osee filii Hela regis Israhel regnavit Ezechias filius Ahaz regis Iuda
2KGS|18|2|viginti quinque annorum erat cum regnare coepisset et viginti et novem annis regnavit in Hierusalem nomen matris eius Abi filia Zacchariae
2KGS|18|3|fecitque quod erat bonum coram Domino iuxta omnia quae fecerat David pater suus
2KGS|18|4|ipse dissipavit excelsa et contrivit statuas et succidit lucos confregitque serpentem aeneum quem fecerat Moses siquidem usque ad illud tempus filii Israhel adolebant ei incensum vocavitque eum Naasthan
2KGS|18|5|in Domino Deo Israhel speravit itaque post eum non fuit similis ei de cunctis regibus Iuda sed neque in his qui ante eum fuerunt
2KGS|18|6|et adhesit Domino et non recessit a vestigiis eius fecitque mandata eius quae praeceperat Dominus Mosi
2KGS|18|7|unde et erat Dominus cum eo et in cunctis ad quae procedebat sapienter se agebat rebellavit quoque contra regem Assyriorum et non servivit ei
2KGS|18|8|ipse percussit Philistheos usque Gazam et omnes terminos eorum a turre custodum usque ad civitatem muratam
2KGS|18|9|anno quarto regis Ezechiae qui erat annus septimus Osee filii Hela regis Israhel ascendit Salmanassar rex Assyriorum Samariam et obpugnavit eam
2KGS|18|10|et cepit nam post annos tres anno sexto Ezechiae id est nono anno Osee regis Israhel capta est Samaria
2KGS|18|11|et transtulit rex Assyriorum Israhel in Assyrios conlocavitque eos in Ala et in Habor fluviis Gozan in civitatibus Medorum
2KGS|18|12|quia non audierunt vocem Domini Dei sui sed praetergressi sunt pactum eius omnia quae praeceperat Moses servus Domini non audierunt neque fecerunt
2KGS|18|13|anno quartodecimo regis Ezechiae ascendit Sennacherib rex Assyriorum ad universas civitates Iuda munitas et cepit eas
2KGS|18|14|tunc misit Ezechias rex Iuda nuntios ad regem Assyriorum Lachis dicens peccavi recede a me et omne quod inposueris mihi feram indixit itaque rex Assyriorum Ezechiae regi Iudae trecenta talenta argenti et triginta talenta auri
2KGS|18|15|deditque Ezechias omne argentum quod reppertum fuerat in domo Domini et in thesauris regis
2KGS|18|16|in tempore illo confregit Ezechias valvas templi Domini et lamminas auri quas ipse adfixerat et dedit eas regi Assyriorum
2KGS|18|17|misit autem rex Assyriorum Tharthan et Rabsaris et Rabsacen de Lachis ad regem Ezechiam cum manu valida Hierusalem qui cum ascendissent venerunt in Hierusalem et steterunt iuxta aquaeductum piscinae superioris quae est in via agri Fullonis
2KGS|18|18|vocaveruntque regem egressus est autem ad eos Eliachim filius Helciae praepositus domus et Sobna scriba et Ioahe filius Asaph a commentariis
2KGS|18|19|dixitque ad eos Rabsaces loquimini Ezechiae haec dicit rex magnus rex Assyriorum quae est ista fiducia qua niteris
2KGS|18|20|forsitan inisti consilium ut praepares te ad proelium in quo confidis ut audeas rebellare
2KGS|18|21|an speras in baculo harundineo atque confracto Aegypto super quem si incubuerit homo comminutus ingreditur manum eius et perforabit eam sic est Pharao rex Aegypti omnibus qui confidunt in se
2KGS|18|22|quod si dixeritis mihi in Domino Deo nostro habemus fiduciam nonne iste est cuius abstulit Ezechias excelsa et altaria et praecepit Iudae et Hierusalem ante altare hoc adorabitis in Hierusalem
2KGS|18|23|nunc igitur transite ad dominum meum regem Assyriorum et dabo vobis duo milia equorum et videte an habere valeatis ascensores eorum
2KGS|18|24|et quomodo potestis resistere ante unum satrapam de servis domini mei minimis an fiduciam habes in Aegypto propter currus et equites
2KGS|18|25|numquid sine Domini voluntate ascendi ad locum istum ut demolirer eum Dominus dixit mihi ascende ad terram hanc et demolire eam
2KGS|18|26|dixerunt autem Eliachim filius Helciae et Sobna et Ioahe Rabsaci precamur ut loquaris nobis servis tuis syriace siquidem intellegimus hanc linguam et non loquaris nobis iudaice audiente populo qui est super murum
2KGS|18|27|responditque eis Rabsaces numquid ad dominum tuum et ad te misit me dominus meus ut loquerer sermones hos et non ad viros qui sedent super murum ut comedant stercora sua et bibant urinam suam vobiscum
2KGS|18|28|stetit itaque Rabsaces et clamavit voce magna iudaice et ait audite verba regis magni regis Assyriorum
2KGS|18|29|haec dicit rex non vos seducat Ezechias non enim poterit eruere vos de manu mea
2KGS|18|30|neque fiduciam vobis tribuat super Domino dicens eruens liberabit nos Dominus et non tradetur civitas haec in manu regis Assyriorum
2KGS|18|31|nolite audire Ezechiam haec enim dicit rex Assyriorum facite mecum quod vobis est utile et egredimini ad me et comedet unusquisque de vinea sua et de ficu sua et bibetis aquas de cisternis vestris
2KGS|18|32|donec veniam et transferam vos in terram quae similis terrae vestrae est in terram fructiferam et fertilem vini terram panis et vinearum terram olivarum et olei ac mellis et vivetis et non moriemini nolite audire Ezechiam qui vos decipit dicens Dominus liberabit nos
2KGS|18|33|numquid liberaverunt dii gentium terram suam de manu regis Assyriorum
2KGS|18|34|ubi est deus Emath et Arfad ubi est deus Sepharvaim Ana et Ava numquid liberaverunt Samariam de manu mea
2KGS|18|35|quinam illi sunt in universis diis terrarum qui eruerunt regionem suam de manu mea ut possit eruere Dominus Hierusalem de manu mea
2KGS|18|36|tacuit itaque populus et non respondit ei quicquam siquidem praeceptum regis acceperant ut non responderent ei
2KGS|18|37|venitque Eliachim filius Helciae praepositus domus et Sobna scriba et Ioahe filius Asaph a commentariis ad Ezechiam scissis vestibus et nuntiaverunt ei verba Rabsacis
2KGS|19|1|quae cum audisset rex Ezechias scidit vestimenta sua et opertus est sacco ingressusque est domum Domini
2KGS|19|2|et misit Eliachim praepositum domus et Sobnam scribam et senes de sacerdotibus opertos saccis ad Esaiam prophetam filium Amos
2KGS|19|3|qui dixerunt haec dicit Ezechias dies tribulationis et increpationis et blasphemiae dies iste venerunt filii usque ad partum et vires non habet parturiens
2KGS|19|4|si forte audiat Dominus Deus tuus universa verba Rabsacis quem misit rex Assyriorum dominus suus ut exprobraret Deum viventem et argueret verbis quae audivit Dominus Deus tuus et fac orationem pro reliquiis quae reppertae sunt
2KGS|19|5|venerunt ergo servi regis Ezechiae ad Esaiam
2KGS|19|6|dixitque eis Esaias haec dicetis domino vestro haec dicit Dominus noli timere a facie sermonum quos audisti quibus blasphemaverunt pueri regis Assyriorum me
2KGS|19|7|ecce ego inmittam ei spiritum et audiet nuntium et revertetur in terram suam et deiciam eum gladio in terra sua
2KGS|19|8|reversus est igitur Rabsaces et invenit regem Assyriorum expugnantem Lobnam audierat enim quod recessisset de Lachis
2KGS|19|9|cumque audisset de Tharaca rege Aethiopiae dicentes ecce egressus est ut pugnet adversum te et iret contra eum misit nuntios ad Ezechiam dicens
2KGS|19|10|haec dicite Ezechiae regi Iudae non te seducat Deus tuus in quo habes fiduciam neque dicas non tradetur Hierusalem in manu regis Assyriorum
2KGS|19|11|tu enim ipse audisti quae fecerint reges Assyriorum universis terris quomodo vastaverint eas num ergo solus poteris liberari
2KGS|19|12|numquid liberaverunt dii gentium singulos quos vastaverunt patres mei Gozan videlicet et Aran et Reseph et filios Eden qui erant in Thelassar
2KGS|19|13|ubi est rex Emath et rex Arfad et rex civitatis Sepharvaim Ana et Ava
2KGS|19|14|itaque cum accepisset Ezechias litteras de manu nuntiorum et legisset eas ascendit in domum Domini et expandit eas coram Domino
2KGS|19|15|et oravit in conspectu eius dicens Domine Deus Israhel qui sedes super cherubin tu es Deus solus regum omnium terrae tu fecisti caelum et terram
2KGS|19|16|inclina aurem tuam et audi aperi Domine oculos tuos et vide et audi omnia verba Sennacherib qui misit ut exprobraret nobis Deum viventem
2KGS|19|17|vere Domine dissipaverunt reges Assyriorum gentes et terras omnium
2KGS|19|18|et miserunt deos eorum in ignem non enim erant dii sed opera manuum hominum e ligno et lapide et perdiderunt eos
2KGS|19|19|nunc igitur Domine Deus noster salvos nos fac de manu eius ut sciant omnia regna terrae quia tu es Dominus Deus solus
2KGS|19|20|misit autem Esaias filius Amos ad Ezechiam dicens haec dicit Dominus Deus Israhel quae deprecatus es me super Sennacherib rege Assyriorum audivi
2KGS|19|21|iste est sermo quem locutus est Dominus de eo sprevit te et subsannavit virgo filia Sion post tergum tuum caput movit filia Hierusalem
2KGS|19|22|cui exprobrasti et quem blasphemasti contra quem exaltasti vocem et elevasti in excelsum oculos tuos contra Sanctum Israhel
2KGS|19|23|per manum servorum tuorum exprobrasti Domino et dixisti in multitudine curruum meorum ascendi excelsa montium in summitate Libani et succidi sublimes cedros eius electas abietes eius et ingressus sum usque ad terminos eius saltum Carmeli eius
2KGS|19|24|ego succidi et bibi aquas alienas et siccavi vestigiis pedum meorum omnes aquas clausas
2KGS|19|25|numquid non audisti quid ab initio fecerim ex diebus antiquis plasmavi illud et nunc adduxi eruntque in ruinam collium pugnantium civitates munitae
2KGS|19|26|et qui sedent in eis humiles manu contremuerunt et confusi sunt facti sunt quasi faenum agri et virens herba tectorum quae arefacta est antequam veniret ad maturitatem
2KGS|19|27|habitaculum tuum et egressum tuum et viam tuam ego praescivi et furorem tuum contra me
2KGS|19|28|insanisti in me et superbia tua ascendit in aures meas ponam itaque circulum in naribus tuis et camum in labris tuis et reducam te in viam per quam venisti
2KGS|19|29|tibi autem Ezechia hoc erit signum comede hoc anno quod reppereris in secundo autem anno quae sponte nascuntur porro in anno tertio seminate et metite plantate vineas et comedite fructum earum
2KGS|19|30|et quodcumque reliquum fuerit de domo Iuda mittet radicem deorsum et faciet fructum sursum
2KGS|19|31|de Hierusalem quippe egredientur reliquiae et quod salvetur de monte Sion zelus Domini exercituum faciet hoc
2KGS|19|32|quam ob rem haec dicit Dominus de rege Assyriorum non ingredietur urbem hanc nec mittet in eam sagittam nec occupabit eam clypeus nec circumdabit eam munitio
2KGS|19|33|per viam qua venit revertetur et civitatem hanc non ingredietur dicit Dominus
2KGS|19|34|protegamque urbem hanc et salvabo eam propter me et propter David servum meum
2KGS|19|35|factum est igitur in nocte illa venit angelus Domini et percussit castra Assyriorum centum octoginta quinque milia cumque diluculo surrexisset vidit omnia corpora mortuorum et recedens abiit
2KGS|19|36|et reversus est Sennacherib rex Assyriorum et mansit in Nineve
2KGS|19|37|cumque adoraret in templo Neserach deum suum Adramelech et Sarasar filii eius percusserunt eum gladio fugeruntque in terram Armeniorum et regnavit Eseraddon filius eius pro eo
2KGS|20|1|in diebus illis aegrotavit Ezechias usque ad mortem et venit ad eum Esaias filius Amos prophetes dixitque ei haec dicit Dominus Deus praecipe domui tuae morieris enim et non vives
2KGS|20|2|qui convertit faciem suam ad parietem et oravit Dominum dicens
2KGS|20|3|obsecro Domine memento quomodo ambulaverim coram te in veritate et in corde perfecto et quod placitum est coram te fecerim flevit itaque Ezechias fletu magno
2KGS|20|4|et antequam egrederetur Esaias mediam partem atrii factus est sermo Domini ad eum dicens
2KGS|20|5|revertere et dic Ezechiae duci populi mei haec dicit Dominus Deus David patris tui audivi orationem tuam vidi lacrimam tuam et ecce sanavi te die tertio ascendes templum Domini
2KGS|20|6|et addam diebus tuis quindecim annos sed et de manu regis Assyriorum liberabo te et civitatem hanc et protegam urbem istam propter me et propter David servum meum
2KGS|20|7|dixitque Esaias adferte massam ficorum quam cum adtulissent et posuissent super ulcus eius curatus est
2KGS|20|8|dixerat autem Ezechias ad Esaiam quod erit signum quia Dominus me sanabit et quia ascensurus sum die tertio templum Domini
2KGS|20|9|cui ait Esaias hoc erit signum a Domino quod facturus sit Dominus sermonem quem locutus est vis ut accedat umbra decem lineis an ut revertatur totidem gradibus
2KGS|20|10|et ait Ezechias facile est umbram crescere decem lineis nec hoc volo ut fiat sed ut revertatur retrorsum decem gradibus
2KGS|20|11|invocavit itaque Esaias propheta Dominum et reduxit umbram per lineas quibus iam descenderat in horologio Ahaz retrorsum decem gradibus
2KGS|20|12|in tempore illo misit Berodach Baladan filius Baladan rex Babyloniorum litteras et munera ad Ezechiam audierat enim quod aegrotasset Ezechias
2KGS|20|13|laetatus est autem in adventum eorum Ezechias et ostendit eis domum aromatum et aurum et argentum et pigmenta varia unguenta quoque et domum vasorum suorum et omnia quae habere potuerat in thesauris suis non fuit quod non monstraret eis Ezechias in domo sua et in omni potestate sua
2KGS|20|14|venit autem Esaias propheta ad regem Ezechiam dixitque ei quid dixerunt viri isti aut unde venerunt ad te cui ait Ezechias de terra longinqua venerunt de Babylone
2KGS|20|15|at ille respondit quid viderunt in domo tua ait Ezechias omnia quae sunt in domo mea viderunt nihil est quod non monstraverim eis in thesauris meis
2KGS|20|16|dixit itaque Esaias Ezechiae audi sermonem Domini
2KGS|20|17|ecce dies venient et auferentur omnia quae sunt in domo tua et quae condiderunt patres tui usque in diem hanc in Babylone non remanebit quicquam ait Dominus
2KGS|20|18|sed et de filiis tuis qui egredientur ex te quos generabis tollentur et erunt eunuchi in palatio regis Babylonis
2KGS|20|19|dixit Ezechias ad Esaiam bonus sermo Domini quem locutus est sit pax et veritas in diebus meis
2KGS|20|20|reliqua autem sermonum Ezechiae et omnis fortitudo eius et quomodo fecerit piscinam et aquaeductum et introduxerit aquas in civitatem nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|20|21|dormivitque Ezechias cum patribus suis et regnavit Manasses filius eius pro eo
2KGS|21|1|duodecim annorum erat Manasses cum regnare coepisset et quinquaginta quinque annis regnavit in Hierusalem nomen matris eius Aphsiba
2KGS|21|2|fecitque malum in conspectu Domini iuxta idola gentium quas delevit Dominus a facie filiorum Israhel
2KGS|21|3|conversusque est et aedificavit excelsa quae dissipaverat Ezechias pater eius et erexit aras Baal et fecit lucos sicut fecerat Ahab rex Israhel et adoravit omnem militiam caeli et coluit eam
2KGS|21|4|extruxitque aras in domo Domini de qua dixit Dominus in Hierusalem ponam nomen meum
2KGS|21|5|et extruxit altaria universae militiae caeli in duobus atriis templi Domini
2KGS|21|6|et transduxit filium suum per ignem et ariolatus est et observavit auguria et fecit pythones et aruspices multiplicavit ut faceret malum coram Domino et inritaret eum
2KGS|21|7|posuit quoque idolum luci quem fecerat in templo Domini super quo locutus est Dominus ad David et ad Salomonem filium eius in templo hoc et in Hierusalem quam elegi de cunctis tribubus Israhel ponam nomen meum in sempiternum
2KGS|21|8|et ultra non faciam commoveri pedem Israhel de terra quam dedi patribus eorum sic tamen si custodierint opere omnia quae praecepi eis et universam legem quam mandavit eis servus meus Moses
2KGS|21|9|illi vero non audierunt sed seducti sunt a Manasse ut facerent malum super gentes quas contrivit Dominus a facie filiorum Israhel
2KGS|21|10|locutusque est Dominus in manu servorum suorum prophetarum dicens
2KGS|21|11|quia fecit Manasses rex Iuda abominationes istas pessimas super omnia quae fecerunt Amorrei ante eum et peccare fecit etiam Iudam in inmunditiis suis
2KGS|21|12|propterea haec dicit Dominus Deus Israhel ecce ego inducam mala super Hierusalem et Iudam ut quicumque audierit tinniant ambae aures eius
2KGS|21|13|et extendam super Hierusalem funiculum Samariae et pondus domus Ahab et delebo Hierusalem sicut deleri solent tabulae delens vertam et ducam crebrius stilum super faciem eius
2KGS|21|14|dimittam vero reliquias hereditatis meae et tradam eas in manu inimicorum eius eruntque in vastitate et rapina cunctis adversariis suis
2KGS|21|15|eo quod fecerint malum coram me et perseveraverint inritantes me ex die qua egressi sunt patres eorum ex Aegypto usque ad diem hanc
2KGS|21|16|insuper et sanguinem innoxium fudit Manasses multum nimis donec impleret Hierusalem usque ad os absque peccatis suis quibus peccare fecit Iudam ut faceret malum coram Domino
2KGS|21|17|reliqua autem sermonum Manasse et universa quae fecit et peccatum eius quod peccavit nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|21|18|dormivitque Manasses cum patribus suis et sepultus est in horto domus suae in horto Aza et regnavit Amon filius eius pro eo
2KGS|21|19|viginti et duo annorum erat Amon cum regnare coepisset duobusque annis regnavit in Hierusalem nomen matris eius Mesallemeth filia Arus de Iethba
2KGS|21|20|fecitque malum in conspectu Domini sicut fecerat Manasses pater eius
2KGS|21|21|et ambulavit in omni via per quam ambulaverat pater eius servivitque inmunditiis quibus servierat pater suus et adoravit eas
2KGS|21|22|et dereliquit Dominum Deum patrum suorum et non ambulavit in via Domini
2KGS|21|23|tetenderuntque ei insidias servi sui et interfecerunt regem in domo sua
2KGS|21|24|percussit autem populus terrae omnes qui coniuraverant contra regem Amon et constituerunt sibi regem Iosiam filium eius pro eo
2KGS|21|25|reliqua autem sermonum Amon quae fecit nonne haec scripta sunt in libro sermonum dierum regum Iuda
2KGS|21|26|sepelieruntque eum in sepulchro suo in horto Aza et regnavit Iosias filius eius pro eo
2KGS|22|1|octo annorum erat Iosias cum regnare coepisset et triginta uno anno regnavit in Hierusalem nomen matris eius Idida filia Phadaia de Besecath
2KGS|22|2|fecitque quod placitum erat coram Domino et ambulavit per omnes vias David patris sui non declinavit ad dextram sive ad sinistram
2KGS|22|3|anno autem octavodecimo regis Iosiae misit rex Saphan filium Aslia filii Mesullam scribam templi Domini dicens ei
2KGS|22|4|vade ad Helciam sacerdotem magnum ut confletur pecunia quae inlata est in templum Domini quam collegerunt ianitores a populo
2KGS|22|5|deturque fabris per praepositos in domo Domini qui et distribuent eam his qui operantur in templo Domini ad instauranda sarta tecta templi
2KGS|22|6|tignariis videlicet et cementariis et his qui interrupta conponunt et ut emantur ligna et lapides de lapidicinis ad instaurandum templum
2KGS|22|7|verumtamen non supputetur eis argentum quod accipiunt sed in potestate habeant et in fide
2KGS|22|8|dixit autem Helcias pontifex ad Saphan scribam librum legis repperi in domo Domini deditque Helcias volumen Saphan qui et legit illud
2KGS|22|9|venit quoque Saphan scriba ad regem et renuntiavit ei quod praeceperat et ait conflaverunt servi tui pecuniam quae repperta est in domo Domini et dederunt ut distribueretur fabris a praefectis operum templi Domini
2KGS|22|10|narravitque Saphan scriba regi dicens librum dedit mihi Helcias sacerdos quem cum legisset Saphan coram rege
2KGS|22|11|et audisset rex verba libri legis Domini scidit vestimenta sua
2KGS|22|12|et praecepit Helciae sacerdoti et Ahicham filio Saphan et Achobor filio Micha et Saphan scribae et Asaiae servo regis dicens
2KGS|22|13|ite et consulite Dominum super me et super populo et super omni Iuda de verbis voluminis istius quod inventum est magna enim ira Domini succensa est contra nos quia non audierunt patres nostri verba libri huius ut facerent omne quod scriptum est nobis
2KGS|22|14|ierunt itaque Helcias sacerdos et Ahicham et Achobor et Saphan et Asaia ad Oldam propheten uxorem Sellum filii Thecue filii Araas custodis vestium quae habitabat in Hierusalem in secunda locutique sunt ad eam
2KGS|22|15|et illa respondit eis haec dicit Dominus Deus Israhel dicite viro qui misit vos ad me
2KGS|22|16|haec dicit Dominus ecce ego adducam mala super locum hunc et super habitatores eius omnia verba legis quae legit rex Iuda
2KGS|22|17|quia dereliquerunt me et sacrificaverunt diis alienis inritantes me in cunctis operibus manuum suarum et succendetur indignatio mea in loco hoc et non extinguetur
2KGS|22|18|regi autem Iuda qui misit vos ut consuleretis Dominum sic dicetis haec dicit Dominus Deus Israhel pro eo quod audisti verba voluminis
2KGS|22|19|et perterritum est cor tuum et humiliatus es coram Domino auditis sermonibus contra locum istum et habitatores eius quo videlicet fierent in stuporem et in maledictum et scidisti vestimenta tua et flevisti coram me et ego audivi ait Dominus
2KGS|22|20|idcirco colligam te ad patres tuos et colligeris ad sepulchrum tuum in pace ut non videant oculi tui omnia mala quae inducturus sum super locum istum
2KGS|23|1|et renuntiaverunt regi quod dixerat qui misit et congregati sunt ad eum omnes senes Iuda et Hierusalem
2KGS|23|2|ascenditque rex templum Domini et omnes viri Iuda universique qui habitant in Hierusalem cum eo sacerdotes et prophetae et omnis populus a parvo usque ad magnum legitque cunctis audientibus omnia verba libri foederis qui inventus est in domo Domini
2KGS|23|3|stetitque rex super gradum et percussit foedus coram Domino ut ambularent post Dominum et custodirent praecepta eius et testimonia et caerimonias in omni corde et in tota anima et suscitarent verba foederis huius quae scripta erant in libro illo adquievitque populus pacto
2KGS|23|4|et praecepit rex Helciae pontifici et sacerdotibus secundi ordinis et ianitoribus ut proicerent de templo Domini omnia vasa quae facta fuerant Baal et in luco et universae militiae caeli et conbusit ea foris Hierusalem in convalle Cedron et tulit pulverem eorum in Bethel
2KGS|23|5|et delevit aruspices quos posuerant reges Iuda ad sacrificandum in excelsis per civitates Iuda et in circuitu Hierusalem et eos qui adolebant incensum Baal et soli et lunae et duodecim signis et omni militiae caeli
2KGS|23|6|et efferri fecit lucum de domo Domini foras Hierusalem in convalle Cedron et conbusit eum ibi et redegit in pulverem et proiecit super sepulchrum vulgi
2KGS|23|7|destruxit quoque aediculas effeminatorum quae erant in domo Domini pro quibus mulieres texebant quasi domunculas luci
2KGS|23|8|congregavitque omnes sacerdotes de civitatibus Iuda et contaminavit excelsa ubi sacrificabant sacerdotes de Gabaa usque Bersabee et destruxit aras portarum in introitu ostii Iosue principis civitatis quod erat ad sinistram portae civitatis
2KGS|23|9|verumtamen non ascendebant sacerdotes excelsorum ad altare Domini in Hierusalem sed tantum comedebant azyma in medio fratrum suorum
2KGS|23|10|contaminavit quoque Thafeth quod est in convalle filii Ennom ut nemo consecraret filium suum aut filiam per ignem Moloch
2KGS|23|11|abstulit quoque equos quos dederant reges Iudae soli in introitu templi Domini iuxta exedram Nathanmelech eunuchi qui erat in Farurim currus autem solis conbusit igni
2KGS|23|12|altaria quoque quae erant super tecta cenaculi Ahaz quae fecerant reges Iuda et altaria quae fecerat Manasses in duobus atriis templi Domini destruxit rex et cucurrit inde et dispersit cinerem eorum in torrentem Cedron
2KGS|23|13|excelsa quoque quae erant in Hierusalem ad dexteram partem montis Offensionis quae aedificaverat Salomon rex Israhel Astharoth idolo Sidoniorum et Chamos offensioni Moab et Melchom abominationi filiorum Ammon polluit rex
2KGS|23|14|et contrivit statuas et succidit lucos replevitque loca eorum ossibus mortuorum
2KGS|23|15|insuper et altare quod erat in Bethel excelsum quod fecerat Hieroboam filius Nabath qui peccare fecit Israhel et altare illud et excelsum destruxit atque conbusit et comminuit in pulverem succenditque etiam lucum
2KGS|23|16|et conversus Iosias vidit ibi sepulchra quae erant in monte misitque et tulit ossa de sepulchris et conbusit ea super altare et polluit illud iuxta verbum Domini quod locutus est vir Dei qui praedixerat verba haec
2KGS|23|17|et ait quis est titulus ille quem video responderuntque ei cives illius urbis sepulchrum est hominis Dei qui venit de Iuda et praedixit verba haec quae fecisti super altare Bethel
2KGS|23|18|et ait dimittite eum nemo commoveat ossa eius et intacta manserunt ossa illius cum ossibus prophetae qui venerat de Samaria
2KGS|23|19|insuper et omnia fana excelsorum quae erant in civitatibus Samariae quae fecerant reges Israhel ad inritandum Dominum abstulit Iosias et fecit eis secundum omnia opera quae fecerat in Bethel
2KGS|23|20|et occidit universos sacerdotes excelsorum qui erant ibi super altaria et conbusit ossa humana super ea reversusque est Hierusalem
2KGS|23|21|et praecepit omni populo dicens facite phase Domino Deo vestro secundum quod scriptum est in libro foederis huius
2KGS|23|22|nec enim factum est phase tale a diebus iudicum qui iudicaverunt Israhel et omnium dierum regum Israhel et regum Iuda
2KGS|23|23|sicut in octavodecimo anno regis Iosiae factum est phase istud Domino in Hierusalem
2KGS|23|24|sed et pythones et ariolos et figuras idolorum et inmunditias abominationesque quae fuerant in terra Iuda et in Hierusalem abstulit Iosias ut statueret verba legis quae scripta sunt in libro quem invenit Helcias sacerdos in templo Domini
2KGS|23|25|similis illi non fuit ante eum rex qui reverteretur ad Dominum in omni corde suo et in tota anima sua et in universa virtute sua iuxta omnem legem Mosi neque post eum surrexit similis illi
2KGS|23|26|verumtamen non est aversus Dominus ab ira furoris sui magni quo iratus est furor eius contra Iudam propter inritationes quibus provocaverat eum Manasses
2KGS|23|27|dixit itaque Dominus etiam Iudam auferam a facie mea sicut abstuli Israhel et proiciam civitatem hanc quam elegi Hierusalem et domum de qua dixi erit nomen meum ibi
2KGS|23|28|reliqua autem verba Iosiae et universa quae fecit nonne haec scripta sunt in libro verborum dierum regum Iuda
2KGS|23|29|in diebus eius ascendit Pharao Necho rex Aegypti contra regem Assyriorum ad flumen Eufraten et abiit Iosias rex in occursum eius et occisus est in Mageddo cum vidisset eum
2KGS|23|30|et portaverunt eum servi sui mortuum de Mageddo et pertulerunt in Hierusalem et sepelierunt eum in sepulchro suo tulitque populus terrae Ioahaz filium Iosiae et unxerunt eum et constituerunt eum regem pro patre suo
2KGS|23|31|viginti trium annorum erat Ioahaz cum regnare coepisset et tribus mensibus regnavit in Hierusalem nomen matris eius Amithal filia Hieremiae de Lobna
2KGS|23|32|et fecit malum coram Domino iuxta omnia quae fecerant patres eius
2KGS|23|33|vinxitque eum Pharao Necho in Rebla quae est in terra Emath ne regnaret in Hierusalem et inposuit multam terrae centum talentis argenti et talento auri
2KGS|23|34|regemque constituit Pharao Necho Eliachim filium Iosiae pro Iosia patre eius vertitque nomen eius Ioiachim porro Ioahaz tulit et duxit in Aegyptum
2KGS|23|35|argentum autem et aurum dedit Ioiachim Pharaoni cum indixisset terrae per singulos ut conferretur iuxta praeceptum Pharaonis et unumquemque secundum vires suas exegit tam argentum quam aurum de populo terrae ut daret Pharaoni Necho
2KGS|23|36|viginti quinque annorum erat Ioiachim cum regnare coepisset et undecim annis regnavit in Hierusalem nomen matris eius Zebida filia Phadaia de Ruma
2KGS|23|37|et fecit malum coram Domino iuxta omnia quae fecerant patres eius
2KGS|24|1|in diebus eius ascendit Nabuchodonosor rex Babylonis et factus est ei Ioiachim servus tribus annis et rursum rebellavit contra eum
2KGS|24|2|inmisitque ei Dominus latrunculos Chaldeorum et latrunculos Syriae latrunculos Moab et latrunculos filiorum Ammon et inmisit eos in Iudam ut disperderent eum iuxta verbum Domini quod locutus erat per servos suos prophetas
2KGS|24|3|factum est autem hoc per verbum Domini contra Iudam ut auferret eum coram se propter peccata Manasse universa quae fecit
2KGS|24|4|et propter sanguinem innoxium quem effudit et implevit Hierusalem cruore innocentium et ob hanc rem noluit Dominus propitiari
2KGS|24|5|reliqua autem sermonum Ioiachim et universa quae fecit nonne haec scripta sunt in libro sermonum dierum regum Iuda et dormivit Ioiachim cum patribus suis
2KGS|24|6|regnavitque Ioiachin filius eius pro eo
2KGS|24|7|et ultra non addidit rex Aegypti ut egrederetur de terra sua tulerat enim rex Babylonis a rivo Aegypti usque ad fluvium Eufraten omnia quae fuerant regis Aegypti
2KGS|24|8|decem et octo annorum erat Ioiachin cum regnare coepisset et tribus mensibus regnavit in Hierusalem nomen matris eius Naestha filia Helnathan de Hierusalem
2KGS|24|9|et fecit malum coram Domino iuxta omnia quae fecerat pater eius
2KGS|24|10|in tempore illo ascenderunt servi Nabuchodonosor regis Babylonis in Hierusalem et circumdata est urbs munitionibus
2KGS|24|11|venitque Nabuchodonosor rex Babylonis ad civitatem cum servi eius obpugnarent eam
2KGS|24|12|egressusque est Ioiachin rex Iuda ad regem Babylonis ipse et mater eius et servi eius et principes eius et eunuchi eius et suscepit eum rex Babylonis anno octavo regni sui
2KGS|24|13|et protulit inde omnes thesauros domus Domini et thesauros domus regiae et concidit universa vasa aurea quae fecerat Salomon rex Israhel in templo Domini iuxta verbum Domini
2KGS|24|14|et transtulit omnem Hierusalem et universos principes et omnes fortes exercitus decem milia in captivitatem et omnem artificem et clusorem nihilque relictum est exceptis pauperibus populi terrae
2KGS|24|15|transtulit quoque Ioiachin in Babylonem et matrem regis et uxores regis et eunuchos eius et iudices terrae duxit in captivitatem de Hierusalem in Babylonem
2KGS|24|16|et omnes viros robustos septem milia et artifices et clusores mille omnes viros fortes et bellatores duxitque eos rex Babylonis captivos in Babylonem
2KGS|24|17|et constituit Matthaniam patruum eius pro eo inposuitque nomen ei Sedeciam
2KGS|24|18|vicesimum et primum annum aetatis habebat Sedecias cum regnare coepisset et undecim annis regnavit in Hierusalem nomen matris eius erat Amithal filia Hieremiae de Lobna
2KGS|24|19|et fecit malum coram Domino iuxta omnia quae fecerat Ioiachim
2KGS|24|20|irascebatur enim Dominus contra Hierusalem et contra Iudam donec proiceret eos a facie sua recessitque Sedecias a rege Babylonis
2KGS|25|1|factum est autem anno nono regni eius mense decimo decima die mensis venit Nabuchodonosor rex Babylonis ipse et omnis exercitus eius in Hierusalem et circumdederunt eam et extruxerunt in circuitu eius munitiones
2KGS|25|2|et clausa est civitas atque vallata usque ad undecimum annum regis Sedeciae
2KGS|25|3|nona die mensis praevaluitque fames in civitate nec erat panis populo terrae
2KGS|25|4|et interrupta est civitas et omnes viri bellatores nocte fugerunt per viam portae quae est inter duplicem murum ad hortum regis porro Chaldei obsidebant in circuitu civitatem fugit itaque per viam quae ducit ad campestria solitudinis
2KGS|25|5|et persecutus est exercitus Chaldeorum regem conprehenditque eum in planitie Hiericho et omnes bellatores qui erant cum eo dispersi sunt et reliquerunt eum
2KGS|25|6|adprehensum ergo regem duxerunt ad regem Babylonis in Reblatha qui locutus est cum eo iudicium
2KGS|25|7|filios autem Sedeciae occidit coram eo et oculos eius effodit vinxitque eum catenis et adduxit in Babylonem
2KGS|25|8|mense quinto septima die mensis ipse est annus nonusdecimus regis Babylonis venit Nabuzardan princeps exercitus servus regis Babylonis Hierusalem
2KGS|25|9|et succendit domum Domini et domum regis et domos Hierusalem omnemque domum conbusit igni
2KGS|25|10|et muros Hierusalem in circuitu destruxit omnis exercitus Chaldeorum qui erat cum principe militum
2KGS|25|11|reliquam autem populi partem qui remanserat in civitate et perfugas qui transfugerant ad regem Babylonis et reliquum vulgus transtulit Nabuzardan princeps militiae
2KGS|25|12|et de pauperibus terrae reliquit vinitores et agricolas
2KGS|25|13|columnas autem aereas quae erant in templo Domini et bases et mare aereum quod erat in domo Domini confregerunt Chaldei et transtulerunt aes omnium in Babylonem
2KGS|25|14|ollas quoque aereas et trullas et tridentes et scyphos et omnia vasa aerea in quibus ministrabant tulerunt
2KGS|25|15|necnon turibula et fialas quae aurea aurea et quae argentea argentea tulit princeps militiae
2KGS|25|16|id est columnas duas mare unum et bases quas fecerat Salomon in templo Domini non erat pondus aeris omnium vasorum
2KGS|25|17|decem et octo cubitos altitudinis habebat columna una et capitellum aereum super se altitudinis trium cubitorum et reticulum et malogranata super capitellum columnae omnia aerea similem et columna secunda habebat ornatum
2KGS|25|18|tulit quoque princeps militiae Seraian sacerdotem primum et Sophoniam sacerdotem secundum et tres ianitores
2KGS|25|19|et de civitate eunuchum unum qui erat praefectus super viros bellatores et quinque viros de his qui steterant coram rege quos repperit in civitate et Sopher principem exercitus qui probabat tirones de populo terrae et sex viros e vulgo qui inventi fuerant in civitate
2KGS|25|20|quos tollens Nabuzardan princeps militum duxit ad regem Babylonis in Reblatha
2KGS|25|21|percussitque eos rex Babylonis et interfecit in Reblatha in terra Emath et translatus est Iuda de terra sua
2KGS|25|22|populo autem qui relictus erat in terra Iuda quem dimiserat Nabuchodonosor rex Babylonis praefecit Godoliam filium Ahicham filii Saphan
2KGS|25|23|quod cum audissent omnes duces militum ipsi et viri qui erant cum eis videlicet quod constituisset rex Babylonis Godoliam venerunt ad Godoliam in Maspha Ismahel filius Nathaniae et Iohanan filius Caree et Sareia filius Thenaameth Nethophathites et Iezonias filius Maachathi ipsi et socii eorum
2KGS|25|24|iuravitque eis Godolias et sociis eorum dicens nolite timere servire Chaldeis manete in terra et servite regi Babylonis et bene erit vobis
2KGS|25|25|factum est autem in mense septimo venit Ismahel filius Nathaniae filii Elisama de semine regio et decem viri cum eo percusseruntque Godoliam qui mortuus est sed et Iudaeos et Chaldeos qui erant cum eo in Maspha
2KGS|25|26|consurgens autem omnis populus a parvo usque ad magnum et principes militum venerunt in Aegyptum timentes Chaldeos
2KGS|25|27|factum est vero anno tricesimo septimo transmigrationis Ioiachin regis Iudae mense duodecimo vicesima septima die mensis sublevavit Evilmerodach rex Babylonis anno quo regnare coeperat caput Ioiachin regis Iuda de carcere
2KGS|25|28|et locutus est ei benigna et posuit thronum eius super thronum regum qui erant cum eo in Babylone
2KGS|25|29|et mutavit vestes eius quas habuerat in carcere et comedebat panem semper in conspectu eius cunctis diebus vitae suae
2KGS|25|30|annonam quoque constituit ei absque intermissione quae et dabatur ei a rege per singulos dies omnibus diebus vitae suae
