LEV|1|1|耶和華從會幕中呼叫 摩西 ，吩咐他說：
LEV|1|2|「你要吩咐 以色列 人，對他們說：你們中間若有人要獻供物給耶和華，可以從牛群羊群中獻牲畜為供物。
LEV|1|3|「他的供物若以牛為燔祭，要獻一頭沒有殘疾的公牛，獻在會幕的門口，他就可以在耶和華面前蒙悅納。
LEV|1|4|他要按手在燔祭牲的頭上，為自己贖罪，就蒙悅納。
LEV|1|5|他要在耶和華面前宰公牛犢； 亞倫 子孫作祭司的要獻上血，把血灑在會幕門口壇的周圍。
LEV|1|6|他要剝去燔祭牲的皮，把燔祭牲切成塊。
LEV|1|7|亞倫 祭司的子孫要在壇上生火，把柴擺在火上。
LEV|1|8|亞倫 子孫作祭司的要把肉塊連頭和脂肪，擺在壇上燒著火的柴上。
LEV|1|9|燔祭牲的內臟與小腿要用水洗淨，祭司要把整隻全燒在壇上，當作燔祭，是獻給耶和華為馨香的火祭。
LEV|1|10|「人的供物若以綿羊或山羊為燔祭，要獻一隻沒有殘疾的公羊。
LEV|1|11|他要在壇的北邊，在耶和華面前宰羊； 亞倫 子孫作祭司的要把血灑在壇的周圍。
LEV|1|12|他要把燔祭牲切成塊，祭司就要把肉塊連頭和脂肪，擺在壇上燒著火的柴上。
LEV|1|13|內臟與小腿要用水洗淨，祭司要把整隻獻上，全燒在壇上。這是燔祭，是獻給耶和華為馨香的火祭。
LEV|1|14|「人獻給耶和華的供物若以鳥為燔祭，就要獻斑鳩或雛鴿為他的供物。
LEV|1|15|祭司要把鳥拿到壇前，扭斷牠的頭，把鳥燒在壇上，鳥的血要流在壇的旁邊；
LEV|1|16|又要把鳥的嗉囊和裏面的髒物 除掉，丟在壇東邊倒灰的地方。
LEV|1|17|他要拿著鳥的兩個翅膀，把鳥撕開，卻不可撕斷；祭司要把牠擺在壇上燒著火的柴上焚燒。這是燔祭，是獻給耶和華為馨香的火祭。」
LEV|2|1|「若有人獻素祭為供物給耶和華，就要獻細麵為供物，把油澆在上面，加上乳香，
LEV|2|2|帶到 亞倫 子孫作祭司的那裏。祭司要從細麵中取出滿滿的一把，又取些油和所有的乳香，把這些作為紀念的燒在壇上，是獻給耶和華為馨香的火祭。
LEV|2|3|素祭所剩的要歸給 亞倫 和他的子孫；在獻給耶和華的火祭中，這是至聖的。
LEV|2|4|「若獻爐中烤的素祭為供物，要用調了油的無酵細麵餅，或抹了油的無酵薄餅。
LEV|2|5|若以鐵盤上的素祭為供物，就要用調了油的無酵細麵，
LEV|2|6|分成小塊，澆上油；這是素祭。
LEV|2|7|若以煎鍋煎的素祭為供物，就要用油與細麵做成。
LEV|2|8|要把這樣做成的素祭帶到耶和華面前，拿給祭司，祭司要帶到壇前。
LEV|2|9|祭司要從素祭中取出作為紀念的燒在壇上，是獻給耶和華為馨香的火祭。
LEV|2|10|素祭所剩的要歸給 亞倫 和他的子孫；在獻給耶和華的火祭中，這是至聖的。
LEV|2|11|「凡獻給耶和華的素祭都不可以有酵，因為你們不可把任何的酵或蜜燒了，當作火祭獻給耶和華。
LEV|2|12|你們可以把這些獻給耶和華當作初熟的供物，但是不可獻在壇上作為馨香的祭。
LEV|2|13|凡獻為素祭的供物都要用鹽調和；在素祭中，不可缺少你與上帝立約的鹽。一切的供物都要加鹽獻上。
LEV|2|14|「你若獻初熟之物給耶和華為素祭，就要獻在火中烘過的新麥穗，就是磨碎的新穀物，當作初熟之物的素祭。
LEV|2|15|你要加上油和乳香；這是素祭。
LEV|2|16|祭司要把供物中作為紀念的，就是一些磨碎的新穀物和一些油，以及所有的乳香，都焚燒，是獻給耶和華的火祭。」
LEV|3|1|「人獻平安祭為供物，若是從牛群中獻，無論是公的母的，要用沒有殘疾的，獻在耶和華面前。
LEV|3|2|他要按手在供物的頭上，在會幕的門口宰了牠。 亞倫 子孫作祭司的，要把血灑在壇的周圍。
LEV|3|3|從平安祭中，他要把火祭獻給耶和華，就是包著內臟的脂肪和內臟上所有的脂肪，
LEV|3|4|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下。
LEV|3|5|亞倫 的子孫要把這些擺在燒著火的柴上，燒在壇的燔祭上，是獻給耶和華為馨香的火祭。
LEV|3|6|「人向耶和華獻平安祭為供物，若是從羊群中獻，無論是公的母的，要用沒有殘疾的。
LEV|3|7|若他獻一隻綿羊為供物，就要把牠獻在耶和華面前。
LEV|3|8|要按手在供物的頭上，在會幕前宰了牠。 亞倫 的子孫要把血灑在壇的周圍。
LEV|3|9|從平安祭中，他要取脂肪當作火祭獻給耶和華，就是靠近脊骨處取下的整條肥尾巴，包著內臟的脂肪和內臟上所有的脂肪，
LEV|3|10|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下。
LEV|3|11|祭司要把這些燒在壇上，是獻給耶和華為食物的火祭。
LEV|3|12|「人的供物若是山羊，就要把牠獻在耶和華面前。
LEV|3|13|要按手在牠的頭上，在會幕前宰了牠。 亞倫 的子孫要把血灑在壇的周圍，
LEV|3|14|又要從供物中把火祭獻給耶和華，就是包著內臟的脂肪和內臟上所有的脂肪，
LEV|3|15|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下。
LEV|3|16|祭司要把這些燒在壇上，作為馨香火祭的食物；所有的脂肪都是耶和華的。
LEV|3|17|在你們一切的住處，脂肪和血都不可吃，這要成為你們世世代代永遠的定例。」
LEV|4|1|耶和華吩咐 摩西 說：
LEV|4|2|「你要吩咐 以色列 人說：若有人無意中犯罪，在任何事上犯了一條耶和華所吩咐的禁令，
LEV|4|3|或是受膏的祭司犯了罪，使百姓陷在罪裏，他就當為自己所犯的罪，把沒有殘疾的公牛犢獻給耶和華為贖罪祭。
LEV|4|4|他要把公牛牽到會幕的門口，在耶和華面前按手在牛的頭上，把牛宰於耶和華面前。
LEV|4|5|受膏的祭司要取些公牛的血，帶到會幕那裏。
LEV|4|6|祭司要把手指蘸在血中，在耶和華面前對著聖所的幔子彈血七次，
LEV|4|7|又要把一些血抹在會幕內，耶和華面前香壇的四個翹角上，再把公牛其餘的血全倒在會幕門口燔祭壇的底座上；
LEV|4|8|又要取出這頭贖罪祭公牛所有的脂肪，就是包著內臟的脂肪和內臟上所有的脂肪，
LEV|4|9|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下，
LEV|4|10|正如從平安祭的牛身上所取的，祭司要把這些燒在燔祭壇上。
LEV|4|11|但公牛的皮和所有的肉，以及頭、腿、內臟、糞，
LEV|4|12|就是全公牛，要搬到營外清潔的地方倒灰之處，放在柴上用火焚燒。
LEV|4|13|「 以色列 全會眾若犯了錯，在任何事上犯了一條耶和華所吩咐的禁令，而有了罪，會眾看不出這隱藏的事；
LEV|4|14|他們一知道犯了罪，就要獻一頭公牛犢為贖罪祭，牽牠到會幕前。
LEV|4|15|會眾的長老要在耶和華面前按手在公牛的頭上，把牛宰於耶和華面前。
LEV|4|16|受膏的祭司要取些公牛的血，帶到會幕那裏。
LEV|4|17|祭司要用手指蘸一些血，在耶和華面前對著幔子彈七次，
LEV|4|18|又要把一些血抹在會幕內，耶和華面前壇的四個翹角上，再把其餘的血全倒在會幕門口燔祭壇的底座上。
LEV|4|19|他要取出公牛所有的脂肪，燒在壇上。
LEV|4|20|他要處理這牛，正如處理那頭贖罪祭的公牛一樣，他要如此去做。祭司要為他們贖罪，他們就蒙赦免。
LEV|4|21|他要把牛搬到營外燒了，像燒前一頭公牛一樣；這是會眾的贖罪祭。
LEV|4|22|「官長若犯罪，在任何事上無意中犯了一條耶和華－他的上帝所吩咐的禁令，而有了罪，
LEV|4|23|他一知道自己犯了罪，就要牽一隻沒有殘疾的公山羊為供物。
LEV|4|24|他要按手在羊的頭上，在耶和華面前宰燔祭牲的地方把牠宰了；這是贖罪祭。
LEV|4|25|祭司要用手指蘸一些贖罪祭牲的血，抹在燔祭壇的四個翹角上，再把其餘的血倒在燔祭壇的底座上。
LEV|4|26|祭牲所有的脂肪都要燒在壇上，正如平安祭的脂肪一樣。祭司要為他的罪贖了他，他就蒙赦免。
LEV|4|27|「這地的百姓若有人無意中犯罪，在任何事上犯了一條耶和華所吩咐的禁令，而有了罪，
LEV|4|28|他一知道自己犯了罪，就要為所犯的罪牽一隻沒有殘疾的母山羊為供物。
LEV|4|29|他要按手在贖罪祭牲的頭上，在燔祭牲的地方把牠宰了。
LEV|4|30|祭司要用手指蘸一些祭牲的血，抹在燔祭壇的四個翹角上，再把其餘的血全倒在壇的底座上；
LEV|4|31|又要把祭牲所有的脂肪都取下，正如取平安祭牲的脂肪一樣。祭司要把脂肪燒在壇上，在耶和華面前作為馨香的祭。祭司要為他贖罪，他就蒙赦免。
LEV|4|32|「人若牽一隻綿羊為贖罪祭作供物，就要牽一隻沒有殘疾的母羊。
LEV|4|33|他要按手在贖罪祭牲的頭上，在宰燔祭牲的地方宰了牠，作為贖罪祭。
LEV|4|34|祭司要用手指蘸一些贖罪祭牲的血，抹在燔祭壇的四個翹角上，再把其餘的血全倒在壇的底座上；
LEV|4|35|又要把祭牲所有的脂肪都取下，正如取平安祭的羊的脂肪一樣。祭司要按獻給耶和華火祭的條例，把脂肪燒在壇上。祭司要為他所犯的罪贖了他，他就蒙赦免。」
LEV|5|1|「若有人犯了罪，就是聽見了誓言，他本來可以作證，卻不把所看見、所知道的說出來，必須擔當他的罪孽。
LEV|5|2|若有人摸了任何不潔之物，無論是野獸的不潔屍體，家畜的不潔屍體，或是群聚動物的不潔屍體，他雖不察覺，也是不潔淨，就有罪了。
LEV|5|3|或是他摸了人的不潔之物，就是任何使人成為不潔的不潔之物，他雖不察覺，但一知道，就有罪了。
LEV|5|4|若有人隨口發誓，或出於惡意，或出於善意，這人無論在甚麼事上隨意發誓，雖不察覺，但一知道，就在這其中的一件事上有罪了。
LEV|5|5|當他在這其中的一件事上有罪的時候，就要承認所犯的罪，
LEV|5|6|並要為所犯的罪，把他的贖愆祭牲，就是羊群中的一隻母綿羊或母山羊，獻給耶和華為贖罪祭，祭司要為他的罪贖了他。
LEV|5|7|「若他的力量不夠獻一隻綿羊，就要為所犯的罪，把兩隻斑鳩或是兩隻雛鴿獻給耶和華為贖愆祭：一隻作贖罪祭，一隻作燔祭。
LEV|5|8|他要把這些帶到祭司那裏，祭司就先把贖罪祭獻上，從鳥的頸項上扭斷牠的頭，但不把鳥撕斷。
LEV|5|9|祭司要把一些贖罪祭牲的血彈在祭壇的邊上，其餘的血要倒在壇的底座上；這是贖罪祭。
LEV|5|10|他要依照條例獻第二隻鳥為燔祭。祭司要為他所犯的罪贖了他，他就蒙赦免。
LEV|5|11|「他的力量若不夠獻兩隻斑鳩或兩隻雛鴿，就要為所犯的罪把供物，就是十分之一伊法細麵，獻上為贖罪祭；不可加上油，也不可加上乳香，因為這是贖罪祭。
LEV|5|12|他要把細麵帶到祭司那裏，祭司要取出滿滿的一把，作為紀念，按照獻火祭給耶和華的條例把它燒在壇上；這是贖罪祭。
LEV|5|13|至於他在這幾件事中所犯的任何罪，祭司要為他贖了，他就蒙赦免。剩下的都歸給祭司，和素祭一樣。」
LEV|5|14|耶和華吩咐 摩西 說：
LEV|5|15|「若有人在耶和華的聖物上無意中犯了罪，有了過犯，就要獻羊群中一隻沒有殘疾的公綿羊給耶和華為贖愆祭，或依聖所的舍客勒所估定的銀子，作為贖愆祭。
LEV|5|16|他要為在聖物上的疏忽賠償，另外加五分之一，把這些都交給祭司。祭司要用贖愆祭的公綿羊為他贖罪，他就蒙赦免。
LEV|5|17|「若有人犯罪，在任何事上犯了一條耶和華所吩咐的禁令，他雖不察覺，仍算有罪，必須擔當自己的罪孽。
LEV|5|18|他要牽羊群中一隻沒有殘疾的公綿羊，或照你所估定的價值，給祭司作贖愆祭。祭司要為他贖他因不知道而無意中所犯的罪，他就蒙赦免。
LEV|5|19|這是贖愆祭；因他確實得罪了耶和華。」
LEV|6|1|耶和華吩咐 摩西 說：
LEV|6|2|「若有人犯罪，得罪了耶和華，就是在鄰舍寄託他的東西或抵押品上行詭詐，或搶奪，或欺壓鄰舍，
LEV|6|3|或是撿了失物行了詭詐，起了假誓，在人所做的任何事上犯了罪；
LEV|6|4|他既犯了罪，有了過犯，就要歸還他所搶奪的，或是因欺壓所得的，或是別人寄託他的，或是他所撿到的失物，
LEV|6|5|或是起假誓得來的任何東西，就要全數歸還，另外再加五分之一。在查出他有罪的日子，就要立刻賠還給原主。
LEV|6|6|他要獻羊群中一隻沒有殘疾的公綿羊，給耶和華為贖愆祭，或照你所估定的價值，給祭司 作贖愆祭。
LEV|6|7|祭司要在耶和華面前為他贖罪；他無論做了甚麼事，以致有了罪，都必蒙赦免。」
LEV|6|8|耶和華吩咐 摩西 說：
LEV|6|9|「你要吩咐 亞倫 和他的子孫說，燔祭的條例是這樣：燔祭要放在壇的底盤上，從晚上到天亮，壇上的火要不斷地燒著。
LEV|6|10|祭司要穿上細麻布衣服，又要把細麻布褲子穿在身上，把在壇上燒剩的燔祭灰收起來，放在壇的旁邊。
LEV|6|11|然後，他要脫去這衣服，穿上別的衣服，把灰拿到營外潔淨之處。
LEV|6|12|壇上的火要不斷地燒著，不可熄滅。每日早晨，祭司要在壇上燒柴，把燔祭擺在壇上，並燒平安祭牲的脂肪。
LEV|6|13|壇上的火要不斷地燒著，不可熄滅。」
LEV|6|14|「素祭的條例是這樣： 亞倫 的子孫要在壇前把這祭獻在耶和華面前。
LEV|6|15|祭司要從素祭中的細麵取出一把，再取些油和素祭上所有的乳香，把這些作為紀念的燒在壇上，是獻給耶和華為馨香的祭。
LEV|6|16|亞倫 和他子孫要吃素祭剩下的；要在聖處吃這無酵餅，在會幕的院子裏吃。
LEV|6|17|烤餅不可加酵。這是從獻給我的火祭中歸給他們的一份；如贖罪祭和贖愆祭一樣，這份是至聖的。
LEV|6|18|亞倫 子孫中的男丁都要吃，因為這是你們世世代代從獻給耶和華的火祭中，他們永遠應得的份。凡摸這些祭物的都要成為聖。」
LEV|6|19|耶和華吩咐 摩西 說：
LEV|6|20|「這是 亞倫 受膏的日子，他和他的子孫所要獻給耶和華的供物：十分之一伊法細麵，如他們經常獻的素祭，早晨一半，晚上一半。
LEV|6|21|要在鐵盤上用油調和，調勻後，就拿去烤。素祭烤熟了要分成小塊，作為獻給耶和華馨香的祭。
LEV|6|22|亞倫 子孫中接續他受膏為祭司的，要把這素祭獻上，全燒給耶和華。這是永遠的定例。
LEV|6|23|祭司一切的素祭要全部燒了，不可以吃。」
LEV|6|24|耶和華吩咐 摩西 說：
LEV|6|25|「你要吩咐 亞倫 和他的子孫說，贖罪祭的條例是這樣：要在耶和華面前宰燔祭牲的地方宰贖罪祭牲；這是至聖的。
LEV|6|26|獻贖罪祭的祭司要吃這祭物；要在聖處，就是在會幕的院子裏吃。
LEV|6|27|凡摸這祭肉的都要成為聖；這祭牲的血若濺在衣服上，你要在聖處洗淨那濺到血的衣服 。
LEV|6|28|煮這祭物的瓦器要打碎；若祭物是在銅器裏煮，要把這銅器擦淨，用水沖洗。
LEV|6|29|祭司中所有的男丁都可以吃；這是至聖的。
LEV|6|30|若將任何贖罪祭的血帶進會幕，為要在聖所贖罪，那肉就不可吃，要用火焚燒。」
LEV|7|1|「贖愆祭的條例是這樣：這祭是至聖的。
LEV|7|2|人在哪裏宰燔祭牲，也要在哪裏宰贖愆祭牲；其血，祭司要灑在壇的周圍。
LEV|7|3|祭司要獻上牠所有的脂肪，把肥尾巴和包著內臟的脂肪，
LEV|7|4|兩個腎和腎上的脂肪，即靠近腎兩旁的脂肪，以及肝上的網油，連同腎一起取下。
LEV|7|5|祭司要把這些燒在壇上，獻給耶和華為火祭，作為贖愆祭。
LEV|7|6|祭司中所有的男丁都可以吃這祭物，要在聖處吃；這是至聖的。
LEV|7|7|贖罪祭怎樣，贖愆祭也是怎樣，都有一樣的條例，用贖愆祭贖罪的祭司要得這祭物。
LEV|7|8|獻燔祭的祭司，無論為誰獻，所獻燔祭牲的皮要歸給那祭司，那是他的。
LEV|7|9|任何素祭，無論是在爐中烤的，用煎鍋或鐵盤做成的，都要歸給獻祭的祭司。
LEV|7|10|任何素祭，無論是用油調和的，是乾的，都要歸 亞倫 的子孫，大家均分。」
LEV|7|11|「獻給耶和華平安祭的條例是這樣：
LEV|7|12|若有人為感謝獻祭，就要把用油調和的無酵餅、抹了油的無酵薄餅，和用油調勻細麵做成的餅，與感謝祭一同獻上。
LEV|7|13|要用有酵的餅，和那為感謝而獻的平安祭，與供物一同獻上。
LEV|7|14|他要從每一種供物中拿一個餅，獻給耶和華為舉祭，是要歸給那灑平安祭牲血的祭司。
LEV|7|15|為感謝而獻的平安祭的肉，要在獻祭當天吃，一點也不可留到早晨。
LEV|7|16|若所獻的是還願祭或甘心祭，要在獻祭當天吃，剩下的，第二天也可以吃。
LEV|7|17|第三天，所剩下的祭肉要用火焚燒。
LEV|7|18|第三天若吃平安祭的肉，必不蒙悅納，所獻的也不算為祭；這祭物是不潔淨的，凡吃這祭物的，必擔當自己的罪孽。
LEV|7|19|「沾了不潔淨之物的肉就不可吃，要用火焚燒。至於其他的肉，凡潔淨的人都可以吃這肉；
LEV|7|20|但不潔淨的人若吃了獻給耶和華平安祭的肉，這人必從民中剪除。
LEV|7|21|若有人摸了不潔之物，無論是人體的不潔淨，或是不潔的牲畜，或是不潔的可憎之物 ，再吃了獻給耶和華平安祭的肉，這人必從民中剪除。」
LEV|7|22|耶和華吩咐 摩西 說：
LEV|7|23|「你要吩咐 以色列 人說：牛、綿羊、山羊的脂肪，你們都不可吃。
LEV|7|24|自然死去的或被野獸撕裂的，那脂肪可以作別的用途，你們卻萬不可吃。
LEV|7|25|任何人吃了獻給耶和華作火祭祭牲的脂肪，這人必從民中剪除。
LEV|7|26|在你們一切的住處，無論是鳥或獸的血，你們都不可吃。
LEV|7|27|無論誰吃了血，這人必從民中剪除。」
LEV|7|28|耶和華吩咐 摩西 說：
LEV|7|29|「你要吩咐 以色列 人說：獻平安祭給耶和華的，要從他的平安祭中取些供物來獻給耶和華。
LEV|7|30|他要親手把獻給耶和華的火祭帶來，要把脂肪和胸帶來，把胸在耶和華面前搖一搖，作為搖祭。
LEV|7|31|祭司要把脂肪燒在壇上，但胸要歸給 亞倫 和他的子孫。
LEV|7|32|你們要從平安祭牲中把右腿作為舉祭，送給祭司。
LEV|7|33|亞倫 子孫中獻平安祭牲的血和脂肪的，要得這右腿，作為他當得的份。
LEV|7|34|因為我從 以色列 人的平安祭中，把這搖祭的胸和這舉祭的腿給 亞倫 祭司和他子孫，作為他們在 以色列 人中永遠當得的份。」
LEV|7|35|這是從耶和華的火祭中取出，作為 亞倫 和他子孫受膏的份，就是 摩西 叫他們前來，給耶和華供祭司職分的那一天開始的。
LEV|7|36|這是在 摩西 膏他們的日子，耶和華吩咐給他們的，作為他們在 以色列 人中世世代代永遠當得的份。
LEV|7|37|這就是燔祭、素祭、贖罪祭、贖愆祭、聖職禮和平安祭的條例，
LEV|7|38|都是耶和華在 西奈山 上吩咐 摩西 的，也是他在 西奈 曠野吩咐 以色列 人獻供物給耶和華的日子所說的。
LEV|8|1|耶和華吩咐 摩西 說：
LEV|8|2|「你領 亞倫 和他兒子前來，並將聖衣、膏油，與贖罪祭的一頭公牛、兩隻公綿羊、一筐無酵餅都一同帶來；
LEV|8|3|又要召集全會眾到會幕的門口。」
LEV|8|4|摩西 就遵照耶和華的吩咐做了，於是會眾聚集在會幕的門口。
LEV|8|5|摩西 對會眾說：「這是耶和華所吩咐當做的事。」
LEV|8|6|摩西 領了 亞倫 和他兒子前來，用水洗他們。
LEV|8|7|他給 亞倫 穿上內袍，束上腰帶，套上外袍，加上以弗得，再束上精緻的帶子，把以弗得繫在他身上。
LEV|8|8|他又給 亞倫 戴上胸袋，把烏陵和土明放在胸袋內。
LEV|8|9|他把禮冠戴在 亞倫 的頭上，禮冠前面安上金牌，成為聖冕，是照耶和華所吩咐 摩西 的。
LEV|8|10|摩西 用膏油抹帳幕和其中所有的，使它們成為聖。
LEV|8|11|他又用膏油在祭壇上彈了七次，抹了壇和壇的一切器皿，以及洗濯盆和盆座，使它們成為聖。
LEV|8|12|他把膏油倒在 亞倫 的頭上膏他，使他成為聖。
LEV|8|13|摩西 帶了 亞倫 的兒子來，給他們穿上內袍，束上腰帶，裹上頭巾，是照耶和華所吩咐 摩西 的。
LEV|8|14|他把贖罪祭的公牛牽來， 亞倫 和他兒子按手在贖罪祭公牛的頭上，
LEV|8|15|就宰了公牛。 摩西 取了血，用指頭抹在祭壇周圍的四個翹角上，使壇潔淨，再把其餘的血倒在壇的底座上，使壇成為聖，為壇贖罪。
LEV|8|16|摩西 把內臟所有的脂肪和肝上的網油，以及兩個腎與腎上的脂肪取出，都燒在壇上。
LEV|8|17|至於公牛，連皮帶肉和糞，他都用火燒在營外，是照耶和華所吩咐 摩西 的。
LEV|8|18|他把燔祭的公綿羊牽來， 亞倫 和他兒子按手在羊的頭上，
LEV|8|19|就宰了公羊。 摩西 把血灑在祭壇的周圍，
LEV|8|20|把羊切成塊，把頭和肉塊，以及脂肪拿去燒，
LEV|8|21|他用水洗了內臟和腿之後，就把全羊燒在壇上，作為馨香的燔祭，是獻給耶和華的火祭，都是照耶和華所吩咐 摩西 的。
LEV|8|22|他又牽來第二隻公綿羊，就是聖職禮的羊， 亞倫 和他兒子按手在羊的頭上，
LEV|8|23|就宰了羊。 摩西 把一些血抹在 亞倫 的右耳垂上，右手的大拇指上和右腳的大腳趾上。
LEV|8|24|他領了 亞倫 的兒子來，把一些血抹在他們的右耳垂上，右手的大拇指上和右腳的大腳趾上。 摩西 把其餘的血灑在壇的周圍。
LEV|8|25|他把脂肪，肥尾巴、內臟所有的脂肪、肝上的網油、兩個腎、腎上的脂肪，和右腿取下，
LEV|8|26|再從耶和華面前那裝無酵餅的籃子中取一個無酵餅、一個油餅和一個薄餅，把這些放在脂肪和右腿上。
LEV|8|27|他把這一切放在 亞倫 和他兒子的手上，在耶和華面前搖一搖，作為搖祭。
LEV|8|28|摩西 從他們的手上把這些祭物拿來，放在壇的燔祭上燒，這就是聖職禮中獻給耶和華馨香的火祭。
LEV|8|29|摩西 拿羊的胸，在耶和華面前搖一搖，作為搖祭，這是聖職禮的羊歸給 摩西 的一份，是照耶和華所吩咐 摩西 的。
LEV|8|30|摩西 取些膏油和壇上的血，彈在 亞倫 和他的衣服上，以及他兒子和他們的衣服上，使 亞倫 和他的衣服，他兒子和他們的衣服都成為聖。
LEV|8|31|摩西 對 亞倫 和他兒子說：「你們要在會幕的門口把肉煮了，在那裏吃這肉和聖職禮中籃子裏的餅，按我所吩咐的說：『這是 亞倫 和他兒子當吃的。』
LEV|8|32|剩下的肉和餅，你們要用火焚燒。
LEV|8|33|這七天，你們不可走出會幕的門口，直等到你們聖職禮的日子滿了，因為授予你們聖職需要七天 。
LEV|8|34|今天所做的，都是耶和華吩咐要做的，好為你們贖罪。
LEV|8|35|這七天，你們要晝夜留在會幕門內，遵守耶和華所吩咐的，免得你們死亡，因為所吩咐我的就是這樣。」
LEV|8|36|於是， 亞倫 和他的兒子就做了耶和華藉著 摩西 所吩咐的一切事。
LEV|9|1|到了第八天， 摩西 召 亞倫 和他兒子，以及 以色列 的眾長老來，
LEV|9|2|對 亞倫 說：「你當取一頭公牛犢作贖罪祭，一隻公綿羊作燔祭，都要沒有殘疾的，獻在耶和華面前。
LEV|9|3|你要對 以色列 人說：『你們當取一隻公山羊作贖罪祭，再取一頭牛犢和一隻小綿羊，都要一歲沒有殘疾的，作燔祭；
LEV|9|4|又當取一頭公牛，一隻公綿羊作平安祭，宰殺獻在耶和華面前，再加上調油的素祭。因為今天耶和華要向你們顯現。』」
LEV|9|5|於是，他們把 摩西 所吩咐的帶到會幕前；全會眾都近前來，站在耶和華面前。
LEV|9|6|摩西 說：「這是耶和華吩咐你們當做的事，耶和華的榮光要向你們顯現。」
LEV|9|7|摩西 對 亞倫 說：「你靠近祭壇前，獻你的贖罪祭和燔祭，為自己與百姓贖罪，再獻上百姓的供物，為他們贖罪，都是照耶和華所吩咐的。」
LEV|9|8|於是， 亞倫 靠近壇前，宰了那頭為自己贖罪的牛犢。
LEV|9|9|亞倫 的兒子把血遞給他，他就把指頭蘸在血中，抹在壇的四個翹角上，再把其餘的血倒在壇的底座上。
LEV|9|10|他把贖罪祭的脂肪和腎，以及肝上的網油，燒在壇上，是照耶和華所吩咐 摩西 的。
LEV|9|11|他用火將肉和皮燒在營外。
LEV|9|12|亞倫 把燔祭牲宰了，他兒子把血遞給他，他就把血灑在壇的周圍。
LEV|9|13|他們又把燔祭一塊一塊地，連頭遞給他，他就燒在壇上。
LEV|9|14|他又洗了內臟和腿，放在壇的燔祭上燒。
LEV|9|15|然後，他奉上百姓的供物。他牽來給百姓作贖罪祭的公山羊，把牠宰了，獻為贖罪祭，和先前的一樣。
LEV|9|16|他也奉上燔祭，按照條例獻上。
LEV|9|17|除了早晨的燔祭以外，他又獻上素祭，用手取了滿滿的一把，燒在壇上。
LEV|9|18|亞倫 宰了那給百姓作平安祭的公牛和公綿羊，他兒子把血遞給他，他就把血灑在壇的周圍；
LEV|9|19|他們把公牛和公綿羊的脂肪、肥尾巴，包著內臟的脂肪，腎和肝上的網油，都遞給他。
LEV|9|20|他們把脂肪放在祭牲的胸上，他就把脂肪燒在壇上。
LEV|9|21|亞倫 把祭牲的胸和右腿在耶和華面前搖一搖，作為搖祭，是照 摩西 所吩咐的。
LEV|9|22|亞倫 向百姓舉手，為他們祝福。他獻了贖罪祭、燔祭、平安祭就下來了。
LEV|9|23|摩西 和 亞倫 進了會幕。他們出來，為百姓祝福；耶和華的榮光向全體百姓顯現。
LEV|9|24|有火從耶和華面前出來，焚燒了壇上的燔祭和脂肪；全體百姓一看見，就都歡呼，臉伏於地。
LEV|10|1|亞倫 的兒子 拿答 和 亞比戶 各拿著自己的香爐，把火放在爐裏，加上香，在耶和華面前獻上凡火，是耶和華沒有吩咐他們的。
LEV|10|2|有火從耶和華面前出來，把他們吞滅，他們就死在耶和華面前。
LEV|10|3|於是， 摩西 對 亞倫 說：「這就是耶和華所吩咐的，說：『我在那親近我的人中要顯為聖；在全體百姓面前，我要得著榮耀。』」 亞倫 就默默不言。
LEV|10|4|摩西 召 亞倫 的叔父 烏薛 的兒子 米沙利 和 以利撒反 前來，對他們說：「過來，把你們的親屬從聖所前抬到營外。」
LEV|10|5|於是，二人過來把屍體連袍子一起抬到營外，是照 摩西 所吩咐的。
LEV|10|6|摩西 對 亞倫 和他兒子 以利亞撒 和 以他瑪 說：「不可蓬頭散髮，也不可撕裂衣服，免得你們死亡，免得耶和華向全會眾發怒。但你們的弟兄 以色列 全家卻要為耶和華發出的火哀哭。
LEV|10|7|你們也不可出會幕的門口，免得你們死亡，因為耶和華的膏油在你們身上。」他們就遵照 摩西 的話去做了。
LEV|10|8|耶和華吩咐 亞倫 說：
LEV|10|9|「你和你兒子進會幕的時候，清酒烈酒都不可喝，免得你們死亡，這要作你們世世代代永遠的定例。
LEV|10|10|你們必須分辨聖的俗的，潔淨的和不潔淨的，
LEV|10|11|也要將耶和華藉 摩西 吩咐 以色列 人的一切律例教導他們。」
LEV|10|12|摩西 對 亞倫 和他剩下的兒子 以利亞撒 和 以他瑪 說：「獻給耶和華的火祭中所剩下的素祭，你們要拿來，在祭壇旁吃這無酵餅，因為它是至聖的。
LEV|10|13|你們要在聖處吃，因為在獻給耶和華的火祭中，這是你和你兒子當得的份；所吩咐我的就是這樣。
LEV|10|14|這搖祭的胸和這舉祭的腿，你要在潔淨的地方和你的兒女一同吃，因為這些是從 以色列 人的平安祭中歸給你，作為你和你兒子當得的份。
LEV|10|15|他們要把舉祭的腿、搖祭的胸和火祭的脂肪一同帶來，在耶和華面前搖一搖，作為搖祭。這些要歸給你和你兒子，作永遠當得的份，都是照耶和華所吩咐的。」
LEV|10|16|那時， 摩西 急切地尋找那隻贖罪祭的公山羊，看哪，牠已經燒掉了。他向 亞倫 剩下的兒子 以利亞撒 和 以他瑪 發怒，說：
LEV|10|17|「你們為何沒有在聖所吃這贖罪祭呢？它是至聖的，是耶和華給你們的，為了除掉會眾的罪孽，在耶和華面前為他們贖罪。
LEV|10|18|看哪，這祭牲的血沒有拿到聖所裏去！你們應當照我所吩咐的，在聖所裏吃這祭肉。」
LEV|10|19|亞倫 對 摩西 說：「看哪，他們今天在耶和華面前獻上贖罪祭和燔祭，但是我卻遭遇這樣的災難。我若今天吃這贖罪祭，耶和華豈能看為美呢？」
LEV|10|20|摩西 聽了，就看為美。
LEV|11|1|耶和華吩咐 摩西 和 亞倫 ，對他們說：
LEV|11|2|「你們要吩咐 以色列 人說，地上一切的走獸中可吃的動物是這些：
LEV|11|3|凡蹄分兩瓣，分趾蹄而又反芻食物的走獸，你們都可以吃。
LEV|11|4|但那反芻或分蹄之中不可吃的是：駱駝，反芻卻不分蹄，對你們是不潔淨的；
LEV|11|5|石獾，反芻卻不分蹄，對你們是不潔淨的；
LEV|11|6|兔子，反芻卻不分蹄，對你們是不潔淨的；
LEV|11|7|豬，蹄分兩瓣，分趾蹄卻不反芻，對你們是不潔淨的。
LEV|11|8|這些獸的肉，你們不可吃；牠們的屍體，你們也不可摸，對你們都是不潔淨的。
LEV|11|9|「水中可吃的是這些：凡在水裏，無論是海或河，有鰭有鱗的，都可以吃。
LEV|11|10|凡在海裏、河裏和水裏滋生的動物，就是在水裏所有的動物，無鰭無鱗的，對你們是可憎的。
LEV|11|11|牠們對你們都是可憎的。你們不可吃牠們的肉；牠們的屍體，也當以為可憎。
LEV|11|12|凡在水裏無鰭無鱗的，對你們是可憎的。
LEV|11|13|「飛鳥中你們當以為可憎，不可吃且可憎的是：鵰、狗頭鵰、紅頭鵰，
LEV|11|14|鷂鷹、小鷹的類群，
LEV|11|15|所有烏鴉的類群，
LEV|11|16|鴕鳥、夜鷹、魚鷹、鷹的類群，
LEV|11|17|鴞鳥、鸕鶿、貓頭鷹，
LEV|11|18|角鴟、鵜鶘、禿鵰，
LEV|11|19|鸛、鷺鷥的類群，戴鵀與蝙蝠。
LEV|11|20|「凡有翅膀卻用四足爬行的群聚動物，對你們是可憎的。
LEV|11|21|只是有翅膀卻用四足爬行的群聚動物中，足上有腿在地上跳的，你們還可以吃；
LEV|11|22|其中你們可以吃的有蝗蟲的類群，螞蚱的類群，蟋蟀的類群和蚱蜢的類群。
LEV|11|23|其餘有翅膀有四足的群聚動物，對你們都是可憎的。
LEV|11|24|「這些都能使你們不潔淨。凡摸牠們屍體的，必不潔淨到晚上。
LEV|11|25|任何人搬動了牠們的屍體，要把衣服洗淨，必不潔淨到晚上。
LEV|11|26|凡蹄分兩瓣卻不分趾或不反芻食物的走獸，對你們是不潔淨的；誰摸了牠們就不潔淨。
LEV|11|27|凡用腳掌行走，四足行走的動物，對你們是不潔淨的；凡摸牠們屍體的，必不潔淨到晚上。
LEV|11|28|誰搬動了牠們的屍體，要把衣服洗淨，必不潔淨到晚上。這些對你們是不潔淨的。
LEV|11|29|「在地上成群的群聚動物中，對你們不潔淨的是這些：鼬鼠、鼫鼠、蜥蜴的類群，
LEV|11|30|壁虎、龍子、守宮、蛇醫、蝘蜓。
LEV|11|31|這些群聚動物對你們都是不潔淨的。在牠們死後，凡摸了牠們屍體的，必不潔淨到晚上。
LEV|11|32|其中死了的，若掉在任何東西上，這東西就不潔淨，無論是木器、衣服、皮革、麻袋，或是任何工作需用的器皿，都要泡在水中，必不潔淨到晚上，然後才是潔淨的。
LEV|11|33|若有一點掉在瓦器裏，裏面的任何東西就不潔淨了； 你們要把這瓦器打破。
LEV|11|34|其中一切可吃的食物，沾到那水的就不潔淨；器皿裏可喝的東西，也必不潔淨。
LEV|11|35|牠們的屍體，只要有一點掉在任何物件上，那物件就不潔淨。無論是烤爐或爐灶，都要打碎；它們不潔淨，而且對你們也不潔淨。
LEV|11|36|但是水泉或池子，就是聚水的地方，仍是潔淨的；凡摸這些屍體的才不潔淨。
LEV|11|37|若牠們的屍體有一點掉在要播的種子上，種子仍是潔淨的；
LEV|11|38|若水已經澆在種子上，牠們的屍體有一點掉在上面，這種子對你們就是不潔淨的了。
LEV|11|39|「你們可吃的走獸中若有死了的，誰摸了牠的屍體，就必不潔淨到晚上。
LEV|11|40|人若吃了那已死的走獸，要把衣服洗淨，必不潔淨到晚上。人若搬動了那已死的牲畜，要把衣服洗淨，必不潔淨到晚上。
LEV|11|41|「凡在地上成群的群聚動物都是可憎的，都不可吃。
LEV|11|42|凡用肚子爬行或用四腳爬行，或是用多足的，地上一切群聚的動物，你們都不可吃，因為是可憎的。
LEV|11|43|你們不可因任何群聚的動物使自己成為可憎的，也不可因牠們成為不潔淨，染了污穢。
LEV|11|44|我是耶和華－你們的上帝。你們要使自己分別為聖，要成為聖，因為我是神聖的。你們不可因地上爬行的群聚動物使自己不潔淨。
LEV|11|45|我是把你們從 埃及 地領出來的耶和華，要作你們的上帝。你們要成為聖，因為我是神聖的。」
LEV|11|46|這是牲畜、飛鳥、水中一切游動的生物和地上一切爬行的動物的條例，
LEV|11|47|為要使你們能分辨潔淨的和不潔淨的，可吃的和不可吃的動物。
LEV|12|1|耶和華吩咐 摩西 說：
LEV|12|2|「你要吩咐 以色列 人說：婦人若懷孕生男孩，就不潔淨七天，像在月經污穢的期間不潔淨一樣。
LEV|12|3|第八天，要給嬰孩行割禮。
LEV|12|4|婦人產後流血的潔淨，要家居三十三天。她潔淨的日子未滿，不可摸聖物，也不可進入聖所。
LEV|12|5|她若生女孩，就不潔淨兩個七天，像經期中一樣。她產後流血的潔淨，要家居六十六天。
LEV|12|6|「潔淨的日子滿了，無論生兒子或女兒，她要把一隻一歲的羔羊作燔祭，一隻雛鴿或一隻斑鳩作贖罪祭，帶到會幕的門口交給祭司。
LEV|12|7|祭司要把這祭物獻在耶和華面前，為她贖罪。這樣，她就從流血中得潔淨了。這是為生男或生女之婦人的條例。
LEV|12|8|婦人的能力若不足，無法獻一隻羔羊，她就要取兩隻斑鳩或兩隻雛鴿，一隻為燔祭，一隻為贖罪祭。祭司要為她贖罪，她就潔淨了。」
LEV|13|1|耶和華吩咐 摩西 和 亞倫 說：
LEV|13|2|「人身上的皮膚若腫脹，或發疹，或有斑點，可能成為痲瘋 的災病，就要把他帶到 亞倫 祭司或 亞倫 的一個作祭司的子孫那裏。
LEV|13|3|祭司要檢查他身上皮膚的患處，若患處的毛已經變白，災病的現象深入身上皮膚內，這就是痲瘋的災病。祭司檢查後，要宣佈他為不潔淨。
LEV|13|4|若這人身上的皮膚有白斑，看起來並沒有深入皮膚內，其上的毛也沒有變白，祭司就要將這病人隔離七天。
LEV|13|5|第七天，祭司要檢查他，看哪，若災病在祭司眼前止住了，沒有在皮膚上擴散，要將他再隔離七天。
LEV|13|6|到了第七天，祭司要再檢查他。看哪，若災病減輕，沒有在皮膚上擴散，祭司就要宣佈他為潔淨，因為他患的不過是疹子。那人要洗自己的衣服，就潔淨了。
LEV|13|7|他給祭司檢查宣佈為潔淨後，疹子若在皮膚上大大擴散，他就要再給祭司檢查。
LEV|13|8|祭司要檢查，看哪，疹子若在皮膚上擴散了，祭司就要宣佈他為不潔淨，是痲瘋病。
LEV|13|9|「人若得了痲瘋的災病，就要把他帶到祭司那裏。
LEV|13|10|祭司要檢查，看哪，若皮膚有白色腫塊，使毛變白，腫塊裏有嫩的新長的肉，
LEV|13|11|這就是他身上皮膚慢性的痲瘋病。祭司要宣佈他為不潔淨，不必將他隔離，因為他已是不潔淨了。
LEV|13|12|若痲瘋在皮膚四處擴散，長滿在患災病之人的皮膚上，據祭司察看，從頭到腳無處不有，
LEV|13|13|祭司就要檢查，看哪，若這病人全身已長滿了痲瘋，就要宣佈他為潔淨；他全身都變白了，他是潔淨的。
LEV|13|14|但他身上一旦出現新長的肉，就不潔淨了。
LEV|13|15|祭司一見新長的肉，就要宣佈他為不潔淨。新長的肉是不潔淨的，這就是痲瘋病。
LEV|13|16|新長的肉若變白了，他就要到祭司那裏。
LEV|13|17|祭司要檢查，看哪，患處若變白了，祭司就要宣佈那患災病的人為潔淨，他就潔淨了。
LEV|13|18|「人身上的皮膚 若長了瘡，卻已經好了，
LEV|13|19|在長瘡之處又發腫變白，或是出現白中帶紅的斑點，就要給祭司檢查。
LEV|13|20|祭司要檢查，看哪，若災病的現象已深入皮膚內，其上的毛也變白了，祭司就要宣佈他為不潔淨，有痲瘋的災病生在瘡中。
LEV|13|21|祭司若檢查，看哪，其上沒有白毛，也沒有深入皮膚內，而且災病減輕，祭司就要將他隔離七天。
LEV|13|22|若在皮膚上大大擴散，祭司就要宣佈他為不潔淨，這是災病。
LEV|13|23|斑點若留在原處，沒有擴散，這就是瘡的疤痕，祭司就要宣佈他為潔淨。
LEV|13|24|「人身上的皮膚若被火燒傷，傷口新長的肉有了斑點，無論是白中帶紅，或是全白，
LEV|13|25|祭司就要檢查，看哪，斑點上的毛若變白了，現象又深入皮膚內，這就是痲瘋長在燒傷處；祭司就要宣佈他為不潔淨，是痲瘋的災病。
LEV|13|26|若祭司檢查，看哪，斑點上沒有白毛，也沒有深入皮膚內，而且災病減輕，祭司就要將他隔離七天。
LEV|13|27|第七天，祭司要檢查他。斑點若在皮膚上大大擴散，祭司就要宣佈他為不潔淨，是患了痲瘋的災病。
LEV|13|28|斑點若留在原處，沒有在皮膚上擴散，並減輕了，它只是燒傷的腫塊，祭司要宣佈他為潔淨，這不過是燒傷後的疤痕。
LEV|13|29|「無論男女，若在頭上或下巴有災病，
LEV|13|30|祭司就要檢查這災病，看哪，若災病的現象深入皮膚內，其上有黃色的細毛，祭司就要宣佈他為不潔淨，這是疥瘡，是頭上或下巴的痲瘋病。
LEV|13|31|祭司要檢查這疥瘡的災病，看哪，現象若未深入皮膚內，其上也沒有黑毛，祭司就要將長疥瘡的人隔離七天。
LEV|13|32|第七天，祭司要檢查這災病，看哪，若疥瘡沒有擴散，其上沒有黃色的毛，疥瘡的現象也沒有深入皮膚內，
LEV|13|33|那人就要剃去鬚髮，但不可剃長疥瘡之處。祭司要將那長疥瘡的人，再隔離七天。
LEV|13|34|第七天，祭司要檢查疥瘡，看哪，疥瘡若沒有在皮膚上擴散，現象也未深入在皮膚內，祭司就要宣佈他為潔淨；那人要洗自己的衣服，就潔淨了。
LEV|13|35|但他被宣佈為潔淨後，疥瘡若在皮膚上大大擴散，
LEV|13|36|祭司就要檢查他。看哪，疥瘡若在皮膚上擴散，祭司就不必找黃色的毛，這人是不潔淨了。
LEV|13|37|若疥瘡在祭司眼前止住了，其上長了黑毛，疥瘡就已痊癒了，那人是潔淨的，祭司要宣佈他為潔淨。
LEV|13|38|「無論男女，身上的皮膚若有斑點，是白色的斑點，
LEV|13|39|祭司就要檢查，看哪，若皮膚的斑點是暗白色的，這是皮膚長了斑；那人是潔淨的。
LEV|13|40|「人的頭髮若掉了，變成禿頭，他是潔淨的。
LEV|13|41|他頭頂的前面若掉了頭髮，以致頂門光禿，他是潔淨的。
LEV|13|42|頭禿處或頂門禿處，若有白中帶紅的災病，這就是痲瘋長在他的頭禿處或頂門禿處。
LEV|13|43|祭司要檢查他，看哪，若頭禿處或頂門禿處的災病腫塊白中帶紅，像身上皮膚痲瘋病的現象一樣，
LEV|13|44|那人就是患了痲瘋病，是不潔淨的。祭司要宣佈他為不潔淨；他的災病是生在頭上。
LEV|13|45|「患有痲瘋災病的人，他的衣服要撕裂，也要蓬頭散髮，遮住上唇，喊著說：『不潔淨！不潔淨！』
LEV|13|46|災病還在他身上的時候，他就是不潔淨的；既然不潔淨，他就要獨居，住在營外。」
LEV|13|47|「衣服若發霉 了，無論是羊毛衣服、麻布衣服，
LEV|13|48|無論是經線、緯線，是麻布的、羊毛的，是皮革，或是任何皮製的物件；
LEV|13|49|若是衣服、皮革、經線、緯線，或是任何皮製的物件呈現綠色或紅色，這就是發霉，必須給祭司檢查。
LEV|13|50|祭司要檢查這霉，把發霉的物件隔離七天。
LEV|13|51|第七天，他要檢查這霉。若霉在衣服上，無論是經線、緯線，或任何用途的皮製物件上擴散，這是侵蝕性的霉，是不潔淨的。
LEV|13|52|發霉的衣服，無論在經線、緯線，羊毛的、麻布的，或是任何皮製物件，都要把它燒掉；因為這是侵蝕性的霉，必須用火焚燒。
LEV|13|53|祭司檢查，看哪，霉若在衣服上，無論是經線、緯線，或在任何的皮製物件上沒有擴散，
LEV|13|54|祭司就要吩咐人把發霉的物件洗了，再隔離七天。
LEV|13|55|洗過之後，祭司要檢查，看哪，若那霉在他眼前沒有變色，霉雖沒有擴散，也是不潔淨的。這是侵蝕性的災病，無論是在正面或反面，都要用火焚燒那物件。
LEV|13|56|祭司若檢查，看哪，那霉在洗過之後已經褪色，他就要從衣服，皮革，或經線、緯線，把發霉的部分撕去。
LEV|13|57|若霉再出現在衣服上，無論是經線、緯線、或在任何皮製物件上，這就是舊霉復發，必須用火將那發霉的物件焚燒。
LEV|13|58|洗過的衣服，或是經線，緯線，或是任何皮製的物件，若霉已經消失了，仍要再洗，這衣服就潔淨了。」
LEV|13|59|這就是衣服發霉的條例。無論是羊毛衣服，麻布衣服，或是經線、緯線，或任何皮製的物件，都按照這條例宣佈為潔淨或不潔淨。
LEV|14|1|耶和華吩咐 摩西 說：
LEV|14|2|「這是患痲瘋病的人得潔淨時的條例：要帶他到祭司那裏，
LEV|14|3|祭司要出到營外，檢查那患痲瘋病的人，看哪，他的痲瘋災病已經痊癒了，
LEV|14|4|祭司就要吩咐人為那求潔淨的人帶兩隻潔淨的活鳥和香柏木、朱紅色紗，以及牛膝草來。
LEV|14|5|祭司要吩咐用瓦器盛清水，把第一隻鳥宰在上面。
LEV|14|6|至於那隻活鳥，祭司要把牠和香柏木、朱紅色紗，以及牛膝草，一同蘸在宰於清水上的鳥血中。
LEV|14|7|他要向那從痲瘋病中得潔淨的人身上彈血七次，宣佈他為潔淨，然後把那活鳥在野地裏放走。
LEV|14|8|求潔淨的人要洗衣服，剃去所有的毛髮，用水洗澡，他就潔淨了。然後，他可以進營，不過仍要在自己的帳棚外居住七天。
LEV|14|9|到了第七天，他要剃所有的毛髮，頭髮、鬍鬚、眼睛的眉毛，他全身的毛都剃了；然後，他要洗衣服，用水洗身，才潔淨了。
LEV|14|10|「第八天，他要取兩隻沒有殘疾的小公羊和一隻沒有殘疾、一歲的小母羊，以及作為素祭的十分之三伊法調了油的細麵和一羅革的油。
LEV|14|11|宣佈潔淨的祭司要將那求潔淨的人，連同這些東西，安置在耶和華面前，會幕的門口。
LEV|14|12|祭司要取一隻小公羊獻為贖愆祭，又取一羅革的油，把它們在耶和華面前搖一搖，作為搖祭；
LEV|14|13|再把小公羊宰於聖處，就是宰贖罪祭牲和燔祭牲的地方。贖愆祭要歸給祭司，與贖罪祭一樣，是至聖的。
LEV|14|14|祭司要取一些贖愆祭牲的血，抹在求潔淨的人的右耳垂上、右手的大拇指上和右腳的大腳趾上。
LEV|14|15|祭司要從那一羅革的油中，取一些倒在自己的左手掌裏，
LEV|14|16|祭司要用右手指蘸在他左手掌的油裏，在耶和華面前用手指彈七次。
LEV|14|17|祭司要把手掌裏剩下的油抹在那求潔淨的人的右耳垂上、右手的大拇指上和右腳的大腳趾上，在贖愆祭牲之血抹過的上面。
LEV|14|18|祭司手掌裏剩下的油要抹在那求潔淨的人的頭上，祭司就在耶和華面前為他贖罪。
LEV|14|19|祭司要獻贖罪祭，為那從不潔淨中得潔淨的人贖罪，然後要宰燔祭牲，
LEV|14|20|祭司要把燔祭和素祭獻在壇上，祭司要為他贖罪，他就潔淨了。
LEV|14|21|「他若貧窮，手頭財力不及，就要取一隻小公羊作贖愆祭，作搖祭為他贖罪。他也要把作為素祭的十分之一伊法調了油的細麵，和一羅革的油，一同取來。
LEV|14|22|他又要照手頭財力所及，取兩隻斑鳩或兩隻雛鴿，一隻作贖罪祭，一隻作燔祭。
LEV|14|23|第八天，為了使自己潔淨，他要把這些祭物帶到耶和華面前，在會幕的門口交給祭司。
LEV|14|24|祭司要把贖愆祭的羔羊和那一羅革的油一同在耶和華面前搖一搖，作為搖祭。
LEV|14|25|祭司要宰贖愆祭的羔羊，取一些贖愆祭牲的血，抹在那求潔淨的人的右耳垂上、右手的大拇指上和右腳的大腳趾上。
LEV|14|26|祭司要把一些油倒在自己的左手掌裏，
LEV|14|27|祭司要用右手指，把他左手掌裏的油在耶和華面前彈七次。
LEV|14|28|祭司要把手掌裏的油抹一些在那求潔淨的人的右耳垂上、右手的大拇指上和右腳的大腳趾上，在贖愆祭牲之血抹過之處的上面。
LEV|14|29|祭司手掌裏剩下的油要抹在那求潔淨的人的頭上，在耶和華面前為他贖罪。
LEV|14|30|那人又要照他手頭財力所及，獻上斑鳩中的一隻或雛鴿中的一隻，
LEV|14|31|照他手頭財力所及，一隻為贖罪祭，一隻為燔祭，與素祭一同獻上。祭司就在耶和華面前為他贖罪。
LEV|14|32|這是為患痲瘋災病，手頭財力不及而求潔淨的人所定的條例。」
LEV|14|33|耶和華吩咐 摩西 和 亞倫 說：
LEV|14|34|「你們到了我所賜給你們為業的 迦南 地，我若使你們所得為業之地的房屋發霉 ，
LEV|14|35|屋主就要去告訴祭司說：『據我看，房屋似乎發霉了。』
LEV|14|36|祭司進去檢查這霉之前，要吩咐把屋內的東西全部搬走，免得屋子裏所有的東西成為不潔淨。然後，祭司要進去檢查房屋。
LEV|14|37|他要檢查這霉，看哪，若屋子牆上的霉有發綠或發紅凹入的斑紋，其現象深入牆內，
LEV|14|38|祭司就要出到屋子的門外，把屋子封鎖七天。
LEV|14|39|第七天，祭司要再去檢查，看哪，霉若在屋子的牆上擴散，
LEV|14|40|祭司要吩咐把發霉的石頭挖出來，扔在城外不潔淨之處。
LEV|14|41|他也要叫人刮屋內的四圍，把刮出來的灰泥倒在城外不潔淨之處。
LEV|14|42|他們要用別的石頭取代挖出來的石頭，用別的灰泥塗抹屋子。
LEV|14|43|「他挖出石頭，刮了屋子，塗抹以後，霉若又在屋子裏出現，
LEV|14|44|祭司就要進去檢查，看哪，霉若在屋子裏擴散，那就是有侵蝕性的霉在屋子裏，是不潔淨的。
LEV|14|45|他要拆毀屋子，把石頭、木料和所有的灰泥都搬到城外不潔淨之處。
LEV|14|46|屋子封鎖的任何時候，進去的人必不潔淨到晚上。
LEV|14|47|在屋子裏躺臥的人必須把衣服洗淨，在屋子裏吃飯的人也必須把衣服洗淨。
LEV|14|48|「屋子塗抹了之後，祭司若進去檢查，看哪，霉沒有在屋內擴散，就要宣佈這房屋為潔淨，因為霉已經消除了。
LEV|14|49|他要為潔淨房屋取兩隻鳥和香柏木、朱紅色紗，以及牛膝草，
LEV|14|50|用瓦器盛清水，把一隻鳥宰在上面。
LEV|14|51|他要把香柏木、牛膝草、朱紅色紗和那一隻活鳥，都蘸在被宰的鳥血和清水中，用來彈屋子七次。
LEV|14|52|他要用鳥血、清水、活鳥、香柏木、牛膝草和朱紅色紗潔淨那房屋。
LEV|14|53|他要把活鳥在城外野地裏放走。他要為房屋贖罪，房屋就潔淨了。」
LEV|14|54|這條例是為痲瘋災病和疥瘡，
LEV|14|55|衣服和房屋發霉，
LEV|14|56|以及皮膚腫脹、發疹、有斑點等，
LEV|14|57|用以分辨何時潔淨，何時不潔淨。這是痲瘋病的條例。
LEV|15|1|耶和華吩咐 摩西 和 亞倫 說：
LEV|15|2|「你們要吩咐 以色列 人，對他們說：人若身體 患了漏症，他因這症就不潔淨了。
LEV|15|3|這就是他因漏症而有的不潔淨：無論是身體流出液體，或身體已經止住不再有液體，他都是不潔淨的。
LEV|15|4|那患漏症的人所躺的床都不潔淨，所坐的任何東西也不潔淨。
LEV|15|5|凡摸他床的人，要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|6|人坐了漏症患者坐過的東西，他要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|7|人摸了漏症患者，他要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|8|若漏症患者吐唾沫在潔淨的人身上，這人要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|9|漏症患者所騎的任何鞍子也不潔淨。
LEV|15|10|凡摸了他坐過的任何東西，必不潔淨到晚上；拿了這些東西的，要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|11|漏症患者若沒有用水沖洗他的手，無論摸了誰，誰就要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|12|漏症患者所摸的瓦器必要打破；他所摸的一切木器必要用水沖洗。
LEV|15|13|「漏症患者的漏症痊癒了，就要為潔淨自己計算七天，也要洗衣服，用清水洗身，就潔淨了。
LEV|15|14|第八天，他要帶兩隻斑鳩或兩隻雛鴿，來到耶和華面前，在會幕門口把鳥交給祭司。
LEV|15|15|祭司要獻上一隻為贖罪祭，一隻為燔祭。祭司要因這人所患的漏症，在耶和華面前為他贖罪。
LEV|15|16|「人若遺精，他要用水洗全身，必不潔淨到晚上。
LEV|15|17|無論是衣服或皮革，若沾染了精液，要用水洗淨，必不潔淨到晚上。
LEV|15|18|女人，若有男人與她同寢，沾染了精液，二人要用水洗澡，必不潔淨到晚上。」
LEV|15|19|「女人月經期間，有血從體內流出，她必不潔淨七天；凡摸她的，必不潔淨到晚上。
LEV|15|20|在不潔淨期間，女人所躺的東西都不潔淨，所坐的任何東西也不潔淨。
LEV|15|21|凡摸她床的，要洗衣服，用水洗澡，必不潔淨到晚上；
LEV|15|22|凡摸她坐過的東西的，要洗衣服，用水洗澡，必不潔淨到晚上；
LEV|15|23|不論是床，或她坐過的東西，人摸了，必不潔淨到晚上。
LEV|15|24|男人若和這女人同寢，沾了她的不潔淨，就不潔淨七天，所躺的床也都不潔淨。
LEV|15|25|「女人若在經期之外仍然流血多日，或是經期過長，她在流血的一切日子都不潔淨，和她在經期的日子不潔淨一樣。
LEV|15|26|在流血的日子，她所躺的床、所坐的任何東西都不潔淨，和在月經期間不潔淨一樣。
LEV|15|27|凡摸這些東西的，就不潔淨；他要洗衣服，用水洗澡，必不潔淨到晚上。
LEV|15|28|這女人的血漏若痊癒了，就要計算七天，然後才潔淨。
LEV|15|29|第八天，她要取兩隻斑鳩或兩隻雛鴿，帶到會幕門口祭司那裏。
LEV|15|30|祭司要獻一隻為贖罪祭，一隻為燔祭。祭司要因這女人血漏的不潔淨，在耶和華面前為她贖罪。
LEV|15|31|「你們要使 以色列 人與他們的不潔淨隔離，免得他們玷污我在他們中間的帳幕，因自己的不潔淨死亡。」
LEV|15|32|這條例是為漏症患者或遺精而不潔淨者，
LEV|15|33|女人經期的不潔，男女患漏症，以及男人與不潔淨女人同寢而立的。
LEV|16|1|亞倫 的兩個兒子靠近耶和華面前，死了。他們死後，耶和華吩咐 摩西 ；
LEV|16|2|耶和華對 摩西 說：「你要吩咐你哥哥 亞倫 ，不可隨時進入聖所的幔子內、到櫃蓋 前，免得他死亡，因為我在櫃蓋上的雲中顯現。
LEV|16|3|亞倫 進聖所要帶這些：一頭公牛犢為贖罪祭，一隻公綿羊為燔祭。
LEV|16|4|他要穿上細麻布聖內袍，把細麻布褲子穿在身上，腰束細麻布帶子，頭戴細麻布禮冠；這些都是聖服。他要用水洗身，然後穿上聖服。
LEV|16|5|他要從 以色列 會眾中取兩隻公山羊為贖罪祭，一隻公綿羊為燔祭。
LEV|16|6|「亞倫要把他自己贖罪祭的公牛獻上，為自己和家人贖罪；
LEV|16|7|也要把兩隻公山羊牽到耶和華面前，安置在會幕的門口。
LEV|16|8|亞倫 要為那兩隻山羊抽籤，一籤歸給耶和華，一籤歸給 阿撒瀉勒 。
LEV|16|9|亞倫 要把那抽中歸給耶和華的山羊牽來獻為贖罪祭，
LEV|16|10|至於抽中歸給 阿撒瀉勒 的山羊，卻要活著安放在耶和華面前，用以贖罪，然後送到曠野去，歸給 阿撒瀉勒 。
LEV|16|11|「 亞倫 要把他自己贖罪祭的公牛獻上，為自己和家人贖罪，他要宰作自己贖罪祭的公牛。
LEV|16|12|他要從耶和華面前的壇上取盛滿火炭的香爐，再拿一捧搗細的香料，把這些都帶入幔子內。
LEV|16|13|在耶和華面前，他要把香放在火上，使香的煙雲遮著法櫃上的蓋子，免得他死亡。
LEV|16|14|他要取一些公牛的血，用手指彈在櫃蓋的前面，就是東面，又在櫃蓋的前面用手指彈血七次。
LEV|16|15|「他要宰那隻為百姓作贖罪祭的公山羊，把羊的血帶入幔子內，把血彈在櫃蓋的上面和前面，好像彈公牛的血一樣。
LEV|16|16|因 以色列 人的不潔淨和過犯，就是他們一切的罪，他要為聖所贖罪；因會幕在他們不潔淨之中，他也要為會幕照樣做。
LEV|16|17|他進聖所贖罪的時候，會幕裏都不准有人，直等到他為自己和家人，以及 以色列 全會眾贖了罪出來。
LEV|16|18|他出來後，要到耶和華面前的祭壇那裏，為壇贖罪。他要取一些公牛的血和公山羊的血，抹在壇周圍的四個翹角上。
LEV|16|19|他也要用手指把血彈在壇上七次，使壇從 以色列 人的不潔淨中得以潔淨，成為聖。」
LEV|16|20|「 亞倫 為聖所和會幕，以及祭壇贖罪後，就要把那隻活的公山羊牽來。
LEV|16|21|他的雙手要按在活的山羊的頭上，承認 以色列 人所有的罪孽過犯，就是他們一切的罪，把這些罪都歸在羊的頭上，再指派一個人把牠送到曠野去。
LEV|16|22|這羊要擔當他們一切的罪孽，帶到無人之地；那人要把羊送到曠野去。
LEV|16|23|「 亞倫 要進入會幕，把他進聖所時所穿的細麻布衣服脫下，放在那裏，
LEV|16|24|又要在聖處用水洗身，穿上衣服出來，把自己的燔祭和百姓的燔祭獻上，為自己和百姓贖罪。
LEV|16|25|贖罪祭牲的脂肪要燒在壇上。
LEV|16|26|那放走山羊歸給 阿撒瀉勒 的人要洗衣服，用水洗身，然後才可以回到營裏。
LEV|16|27|作贖罪祭的公牛和作贖罪祭的公山羊的血被帶入聖所贖罪之後，就要把這牛羊搬到營外，皮、肉、糞都用火焚燒。
LEV|16|28|焚燒的人要洗衣服，用水洗身，然後才可以回到營裏。」
LEV|16|29|「這是你們永遠的定例：每年七月初十，你們要刻苦己心；無論是本地人，是寄居在你們中間的外人，任何工都不可做。
LEV|16|30|因為這日要為你們贖罪，潔淨你們，使你們脫離一切的罪，在耶和華面前得以潔淨。
LEV|16|31|這日你們要守完全安息的安息日，刻苦己心；這是永遠的定例。
LEV|16|32|那受膏接續他父親擔任聖職的祭司要贖罪，穿上細麻布衣服，就是聖衣，
LEV|16|33|為至聖所和會幕贖罪，為祭壇贖罪，並要為祭司和會眾的全體百姓贖罪。
LEV|16|34|這要作你們永遠的定例：因 以色列 人一切的罪，要一年一次為他們贖罪。」於是， 亞倫 照耶和華所吩咐 摩西 的做了 。
LEV|17|1|耶和華吩咐 摩西 說：
LEV|17|2|「你要吩咐 亞倫 和他兒子，以及 以色列 眾人，對他們說，耶和華所吩咐的話是這樣：
LEV|17|3|凡 以色列 家中的人宰公牛，或小綿羊，或山羊，無論是在營內或營外，
LEV|17|4|若不把牲畜牽到會幕門口耶和華的帳幕前，獻給耶和華為供物，所流的血必歸到那人身上。他既使血流出，就要從百姓中剪除。
LEV|17|5|這是為要使 以色列 人把他們在野地裏所宰的祭牲帶來，帶到耶和華前，會幕門口祭司那裏，宰殺這些祭牲，把牠們獻給耶和華為平安祭。
LEV|17|6|祭司要在會幕門口，把血灑在耶和華的祭壇上，把脂肪焚燒，獻給耶和華為馨香的祭。
LEV|17|7|他們不可再宰殺祭牲獻給他們行淫所隨從的山羊鬼魔。這要作他們世世代代永遠的定例。
LEV|17|8|「你要對他們說：凡 以色列 家中的任何人，或寄居在他們中間的外人獻燔祭或祭物，
LEV|17|9|若不帶到會幕門口獻給耶和華，那人必從百姓中剪除。
LEV|17|10|「凡 以色列 家中的任何人，或寄居在他們中間的外人，吃任何的血，我必向那吃血的人變臉，把他從百姓中剪除。
LEV|17|11|因為動物的生命是在血中。我把這血賜給你們，可以在祭壇上為你們的生命贖罪；因為血就是生命，能夠贖罪。
LEV|17|12|因此，我對 以色列 人說：你們都不可吃血；寄居在你們中間的外人也不可吃血。
LEV|17|13|凡 以色列 人，或寄居在他們中間的外人，獵取了可吃的飛禽走獸，必須把牠的血放出來，用土掩蓋。
LEV|17|14|「因一切動物的生命，牠的血就是牠的生命。所以我對 以色列 人說：無論甚麼動物的血，你們都不可吃，因為一切動物的生命就是牠的血。凡吃血的必被剪除。
LEV|17|15|無論是本地人，是寄居的，若吃了自然死去或被野獸撕裂的動物，要洗衣服，用水洗澡，必不潔淨到晚上，晚上就潔淨了。
LEV|17|16|但他若不洗衣服，也不洗身，就要擔當自己的罪孽。」
LEV|18|1|耶和華吩咐 摩西 說：
LEV|18|2|「你要吩咐 以色列 人，對他們說：我是耶和華－你們的上帝。
LEV|18|3|你們不可做你們從前住 埃及 地的人所做的，也不可做我要領你們去的 迦南 地的人所做的。你們不可照他們的習俗行。
LEV|18|4|你們要遵行我的典章，謹守我的律例，按此而行。我是耶和華－你們的上帝。
LEV|18|5|你們要謹守我的律例典章；遵行的人就必因此得生。我是耶和華。
LEV|18|6|「任何人都不可親近骨肉之親，露其下體。我是耶和華。
LEV|18|7|你父親的下體，就是你母親的下體，你不可露；她是你的母親，不可露她的下體。
LEV|18|8|不可露你繼母的下體，就是你父親的下體。
LEV|18|9|你姊妹的下體，或是同父異母的，或是同母異父的，無論生在家或生在外的，都不可露她們的下體。
LEV|18|10|不可露你孫女或外孫女的下體，因為她們的下體就是你自己的下體。
LEV|18|11|你繼母為你父親所生的女兒是你的姊妹，不可露她的下體。
LEV|18|12|不可露你姑母的下體；她是你父親的骨肉之親。
LEV|18|13|不可露你姨母的下體；她是你母親的骨肉之親。
LEV|18|14|不可露你叔伯的下體，不可親近他的妻子；她是你的叔母、伯母。
LEV|18|15|不可露你媳婦的下體，她是你兒子的妻，不可露她的下體。
LEV|18|16|不可露你兄弟妻子的下體，這是你兄弟的下體。
LEV|18|17|不可露婦人的下體，又露她女兒的下體，也不可娶她的孫女或外孫女，露她們的下體；她們是骨肉之親 。這是邪惡的事。
LEV|18|18|你妻子還活著的時候，不可另娶她的姊妹與她作對，露她姊妹的下體。
LEV|18|19|「不可親近經期中不潔淨的女人，露她的下體。
LEV|18|20|不可跟鄰舍的妻交合，因她玷污自己。
LEV|18|21|不可使你兒女經火獻給 摩洛 ，也不可褻瀆你上帝的名。我是耶和華。
LEV|18|22|不可跟男人同寢，像跟女人同寢；這是可憎惡的事。
LEV|18|23|不可跟獸交合，因牠玷污自己。女人也不可站在獸前，與牠交合；這是逆性的事。
LEV|18|24|「在這一切的事上，你們都不可玷污自己，因為我在你們面前所逐出的列國，在這一切的事上玷污了自己。
LEV|18|25|連地也玷污了，我懲罰那地的罪孽，地就吐出它的居民來。
LEV|18|26|但你們要遵守我的律例典章。這一切可憎惡的事，無論是本地人或寄居在你們中間的外人，都不可以做。
LEV|18|27|在你們之前居住那地的人做了這一切可憎惡的事，地就玷污了。
LEV|18|28|不要讓地因你們玷污了它而把你們吐出來，像吐出在你們之前的國一樣。
LEV|18|29|無論是誰，若做了這其中一件可憎惡的事，必從百姓中剪除。
LEV|18|30|你們要遵守我的吩咐，免得你們隨從那些可憎的習俗，就是在你們之前的人所做的，玷污了自己。我是耶和華－你們的上帝。」
LEV|19|1|耶和華吩咐 摩西 說：
LEV|19|2|「你要吩咐 以色列 全會眾，對他們說：你們要成為聖，因為我耶和華－你們的上帝是神聖的。
LEV|19|3|你們各人都當孝敬父母，也要守我的安息日。我是耶和華－你們的上帝。
LEV|19|4|你們不可轉向虛無的神明，也不可為自己鑄造神像。我是耶和華－你們的上帝。
LEV|19|5|「你們宰殺祭牲獻平安祭給耶和華的時候，要獻得使你們可蒙悅納。
LEV|19|6|這祭物要在獻的當天或第二天吃；若有剩到第三天的，就要用火焚燒。
LEV|19|7|第三天若再吃，這祭物是不潔淨的，必不蒙悅納。
LEV|19|8|吃的人必擔當自己的罪孽，因為他褻瀆了耶和華的聖物，這人必從百姓中剪除。
LEV|19|9|「你們在自己的地收割莊稼時，不可割盡田的角落，也不可拾取莊稼所掉落的。
LEV|19|10|不可摘盡葡萄園的葡萄，也不可拾取葡萄園中掉落的葡萄，要把它們留給窮人和寄居的。我是耶和華－你們的上帝。
LEV|19|11|「你們不可偷盜，不可欺騙，也不可彼此說謊。
LEV|19|12|不可指著我的名起假誓，褻瀆你上帝的名。我是耶和華。
LEV|19|13|「不可欺壓你的鄰舍，也不可偷盜。雇工的工錢不可在你那裏過夜，留到早晨。
LEV|19|14|不可咒罵聾子，也不可將絆腳石放在盲人面前。你要敬畏你的上帝。我是耶和華。
LEV|19|15|「你們審判的時候，不可不公正；不可偏護貧窮人，也不可看重有權勢人的臉，總要公平審判你的鄰舍。
LEV|19|16|不可在百姓中到處搬弄是非，不可陷害鄰舍的性命 。我是耶和華。
LEV|19|17|「不可心裏恨你的弟兄；要指摘你的鄰舍，免得因他承擔罪過。
LEV|19|18|不可報仇，也不可埋怨你本國的子民。你要愛鄰如己。我是耶和華。
LEV|19|19|「你們要遵守我的律例。不可使你的牲畜與異類交配；不可在你的田地播下兩樣的種子；也不可穿兩種原料做成的衣服。
LEV|19|20|「若有人與女子同寢交合，而她是婢女，許配了丈夫，尚未被贖或得自由，就要受到懲罰，卻不可把他們處死，因為婢女還沒有得自由。
LEV|19|21|男的要把贖愆祭，就是一隻公綿羊牽到耶和華面前，會幕的門口。
LEV|19|22|祭司要用贖愆祭的羊在耶和華面前為他所犯的罪贖罪，他所犯的罪就必蒙赦免。
LEV|19|23|「你們到了 迦南 地，栽種各樣的果樹，就要把所結的果子當作不潔淨的 ；三年之內，你們要把它視為不潔淨，是不可吃的。
LEV|19|24|但第四年所結的果子全是聖的，用以讚美耶和華 。
LEV|19|25|第五年，你們就可以吃樹上的果子，使樹給你們結出更多的果子。我是耶和華－你們的上帝。
LEV|19|26|「你們不可吃帶血的食物。不可占卜，也不可觀星象。
LEV|19|27|頭的周圍 不可剃，鬍鬚的周圍不可損壞。
LEV|19|28|不可為死人割劃自己的身體，也不可在身上刺花紋。我是耶和華。
LEV|19|29|「不可侮辱你的女兒，使她淪為娼妓，免得這地行淫亂，地就充滿了邪惡。
LEV|19|30|你們要謹守我的安息日，敬畏我的聖所。我是耶和華。
LEV|19|31|「不可轉向招魂的，也不可求問行巫術的，免得被他們玷污。我是耶和華－你們的上帝。
LEV|19|32|「在白髮的人面前，你要站起來，要尊敬老人；要敬畏你的上帝，我是耶和華。
LEV|19|33|「若有外人寄居在你們的地上和你同住，不可欺負他。
LEV|19|34|寄居在你們那裏的外人，你們要看他如本地人，並要愛他如己，因為你們在 埃及 地也作過寄居的。我是耶和華－你們的上帝。
LEV|19|35|「你們審判的時候，不可用不公正的度量衡。
LEV|19|36|你們要用公正的天平、公正的法碼、公正的伊法和公正的欣。我是耶和華－你們的上帝，曾把你們從 埃及 地領出來。
LEV|19|37|你們要謹守我一切的律例典章，遵行它們。我是耶和華。」
LEV|20|1|耶和華吩咐 摩西 說：
LEV|20|2|「你要對 以色列 人說：凡 以色列 人，或是寄居在 以色列 的外人，把自己兒女獻給 摩洛 的，必被處死；本地的百姓要用石頭打死他。
LEV|20|3|我也要向那人變臉，把他從百姓中剪除，因為他把兒女獻給 摩洛 ，玷污了我的聖所，褻瀆了我的聖名。
LEV|20|4|那人把兒女獻給 摩洛 ，本地的百姓若假裝沒看見，不把他處死，
LEV|20|5|我就要向這人和他的家人變臉，把他和所有跟隨他與 摩洛 行淫的人都從百姓中剪除。
LEV|20|6|「人若轉向招魂的和行巫術的，隨從他們行淫，我就要向這人變臉，把他從百姓中剪除。
LEV|20|7|你們要使自己分別為聖，要成為聖，因為我是耶和華－你們的上帝。
LEV|20|8|你們要謹守我的律例，遵行它們；我是使你們分別為聖的耶和華。
LEV|20|9|凡咒罵父母的，必被處死；他咒罵了父母，他的血要歸在他身上。
LEV|20|10|「凡與有夫之婦行姦淫，就是與鄰舍的妻子行姦淫的，姦夫淫婦必被處死。
LEV|20|11|人若與繼母同寢，就是露了父親的下體，二人必被處死，血要歸在他們身上。
LEV|20|12|人若與媳婦同寢，二人必被處死；他們行了亂倫的事，血要歸在他們身上。
LEV|20|13|男人若跟男人同寢，像跟女人同寢，他們二人行了可憎惡的事，必被處死，血要歸在他們身上。
LEV|20|14|人若娶妻，又娶妻子的母親，這是邪惡的事；要把這三人用火焚燒，在你們中間除去這邪惡。
LEV|20|15|人若與獸交合，必被處死；你們也要殺死那獸。
LEV|20|16|女人若與獸親近，與牠交合，你要把那女人和獸殺死；他們必被處死，血要歸在他們身上。
LEV|20|17|「人若娶自己的姊妹，或是同父異母的，或是同母異父的，彼此見了下體，這是可恥的事；他們必在自己百姓眼前被剪除。他露了姊妹的下體，必擔當自己的罪孽。
LEV|20|18|若有人跟經期中的婦人同寢，露了她的下體，暴露婦人的血源，婦人也露了自己的血源，二人必從百姓中剪除。
LEV|20|19|不可露姨母或姑母的下體，因為這是露了骨肉之親的下體，他們必擔當自己的罪孽。
LEV|20|20|人若與叔伯之妻同寢，就露了他叔伯的下體，他們必擔當自己的罪，必沒有子女而死。
LEV|20|21|人若娶了自己兄弟的妻子，就露了他兄弟的下體，這是不潔淨的事，他們必沒有子女。
LEV|20|22|「你們要謹守我一切的律例典章，遵行它們，免得我領你們去住的那地把你們吐出來。
LEV|20|23|我在你們面前所逐出的國民，你們不可隨從他們的風俗。因為他們行了這一切的事，所以我厭惡他們。
LEV|20|24|但我對你們說過，你們要承受他們的土地；我要把這流奶與蜜之地賜給你們，作為你們的產業。我是耶和華－你們的上帝，是把你們從萬民中分別出來的。
LEV|20|25|你們要分辨潔淨和不潔淨的飛禽走獸；不可因我定為不潔淨的飛禽走獸，或爬行在土地上的任何生物，使自己成為可憎惡的。
LEV|20|26|你們要歸我為聖，因為－我耶和華是神聖的；我把你們從萬民中分別出來，作我的子民。
LEV|20|27|「無論男女，是招魂的或行巫術的，他們必被處死。人要用石頭打死他們，血要歸在他們身上。」
LEV|21|1|耶和華對 摩西 說：「你要告訴 亞倫 子孫作祭司的，對他們說：祭司不可為自己百姓中的死人玷污自己，
LEV|21|2|除非是他的骨肉之親，他的父母、兒女、兄弟、
LEV|21|3|或未出嫁還是處女的姊妹，因她是至親，才可以玷污自己。
LEV|21|4|祭司既然在自己百姓中為首，就不可從俗玷污自己 。
LEV|21|5|「不可使頭光禿，不可剃除鬍鬚的邊緣，也不可割劃自己的身體。
LEV|21|6|他們要歸上帝為聖，不可褻瀆他們上帝的名，因為耶和華的火祭，就是上帝的食物，是他們獻的，所以他們要成為聖。
LEV|21|7|「祭司不可娶妓女，或被玷污的女人為妻，也不可娶被休的婦人為妻，因為他是歸上帝為聖的。
LEV|21|8|你要使祭司分別為聖，因為他獻你上帝的食物。你要以他為聖，因為我是使你們分別為聖 的耶和華，是神聖的。
LEV|21|9|「祭司的女兒若行淫玷污自己，就侮辱了父親，要用火將她焚燒。
LEV|21|10|「在弟兄中作大祭司的，頭上倒了膏油，承接聖職，穿了聖衣，不可蓬頭散髮，也不可撕裂衣服；
LEV|21|11|不可挨近任何死屍，即使為了父母也不可玷污自己。
LEV|21|12|他不可出聖所，免得褻瀆了上帝的聖所，因為在他身上有上帝的膏油為聖冕。我是耶和華。
LEV|21|13|他要娶處女為妻。
LEV|21|14|大祭司不可娶寡婦，被休的婦人，或被玷污的妓女為妻；他只可以娶自己百姓中的處女為妻。
LEV|21|15|他不可在自己百姓中侮辱他的兒女，因為我是使他分別為聖的耶和華。」
LEV|21|16|耶和華吩咐 摩西 說：
LEV|21|17|「你吩咐 亞倫 說：你世世代代的後裔，凡有殘疾的都不可近前來獻上帝的食物。
LEV|21|18|因為凡有殘疾的，無論是失明的、瘸腿的、五官不正的、肢體之一過長的、
LEV|21|19|斷腳的、斷手的、
LEV|21|20|駝背的、侏儒的、有眼疾的、長癬的、長疥的，或是睪丸壓傷的，都不可近前來。
LEV|21|21|亞倫 祭司的後裔，凡有殘疾的都不可近前來獻耶和華的火祭。他有殘疾，不可近前來獻上帝的食物。
LEV|21|22|上帝的食物，無論是聖的，或是至聖的，他都可以吃。
LEV|21|23|但他不可進到幔子前，也不可挨近祭壇前，因為他有殘疾，免得他褻瀆我的聖所。我是使他們分別為聖的耶和華。」
LEV|21|24|於是， 摩西 吩咐了 亞倫 和他的兒子，以及 以色列 眾人。
LEV|22|1|耶和華吩咐 摩西 說：
LEV|22|2|「你要吩咐 亞倫 和他子孫說：你們要謹慎處理 以色列 人所分別為聖，歸給我的聖物，免得褻瀆我的聖名。我是耶和華。
LEV|22|3|你要對他們說：你們世世代代的後裔，凡不潔淨，卻挨近 以色列 人所分別為聖，歸給耶和華的聖物，那人必從我面前剪除。我是耶和華。
LEV|22|4|亞倫 的後裔中，凡有痲瘋病的，或患漏症的，都不可吃聖物，直等他潔淨了。無論誰摸了那因屍體而不潔淨的東西，或遺精的人，
LEV|22|5|或摸到任何使他不潔淨的群聚動物或使他不潔淨的人，無論那人有甚麼不潔淨，
LEV|22|6|摸了這些的人必不潔淨到晚上；若不用水洗身，就不可吃聖物。
LEV|22|7|日落的時候，他就潔淨了，然後可以吃聖物，因為這是他的食物。
LEV|22|8|自然死去的或被野獸撕裂的，他不可吃，免得玷污自己。我是耶和華。
LEV|22|9|他們要遵守我的吩咐，免得因褻瀆聖物 ，擔當自己的罪而死。我是使他們分別為聖的耶和華。
LEV|22|10|「任何外人都不可吃聖物；寄居在祭司家的，或雇工，都不可吃聖物。
LEV|22|11|若是祭司用自己的銀錢買來的人，就可以吃聖物；在他家出生的人也可以吃他的食物。
LEV|22|12|祭司的女兒若嫁給外人，就不可吃舉祭的聖物。
LEV|22|13|但祭司的女兒若成為寡婦或被休，又沒有後裔，她回到父家，好像年輕的時候，就可以吃她父親的食物。只是任何外人都不可吃它。
LEV|22|14|若有人誤吃了聖物，要把聖物加上五分之一交給祭司。
LEV|22|15|祭司不可褻瀆 以色列 人獻給耶和華的聖物，
LEV|22|16|免得他們因吃聖物而自取罪孽。我是使他們分別為聖的耶和華。」
LEV|22|17|耶和華吩咐 摩西 說：
LEV|22|18|「你要吩咐 亞倫 和他子孫，以及 以色列 眾人，對他們說： 以色列 家中的人，或在 以色列 中寄居的 ，若要獻供物給耶和華作燔祭，無論是為所許的願或是甘心獻的，
LEV|22|19|就要將一頭公的，沒有殘疾的牛，或綿羊，或山羊獻上，這樣你們才蒙悅納。
LEV|22|20|凡有殘疾的，你們不可獻上，因為這樣你們必不蒙悅納。
LEV|22|21|若有人從牛群或羊群中，將平安祭獻給耶和華，無論是為還所許特別的願，或是甘心獻的，所獻的必須是健康、無任何殘疾的，才蒙悅納。
LEV|22|22|凡瞎眼的、受傷的、斷腿的、潰爛的、長癬的、長疥的，都不可獻給耶和華，不可在壇上作為火祭獻給耶和華。
LEV|22|23|無論是公牛或小綿羊，若一條腿太長或太短，只可作甘心祭獻上；若用來還願，就不蒙悅納。
LEV|22|24|凡睪丸損傷，或壓碎，或破裂，或閹割的，都不可獻給耶和華；不可在你們的地上行這事。
LEV|22|25|從外人的手裏得到任何這類的動物，也不可獻上作你們上帝的食物；因為牠們有缺陷，有殘疾，牠們必不為你們而蒙悅納。」
LEV|22|26|耶和華吩咐 摩西 說：
LEV|22|27|「剛出生的公牛，或綿羊，或山羊，七天當跟著牠的母親；從第八天起，可以當供物作為耶和華的火祭，這是蒙悅納的。
LEV|22|28|無論是牛或羊，不可在同一日宰牠和牠的小牛小羊。
LEV|22|29|你們宰殺祭牲獻感謝祭給耶和華，要獻得使你們可蒙悅納；
LEV|22|30|要在當天吃，一點也不可留到早晨。我是耶和華。
LEV|22|31|「你們要謹守我的誡命，遵行它們。我是耶和華。
LEV|22|32|你們不可褻瀆我的聖名；我在 以色列 人中要被尊為聖。我是使你們分別為聖的耶和華，
LEV|22|33|曾把你們從 埃及 地領出來，作你們的上帝。我是耶和華。」
LEV|23|1|耶和華吩咐 摩西 說：
LEV|23|2|「你要吩咐 以色列 人，對他們說：以下是我的節期，是你們要宣告為聖會的耶和華的節期。」
LEV|23|3|「六日要做工，第七日是完全安息的安息日，要有聖會；你們任何工都不可做。這是在你們一切的住處向耶和華當守的安息日。」
LEV|23|4|「以下是你們要按時宣告為聖會的耶和華的節期。」
LEV|23|5|「正月十四日黃昏的時候 ，是向耶和華守的逾越節。
LEV|23|6|這月的十五日是向耶和華守的除酵節；你們要吃無酵餅七日。
LEV|23|7|第一日要有聖會，任何勞動的工都不可做；
LEV|23|8|要將火祭獻給耶和華七日。第七日要有聖會，任何勞動的工都不可做。」
LEV|23|9|耶和華吩咐 摩西 說：
LEV|23|10|「你要吩咐 以色列 人，對他們說：你們到了我賜給你們的地，收割莊稼的時候，要把初熟莊稼中的一捆拿來給祭司。
LEV|23|11|他要把這捆在耶和華面前搖一搖，使你們蒙悅納。祭司要在安息日的次日把這捆搖一搖。
LEV|23|12|搖這捆的那一日，你們要獻一隻一歲沒有殘疾的小公綿羊，給耶和華作燔祭。
LEV|23|13|同獻的素祭是十分之二伊法調了油的細麵，作為獻給耶和華馨香的火祭；同獻的澆酒祭是四分之一欣酒。
LEV|23|14|無論是餅，是烘熟的穀物，是新穗子，你們都不可吃；直等到你們把這供物帶來獻給你們上帝的那一天，才可以吃。在你們一切的住處，這要成為你們世世代代永遠的定例。」
LEV|23|15|「你們要從安息日的次日，就是獻那捆莊稼為搖祭的那日起，計算足足的七個安息日。
LEV|23|16|到第七個安息日的次日，共計五十天，你們要將新的素祭獻給耶和華。
LEV|23|17|要從你們的住處取十分之二伊法細麵，加酵烤成兩個搖祭的餅，作為初熟之物獻給耶和華。
LEV|23|18|又要將七隻一歲沒有殘疾的羔羊、一頭公牛犢、兩隻公綿羊和餅一同奉上。這些要和素祭和澆酒祭一同作為燔祭獻給耶和華，作馨香的火祭獻給耶和華。
LEV|23|19|你們要獻一隻公山羊為贖罪祭，兩隻一歲的小公綿羊為平安祭。
LEV|23|20|祭司要把這些和初熟莊稼做成的餅，與兩隻小公綿羊一同在耶和華面前搖一搖，作為搖祭。這些獻給耶和華的聖物是歸給祭司的。
LEV|23|21|在這一日，你們要宣告聖會；任何勞動的工都不可做。在你們一切的住處，這要成為你們世世代代永遠的定例。
LEV|23|22|「你們在自己的地收割莊稼時，不可割盡田的角落，也不可拾取莊稼所掉落的，要把它們留給窮人和寄居的。我是耶和華－你們的上帝。」
LEV|23|23|耶和華吩咐 摩西 說：
LEV|23|24|「你要吩咐 以色列 人說：七月初一，你們要守為完全安息的日子，要吹角作紀念，當有聖會。
LEV|23|25|任何勞動的工都不可做；要將火祭獻給耶和華。」
LEV|23|26|耶和華吩咐 摩西 說：
LEV|23|27|「但是，七月初十是贖罪日；你們要守為聖會，刻苦己心，並要將火祭獻給耶和華。
LEV|23|28|在這一日，任何工都不可做；因為這是贖罪日，要在耶和華－你們的上帝面前贖罪。
LEV|23|29|在這一日，凡不刻苦己心的，必從百姓中剪除。
LEV|23|30|凡在這一日做任何工的，我必將他從百姓中除滅。
LEV|23|31|任何工你們都不可做。在你們一切的住處，這要成為你們世世代代永遠的定例。
LEV|23|32|你們要守這日為完全安息的安息日，刻苦己心；從這月初九晚上到次日晚上，你們要守為安息日。」
LEV|23|33|耶和華吩咐 摩西 說：
LEV|23|34|「你要吩咐 以色列 人說：這七月十五日是住棚節，要向耶和華守這節七日。
LEV|23|35|第一日當有聖會，任何勞動的工都不可做。
LEV|23|36|要將火祭獻給耶和華七日。第八日當守聖會，並要獻火祭給耶和華。這是嚴肅會，任何勞動的工都不可做。
LEV|23|37|「這是耶和華的節期，就是你們要宣告為聖會的節期；要將火祭，就是燔祭、素祭、祭物和澆酒祭，按照每日的規定獻給耶和華。
LEV|23|38|除此之外，還有耶和華的安息日，你們獻給耶和華的供物，一切的還願祭，和一切的甘心祭。
LEV|23|39|「但是，從七月十五日起，你們收藏了地的出產之後，要守耶和華的節期七日。第一日為要完全安息，第八日也要完全安息。
LEV|23|40|第一日，你們要拿美好樹上的果子、棕樹枝、樹葉茂密的枝條和河邊的柳枝，在耶和華－你們的上帝面前歡樂七日。
LEV|23|41|每年你們要向耶和華守這節七日。你們在七月裏所守的節，要成為世世代代永遠的定例。
LEV|23|42|你們要住在棚裏七日；凡 以色列 家出生的人都要住在棚裏，
LEV|23|43|好叫你們世世代代知道，我領 以色列 人出 埃及 地的時候，曾使他們住在棚裏。我是耶和華－你們的上帝。」
LEV|23|44|於是， 摩西 向 以色列 人頒佈了耶和華的節期。
LEV|24|1|耶和華吩咐 摩西 說：
LEV|24|2|「你要吩咐 以色列 人，把那搗成的純橄欖油拿來給你，用以點燈，使燈經常點著。
LEV|24|3|在會幕中法櫃前的幔子外， 亞倫 從晚上到早晨要在耶和華面前照管這燈。這要成為你們世世代代永遠的定例。
LEV|24|4|他要在耶和華面前經常照管純金 燈臺上的燈。」
LEV|24|5|「你要取細麵，烤成十二個餅，每個用十分之二伊法。
LEV|24|6|要把餅排成兩行 ，每行六個，供在耶和華面前的純金桌子上。
LEV|24|7|再把純乳香撒在每行餅上，作為紀念，是獻給耶和華為食物的火祭。
LEV|24|8|每個安息日， 亞倫 要把餅不間斷地供在耶和華面前。這是 以色列 人永遠的約。
LEV|24|9|這餅要歸給 亞倫 和他的子孫。他們要在聖處吃這餅，因為在獻給耶和華的火祭中，這餅是至聖的，歸給他作永遠當得的份。」
LEV|24|10|有一個 以色列 婦人的兒子，他父親是 埃及 人。有一日他出去，到 以色列 人中。這 以色列 婦人的兒子和一個 以色列 人在營裏爭吵。
LEV|24|11|以色列 婦人的兒子詛咒，褻瀆了聖名。有人把他送到 摩西 那裏。他的母親名叫 示羅密 ，是 但 支派 底伯利 的女兒。
LEV|24|12|他們把這人收押在監裏，等候耶和華指示的話。
LEV|24|13|耶和華吩咐 摩西 說：
LEV|24|14|「把那詛咒的人帶到營外。凡聽見的人都要把手放在他頭上，全會眾要用石頭打死他。
LEV|24|15|你要吩咐 以色列 人說：凡詛咒上帝的，必要擔當自己的罪。
LEV|24|16|褻瀆耶和華名的，必被處死；全會眾必須用石頭打死他。無論是寄居的，是本地人，他褻瀆聖名的時候必被處死。
LEV|24|17|「打死人的，必被處死；
LEV|24|18|打死牲畜的，必賠上牲畜，以命償命。
LEV|24|19|人若傷害鄰舍以致殘疾，他怎樣做，也要照樣向他做：
LEV|24|20|以傷還傷，以眼還眼，以牙還牙。他怎樣使人有殘疾，也要照樣向他做。
LEV|24|21|打死牲畜的，必賠上牲畜；打死人的，必被處死。
LEV|24|22|無論是寄居的，是本地人，都依照同一條例。我是耶和華－你們的上帝。」
LEV|24|23|於是， 摩西 吩咐 以色列 人，他們就把那詛咒的人帶到營外，用石頭打死。 以色列 人就照耶和華所吩咐 摩西 的做了。
LEV|25|1|耶和華在 西奈山 吩咐 摩西 說：
LEV|25|2|「你要吩咐 以色列 人，對他們說：你們到了我所賜你們那地的時候，地要休耕，向耶和華守安息。
LEV|25|3|你們六年要耕種田地，六年要修整葡萄園，收藏地的出產。
LEV|25|4|第七年，地要守完全安息的安息年，就是向耶和華守安息。你們不可耕種田地，也不可修整葡萄園。
LEV|25|5|不可收割自然生長的莊稼，也不可摘取沒有修剪的葡萄樹上的葡萄。這年，地要完全安息。
LEV|25|6|地在安息年所長出的，要給你和你的奴僕、使女、雇工，以及寄居在你那裏的外人作食物。
LEV|25|7|所有的出產也要給你的牲畜和你地上的走獸作食物。」
LEV|25|8|「你要計算七個安息年，就是七個七年。這就成為你的七個安息年，一共四十九年。
LEV|25|9|七月初十，你要大聲吹角；這是贖罪日，你要在全地吹角。
LEV|25|10|你們要以第五十年為聖年，在全地向所有的居民宣告自由。這是你們的禧年，各人的產業要歸還自己，各人要歸回自己的家。
LEV|25|11|第五十年要作為你們的禧年。你們不可耕種，不可收割自然生長的莊稼，也不可摘取沒有修剪的葡萄樹上的葡萄。
LEV|25|12|因為這是禧年，是你們的聖年；你們要吃地中自然生長的農作物。
LEV|25|13|「這禧年，你們各人的產業要歸還自己。
LEV|25|14|無論你賣甚麼給鄰舍，或從鄰舍的手中買甚麼，彼此不可虧負。
LEV|25|15|你要按照禧年後的年數向鄰舍買；他要按照可收成的年數賣給你；
LEV|25|16|年數越多，價錢就越高；年數越少，價錢就越低，因為他賣給你的是收成的數量。
LEV|25|17|你們彼此不可虧負，只要敬畏你的上帝，因為我是耶和華－你們的上帝。」
LEV|25|18|「你們要遵行我的律例，謹守我的典章，遵行它們，就可以在那地上安然居住。
LEV|25|19|地必出產果實，你們可以吃飽，在那地上安然居住。
LEV|25|20|你們若說：『看哪，第七年我們不耕種，也不收藏農作物，我們吃甚麼呢？』
LEV|25|21|我必在第六年發令賜福給你們，地就長出三年的農作物來。
LEV|25|22|第八年你們要耕種，也要吃陳糧；等到第九年農作物收成的時候，你們還有陳糧吃。」
LEV|25|23|「地不可以賣斷，因為地是我的；你們在我面前是客旅，是寄居的。
LEV|25|24|在你們所得為業的全地，要准許人有權將地贖回。
LEV|25|25|「你的弟兄若漸漸貧窮，賣了他的一些產業，他的至親就要來把弟兄所賣的贖回。
LEV|25|26|若沒有人能為他贖回，他的手頭漸漸寬裕，能夠贖回，
LEV|25|27|就要計算賣後的年數，把剩餘年數的價錢歸還給那買主，他的地業便歸還自己。
LEV|25|28|若他手頭的財力不夠贖回，所賣的地就要留在買主的手裏，直到禧年。到了禧年，地業要歸還賣主。
LEV|25|29|「人若賣城牆內的住宅，賣了以後，一整年內他有權贖回；這是他可以贖回的期限。
LEV|25|30|若他在一整年內不贖回，這有牆之城的房屋就確定永歸買主，直到世世代代；在禧年也不必歸還。
LEV|25|31|但周圍無城牆之村莊的房屋，要看為鄉下的田地，可以贖回；到了禧年就要歸還。
LEV|25|32|至於 利未 人所得為業的城鎮， 利未 人可以隨時贖回他們城鎮中的房屋。
LEV|25|33|在所得為業的城鎮， 利未 人若賣了房屋，又不贖回，到了禧年仍要歸還原主，因為 利未 人城鎮的房屋是他們在 以色列 人中的產業。
LEV|25|34|但是 利未 人各城郊外之地是不可賣的，因為這是他們永遠的產業。」
LEV|25|35|「你的弟兄在你那裏若漸漸貧窮，手頭缺乏，你就要幫補他，使他與你一同生活，像外人和寄居的一樣。
LEV|25|36|不可向他取利息，也不可向他索取高利；要敬畏你的上帝，使你的弟兄與你一同生活。
LEV|25|37|你不可為了利息借錢給他，也不可為了高利而借糧。
LEV|25|38|我是耶和華－你們的上帝，曾領你們從 埃及 地出來，為要把 迦南 地賜給你們，要作你們的上帝。
LEV|25|39|「你的弟兄在你那裏若漸漸貧窮，將自己賣給你，你不可叫他像奴僕服事你。
LEV|25|40|他在你那裏要像雇工和寄居的，服事你直到禧年。
LEV|25|41|他和他兒女要離開你，一同出去，歸回自己的家，回到他祖宗的地業去。
LEV|25|42|因為他們是我的僕人，是我從 埃及 地領出來的。他們不可被賣為奴僕。
LEV|25|43|不可苛刻管轄他，只要敬畏你的上帝。
LEV|25|44|至於你所要的奴僕和使女，可以來自你們四圍的列國，你們可以從他們中買奴僕和使女。
LEV|25|45|那些寄居在你們中間的外人和他們的家屬，就是在你們地上所生的，你們可以從其中買人；他們要作你們的產業。
LEV|25|46|你們可以把他們遺留給你們後代的子孫，作為永遠繼承的產業；你們可以使他們作奴僕。至於你們的弟兄 以色列 人，你們彼此不可苛刻管轄。
LEV|25|47|「住在你那裏的外人或寄居的，若手頭漸漸寬裕，你的弟兄卻漸漸貧窮，將自己賣給那外人或寄居的，或外人家族的一支，
LEV|25|48|賣了以後，有權把自己贖回。他弟兄中的一位可以把他贖回。
LEV|25|49|他的叔伯或叔伯的兒子可以贖他。他家族中的骨肉之親也可以贖他。他自己若手頭漸漸寬裕，也可以贖回自己。
LEV|25|50|他要跟買主計算，從賣自己的那年起，算到禧年；所賣的價錢要按照年數計算，就是雇工跟買主在一起的日子。
LEV|25|51|若剩餘的年數多，就要按著年數從買價中償還他的贖價。
LEV|25|52|若到禧年只剩下幾年，就要按著年數跟買主計算，償還他的贖價。
LEV|25|53|他和買主同住，要像按年雇用的工人，買主不可苛刻管轄他。
LEV|25|54|他若不這樣被贖，到了禧年，仍要和他的兒女一同出去。
LEV|25|55|因為 以色列 人都是我的僕人，他們是我的僕人，是我領他們從 埃及 地出來的。我是耶和華－你們的上帝。」
LEV|26|1|「你們不可為自己造虛無的神明，不可豎立雕刻的偶像或柱像，也不可在你們的地上安放石像，向它跪拜，因為我是耶和華－你們的上帝。
LEV|26|2|你們要謹守我的安息日，敬畏我的聖所。我是耶和華。
LEV|26|3|「你們若遵行我的律例，謹守我的誡命，實行它們，
LEV|26|4|我必按時降雨給你們，使地長出農作物，田野的樹結出果實。
LEV|26|5|你們打穀物要打到摘葡萄的時候，摘葡萄要摘到播種的時候。你們要吃糧食得飽足，在你們的地上安然居住。
LEV|26|6|我要賜平安在地上；你們躺臥，無人驚嚇。我要使你們地上的惡獸消滅，刀劍必不穿越你們的地。
LEV|26|7|你們要追趕仇敵，他們必倒在你們刀下。
LEV|26|8|你們五個人要追趕一百人，一百人要追趕一萬人；仇敵必在你們面前倒在刀下。
LEV|26|9|我要眷顧你們，使你們生養眾多，也要與你們堅立我的約。
LEV|26|10|你們要吃儲存的陳糧，又要為新糧清理陳糧。
LEV|26|11|我要在你們中間立我的帳幕，我的心也不厭惡你們。
LEV|26|12|我要行走在你們中間，作你們的上帝，你們要作我的子民。
LEV|26|13|我是耶和華－你們的上帝，曾將你們從 埃及 地領出來，使你們不再作 埃及 人的奴僕；我曾折斷你們所負的軛，使你們挺身前行。」
LEV|26|14|「你們若不聽從我，不遵行我這一切的誡命，
LEV|26|15|厭棄我的律例，心中厭惡我的典章，不遵行我一切的誡命，背棄了我的約，
LEV|26|16|我就要這樣對待你們：我必使驚惶臨到你們，使你們患癆病，害熱病，以致眼睛失明，身體衰弱。你們要白白撒種，因為仇敵要吃盡你們所種的。
LEV|26|17|我要向你們變臉，使你們敗在仇敵的面前。恨惡你們的必管轄你們；無人追趕，你們卻要逃跑。
LEV|26|18|如果這樣，你們還不聽從我，我就要因你們的罪，加重七倍懲罰你們。
LEV|26|19|我必粉碎你們因勢力而有的驕傲，又要使你們的天堅如鐵，地硬如銅。
LEV|26|20|你們勞力卻白費，因為你們的地沒有出產，地上的樹也不結果實。
LEV|26|21|「你們行事若與我作對，不肯聽從我，我就要因你們的罪，加重七倍災禍擊打你們。
LEV|26|22|我要打發野地的走獸到你們中間，奪去你們的兒女，吞滅你們的牲畜，使你們人數減少，道路荒涼。
LEV|26|23|「如果這樣，你們還不接受管教歸向我，行事與我作對，
LEV|26|24|我就要行事與你們作對，因你們的罪，加重七倍擊打你們。
LEV|26|25|我要使刀劍臨到你們，報復你們的背約。你們若被趕入城中，我要降瘟疫在你們中間，把你們交在仇敵手中。
LEV|26|26|我要斷絕你們糧食的供應 ，使十個女人用一個烤爐給你們烤餅，按配給的定量秤給你們。你們要吃，卻吃不飽。
LEV|26|27|「如果這樣，你們還不聽從我，行事與我作對，
LEV|26|28|我就要向你們發烈怒，行事與你們作對，因你們的罪，加重七倍懲罰你們。
LEV|26|29|你們要吃你們兒子的肉，也要吃你們女兒的肉。
LEV|26|30|我要摧毀你們的丘壇，砍掉你們的香壇，把你們的屍首扔在你們偶像的殘骸上。我的心也必厭惡你們，
LEV|26|31|使你們的城鎮變成廢墟，你們的眾聖所變荒涼，我也不聞你們芬芳的香氣。
LEV|26|32|我要使這地變荒涼，甚至佔領這地的敵人都驚訝。
LEV|26|33|我要把你們驅散到列國中，也要拔刀追趕你們。你們的地要成為荒涼，你們的城鎮要變成廢墟。
LEV|26|34|「當你們在敵人之地的時候，你們的地要在一切荒涼的日子重享安息；在那時候，地要休息，重享安息。
LEV|26|35|地在一切荒涼的日子都要安息，這是你們住在其上的時候所不能得的安息。
LEV|26|36|至於你們倖存的人，我要使他們在敵人之地心中驚慌，甚至風吹落葉的聲音也把他們嚇跑。他們要逃避，像人逃避刀劍，雖無人追趕，卻要跌倒。
LEV|26|37|雖然無人追趕，他們卻要彼此絆倒，像逃避刀劍一樣。你們在仇敵面前必站立不住。
LEV|26|38|你們要在列國中滅亡，敵人之地要吞滅你們，
LEV|26|39|你們倖存的人必因自己的罪孽在敵人之地衰殘，也要因祖先的罪孽衰殘。
LEV|26|40|「他們要承認自己的罪孽和祖先的罪孽，就是背叛我，行事與我作對的過犯。
LEV|26|41|我也行事與他們作對，把他們遣送到敵人之地。那時，他們未受割禮的心若肯謙卑，也服了罪孽的懲罰，
LEV|26|42|我就要記念我與 雅各 的約，記念我與 以撒 的約，與 亞伯拉罕 的約；我也要記念這地。
LEV|26|43|地被他們離棄，因他們不在而荒涼的時候，就要重享安息。他們服了罪孽的懲罰，因為他們厭棄我的典章，心中厭惡我的律例。
LEV|26|44|雖然如此，當他們在敵人之地時，我卻不厭棄他們，不厭惡他們，將他們全然滅絕，也不背棄我與他們的約，因為我是耶和華－他們的上帝。
LEV|26|45|我要為他們的緣故記念我與他們祖先的約；我在列國眼前曾把他們的祖先從 埃及 地領出來，為要作他們的上帝。我是耶和華。」
LEV|26|46|這些律例、典章和法度是耶和華在 西奈山 上藉著 摩西 與 以色列 人立的。
LEV|27|1|耶和華吩咐 摩西 說：
LEV|27|2|「你要吩咐 以色列 人，對他們說：人向耶和華許特別的願，要按照你所估一個人的價錢。
LEV|27|3|你所估的是：二十歲到六十歲男的，按照聖所的舍客勒，估價是五十舍客勒銀子。
LEV|27|4|若是女的，估價是三十舍客勒。
LEV|27|5|五歲到二十歲男的，估價是二十舍客勒，女的十舍客勒。
LEV|27|6|一個月到五歲男的，估價是五舍客勒，女的三舍客勒。
LEV|27|7|六十歲以上男的，估價是十五舍客勒，女的十舍客勒。
LEV|27|8|他若貧窮，不能按照你的估價，就要把他帶到祭司面前，讓祭司為他估價；祭司要按許願者手頭財力所及估價。
LEV|27|9|「許願要獻給耶和華的供物若是牲畜，凡這類獻給耶和華的都要成為聖。
LEV|27|10|不可更換，也不可用另一隻取代，無論是好的換壞的，或是壞的換好的，都不可。若一定要以牲畜取代牲畜，所許的與所取代的都要成為聖。
LEV|27|11|若牲畜不潔淨，不可獻給耶和華為供物，就要把牲畜帶到祭司面前。
LEV|27|12|祭司要估價；牲畜是好是壞，祭司怎樣估定，就是你的估價。
LEV|27|13|許願者若一定要把牠贖回，就要在你的估價上加五分之一。
LEV|27|14|「人將房屋分別為聖，歸給耶和華為聖，祭司就要估價。房屋是好是壞，祭司怎樣估定，就要以他的估價為準。
LEV|27|15|將房屋分別為聖的人，若要贖回房屋，必須付你所估定的價錢，再加上五分之一，房屋才可以歸還給他。
LEV|27|16|「人若將所繼承的一塊田地分別為聖，歸給耶和華，就要按照這地撒種多少來估價；能撒一賀梅珥大麥種子的，是五十舍客勒銀子。
LEV|27|17|他若從禧年起將地分別為聖，就要以你的估價為準。
LEV|27|18|倘若他在禧年以後將地分別為聖，祭司就要按照從那時到下一個禧年所剩的年數推算，從你的估價中減掉。
LEV|27|19|將地分別為聖的人若要把地贖回，必須付你所估定的價錢，再加上五分之一，地才可以歸還給他。
LEV|27|20|他若不贖回那地，或是將地賣給別人，就不能再贖了。
LEV|27|21|到了禧年，那田地要從買主手中退還，歸耶和華為聖，和永獻的地一樣，要歸祭司為業。
LEV|27|22|若分別為聖歸耶和華的田地不是繼承的，而是買來的，
LEV|27|23|祭司就要依照你的估價，推算到禧年。當天，這人要將你所估的歸給耶和華為聖。
LEV|27|24|到了禧年，那田地要退還給賣主，就是繼承那地的原主。
LEV|27|25|凡你所估的價錢都要按照聖所的舍客勒：二十季拉是一舍客勒。
LEV|27|26|「頭生的，就是牲畜中頭生屬耶和華的，人不可再將牠分別為聖，無論是牛是羊都是耶和華的。
LEV|27|27|頭生的牲畜若是不潔淨的，就要按照所估定的價錢，再加上五分之一，把牠贖回。若不贖回，就要按照你的估價把牠賣了。
LEV|27|28|「但一切永獻作當滅的，就是人從他所有永獻給耶和華作當滅的，無論是人，是牲畜，是他繼承的田地，都不可賣，也不可贖。凡永獻作當滅的都歸耶和華為至聖。
LEV|27|29|凡從人中永獻作當滅的都不可贖，必被處死。
LEV|27|30|「地上所有的，無論是地上的種子，是樹上的果子，十分之一是耶和華的，是歸耶和華為聖的。
LEV|27|31|人若要贖回這十分之一，就要另加五分之一。
LEV|27|32|凡牛群羊群中的十分之一，就是一切從牧人杖下經過的，每第十隻要歸耶和華為聖。
LEV|27|33|不可追究是好是壞，也不可取代；若一定要取代，所取代的和本來當獻的牲畜都要成為聖，不可贖回。」
LEV|27|34|這些是耶和華在 西奈山 為 以色列 人所吩咐 摩西 的命令。
