EPH|1|1|Павло, з волі Божої апостол Христа Ісуса, святим, що в Ефесі, і вірним у Христі Ісусі,
EPH|1|2|нехай буде вам благодать та мир від Бога, Отця нашого, і Господа Ісуса Христа!
EPH|1|3|Благословенний Бог і Отець Господа нашого Ісуса Христа, що нас у Христі поблагословив усяким благословенням духовним у небесах,
EPH|1|4|так як вибрав у Ньому Він нас перше заложення світу, щоб були перед Ним ми святі й непорочні, у любові,
EPH|1|5|призначивши наперед, щоб нас усиновити для Себе Ісусом Христом, за вподобанням волі Своєї,
EPH|1|6|на хвалу слави благодаті Своєї, якою Він обдарував нас в Улюбленім,
EPH|1|7|що маємо в Ньому відкуплення кров'ю Його, прощення провин, через багатство благодаті Його,
EPH|1|8|яку Він намножив у нас у всякій премудрості й розважності,
EPH|1|9|об'явивши нам таємницю волі Своєї за Своїм уподобанням, яке постановив у Самому Собі,
EPH|1|10|для урядження виповнення часів, щоб усе об'єднати в Христі, що на небі, і що на землі.
EPH|1|11|У Нім, що в Нім стали ми й спадкоємцями, бувши призначені наперед постановою Того, Хто все чинить за радою волі Своєї,
EPH|1|12|щоб на хвалу Його слави були ми, що перше надіялися на Христа.
EPH|1|13|У Ньому й ви, як почули були слово істини, Євангелію спасіння свого, та в Нього й увірували, запечатані стали Святим Духом обітниці,
EPH|1|14|Який є завдаток нашого спадку, на викуп здобутого, на хвалу Його слави!
EPH|1|15|Тому й я, прочувши про вашу віру в Господа Ісуса, і про любов до всіх святих,
EPH|1|16|не перестаю за вас дякувати, і в молитвах своїх за вас згадую,
EPH|1|17|щоб Бог Господа нашого Ісуса Христа, Отець слави, дав вам Духа премудрости та відкриття для пізнання Його,
EPH|1|18|просвітив очі вашого серця, щоб ви зрозуміли, до якої надії Він вас закликає, і який багатий Його славний спадок у святих,
EPH|1|19|і яка безмірна велич Його сили в нас, що віруємо за виявленням потужної сили Його,
EPH|1|20|яку виявив Він у Христі, воскресивши із мертвих Його, і посадивши на небі праворуч Себе,
EPH|1|21|вище від усякого уряду, і влади, і сили, і панування, і всякого ймення, що назване не тільки в цім віці, але й у майбутньому.
EPH|1|22|І все впокорив Він під ноги Йому, і Його дав найвище за все за Голову Церкви,
EPH|1|23|а вона Його тіло, повня Того, що все всім наповняє!
EPH|2|1|І вас, що мертві були через ваші провини й гріхи,
EPH|2|2|в яких ви колись проживали за звичаєм віку цього, за волею князя, що панує в повітрі, духа, що працює тепер у неслухняних,
EPH|2|3|між якими й усі ми проживали колись у пожадливостях нашого тіла, як чинили волю тіла й думок, і з природи були дітьми гніву, як і інші,
EPH|2|4|Бог же, багатий на милосердя, через Свою превелику любов, що нею Він нас полюбив,
EPH|2|5|і нас, що мертві були через прогріхи, оживив разом із Христом, спасені ви благодаттю,
EPH|2|6|і разом із Ним воскресив, і разом із Ним посадив на небесних місцях у Христі Ісусі,
EPH|2|7|щоб у наступних віках показати безмірне багатство благодаті Своєї в добрості до нас у Христі Ісусі.
EPH|2|8|Бо спасені ви благодаттю через віру, а це не від вас, то дар Божий,
EPH|2|9|не від діл, щоб ніхто не хвалився.
EPH|2|10|Бо ми Його твориво, створені в Христі Ісусі на добрі діла, які Бог наперед приготував, щоб ми в них перебували.
EPH|2|11|Отож, пам'ятайте, що ви, колись тілом погани, що вас так звані рукотворно обрізані на тілі звуть необрізаними,
EPH|2|12|що ви того часу були без Христа, відлучені від громади ізраїльської, і чужі заповітам обітниці, не мавши надії й без Бога на світі.
EPH|2|13|А тепер у Христі Ісусі ви, що колись далекі були, стали близькі Христовою кров'ю.
EPH|2|14|Він бо наш мир, що вчинив із двох одне й зруйнував серединну перегороду, ворожнечу, Своїм тілом,
EPH|2|15|Він Своєю наукою знищив Закона заповідей, щоб з обох збудувати Собою одного нового чоловіка, мир чинивши,
EPH|2|16|і хрестом примирити із Богом обох в однім тілі, ворожнечу на ньому забивши.
EPH|2|17|І, прийшовши, Він благовістив мир вам, далеким, і мир близьким,
EPH|2|18|бо обоє Ним маємо приступ у Дусі однім до Отця.
EPH|2|19|Отже, ви вже не чужі й не приходьки, а співгорожани святим, і домашні для Бога,
EPH|2|20|збудовані на основі апостолів і пророків, де наріжним каменем є Сам Ісус Христос,
EPH|2|21|що на ньому вся будівля, улад побудована, росте в святий храм у Господі,
EPH|2|22|що на ньому і ви разом будуєтеся Духом на оселю Божу.
EPH|3|1|Через це я, Павло, є в'язень Ісуса Христа за вас, поган,
EPH|3|2|якщо ви тільки чули про зарядження Божої благодаті, що для вас мені дана.
EPH|3|3|Бо мені відкриттям об'явилась була таємниця, як писав я вам коротко вище,
EPH|3|4|з чого можете ви, читаючи, пізнати моє розуміння таємниці Христової.
EPH|3|5|А вона за інших поколінь не була оголошена людським синам, як відкрилась тепер через Духа Його святим апостолам і пророкам,
EPH|3|6|що погани співспадкоємці, і одне тіло, і співучасники Його обітниці в Христі Ісусі через Євангелію,
EPH|3|7|якій служителем я став через дар благодаті Божої, що дана мені чином сили Його.
EPH|3|8|Мені, найменшому від усіх святих, дана була оця благодать, благовістити поганам недосліджене багатство Христове,
EPH|3|9|та висвітлити, що то є зарядження таємниці, яка від віків захована в Бозі, Який створив усе,
EPH|3|10|щоб тепер через Церкву була оголошена початкам та владам на небі найрізніша мудрість Божа,
EPH|3|11|за відвічної постанови, яку Він учинив у Христі Ісусі, Господі нашім,
EPH|3|12|в Якім маємо відвагу та доступ у надії через віру в Нього.
EPH|3|13|Тому то благаю я вас не занепадати духом через терпіння моє через вас, бо воно ваша слава.
EPH|3|14|Для того схиляю коліна свої перед Отцем,
EPH|3|15|що від Нього має ймення кожен рід на небі й на землі,
EPH|3|16|щоб Він дав вам за багатством слави Своєї силою зміцнитися через Духа Його в чоловікові внутрішнім,
EPH|3|17|щоб Христос через віру замешкав у ваших серцях, щоб ви, закорінені й основані в любові,
EPH|3|18|змогли зрозуміти зо всіма святими, що то ширина й довжина, і глибина й вишина,
EPH|3|19|і пізнати Христову любов, яка перевищує знання, щоб були ви наповнені всякою повнотою Божою.
EPH|3|20|А Тому, Хто може зробити значно більш над усе, чого просимо або думаємо, силою, що діє в нас,
EPH|3|21|Тому слава в Церкві та в Христі Ісусі на всі покоління на вічні віки. Амінь.
EPH|4|1|Отож, благаю вас я, в'язень у Господі, щоб ви поводилися гідно покликання, що до нього покликано вас,
EPH|4|2|зо всякою покорою та лагідністю, з довготерпінням, у любові терплячи один одного,
EPH|4|3|пильнуючи зберігати єдність духа в союзі миру.
EPH|4|4|Одне тіло, один дух, як і були ви покликані в одній надії вашого покликання.
EPH|4|5|Один Господь, одна віра, одне хрищення,
EPH|4|6|один Бог і Отець усіх, що Він над усіма, і через усіх, і в усіх.
EPH|4|7|А кожному з нас дана благодать у міру дару Христового.
EPH|4|8|Тому й сказано: Піднявшися на висоту, Ти полонених набрав і людям дав дари!
EPH|4|9|А те, що піднявся був, що то, як не те, що перше й зійшов був до найнижчих місць землі?
EPH|4|10|Хто зійшов був, Той саме й піднявся високо над усі небеса, щоб наповнити все.
EPH|4|11|І Він, отож, настановив одних за апостолів, одних за пророків, а тих за благовісників, а тих за пастирів та вчителів,
EPH|4|12|щоб приготувати святих на діло служби для збудування тіла Христового,
EPH|4|13|аж поки ми всі не досягнемо з'єднання віри й пізнання Сина Божого, Мужа досконалого, у міру зросту Христової повноти,
EPH|4|14|щоб більш не були ми малолітками, що хитаються й захоплюються від усякого вітру науки за людською оманою та за лукавством до хитрого блуду,
EPH|4|15|щоб були ми правдомовні в любові, і в усьому зростали в Нього, а Він Голова, Христос.
EPH|4|16|А з Нього все тіло, складене й зв'язане всяким допомічним суглобом, у міру чинности кожного окремого члена, чинить зріст тіла на будування самого себе любов'ю.
EPH|4|17|Отже, говорю я це й свідкую в Господі, щоб ви більш не поводилися, як поводяться погани в марноті свого розуму,
EPH|4|18|вони запаморочені розумом, відчужені від життя Божого за неуцтво, що в них, за стверділість їхніх сердець,
EPH|4|19|вони отупіли й віддалися розпусті, щоб чинити всяку нечисть із зажерливістю.
EPH|4|20|Але ви не так пізнали Христа,
EPH|4|21|якщо ви чули про Нього, і навчилися в Нім, бо правда в Ісусі,
EPH|4|22|щоб відкинути, за першим поступованням, старого чоловіка, який зотліває в звабливих пожадливостях,
EPH|4|23|та відновлятися духом вашого розуму,
EPH|4|24|і зодягнутися в нового чоловіка, створеного за Богом у справедливості й святості правди.
EPH|4|25|Тому то, неправду відкинувши, говоріть кожен правду до свого ближнього, бо ми члени один для одного.
EPH|4|26|Гнівайтеся, та не грішіть, сонце нехай не заходить у вашому гніві,
EPH|4|27|і місця дияволові не давайте!
EPH|4|28|Хто крав, нехай більше не краде, а краще нехай працює та чинить руками своїми добро, щоб мати подати нужденному.
EPH|4|29|Нехай жадне слово гниле не виходить із уст ваших, але тільки таке, що добре на потрібне збудування, щоб воно подало благодать тим, хто чує.
EPH|4|30|І не засмучуйте Духа Святого Божого, Яким ви запечатані на день викупу.
EPH|4|31|Усяке подратування, і гнів, і лютість, і крик, і лайка нехай буде взято від вас разом із усякою злобою.
EPH|4|32|А ви один до одного будьте ласкаві, милостиві, прощаючи один одному, як і Бог через Христа вам простив!
EPH|5|1|Отже, будьте наслідувачами Богові, як улюблені діти,
EPH|5|2|і поводьтеся в любові, як і Христос полюбив вас, і видав за нас Самого Себе, як дар і жертву Богові на приємні пахощі.
EPH|5|3|А розпуста та нечисть усяка й зажерливість нехай навіть не згадуються поміж вами, як личить святим,
EPH|5|4|і гидота, і марнословство або жарти, що непристойні вам, але краще дякування.
EPH|5|5|Знайте бо це, що жаден розпусник, чи нечистий, або зажерливий, що він ідолянин, не має спадку в Христовому й Божому Царстві!
EPH|5|6|Нехай вас не зводить ніхто словами марнотними, бо гнів Божий приходить за них на неслухняних,
EPH|5|7|тож не будьте їм спільниками!
EPH|5|8|Ви бо були колись темрявою, тепер же ви світло в Господі, поводьтеся, як діти світла,
EPH|5|9|бо плід світла знаходиться в кожній добрості, і праведності, і правді.
EPH|5|10|Допевняйтеся, що приємне для Господа,
EPH|5|11|і не беріть участи в неплідних ділах темряви, а краще й докоряйте.
EPH|5|12|Бо соромно навіть казати про те, що роблять вони потаємно!
EPH|5|13|Усе ж те, що світлом докоряється, стає явне, бо все, що явне стає, то світло.
EPH|5|14|Через це то й говорить: Сплячий, вставай, і воскресни із мертвих, і Христос освітлить тебе!
EPH|5|15|Отож, уважайте, щоб поводитися обережно, не як немудрі, але як мудрі,
EPH|5|16|використовуючи час, дні бо лукаві!
EPH|5|17|Через це не будьте нерозумні, але розумійте, що є воля Господня.
EPH|5|18|І не впивайтесь вином, в якому розпуста, але краще наповнюйтесь Духом,
EPH|5|19|розмовляючи поміж собою псалмами, і гімнами, і піснями духовними, співаючи й граючи в серці своєму для Господа,
EPH|5|20|дякуючи завжди за все Богові й Отцеві в Ім'я Господа нашого Ісуса Христа,
EPH|5|21|корячися один одному у Христовім страху.
EPH|5|22|Дружини, коріться своїм чоловікам, як Господеві,
EPH|5|23|бо чоловік голова дружини, як і Христос Голова Церкви, Сам Спаситель тіла!
EPH|5|24|І як кориться Церква Христові, так і дружини своїм чоловікам у всьому.
EPH|5|25|Чоловіки, любіть своїх дружин, як і Христос полюбив Церкву, і віддав за неї Себе,
EPH|5|26|щоб її освятити, очистивши водяним купелем у слові,
EPH|5|27|щоб поставити її Собі славною Церквою, що не має плями чи вади, чи чогось такого, але щоб була свята й непорочна!
EPH|5|28|Чоловіки повинні любити дружин своїх так, як власні тіла, бо хто любить дружину свою, той любить самого себе.
EPH|5|29|Бо ніколи ніхто не зненавидів власного тіла, а годує та гріє його, як і Христос Церкву,
EPH|5|30|бо ми члени Тіла Його від тіла Його й від костей Його!
EPH|5|31|Покине тому чоловік батька й матір, і пристане до дружини своєї, і будуть обоє вони одним тілом.
EPH|5|32|Ця таємниця велика, а я говорю про Христа та про Церкву!
EPH|5|33|Отже, нехай кожен зокрема із вас любить так свою дружину, як самого себе, а дружина нехай боїться свого чоловіка!
EPH|6|1|Діти, слухайтеся своїх батьків у Господі, бо це справедливе!
EPH|6|2|Шануй свого батька та матір це перша заповідь з обітницею,
EPH|6|3|щоб добре велося тобі, і щоб ти був на землі довголітній!
EPH|6|4|А батьки, не дратуйте дітей своїх, а виховуйте їх в напоминанні й остереженні Божому!
EPH|6|5|Раби, слухайтеся тілесних панів зо страхом і тремтінням у простоті серця вашого, як Христа!
EPH|6|6|Не працюйте тільки про людське око, немов чоловіковгодники, а як раби Христові, чиніть від душі волю Божу,
EPH|6|7|служіть із зичливістю, немов Господеві, а не людям!
EPH|6|8|Знайте, що кожен, коли зробить що добре, те саме одержить від Господа, чи то раб, чи то вільний.
EPH|6|9|А пани, чиніть їм те саме, занехаюйте погрози, знайте, що для вас і для них є на небі Господь, а Він на обличчя не дивиться!
EPH|6|10|Нарешті, мої брати, зміцняйтеся Господом та могутністю сили Його!
EPH|6|11|Зодягніться в повну Божу зброю, щоб могли ви стати проти хитрощів диявольських.
EPH|6|12|Бо ми не маємо боротьби проти крови та тіла, але проти початків, проти влади, проти світоправителів цієї темряви, проти піднебесних духів злоби.
EPH|6|13|Через це візьміть повну Божу зброю, щоб могли ви дати опір дня злого, і, все виконавши, витримати.
EPH|6|14|Отже, стійте, підперезавши стегна свої правдою, і зодягнувшись у броню праведности,
EPH|6|15|і взувши ноги в готовість Євангелії миру.
EPH|6|16|А найбільш над усе візьміть щита віри, яким зможете погасити всі огненні стріли лукавого.
EPH|6|17|Візьміть і шолома спасіння, і меча духовного, який є Слово Боже.
EPH|6|18|Усякою молитвою й благанням кожного часу моліться духом, а для того пильнуйте з повною витривалістю та молитвою за всіх святих,
EPH|6|19|і за мене, щоб дане було мені слово відкрити уста свої, і зо сміливістю провіщати таємницю Євангелії,
EPH|6|20|для якої посол я в кайданах, щоб сміливо про неї звіщати, як належить мені.
EPH|6|21|А щоб знали і ви щось про мене, та що я роблю, то все вам розповість Тихик, улюблений брат і в Господі вірний служитель,
EPH|6|22|якого послав я до вас на це саме, щоб довідалися ви про нас, і щоб ваші серця він потішив.
EPH|6|23|Мир братам і любов із вірою від Бога Отця й Господа Ісуса Христа!
EPH|6|24|Благодать зо всіма, що незмінно люблять Господа нашого Ісуса Христа! Амінь.
