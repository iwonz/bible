RUTH|1|1|In the days when the judges ruled, there was a famine in the land, and a man from Bethlehem in Judah, together with his wife and two sons, went to live for a while in the country of Moab.
RUTH|1|2|The man's name was Elimelech, his wife's name Naomi, and the names of his two sons were Mahlon and Kilion. They were Ephrathites from Bethlehem, Judah. And they went to Moab and lived there.
RUTH|1|3|Now Elimelech, Naomi's husband, died, and she was left with her two sons.
RUTH|1|4|They married Moabite women, one named Orpah and the other Ruth. After they had lived there about ten years,
RUTH|1|5|both Mahlon and Kilion also died, and Naomi was left without her two sons and her husband.
RUTH|1|6|When she heard in Moab that the LORD had come to the aid of his people by providing food for them, Naomi and her daughters-in-law prepared to return home from there.
RUTH|1|7|With her two daughters-in-law she left the place where she had been living and set out on the road that would take them back to the land of Judah.
RUTH|1|8|Then Naomi said to her two daughters-in-law, "Go back, each of you, to your mother's home. May the LORD show kindness to you, as you have shown to your dead and to me.
RUTH|1|9|May the LORD grant that each of you will find rest in the home of another husband." Then she kissed them and they wept aloud
RUTH|1|10|and said to her, "We will go back with you to your people."
RUTH|1|11|But Naomi said, "Return home, my daughters. Why would you come with me? Am I going to have any more sons, who could become your husbands?
RUTH|1|12|Return home, my daughters; I am too old to have another husband. Even if I thought there was still hope for me-even if I had a husband tonight and then gave birth to sons-
RUTH|1|13|would you wait until they grew up? Would you remain unmarried for them? No, my daughters. It is more bitter for me than for you, because the LORD's hand has gone out against me!"
RUTH|1|14|At this they wept again. Then Orpah kissed her mother-in-law good-by, but Ruth clung to her.
RUTH|1|15|"Look," said Naomi, "your sister-in-law is going back to her people and her gods. Go back with her."
RUTH|1|16|But Ruth replied, "Don't urge me to leave you or to turn back from you. Where you go I will go, and where you stay I will stay. Your people will be my people and your God my God.
RUTH|1|17|Where you die I will die, and there I will be buried. May the LORD deal with me, be it ever so severely, if anything but death separates you and me."
RUTH|1|18|When Naomi realized that Ruth was determined to go with her, she stopped urging her.
RUTH|1|19|So the two women went on until they came to Bethlehem. When they arrived in Bethlehem, the whole town was stirred because of them, and the women exclaimed, "Can this be Naomi?"
RUTH|1|20|"Don't call me Naomi, "she told them. "Call me Mara, because the Almighty has made my life very bitter.
RUTH|1|21|I went away full, but the LORD has brought me back empty. Why call me Naomi? The LORD has afflicted me; the Almighty has brought misfortune upon me."
RUTH|1|22|So Naomi returned from Moab accompanied by Ruth the Moabitess, her daughter-in-law, arriving in Bethlehem as the barley harvest was beginning.
RUTH|2|1|Now Naomi had a relative on her husband's side, from the clan of Elimelech, a man of standing, whose name was Boaz.
RUTH|2|2|And Ruth the Moabitess said to Naomi, "Let me go to the fields and pick up the leftover grain behind anyone in whose eyes I find favor." Naomi said to her, "Go ahead, my daughter."
RUTH|2|3|So she went out and began to glean in the fields behind the harvesters. As it turned out, she found herself working in a field belonging to Boaz, who was from the clan of Elimelech.
RUTH|2|4|Just then Boaz arrived from Bethlehem and greeted the harvesters, "The LORD be with you!The LORD bless you!" they called back.
RUTH|2|5|Boaz asked the foreman of his harvesters, "Whose young woman is that?"
RUTH|2|6|The foreman replied, "She is the Moabitess who came back from Moab with Naomi.
RUTH|2|7|She said, 'Please let me glean and gather among the sheaves behind the harvesters.' She went into the field and has worked steadily from morning till now, except for a short rest in the shelter."
RUTH|2|8|So Boaz said to Ruth, "My daughter, listen to me. Don't go and glean in another field and don't go away from here. Stay here with my servant girls.
RUTH|2|9|Watch the field where the men are harvesting, and follow along after the girls. I have told the men not to touch you. And whenever you are thirsty, go and get a drink from the water jars the men have filled."
RUTH|2|10|At this, she bowed down with her face to the ground. She exclaimed, "Why have I found such favor in your eyes that you notice me-a foreigner?"
RUTH|2|11|Boaz replied, "I've been told all about what you have done for your mother-in-law since the death of your husband-how you left your father and mother and your homeland and came to live with a people you did not know before.
RUTH|2|12|May the LORD repay you for what you have done. May you be richly rewarded by the LORD, the God of Israel, under whose wings you have come to take refuge."
RUTH|2|13|"May I continue to find favor in your eyes, my lord," she said. "You have given me comfort and have spoken kindly to your servant-though I do not have the standing of one of your servant girls."
RUTH|2|14|At mealtime Boaz said to her, "Come over here. Have some bread and dip it in the wine vinegar." When she sat down with the harvesters, he offered her some roasted grain. She ate all she wanted and had some left over.
RUTH|2|15|As she got up to glean, Boaz gave orders to his men, "Even if she gathers among the sheaves, don't embarrass her.
RUTH|2|16|Rather, pull out some stalks for her from the bundles and leave them for her to pick up, and don't rebuke her."
RUTH|2|17|So Ruth gleaned in the field until evening. Then she threshed the barley she had gathered, and it amounted to about an ephah.
RUTH|2|18|She carried it back to town, and her mother-in-law saw how much she had gathered. Ruth also brought out and gave her what she had left over after she had eaten enough.
RUTH|2|19|Her mother-in-law asked her, "Where did you glean today? Where did you work? Blessed be the man who took notice of you!" Then Ruth told her mother-in-law about the one at whose place she had been working. "The name of the man I worked with today is Boaz," she said.
RUTH|2|20|"The LORD bless him!" Naomi said to her daughter-in-law. "He has not stopped showing his kindness to the living and the dead." She added, "That man is our close relative; he is one of our kinsman-redeemers."
RUTH|2|21|Then Ruth the Moabitess said, "He even said to me, 'Stay with my workers until they finish harvesting all my grain.'"
RUTH|2|22|Naomi said to Ruth her daughter-in-law, "It will be good for you, my daughter, to go with his girls, because in someone else's field you might be harmed."
RUTH|2|23|So Ruth stayed close to the servant girls of Boaz to glean until the barley and wheat harvests were finished. And she lived with her mother-in-law.
RUTH|3|1|One day Naomi her mother-in-law said to her, "My daughter, should I not try to find a home for you, where you will be well provided for?
RUTH|3|2|Is not Boaz, with whose servant girls you have been, a kinsman of ours? Tonight he will be winnowing barley on the threshing floor.
RUTH|3|3|Wash and perfume yourself, and put on your best clothes. Then go down to the threshing floor, but don't let him know you are there until he has finished eating and drinking.
RUTH|3|4|When he lies down, note the place where he is lying. Then go and uncover his feet and lie down. He will tell you what to do."
RUTH|3|5|"I will do whatever you say," Ruth answered.
RUTH|3|6|So she went down to the threshing floor and did everything her mother-in-law told her to do.
RUTH|3|7|When Boaz had finished eating and drinking and was in good spirits, he went over to lie down at the far end of the grain pile. Ruth approached quietly, uncovered his feet and lay down.
RUTH|3|8|In the middle of the night something startled the man, and he turned and discovered a woman lying at his feet.
RUTH|3|9|"Who are you?" he asked. "I am your servant Ruth," she said. "Spread the corner of your garment over me, since you are a kinsman-redeemer."
RUTH|3|10|"The LORD bless you, my daughter," he replied. "This kindness is greater than that which you showed earlier: You have not run after the younger men, whether rich or poor.
RUTH|3|11|And now, my daughter, don't be afraid. I will do for you all you ask. All my fellow townsmen know that you are a woman of noble character.
RUTH|3|12|Although it is true that I am near of kin, there is a kinsman-redeemer nearer than I.
RUTH|3|13|Stay here for the night, and in the morning if he wants to redeem, good; let him redeem. But if he is not willing, as surely as the LORD lives I will do it. Lie here until morning."
RUTH|3|14|So she lay at his feet until morning, but got up before anyone could be recognized; and he said, "Don't let it be known that a woman came to the threshing floor."
RUTH|3|15|He also said, "Bring me the shawl you are wearing and hold it out." When she did so, he poured into it six measures of barley and put it on her. Then he went back to town.
RUTH|3|16|When Ruth came to her mother-in-law, Naomi asked, "How did it go, my daughter?" Then she told her everything Boaz had done for her
RUTH|3|17|and added, "He gave me these six measures of barley, saying, 'Don't go back to your mother-in-law empty-handed.'"
RUTH|3|18|Then Naomi said, "Wait, my daughter, until you find out what happens. For the man will not rest until the matter is settled today."
RUTH|4|1|Meanwhile Boaz went up to the town gate and sat there. When the kinsman-redeemer he had mentioned came along, Boaz said, "Come over here, my friend, and sit down." So he went over and sat down.
RUTH|4|2|Boaz took ten of the elders of the town and said, "Sit here," and they did so.
RUTH|4|3|Then he said to the kinsman-redeemer, "Naomi, who has come back from Moab, is selling the piece of land that belonged to our brother Elimelech.
RUTH|4|4|I thought I should bring the matter to your attention and suggest that you buy it in the presence of these seated here and in the presence of the elders of my people. If you will redeem it, do so. But if you will not, tell me, so I will know. For no one has the right to do it except you, and I am next in line.I will redeem it," he said.
RUTH|4|5|Then Boaz said, "On the day you buy the land from Naomi and from Ruth the Moabitess, you acquire the dead man's widow, in order to maintain the name of the dead with his property."
RUTH|4|6|At this, the kinsman-redeemer said, "Then I cannot redeem it because I might endanger my own estate. You redeem it yourself. I cannot do it."
RUTH|4|7|(Now in earlier times in Israel, for the redemption and transfer of property to become final, one party took off his sandal and gave it to the other. This was the method of legalizing transactions in Israel.)
RUTH|4|8|So the kinsman-redeemer said to Boaz, "Buy it yourself." And he removed his sandal.
RUTH|4|9|Then Boaz announced to the elders and all the people, "Today you are witnesses that I have bought from Naomi all the property of Elimelech, Kilion and Mahlon.
RUTH|4|10|I have also acquired Ruth the Moabitess, Mahlon's widow, as my wife, in order to maintain the name of the dead with his property, so that his name will not disappear from among his family or from the town records. Today you are witnesses!"
RUTH|4|11|Then the elders and all those at the gate said, "We are witnesses. May the LORD make the woman who is coming into your home like Rachel and Leah, who together built up the house of Israel. May you have standing in Ephrathah and be famous in Bethlehem.
RUTH|4|12|Through the offspring the LORD gives you by this young woman, may your family be like that of Perez, whom Tamar bore to Judah."
RUTH|4|13|So Boaz took Ruth and she became his wife. Then he went to her, and the LORD enabled her to conceive, and she gave birth to a son.
RUTH|4|14|The women said to Naomi: "Praise be to the LORD, who this day has not left you without a kinsman-redeemer. May he become famous throughout Israel!
RUTH|4|15|He will renew your life and sustain you in your old age. For your daughter-in-law, who loves you and who is better to you than seven sons, has given him birth."
RUTH|4|16|Then Naomi took the child, laid him in her lap and cared for him.
RUTH|4|17|The women living there said, "Naomi has a son." And they named him Obed. He was the father of Jesse, the father of David.
RUTH|4|18|This, then, is the family line of Perez: Perez was the father of Hezron,
RUTH|4|19|Hezron the father of Ram, Ram the father of Amminadab,
RUTH|4|20|Amminadab the father of Nahshon, Nahshon the father of Salmon,
RUTH|4|21|Salmon the father of Boaz, Boaz the father of Obed,
RUTH|4|22|Obed the father of Jesse, and Jesse the father of David.
