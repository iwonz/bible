EXOD|1|1|Now these are the names of the children of Israel, which came into Egypt; every man and his household came with Jacob.
EXOD|1|2|Reuben, Simeon, Levi, and Judah,
EXOD|1|3|Issachar, Zebulun, and Benjamin,
EXOD|1|4|Dan, and Naphtali, Gad, and Asher.
EXOD|1|5|And all the souls that came out of the loins of Jacob were seventy souls: for Joseph was in Egypt already.
EXOD|1|6|And Joseph died, and all his brethren, and all that generation.
EXOD|1|7|And the children of Israel were fruitful, and increased abundantly, and multiplied, and waxed exceeding mighty; and the land was filled with them.
EXOD|1|8|Now there arose up a new king over Egypt, which knew not Joseph.
EXOD|1|9|And he said unto his people, Behold, the people of the children of Israel are more and mightier than we:
EXOD|1|10|Come on, let us deal wisely with them; lest they multiply, and it come to pass, that, when there falleth out any war, they join also unto our enemies, and fight against us, and so get them up out of the land.
EXOD|1|11|Therefore they did set over them taskmasters to afflict them with their burdens. And they built for Pharaoh treasure cities, Pithom and Raamses.
EXOD|1|12|But the more they afflicted them, the more they multiplied and grew. And they were grieved because of the children of Israel.
EXOD|1|13|And the Egyptians made the children of Israel to serve with rigor:
EXOD|1|14|And they made their lives bitter with hard bondage, in mortar, and in brick, and in all manner of service in the field: all their service, wherein they made them serve, was with rigor.
EXOD|1|15|And the king of Egypt spake to the Hebrew midwives, of which the name of the one was Shiphrah, and the name of the other Puah:
EXOD|1|16|And he said, When ye do the office of a midwife to the Hebrew women, and see them upon the stools; if it be a son, then ye shall kill him: but if it be a daughter, then she shall live.
EXOD|1|17|But the midwives feared God, and did not as the king of Egypt commanded them, but saved the men children alive.
EXOD|1|18|And the king of Egypt called for the midwives, and said unto them, Why have ye done this thing, and have saved the men children alive?
EXOD|1|19|And the midwives said unto Pharaoh, Because the Hebrew women are not as the Egyptian women; for they are lively, and are delivered ere the midwives come in unto them.
EXOD|1|20|Therefore God dealt well with the midwives: and the people multiplied, and waxed very mighty.
EXOD|1|21|And it came to pass, because the midwives feared God, that he made them houses.
EXOD|1|22|And Pharaoh charged all his people, saying, Every son that is born ye shall cast into the river, and every daughter ye shall save alive.
EXOD|2|1|And there went a man of the house of Levi, and took to wife a daughter of Levi.
EXOD|2|2|And the woman conceived, and bare a son: and when she saw him that he was a goodly child, she hid him three months.
EXOD|2|3|And when she could not longer hide him, she took for him an ark of bulrushes, and daubed it with slime and with pitch, and put the child therein; and she laid it in the flags by the river's brink.
EXOD|2|4|And his sister stood afar off, to wit what would be done to him.
EXOD|2|5|And the daughter of Pharaoh came down to wash herself at the river; and her maidens walked along by the river's side; and when she saw the ark among the flags, she sent her maid to fetch it.
EXOD|2|6|And when she had opened it, she saw the child: and, behold, the babe wept. And she had compassion on him, and said, This is one of the Hebrews' children.
EXOD|2|7|Then said his sister to Pharaoh's daughter, Shall I go and call to thee a nurse of the Hebrew women, that she may nurse the child for thee?
EXOD|2|8|And Pharaoh's daughter said to her, Go. And the maid went and called the child's mother.
EXOD|2|9|And Pharaoh's daughter said unto her, Take this child away, and nurse it for me, and I will give thee thy wages. And the women took the child, and nursed it.
EXOD|2|10|And the child grew, and she brought him unto Pharaoh's daughter, and he became her son. And she called his name Moses: and she said, Because I drew him out of the water.
EXOD|2|11|And it came to pass in those days, when Moses was grown, that he went out unto his brethren, and looked on their burdens: and he spied an Egyptian smiting an Hebrew, one of his brethren.
EXOD|2|12|And he looked this way and that way, and when he saw that there was no man, he slew the Egyptian, and hid him in the sand.
EXOD|2|13|And when he went out the second day, behold, two men of the Hebrews strove together: and he said to him that did the wrong, Wherefore smitest thou thy fellow?
EXOD|2|14|And he said, Who made thee a prince and a judge over us? intendest thou to kill me, as thou killedst the Egyptian? And Moses feared, and said, Surely this thing is known.
EXOD|2|15|Now when Pharaoh heard this thing, he sought to slay Moses. But Moses fled from the face of Pharaoh, and dwelt in the land of Midian: and he sat down by a well.
EXOD|2|16|Now the priest of Midian had seven daughters: and they came and drew water, and filled the troughs to water their father's flock.
EXOD|2|17|And the shepherds came and drove them away: but Moses stood up and helped them, and watered their flock.
EXOD|2|18|And when they came to Reuel their father, he said, How is it that ye are come so soon to day?
EXOD|2|19|And they said, An Egyptian delivered us out of the hand of the shepherds, and also drew water enough for us, and watered the flock.
EXOD|2|20|And he said unto his daughters, And where is he? why is it that ye have left the man? call him, that he may eat bread.
EXOD|2|21|And Moses was content to dwell with the man: and he gave Moses Zipporah his daughter.
EXOD|2|22|And she bare him a son, and he called his name Gershom: for he said, I have been a stranger in a strange land.
EXOD|2|23|And it came to pass in process of time, that the king of Egypt died: and the children of Israel sighed by reason of the bondage, and they cried, and their cry came up unto God by reason of the bondage.
EXOD|2|24|And God heard their groaning, and God remembered his covenant with Abraham, with Isaac, and with Jacob.
EXOD|2|25|And God looked upon the children of Israel, and God had respect unto them.
EXOD|3|1|Now Moses kept the flock of Jethro his father in law, the priest of Midian: and he led the flock to the backside of the desert, and came to the mountain of God, even to Horeb.
EXOD|3|2|And the angel of the LORD appeared unto him in a flame of fire out of the midst of a bush: and he looked, and, behold, the bush burned with fire, and the bush was not consumed.
EXOD|3|3|And Moses said, I will now turn aside, and see this great sight, why the bush is not burnt.
EXOD|3|4|And when the LORD saw that he turned aside to see, God called unto him out of the midst of the bush, and said, Moses, Moses. And he said, Here am I.
EXOD|3|5|And he said, Draw not nigh hither: put off thy shoes from off thy feet, for the place whereon thou standest is holy ground.
EXOD|3|6|Moreover he said, I am the God of thy father, the God of Abraham, the God of Isaac, and the God of Jacob. And Moses hid his face; for he was afraid to look upon God.
EXOD|3|7|And the LORD said, I have surely seen the affliction of my people which are in Egypt, and have heard their cry by reason of their taskmasters; for I know their sorrows;
EXOD|3|8|And I am come down to deliver them out of the hand of the Egyptians, and to bring them up out of that land unto a good land and a large, unto a land flowing with milk and honey; unto the place of the Canaanites, and the Hittites, and the Amorites, and the Perizzites, and the Hivites, and the Jebusites.
EXOD|3|9|Now therefore, behold, the cry of the children of Israel is come unto me: and I have also seen the oppression wherewith the Egyptians oppress them.
EXOD|3|10|Come now therefore, and I will send thee unto Pharaoh, that thou mayest bring forth my people the children of Israel out of Egypt.
EXOD|3|11|And Moses said unto God, Who am I, that I should go unto Pharaoh, and that I should bring forth the children of Israel out of Egypt?
EXOD|3|12|And he said, Certainly I will be with thee; and this shall be a token unto thee, that I have sent thee: When thou hast brought forth the people out of Egypt, ye shall serve God upon this mountain.
EXOD|3|13|And Moses said unto God, Behold, when I come unto the children of Israel, and shall say unto them, The God of your fathers hath sent me unto you; and they shall say to me, What is his name? what shall I say unto them?
EXOD|3|14|And God said unto Moses, I AM THAT I AM: and he said, Thus shalt thou say unto the children of Israel, I AM hath sent me unto you.
EXOD|3|15|And God said moreover unto Moses, Thus shalt thou say unto the children of Israel, the LORD God of your fathers, the God of Abraham, the God of Isaac, and the God of Jacob, hath sent me unto you: this is my name for ever, and this is my memorial unto all generations.
EXOD|3|16|Go, and gather the elders of Israel together, and say unto them, The LORD God of your fathers, the God of Abraham, of Isaac, and of Jacob, appeared unto me, saying, I have surely visited you, and seen that which is done to you in Egypt:
EXOD|3|17|And I have said, I will bring you up out of the affliction of Egypt unto the land of the Canaanites, and the Hittites, and the Amorites, and the Perizzites, and the Hivites, and the Jebusites, unto a land flowing with milk and honey.
EXOD|3|18|And they shall hearken to thy voice: and thou shalt come, thou and the elders of Israel, unto the king of Egypt, and ye shall say unto him, The LORD God of the Hebrews hath met with us: and now let us go, we beseech thee, three days' journey into the wilderness, that we may sacrifice to the LORD our God.
EXOD|3|19|And I am sure that the king of Egypt will not let you go, no, not by a mighty hand.
EXOD|3|20|And I will stretch out my hand, and smite Egypt with all my wonders which I will do in the midst thereof: and after that he will let you go.
EXOD|3|21|And I will give this people favor in the sight of the Egyptians: and it shall come to pass, that, when ye go, ye shall not go empty.
EXOD|3|22|But every woman shall borrow of her neighbor, and of her that sojourneth in her house, jewels of silver, and jewels of gold, and raiment: and ye shall put them upon your sons, and upon your daughters; and ye shall spoil the Egyptians.
EXOD|4|1|And Moses answered and said, But, behold, they will not believe me, nor hearken unto my voice: for they will say, The LORD hath not appeared unto thee.
EXOD|4|2|And the LORD said unto him, What is that in thine hand? And he said, A rod.
EXOD|4|3|And he said, Cast it on the ground. And he cast it on the ground, and it became a serpent; and Moses fled from before it.
EXOD|4|4|And the LORD said unto Moses, Put forth thine hand, and take it by the tail. And he put forth his hand, and caught it, and it became a rod in his hand:
EXOD|4|5|That they may believe that the LORD God of their fathers, the God of Abraham, the God of Isaac, and the God of Jacob, hath appeared unto thee.
EXOD|4|6|And the LORD said furthermore unto him, Put now thine hand into thy bosom. And he put his hand into his bosom: and when he took it out, behold, his hand was leprous as snow.
EXOD|4|7|And he said, Put thine hand into thy bosom again. And he put his hand into his bosom again; and plucked it out of his bosom, and, behold, it was turned again as his other flesh.
EXOD|4|8|And it shall come to pass, if they will not believe thee, neither hearken to the voice of the first sign, that they will believe the voice of the latter sign.
EXOD|4|9|And it shall come to pass, if they will not believe also these two signs, neither hearken unto thy voice, that thou shalt take of the water of the river, and pour it upon the dry land: and the water which thou takest out of the river shall become blood upon the dry land.
EXOD|4|10|And Moses said unto the LORD, O my LORD, I am not eloquent, neither heretofore, nor since thou hast spoken unto thy servant: but I am slow of speech, and of a slow tongue.
EXOD|4|11|And the LORD said unto him, Who hath made man's mouth? or who maketh the dumb, or deaf, or the seeing, or the blind? have not I the LORD?
EXOD|4|12|Now therefore go, and I will be with thy mouth, and teach thee what thou shalt say.
EXOD|4|13|And he said, O my LORD, send, I pray thee, by the hand of him whom thou wilt send.
EXOD|4|14|And the anger of the LORD was kindled against Moses, and he said, Is not Aaron the Levite thy brother? I know that he can speak well. And also, behold, he cometh forth to meet thee: and when he seeth thee, he will be glad in his heart.
EXOD|4|15|And thou shalt speak unto him, and put words in his mouth: and I will be with thy mouth, and with his mouth, and will teach you what ye shall do.
EXOD|4|16|And he shall be thy spokesman unto the people: and he shall be, even he shall be to thee instead of a mouth, and thou shalt be to him instead of God.
EXOD|4|17|And thou shalt take this rod in thine hand, wherewith thou shalt do signs.
EXOD|4|18|And Moses went and returned to Jethro his father in law, and said unto him, Let me go, I pray thee, and return unto my brethren which are in Egypt, and see whether they be yet alive. And Jethro said to Moses, Go in peace.
EXOD|4|19|And the LORD said unto Moses in Midian, Go, return into Egypt: for all the men are dead which sought thy life.
EXOD|4|20|And Moses took his wife and his sons, and set them upon an ass, and he returned to the land of Egypt: and Moses took the rod of God in his hand.
EXOD|4|21|And the LORD said unto Moses, When thou goest to return into Egypt, see that thou do all those wonders before Pharaoh, which I have put in thine hand: but I will harden his heart, that he shall not let the people go.
EXOD|4|22|And thou shalt say unto Pharaoh, Thus saith the LORD, Israel is my son, even my firstborn:
EXOD|4|23|And I say unto thee, Let my son go, that he may serve me: and if thou refuse to let him go, behold, I will slay thy son, even thy firstborn.
EXOD|4|24|And it came to pass by the way in the inn, that the LORD met him, and sought to kill him.
EXOD|4|25|Then Zipporah took a sharp stone, and cut off the foreskin of her son, and cast it at his feet, and said, Surely a bloody husband art thou to me.
EXOD|4|26|So he let him go: then she said, A bloody husband thou art, because of the circumcision.
EXOD|4|27|And the LORD said to Aaron, Go into the wilderness to meet Moses. And he went, and met him in the mount of God, and kissed him.
EXOD|4|28|And Moses told Aaron all the words of the LORD who had sent him, and all the signs which he had commanded him.
EXOD|4|29|And Moses and Aaron went and gathered together all the elders of the children of Israel:
EXOD|4|30|And Aaron spake all the words which the LORD had spoken unto Moses, and did the signs in the sight of the people.
EXOD|4|31|And the people believed: and when they heard that the LORD had visited the children of Israel, and that he had looked upon their affliction, then they bowed their heads and worshipped.
EXOD|5|1|And afterward Moses and Aaron went in, and told Pharaoh, Thus saith the LORD God of Israel, Let my people go, that they may hold a feast unto me in the wilderness.
EXOD|5|2|And Pharaoh said, Who is the LORD, that I should obey his voice to let Israel go? I know not the LORD, neither will I let Israel go.
EXOD|5|3|And they said, The God of the Hebrews hath met with us: let us go, we pray thee, three days' journey into the desert, and sacrifice unto the LORD our God; lest he fall upon us with pestilence, or with the sword.
EXOD|5|4|And the king of Egypt said unto them, Wherefore do ye, Moses and Aaron, let the people from their works? get you unto your burdens.
EXOD|5|5|And Pharaoh said, Behold, the people of the land now are many, and ye make them rest from their burdens.
EXOD|5|6|And Pharaoh commanded the same day the taskmasters of the people, and their officers, saying,
EXOD|5|7|Ye shall no more give the people straw to make brick, as heretofore: let them go and gather straw for themselves.
EXOD|5|8|And the tale of the bricks, which they did make heretofore, ye shall lay upon them; ye shall not diminish ought thereof: for they be idle; therefore they cry, saying, Let us go and sacrifice to our God.
EXOD|5|9|Let there more work be laid upon the men, that they may labor therein; and let them not regard vain words.
EXOD|5|10|And the taskmasters of the people went out, and their officers, and they spake to the people, saying, Thus saith Pharaoh, I will not give you straw.
EXOD|5|11|Go ye, get you straw where ye can find it: yet not ought of your work shall be diminished.
EXOD|5|12|So the people were scattered abroad throughout all the land of Egypt to gather stubble instead of straw.
EXOD|5|13|And the taskmasters hasted them, saying, Fulfil your works, your daily tasks, as when there was straw.
EXOD|5|14|And the officers of the children of Israel, which Pharaoh's taskmasters had set over them, were beaten, and demanded, Wherefore have ye not fulfilled your task in making brick both yesterday and to day, as heretofore?
EXOD|5|15|Then the officers of the children of Israel came and cried unto Pharaoh, saying, Wherefore dealest thou thus with thy servants?
EXOD|5|16|There is no straw given unto thy servants, and they say to us, Make brick: and, behold, thy servants are beaten; but the fault is in thine own people.
EXOD|5|17|But he said, Ye are idle, ye are idle: therefore ye say, Let us go and do sacrifice to the LORD.
EXOD|5|18|Go therefore now, and work; for there shall no straw be given you, yet shall ye deliver the tale of bricks.
EXOD|5|19|And the officers of the children of Israel did see that they were in evil case, after it was said, Ye shall not minish ought from your bricks of your daily task.
EXOD|5|20|And they met Moses and Aaron, who stood in the way, as they came forth from Pharaoh:
EXOD|5|21|And they said unto them, The LORD look upon you, and judge; because ye have made our savor to be abhorred in the eyes of Pharaoh, and in the eyes of his servants, to put a sword in their hand to slay us.
EXOD|5|22|And Moses returned unto the LORD, and said, LORD, wherefore hast thou so evil entreated this people? why is it that thou hast sent me?
EXOD|5|23|For since I came to Pharaoh to speak in thy name, he hath done evil to this people; neither hast thou delivered thy people at all.
EXOD|6|1|Then the LORD said unto Moses, Now shalt thou see what I will do to Pharaoh: for with a strong hand shall he let them go, and with a strong hand shall he drive them out of his land.
EXOD|6|2|And God spake unto Moses, and said unto him, I am the LORD:
EXOD|6|3|And I appeared unto Abraham, unto Isaac, and unto Jacob, by the name of God Almighty, but by my name JEHOVAH was I not known to them.
EXOD|6|4|And I have also established my covenant with them, to give them the land of Canaan, the land of their pilgrimage, wherein they were strangers.
EXOD|6|5|And I have also heard the groaning of the children of Israel, whom the Egyptians keep in bondage; and I have remembered my covenant.
EXOD|6|6|Wherefore say unto the children of Israel, I am the LORD, and I will bring you out from under the burdens of the Egyptians, and I will rid you out of their bondage, and I will redeem you with a stretched out arm, and with great judgments:
EXOD|6|7|And I will take you to me for a people, and I will be to you a God: and ye shall know that I am the LORD your God, which bringeth you out from under the burdens of the Egyptians.
EXOD|6|8|And I will bring you in unto the land, concerning the which I did swear to give it to Abraham, to Isaac, and to Jacob; and I will give it you for an heritage: I am the LORD.
EXOD|6|9|And Moses spake so unto the children of Israel: but they hearkened not unto Moses for anguish of spirit, and for cruel bondage.
EXOD|6|10|And the LORD spake unto Moses, saying,
EXOD|6|11|Go in, speak unto Pharaoh king of Egypt, that he let the children of Israel go out of his land.
EXOD|6|12|And Moses spake before the LORD, saying, Behold, the children of Israel have not hearkened unto me; how then shall Pharaoh hear me, who am of uncircumcised lips?
EXOD|6|13|And the LORD spake unto Moses and unto Aaron, and gave them a charge unto the children of Israel, and unto Pharaoh king of Egypt, to bring the children of Israel out of the land of Egypt.
EXOD|6|14|These be the heads of their fathers' houses: The sons of Reuben the firstborn of Israel; Hanoch, and Pallu, Hezron, and Carmi: these be the families of Reuben.
EXOD|6|15|And the sons of Simeon; Jemuel, and Jamin, and Ohad, and Jachin, and Zohar, and Shaul the son of a Canaanitish woman: these are the families of Simeon.
EXOD|6|16|And these are the names of the sons of Levi according to their generations; Gershon, and Kohath, and Merari: and the years of the life of Levi were an hundred thirty and seven years.
EXOD|6|17|The sons of Gershon; Libni, and Shimi, according to their families.
EXOD|6|18|And the sons of Kohath; Amram, and Izhar, and Hebron, and Uzziel: and the years of the life of Kohath were an hundred thirty and three years.
EXOD|6|19|And the sons of Merari; Mahali and Mushi: these are the families of Levi according to their generations.
EXOD|6|20|And Amram took him Jochebed his father's sister to wife; and she bare him Aaron and Moses: and the years of the life of Amram were an hundred and thirty and seven years.
EXOD|6|21|And the sons of Izhar; Korah, and Nepheg, and Zichri.
EXOD|6|22|And the sons of Uzziel; Mishael, and Elzaphan, and Zithri.
EXOD|6|23|And Aaron took him Elisheba, daughter of Amminadab, sister of Naashon, to wife; and she bare him Nadab, and Abihu, Eleazar, and Ithamar.
EXOD|6|24|And the sons of Korah; Assir, and Elkanah, and Abiasaph: these are the families of the Korhites.
EXOD|6|25|And Eleazar Aaron's son took him one of the daughters of Putiel to wife; and she bare him Phinehas: these are the heads of the fathers of the Levites according to their families.
EXOD|6|26|These are that Aaron and Moses, to whom the LORD said, Bring out the children of Israel from the land of Egypt according to their armies.
EXOD|6|27|These are they which spake to Pharaoh king of Egypt, to bring out the children of Israel from Egypt: these are that Moses and Aaron.
EXOD|6|28|And it came to pass on the day when the LORD spake unto Moses in the land of Egypt,
EXOD|6|29|That the LORD spake unto Moses, saying, I am the LORD: speak thou unto Pharaoh king of Egypt all that I say unto thee.
EXOD|6|30|And Moses said before the LORD, Behold, I am of uncircumcised lips, and how shall Pharaoh hearken unto me?
EXOD|7|1|And the LORD said unto Moses, See, I have made thee a god to Pharaoh: and Aaron thy brother shall be thy prophet.
EXOD|7|2|Thou shalt speak all that I command thee: and Aaron thy brother shall speak unto Pharaoh, that he send the children of Israel out of his land.
EXOD|7|3|And I will harden Pharaoh's heart, and multiply my signs and my wonders in the land of Egypt.
EXOD|7|4|But Pharaoh shall not hearken unto you, that I may lay my hand upon Egypt, and bring forth mine armies, and my people the children of Israel, out of the land of Egypt by great judgments.
EXOD|7|5|And the Egyptians shall know that I am the LORD, when I stretch forth mine hand upon Egypt, and bring out the children of Israel from among them.
EXOD|7|6|And Moses and Aaron did as the LORD commanded them, so did they.
EXOD|7|7|And Moses was fourscore years old, and Aaron fourscore and three years old, when they spake unto Pharaoh.
EXOD|7|8|And the LORD spake unto Moses and unto Aaron, saying,
EXOD|7|9|When Pharaoh shall speak unto you, saying, Show a miracle for you: then thou shalt say unto Aaron, Take thy rod, and cast it before Pharaoh, and it shall become a serpent.
EXOD|7|10|And Moses and Aaron went in unto Pharaoh, and they did so as the LORD had commanded: and Aaron cast down his rod before Pharaoh, and before his servants, and it became a serpent.
EXOD|7|11|Then Pharaoh also called the wise men and the sorcerers: now the magicians of Egypt, they also did in like manner with their enchantments.
EXOD|7|12|For they cast down every man his rod, and they became serpents: but Aaron's rod swallowed up their rods.
EXOD|7|13|And he hardened Pharaoh's heart, that he hearkened not unto them; as the LORD had said.
EXOD|7|14|And the LORD said unto Moses, Pharaoh's heart is hardened, he refuseth to let the people go.
EXOD|7|15|Get thee unto Pharaoh in the morning; lo, he goeth out unto the water; and thou shalt stand by the river's brink against he come; and the rod which was turned to a serpent shalt thou take in thine hand.
EXOD|7|16|And thou shalt say unto him, The LORD God of the Hebrews hath sent me unto thee, saying, Let my people go, that they may serve me in the wilderness: and, behold, hitherto thou wouldest not hear.
EXOD|7|17|Thus saith the LORD, In this thou shalt know that I am the LORD: behold, I will smite with the rod that is in mine hand upon the waters which are in the river, and they shall be turned to blood.
EXOD|7|18|And the fish that is in the river shall die, and the river shall stink; and the Egyptians shall loathe to drink of the water of the river.
EXOD|7|19|And the LORD spake unto Moses, Say unto Aaron, Take thy rod, and stretch out thine hand upon the waters of Egypt, upon their streams, upon their rivers, and upon their ponds, and upon all their pools of water, that they may become blood; and that there may be blood throughout all the land of Egypt, both in vessels of wood, and in vessels of stone.
EXOD|7|20|And Moses and Aaron did so, as the LORD commanded; and he lifted up the rod, and smote the waters that were in the river, in the sight of Pharaoh, and in the sight of his servants; and all the waters that were in the river were turned to blood.
EXOD|7|21|And the fish that was in the river died; and the river stank, and the Egyptians could not drink of the water of the river; and there was blood throughout all the land of Egypt.
EXOD|7|22|And the magicians of Egypt did so with their enchantments: and Pharaoh's heart was hardened, neither did he hearken unto them; as the LORD had said.
EXOD|7|23|And Pharaoh turned and went into his house, neither did he set his heart to this also.
EXOD|7|24|And all the Egyptians digged round about the river for water to drink; for they could not drink of the water of the river.
EXOD|7|25|And seven days were fulfilled, after that the LORD had smitten the river.
EXOD|8|1|And the LORD spake unto Moses, Go unto Pharaoh, and say unto him, Thus saith the LORD, Let my people go, that they may serve me.
EXOD|8|2|And if thou refuse to let them go, behold, I will smite all thy borders with frogs:
EXOD|8|3|And the river shall bring forth frogs abundantly, which shall go up and come into thine house, and into thy bedchamber, and upon thy bed, and into the house of thy servants, and upon thy people, and into thine ovens, and into thy kneadingtroughs:
EXOD|8|4|And the frogs shall come up both on thee, and upon thy people, and upon all thy servants.
EXOD|8|5|And the LORD spake unto Moses, Say unto Aaron, Stretch forth thine hand with thy rod over the streams, over the rivers, and over the ponds, and cause frogs to come up upon the land of Egypt.
EXOD|8|6|And Aaron stretched out his hand over the waters of Egypt; and the frogs came up, and covered the land of Egypt.
EXOD|8|7|And the magicians did so with their enchantments, and brought up frogs upon the land of Egypt.
EXOD|8|8|Then Pharaoh called for Moses and Aaron, and said, Entreat the LORD, that he may take away the frogs from me, and from my people; and I will let the people go, that they may do sacrifice unto the LORD.
EXOD|8|9|And Moses said unto Pharaoh, Glory over me: when shall I entreat for thee, and for thy servants, and for thy people, to destroy the frogs from thee and thy houses, that they may remain in the river only?
EXOD|8|10|And he said, To morrow. And he said, Be it according to thy word: that thou mayest know that there is none like unto the LORD our God.
EXOD|8|11|And the frogs shall depart from thee, and from thy houses, and from thy servants, and from thy people; they shall remain in the river only.
EXOD|8|12|And Moses and Aaron went out from Pharaoh: and Moses cried unto the LORD because of the frogs which he had brought against Pharaoh.
EXOD|8|13|And the LORD did according to the word of Moses; and the frogs died out of the houses, out of the villages, and out of the fields.
EXOD|8|14|And they gathered them together upon heaps: and the land stank.
EXOD|8|15|But when Pharaoh saw that there was respite, he hardened his heart, and hearkened not unto them; as the LORD had said.
EXOD|8|16|And the LORD said unto Moses, Say unto Aaron, Stretch out thy rod, and smite the dust of the land, that it may become lice throughout all the land of Egypt.
EXOD|8|17|And they did so; for Aaron stretched out his hand with his rod, and smote the dust of the earth, and it became lice in man, and in beast; all the dust of the land became lice throughout all the land of Egypt.
EXOD|8|18|And the magicians did so with their enchantments to bring forth lice, but they could not: so there were lice upon man, and upon beast.
EXOD|8|19|Then the magicians said unto Pharaoh, This is the finger of God: and Pharaoh's heart was hardened, and he hearkened not unto them; as the LORD had said.
EXOD|8|20|And the LORD said unto Moses, Rise up early in the morning, and stand before Pharaoh; lo, he cometh forth to the water; and say unto him, Thus saith the LORD, Let my people go, that they may serve me.
EXOD|8|21|Else, if thou wilt not let my people go, behold, I will send swarms of flies upon thee, and upon thy servants, and upon thy people, and into thy houses: and the houses of the Egyptians shall be full of swarms of flies, and also the ground whereon they are.
EXOD|8|22|And I will sever in that day the land of Goshen, in which my people dwell, that no swarms of flies shall be there; to the end thou mayest know that I am the LORD in the midst of the earth.
EXOD|8|23|And I will put a division between my people and thy people: to morrow shall this sign be.
EXOD|8|24|And the LORD did so; and there came a grievous swarm of flies into the house of Pharaoh, and into his servants' houses, and into all the land of Egypt: the land was corrupted by reason of the swarm of flies.
EXOD|8|25|And Pharaoh called for Moses and for Aaron, and said, Go ye, sacrifice to your God in the land.
EXOD|8|26|And Moses said, It is not meet so to do; for we shall sacrifice the abomination of the Egyptians to the LORD our God: lo, shall we sacrifice the abomination of the Egyptians before their eyes, and will they not stone us?
EXOD|8|27|We will go three days' journey into the wilderness, and sacrifice to the LORD our God, as he shall command us.
EXOD|8|28|And Pharaoh said, I will let you go, that ye may sacrifice to the LORD your God in the wilderness; only ye shall not go very far away: entreat for me.
EXOD|8|29|And Moses said, Behold, I go out from thee, and I will entreat the LORD that the swarms of flies may depart from Pharaoh, from his servants, and from his people, to morrow: but let not Pharaoh deal deceitfully any more in not letting the people go to sacrifice to the LORD.
EXOD|8|30|And Moses went out from Pharaoh, and entreated the LORD.
EXOD|8|31|And the LORD did according to the word of Moses; and he removed the swarms of flies from Pharaoh, from his servants, and from his people; there remained not one.
EXOD|8|32|And Pharaoh hardened his heart at this time also, neither would he let the people go.
EXOD|9|1|Then the LORD said unto Moses, Go in unto Pharaoh, and tell him, Thus saith the LORD God of the Hebrews, Let my people go, that they may serve me.
EXOD|9|2|For if thou refuse to let them go, and wilt hold them still,
EXOD|9|3|Behold, the hand of the LORD is upon thy cattle which is in the field, upon the horses, upon the asses, upon the camels, upon the oxen, and upon the sheep: there shall be a very grievous murrain.
EXOD|9|4|And the LORD shall sever between the cattle of Israel and the cattle of Egypt: and there shall nothing die of all that is the children's of Israel.
EXOD|9|5|And the LORD appointed a set time, saying, To morrow the LORD shall do this thing in the land.
EXOD|9|6|And the LORD did that thing on the morrow, and all the cattle of Egypt died: but of the cattle of the children of Israel died not one.
EXOD|9|7|And Pharaoh sent, and, behold, there was not one of the cattle of the Israelites dead. And the heart of Pharaoh was hardened, and he did not let the people go.
EXOD|9|8|And the LORD said unto Moses and unto Aaron, Take to you handfuls of ashes of the furnace, and let Moses sprinkle it toward the heaven in the sight of Pharaoh.
EXOD|9|9|And it shall become small dust in all the land of Egypt, and shall be a boil breaking forth with blains upon man, and upon beast, throughout all the land of Egypt.
EXOD|9|10|And they took ashes of the furnace, and stood before Pharaoh; and Moses sprinkled it up toward heaven; and it became a boil breaking forth with blains upon man, and upon beast.
EXOD|9|11|And the magicians could not stand before Moses because of the boils; for the boil was upon the magicians, and upon all the Egyptians.
EXOD|9|12|And the LORD hardened the heart of Pharaoh, and he hearkened not unto them; as the LORD had spoken unto Moses.
EXOD|9|13|And the LORD said unto Moses, Rise up early in the morning, and stand before Pharaoh, and say unto him, Thus saith the LORD God of the Hebrews, Let my people go, that they may serve me.
EXOD|9|14|For I will at this time send all my plagues upon thine heart, and upon thy servants, and upon thy people; that thou mayest know that there is none like me in all the earth.
EXOD|9|15|For now I will stretch out my hand, that I may smite thee and thy people with pestilence; and thou shalt be cut off from the earth.
EXOD|9|16|And in very deed for this cause have I raised thee up, for to show in thee my power; and that my name may be declared throughout all the earth.
EXOD|9|17|As yet exaltest thou thyself against my people, that thou wilt not let them go?
EXOD|9|18|Behold, to morrow about this time I will cause it to rain a very grievous hail, such as hath not been in Egypt since the foundation thereof even until now.
EXOD|9|19|Send therefore now, and gather thy cattle, and all that thou hast in the field; for upon every man and beast which shall be found in the field, and shall not be brought home, the hail shall come down upon them, and they shall die.
EXOD|9|20|He that feared the word of the LORD among the servants of Pharaoh made his servants and his cattle flee into the houses:
EXOD|9|21|And he that regarded not the word of the LORD left his servants and his cattle in the field.
EXOD|9|22|And the LORD said unto Moses, Stretch forth thine hand toward heaven, that there may be hail in all the land of Egypt, upon man, and upon beast, and upon every herb of the field, throughout the land of Egypt.
EXOD|9|23|And Moses stretched forth his rod toward heaven: and the LORD sent thunder and hail, and the fire ran along upon the ground; and the LORD rained hail upon the land of Egypt.
EXOD|9|24|So there was hail, and fire mingled with the hail, very grievous, such as there was none like it in all the land of Egypt since it became a nation.
EXOD|9|25|And the hail smote throughout all the land of Egypt all that was in the field, both man and beast; and the hail smote every herb of the field, and brake every tree of the field.
EXOD|9|26|Only in the land of Goshen, where the children of Israel were, was there no hail.
EXOD|9|27|And Pharaoh sent, and called for Moses and Aaron, and said unto them, I have sinned this time: the LORD is righteous, and I and my people are wicked.
EXOD|9|28|Entreat the LORD (for it is enough) that there be no more mighty thunderings and hail; and I will let you go, and ye shall stay no longer.
EXOD|9|29|And Moses said unto him, As soon as I am gone out of the city, I will spread abroad my hands unto the LORD; and the thunder shall cease, neither shall there be any more hail; that thou mayest know how that the earth is the LORD's.
EXOD|9|30|But as for thee and thy servants, I know that ye will not yet fear the LORD God.
EXOD|9|31|And the flax and the barley was smitten: for the barley was in the ear, and the flax was bolled.
EXOD|9|32|But the wheat and the rye were not smitten: for they were not grown up.
EXOD|9|33|And Moses went out of the city from Pharaoh, and spread abroad his hands unto the LORD: and the thunders and hail ceased, and the rain was not poured upon the earth.
EXOD|9|34|And when Pharaoh saw that the rain and the hail and the thunders were ceased, he sinned yet more, and hardened his heart, he and his servants.
EXOD|9|35|And the heart of Pharaoh was hardened, neither would he let the children of Israel go; as the LORD had spoken by Moses.
EXOD|10|1|And the LORD said unto Moses, Go in unto Pharaoh: for I have hardened his heart, and the heart of his servants, that I might show these my signs before him:
EXOD|10|2|And that thou mayest tell in the ears of thy son, and of thy son's son, what things I have wrought in Egypt, and my signs which I have done among them; that ye may know how that I am the LORD.
EXOD|10|3|And Moses and Aaron came in unto Pharaoh, and said unto him, Thus saith the LORD God of the Hebrews, How long wilt thou refuse to humble thyself before me? let my people go, that they may serve me.
EXOD|10|4|Else, if thou refuse to let my people go, behold, to morrow will I bring the locusts into thy coast:
EXOD|10|5|And they shall cover the face of the earth, that one cannot be able to see the earth: and they shall eat the residue of that which is escaped, which remaineth unto you from the hail, and shall eat every tree which groweth for you out of the field:
EXOD|10|6|And they shall fill thy houses, and the houses of all thy servants, and the houses of all the Egyptians; which neither thy fathers, nor thy fathers' fathers have seen, since the day that they were upon the earth unto this day. And he turned himself, and went out from Pharaoh.
EXOD|10|7|And Pharaoh's servants said unto him, How long shall this man be a snare unto us? let the men go, that they may serve the LORD their God: knowest thou not yet that Egypt is destroyed?
EXOD|10|8|And Moses and Aaron were brought again unto Pharaoh: and he said unto them, Go, serve the LORD your God: but who are they that shall go?
EXOD|10|9|And Moses said, We will go with our young and with our old, with our sons and with our daughters, with our flocks and with our herds will we go; for we must hold a feast unto the LORD.
EXOD|10|10|And he said unto them, Let the LORD be so with you, as I will let you go, and your little ones: look to it; for evil is before you.
EXOD|10|11|Not so: go now ye that are men, and serve the LORD; for that ye did desire. And they were driven out from Pharaoh's presence.
EXOD|10|12|And the LORD said unto Moses, Stretch out thine hand over the land of Egypt for the locusts, that they may come up upon the land of Egypt, and eat every herb of the land, even all that the hail hath left.
EXOD|10|13|And Moses stretched forth his rod over the land of Egypt, and the LORD brought an east wind upon the land all that day, and all that night; and when it was morning, the east wind brought the locusts.
EXOD|10|14|And the locust went up over all the land of Egypt, and rested in all the coasts of Egypt: very grievous were they; before them there were no such locusts as they, neither after them shall be such.
EXOD|10|15|For they covered the face of the whole earth, so that the land was darkened; and they did eat every herb of the land, and all the fruit of the trees which the hail had left: and there remained not any green thing in the trees, or in the herbs of the field, through all the land of Egypt.
EXOD|10|16|Then Pharaoh called for Moses and Aaron in haste; and he said, I have sinned against the LORD your God, and against you.
EXOD|10|17|Now therefore forgive, I pray thee, my sin only this once, and entreat the LORD your God, that he may take away from me this death only.
EXOD|10|18|And he went out from Pharaoh, and entreated the LORD.
EXOD|10|19|And the LORD turned a mighty strong west wind, which took away the locusts, and cast them into the Red sea; there remained not one locust in all the coasts of Egypt.
EXOD|10|20|But the LORD hardened Pharaoh's heart, so that he would not let the children of Israel go.
EXOD|10|21|And the LORD said unto Moses, Stretch out thine hand toward heaven, that there may be darkness over the land of Egypt, even darkness which may be felt.
EXOD|10|22|And Moses stretched forth his hand toward heaven; and there was a thick darkness in all the land of Egypt three days:
EXOD|10|23|They saw not one another, neither rose any from his place for three days: but all the children of Israel had light in their dwellings.
EXOD|10|24|And Pharaoh called unto Moses, and said, Go ye, serve the LORD; only let your flocks and your herds be stayed: let your little ones also go with you.
EXOD|10|25|And Moses said, Thou must give us also sacrifices and burnt offerings, that we may sacrifice unto the LORD our God.
EXOD|10|26|Our cattle also shall go with us; there shall not an hoof be left behind; for thereof must we take to serve the LORD our God; and we know not with what we must serve the LORD, until we come thither.
EXOD|10|27|But the LORD hardened Pharaoh's heart, and he would not let them go.
EXOD|10|28|And Pharaoh said unto him, Get thee from me, take heed to thyself, see my face no more; for in that day thou seest my face thou shalt die.
EXOD|10|29|And Moses said, Thou hast spoken well, I will see thy face again no more.
EXOD|11|1|And the LORD said unto Moses, Yet will I bring one plague more upon Pharaoh, and upon Egypt; afterwards he will let you go hence: when he shall let you go, he shall surely thrust you out hence altogether.
EXOD|11|2|Speak now in the ears of the people, and let every man borrow of his neighbor, and every woman of her neighbor, jewels of silver and jewels of gold.
EXOD|11|3|And the LORD gave the people favor in the sight of the Egyptians. Moreover the man Moses was very great in the land of Egypt, in the sight of Pharaoh's servants, and in the sight of the people.
EXOD|11|4|And Moses said, Thus saith the LORD, About midnight will I go out into the midst of Egypt:
EXOD|11|5|And all the firstborn in the land of Egypt shall die, from the first born of Pharaoh that sitteth upon his throne, even unto the firstborn of the maidservant that is behind the mill; and all the firstborn of beasts.
EXOD|11|6|And there shall be a great cry throughout all the land of Egypt, such as there was none like it, nor shall be like it any more.
EXOD|11|7|But against any of the children of Israel shall not a dog move his tongue, against man or beast: that ye may know how that the LORD doth put a difference between the Egyptians and Israel.
EXOD|11|8|And all these thy servants shall come down unto me, and bow down themselves unto me, saying, Get thee out, and all the people that follow thee: and after that I will go out. And he went out from Pharaoh in a great anger.
EXOD|11|9|And the LORD said unto Moses, Pharaoh shall not hearken unto you; that my wonders may be multiplied in the land of Egypt.
EXOD|11|10|And Moses and Aaron did all these wonders before Pharaoh: and the LORD hardened Pharaoh's heart, so that he would not let the children of Israel go out of his land.
EXOD|12|1|And the LORD spake unto Moses and Aaron in the land of Egypt saying,
EXOD|12|2|This month shall be unto you the beginning of months: it shall be the first month of the year to you.
EXOD|12|3|Speak ye unto all the congregation of Israel, saying, In the tenth day of this month they shall take to them every man a lamb, according to the house of their fathers, a lamb for an house:
EXOD|12|4|And if the household be too little for the lamb, let him and his neighbor next unto his house take it according to the number of the souls; every man according to his eating shall make your count for the lamb.
EXOD|12|5|Your lamb shall be without blemish, a male of the first year: ye shall take it out from the sheep, or from the goats:
EXOD|12|6|And ye shall keep it up until the fourteenth day of the same month: and the whole assembly of the congregation of Israel shall kill it in the evening.
EXOD|12|7|And they shall take of the blood, and strike it on the two side posts and on the upper door post of the houses, wherein they shall eat it.
EXOD|12|8|And they shall eat the flesh in that night, roast with fire, and unleavened bread; and with bitter herbs they shall eat it.
EXOD|12|9|Eat not of it raw, nor sodden at all with water, but roast with fire; his head with his legs, and with the purtenance thereof.
EXOD|12|10|And ye shall let nothing of it remain until the morning; and that which remaineth of it until the morning ye shall burn with fire.
EXOD|12|11|And thus shall ye eat it; with your loins girded, your shoes on your feet, and your staff in your hand; and ye shall eat it in haste: it is the LORD's passover.
EXOD|12|12|For I will pass through the land of Egypt this night, and will smite all the firstborn in the land of Egypt, both man and beast; and against all the gods of Egypt I will execute judgment: I am the LORD.
EXOD|12|13|And the blood shall be to you for a token upon the houses where ye are: and when I see the blood, I will pass over you, and the plague shall not be upon you to destroy you, when I smite the land of Egypt.
EXOD|12|14|And this day shall be unto you for a memorial; and ye shall keep it a feast to the LORD throughout your generations; ye shall keep it a feast by an ordinance for ever.
EXOD|12|15|Seven days shall ye eat unleavened bread; even the first day ye shall put away leaven out of your houses: for whosoever eateth leavened bread from the first day until the seventh day, that soul shall be cut off from Israel.
EXOD|12|16|And in the first day there shall be an holy convocation, and in the seventh day there shall be an holy convocation to you; no manner of work shall be done in them, save that which every man must eat, that only may be done of you.
EXOD|12|17|And ye shall observe the feast of unleavened bread; for in this selfsame day have I brought your armies out of the land of Egypt: therefore shall ye observe this day in your generations by an ordinance for ever.
EXOD|12|18|In the first month, on the fourteenth day of the month at even, ye shall eat unleavened bread, until the one and twentieth day of the month at even.
EXOD|12|19|Seven days shall there be no leaven found in your houses: for whosoever eateth that which is leavened, even that soul shall be cut off from the congregation of Israel, whether he be a stranger, or born in the land.
EXOD|12|20|Ye shall eat nothing leavened; in all your habitations shall ye eat unleavened bread.
EXOD|12|21|Then Moses called for all the elders of Israel, and said unto them, Draw out and take you a lamb according to your families, and kill the passover.
EXOD|12|22|And ye shall take a bunch of hyssop, and dip it in the blood that is in the basin, and strike the lintel and the two side posts with the blood that is in the basin; and none of you shall go out at the door of his house until the morning.
EXOD|12|23|For the LORD will pass through to smite the Egyptians; and when he seeth the blood upon the lintel, and on the two side posts, the LORD will pass over the door, and will not suffer the destroyer to come in unto your houses to smite you.
EXOD|12|24|And ye shall observe this thing for an ordinance to thee and to thy sons for ever.
EXOD|12|25|And it shall come to pass, when ye be come to the land which the LORD will give you, according as he hath promised, that ye shall keep this service.
EXOD|12|26|And it shall come to pass, when your children shall say unto you, What mean ye by this service?
EXOD|12|27|That ye shall say, It is the sacrifice of the LORD's passover, who passed over the houses of the children of Israel in Egypt, when he smote the Egyptians, and delivered our houses. And the people bowed the head and worshipped.
EXOD|12|28|And the children of Israel went away, and did as the LORD had commanded Moses and Aaron, so did they.
EXOD|12|29|And it came to pass, that at midnight the LORD smote all the firstborn in the land of Egypt, from the firstborn of Pharaoh that sat on his throne unto the firstborn of the captive that was in the dungeon; and all the firstborn of cattle.
EXOD|12|30|And Pharaoh rose up in the night, he, and all his servants, and all the Egyptians; and there was a great cry in Egypt; for there was not a house where there was not one dead.
EXOD|12|31|And he called for Moses and Aaron by night, and said, Rise up, and get you forth from among my people, both ye and the children of Israel; and go, serve the LORD, as ye have said.
EXOD|12|32|Also take your flocks and your herds, as ye have said, and be gone; and bless me also.
EXOD|12|33|And the Egyptians were urgent upon the people, that they might send them out of the land in haste; for they said, We be all dead men.
EXOD|12|34|And the people took their dough before it was leavened, their kneadingtroughs being bound up in their clothes upon their shoulders.
EXOD|12|35|And the children of Israel did according to the word of Moses; and they borrowed of the Egyptians jewels of silver, and jewels of gold, and raiment:
EXOD|12|36|And the LORD gave the people favor in the sight of the Egyptians, so that they lent unto them such things as they required. And they spoiled the Egyptians.
EXOD|12|37|And the children of Israel journeyed from Rameses to Succoth, about six hundred thousand on foot that were men, beside children.
EXOD|12|38|And a mixed multitude went up also with them; and flocks, and herds, even very much cattle.
EXOD|12|39|And they baked unleavened cakes of the dough which they brought forth out of Egypt, for it was not leavened; because they were thrust out of Egypt, and could not tarry, neither had they prepared for themselves any victual.
EXOD|12|40|Now the sojourning of the children of Israel, who dwelt in Egypt, was four hundred and thirty years.
EXOD|12|41|And it came to pass at the end of the four hundred and thirty years, even the selfsame day it came to pass, that all the hosts of the LORD went out from the land of Egypt.
EXOD|12|42|It is a night to be much observed unto the LORD for bringing them out from the land of Egypt: this is that night of the LORD to be observed of all the children of Israel in their generations.
EXOD|12|43|And the LORD said unto Moses and Aaron, This is the ordinance of the passover: There shall no stranger eat thereof:
EXOD|12|44|But every man's servant that is bought for money, when thou hast circumcised him, then shall he eat thereof.
EXOD|12|45|A foreigner and an hired servant shall not eat thereof.
EXOD|12|46|In one house shall it be eaten; thou shalt not carry forth ought of the flesh abroad out of the house; neither shall ye break a bone thereof.
EXOD|12|47|All the congregation of Israel shall keep it.
EXOD|12|48|And when a stranger shall sojourn with thee, and will keep the passover to the LORD, let all his males be circumcised, and then let him come near and keep it; and he shall be as one that is born in the land: for no uncircumcised person shall eat thereof.
EXOD|12|49|One law shall be to him that is homeborn, and unto the stranger that sojourneth among you.
EXOD|12|50|Thus did all the children of Israel; as the LORD commanded Moses and Aaron, so did they.
EXOD|12|51|And it came to pass the selfsame day, that the LORD did bring the children of Israel out of the land of Egypt by their armies.
EXOD|13|1|And the LORD spake unto Moses, saying,
EXOD|13|2|Sanctify unto me all the firstborn, whatsoever openeth the womb among the children of Israel, both of man and of beast: it is mine.
EXOD|13|3|And Moses said unto the people, Remember this day, in which ye came out from Egypt, out of the house of bondage; for by strength of hand the LORD brought you out from this place: there shall no leavened bread be eaten.
EXOD|13|4|This day came ye out in the month Abib.
EXOD|13|5|And it shall be when the LORD shall bring thee into the land of the Canaanites, and the Hittites, and the Amorites, and the Hivites, and the Jebusites, which he sware unto thy fathers to give thee, a land flowing with milk and honey, that thou shalt keep this service in this month.
EXOD|13|6|Seven days thou shalt eat unleavened bread, and in the seventh day shall be a feast to the LORD.
EXOD|13|7|Unleavened bread shall be eaten seven days; and there shall no leavened bread be seen with thee, neither shall there be leaven seen with thee in all thy quarters.
EXOD|13|8|And thou shalt show thy son in that day, saying, This is done because of that which the LORD did unto me when I came forth out of Egypt.
EXOD|13|9|And it shall be for a sign unto thee upon thine hand, and for a memorial between thine eyes, that the LORD's law may be in thy mouth: for with a strong hand hath the LORD brought thee out of Egypt.
EXOD|13|10|Thou shalt therefore keep this ordinance in his season from year to year.
EXOD|13|11|And it shall be when the LORD shall bring thee into the land of the Canaanites, as he sware unto thee and to thy fathers, and shall give it thee,
EXOD|13|12|That thou shalt set apart unto the LORD all that openeth the matrix, and every firstling that cometh of a beast which thou hast; the males shall be the LORD's.
EXOD|13|13|And every firstling of an ass thou shalt redeem with a lamb; and if thou wilt not redeem it, then thou shalt break his neck: and all the firstborn of man among thy children shalt thou redeem.
EXOD|13|14|And it shall be when thy son asketh thee in time to come, saying, What is this? that thou shalt say unto him, By strength of hand the LORD brought us out from Egypt, from the house of bondage:
EXOD|13|15|And it came to pass, when Pharaoh would hardly let us go, that the LORD slew all the firstborn in the land of Egypt, both the firstborn of man, and the firstborn of beast: therefore I sacrifice to the LORD all that openeth the matrix, being males; but all the firstborn of my children I redeem.
EXOD|13|16|And it shall be for a token upon thine hand, and for frontlets between thine eyes: for by strength of hand the LORD brought us forth out of Egypt.
EXOD|13|17|And it came to pass, when Pharaoh had let the people go, that God led them not through the way of the land of the Philistines, although that was near; for God said, Lest peradventure the people repent when they see war, and they return to Egypt:
EXOD|13|18|But God led the people about, through the way of the wilderness of the Red sea: and the children of Israel went up harnessed out of the land of Egypt.
EXOD|13|19|And Moses took the bones of Joseph with him: for he had straitly sworn the children of Israel, saying, God will surely visit you; and ye shall carry up my bones away hence with you.
EXOD|13|20|And they took their journey from Succoth, and encamped in Etham, in the edge of the wilderness.
EXOD|13|21|And the LORD went before them by day in a pillar of a cloud, to lead them the way; and by night in a pillar of fire, to give them light; to go by day and night:
EXOD|13|22|He took not away the pillar of the cloud by day, nor the pillar of fire by night, from before the people.
EXOD|14|1|And the LORD spake unto Moses, saying,
EXOD|14|2|Speak unto the children of Israel, that they turn and encamp before Pihahiroth, between Migdol and the sea, over against Baalzephon: before it shall ye encamp by the sea.
EXOD|14|3|For Pharaoh will say of the children of Israel, They are entangled in the land, the wilderness hath shut them in.
EXOD|14|4|And I will harden Pharaoh's heart, that he shall follow after them; and I will be honored upon Pharaoh, and upon all his host; that the Egyptians may know that I am the LORD. And they did so.
EXOD|14|5|And it was told the king of Egypt that the people fled: and the heart of Pharaoh and of his servants was turned against the people, and they said, Why have we done this, that we have let Israel go from serving us?
EXOD|14|6|And he made ready his chariot, and took his people with him:
EXOD|14|7|And he took six hundred chosen chariots, and all the chariots of Egypt, and captains over every one of them.
EXOD|14|8|And the LORD hardened the heart of Pharaoh king of Egypt, and he pursued after the children of Israel: and the children of Israel went out with an high hand.
EXOD|14|9|But the Egyptians pursued after them, all the horses and chariots of Pharaoh, and his horsemen, and his army, and overtook them encamping by the sea, beside Pihahiroth, before Baalzephon.
EXOD|14|10|And when Pharaoh drew nigh, the children of Israel lifted up their eyes, and, behold, the Egyptians marched after them; and they were sore afraid: and the children of Israel cried out unto the LORD.
EXOD|14|11|And they said unto Moses, Because there were no graves in Egypt, hast thou taken us away to die in the wilderness? wherefore hast thou dealt thus with us, to carry us forth out of Egypt?
EXOD|14|12|Is not this the word that we did tell thee in Egypt, saying, Let us alone, that we may serve the Egyptians? For it had been better for us to serve the Egyptians, than that we should die in the wilderness.
EXOD|14|13|And Moses said unto the people, Fear ye not, stand still, and see the salvation of the LORD, which he will show to you to day: for the Egyptians whom ye have seen to day, ye shall see them again no more for ever.
EXOD|14|14|The LORD shall fight for you, and ye shall hold your peace.
EXOD|14|15|And the LORD said unto Moses, Wherefore criest thou unto me? speak unto the children of Israel, that they go forward:
EXOD|14|16|But lift thou up thy rod, and stretch out thine hand over the sea, and divide it: and the children of Israel shall go on dry ground through the midst of the sea.
EXOD|14|17|And I, behold, I will harden the hearts of the Egyptians, and they shall follow them: and I will get me honor upon Pharaoh, and upon all his host, upon his chariots, and upon his horsemen.
EXOD|14|18|And the Egyptians shall know that I am the LORD, when I have gotten me honor upon Pharaoh, upon his chariots, and upon his horsemen.
EXOD|14|19|And the angel of God, which went before the camp of Israel, removed and went behind them; and the pillar of the cloud went from before their face, and stood behind them:
EXOD|14|20|And it came between the camp of the Egyptians and the camp of Israel; and it was a cloud and darkness to them, but it gave light by night to these: so that the one came not near the other all the night.
EXOD|14|21|And Moses stretched out his hand over the sea; and the LORD caused the sea to go back by a strong east wind all that night, and made the sea dry land, and the waters were divided.
EXOD|14|22|And the children of Israel went into the midst of the sea upon the dry ground: and the waters were a wall unto them on their right hand, and on their left.
EXOD|14|23|And the Egyptians pursued, and went in after them to the midst of the sea, even all Pharaoh's horses, his chariots, and his horsemen.
EXOD|14|24|And it came to pass, that in the morning watch the LORD looked unto the host of the Egyptians through the pillar of fire and of the cloud, and troubled the host of the Egyptians,
EXOD|14|25|And took off their chariot wheels, that they drave them heavily: so that the Egyptians said, Let us flee from the face of Israel; for the LORD fighteth for them against the Egyptians.
EXOD|14|26|And the LORD said unto Moses, Stretch out thine hand over the sea, that the waters may come again upon the Egyptians, upon their chariots, and upon their horsemen.
EXOD|14|27|And Moses stretched forth his hand over the sea, and the sea returned to his strength when the morning appeared; and the Egyptians fled against it; and the LORD overthrew the Egyptians in the midst of the sea.
EXOD|14|28|And the waters returned, and covered the chariots, and the horsemen, and all the host of Pharaoh that came into the sea after them; there remained not so much as one of them.
EXOD|14|29|But the children of Israel walked upon dry land in the midst of the sea; and the waters were a wall unto them on their right hand, and on their left.
EXOD|14|30|Thus the LORD saved Israel that day out of the hand of the Egyptians; and Israel saw the Egyptians dead upon the sea shore.
EXOD|14|31|And Israel saw that great work which the LORD did upon the Egyptians: and the people feared the LORD, and believed the LORD, and his servant Moses.
EXOD|15|1|Then sang Moses and the children of Israel this song unto the LORD, and spake, saying, I will sing unto the LORD, for he hath triumphed gloriously: the horse and his rider hath he thrown into the sea.
EXOD|15|2|The LORD is my strength and song, and he is become my salvation: he is my God, and I will prepare him an habitation; my father's God, and I will exalt him.
EXOD|15|3|The LORD is a man of war: the LORD is his name.
EXOD|15|4|Pharaoh's chariots and his host hath he cast into the sea: his chosen captains also are drowned in the Red sea.
EXOD|15|5|The depths have covered them: they sank into the bottom as a stone.
EXOD|15|6|Thy right hand, O LORD, is become glorious in power: thy right hand, O LORD, hath dashed in pieces the enemy.
EXOD|15|7|And in the greatness of thine excellency thou hast overthrown them that rose up against thee: thou sentest forth thy wrath, which consumed them as stubble.
EXOD|15|8|And with the blast of thy nostrils the waters were gathered together, the floods stood upright as an heap, and the depths were congealed in the heart of the sea.
EXOD|15|9|The enemy said, I will pursue, I will overtake, I will divide the spoil; my lust shall be satisfied upon them; I will draw my sword, my hand shall destroy them.
EXOD|15|10|Thou didst blow with thy wind, the sea covered them: they sank as lead in the mighty waters.
EXOD|15|11|Who is like unto thee, O LORD, among the gods? who is like thee, glorious in holiness, fearful in praises, doing wonders?
EXOD|15|12|Thou stretchedst out thy right hand, the earth swallowed them.
EXOD|15|13|Thou in thy mercy hast led forth the people which thou hast redeemed: thou hast guided them in thy strength unto thy holy habitation.
EXOD|15|14|The people shall hear, and be afraid: sorrow shall take hold on the inhabitants of Palestina.
EXOD|15|15|Then the dukes of Edom shall be amazed; the mighty men of Moab, trembling shall take hold upon them; all the inhabitants of Canaan shall melt away.
EXOD|15|16|Fear and dread shall fall upon them; by the greatness of thine arm they shall be as still as a stone; till thy people pass over, O LORD, till the people pass over, which thou hast purchased.
EXOD|15|17|Thou shalt bring them in, and plant them in the mountain of thine inheritance, in the place, O LORD, which thou hast made for thee to dwell in, in the Sanctuary, O LORD, which thy hands have established.
EXOD|15|18|The LORD shall reign for ever and ever.
EXOD|15|19|For the horse of Pharaoh went in with his chariots and with his horsemen into the sea, and the LORD brought again the waters of the sea upon them; but the children of Israel went on dry land in the midst of the sea.
EXOD|15|20|And Miriam the prophetess, the sister of Aaron, took a timbrel in her hand; and all the women went out after her with timbrels and with dances.
EXOD|15|21|And Miriam answered them, Sing ye to the LORD, for he hath triumphed gloriously; the horse and his rider hath he thrown into the sea.
EXOD|15|22|So Moses brought Israel from the Red sea, and they went out into the wilderness of Shur; and they went three days in the wilderness, and found no water.
EXOD|15|23|And when they came to Marah, they could not drink of the waters of Marah, for they were bitter: therefore the name of it was called Marah.
EXOD|15|24|And the people murmured against Moses, saying, What shall we drink?
EXOD|15|25|And he cried unto the LORD; and the LORD showed him a tree, which when he had cast into the waters, the waters were made sweet: there he made for them a statute and an ordinance, and there he proved them,
EXOD|15|26|And said, If thou wilt diligently hearken to the voice of the LORD thy God, and wilt do that which is right in his sight, and wilt give ear to his commandments, and keep all his statutes, I will put none of these diseases upon thee, which I have brought upon the Egyptians: for I am the LORD that healeth thee.
EXOD|15|27|And they came to Elim, where were twelve wells of water, and threescore and ten palm trees: and they encamped there by the waters.
EXOD|16|1|And they took their journey from Elim, and all the congregation of the children of Israel came unto the wilderness of Sin, which is between Elim and Sinai, on the fifteenth day of the second month after their departing out of the land of Egypt.
EXOD|16|2|And the whole congregation of the children of Israel murmured against Moses and Aaron in the wilderness:
EXOD|16|3|And the children of Israel said unto them, Would to God we had died by the hand of the LORD in the land of Egypt, when we sat by the flesh pots, and when we did eat bread to the full; for ye have brought us forth into this wilderness, to kill this whole assembly with hunger.
EXOD|16|4|Then said the LORD unto Moses, Behold, I will rain bread from heaven for you; and the people shall go out and gather a certain rate every day, that I may prove them, whether they will walk in my law, or no.
EXOD|16|5|And it shall come to pass, that on the sixth day they shall prepare that which they bring in; and it shall be twice as much as they gather daily.
EXOD|16|6|And Moses and Aaron said unto all the children of Israel, At even, then ye shall know that the LORD hath brought you out from the land of Egypt:
EXOD|16|7|And in the morning, then ye shall see the glory of the LORD; for that he heareth your murmurings against the LORD: and what are we, that ye murmur against us?
EXOD|16|8|And Moses said, This shall be, when the LORD shall give you in the evening flesh to eat, and in the morning bread to the full; for that the LORD heareth your murmurings which ye murmur against him: and what are we? your murmurings are not against us, but against the LORD.
EXOD|16|9|And Moses spake unto Aaron, Say unto all the congregation of the children of Israel, Come near before the LORD: for he hath heard your murmurings.
EXOD|16|10|And it came to pass, as Aaron spake unto the whole congregation of the children of Israel, that they looked toward the wilderness, and, behold, the glory of the LORD appeared in the cloud.
EXOD|16|11|And the LORD spake unto Moses, saying,
EXOD|16|12|I have heard the murmurings of the children of Israel: speak unto them, saying, At even ye shall eat flesh, and in the morning ye shall be filled with bread; and ye shall know that I am the LORD your God.
EXOD|16|13|And it came to pass, that at even the quails came up, and covered the camp: and in the morning the dew lay round about the host.
EXOD|16|14|And when the dew that lay was gone up, behold, upon the face of the wilderness there lay a small round thing, as small as the hoar frost on the ground.
EXOD|16|15|And when the children of Israel saw it, they said one to another, It is manna: for they wist not what it was. And Moses said unto them, This is the bread which the LORD hath given you to eat.
EXOD|16|16|This is the thing which the LORD hath commanded, Gather of it every man according to his eating, an omer for every man, according to the number of your persons; take ye every man for them which are in his tents.
EXOD|16|17|And the children of Israel did so, and gathered, some more, some less.
EXOD|16|18|And when they did mete it with an omer, he that gathered much had nothing over, and he that gathered little had no lack; they gathered every man according to his eating.
EXOD|16|19|And Moses said, Let no man leave of it till the morning.
EXOD|16|20|Notwithstanding they hearkened not unto Moses; but some of them left of it until the morning, and it bred worms, and stank: and Moses was wroth with them.
EXOD|16|21|And they gathered it every morning, every man according to his eating: and when the sun waxed hot, it melted.
EXOD|16|22|And it came to pass, that on the sixth day they gathered twice as much bread, two omers for one man: and all the rulers of the congregation came and told Moses.
EXOD|16|23|And he said unto them, This is that which the LORD hath said, To morrow is the rest of the holy sabbath unto the LORD: bake that which ye will bake to day, and seethe that ye will seethe; and that which remaineth over lay up for you to be kept until the morning.
EXOD|16|24|And they laid it up till the morning, as Moses bade: and it did not stink, neither was there any worm therein.
EXOD|16|25|And Moses said, Eat that to day; for to day is a sabbath unto the LORD: to day ye shall not find it in the field.
EXOD|16|26|Six days ye shall gather it; but on the seventh day, which is the sabbath, in it there shall be none.
EXOD|16|27|And it came to pass, that there went out some of the people on the seventh day for to gather, and they found none.
EXOD|16|28|And the LORD said unto Moses, How long refuse ye to keep my commandments and my laws?
EXOD|16|29|See, for that the LORD hath given you the sabbath, therefore he giveth you on the sixth day the bread of two days; abide ye every man in his place, let no man go out of his place on the seventh day.
EXOD|16|30|So the people rested on the seventh day.
EXOD|16|31|And the house of Israel called the name thereof Manna: and it was like coriander seed, white; and the taste of it was like wafers made with honey.
EXOD|16|32|And Moses said, This is the thing which the LORD commandeth, Fill an omer of it to be kept for your generations; that they may see the bread wherewith I have fed you in the wilderness, when I brought you forth from the land of Egypt.
EXOD|16|33|And Moses said unto Aaron, Take a pot, and put an omer full of manna therein, and lay it up before the LORD, to be kept for your generations.
EXOD|16|34|As the LORD commanded Moses, so Aaron laid it up before the Testimony, to be kept.
EXOD|16|35|And the children of Israel did eat manna forty years, until they came to a land inhabited; they did eat manna, until they came unto the borders of the land of Canaan.
EXOD|16|36|Now an omer is the tenth part of an ephah.
EXOD|17|1|And all the congregation of the children of Israel journeyed from the wilderness of Sin, after their journeys, according to the commandment of the LORD, and pitched in Rephidim: and there was no water for the people to drink.
EXOD|17|2|Wherefore the people did chide with Moses, and said, Give us water that we may drink. And Moses said unto them, Why chide ye with me? wherefore do ye tempt the LORD?
EXOD|17|3|And the people thirsted there for water; and the people murmured against Moses, and said, Wherefore is this that thou hast brought us up out of Egypt, to kill us and our children and our cattle with thirst?
EXOD|17|4|And Moses cried unto the LORD, saying, What shall I do unto this people? they be almost ready to stone me.
EXOD|17|5|And the LORD said unto Moses, Go on before the people, and take with thee of the elders of Israel; and thy rod, wherewith thou smotest the river, take in thine hand, and go.
EXOD|17|6|Behold, I will stand before thee there upon the rock in Horeb; and thou shalt smite the rock, and there shall come water out of it, that the people may drink. And Moses did so in the sight of the elders of Israel.
EXOD|17|7|And he called the name of the place Massah, and Meribah, because of the chiding of the children of Israel, and because they tempted the LORD, saying, Is the LORD among us, or not?
EXOD|17|8|Then came Amalek, and fought with Israel in Rephidim.
EXOD|17|9|And Moses said unto Joshua, Choose us out men, and go out, fight with Amalek: to morrow I will stand on the top of the hill with the rod of God in mine hand.
EXOD|17|10|So Joshua did as Moses had said to him, and fought with Amalek: and Moses, Aaron, and Hur went up to the top of the hill.
EXOD|17|11|And it came to pass, when Moses held up his hand, that Israel prevailed: and when he let down his hand, Amalek prevailed.
EXOD|17|12|But Moses hands were heavy; and they took a stone, and put it under him, and he sat thereon; and Aaron and Hur stayed up his hands, the one on the one side, and the other on the other side; and his hands were steady until the going down of the sun.
EXOD|17|13|And Joshua discomfited Amalek and his people with the edge of the sword.
EXOD|17|14|And the LORD said unto Moses, Write this for a memorial in a book, and rehearse it in the ears of Joshua: for I will utterly put out the remembrance of Amalek from under heaven.
EXOD|17|15|And Moses built an altar, and called the name of it Jehovahnissi:
EXOD|17|16|For he said, Because the LORD hath sworn that the LORD will have war with Amalek from generation to generation.
EXOD|18|1|When Jethro, the priest of Midian, Moses' father in law, heard of all that God had done for Moses, and for Israel his people, and that the LORD had brought Israel out of Egypt;
EXOD|18|2|Then Jethro, Moses' father in law, took Zipporah, Moses' wife, after he had sent her back,
EXOD|18|3|And her two sons; of which the name of the one was Gershom; for he said, I have been an alien in a strange land:
EXOD|18|4|And the name of the other was Eliezer; for the God of my father, said he, was mine help, and delivered me from the sword of Pharaoh:
EXOD|18|5|And Jethro, Moses' father in law, came with his sons and his wife unto Moses into the wilderness, where he encamped at the mount of God:
EXOD|18|6|And he said unto Moses, I thy father in law Jethro am come unto thee, and thy wife, and her two sons with her.
EXOD|18|7|And Moses went out to meet his father in law, and did obeisance, and kissed him; and they asked each other of their welfare; and they came into the tent.
EXOD|18|8|And Moses told his father in law all that the LORD had done unto Pharaoh and to the Egyptians for Israel's sake, and all the travail that had come upon them by the way, and how the LORD delivered them.
EXOD|18|9|And Jethro rejoiced for all the goodness which the LORD had done to Israel, whom he had delivered out of the hand of the Egyptians.
EXOD|18|10|And Jethro said, Blessed be the LORD, who hath delivered you out of the hand of the Egyptians, and out of the hand of Pharaoh, who hath delivered the people from under the hand of the Egyptians.
EXOD|18|11|Now I know that the LORD is greater than all gods: for in the thing wherein they dealt proudly he was above them.
EXOD|18|12|And Jethro, Moses' father in law, took a burnt offering and sacrifices for God: and Aaron came, and all the elders of Israel, to eat bread with Moses' father in law before God.
EXOD|18|13|And it came to pass on the morrow, that Moses sat to judge the people: and the people stood by Moses from the morning unto the evening.
EXOD|18|14|And when Moses' father in law saw all that he did to the people, he said, What is this thing that thou doest to the people? why sittest thou thyself alone, and all the people stand by thee from morning unto even?
EXOD|18|15|And Moses said unto his father in law, Because the people come unto me to inquire of God:
EXOD|18|16|When they have a matter, they come unto me; and I judge between one and another, and I do make them know the statutes of God, and his laws.
EXOD|18|17|And Moses' father in law said unto him, The thing that thou doest is not good.
EXOD|18|18|Thou wilt surely wear away, both thou, and this people that is with thee: for this thing is too heavy for thee; thou art not able to perform it thyself alone.
EXOD|18|19|Hearken now unto my voice, I will give thee counsel, and God shall be with thee: Be thou for the people to God-ward, that thou mayest bring the causes unto God:
EXOD|18|20|And thou shalt teach them ordinances and laws, and shalt show them the way wherein they must walk, and the work that they must do.
EXOD|18|21|Moreover thou shalt provide out of all the people able men, such as fear God, men of truth, hating covetousness; and place such over them, to be rulers of thousands, and rulers of hundreds, rulers of fifties, and rulers of tens:
EXOD|18|22|And let them judge the people at all seasons: and it shall be, that every great matter they shall bring unto thee, but every small matter they shall judge: so shall it be easier for thyself, and they shall bear the burden with thee.
EXOD|18|23|If thou shalt do this thing, and God command thee so, then thou shalt be able to endure, and all this people shall also go to their place in peace.
EXOD|18|24|So Moses hearkened to the voice of his father in law, and did all that he had said.
EXOD|18|25|And Moses chose able men out of all Israel, and made them heads over the people, rulers of thousands, rulers of hundreds, rulers of fifties, and rulers of tens.
EXOD|18|26|And they judged the people at all seasons: the hard causes they brought unto Moses, but every small matter they judged themselves.
EXOD|18|27|And Moses let his father in law depart; and he went his way into his own land.
EXOD|19|1|In the third month, when the children of Israel were gone forth out of the land of Egypt, the same day came they into the wilderness of Sinai.
EXOD|19|2|For they were departed from Rephidim, and were come to the desert of Sinai, and had pitched in the wilderness; and there Israel camped before the mount.
EXOD|19|3|And Moses went up unto God, and the LORD called unto him out of the mountain, saying, Thus shalt thou say to the house of Jacob, and tell the children of Israel;
EXOD|19|4|Ye have seen what I did unto the Egyptians, and how I bare you on eagles' wings, and brought you unto myself.
EXOD|19|5|Now therefore, if ye will obey my voice indeed, and keep my covenant, then ye shall be a peculiar treasure unto me above all people: for all the earth is mine:
EXOD|19|6|And ye shall be unto me a kingdom of priests, and an holy nation. These are the words which thou shalt speak unto the children of Israel.
EXOD|19|7|And Moses came and called for the elders of the people, and laid before their faces all these words which the LORD commanded him.
EXOD|19|8|And all the people answered together, and said, All that the LORD hath spoken we will do. And Moses returned the words of the people unto the LORD.
EXOD|19|9|And the LORD said unto Moses, Lo, I come unto thee in a thick cloud, that the people may hear when I speak with thee, and believe thee for ever. And Moses told the words of the people unto the LORD.
EXOD|19|10|And the LORD said unto Moses, Go unto the people, and sanctify them to day and to morrow, and let them wash their clothes,
EXOD|19|11|And be ready against the third day: for the third day the LORD will come down in the sight of all the people upon mount Sinai.
EXOD|19|12|And thou shalt set bounds unto the people round about, saying, Take heed to yourselves, that ye go not up into the mount, or touch the border of it: whosoever toucheth the mount shall be surely put to death:
EXOD|19|13|There shall not an hand touch it, but he shall surely be stoned, or shot through; whether it be beast or man, it shall not live: when the trumpet soundeth long, they shall come up to the mount.
EXOD|19|14|And Moses went down from the mount unto the people, and sanctified the people; and they washed their clothes.
EXOD|19|15|And he said unto the people, Be ready against the third day: come not at your wives.
EXOD|19|16|And it came to pass on the third day in the morning, that there were thunders and lightnings, and a thick cloud upon the mount, and the voice of the trumpet exceeding loud; so that all the people that was in the camp trembled.
EXOD|19|17|And Moses brought forth the people out of the camp to meet with God; and they stood at the nether part of the mount.
EXOD|19|18|And mount Sinai was altogether on a smoke, because the LORD descended upon it in fire: and the smoke thereof ascended as the smoke of a furnace, and the whole mount quaked greatly.
EXOD|19|19|And when the voice of the trumpet sounded long, and waxed louder and louder, Moses spake, and God answered him by a voice.
EXOD|19|20|And the LORD came down upon mount Sinai, on the top of the mount: and the LORD called Moses up to the top of the mount; and Moses went up.
EXOD|19|21|And the LORD said unto Moses, Go down, charge the people, lest they break through unto the LORD to gaze, and many of them perish.
EXOD|19|22|And let the priests also, which come near to the LORD, sanctify themselves, lest the LORD break forth upon them.
EXOD|19|23|And Moses said unto the LORD, The people cannot come up to mount Sinai: for thou chargedst us, saying, Set bounds about the mount, and sanctify it.
EXOD|19|24|And the LORD said unto him, Away, get thee down, and thou shalt come up, thou, and Aaron with thee: but let not the priests and the people break through to come up unto the LORD, lest he break forth upon them.
EXOD|19|25|So Moses went down unto the people, and spake unto them.
EXOD|20|1|And God spake all these words, saying,
EXOD|20|2|I am the LORD thy God, which have brought thee out of the land of Egypt, out of the house of bondage.
EXOD|20|3|Thou shalt have no other gods before me.
EXOD|20|4|Thou shalt not make unto thee any graven image, or any likeness of any thing that is in heaven above, or that is in the earth beneath, or that is in the water under the earth.
EXOD|20|5|Thou shalt not bow down thyself to them, nor serve them: for I the LORD thy God am a jealous God, visiting the iniquity of the fathers upon the children unto the third and fourth generation of them that hate me;
EXOD|20|6|And showing mercy unto thousands of them that love me, and keep my commandments.
EXOD|20|7|Thou shalt not take the name of the LORD thy God in vain; for the LORD will not hold him guiltless that taketh his name in vain.
EXOD|20|8|Remember the sabbath day, to keep it holy.
EXOD|20|9|Six days shalt thou labor, and do all thy work:
EXOD|20|10|But the seventh day is the sabbath of the LORD thy God: in it thou shalt not do any work, thou, nor thy son, nor thy daughter, thy manservant, nor thy maidservant, nor thy cattle, nor thy stranger that is within thy gates:
EXOD|20|11|For in six days the LORD made heaven and earth, the sea, and all that in them is, and rested the seventh day: wherefore the LORD blessed the sabbath day, and hallowed it.
EXOD|20|12|Honor thy father and thy mother: that thy days may be long upon the land which the LORD thy God giveth thee.
EXOD|20|13|Thou shalt not kill.
EXOD|20|14|Thou shalt not commit adultery.
EXOD|20|15|Thou shalt not steal.
EXOD|20|16|Thou shalt not bear false witness against thy neighbor.
EXOD|20|17|Thou shalt not covet thy neighbor's house, thou shalt not covet thy neighbor's wife, nor his manservant, nor his maidservant, nor his ox, nor his ass, nor any thing that is thy neighbor's.
EXOD|20|18|And all the people saw the thunderings, and the lightnings, and the noise of the trumpet, and the mountain smoking: and when the people saw it, they removed, and stood afar off.
EXOD|20|19|And they said unto Moses, Speak thou with us, and we will hear: but let not God speak with us, lest we die.
EXOD|20|20|And Moses said unto the people, Fear not: for God is come to prove you, and that his fear may be before your faces, that ye sin not.
EXOD|20|21|And the people stood afar off, and Moses drew near unto the thick darkness where God was.
EXOD|20|22|And the LORD said unto Moses, Thus thou shalt say unto the children of Israel, Ye have seen that I have talked with you from heaven.
EXOD|20|23|Ye shall not make with me gods of silver, neither shall ye make unto you gods of gold.
EXOD|20|24|An altar of earth thou shalt make unto me, and shalt sacrifice thereon thy burnt offerings, and thy peace offerings, thy sheep, and thine oxen: in all places where I record my name I will come unto thee, and I will bless thee.
EXOD|20|25|And if thou wilt make me an altar of stone, thou shalt not build it of hewn stone: for if thou lift up thy tool upon it, thou hast polluted it.
EXOD|20|26|Neither shalt thou go up by steps unto mine altar, that thy nakedness be not discovered thereon.
EXOD|21|1|Now these are the judgments which thou shalt set before them.
EXOD|21|2|If thou buy an Hebrew servant, six years he shall serve: and in the seventh he shall go out free for nothing.
EXOD|21|3|If he came in by himself, he shall go out by himself: if he were married, then his wife shall go out with him.
EXOD|21|4|If his master have given him a wife, and she have born him sons or daughters; the wife and her children shall be her master's, and he shall go out by himself.
EXOD|21|5|And if the servant shall plainly say, I love my master, my wife, and my children; I will not go out free:
EXOD|21|6|Then his master shall bring him unto the judges; he shall also bring him to the door, or unto the door post; and his master shall bore his ear through with an awl; and he shall serve him for ever.
EXOD|21|7|And if a man sell his daughter to be a maidservant, she shall not go out as the menservants do.
EXOD|21|8|If she please not her master, who hath betrothed her to himself, then shall he let her be redeemed: to sell her unto a strange nation he shall have no power, seeing he hath dealt deceitfully with her.
EXOD|21|9|And if he have betrothed her unto his son, he shall deal with her after the manner of daughters.
EXOD|21|10|If he take him another wife; her food, her raiment, and her duty of marriage, shall he not diminish.
EXOD|21|11|And if he do not these three unto her, then shall she go out free without money.
EXOD|21|12|He that smiteth a man, so that he die, shall be surely put to death.
EXOD|21|13|And if a man lie not in wait, but God deliver him into his hand; then I will appoint thee a place whither he shall flee.
EXOD|21|14|But if a man come presumptuously upon his neighbor, to slay him with guile; thou shalt take him from mine altar, that he may die.
EXOD|21|15|And he that smiteth his father, or his mother, shall be surely put to death.
EXOD|21|16|And he that stealeth a man, and selleth him, or if he be found in his hand, he shall surely be put to death.
EXOD|21|17|And he that curseth his father, or his mother, shall surely be put to death.
EXOD|21|18|And if men strive together, and one smite another with a stone, or with his fist, and he die not, but keepeth his bed:
EXOD|21|19|If he rise again, and walk abroad upon his staff, then shall he that smote him be quit: only he shall pay for the loss of his time, and shall cause him to be thoroughly healed.
EXOD|21|20|And if a man smite his servant, or his maid, with a rod, and he die under his hand; he shall be surely punished.
EXOD|21|21|Notwithstanding, if he continue a day or two, he shall not be punished: for he is his money.
EXOD|21|22|If men strive, and hurt a woman with child, so that her fruit depart from her, and yet no mischief follow: he shall be surely punished, according as the woman's husband will lay upon him; and he shall pay as the judges determine.
EXOD|21|23|And if any mischief follow, then thou shalt give life for life,
EXOD|21|24|Eye for eye, tooth for tooth, hand for hand, foot for foot,
EXOD|21|25|Burning for burning, wound for wound, stripe for stripe.
EXOD|21|26|And if a man smite the eye of his servant, or the eye of his maid, that it perish; he shall let him go free for his eye's sake.
EXOD|21|27|And if he smite out his manservant's tooth, or his maidservant's tooth; he shall let him go free for his tooth's sake.
EXOD|21|28|If an ox gore a man or a woman, that they die: then the ox shall be surely stoned, and his flesh shall not be eaten; but the owner of the ox shall be quit.
EXOD|21|29|But if the ox were wont to push with his horn in time past, and it hath been testified to his owner, and he hath not kept him in, but that he hath killed a man or a woman; the ox shall be stoned, and his owner also shall be put to death.
EXOD|21|30|If there be laid on him a sum of money, then he shall give for the ransom of his life whatsoever is laid upon him.
EXOD|21|31|Whether he have gored a son, or have gored a daughter, according to this judgment shall it be done unto him.
EXOD|21|32|If the ox shall push a manservant or a maidservant; he shall give unto their master thirty shekels of silver, and the ox shall be stoned.
EXOD|21|33|And if a man shall open a pit, or if a man shall dig a pit, and not cover it, and an ox or an ass fall therein;
EXOD|21|34|The owner of the pit shall make it good, and give money unto the owner of them; and the dead beast shall be his.
EXOD|21|35|And if one man's ox hurt another's, that he die; then they shall sell the live ox, and divide the money of it; and the dead ox also they shall divide.
EXOD|21|36|Or if it be known that the ox hath used to push in time past, and his owner hath not kept him in; he shall surely pay ox for ox; and the dead shall be his own.
EXOD|22|1|If a man shall steal an ox, or a sheep, and kill it, or sell it; he shall restore five oxen for an ox, and four sheep for a sheep.
EXOD|22|2|If a thief be found breaking up, and be smitten that he die, there shall no blood be shed for him.
EXOD|22|3|If the sun be risen upon him, there shall be blood shed for him; for he should make full restitution; if he have nothing, then he shall be sold for his theft.
EXOD|22|4|If the theft be certainly found in his hand alive, whether it be ox, or ass, or sheep; he shall restore double.
EXOD|22|5|If a man shall cause a field or vineyard to be eaten, and shall put in his beast, and shall feed in another man's field; of the best of his own field, and of the best of his own vineyard, shall he make restitution.
EXOD|22|6|If fire break out, and catch in thorns, so that the stacks of corn, or the standing corn, or the field, be consumed therewith; he that kindled the fire shall surely make restitution.
EXOD|22|7|If a man shall deliver unto his neighbor money or stuff to keep, and it be stolen out of the man's house; if the thief be found, let him pay double.
EXOD|22|8|If the thief be not found, then the master of the house shall be brought unto the judges, to see whether he have put his hand unto his neighbor's goods.
EXOD|22|9|For all manner of trespass, whether it be for ox, for ass, for sheep, for raiment, or for any manner of lost thing which another challengeth to be his, the cause of both parties shall come before the judges; and whom the judges shall condemn, he shall pay double unto his neighbor.
EXOD|22|10|If a man deliver unto his neighbor an ass, or an ox, or a sheep, or any beast, to keep; and it die, or be hurt, or driven away, no man seeing it:
EXOD|22|11|Then shall an oath of the LORD be between them both, that he hath not put his hand unto his neighbor's goods; and the owner of it shall accept thereof, and he shall not make it good.
EXOD|22|12|And if it be stolen from him, he shall make restitution unto the owner thereof.
EXOD|22|13|If it be torn in pieces, then let him bring it for witness, and he shall not make good that which was torn.
EXOD|22|14|And if a man borrow ought of his neighbor, and it be hurt, or die, the owner thereof being not with it, he shall surely make it good.
EXOD|22|15|But if the owner thereof be with it, he shall not make it good: if it be an hired thing, it came for his hire.
EXOD|22|16|And if a man entice a maid that is not betrothed, and lie with her, he shall surely endow her to be his wife.
EXOD|22|17|If her father utterly refuse to give her unto him, he shall pay money according to the dowry of virgins.
EXOD|22|18|Thou shalt not suffer a witch to live.
EXOD|22|19|Whosoever lieth with a beast shall surely be put to death.
EXOD|22|20|He that sacrificeth unto any god, save unto the LORD only, he shall be utterly destroyed.
EXOD|22|21|Thou shalt neither vex a stranger, nor oppress him: for ye were strangers in the land of Egypt.
EXOD|22|22|Ye shall not afflict any widow, or fatherless child.
EXOD|22|23|If thou afflict them in any wise, and they cry at all unto me, I will surely hear their cry;
EXOD|22|24|And my wrath shall wax hot, and I will kill you with the sword; and your wives shall be widows, and your children fatherless.
EXOD|22|25|If thou lend money to any of my people that is poor by thee, thou shalt not be to him as an usurer, neither shalt thou lay upon him usury.
EXOD|22|26|If thou at all take thy neighbor's raiment to pledge, thou shalt deliver it unto him by that the sun goeth down:
EXOD|22|27|For that is his covering only, it is his raiment for his skin: wherein shall he sleep? and it shall come to pass, when he crieth unto me, that I will hear; for I am gracious.
EXOD|22|28|Thou shalt not revile the gods, nor curse the ruler of thy people.
EXOD|22|29|Thou shalt not delay to offer the first of thy ripe fruits, and of thy liquors: the firstborn of thy sons shalt thou give unto me.
EXOD|22|30|Likewise shalt thou do with thine oxen, and with thy sheep: seven days it shall be with his dam; on the eighth day thou shalt give it me.
EXOD|22|31|And ye shall be holy men unto me: neither shall ye eat any flesh that is torn of beasts in the field; ye shall cast it to the dogs.
EXOD|23|1|Thou shalt not raise a false report: put not thine hand with the wicked to be an unrighteous witness.
EXOD|23|2|Thou shalt not follow a multitude to do evil; neither shalt thou speak in a cause to decline after many to wrest judgment:
EXOD|23|3|Neither shalt thou countenance a poor man in his cause.
EXOD|23|4|If thou meet thine enemy's ox or his ass going astray, thou shalt surely bring it back to him again.
EXOD|23|5|If thou see the ass of him that hateth thee lying under his burden, and wouldest forbear to help him, thou shalt surely help with him.
EXOD|23|6|Thou shalt not wrest the judgment of thy poor in his cause.
EXOD|23|7|Keep thee far from a false matter; and the innocent and righteous slay thou not: for I will not justify the wicked.
EXOD|23|8|And thou shalt take no gift: for the gift blindeth the wise, and perverteth the words of the righteous.
EXOD|23|9|Also thou shalt not oppress a stranger: for ye know the heart of a stranger, seeing ye were strangers in the land of Egypt.
EXOD|23|10|And six years thou shalt sow thy land, and shalt gather in the fruits thereof:
EXOD|23|11|But the seventh year thou shalt let it rest and lie still; that the poor of thy people may eat: and what they leave the beasts of the field shall eat. In like manner thou shalt deal with thy vineyard, and with thy oliveyard.
EXOD|23|12|Six days thou shalt do thy work, and on the seventh day thou shalt rest: that thine ox and thine ass may rest, and the son of thy handmaid, and the stranger, may be refreshed.
EXOD|23|13|And in all things that I have said unto you be circumspect: and make no mention of the name of other gods, neither let it be heard out of thy mouth.
EXOD|23|14|Three times thou shalt keep a feast unto me in the year.
EXOD|23|15|Thou shalt keep the feast of unleavened bread: (thou shalt eat unleavened bread seven days, as I commanded thee, in the time appointed of the month Abib; for in it thou camest out from Egypt: and none shall appear before me empty:)
EXOD|23|16|And the feast of harvest, the firstfruits of thy labors, which thou hast sown in the field: and the feast of ingathering, which is in the end of the year, when thou hast gathered in thy labors out of the field.
EXOD|23|17|Three items in the year all thy males shall appear before the LORD God.
EXOD|23|18|Thou shalt not offer the blood of my sacrifice with leavened bread; neither shall the fat of my sacrifice remain until the morning.
EXOD|23|19|The first of the firstfruits of thy land thou shalt bring into the house of the LORD thy God. Thou shalt not seethe a kid in his mother's milk.
EXOD|23|20|Behold, I send an Angel before thee, to keep thee in the way, and to bring thee into the place which I have prepared.
EXOD|23|21|Beware of him, and obey his voice, provoke him not; for he will not pardon your transgressions: for my name is in him.
EXOD|23|22|But if thou shalt indeed obey his voice, and do all that I speak; then I will be an enemy unto thine enemies, and an adversary unto thine adversaries.
EXOD|23|23|For mine Angel shall go before thee, and bring thee in unto the Amorites, and the Hittites, and the Perizzites, and the Canaanites, the Hivites, and the Jebusites: and I will cut them off.
EXOD|23|24|Thou shalt not bow down to their gods, nor serve them, nor do after their works: but thou shalt utterly overthrow them, and quite break down their images.
EXOD|23|25|And ye shall serve the LORD your God, and he shall bless thy bread, and thy water; and I will take sickness away from the midst of thee.
EXOD|23|26|There shall nothing cast their young, nor be barren, in thy land: the number of thy days I will fulfil.
EXOD|23|27|I will send my fear before thee, and will destroy all the people to whom thou shalt come, and I will make all thine enemies turn their backs unto thee.
EXOD|23|28|And I will send hornets before thee, which shall drive out the Hivite, the Canaanite, and the Hittite, from before thee.
EXOD|23|29|I will not drive them out from before thee in one year; lest the land become desolate, and the beast of the field multiply against thee.
EXOD|23|30|By little and little I will drive them out from before thee, until thou be increased, and inherit the land.
EXOD|23|31|And I will set thy bounds from the Red sea even unto the sea of the Philistines, and from the desert unto the river: for I will deliver the inhabitants of the land into your hand; and thou shalt drive them out before thee.
EXOD|23|32|Thou shalt make no covenant with them, nor with their gods.
EXOD|23|33|They shall not dwell in thy land, lest they make thee sin against me: for if thou serve their gods, it will surely be a snare unto thee.
EXOD|24|1|And he said unto Moses, Come up unto the LORD, thou, and Aaron, Nadab, and Abihu, and seventy of the elders of Israel; and worship ye afar off.
EXOD|24|2|And Moses alone shall come near the LORD: but they shall not come nigh; neither shall the people go up with him.
EXOD|24|3|And Moses came and told the people all the words of the LORD, and all the judgments: and all the people answered with one voice, and said, All the words which the LORD hath said will we do.
EXOD|24|4|And Moses wrote all the words of the LORD, and rose up early in the morning, and builded an altar under the hill, and twelve pillars, according to the twelve tribes of Israel.
EXOD|24|5|And he sent young men of the children of Israel, which offered burnt offerings, and sacrificed peace offerings of oxen unto the LORD.
EXOD|24|6|And Moses took half of the blood, and put it in basins; and half of the blood he sprinkled on the altar.
EXOD|24|7|And he took the book of the covenant, and read in the audience of the people: and they said, All that the LORD hath said will we do, and be obedient.
EXOD|24|8|And Moses took the blood, and sprinkled it on the people, and said, Behold the blood of the covenant, which the LORD hath made with you concerning all these words.
EXOD|24|9|Then went up Moses, and Aaron, Nadab, and Abihu, and seventy of the elders of Israel:
EXOD|24|10|And they saw the God of Israel: and there was under his feet as it were a paved work of a sapphire stone, and as it were the body of heaven in his clearness.
EXOD|24|11|And upon the nobles of the children of Israel he laid not his hand: also they saw God, and did eat and drink.
EXOD|24|12|And the LORD said unto Moses, Come up to me into the mount, and be there: and I will give thee tables of stone, and a law, and commandments which I have written; that thou mayest teach them.
EXOD|24|13|And Moses rose up, and his minister Joshua: and Moses went up into the mount of God.
EXOD|24|14|And he said unto the elders, Tarry ye here for us, until we come again unto you: and, behold, Aaron and Hur are with you: if any man have any matters to do, let him come unto them.
EXOD|24|15|And Moses went up into the mount, and a cloud covered the mount.
EXOD|24|16|And the glory of the LORD abode upon mount Sinai, and the cloud covered it six days: and the seventh day he called unto Moses out of the midst of the cloud.
EXOD|24|17|And the sight of the glory of the LORD was like devouring fire on the top of the mount in the eyes of the children of Israel.
EXOD|24|18|And Moses went into the midst of the cloud, and gat him up into the mount: and Moses was in the mount forty days and forty nights.
EXOD|25|1|And the LORD spake unto Moses, saying,
EXOD|25|2|Speak unto the children of Israel, that they bring me an offering: of every man that giveth it willingly with his heart ye shall take my offering.
EXOD|25|3|And this is the offering which ye shall take of them; gold, and silver, and brass,
EXOD|25|4|And blue, and purple, and scarlet, and fine linen, and goats' hair,
EXOD|25|5|And rams' skins dyed red, and badgers' skins, and shittim wood,
EXOD|25|6|Oil for the light, spices for anointing oil, and for sweet incense,
EXOD|25|7|Onyx stones, and stones to be set in the ephod, and in the breastplate.
EXOD|25|8|And let them make me a sanctuary; that I may dwell among them.
EXOD|25|9|According to all that I show thee, after the pattern of the tabernacle, and the pattern of all the instruments thereof, even so shall ye make it.
EXOD|25|10|And they shall make an ark of shittim wood: two cubits and a half shall be the length thereof, and a cubit and a half the breadth thereof, and a cubit and a half the height thereof.
EXOD|25|11|And thou shalt overlay it with pure gold, within and without shalt thou overlay it, and shalt make upon it a crown of gold round about.
EXOD|25|12|And thou shalt cast four rings of gold for it, and put them in the four corners thereof; and two rings shall be in the one side of it, and two rings in the other side of it.
EXOD|25|13|And thou shalt make staves of shittim wood, and overlay them with gold.
EXOD|25|14|And thou shalt put the staves into the rings by the sides of the ark, that the ark may be borne with them.
EXOD|25|15|The staves shall be in the rings of the ark: they shall not be taken from it.
EXOD|25|16|And thou shalt put into the ark the testimony which I shall give thee.
EXOD|25|17|And thou shalt make a mercy seat of pure gold: two cubits and a half shall be the length thereof, and a cubit and a half the breadth thereof.
EXOD|25|18|And thou shalt make two cherubim of gold, of beaten work shalt thou make them, in the two ends of the mercy seat.
EXOD|25|19|And make one cherub on the one end, and the other cherub on the other end: even of the mercy seat shall ye make the cherubim on the two ends thereof.
EXOD|25|20|And the cherubim shall stretch forth their wings on high, covering the mercy seat with their wings, and their faces shall look one to another; toward the mercy seat shall the faces of the cherubim be.
EXOD|25|21|And thou shalt put the mercy seat above upon the ark; and in the ark thou shalt put the testimony that I shall give thee.
EXOD|25|22|And there I will meet with thee, and I will commune with thee from above the mercy seat, from between the two cherubim which are upon the ark of the testimony, of all things which I will give thee in commandment unto the children of Israel.
EXOD|25|23|Thou shalt also make a table of shittim wood: two cubits shall be the length thereof, and a cubit the breadth thereof, and a cubit and a half the height thereof.
EXOD|25|24|And thou shalt overlay it with pure gold, and make thereto a crown of gold round about.
EXOD|25|25|And thou shalt make unto it a border of an hand breadth round about, and thou shalt make a golden crown to the border thereof round about.
EXOD|25|26|And thou shalt make for it four rings of gold, and put the rings in the four corners that are on the four feet thereof.
EXOD|25|27|Over against the border shall the rings be for places of the staves to bear the table.
EXOD|25|28|And thou shalt make the staves of shittim wood, and overlay them with gold, that the table may be borne with them.
EXOD|25|29|And thou shalt make the dishes thereof, and spoons thereof, and covers thereof, and bowls thereof, to cover withal: of pure gold shalt thou make them.
EXOD|25|30|And thou shalt set upon the table showbread before me always.
EXOD|25|31|And thou shalt make a candlestick of pure gold: of beaten work shall the candlestick be made: his shaft, and his branches, his bowls, his knops, and his flowers, shall be of the same.
EXOD|25|32|And six branches shall come out of the sides of it; three branches of the candlestick out of the one side, and three branches of the candlestick out of the other side:
EXOD|25|33|Three bowls made like unto almonds, with a knop and a flower in one branch; and three bowls made like almonds in the other branch, with a knop and a flower: so in the six branches that come out of the candlestick.
EXOD|25|34|And in the candlesticks shall be four bowls made like unto almonds, with their knops and their flowers.
EXOD|25|35|And there shall be a knop under two branches of the same, and a knop under two branches of the same, and a knop under two branches of the same, according to the six branches that proceed out of the candlestick.
EXOD|25|36|Their knops and their branches shall be of the same: all it shall be one beaten work of pure gold.
EXOD|25|37|And thou shalt make the seven lamps thereof: and they shall light the lamps thereof, that they may give light over against it.
EXOD|25|38|And the tongs thereof, and the snuffdishes thereof, shall be of pure gold.
EXOD|25|39|Of a talent of pure gold shall he make it, with all these vessels.
EXOD|25|40|And look that thou make them after their pattern, which was showed thee in the mount.
EXOD|26|1|Moreover thou shalt make the tabernacle with ten curtains of fine twined linen, and blue, and purple, and scarlet: with cherubim of cunning work shalt thou make them.
EXOD|26|2|The length of one curtain shall be eight and twenty cubits, and the breadth of one curtain four cubits: and every one of the curtains shall have one measure.
EXOD|26|3|The five curtains shall be coupled together one to another; and other five curtains shall be coupled one to another.
EXOD|26|4|And thou shalt make loops of blue upon the edge of the one curtain from the selvedge in the coupling; and likewise shalt thou make in the uttermost edge of another curtain, in the coupling of the second.
EXOD|26|5|Fifty loops shalt thou make in the one curtain, and fifty loops shalt thou make in the edge of the curtain that is in the coupling of the second; that the loops may take hold one of another.
EXOD|26|6|And thou shalt make fifty taches of gold, and couple the curtains together with the taches: and it shall be one tabernacle.
EXOD|26|7|And thou shalt make curtains of goats' hair to be a covering upon the tabernacle: eleven curtains shalt thou make.
EXOD|26|8|The length of one curtain shall be thirty cubits, and the breadth of one curtain four cubits: and the eleven curtains shall be all of one measure.
EXOD|26|9|And thou shalt couple five curtains by themselves, and six curtains by themselves, and shalt double the sixth curtain in the forefront of the tabernacle.
EXOD|26|10|And thou shalt make fifty loops on the edge of the one curtain that is outmost in the coupling, and fifty loops in the edge of the curtain which coupleth the second.
EXOD|26|11|And thou shalt make fifty taches of brass, and put the taches into the loops, and couple the tent together, that it may be one.
EXOD|26|12|And the remnant that remaineth of the curtains of the tent, the half curtain that remaineth, shall hang over the backside of the tabernacle.
EXOD|26|13|And a cubit on the one side, and a cubit on the other side of that which remaineth in the length of the curtains of the tent, it shall hang over the sides of the tabernacle on this side and on that side, to cover it.
EXOD|26|14|And thou shalt make a covering for the tent of rams' skins dyed red, and a covering above of badgers' skins.
EXOD|26|15|And thou shalt make boards for the tabernacle of shittim wood standing up.
EXOD|26|16|Ten cubits shall be the length of a board, and a cubit and a half shall be the breadth of one board.
EXOD|26|17|Two tenons shall there be in one board, set in order one against another: thus shalt thou make for all the boards of the tabernacle.
EXOD|26|18|And thou shalt make the boards for the tabernacle, twenty boards on the south side southward.
EXOD|26|19|And thou shalt make forty sockets of silver under the twenty boards; two sockets under one board for his two tenons, and two sockets under another board for his two tenons.
EXOD|26|20|And for the second side of the tabernacle on the north side there shall be twenty boards:
EXOD|26|21|And their forty sockets of silver; two sockets under one board, and two sockets under another board.
EXOD|26|22|And for the sides of the tabernacle westward thou shalt make six boards.
EXOD|26|23|And two boards shalt thou make for the corners of the tabernacle in the two sides.
EXOD|26|24|And they shall be coupled together beneath, and they shall be coupled together above the head of it unto one ring: thus shall it be for them both; they shall be for the two corners.
EXOD|26|25|And they shall be eight boards, and their sockets of silver, sixteen sockets; two sockets under one board, and two sockets under another board.
EXOD|26|26|And thou shalt make bars of shittim wood; five for the boards of the one side of the tabernacle,
EXOD|26|27|And five bars for the boards of the other side of the tabernacle, and five bars for the boards of the side of the tabernacle, for the two sides westward.
EXOD|26|28|And the middle bar in the midst of the boards shall reach from end to end.
EXOD|26|29|And thou shalt overlay the boards with gold, and make their rings of gold for places for the bars: and thou shalt overlay the bars with gold.
EXOD|26|30|And thou shalt rear up the tabernacle according to the fashion thereof which was showed thee in the mount.
EXOD|26|31|And thou shalt make a vail of blue, and purple, and scarlet, and fine twined linen of cunning work: with cherubim shall it be made:
EXOD|26|32|And thou shalt hang it upon four pillars of shittim wood overlaid with gold: their hooks shall be of gold, upon the four sockets of silver.
EXOD|26|33|And thou shalt hang up the vail under the taches, that thou mayest bring in thither within the vail the ark of the testimony: and the vail shall divide unto you between the holy place and the most holy.
EXOD|26|34|And thou shalt put the mercy seat upon the ark of the testimony in the most holy place.
EXOD|26|35|And thou shalt set the table without the vail, and the candlestick over against the table on the side of the tabernacle toward the south: and thou shalt put the table on the north side.
EXOD|26|36|And thou shalt make an hanging for the door of the tent, of blue, and purple, and scarlet, and fine twined linen, wrought with needlework.
EXOD|26|37|And thou shalt make for the hanging five pillars of shittim wood, and overlay them with gold, and their hooks shall be of gold: and thou shalt cast five sockets of brass for them.
EXOD|27|1|And thou shalt make an altar of shittim wood, five cubits long, and five cubits broad; the altar shall be foursquare: and the height thereof shall be three cubits.
EXOD|27|2|And thou shalt make the horns of it upon the four corners thereof: his horns shall be of the same: and thou shalt overlay it with brass.
EXOD|27|3|And thou shalt make his pans to receive his ashes, and his shovels, and his basins, and his fleshhooks, and his firepans: all the vessels thereof thou shalt make of brass.
EXOD|27|4|And thou shalt make for it a grate of network of brass; and upon the net shalt thou make four brazen rings in the four corners thereof.
EXOD|27|5|And thou shalt put it under the compass of the altar beneath, that the net may be even to the midst of the altar.
EXOD|27|6|And thou shalt make staves for the altar, staves of shittim wood, and overlay them with brass.
EXOD|27|7|And the staves shall be put into the rings, and the staves shall be upon the two sides of the altar, to bear it.
EXOD|27|8|Hollow with boards shalt thou make it: as it was showed thee in the mount, so shall they make it.
EXOD|27|9|And thou shalt make the court of the tabernacle: for the south side southward there shall be hangings for the court of fine twined linen of an hundred cubits long for one side:
EXOD|27|10|And the twenty pillars thereof and their twenty sockets shall be of brass; the hooks of the pillars and their fillets shall be of silver.
EXOD|27|11|And likewise for the north side in length there shall be hangings of an hundred cubits long, and his twenty pillars and their twenty sockets of brass; the hooks of the pillars and their fillets of silver.
EXOD|27|12|And for the breadth of the court on the west side shall be hangings of fifty cubits: their pillars ten, and their sockets ten.
EXOD|27|13|And the breadth of the court on the east side eastward shall be fifty cubits.
EXOD|27|14|The hangings of one side of the gate shall be fifteen cubits: their pillars three, and their sockets three.
EXOD|27|15|And on the other side shall be hangings fifteen cubits: their pillars three, and their sockets three.
EXOD|27|16|And for the gate of the court shall be an hanging of twenty cubits, of blue, and purple, and scarlet, and fine twined linen, wrought with needlework: and their pillars shall be four, and their sockets four.
EXOD|27|17|All the pillars round about the court shall be filleted with silver; their hooks shall be of silver, and their sockets of brass.
EXOD|27|18|The length of the court shall be an hundred cubits, and the breadth fifty every where, and the height five cubits of fine twined linen, and their sockets of brass.
EXOD|27|19|All the vessels of the tabernacle in all the service thereof, and all the pins thereof, and all the pins of the court, shall be of brass.
EXOD|27|20|And thou shalt command the children of Israel, that they bring thee pure oil olive beaten for the light, to cause the lamp to burn always.
EXOD|27|21|In the tabernacle of the congregation without the vail, which is before the testimony, Aaron and his sons shall order it from evening to morning before the LORD: it shall be a statute for ever unto their generations on the behalf of the children of Israel.
EXOD|28|1|And take thou unto thee Aaron thy brother, and his sons with him, from among the children of Israel, that he may minister unto me in the priest's office, even Aaron, Nadab and Abihu, Eleazar and Ithamar, Aaron's sons.
EXOD|28|2|And thou shalt make holy garments for Aaron thy brother for glory and for beauty.
EXOD|28|3|And thou shalt speak unto all that are wise hearted, whom I have filled with the spirit of wisdom, that they may make Aaron's garments to consecrate him, that he may minister unto me in the priest's office.
EXOD|28|4|And these are the garments which they shall make; a breastplate, and an ephod, and a robe, and a broidered coat, a mitre, and a girdle: and they shall make holy garments for Aaron thy brother, and his sons, that he may minister unto me in the priest's office.
EXOD|28|5|And they shall take gold, and blue, and purple, and scarlet, and fine linen.
EXOD|28|6|And they shall make the ephod of gold, of blue, and of purple, of scarlet, and fine twined linen, with cunning work.
EXOD|28|7|It shall have the two shoulderpieces thereof joined at the two edges thereof; and so it shall be joined together.
EXOD|28|8|And the curious girdle of the ephod, which is upon it, shall be of the same, according to the work thereof; even of gold, of blue, and purple, and scarlet, and fine twined linen.
EXOD|28|9|And thou shalt take two onyx stones, and grave on them the names of the children of Israel:
EXOD|28|10|Six of their names on one stone, and the other six names of the rest on the other stone, according to their birth.
EXOD|28|11|With the work of an engraver in stone, like the engravings of a signet, shalt thou engrave the two stones with the names of the children of Israel: thou shalt make them to be set in ouches of gold.
EXOD|28|12|And thou shalt put the two stones upon the shoulders of the ephod for stones of memorial unto the children of Israel: and Aaron shall bear their names before the LORD upon his two shoulders for a memorial.
EXOD|28|13|And thou shalt make ouches of gold;
EXOD|28|14|And two chains of pure gold at the ends; of wreathed work shalt thou make them, and fasten the wreathed chains to the ouches.
EXOD|28|15|And thou shalt make the breastplate of judgment with cunning work; after the work of the ephod thou shalt make it; of gold, of blue, and of purple, and of scarlet, and of fine twined linen, shalt thou make it.
EXOD|28|16|Foursquare it shall be being doubled; a span shall be the length thereof, and a span shall be the breadth thereof.
EXOD|28|17|And thou shalt set in it settings of stones, even four rows of stones: the first row shall be a sardius, a topaz, and a carbuncle: this shall be the first row.
EXOD|28|18|And the second row shall be an emerald, a sapphire, and a diamond.
EXOD|28|19|And the third row a ligure, an agate, and an amethyst.
EXOD|28|20|And the fourth row a beryl, and an onyx, and a jasper: they shall be set in gold in their inclosings.
EXOD|28|21|And the stones shall be with the names of the children of Israel, twelve, according to their names, like the engravings of a signet; every one with his name shall they be according to the twelve tribes.
EXOD|28|22|And thou shalt make upon the breastplate chains at the ends of wreathed work of pure gold.
EXOD|28|23|And thou shalt make upon the breastplate two rings of gold, and shalt put the two rings on the two ends of the breastplate.
EXOD|28|24|And thou shalt put the two wreathed chains of gold in the two rings which are on the ends of the breastplate.
EXOD|28|25|And the other two ends of the two wreathed chains thou shalt fasten in the two ouches, and put them on the shoulderpieces of the ephod before it.
EXOD|28|26|And thou shalt make two rings of gold, and thou shalt put them upon the two ends of the breastplate in the border thereof, which is in the side of the ephod inward.
EXOD|28|27|And two other rings of gold thou shalt make, and shalt put them on the two sides of the ephod underneath, toward the forepart thereof, over against the other coupling thereof, above the curious girdle of the ephod.
EXOD|28|28|And they shall bind the breastplate by the rings thereof unto the rings of the ephod with a lace of blue, that it may be above the curious girdle of the ephod, and that the breastplate be not loosed from the ephod.
EXOD|28|29|And Aaron shall bear the names of the children of Israel in the breastplate of judgment upon his heart, when he goeth in unto the holy place, for a memorial before the LORD continually.
EXOD|28|30|And thou shalt put in the breastplate of judgment the Urim and the Thummim; and they shall be upon Aaron's heart, when he goeth in before the LORD: and Aaron shall bear the judgment of the children of Israel upon his heart before the LORD continually.
EXOD|28|31|And thou shalt make the robe of the ephod all of blue.
EXOD|28|32|And there shall be an hole in the top of it, in the midst thereof: it shall have a binding of woven work round about the hole of it, as it were the hole of an habergeon, that it be not rent.
EXOD|28|33|And beneath upon the hem of it thou shalt make pomegranates of blue, and of purple, and of scarlet, round about the hem thereof; and bells of gold between them round about:
EXOD|28|34|A golden bell and a pomegranate, a golden bell and a pomegranate, upon the hem of the robe round about.
EXOD|28|35|And it shall be upon Aaron to minister: and his sound shall be heard when he goeth in unto the holy place before the LORD, and when he cometh out, that he die not.
EXOD|28|36|And thou shalt make a plate of pure gold, and grave upon it, like the engravings of a signet, HOLINESS TO THE LORD.
EXOD|28|37|And thou shalt put it on a blue lace, that it may be upon the mitre; upon the forefront of the mitre it shall be.
EXOD|28|38|And it shall be upon Aaron's forehead, that Aaron may bear the iniquity of the holy things, which the children of Israel shall hallow in all their holy gifts; and it shall be always upon his forehead, that they may be accepted before the LORD.
EXOD|28|39|And thou shalt embroider the coat of fine linen, and thou shalt make the mitre of fine linen, and thou shalt make the girdle of needlework.
EXOD|28|40|And for Aaron's sons thou shalt make coats, and thou shalt make for them girdles, and bonnets shalt thou make for them, for glory and for beauty.
EXOD|28|41|And thou shalt put them upon Aaron thy brother, and his sons with him; and shalt anoint them, and consecrate them, and sanctify them, that they may minister unto me in the priest's office.
EXOD|28|42|And thou shalt make them linen breeches to cover their nakedness; from the loins even unto the thighs they shall reach:
EXOD|28|43|And they shall be upon Aaron, and upon his sons, when they come in unto the tabernacle of the congregation, or when they come near unto the altar to minister in the holy place; that they bear not iniquity, and die: it shall be a statute for ever unto him and his seed after him.
EXOD|29|1|And this is the thing that thou shalt do unto them to hallow them, to minister unto me in the priest's office: Take one young bullock, and two rams without blemish,
EXOD|29|2|And unleavened bread, and cakes unleavened tempered with oil, and wafers unleavened anointed with oil: of wheaten flour shalt thou make them.
EXOD|29|3|And thou shalt put them into one basket, and bring them in the basket, with the bullock and the two rams.
EXOD|29|4|And Aaron and his sons thou shalt bring unto the door of the tabernacle of the congregation, and shalt wash them with water.
EXOD|29|5|And thou shalt take the garments, and put upon Aaron the coat, and the robe of the ephod, and the ephod, and the breastplate, and gird him with the curious girdle of the ephod:
EXOD|29|6|And thou shalt put the mitre upon his head, and put the holy crown upon the mitre.
EXOD|29|7|Then shalt thou take the anointing oil, and pour it upon his head, and anoint him.
EXOD|29|8|And thou shalt bring his sons, and put coats upon them.
EXOD|29|9|And thou shalt gird them with girdles, Aaron and his sons, and put the bonnets on them: and the priest's office shall be theirs for a perpetual statute: and thou shalt consecrate Aaron and his sons.
EXOD|29|10|And thou shalt cause a bullock to be brought before the tabernacle of the congregation: and Aaron and his sons shall put their hands upon the head of the bullock.
EXOD|29|11|And thou shalt kill the bullock before the LORD, by the door of the tabernacle of the congregation.
EXOD|29|12|And thou shalt take of the blood of the bullock, and put it upon the horns of the altar with thy finger, and pour all the blood beside the bottom of the altar.
EXOD|29|13|And thou shalt take all the fat that covereth the inwards, and the caul that is above the liver, and the two kidneys, and the fat that is upon them, and burn them upon the altar.
EXOD|29|14|But the flesh of the bullock, and his skin, and his dung, shalt thou burn with fire without the camp: it is a sin offering.
EXOD|29|15|Thou shalt also take one ram; and Aaron and his sons shall put their hands upon the head of the ram.
EXOD|29|16|And thou shalt slay the ram, and thou shalt take his blood, and sprinkle it round about upon the altar.
EXOD|29|17|And thou shalt cut the ram in pieces, and wash the inwards of him, and his legs, and put them unto his pieces, and unto his head.
EXOD|29|18|And thou shalt burn the whole ram upon the altar: it is a burnt offering unto the LORD: it is a sweet savor, an offering made by fire unto the LORD.
EXOD|29|19|And thou shalt take the other ram; and Aaron and his sons shall put their hands upon the head of the ram.
EXOD|29|20|Then shalt thou kill the ram, and take of his blood, and put it upon the tip of the right ear of Aaron, and upon the tip of the right ear of his sons, and upon the thumb of their right hand, and upon the great toe of their right foot, and sprinkle the blood upon the altar round about.
EXOD|29|21|And thou shalt take of the blood that is upon the altar, and of the anointing oil, and sprinkle it upon Aaron, and upon his garments, and upon his sons, and upon the garments of his sons with him: and he shall be hallowed, and his garments, and his sons, and his sons' garments with him.
EXOD|29|22|Also thou shalt take of the ram the fat and the rump, and the fat that covereth the inwards, and the caul above the liver, and the two kidneys, and the fat that is upon them, and the right shoulder; for it is a ram of consecration:
EXOD|29|23|And one loaf of bread, and one cake of oiled bread, and one wafer out of the basket of the unleavened bread that is before the LORD:
EXOD|29|24|And thou shalt put all in the hands of Aaron, and in the hands of his sons; and shalt wave them for a wave offering before the LORD.
EXOD|29|25|And thou shalt receive them of their hands, and burn them upon the altar for a burnt offering, for a sweet savor before the LORD: it is an offering made by fire unto the LORD.
EXOD|29|26|And thou shalt take the breast of the ram of Aaron's consecration, and wave it for a wave offering before the LORD: and it shall be thy part.
EXOD|29|27|And thou shalt sanctify the breast of the wave offering, and the shoulder of the heave offering, which is waved, and which is heaved up, of the ram of the consecration, even of that which is for Aaron, and of that which is for his sons:
EXOD|29|28|And it shall be Aaron's and his sons' by a statute for ever from the children of Israel: for it is an heave offering: and it shall be an heave offering from the children of Israel of the sacrifice of their peace offerings, even their heave offering unto the LORD.
EXOD|29|29|And the holy garments of Aaron shall be his sons' after him, to be anointed therein, and to be consecrated in them.
EXOD|29|30|And that son that is priest in his stead shall put them on seven days, when he cometh into the tabernacle of the congregation to minister in the holy place.
EXOD|29|31|And thou shalt take the ram of the consecration, and seethe his flesh in the holy place.
EXOD|29|32|And Aaron and his sons shall eat the flesh of the ram, and the bread that is in the basket by the door of the tabernacle of the congregation.
EXOD|29|33|And they shall eat those things wherewith the atonement was made, to consecrate and to sanctify them: but a stranger shall not eat thereof, because they are holy.
EXOD|29|34|And if ought of the flesh of the consecrations, or of the bread, remain unto the morning, then thou shalt burn the remainder with fire: it shall not be eaten, because it is holy.
EXOD|29|35|And thus shalt thou do unto Aaron, and to his sons, according to all things which I have commanded thee: seven days shalt thou consecrate them.
EXOD|29|36|And thou shalt offer every day a bullock for a sin offering for atonement: and thou shalt cleanse the altar, when thou hast made an atonement for it, and thou shalt anoint it, to sanctify it.
EXOD|29|37|Seven days thou shalt make an atonement for the altar, and sanctify it; and it shall be an altar most holy: whatsoever toucheth the altar shall be holy.
EXOD|29|38|Now this is that which thou shalt offer upon the altar; two lambs of the first year day by day continually.
EXOD|29|39|The one lamb thou shalt offer in the morning; and the other lamb thou shalt offer at even:
EXOD|29|40|And with the one lamb a tenth deal of flour mingled with the fourth part of an hin of beaten oil; and the fourth part of an hin of wine for a drink offering.
EXOD|29|41|And the other lamb thou shalt offer at even, and shalt do thereto according to the meat offering of the morning, and according to the drink offering thereof, for a sweet savor, an offering made by fire unto the LORD.
EXOD|29|42|This shall be a continual burnt offering throughout your generations at the door of the tabernacle of the congregation before the LORD: where I will meet you, to speak there unto thee.
EXOD|29|43|And there I will meet with the children of Israel, and the tabernacle shall be sanctified by my glory.
EXOD|29|44|And I will sanctify the tabernacle of the congregation, and the altar: I will sanctify also both Aaron and his sons, to minister to me in the priest's office.
EXOD|29|45|And I will dwell among the children of Israel, and will be their God.
EXOD|29|46|And they shall know that I am the LORD their God, that brought them forth out of the land of Egypt, that I may dwell among them: I am the LORD their God.
EXOD|30|1|And thou shalt make an altar to burn incense upon: of shittim wood shalt thou make it.
EXOD|30|2|A cubit shall be the length thereof, and a cubit the breadth thereof; foursquare shall it be: and two cubits shall be the height thereof: the horns thereof shall be of the same.
EXOD|30|3|And thou shalt overlay it with pure gold, the top thereof, and the sides thereof round about, and the horns thereof; and thou shalt make unto it a crown of gold round about.
EXOD|30|4|And two golden rings shalt thou make to it under the crown of it, by the two corners thereof, upon the two sides of it shalt thou make it; and they shall be for places for the staves to bear it withal.
EXOD|30|5|And thou shalt make the staves of shittim wood, and overlay them with gold.
EXOD|30|6|And thou shalt put it before the vail that is by the ark of the testimony, before the mercy seat that is over the testimony, where I will meet with thee.
EXOD|30|7|And Aaron shall burn thereon sweet incense every morning: when he dresseth the lamps, he shall burn incense upon it.
EXOD|30|8|And when Aaron lighteth the lamps at even, he shall burn incense upon it, a perpetual incense before the LORD throughout your generations.
EXOD|30|9|Ye shall offer no strange incense thereon, nor burnt sacrifice, nor meat offering; neither shall ye pour drink offering thereon.
EXOD|30|10|And Aaron shall make an atonement upon the horns of it once in a year with the blood of the sin offering of atonements: once in the year shall he make atonement upon it throughout your generations: it is most holy unto the LORD.
EXOD|30|11|And the LORD spake unto Moses, saying,
EXOD|30|12|When thou takest the sum of the children of Israel after their number, then shall they give every man a ransom for his soul unto the LORD, when thou numberest them; that there be no plague among them, when thou numberest them.
EXOD|30|13|This they shall give, every one that passeth among them that are numbered, half a shekel after the shekel of the sanctuary: (a shekel is twenty gerahs:) an half shekel shall be the offering of the LORD.
EXOD|30|14|Every one that passeth among them that are numbered, from twenty years old and above, shall give an offering unto the LORD.
EXOD|30|15|The rich shall not give more, and the poor shall not give less than half a shekel, when they give an offering unto the LORD, to make an atonement for your souls.
EXOD|30|16|And thou shalt take the atonement money of the children of Israel, and shalt appoint it for the service of the tabernacle of the congregation; that it may be a memorial unto the children of Israel before the LORD, to make an atonement for your souls.
EXOD|30|17|And the LORD spake unto Moses, saying,
EXOD|30|18|Thou shalt also make a laver of brass, and his foot also of brass, to wash withal: and thou shalt put it between the tabernacle of the congregation and the altar, and thou shalt put water therein.
EXOD|30|19|For Aaron and his sons shall wash their hands and their feet thereat:
EXOD|30|20|When they go into the tabernacle of the congregation, they shall wash with water, that they die not; or when they come near to the altar to minister, to burn offering made by fire unto the LORD:
EXOD|30|21|So they shall wash their hands and their feet, that they die not: and it shall be a statute for ever to them, even to him and to his seed throughout their generations.
EXOD|30|22|Moreover the LORD spake unto Moses, saying,
EXOD|30|23|Take thou also unto thee principal spices, of pure myrrh five hundred shekels, and of sweet cinnamon half so much, even two hundred and fifty shekels, and of sweet calamus two hundred and fifty shekels,
EXOD|30|24|And of cassia five hundred shekels, after the shekel of the sanctuary, and of oil olive an hin:
EXOD|30|25|And thou shalt make it an oil of holy ointment, an ointment compound after the art of the apothecary: it shall be an holy anointing oil.
EXOD|30|26|And thou shalt anoint the tabernacle of the congregation therewith, and the ark of the testimony,
EXOD|30|27|And the table and all his vessels, and the candlestick and his vessels, and the altar of incense,
EXOD|30|28|And the altar of burnt offering with all his vessels, and the laver and his foot.
EXOD|30|29|And thou shalt sanctify them, that they may be most holy: whatsoever toucheth them shall be holy.
EXOD|30|30|And thou shalt anoint Aaron and his sons, and consecrate them, that they may minister unto me in the priest's office.
EXOD|30|31|And thou shalt speak unto the children of Israel, saying, This shall be an holy anointing oil unto me throughout your generations.
EXOD|30|32|Upon man's flesh shall it not be poured, neither shall ye make any other like it, after the composition of it: it is holy, and it shall be holy unto you.
EXOD|30|33|Whosoever compoundeth any like it, or whosoever putteth any of it upon a stranger, shall even be cut off from his people.
EXOD|30|34|And the LORD said unto Moses, Take unto thee sweet spices, stacte, and onycha, and galbanum; these sweet spices with pure frankincense: of each shall there be a like weight:
EXOD|30|35|And thou shalt make it a perfume, a confection after the art of the apothecary, tempered together, pure and holy:
EXOD|30|36|And thou shalt beat some of it very small, and put of it before the testimony in the tabernacle of the congregation, where I will meet with thee: it shall be unto you most holy.
EXOD|30|37|And as for the perfume which thou shalt make, ye shall not make to yourselves according to the composition thereof: it shall be unto thee holy for the LORD.
EXOD|30|38|Whosoever shall make like unto that, to smell thereto, shall even be cut off from his people.
EXOD|31|1|And the LORD spake unto Moses, saying,
EXOD|31|2|See, I have called by name Bezaleel the son of Uri, the son of Hur, of the tribe of Judah:
EXOD|31|3|And I have filled him with the spirit of God, in wisdom, and in understanding, and in knowledge, and in all manner of workmanship,
EXOD|31|4|To devise cunning works, to work in gold, and in silver, and in brass,
EXOD|31|5|And in cutting of stones, to set them, and in carving of timber, to work in all manner of workmanship.
EXOD|31|6|And I, behold, I have given with him Aholiab, the son of Ahisamach, of the tribe of Dan: and in the hearts of all that are wise hearted I have put wisdom, that they may make all that I have commanded thee;
EXOD|31|7|The tabernacle of the congregation, and the ark of the testimony, and the mercy seat that is thereupon, and all the furniture of the tabernacle,
EXOD|31|8|And the table and his furniture, and the pure candlestick with all his furniture, and the altar of incense,
EXOD|31|9|And the altar of burnt offering with all his furniture, and the laver and his foot,
EXOD|31|10|And the cloths of service, and the holy garments for Aaron the priest, and the garments of his sons, to minister in the priest's office,
EXOD|31|11|And the anointing oil, and sweet incense for the holy place: according to all that I have commanded thee shall they do.
EXOD|31|12|And the LORD spake unto Moses, saying,
EXOD|31|13|Speak thou also unto the children of Israel, saying, Verily my sabbaths ye shall keep: for it is a sign between me and you throughout your generations; that ye may know that I am the LORD that doth sanctify you.
EXOD|31|14|Ye shall keep the sabbath therefore; for it is holy unto you: every one that defileth it shall surely be put to death: for whosoever doeth any work therein, that soul shall be cut off from among his people.
EXOD|31|15|Six days may work be done; but in the seventh is the sabbath of rest, holy to the LORD: whosoever doeth any work in the sabbath day, he shall surely be put to death.
EXOD|31|16|Wherefore the children of Israel shall keep the sabbath, to observe the sabbath throughout their generations, for a perpetual covenant.
EXOD|31|17|It is a sign between me and the children of Israel for ever: for in six days the LORD made heaven and earth, and on the seventh day he rested, and was refreshed.
EXOD|31|18|And he gave unto Moses, when he had made an end of communing with him upon mount Sinai, two tables of testimony, tables of stone, written with the finger of God.
EXOD|32|1|And when the people saw that Moses delayed to come down out of the mount, the people gathered themselves together unto Aaron, and said unto him, Up, make us gods, which shall go before us; for as for this Moses, the man that brought us up out of the land of Egypt, we wot not what is become of him.
EXOD|32|2|And Aaron said unto them, Break off the golden earrings, which are in the ears of your wives, of your sons, and of your daughters, and bring them unto me.
EXOD|32|3|And all the people brake off the golden earrings which were in their ears, and brought them unto Aaron.
EXOD|32|4|And he received them at their hand, and fashioned it with a graving tool, after he had made it a molten calf: and they said, These be thy gods, O Israel, which brought thee up out of the land of Egypt.
EXOD|32|5|And when Aaron saw it, he built an altar before it; and Aaron made proclamation, and said, To morrow is a feast to the LORD.
EXOD|32|6|And they rose up early on the morrow, and offered burnt offerings, and brought peace offerings; and the people sat down to eat and to drink, and rose up to play.
EXOD|32|7|And the LORD said unto Moses, Go, get thee down; for thy people, which thou broughtest out of the land of Egypt, have corrupted themselves:
EXOD|32|8|They have turned aside quickly out of the way which I commanded them: they have made them a molten calf, and have worshipped it, and have sacrificed thereunto, and said, These be thy gods, O Israel, which have brought thee up out of the land of Egypt.
EXOD|32|9|And the LORD said unto Moses, I have seen this people, and, behold, it is a stiffnecked people:
EXOD|32|10|Now therefore let me alone, that my wrath may wax hot against them, and that I may consume them: and I will make of thee a great nation.
EXOD|32|11|And Moses besought the LORD his God, and said, LORD, why doth thy wrath wax hot against thy people, which thou hast brought forth out of the land of Egypt with great power, and with a mighty hand?
EXOD|32|12|Wherefore should the Egyptians speak, and say, For mischief did he bring them out, to slay them in the mountains, and to consume them from the face of the earth? Turn from thy fierce wrath, and repent of this evil against thy people.
EXOD|32|13|Remember Abraham, Isaac, and Israel, thy servants, to whom thou swarest by thine own self, and saidst unto them, I will multiply your seed as the stars of heaven, and all this land that I have spoken of will I give unto your seed, and they shall inherit it for ever.
EXOD|32|14|And the LORD repented of the evil which he thought to do unto his people.
EXOD|32|15|And Moses turned, and went down from the mount, and the two tables of the testimony were in his hand: the tables were written on both their sides; on the one side and on the other were they written.
EXOD|32|16|And the tables were the work of God, and the writing was the writing of God, graven upon the tables.
EXOD|32|17|And when Joshua heard the noise of the people as they shouted, he said unto Moses, There is a noise of war in the camp.
EXOD|32|18|And he said, It is not the voice of them that shout for mastery, neither is it the voice of them that cry for being overcome: but the noise of them that sing do I hear.
EXOD|32|19|And it came to pass, as soon as he came nigh unto the camp, that he saw the calf, and the dancing: and Moses' anger waxed hot, and he cast the tables out of his hands, and brake them beneath the mount.
EXOD|32|20|And he took the calf which they had made, and burnt it in the fire, and ground it to powder, and strewed it upon the water, and made the children of Israel drink of it.
EXOD|32|21|And Moses said unto Aaron, What did this people unto thee, that thou hast brought so great a sin upon them?
EXOD|32|22|And Aaron said, Let not the anger of my lord wax hot: thou knowest the people, that they are set on mischief.
EXOD|32|23|For they said unto me, Make us gods, which shall go before us: for as for this Moses, the man that brought us up out of the land of Egypt, we wot not what is become of him.
EXOD|32|24|And I said unto them, Whosoever hath any gold, let them break it off. So they gave it me: then I cast it into the fire, and there came out this calf.
EXOD|32|25|And when Moses saw that the people were naked; (for Aaron had made them naked unto their shame among their enemies:)
EXOD|32|26|Then Moses stood in the gate of the camp, and said, Who is on the LORD's side? let him come unto me. And all the sons of Levi gathered themselves together unto him.
EXOD|32|27|And he said unto them, Thus saith the LORD God of Israel, Put every man his sword by his side, and go in and out from gate to gate throughout the camp, and slay every man his brother, and every man his companion, and every man his neighbor.
EXOD|32|28|And the children of Levi did according to the word of Moses: and there fell of the people that day about three thousand men.
EXOD|32|29|For Moses had said, Consecrate yourselves today to the LORD, even every man upon his son, and upon his brother; that he may bestow upon you a blessing this day.
EXOD|32|30|And it came to pass on the morrow, that Moses said unto the people, Ye have sinned a great sin: and now I will go up unto the LORD; peradventure I shall make an atonement for your sin.
EXOD|32|31|And Moses returned unto the LORD, and said, Oh, this people have sinned a great sin, and have made them gods of gold.
EXOD|32|32|Yet now, if thou wilt forgive their sin--; and if not, blot me, I pray thee, out of thy book which thou hast written.
EXOD|32|33|And the LORD said unto Moses, Whosoever hath sinned against me, him will I blot out of my book.
EXOD|32|34|Therefore now go, lead the people unto the place of which I have spoken unto thee: behold, mine Angel shall go before thee: nevertheless in the day when I visit I will visit their sin upon them.
EXOD|32|35|And the LORD plagued the people, because they made the calf, which Aaron made.
EXOD|33|1|And the LORD said unto Moses, Depart, and go up hence, thou and the people which thou hast brought up out of the land of Egypt, unto the land which I sware unto Abraham, to Isaac, and to Jacob, saying, Unto thy seed will I give it:
EXOD|33|2|And I will send an angel before thee; and I will drive out the Canaanite, the Amorite, and the Hittite, and the Perizzite, the Hivite, and the Jebusite:
EXOD|33|3|Unto a land flowing with milk and honey: for I will not go up in the midst of thee; for thou art a stiffnecked people: lest I consume thee in the way.
EXOD|33|4|And when the people heard these evil tidings, they mourned: and no man did put on him his ornaments.
EXOD|33|5|For the LORD had said unto Moses, Say unto the children of Israel, Ye are a stiffnecked people: I will come up into the midst of thee in a moment, and consume thee: therefore now put off thy ornaments from thee, that I may know what to do unto thee.
EXOD|33|6|And the children of Israel stripped themselves of their ornaments by the mount Horeb.
EXOD|33|7|And Moses took the tabernacle, and pitched it without the camp, afar off from the camp, and called it the Tabernacle of the congregation. And it came to pass, that every one which sought the LORD went out unto the tabernacle of the congregation, which was without the camp.
EXOD|33|8|And it came to pass, when Moses went out unto the tabernacle, that all the people rose up, and stood every man at his tent door, and looked after Moses, until he was gone into the tabernacle.
EXOD|33|9|And it came to pass, as Moses entered into the tabernacle, the cloudy pillar descended, and stood at the door of the tabernacle, and the Lord talked with Moses.
EXOD|33|10|And all the people saw the cloudy pillar stand at the tabernacle door: and all the people rose up and worshipped, every man in his tent door.
EXOD|33|11|And the LORD spake unto Moses face to face, as a man speaketh unto his friend. And he turned again into the camp: but his servant Joshua, the son of Nun, a young man, departed not out of the tabernacle.
EXOD|33|12|And Moses said unto the LORD, See, thou sayest unto me, Bring up this people: and thou hast not let me know whom thou wilt send with me. Yet thou hast said, I know thee by name, and thou hast also found grace in my sight.
EXOD|33|13|Now therefore, I pray thee, if I have found grace in thy sight, show me now thy way, that I may know thee, that I may find grace in thy sight: and consider that this nation is thy people.
EXOD|33|14|And he said, My presence shall go with thee, and I will give thee rest.
EXOD|33|15|And he said unto him, If thy presence go not with me, carry us not up hence.
EXOD|33|16|For wherein shall it be known here that I and thy people have found grace in thy sight? is it not in that thou goest with us? so shall we be separated, I and thy people, from all the people that are upon the face of the earth.
EXOD|33|17|And the LORD said unto Moses, I will do this thing also that thou hast spoken: for thou hast found grace in my sight, and I know thee by name.
EXOD|33|18|And he said, I beseech thee, show me thy glory.
EXOD|33|19|And he said, I will make all my goodness pass before thee, and I will proclaim the name of the LORD before thee; and will be gracious to whom I will be gracious, and will show mercy on whom I will show mercy.
EXOD|33|20|And he said, Thou canst not see my face: for there shall no man see me, and live.
EXOD|33|21|And the LORD said, Behold, there is a place by me, and thou shalt stand upon a rock:
EXOD|33|22|And it shall come to pass, while my glory passeth by, that I will put thee in a cleft of the rock, and will cover thee with my hand while I pass by:
EXOD|33|23|And I will take away mine hand, and thou shalt see my back parts: but my face shall not be seen.
EXOD|34|1|And the LORD said unto Moses, Hew thee two tables of stone like unto the first: and I will write upon these tables the words that were in the first tables, which thou brakest.
EXOD|34|2|And be ready in the morning, and come up in the morning unto mount Sinai, and present thyself there to me in the top of the mount.
EXOD|34|3|And no man shall come up with thee, neither let any man be seen throughout all the mount; neither let the flocks nor herds feed before that mount.
EXOD|34|4|And he hewed two tables of stone like unto the first; and Moses rose up early in the morning, and went up unto mount Sinai, as the LORD had commanded him, and took in his hand the two tables of stone.
EXOD|34|5|And the LORD descended in the cloud, and stood with him there, and proclaimed the name of the LORD.
EXOD|34|6|And the LORD passed by before him, and proclaimed, The LORD, The LORD God, merciful and gracious, long-suffering, and abundant in goodness and truth,
EXOD|34|7|Keeping mercy for thousands, forgiving iniquity and transgression and sin, and that will by no means clear the guilty; visiting the iniquity of the fathers upon the children, and upon the children's children, unto the third and to the fourth generation.
EXOD|34|8|And Moses made haste, and bowed his head toward the earth, and worshipped.
EXOD|34|9|And he said, If now I have found grace in thy sight, O LORD, let my LORD, I pray thee, go among us; for it is a stiffnecked people; and pardon our iniquity and our sin, and take us for thine inheritance.
EXOD|34|10|And he said, Behold, I make a covenant: before all thy people I will do marvels, such as have not been done in all the earth, nor in any nation: and all the people among which thou art shall see the work of the LORD: for it is a terrible thing that I will do with thee.
EXOD|34|11|Observe thou that which I command thee this day: behold, I drive out before thee the Amorite, and the Canaanite, and the Hittite, and the Perizzite, and the Hivite, and the Jebusite.
EXOD|34|12|Take heed to thyself, lest thou make a covenant with the inhabitants of the land whither thou goest, lest it be for a snare in the midst of thee:
EXOD|34|13|But ye shall destroy their altars, break their images, and cut down their groves:
EXOD|34|14|For thou shalt worship no other god: for the LORD, whose name is Jealous, is a jealous God:
EXOD|34|15|Lest thou make a covenant with the inhabitants of the land, and they go a whoring after their gods, and do sacrifice unto their gods, and one call thee, and thou eat of his sacrifice;
EXOD|34|16|And thou take of their daughters unto thy sons, and their daughters go a whoring after their gods, and make thy sons go a whoring after their gods.
EXOD|34|17|Thou shalt make thee no molten gods.
EXOD|34|18|The feast of unleavened bread shalt thou keep. Seven days thou shalt eat unleavened bread, as I commanded thee, in the time of the month Abib: for in the month Abib thou camest out from Egypt.
EXOD|34|19|All that openeth the matrix is mine; and every firstling among thy cattle, whether ox or sheep, that is male.
EXOD|34|20|But the firstling of an ass thou shalt redeem with a lamb: and if thou redeem him not, then shalt thou break his neck. All the firstborn of thy sons thou shalt redeem. And none shall appear before me empty.
EXOD|34|21|Six days thou shalt work, but on the seventh day thou shalt rest: in earing time and in harvest thou shalt rest.
EXOD|34|22|And thou shalt observe the feast of weeks, of the firstfruits of wheat harvest, and the feast of ingathering at the year's end.
EXOD|34|23|Thrice in the year shall all your men children appear before the LORD God, the God of Israel.
EXOD|34|24|For I will cast out the nations before thee, and enlarge thy borders: neither shall any man desire thy land, when thou shalt go up to appear before the LORD thy God thrice in the year.
EXOD|34|25|Thou shalt not offer the blood of my sacrifice with leaven; neither shall the sacrifice of the feast of the passover be left unto the morning.
EXOD|34|26|The first of the firstfruits of thy land thou shalt bring unto the house of the LORD thy God. Thou shalt not seethe a kid in his mother's milk.
EXOD|34|27|And the LORD said unto Moses, Write thou these words: for after the tenor of these words I have made a covenant with thee and with Israel.
EXOD|34|28|And he was there with the LORD forty days and forty nights; he did neither eat bread, nor drink water. And he wrote upon the tables the words of the covenant, the ten commandments.
EXOD|34|29|And it came to pass, when Moses came down from mount Sinai with the two tables of testimony in Moses' hand, when he came down from the mount, that Moses wist not that the skin of his face shone while he talked with him.
EXOD|34|30|And when Aaron and all the children of Israel saw Moses, behold, the skin of his face shone; and they were afraid to come nigh him.
EXOD|34|31|And Moses called unto them; and Aaron and all the rulers of the congregation returned unto him: and Moses talked with them.
EXOD|34|32|And afterward all the children of Israel came nigh: and he gave them in commandment all that the LORD had spoken with him in mount Sinai.
EXOD|34|33|And till Moses had done speaking with them, he put a vail on his face.
EXOD|34|34|But when Moses went in before the LORD to speak with him, he took the vail off, until he came out. And he came out, and spake unto the children of Israel that which he was commanded.
EXOD|34|35|And the children of Israel saw the face of Moses, that the skin of Moses' face shone: and Moses put the vail upon his face again, until he went in to speak with him.
EXOD|35|1|And Moses gathered all the congregation of the children of Israel together, and said unto them, These are the words which the LORD hath commanded, that ye should do them.
EXOD|35|2|Six days shall work be done, but on the seventh day there shall be to you an holy day, a sabbath of rest to the LORD: whosoever doeth work therein shall be put to death.
EXOD|35|3|Ye shall kindle no fire throughout your habitations upon the sabbath day.
EXOD|35|4|And Moses spake unto all the congregation of the children of Israel, saying, This is the thing which the LORD commanded, saying,
EXOD|35|5|Take ye from among you an offering unto the LORD: whosoever is of a willing heart, let him bring it, an offering of the LORD; gold, and silver, and brass,
EXOD|35|6|And blue, and purple, and scarlet, and fine linen, and goats' hair,
EXOD|35|7|And rams' skins dyed red, and badgers' skins, and shittim wood,
EXOD|35|8|And oil for the light, and spices for anointing oil, and for the sweet incense,
EXOD|35|9|And onyx stones, and stones to be set for the ephod, and for the breastplate.
EXOD|35|10|And every wise hearted among you shall come, and make all that the LORD hath commanded;
EXOD|35|11|The tabernacle, his tent, and his covering, his taches, and his boards, his bars, his pillars, and his sockets,
EXOD|35|12|The ark, and the staves thereof, with the mercy seat, and the vail of the covering,
EXOD|35|13|The table, and his staves, and all his vessels, and the showbread,
EXOD|35|14|The candlestick also for the light, and his furniture, and his lamps, with the oil for the light,
EXOD|35|15|And the incense altar, and his staves, and the anointing oil, and the sweet incense, and the hanging for the door at the entering in of the tabernacle,
EXOD|35|16|The altar of burnt offering, with his brazen grate, his staves, and all his vessels, the laver and his foot,
EXOD|35|17|The hangings of the court, his pillars, and their sockets, and the hanging for the door of the court,
EXOD|35|18|The pins of the tabernacle, and the pins of the court, and their cords,
EXOD|35|19|The cloths of service, to do service in the holy place, the holy garments for Aaron the priest, and the garments of his sons, to minister in the priest's office.
EXOD|35|20|And all the congregation of the children of Israel departed from the presence of Moses.
EXOD|35|21|And they came, every one whose heart stirred him up, and every one whom his spirit made willing, and they brought the LORD's offering to the work of the tabernacle of the congregation, and for all his service, and for the holy garments.
EXOD|35|22|And they came, both men and women, as many as were willing hearted, and brought bracelets, and earrings, and rings, and tablets, all jewels of gold: and every man that offered, offered an offering of gold unto the LORD.
EXOD|35|23|And every man, with whom was found blue, and purple, and scarlet, and fine linen, and goats' hair, and red skins of rams, and badgers' skins, brought them.
EXOD|35|24|Every one that did offer an offering of silver and brass brought the LORD's offering: and every man, with whom was found shittim wood for any work of the service, brought it.
EXOD|35|25|And all the women that were wise hearted did spin with their hands, and brought that which they had spun, both of blue, and of purple, and of scarlet, and of fine linen.
EXOD|35|26|And all the women whose heart stirred them up in wisdom spun goats' hair.
EXOD|35|27|And the rulers brought onyx stones, and stones to be set, for the ephod, and for the breastplate;
EXOD|35|28|And spice, and oil for the light, and for the anointing oil, and for the sweet incense.
EXOD|35|29|The children of Israel brought a willing offering unto the LORD, every man and woman, whose heart made them willing to bring for all manner of work, which the LORD had commanded to be made by the hand of Moses.
EXOD|35|30|And Moses said unto the children of Israel, See, the LORD hath called by name Bezaleel the son of Uri, the son of Hur, of the tribe of Judah;
EXOD|35|31|And he hath filled him with the spirit of God, in wisdom, in understanding, and in knowledge, and in all manner of workmanship;
EXOD|35|32|And to devise curious works, to work in gold, and in silver, and in brass,
EXOD|35|33|And in the cutting of stones, to set them, and in carving of wood, to make any manner of cunning work.
EXOD|35|34|And he hath put in his heart that he may teach, both he, and Aholiab, the son of Ahisamach, of the tribe of Dan.
EXOD|35|35|Them hath he filled with wisdom of heart, to work all manner of work, of the engraver, and of the cunning workman, and of the embroiderer, in blue, and in purple, in scarlet, and in fine linen, and of the weaver, even of them that do any work, and of those that devise cunning work.
EXOD|36|1|Then wrought Bezaleel and Aholiab, and every wise hearted man, in whom the LORD put wisdom and understanding to know how to work all manner of work for the service of the sanctuary, according to all that the LORD had commanded.
EXOD|36|2|And Moses called Bezaleel and Aholiab, and every wise hearted man, in whose heart the LORD had put wisdom, even every one whose heart stirred him up to come unto the work to do it:
EXOD|36|3|And they received of Moses all the offering, which the children of Israel had brought for the work of the service of the sanctuary, to make it withal. And they brought yet unto him free offerings every morning.
EXOD|36|4|And all the wise men, that wrought all the work of the sanctuary, came every man from his work which they made;
EXOD|36|5|And they spake unto Moses, saying, The people bring much more than enough for the service of the work, which the LORD commanded to make.
EXOD|36|6|And Moses gave commandment, and they caused it to be proclaimed throughout the camp, saying, Let neither man nor woman make any more work for the offering of the sanctuary. So the people were restrained from bringing.
EXOD|36|7|For the stuff they had was sufficient for all the work to make it, and too much.
EXOD|36|8|And every wise hearted man among them that wrought the work of the tabernacle made ten curtains of fine twined linen, and blue, and purple, and scarlet: with cherubim of cunning work made he them.
EXOD|36|9|The length of one curtain was twenty and eight cubits, and the breadth of one curtain four cubits: the curtains were all of one size.
EXOD|36|10|And he coupled the five curtains one unto another: and the other five curtains he coupled one unto another.
EXOD|36|11|And he made loops of blue on the edge of one curtain from the selvedge in the coupling: likewise he made in the uttermost side of another curtain, in the coupling of the second.
EXOD|36|12|Fifty loops made he in one curtain, and fifty loops made he in the edge of the curtain which was in the coupling of the second: the loops held one curtain to another.
EXOD|36|13|And he made fifty taches of gold, and coupled the curtains one unto another with the taches: so it became one tabernacle.
EXOD|36|14|And he made curtains of goats' hair for the tent over the tabernacle: eleven curtains he made them.
EXOD|36|15|The length of one curtain was thirty cubits, and four cubits was the breadth of one curtain: the eleven curtains were of one size.
EXOD|36|16|And he coupled five curtains by themselves, and six curtains by themselves.
EXOD|36|17|And he made fifty loops upon the uttermost edge of the curtain in the coupling, and fifty loops made he upon the edge of the curtain which coupleth the second.
EXOD|36|18|And he made fifty taches of brass to couple the tent together, that it might be one.
EXOD|36|19|And he made a covering for the tent of rams' skins dyed red, and a covering of badgers' skins above that.
EXOD|36|20|And he made boards for the tabernacle of shittim wood, standing up.
EXOD|36|21|The length of a board was ten cubits, and the breadth of a board one cubit and a half.
EXOD|36|22|One board had two tenons, equally distant one from another: thus did he make for all the boards of the tabernacle.
EXOD|36|23|And he made boards for the tabernacle; twenty boards for the south side southward:
EXOD|36|24|And forty sockets of silver he made under the twenty boards; two sockets under one board for his two tenons, and two sockets under another board for his two tenons.
EXOD|36|25|And for the other side of the tabernacle, which is toward the north corner, he made twenty boards,
EXOD|36|26|And their forty sockets of silver; two sockets under one board, and two sockets under another board.
EXOD|36|27|And for the sides of the tabernacle westward he made six boards.
EXOD|36|28|And two boards made he for the corners of the tabernacle in the two sides.
EXOD|36|29|And they were coupled beneath, and coupled together at the head thereof, to one ring: thus he did to both of them in both the corners.
EXOD|36|30|And there were eight boards; and their sockets were sixteen sockets of silver, under every board two sockets.
EXOD|36|31|And he made bars of shittim wood; five for the boards of the one side of the tabernacle,
EXOD|36|32|And five bars for the boards of the other side of the tabernacle, and five bars for the boards of the tabernacle for the sides westward.
EXOD|36|33|And he made the middle bar to shoot through the boards from the one end to the other.
EXOD|36|34|And he overlaid the boards with gold, and made their rings of gold to be places for the bars, and overlaid the bars with gold.
EXOD|36|35|And he made a vail of blue, and purple, and scarlet, and fine twined linen: with cherubim made he it of cunning work.
EXOD|36|36|And he made thereunto four pillars of shittim wood, and overlaid them with gold: their hooks were of gold; and he cast for them four sockets of silver.
EXOD|36|37|And he made an hanging for the tabernacle door of blue, and purple, and scarlet, and fine twined linen, of needlework;
EXOD|36|38|And the five pillars of it with their hooks: and he overlaid their chapiters and their fillets with gold: but their five sockets were of brass.
EXOD|37|1|And Bezaleel made the ark of shittim wood: two cubits and a half was the length of it, and a cubit and a half the breadth of it, and a cubit and a half the height of it:
EXOD|37|2|And he overlaid it with pure gold within and without, and made a crown of gold to it round about.
EXOD|37|3|And he cast for it four rings of gold, to be set by the four corners of it; even two rings upon the one side of it, and two rings upon the other side of it.
EXOD|37|4|And he made staves of shittim wood, and overlaid them with gold.
EXOD|37|5|And he put the staves into the rings by the sides of the ark, to bear the ark.
EXOD|37|6|And he made the mercy seat of pure gold: two cubits and a half was the length thereof, and one cubit and a half the breadth thereof.
EXOD|37|7|And he made two cherubim of gold, beaten out of one piece made he them, on the two ends of the mercy seat;
EXOD|37|8|One cherub on the end on this side, and another cherub on the other end on that side: out of the mercy seat made he the cherubim on the two ends thereof.
EXOD|37|9|And the cherubim spread out their wings on high, and covered with their wings over the mercy seat, with their faces one to another; even to the mercy seatward were the faces of the cherubim.
EXOD|37|10|And he made the table of shittim wood: two cubits was the length thereof, and a cubit the breadth thereof, and a cubit and a half the height thereof:
EXOD|37|11|And he overlaid it with pure gold, and made thereunto a crown of gold round about.
EXOD|37|12|Also he made thereunto a border of an handbreadth round about; and made a crown of gold for the border thereof round about.
EXOD|37|13|And he cast for it four rings of gold, and put the rings upon the four corners that were in the four feet thereof.
EXOD|37|14|Over against the border were the rings, the places for the staves to bear the table.
EXOD|37|15|And he made the staves of shittim wood, and overlaid them with gold, to bear the table.
EXOD|37|16|And he made the vessels which were upon the table, his dishes, and his spoons, and his bowls, and his covers to cover withal, of pure gold.
EXOD|37|17|And he made the candlestick of pure gold: of beaten work made he the candlestick; his shaft, and his branch, his bowls, his knops, and his flowers, were of the same:
EXOD|37|18|And six branches going out of the sides thereof; three branches of the candlestick out of the one side thereof, and three branches of the candlestick out of the other side thereof:
EXOD|37|19|Three bowls made after the fashion of almonds in one branch, a knop and a flower; and three bowls made like almonds in another branch, a knop and a flower: so throughout the six branches going out of the candlestick.
EXOD|37|20|And in the candlestick were four bowls made like almonds, his knops, and his flowers:
EXOD|37|21|And a knop under two branches of the same, and a knop under two branches of the same, and a knop under two branches of the same, according to the six branches going out of it.
EXOD|37|22|Their knops and their branches were of the same: all of it was one beaten work of pure gold.
EXOD|37|23|And he made his seven lamps, and his snuffers, and his snuffdishes, of pure gold.
EXOD|37|24|Of a talent of pure gold made he it, and all the vessels thereof.
EXOD|37|25|And he made the incense altar of shittim wood: the length of it was a cubit, and the breadth of it a cubit; it was foursquare; and two cubits was the height of it; the horns thereof were of the same.
EXOD|37|26|And he overlaid it with pure gold, both the top of it, and the sides thereof round about, and the horns of it: also he made unto it a crown of gold round about.
EXOD|37|27|And he made two rings of gold for it under the crown thereof, by the two corners of it, upon the two sides thereof, to be places for the staves to bear it withal.
EXOD|37|28|And he made the staves of shittim wood, and overlaid them with gold.
EXOD|37|29|And he made the holy anointing oil, and the pure incense of sweet spices, according to the work of the apothecary.
EXOD|38|1|And he made the altar of burnt offering of shittim wood: five cubits was the length thereof, and five cubits the breadth thereof; it was foursquare; and three cubits the height thereof.
EXOD|38|2|And he made the horns thereof on the four corners of it; the horns thereof were of the same: and he overlaid it with brass.
EXOD|38|3|And he made all the vessels of the altar, the pots, and the shovels, and the basins, and the fleshhooks, and the firepans: all the vessels thereof made he of brass.
EXOD|38|4|And he made for the altar a brazen grate of network under the compass thereof beneath unto the midst of it.
EXOD|38|5|And he cast four rings for the four ends of the grate of brass, to be places for the staves.
EXOD|38|6|And he made the staves of shittim wood, and overlaid them with brass.
EXOD|38|7|And he put the staves into the rings on the sides of the altar, to bear it withal; he made the altar hollow with boards.
EXOD|38|8|And he made the laver of brass, and the foot of it of brass, of the lookingglasses of the women assembling, which assembled at the door of the tabernacle of the congregation.
EXOD|38|9|And he made the court: on the south side southward the hangings of the court were of fine twined linen, an hundred cubits:
EXOD|38|10|Their pillars were twenty, and their brazen sockets twenty; the hooks of the pillars and their fillets were of silver.
EXOD|38|11|And for the north side the hangings were an hundred cubits, their pillars were twenty, and their sockets of brass twenty; the hooks of the pillars and their fillets of silver.
EXOD|38|12|And for the west side were hangings of fifty cubits, their pillars ten, and their sockets ten; the hooks of the pillars and their fillets of silver.
EXOD|38|13|And for the east side eastward fifty cubits.
EXOD|38|14|The hangings of the one side of the gate were fifteen cubits; their pillars three, and their sockets three.
EXOD|38|15|And for the other side of the court gate, on this hand and that hand, were hangings of fifteen cubits; their pillars three, and their sockets three.
EXOD|38|16|All the hangings of the court round about were of fine twined linen.
EXOD|38|17|And the sockets for the pillars were of brass; the hooks of the pillars and their fillets of silver; and the overlaying of their chapiters of silver; and all the pillars of the court were filleted with silver.
EXOD|38|18|And the hanging for the gate of the court was needlework, of blue, and purple, and scarlet, and fine twined linen: and twenty cubits was the length, and the height in the breadth was five cubits, answerable to the hangings of the court.
EXOD|38|19|And their pillars were four, and their sockets of brass four; their hooks of silver, and the overlaying of their chapiters and their fillets of silver.
EXOD|38|20|And all the pins of the tabernacle, and of the court round about, were of brass.
EXOD|38|21|This is the sum of the tabernacle, even of the tabernacle of testimony, as it was counted, according to the commandment of Moses, for the service of the Levites, by the hand of Ithamar, son to Aaron the priest.
EXOD|38|22|And Bezaleel the son Uri, the son of Hur, of the tribe of Judah, made all that the LORD commanded Moses.
EXOD|38|23|And with him was Aholiab, son of Ahisamach, of the tribe of Dan, an engraver, and a cunning workman, and an embroiderer in blue, and in purple, and in scarlet, and fine linen.
EXOD|38|24|All the gold that was occupied for the work in all the work of the holy place, even the gold of the offering, was twenty and nine talents, and seven hundred and thirty shekels, after the shekel of the sanctuary.
EXOD|38|25|And the silver of them that were numbered of the congregation was an hundred talents, and a thousand seven hundred and threescore and fifteen shekels, after the shekel of the sanctuary:
EXOD|38|26|A bekah for every man, that is, half a shekel, after the shekel of the sanctuary, for every one that went to be numbered, from twenty years old and upward, for six hundred thousand and three thousand and five hundred and fifty men.
EXOD|38|27|And of the hundred talents of silver were cast the sockets of the sanctuary, and the sockets of the vail; an hundred sockets of the hundred talents, a talent for a socket.
EXOD|38|28|And of the thousand seven hundred seventy and five shekels he made hooks for the pillars, and overlaid their chapiters, and filleted them.
EXOD|38|29|And the brass of the offering was seventy talents, and two thousand and four hundred shekels.
EXOD|38|30|And therewith he made the sockets to the door of the tabernacle of the congregation, and the brazen altar, and the brazen grate for it, and all the vessels of the altar,
EXOD|38|31|And the sockets of the court round about, and the sockets of the court gate, and all the pins of the tabernacle, and all the pins of the court round about.
EXOD|39|1|And of the blue, and purple, and scarlet, they made cloths of service, to do service in the holy place, and made the holy garments for Aaron; as the LORD commanded Moses.
EXOD|39|2|And he made the ephod of gold, blue, and purple, and scarlet, and fine twined linen.
EXOD|39|3|And they did beat the gold into thin plates, and cut it into wires, to work it in the blue, and in the purple, and in the scarlet, and in the fine linen, with cunning work.
EXOD|39|4|They made shoulderpieces for it, to couple it together: by the two edges was it coupled together.
EXOD|39|5|And the curious girdle of his ephod, that was upon it, was of the same, according to the work thereof; of gold, blue, and purple, and scarlet, and fine twined linen; as the LORD commanded Moses.
EXOD|39|6|And they wrought onyx stones inclosed in ouches of gold, graven, as signets are graven, with the names of the children of Israel.
EXOD|39|7|And he put them on the shoulders of the ephod, that they should be stones for a memorial to the children of Israel; as the LORD commanded Moses.
EXOD|39|8|And he made the breastplate of cunning work, like the work of the ephod; of gold, blue, and purple, and scarlet, and fine twined linen.
EXOD|39|9|It was foursquare; they made the breastplate double: a span was the length thereof, and a span the breadth thereof, being doubled.
EXOD|39|10|And they set in it four rows of stones: the first row was a sardius, a topaz, and a carbuncle: this was the first row.
EXOD|39|11|And the second row, an emerald, a sapphire, and a diamond.
EXOD|39|12|And the third row, a ligure, an agate, and an amethyst.
EXOD|39|13|And the fourth row, a beryl, an onyx, and a jasper: they were inclosed in ouches of gold in their inclosings.
EXOD|39|14|And the stones were according to the names of the children of Israel, twelve, according to their names, like the engravings of a signet, every one with his name, according to the twelve tribes.
EXOD|39|15|And they made upon the breastplate chains at the ends, of wreathed work of pure gold.
EXOD|39|16|And they made two ouches of gold, and two gold rings; and put the two rings in the two ends of the breastplate.
EXOD|39|17|And they put the two wreathed chains of gold in the two rings on the ends of the breastplate.
EXOD|39|18|And the two ends of the two wreathed chains they fastened in the two ouches, and put them on the shoulderpieces of the ephod, before it.
EXOD|39|19|And they made two rings of gold, and put them on the two ends of the breastplate, upon the border of it, which was on the side of the ephod inward.
EXOD|39|20|And they made two other golden rings, and put them on the two sides of the ephod underneath, toward the forepart of it, over against the other coupling thereof, above the curious girdle of the ephod.
EXOD|39|21|And they did bind the breastplate by his rings unto the rings of the ephod with a lace of blue, that it might be above the curious girdle of the ephod, and that the breastplate might not be loosed from the ephod; as the LORD commanded Moses.
EXOD|39|22|And he made the robe of the ephod of woven work, all of blue.
EXOD|39|23|And there was an hole in the midst of the robe, as the hole of an habergeon, with a band round about the hole, that it should not rend.
EXOD|39|24|And they made upon the hems of the robe pomegranates of blue, and purple, and scarlet, and twined linen.
EXOD|39|25|And they made bells of pure gold, and put the bells between the pomegranates upon the hem of the robe, round about between the pomegranates;
EXOD|39|26|A bell and a pomegranate, a bell and a pomegranate, round about the hem of the robe to minister in; as the LORD commanded Moses.
EXOD|39|27|And they made coats of fine linen of woven work for Aaron, and for his sons,
EXOD|39|28|And a mitre of fine linen, and goodly bonnets of fine linen, and linen breeches of fine twined linen,
EXOD|39|29|And a girdle of fine twined linen, and blue, and purple, and scarlet, of needlework; as the LORD commanded Moses.
EXOD|39|30|And they made the plate of the holy crown of pure gold, and wrote upon it a writing, like to the engravings of a signet, HOLINESS TO THE LORD.
EXOD|39|31|And they tied unto it a lace of blue, to fasten it on high upon the mitre; as the LORD commanded Moses.
EXOD|39|32|Thus was all the work of the tabernacle of the tent of the congregation finished: and the children of Israel did according to all that the LORD commanded Moses, so did they.
EXOD|39|33|And they brought the tabernacle unto Moses, the tent, and all his furniture, his taches, his boards, his bars, and his pillars, and his sockets,
EXOD|39|34|And the covering of rams' skins dyed red, and the covering of badgers' skins, and the vail of the covering,
EXOD|39|35|The ark of the testimony, and the staves thereof, and the mercy seat,
EXOD|39|36|The table, and all the vessels thereof, and the showbread,
EXOD|39|37|The pure candlestick, with the lamps thereof, even with the lamps to be set in order, and all the vessels thereof, and the oil for light,
EXOD|39|38|And the golden altar, and the anointing oil, and the sweet incense, and the hanging for the tabernacle door,
EXOD|39|39|The brazen altar, and his grate of brass, his staves, and all his vessels, the laver and his foot,
EXOD|39|40|The hangings of the court, his pillars, and his sockets, and the hanging for the court gate, his cords, and his pins, and all the vessels of the service of the tabernacle, for the tent of the congregation,
EXOD|39|41|The cloths of service to do service in the holy place, and the holy garments for Aaron the priest, and his sons' garments, to minister in the priest's office.
EXOD|39|42|According to all that the LORD commanded Moses, so the children of Israel made all the work.
EXOD|39|43|And Moses did look upon all the work, and, behold, they had done it as the LORD had commanded, even so had they done it: and Moses blessed them.
EXOD|40|1|And the LORD spake unto Moses, saying,
EXOD|40|2|On the first day of the first month shalt thou set up the tabernacle of the tent of the congregation.
EXOD|40|3|And thou shalt put therein the ark of the testimony, and cover the ark with the vail.
EXOD|40|4|And thou shalt bring in the table, and set in order the things that are to be set in order upon it; and thou shalt bring in the candlestick, and light the lamps thereof.
EXOD|40|5|And thou shalt set the altar of gold for the incense before the ark of the testimony, and put the hanging of the door to the tabernacle.
EXOD|40|6|And thou shalt set the altar of the burnt offering before the door of the tabernacle of the tent of the congregation.
EXOD|40|7|And thou shalt set the laver between the tent of the congregation and the altar, and shalt put water therein.
EXOD|40|8|And thou shalt set up the court round about, and hang up the hanging at the court gate.
EXOD|40|9|And thou shalt take the anointing oil, and anoint the tabernacle, and all that is therein, and shalt hallow it, and all the vessels thereof: and it shall be holy.
EXOD|40|10|And thou shalt anoint the altar of the burnt offering, and all his vessels, and sanctify the altar: and it shall be an altar most holy.
EXOD|40|11|And thou shalt anoint the laver and his foot, and sanctify it.
EXOD|40|12|And thou shalt bring Aaron and his sons unto the door of the tabernacle of the congregation, and wash them with water.
EXOD|40|13|And thou shalt put upon Aaron the holy garments, and anoint him, and sanctify him; that he may minister unto me in the priest's office.
EXOD|40|14|And thou shalt bring his sons, and clothe them with coats:
EXOD|40|15|And thou shalt anoint them, as thou didst anoint their father, that they may minister unto me in the priest's office: for their anointing shall surely be an everlasting priesthood throughout their generations.
EXOD|40|16|Thus did Moses: according to all that the LORD commanded him, so did he.
EXOD|40|17|And it came to pass in the first month in the second year, on the first day of the month, that the tabernacle was reared up.
EXOD|40|18|And Moses reared up the tabernacle, and fastened his sockets, and set up the boards thereof, and put in the bars thereof, and reared up his pillars.
EXOD|40|19|And he spread abroad the tent over the tabernacle, and put the covering of the tent above upon it; as the LORD commanded Moses.
EXOD|40|20|And he took and put the testimony into the ark, and set the staves on the ark, and put the mercy seat above upon the ark:
EXOD|40|21|And he brought the ark into the tabernacle, and set up the vail of the covering, and covered the ark of the testimony; as the LORD commanded Moses.
EXOD|40|22|And he put the table in the tent of the congregation, upon the side of the tabernacle northward, without the vail.
EXOD|40|23|And he set the bread in order upon it before the LORD; as the LORD had commanded Moses.
EXOD|40|24|And he put the candlestick in the tent of the congregation, over against the table, on the side of the tabernacle southward.
EXOD|40|25|And he lighted the lamps before the LORD; as the LORD commanded Moses.
EXOD|40|26|And he put the golden altar in the tent of the congregation before the vail:
EXOD|40|27|And he burnt sweet incense thereon; as the LORD commanded Moses.
EXOD|40|28|And he set up the hanging at the door of the tabernacle.
EXOD|40|29|And he put the altar of burnt offering by the door of the tabernacle of the tent of the congregation, and offered upon it the burnt offering and the meat offering; as the LORD commanded Moses.
EXOD|40|30|And he set the laver between the tent of the congregation and the altar, and put water there, to wash withal.
EXOD|40|31|And Moses and Aaron and his sons washed their hands and their feet thereat:
EXOD|40|32|When they went into the tent of the congregation, and when they came near unto the altar, they washed; as the LORD commanded Moses.
EXOD|40|33|And he reared up the court round about the tabernacle and the altar, and set up the hanging of the court gate. So Moses finished the work.
EXOD|40|34|Then a cloud covered the tent of the congregation, and the glory of the LORD filled the tabernacle.
EXOD|40|35|And Moses was not able to enter into the tent of the congregation, because the cloud abode thereon, and the glory of the LORD filled the tabernacle.
EXOD|40|36|And when the cloud was taken up from over the tabernacle, the children of Israel went onward in all their journeys:
EXOD|40|37|But if the cloud were not taken up, then they journeyed not till the day that it was taken up.
EXOD|40|38|For the cloud of the LORD was upon the tabernacle by day, and fire was on it by night, in the sight of all the house of Israel, throughout all their journeys.
