PHIL|1|1|Paul and Timotheus, the servants of Jesus Christ, to all the saints in Christ Jesus which are at Philippi, with the bishops and deacons:
PHIL|1|2|Grace be unto you, and peace, from God our Father, and from the Lord Jesus Christ.
PHIL|1|3|I thank my God upon every remembrance of you,
PHIL|1|4|Always in every prayer of mine for you all making request with joy,
PHIL|1|5|For your fellowship in the gospel from the first day until now;
PHIL|1|6|Being confident of this very thing, that he which hath begun a good work in you will perform it until the day of Jesus Christ:
PHIL|1|7|Even as it is meet for me to think this of you all, because I have you in my heart; inasmuch as both in my bonds, and in the defence and confirmation of the gospel, ye all are partakers of my grace.
PHIL|1|8|For God is my record, how greatly I long after you all in the bowels of Jesus Christ.
PHIL|1|9|And this I pray, that your love may abound yet more and more in knowledge and in all judgment;
PHIL|1|10|That ye may approve things that are excellent; that ye may be sincere and without offence till the day of Christ.
PHIL|1|11|Being filled with the fruits of righteousness, which are by Jesus Christ, unto the glory and praise of God.
PHIL|1|12|But I would ye should understand, brethren, that the things which happened unto me have fallen out rather unto the furtherance of the gospel;
PHIL|1|13|So that my bonds in Christ are manifest in all the palace, and in all other places;
PHIL|1|14|And many of the brethren in the Lord, waxing confident by my bonds, are much more bold to speak the word without fear.
PHIL|1|15|Some indeed preach Christ even of envy and strife; and some also of good will:
PHIL|1|16|The one preach Christ of contention, not sincerely, supposing to add affliction to my bonds:
PHIL|1|17|But the other of love, knowing that I am set for the defence of the gospel.
PHIL|1|18|What then? notwithstanding, every way, whether in pretence, or in truth, Christ is preached; and I therein do rejoice, yea, and will rejoice.
PHIL|1|19|For I know that this shall turn to my salvation through your prayer, and the supply of the Spirit of Jesus Christ,
PHIL|1|20|According to my earnest expectation and my hope, that in nothing I shall be ashamed, but that with all boldness, as always, so now also Christ shall be magnified in my body, whether it be by life, or by death.
PHIL|1|21|For to me to live is Christ, and to die is gain.
PHIL|1|22|But if I live in the flesh, this is the fruit of my labour: yet what I shall choose I wot not.
PHIL|1|23|For I am in a strait betwixt two, having a desire to depart, and to be with Christ; which is far better:
PHIL|1|24|Nevertheless to abide in the flesh is more needful for you.
PHIL|1|25|And having this confidence, I know that I shall abide and continue with you all for your furtherance and joy of faith;
PHIL|1|26|That your rejoicing may be more abundant in Jesus Christ for me by my coming to you again.
PHIL|1|27|Only let your conversation be as it becometh the gospel of Christ: that whether I come and see you, or else be absent, I may hear of your affairs, that ye stand fast in one spirit, with one mind striving together for the faith of the gospel;
PHIL|1|28|And in nothing terrified by your adversaries: which is to them an evident token of perdition, but to you of salvation, and that of God.
PHIL|1|29|For unto you it is given in the behalf of Christ, not only to believe on him, but also to suffer for his sake;
PHIL|1|30|Having the same conflict which ye saw in me, and now hear to be in me.
PHIL|2|1|If there be therefore any consolation in Christ, if any comfort of love, if any fellowship of the Spirit, if any bowels and mercies,
PHIL|2|2|Fulfil ye my joy, that ye be likeminded, having the same love, being of one accord, of one mind.
PHIL|2|3|Let nothing be done through strife or vainglory; but in lowliness of mind let each esteem other better than themselves.
PHIL|2|4|Look not every man on his own things, but every man also on the things of others.
PHIL|2|5|Let this mind be in you, which was also in Christ Jesus:
PHIL|2|6|Who, being in the form of God, thought it not robbery to be equal with God:
PHIL|2|7|But made himself of no reputation, and took upon him the form of a servant, and was made in the likeness of men:
PHIL|2|8|And being found in fashion as a man, he humbled himself, and became obedient unto death, even the death of the cross.
PHIL|2|9|Wherefore God also hath highly exalted him, and given him a name which is above every name:
PHIL|2|10|That at the name of Jesus every knee should bow, of things in heaven, and things in earth, and things under the earth;
PHIL|2|11|And that every tongue should confess that Jesus Christ is Lord, to the glory of God the Father.
PHIL|2|12|Wherefore, my beloved, as ye have always obeyed, not as in my presence only, but now much more in my absence, work out your own salvation with fear and trembling.
PHIL|2|13|For it is God which worketh in you both to will and to do of his good pleasure.
PHIL|2|14|Do all things without murmurings and disputings:
PHIL|2|15|That ye may be blameless and harmless, the sons of God, without rebuke, in the midst of a crooked and perverse nation, among whom ye shine as lights in the world;
PHIL|2|16|Holding forth the word of life; that I may rejoice in the day of Christ, that I have not run in vain, neither laboured in vain.
PHIL|2|17|Yea, and if I be offered upon the sacrifice and service of your faith, I joy, and rejoice with you all.
PHIL|2|18|For the same cause also do ye joy, and rejoice with me.
PHIL|2|19|But I trust in the Lord Jesus to send Timotheus shortly unto you, that I also may be of good comfort, when I know your state.
PHIL|2|20|For I have no man likeminded, who will naturally care for your state.
PHIL|2|21|For all seek their own, not the things which are Jesus Christ's.
PHIL|2|22|But ye know the proof of him, that, as a son with the father, he hath served with me in the gospel.
PHIL|2|23|Him therefore I hope to send presently, so soon as I shall see how it will go with me.
PHIL|2|24|But I trust in the Lord that I also myself shall come shortly.
PHIL|2|25|Yet I supposed it necessary to send to you Epaphroditus, my brother, and companion in labour, and fellowsoldier, but your messenger, and he that ministered to my wants.
PHIL|2|26|For he longed after you all, and was full of heaviness, because that ye had heard that he had been sick.
PHIL|2|27|For indeed he was sick nigh unto death: but God had mercy on him; and not on him only, but on me also, lest I should have sorrow upon sorrow.
PHIL|2|28|I sent him therefore the more carefully, that, when ye see him again, ye may rejoice, and that I may be the less sorrowful.
PHIL|2|29|Receive him therefore in the Lord with all gladness; and hold such in reputation:
PHIL|2|30|Because for the work of Christ he was nigh unto death, not regarding his life, to supply your lack of service toward me.
PHIL|3|1|Finally, my brethren, rejoice in the Lord. To write the same things to you, to me indeed is not grievous, but for you it is safe.
PHIL|3|2|Beware of dogs, beware of evil workers, beware of the concision.
PHIL|3|3|For we are the circumcision, which worship God in the spirit, and rejoice in Christ Jesus, and have no confidence in the flesh.
PHIL|3|4|Though I might also have confidence in the flesh. If any other man thinketh that he hath whereof he might trust in the flesh, I more:
PHIL|3|5|Circumcised the eighth day, of the stock of Israel, of the tribe of Benjamin, an Hebrew of the Hebrews; as touching the law, a Pharisee;
PHIL|3|6|Concerning zeal, persecuting the church; touching the righteousness which is in the law, blameless.
PHIL|3|7|But what things were gain to me, those I counted loss for Christ.
PHIL|3|8|Yea doubtless, and I count all things but loss for the excellency of the knowledge of Christ Jesus my Lord: for whom I have suffered the loss of all things, and do count them but dung, that I may win Christ,
PHIL|3|9|And be found in him, not having mine own righteousness, which is of the law, but that which is through the faith of Christ, the righteousness which is of God by faith:
PHIL|3|10|That I may know him, and the power of his resurrection, and the fellowship of his sufferings, being made conformable unto his death;
PHIL|3|11|If by any means I might attain unto the resurrection of the dead.
PHIL|3|12|Not as though I had already attained, either were already perfect: but I follow after, if that I may apprehend that for which also I am apprehended of Christ Jesus.
PHIL|3|13|Brethren, I count not myself to have apprehended: but this one thing I do, forgetting those things which are behind, and reaching forth unto those things which are before,
PHIL|3|14|I press toward the mark for the prize of the high calling of God in Christ Jesus.
PHIL|3|15|Let us therefore, as many as be perfect, be thus minded: and if in any thing ye be otherwise minded, God shall reveal even this unto you.
PHIL|3|16|Nevertheless, whereto we have already attained, let us walk by the same rule, let us mind the same thing.
PHIL|3|17|Brethren, be followers together of me, and mark them which walk so as ye have us for an ensample.
PHIL|3|18|(For many walk, of whom I have told you often, and now tell you even weeping, that they are the enemies of the cross of Christ:
PHIL|3|19|Whose end is destruction, whose God is their belly, and whose glory is in their shame, who mind earthly things.)
PHIL|3|20|For our conversation is in heaven; from whence also we look for the Saviour, the Lord Jesus Christ:
PHIL|3|21|Who shall change our vile body, that it may be fashioned like unto his glorious body, according to the working whereby he is able even to subdue all things unto himself.
PHIL|4|1|Therefore, my brethren dearly beloved and longed for, my joy and crown, so stand fast in the Lord, my dearly beloved.
PHIL|4|2|I beseech Euodias, and beseech Syntyche, that they be of the same mind in the Lord.
PHIL|4|3|And I intreat thee also, true yokefellow, help those women which laboured with me in the gospel, with Clement also, and with other my fellowlabourers, whose names are in the book of life.
PHIL|4|4|Rejoice in the Lord alway: and again I say, Rejoice.
PHIL|4|5|Let your moderation be known unto all men. The Lord is at hand.
PHIL|4|6|Be careful for nothing; but in every thing by prayer and supplication with thanksgiving let your requests be made known unto God.
PHIL|4|7|And the peace of God, which passeth all understanding, shall keep your hearts and minds through Christ Jesus.
PHIL|4|8|Finally, brethren, whatsoever things are true, whatsoever things are honest, whatsoever things are just, whatsoever things are pure, whatsoever things are lovely, whatsoever things are of good report; if there be any virtue, and if there be any praise, think on these things.
PHIL|4|9|Those things, which ye have both learned, and received, and heard, and seen in me, do: and the God of peace shall be with you.
PHIL|4|10|But I rejoiced in the Lord greatly, that now at the last your care of me hath flourished again; wherein ye were also careful, but ye lacked opportunity.
PHIL|4|11|Not that I speak in respect of want: for I have learned, in whatsoever state I am, therewith to be content.
PHIL|4|12|I know both how to be abased, and I know how to abound: every where and in all things I am instructed both to be full and to be hungry, both to abound and to suffer need.
PHIL|4|13|I can do all things through Christ which strengtheneth me.
PHIL|4|14|Notwithstanding ye have well done, that ye did communicate with my affliction.
PHIL|4|15|Now ye Philippians know also, that in the beginning of the gospel, when I departed from Macedonia, no church communicated with me as concerning giving and receiving, but ye only.
PHIL|4|16|For even in Thessalonica ye sent once and again unto my necessity.
PHIL|4|17|Not because I desire a gift: but I desire fruit that may abound to your account.
PHIL|4|18|But I have all, and abound: I am full, having received of Epaphroditus the things which were sent from you, an odour of a sweet smell, a sacrifice acceptable, wellpleasing to God.
PHIL|4|19|But my God shall supply all your need according to his riches in glory by Christ Jesus.
PHIL|4|20|Now unto God and our Father be glory for ever and ever. Amen.
PHIL|4|21|Salute every saint in Christ Jesus. The brethren which are with me greet you.
PHIL|4|22|All the saints salute you, chiefly they that are of Caesar's household.
PHIL|4|23|The grace of our Lord Jesus Christ be with you all. Amen.
