ZEPH|1|1|The word of the LORD that came to Zephaniah son of Cushi, the son of Gedaliah, the son of Amariah, the son of Hezekiah, during the reign of Josiah son of Amon king of Judah:
ZEPH|1|2|"I will sweep away everything from the face of the earth," declares the LORD.
ZEPH|1|3|"I will sweep away both men and animals; I will sweep away the birds of the air and the fish of the sea. The wicked will have only heaps of rubble when I cut off man from the face of the earth," declares the LORD.
ZEPH|1|4|"I will stretch out my hand against Judah and against all who live in Jerusalem. I will cut off from this place every remnant of Baal, the names of the pagan and the idolatrous priests-
ZEPH|1|5|those who bow down on the roofs to worship the starry host, those who bow down and swear by the LORD and who also swear by Molech,
ZEPH|1|6|those who turn back from following the LORD and neither seek the LORD nor inquire of him.
ZEPH|1|7|Be silent before the Sovereign LORD, for the day of the LORD is near. The LORD has prepared a sacrifice; he has consecrated those he has invited.
ZEPH|1|8|On the day of the LORD's sacrifice I will punish the princes and the king's sons and all those clad in foreign clothes.
ZEPH|1|9|On that day I will punish all who avoid stepping on the threshold, who fill the temple of their gods with violence and deceit.
ZEPH|1|10|"On that day," declares the LORD, "a cry will go up from the Fish Gate, wailing from the New Quarter, and a loud crash from the hills.
ZEPH|1|11|Wail, you who live in the market district; all your merchants will be wiped out, all who trade with silver will be ruined.
ZEPH|1|12|At that time I will search Jerusalem with lamps and punish those who are complacent, who are like wine left on its dregs, who think, 'The LORD will do nothing, either good or bad.'
ZEPH|1|13|Their wealth will be plundered, their houses demolished. They will build houses but not live in them; they will plant vineyards but not drink the wine.
ZEPH|1|14|"The great day of the LORD is near- near and coming quickly. Listen! The cry on the day of the LORD will be bitter, the shouting of the warrior there.
ZEPH|1|15|That day will be a day of wrath, a day of distress and anguish, a day of trouble and ruin, a day of darkness and gloom, a day of clouds and blackness,
ZEPH|1|16|a day of trumpet and battle cry against the fortified cities and against the corner towers.
ZEPH|1|17|I will bring distress on the people and they will walk like blind men, because they have sinned against the LORD. Their blood will be poured out like dust and their entrails like filth.
ZEPH|1|18|Neither their silver nor their gold will be able to save them on the day of the LORD's wrath. In the fire of his jealousy the whole world will be consumed, for he will make a sudden end of all who live in the earth."
ZEPH|2|1|Gather together, gather together, O shameful nation,
ZEPH|2|2|before the appointed time arrives and that day sweeps on like chaff, before the fierce anger of the LORD comes upon you, before the day of the LORD's wrath comes upon you.
ZEPH|2|3|Seek the LORD, all you humble of the land, you who do what he commands. Seek righteousness, seek humility; perhaps you will be sheltered on the day of the LORD's anger.
ZEPH|2|4|Gaza will be abandoned and Ashkelon left in ruins. At midday Ashdod will be emptied and Ekron uprooted.
ZEPH|2|5|Woe to you who live by the sea, O Kerethite people; the word of the LORD is against you, O Canaan, land of the Philistines. "I will destroy you, and none will be left."
ZEPH|2|6|The land by the sea, where the Kerethites dwell, will be a place for shepherds and sheep pens.
ZEPH|2|7|It will belong to the remnant of the house of Judah; there they will find pasture. In the evening they will lie down in the houses of Ashkelon. The LORD their God will care for them; he will restore their fortunes.
ZEPH|2|8|"I have heard the insults of Moab and the taunts of the Ammonites, who insulted my people and made threats against their land.
ZEPH|2|9|Therefore, as surely as I live," declares the LORD Almighty, the God of Israel, "surely Moab will become like Sodom, the Ammonites like Gomorrah- a place of weeds and salt pits, a wasteland forever. The remnant of my people will plunder them; the survivors of my nation will inherit their land."
ZEPH|2|10|This is what they will get in return for their pride, for insulting and mocking the people of the LORD Almighty.
ZEPH|2|11|The LORD will be awesome to them when he destroys all the gods of the land. The nations on every shore will worship him, every one in its own land.
ZEPH|2|12|"You too, O Cushites, will be slain by my sword."
ZEPH|2|13|He will stretch out his hand against the north and destroy Assyria, leaving Nineveh utterly desolate and dry as the desert.
ZEPH|2|14|Flocks and herds will lie down there, creatures of every kind. The desert owl and the screech owl will roost on her columns. Their calls will echo through the windows, rubble will be in the doorways, the beams of cedar will be exposed.
ZEPH|2|15|This is the carefree city that lived in safety. She said to herself, "I am, and there is none besides me." What a ruin she has become, a lair for wild beasts! All who pass by her scoff and shake their fists.
ZEPH|3|1|Woe to the city of oppressors, rebellious and defiled!
ZEPH|3|2|She obeys no one, she accepts no correction. She does not trust in the LORD, she does not draw near to her God.
ZEPH|3|3|Her officials are roaring lions, her rulers are evening wolves, who leave nothing for the morning.
ZEPH|3|4|Her prophets are arrogant; they are treacherous men. Her priests profane the sanctuary and do violence to the law.
ZEPH|3|5|The LORD within her is righteous; he does no wrong. Morning by morning he dispenses his justice, and every new day he does not fail, yet the unrighteous know no shame.
ZEPH|3|6|"I have cut off nations; their strongholds are demolished. I have left their streets deserted, with no one passing through. Their cities are destroyed; no one will be left-no one at all.
ZEPH|3|7|I said to the city, 'Surely you will fear me and accept correction!' Then her dwelling would not be cut off, nor all my punishments come upon her. But they were still eager to act corruptly in all they did.
ZEPH|3|8|Therefore wait for me," declares the LORD, "for the day I will stand up to testify. I have decided to assemble the nations, to gather the kingdoms and to pour out my wrath on them- all my fierce anger. The whole world will be consumed by the fire of my jealous anger.
ZEPH|3|9|"Then will I purify the lips of the peoples, that all of them may call on the name of the LORD and serve him shoulder to shoulder.
ZEPH|3|10|From beyond the rivers of Cush my worshipers, my scattered people, will bring me offerings.
ZEPH|3|11|On that day you will not be put to shame for all the wrongs you have done to me, because I will remove from this city those who rejoice in their pride. Never again will you be haughty on my holy hill.
ZEPH|3|12|But I will leave within you the meek and humble, who trust in the name of the LORD.
ZEPH|3|13|The remnant of Israel will do no wrong; they will speak no lies, nor will deceit be found in their mouths. They will eat and lie down and no one will make them afraid."
ZEPH|3|14|Sing, O Daughter of Zion; shout aloud, O Israel! Be glad and rejoice with all your heart, O Daughter of Jerusalem!
ZEPH|3|15|The LORD has taken away your punishment, he has turned back your enemy. The LORD, the King of Israel, is with you; never again will you fear any harm.
ZEPH|3|16|On that day they will say to Jerusalem, "Do not fear, O Zion; do not let your hands hang limp.
ZEPH|3|17|The LORD your God is with you, he is mighty to save. He will take great delight in you, he will quiet you with his love, he will rejoice over you with singing."
ZEPH|3|18|"The sorrows for the appointed feasts I will remove from you; they are a burden and a reproach to you.
ZEPH|3|19|At that time I will deal with all who oppressed you; I will rescue the lame and gather those who have been scattered. I will give them praise and honor in every land where they were put to shame.
ZEPH|3|20|At that time I will gather you; at that time I will bring you home. I will give you honor and praise among all the peoples of the earth when I restore your fortunes before your very eyes," says the LORD.
