1SAM|1|1|There was a certain man of Ramathaim-zophim of the hill country of Ephraim whose name was Elkanah the son of Jeroham, son of Elihu, son of Tohu, son of Zuph, an Ephrathite.
1SAM|1|2|He had two wives. The name of the one was Hannah, and the name of the other, Peninnah. And Peninnah had children, but Hannah had no children.
1SAM|1|3|Now this man used to go up year by year from his city to worship and to sacrifice to the LORD of hosts at Shiloh, where the two sons of Eli, Hophni and Phinehas, were priests of the LORD.
1SAM|1|4|On the day when Elkanah sacrificed, he would give portions to Peninnah his wife and to all her sons and daughters.
1SAM|1|5|But to Hannah he gave a double portion, because he loved her, though the LORD had closed her womb.
1SAM|1|6|And her rival used to provoke her grievously to irritate her, because the LORD had closed her womb.
1SAM|1|7|So it went on year by year. As often as she went up to the house of the LORD, she used to provoke her. Therefore Hannah wept and would not eat.
1SAM|1|8|And Elkanah, her husband, said to her, "Hannah, why do you weep? And why do you not eat? And why is your heart sad? Am I not more to you than ten sons?"
1SAM|1|9|After they had eaten and drunk in Shiloh, Hannah rose. Now Eli the priest was sitting on the seat beside the doorpost of the temple of the LORD.
1SAM|1|10|She was deeply distressed and prayed to the LORD and wept bitterly.
1SAM|1|11|And she vowed a vow and said, "O LORD of hosts, if you will indeed look on the affliction of your servant and remember me and not forget your servant, but will give to your servant a son, then I will give him to the LORD all the days of his life, and no razor shall touch his head."
1SAM|1|12|As she continued praying before the LORD, Eli observed her mouth.
1SAM|1|13|Hannah was speaking in her heart; only her lips moved, and her voice was not heard. Therefore Eli took her to be a drunken woman.
1SAM|1|14|And Eli said to her, "How long will you go on being drunk? Put away your wine from you."
1SAM|1|15|But Hannah answered, "No, my lord, I am a woman troubled in spirit. I have drunk neither wine nor strong drink, but I have been pouring out my soul before the LORD.
1SAM|1|16|Do not regard your servant as a worthless woman, for all along I have been speaking out of my great anxiety and vexation."
1SAM|1|17|Then Eli answered, "Go in peace, and the God of Israel grant your petition that you have made to him."
1SAM|1|18|And she said, "Let your servant find favor in your eyes." Then the woman went her way and ate, and her face was no longer sad.
1SAM|1|19|They rose early in the morning and worshiped before the LORD; then they went back to their house at Ramah. And Elkanah knew Hannah his wife, and the LORD remembered her.
1SAM|1|20|And in due time Hannah conceived and bore a son, and she called his name Samuel, for she said, "I have asked for him from the LORD."
1SAM|1|21|The man Elkanah and all his house went up to offer to the LORD the yearly sacrifice and to pay his vow.
1SAM|1|22|But Hannah did not go up, for she said to her husband, "As soon as the child is weaned, I will bring him, so that he may appear in the presence of the LORD and dwell there forever."
1SAM|1|23|Elkanah her husband said to her, "Do what seems best to you; wait until you have weaned him; only, may the LORD establish his word." So the woman remained and nursed her son until she weaned him.
1SAM|1|24|And when she had weaned him, she took him up with her, along with a three-year-old bull, an ephah of flour, and a skin of wine, and she brought him to the house of the LORD at Shiloh. And the child was young.
1SAM|1|25|Then they slaughtered the bull, and they brought the child to Eli.
1SAM|1|26|And she said, "Oh, my lord! As you live, my lord, I am the woman who was standing here in your presence, praying to the LORD.
1SAM|1|27|For this child I prayed, and the LORD has granted me my petition that I made to him.
1SAM|1|28|Therefore I have lent him to the LORD. As long as he lives, he is lent to the LORD." And he worshiped the LORD there.
1SAM|2|1|And Hannah prayed and said, "My heart exults in the LORD; my strength is exalted in the LORD. My mouth derides my enemies, because I rejoice in your salvation.
1SAM|2|2|"There is none holy like the LORD; there is none besides you; there is no rock like our God.
1SAM|2|3|Talk no more so very proudly, let not arrogance come from your mouth; for the LORD is a God of knowledge, and by him actions are weighed.
1SAM|2|4|The bows of the mighty are broken, but the feeble bind on strength.
1SAM|2|5|Those who were full have hired themselves out for bread, but those who were hungry have ceased to hunger. The barren has borne seven, but she who has many children is forlorn.
1SAM|2|6|The LORD kills and brings to life; he brings down to Sheol and raises up.
1SAM|2|7|The LORD makes poor and makes rich; he brings low and he exalts.
1SAM|2|8|He raises up the poor from the dust; he lifts the needy from the ash heap to make them sit with princes and inherit a seat of honor. For the pillars of the earth are the LORD's, and on them he has set the world.
1SAM|2|9|"He will guard the feet of his faithful ones, but the wicked shall be cut off in darkness, for not by might shall a man prevail.
1SAM|2|10|The adversaries of the LORD shall be broken to pieces; against them he will thunder in heaven. The LORD will judge the ends of the earth; he will give strength to his king and exalt the power of his anointed."
1SAM|2|11|Then Elkanah went home to Ramah. And the boy ministered to the LORD in the presence of Eli the priest.
1SAM|2|12|Now the sons of Eli were worthless men. They did not know the LORD.
1SAM|2|13|The custom of the priests with the people was that when any man offered sacrifice, the priest's servant would come, while the meat was boiling, with a three-pronged fork in his hand,
1SAM|2|14|and he would thrust it into the pan or kettle or cauldron or pot. All that the fork brought up the priest would take for himself. This is what they did at Shiloh to all the Israelites who came there.
1SAM|2|15|Moreover, before the fat was burned, the priest's servant would come and say to the man who was sacrificing, "Give meat for the priest to roast, for he will not accept boiled meat from you but only raw."
1SAM|2|16|And if the man said to him, "Let them burn the fat first, and then take as much as you wish," he would say, "No, you must give it now, and if not, I will take it by force."
1SAM|2|17|Thus the sin of the young men was very great in the sight of the LORD, for the men treated the offering of the LORD with contempt.
1SAM|2|18|Samuel was ministering before the LORD, a boy clothed with a linen ephod.
1SAM|2|19|And his mother used to make for him a little robe and take it to him each year when she went up with her husband to offer the yearly sacrifice.
1SAM|2|20|Then Eli would bless Elkanah and his wife, and say, "May the LORD give you children by this woman for the petition she asked of the LORD." So then they would return to their home.
1SAM|2|21|Indeed the LORD visited Hannah, and she conceived and bore three sons and two daughters. And the young man Samuel grew in the presence of the LORD.
1SAM|2|22|Now Eli was very old, and he kept hearing all that his sons were doing to all Israel, and how they lay with the women who were serving at the entrance to the tent of meeting.
1SAM|2|23|And he said to them, "Why do you do such things? For I hear of your evil dealings from all the people.
1SAM|2|24|No, my sons; it is no good report that I hear the people of the LORD spreading abroad.
1SAM|2|25|If someone sins against a man, God will mediate for him, but if someone sins against the LORD, who can intercede for him?" But they would not listen to the voice of their father, for it was the will of the LORD to put them to death.
1SAM|2|26|Now the young man Samuel continued to grow both in stature and in favor with the LORD and also with man.
1SAM|2|27|And there came a man of God to Eli and said to him, "Thus the LORD has said, 'Did I indeed reveal myself to the house of your father when they were in Egypt subject to the house of Pharaoh?
1SAM|2|28|Did I choose him out of all the tribes of Israel to be my priest, to go up to my altar, to burn incense, to wear an ephod before me? I gave to the house of your father all my offerings by fire from the people of Israel.
1SAM|2|29|Why then do you scorn my sacrifices and my offerings that I commanded, and honor your sons above me by fattening yourselves on the choicest parts of every offering of my people Israel?'
1SAM|2|30|Therefore the LORD the God of Israel declares: 'I promised that your house and the house of your father should go in and out before me forever,' but now the LORD declares: 'Far be it from me, for those who honor me I will honor, and those who despise me shall be lightly esteemed.
1SAM|2|31|Behold, the days are coming when I will cut off your strength and the strength of your father's house, so that there will not be an old man in your house.
1SAM|2|32|Then in distress you will look with envious eye on all the prosperity that shall be bestowed on Israel, and there shall not be an old man in your house forever.
1SAM|2|33|The only one of you whom I shall not cut off from my altar shall be spared to weep his eyes out to grieve his heart, and all the descendants of your house shall die by the sword of men.
1SAM|2|34|And this that shall come upon your two sons, Hophni and Phinehas, shall be the sign to you: both of them shall die on the same day.
1SAM|2|35|And I will raise up for myself a faithful priest, who shall do according to what is in my heart and in my mind. And I will build him a sure house, and he shall go in and out before my anointed forever.
1SAM|2|36|And everyone who is left in your house shall come to implore him for a piece of silver or a loaf of bread and shall say, "Please put me in one of the priests' places, that I may eat a morsel of bread."'"
1SAM|3|1|Now the young man Samuel was ministering to the LORD under Eli. And the word of the LORD was rare in those days; there was no frequent vision.
1SAM|3|2|At that time Eli, whose eyesight had begun to grow dim so that he could not see, was lying down in his own place.
1SAM|3|3|The lamp of God had not yet gone out, and Samuel was lying down in the temple of the LORD, where the ark of God was.
1SAM|3|4|Then the LORD called Samuel, and he said, "Here I am!"
1SAM|3|5|and ran to Eli and said, "Here I am, for you called me." But he said, "I did not call; lie down again." So he went and lay down.
1SAM|3|6|And the LORD called again, "Samuel!" and Samuel arose and went to Eli and said, "Here I am, for you called me." But he said, "I did not call, my son; lie down again."
1SAM|3|7|Now Samuel did not yet know the LORD, and the word of the LORD had not yet been revealed to him.
1SAM|3|8|And the LORD called Samuel again the third time. And he arose and went to Eli and said, "Here I am, for you called me." Then Eli perceived that the LORD was calling the young man.
1SAM|3|9|Therefore Eli said to Samuel, "Go, lie down, and if he calls you, you shall say, 'Speak, LORD, for your servant hears.'"So Samuel went and lay down in his place.
1SAM|3|10|And the LORD came and stood, calling as at other times, "Samuel! Samuel!" And Samuel said, "Speak, for your servant hears."
1SAM|3|11|Then the LORD said to Samuel, "Behold, I am about to do a thing in Israel at which the two ears of everyone who hears it will tingle.
1SAM|3|12|On that day I will fulfill against Eli all that I have spoken concerning his house, from beginning to end.
1SAM|3|13|And I declare to him that I am about to punish his house forever, for the iniquity that he knew, because his sons were blaspheming God, and he did not restrain them.
1SAM|3|14|Therefore I swear to the house of Eli that the iniquity of Eli's house shall not be atoned for by sacrifice or offering forever."
1SAM|3|15|Samuel lay until morning; then he opened the doors of the house of the LORD. And Samuel was afraid to tell the vision to Eli.
1SAM|3|16|But Eli called Samuel and said, "Samuel, my son." And he said, "Here I am."
1SAM|3|17|And Eli said, "What was it that he told you? Do not hide it from me. May God do so to you and more also if you hide anything from me of all that he told you."
1SAM|3|18|So Samuel told him everything and hid nothing from him. And he said, "It is the LORD. Let him do what seems good to him."
1SAM|3|19|And Samuel grew, and the LORD was with him and let none of his words fall to the ground.
1SAM|3|20|And all Israel from Dan to Beersheba knew that Samuel was established as a prophet of the LORD.
1SAM|3|21|And the LORD appeared again at Shiloh, for the LORD revealed himself to Samuel at Shiloh by the word of the LORD.
1SAM|4|1|And the word of Samuel came to all Israel. Now Israel went out to battle against the Philistines. They encamped at Ebenezer, and the Philistines encamped at Aphek.
1SAM|4|2|The Philistines drew up in line against Israel, and when the battle spread, Israel was defeated by the Philistines, who killed about four thousand men on the field of battle.
1SAM|4|3|And when the troops came to the camp, the elders of Israel said, "Why has the LORD defeated us today before the Philistines? Let us bring the ark of the covenant of the LORD here from Shiloh, that it may come among us and save us from the power of our enemies."
1SAM|4|4|So the people sent to Shiloh and brought from there the ark of the covenant of the LORD of hosts, who is enthroned on the cherubim. And the two sons of Eli, Hophni and Phinehas, were there with the ark of the covenant of God.
1SAM|4|5|As soon as the ark of the covenant of the LORD came into the camp, all Israel gave a mighty shout, so that the earth resounded.
1SAM|4|6|And when the Philistines heard the noise of the shouting, they said, "What does this great shouting in the camp of the Hebrews mean?" And when they learned that the ark of the LORD had come to the camp,
1SAM|4|7|the Philistines were afraid, for they said, "A god has come into the camp." And they said, "Woe to us! For nothing like this has happened before.
1SAM|4|8|Woe to us! Who can deliver us from the power of these mighty gods? These are the gods who struck the Egyptians with every sort of plague in the wilderness.
1SAM|4|9|Take courage, and be men, O Philistines, lest you become slaves to the Hebrews as they have been to you; be men and fight."
1SAM|4|10|So the Philistines fought, and Israel was defeated, and they fled, every man to his home. And there was a very great slaughter, for there fell of Israel thirty thousand foot soldiers.
1SAM|4|11|And the ark of God was captured, and the two sons of Eli, Hophni and Phinehas, died.
1SAM|4|12|A man of Benjamin ran from the battle line and came to Shiloh the same day, with his clothes torn and with dirt on his head.
1SAM|4|13|When he arrived, Eli was sitting on his seat by the road watching, for his heart trembled for the ark of God. And when the man came into the city and told the news, all the city cried out.
1SAM|4|14|When Eli heard the sound of the outcry, he said, "What is this uproar?" Then the man hurried and came and told Eli.
1SAM|4|15|Now Eli was ninety-eight years old and his eyes were set so that he could not see.
1SAM|4|16|And the man said to Eli, "I am he who has come from the battle; I fled from the battle today." And he said, "How did it go, my son?"
1SAM|4|17|He who brought the news answered and said, "Israel has fled before the Philistines, and there has also been a great defeat among the people. Your two sons also, Hophni and Phinehas, are dead, and the ark of God has been captured."
1SAM|4|18|As soon as he mentioned the ark of God, Eli fell over backward from his seat by the side of the gate, and his neck was broken and he died, for the man was old and heavy. He had judged Israel forty years.
1SAM|4|19|Now his daughter-in-law, the wife of Phinehas, was pregnant, about to give birth. And when she heard the news that the ark of God was captured, and that her father-in-law and her husband were dead, she bowed and gave birth, for her pains came upon her.
1SAM|4|20|And about the time of her death the women attending her said to her, "Do not be afraid, for you have borne a son." But she did not answer or pay attention.
1SAM|4|21|And she named the child Ichabod, saying, "The glory has departed from Israel!" because the ark of God had been captured and because of her father-in-law and her husband.
1SAM|4|22|And she said, "The glory has departed from Israel, for the ark of God has been captured."
1SAM|5|1|When the Philistines captured the ark of God, they brought it from Ebenezer to Ashdod.
1SAM|5|2|Then the Philistines took the ark of God and brought it into the house of Dagon and set it up beside Dagon.
1SAM|5|3|And when the people of Ashdod rose early the next day, behold, Dagon had fallen face downward on the ground before the ark of the LORD. So they took Dagon and put him back in his place.
1SAM|5|4|But when they rose early on the next morning, behold, Dagon had fallen face downward on the ground before the ark of the LORD, and the head of Dagon and both his hands were lying cut off on the threshold. Only the trunk of Dagon was left to him.
1SAM|5|5|This is why the priests of Dagon and all who enter the house of Dagon do not tread on the threshold of Dagon in Ashdod to this day.
1SAM|5|6|The hand of the LORD was heavy against the people of Ashdod, and he terrified and afflicted them with tumors, both Ashdod and its territory.
1SAM|5|7|And when the men of Ashdod saw how things were, they said, "The ark of the God of Israel must not remain with us, for his hand is hard against us and against Dagon our god."
1SAM|5|8|So they sent and gathered together all the lords of the Philistines and said, "What shall we do with the ark of the God of Israel?" They answered, "Let the ark of the God of Israel be brought around to Gath." So they brought the ark of the God of Israel there.
1SAM|5|9|But after they had brought it around, the hand of the LORD was against the city, causing a very great panic, and he afflicted the men of the city, both young and old, so that tumors broke out on them.
1SAM|5|10|So they sent the ark of God to Ekron. But as soon as the ark of God came to Ekron, the people of Ekron cried out, "They have brought around to us the ark of the God of Israel to kill us and our people."
1SAM|5|11|They sent therefore and gathered together all the lords of the Philistines and said, "Send away the ark of the God of Israel, and let it return to its own place, that it may not kill us and our people." For there was a deathly panic throughout the whole city. The hand of God was very heavy there.
1SAM|5|12|The men who did not die were struck with tumors, and the cry of the city went up to heaven.
1SAM|6|1|The ark of the LORD was in the country of the Philistines seven months.
1SAM|6|2|And the Philistines called for the priests and the diviners and said, "What shall we do with the ark of the LORD? Tell us with what we shall send it to its place."
1SAM|6|3|They said, "If you send away the ark of the God of Israel, do not send it empty, but by all means return him a guilt offering. Then you will be healed, and it will be known to you why his hand does not turn away from you."
1SAM|6|4|And they said, "What is the guilt offering that we shall return to him?" They answered, "Five golden tumors and five golden mice, according to the number of the lords of the Philistines, for the same plague was on all of you and on your lords.
1SAM|6|5|So you must make images of your tumors and images of your mice that ravage the land, and give glory to the God of Israel. Perhaps he will lighten his hand from off you and your gods and your land.
1SAM|6|6|Why should you harden your hearts as the Egyptians and Pharaoh hardened their hearts? After he had dealt severely with them, did they not send the people away, and they departed?
1SAM|6|7|Now then, take and prepare a new cart and two milk cows on which there has never come a yoke, and yoke the cows to the cart, but take their calves home, away from them.
1SAM|6|8|And take the ark of the LORD and place it on the cart and put in a box at its side the figures of gold, which you are returning to him as a guilt offering. Then send it off and let it go its way
1SAM|6|9|and watch. If it goes up on the way to its own land, to Beth-shemesh, then it is he who has done us this great harm, but if not, then we shall know that it is not his hand that struck us; it happened to us by coincidence."
1SAM|6|10|The men did so, and took two milk cows and yoked them to the cart and shut up their calves at home.
1SAM|6|11|And they put the ark of the LORD on the cart and the box with the golden mice and the images of their tumors.
1SAM|6|12|And the cows went straight in the direction of Beth-shemesh along one highway, lowing as they went. They turned neither to the right nor to the left, and the lords of the Philistines went after them as far as the border of Beth-shemesh.
1SAM|6|13|Now the people of Beth-shemesh were reaping their wheat harvest in the valley. And when they lifted up their eyes and saw the ark, they rejoiced to see it.
1SAM|6|14|The cart came into the field of Joshua of Beth-shemesh and stopped there. A great stone was there. And they split up the wood of the cart and offered the cows as a burnt offering to the LORD.
1SAM|6|15|And the Levites took down the ark of the LORD and the box that was beside it, in which were the golden figures, and set them upon the great stone. And the men of Beth-shemesh offered burnt offerings and sacrificed sacrifices on that day to the LORD.
1SAM|6|16|And when the five lords of the Philistines saw it, they returned that day to Ekron.
1SAM|6|17|These are the golden tumors that the Philistines returned as a guilt offering to the LORD: one for Ashdod, one for Gaza, one for Ashkelon, one for Gath, one for Ekron,
1SAM|6|18|and the golden mice, according to the number of all the cities of the Philistines belonging to the five lords, both fortified cities and unwalled villages. The great stone beside which they set down the ark of the LORD is a witness to this day in the field of Joshua of Beth-shemesh.
1SAM|6|19|And he struck some of the men of Beth-shemesh, because they looked upon the ark of the LORD. He struck seventy men of them, and the people mourned because the LORD had struck the people with a great blow.
1SAM|6|20|Then the men of Beth-shemesh said, "Who is able to stand before the LORD, this holy God? And to whom shall he go up away from us?"
1SAM|6|21|So they sent messengers to the inhabitants of Kiriath-jearim, saying, "The Philistines have returned the ark of the LORD. Come down and take it up to you."
1SAM|7|1|And the men of Kiriath-jearim came and took up the ark of the LORD and brought it to the house of Abinadab on the hill. And they consecrated his son Eleazar to have charge of the ark of the LORD.
1SAM|7|2|From the day that the ark was lodged at Kiriath-jearim, a long time passed, some twenty years, and all the house of Israel lamented after the LORD.
1SAM|7|3|And Samuel said to all the house of Israel, "If you are returning to the LORD with all your heart, then put away the foreign gods and the Ashtaroth from among you and direct your heart to the LORD and serve him only, and he will deliver you out of the hand of the Philistines."
1SAM|7|4|So the people of Israel put away the Baals and the Ashtaroth, and they served the LORD only.
1SAM|7|5|Then Samuel said, "Gather all Israel at Mizpah, and I will pray to the LORD for you."
1SAM|7|6|So they gathered at Mizpah and drew water and poured it out before the LORD and fasted on that day and said there, "We have sinned against the LORD." And Samuel judged the people of Israel at Mizpah.
1SAM|7|7|Now when the Philistines heard that the people of Israel had gathered at Mizpah, the lords of the Philistines went up against Israel. And when the people of Israel heard of it, they were afraid of the Philistines.
1SAM|7|8|And the people of Israel said to Samuel, "Do not cease to cry out to the LORD our God for us, that he may save us from the hand of the Philistines."
1SAM|7|9|So Samuel took a nursing lamb and offered it as a whole burnt offering to the LORD. And Samuel cried out to the LORD for Israel, and the LORD answered him.
1SAM|7|10|As Samuel was offering up the burnt offering, the Philistines drew near to attack Israel. But the LORD thundered with a mighty sound that day against the Philistines and threw them into confusion, and they were routed before Israel.
1SAM|7|11|And the men of Israel went out from Mizpah and pursued the Philistines and struck them, as far as below Beth-car.
1SAM|7|12|Then Samuel took a stone and set it up between Mizpah and Shen and called its name Ebenezer; for he said, "Till now the LORD has helped us."
1SAM|7|13|So the Philistines were subdued and did not again enter the territory of Israel. And the hand of the LORD was against the Philistines all the days of Samuel.
1SAM|7|14|The cities that the Philistines had taken from Israel were restored to Israel, from Ekron to Gath, and Israel delivered their territory from the hand of the Philistines. There was peace also between Israel and the Amorites.
1SAM|7|15|Samuel judged Israel all the days of his life.
1SAM|7|16|And he went on a circuit year by year to Bethel, Gilgal, and Mizpah. And he judged Israel in all these places.
1SAM|7|17|Then he would return to Ramah, for his home was there, and there also he judged Israel. And he built there an altar to the LORD.
1SAM|8|1|When Samuel became old, he made his sons judges over Israel.
1SAM|8|2|The name of his firstborn son was Joel, and the name of his second, Abijah; they were judges in Beersheba.
1SAM|8|3|Yet his sons did not walk in his ways but turned aside after gain. They took bribes and perverted justice.
1SAM|8|4|Then all the elders of Israel gathered together and came to Samuel at Ramah
1SAM|8|5|and said to him, "Behold, you are old and your sons do not walk in your ways. Now appoint for us a king to judge us like all the nations."
1SAM|8|6|But the thing displeased Samuel when they said, "Give us a king to judge us." And Samuel prayed to the LORD.
1SAM|8|7|And the LORD said to Samuel, "Obey the voice of the people in all that they say to you, for they have not rejected you, but they have rejected me from being king over them.
1SAM|8|8|According to all the deeds that they have done, from the day I brought them up out of Egypt even to this day, forsaking me and serving other gods, so they are also doing to you.
1SAM|8|9|Now then, obey their voice; only you shall solemnly warn them and show them the ways of the king who shall reign over them."
1SAM|8|10|So Samuel told all the words of the LORD to the people who were asking for a king from him.
1SAM|8|11|He said, "These will be the ways of the king who will reign over you: he will take your sons and appoint them to his chariots and to be his horsemen and to run before his chariots.
1SAM|8|12|And he will appoint for himself commanders of thousands and commanders of fifties, and some to plow his ground and to reap his harvest, and to make his implements of war and the equipment of his chariots.
1SAM|8|13|He will take your daughters to be perfumers and cooks and bakers.
1SAM|8|14|He will take the best of your fields and vineyards and olive orchards and give them to his servants.
1SAM|8|15|He will take the tenth of your grain and of your vineyards and give it to his officers and to his servants.
1SAM|8|16|He will take your male servants and female servants and the best of your young men and your donkeys, and put them to his work.
1SAM|8|17|He will take the tenth of your flocks, and you shall be his slaves.
1SAM|8|18|And in that day you will cry out because of your king, whom you have chosen for yourselves, but the LORD will not answer you in that day."
1SAM|8|19|But the people refused to obey the voice of Samuel. And they said, "No! But there shall be a king over us,
1SAM|8|20|that we also may be like all the nations, and that our king may judge us and go out before us and fight our battles."
1SAM|8|21|And when Samuel had heard all the words of the people, he repeated them in the ears of the LORD.
1SAM|8|22|And the LORD said to Samuel, "Obey their voice and make them a king." Samuel then said to the men of Israel, "Go every man to his city."
1SAM|9|1|There was a man of Benjamin whose name was Kish, the son of Abiel, son of Zeror, son of Becorath, son of Aphiah, a Benjaminite, a man of wealth.
1SAM|9|2|And he had a son whose name was Saul, a handsome young man. There was not a man among the people of Israel more handsome than he. From his shoulders upward he was taller than any of the people.
1SAM|9|3|Now the donkeys of Kish, Saul's father, were lost. So Kish said to Saul his son, "Take one of the young men with you, and arise, go and look for the donkeys."
1SAM|9|4|And he passed through the hill country of Ephraim and passed through the land of Shalishah, but they did not find them. And they passed through the land of Shaalim, but they were not there. Then they passed through the land of Benjamin, but did not find them.
1SAM|9|5|When they came to the land of Zuph, Saul said to his servant who was with him, "Come, let us go back, lest my father cease to care about the donkeys and become anxious about us."
1SAM|9|6|But he said to him, "Behold, there is a man of God in this city, and he is a man who is held in honor; all that he says comes true. So now let us go there. Perhaps he can tell us the way we should go."
1SAM|9|7|Then Saul said to his servant, "But if we go, what can we bring the man? For the bread in our sacks is gone, and there is no present to bring to the man of God. What do we have?"
1SAM|9|8|The servant answered Saul again, "Here, I have with me a quarter of a shekel of silver, and I will give it to the man of God to tell us our way."
1SAM|9|9|(Formerly in Israel, when a man went to inquire of God, he said, "Come, let us go to the seer," for today's "prophet" was formerly called a seer.)
1SAM|9|10|And Saul said to his servant, "Well said; come, let us go." So they went to the city where the man of God was.
1SAM|9|11|As they went up the hill to the city, they met young women coming out to draw water and said to them, "Is the seer here?"
1SAM|9|12|They answered, "He is; behold, he is just ahead of you. Hurry. He has come just now to the city, because the people have a sacrifice today on the high place.
1SAM|9|13|As soon as you enter the city you will find him, before he goes up to the high place to eat. For the people will not eat till he comes, since he must bless the sacrifice; afterward those who are invited will eat. Now go up, for you will meet him immediately."
1SAM|9|14|So they went up to the city. As they were entering the city, they saw Samuel coming out toward them on his way up to the high place.
1SAM|9|15|Now the day before Saul came, the LORD had revealed to Samuel:
1SAM|9|16|"Tomorrow about this time I will send to you a man from the land of Benjamin, and you shall anoint him to be prince over my people Israel. He shall save my people from the hand of the Philistines. For I have seen my people, because their cry has come to me."
1SAM|9|17|When Samuel saw Saul, the LORD told him, "Here is the man of whom I spoke to you! He it is who shall restrain my people."
1SAM|9|18|Then Saul approached Samuel in the gate and said, "Tell me where is the house of the seer?"
1SAM|9|19|Samuel answered Saul, "I am the seer. Go up before me to the high place, for today you shall eat with me, and in the morning I will let you go and will tell you all that is on your mind.
1SAM|9|20|As for your donkeys that were lost three days ago, do not set your mind on them, for they have been found. And for whom is all that is desirable in Israel? Is it not for you and for all your father's house?"
1SAM|9|21|Saul answered, "Am I not a Benjaminite, from the least of the tribes of Israel? And is not my clan the humblest of all the clans of the tribe of Benjamin? Why then have you spoken to me in this way?"
1SAM|9|22|Then Samuel took Saul and his young man and brought them into the hall and gave them a place at the head of those who had been invited, who were about thirty persons.
1SAM|9|23|And Samuel said to the cook, "Bring the portion I gave you, of which I said to you, 'Put it aside.'"
1SAM|9|24|So the cook took up the leg and what was on it and set them before Saul. And Samuel said, "See, what was kept is set before you. Eat, because it was kept for you until the hour appointed, that you might eat with the guests." So Saul ate with Samuel that day.
1SAM|9|25|And when they came down from the high place into the city, a bed was spread for Saul on the roof, and he lay down to sleep.
1SAM|9|26|Then at the break of dawn Samuel called to Saul on the roof, "Up, that I may send you on your way." So Saul arose, and both he and Samuel went out into the street.
1SAM|9|27|As they were going down to the outskirts of the city, Samuel said to Saul, "Tell the servant to pass on before us, and when he has passed on, stop here yourself for a while, that I may make known to you the word of God."
1SAM|10|1|Then Samuel took a flask of oil and poured it on his head and kissed him and said, "Has not the LORD anointed you to be prince over his people Israel? And you shall reign over the people of the LORD and you will save them from the hand of their surrounding enemies. And this shall be the sign to you that the LORD has anointed you to be prince over his heritage.
1SAM|10|2|When you depart from me today, you will meet two men by Rachel's tomb in the territory of Benjamin at Zelzah, and they will say to you, 'The donkeys that you went to seek are found, and now your father has ceased to care about the donkeys and is anxious about you, saying, "What shall I do about my son?"'
1SAM|10|3|Then you shall go on from there further and come to the oak of Tabor. Three men going up to God at Bethel will meet you there, one carrying three young goats, another carrying three loaves of bread, and another carrying a skin of wine.
1SAM|10|4|And they will greet you and give you two loaves of bread, which you shall accept from their hand.
1SAM|10|5|After that you shall come to Gibeath-elohim, where there is a garrison of the Philistines. And there, as soon as you come to the city, you will meet a group of prophets coming down from the high place with harp, tambourine, flute, and lyre before them, prophesying.
1SAM|10|6|Then the Spirit of the LORD will rush upon you, and you will prophesy with them and be turned into another man.
1SAM|10|7|Now when these signs meet you, do what your hand finds to do, for God is with you.
1SAM|10|8|Then go down before me to Gilgal. And behold, I am coming to you to offer burnt offerings and to sacrifice peace offerings. Seven days you shall wait, until I come to you and show you what you shall do."
1SAM|10|9|When he turned his back to leave Samuel, God gave him another heart. And all these signs came to pass that day.
1SAM|10|10|When they came to Gibeah, behold, a group of prophets met him, and the Spirit of God rushed upon him, and he prophesied among them.
1SAM|10|11|And when all who knew him previously saw how he prophesied with the prophets, the people said to one another, "What has come over the son of Kish? Is Saul also among the prophets?"
1SAM|10|12|And a man of the place answered, "And who is their father?" Therefore it became a proverb, "Is Saul also among the prophets?"
1SAM|10|13|When he had finished prophesying, he came to the high place.
1SAM|10|14|Saul's uncle said to him and to his servant, "Where did you go?" And he said, "To seek the donkeys. And when we saw they were not to be found, we went to Samuel."
1SAM|10|15|And Saul's uncle said, "Please tell me what Samuel said to you."
1SAM|10|16|And Saul said to his uncle, "He told us plainly that the donkeys had been found." But about the matter of the kingdom, of which Samuel had spoken, he did not tell him anything.
1SAM|10|17|Now Samuel called the people together to the LORD at Mizpah.
1SAM|10|18|And he said to the people of Israel, "Thus says the LORD, the God of Israel, 'I brought up Israel out of Egypt, and I delivered you from the hand of the Egyptians and from the hand of all the kingdoms that were oppressing you.'
1SAM|10|19|But today you have rejected your God, who saves you from all your calamities and your distresses, and you have said to him, 'Set a king over us.' Now therefore present yourselves before the LORD by your tribes and by your thousands."
1SAM|10|20|Then Samuel brought all the tribes of Israel near, and the tribe of Benjamin was taken by lot.
1SAM|10|21|He brought the tribe of Benjamin near by its clans, and the clan of the Matrites was taken by lot; and Saul the son of Kish was taken by lot. But when they sought him, he could not be found.
1SAM|10|22|So they inquired again of the LORD, "Is there a man still to come?" and the LORD said, "Behold, he has hidden himself among the baggage."
1SAM|10|23|Then they ran and took him from there. And when he stood among the people, he was taller than any of the people from his shoulders upward.
1SAM|10|24|And Samuel said to all the people, "Do you see him whom the LORD has chosen? There is none like him among all the people." And all the people shouted, "Long live the king!"
1SAM|10|25|Then Samuel told the people the rights and duties of the kingship, and he wrote them in a book and laid it up before the LORD. Then Samuel sent all the people away, each one to his home.
1SAM|10|26|Saul also went to his home at Gibeah, and with him went men of valor whose hearts God had touched.
1SAM|10|27|But some worthless fellows said, "How can this man save us?" And they despised him and brought him no present. But he held his peace.
1SAM|11|1|Then Nahash the Ammonite went up and besieged Jabesh-gilead, and all the men of Jabesh said to Nahash, "Make a treaty with us, and we will serve you."
1SAM|11|2|But Nahash the Ammonite said to them, "On this condition I will make a treaty with you, that I gouge out all your right eyes, and thus bring disgrace on all Israel."
1SAM|11|3|The elders of Jabesh said to him, "Give us seven days respite that we may send messengers through all the territory of Israel. Then, if there is no one to save us, we will give ourselves up to you."
1SAM|11|4|When the messengers came to Gibeah of Saul, they reported the matter in the ears of the people, and all the people wept aloud.
1SAM|11|5|Now, behold, Saul was coming from the field behind the oxen. And Saul said, "What is wrong with the people, that they are weeping?" So they told him the news of the men of Jabesh.
1SAM|11|6|And the Spirit of God rushed upon Saul when he heard these words, and his anger was greatly kindled.
1SAM|11|7|He took a yoke of oxen and cut them in pieces and sent them throughout all the territory of Israel by the hand of messengers, saying, "Whoever does not come out after Saul and Samuel, so shall it be done to his oxen!" Then the dread of the LORD fell upon the people, and they came out as one man.
1SAM|11|8|When he mustered them at Bezek, the people of Israel were three hundred thousand, and the men of Judah thirty thousand.
1SAM|11|9|And they said to the messengers who had come, "Thus shall you say to the men of Jabesh-gilead: 'Tomorrow, by the time the sun is hot, you shall have deliverance.'"When the messengers came and told the men of Jabesh, they were glad.
1SAM|11|10|Therefore the men of Jabesh said, "Tomorrow we will give ourselves up to you, and you may do to us whatever seems good to you."
1SAM|11|11|And the next day Saul put the people in three companies. And they came into the midst of the camp in the morning watch and struck down the Ammonites until the heat of the day. And those who survived were scattered, so that no two of them were left together.
1SAM|11|12|Then the people said to Samuel, "Who is it that said, 'Shall Saul reign over us?' Bring the men, that we may put them to death."
1SAM|11|13|But Saul said, "Not a man shall be put to death this day, for today the LORD has worked salvation in Israel."
1SAM|11|14|Then Samuel said to the people, "Come, let us go to Gilgal and there renew the kingdom."
1SAM|11|15|So all the people went to Gilgal, and there they made Saul king before the LORD in Gilgal. There they sacrificed peace offerings before the LORD, and there Saul and all the men of Israel rejoiced greatly.
1SAM|12|1|And Samuel said to all Israel, "Behold, I have obeyed your voice in all that you have said to me and have made a king over you.
1SAM|12|2|And now, behold, the king walks before you, and I am old and gray; and behold, my sons are with you. I have walked before you from my youth until this day.
1SAM|12|3|Here I am; testify against me before the LORD and before his anointed. Whose ox have I taken? Or whose donkey have I taken? Or whom have I defrauded? Whom have I oppressed? Or from whose hand have I taken a bribe to blind my eyes with it? Testify against me and I will restore it to you."
1SAM|12|4|They said, "You have not defrauded us or oppressed us or taken anything from any man's hand."
1SAM|12|5|And he said to them, "The LORD is witness against you, and his anointed is witness this day, that you have not found anything in my hand." And they said, "He is witness."
1SAM|12|6|And Samuel said to the people, "The LORD is witness, who appointed Moses and Aaron and brought your fathers up out of the land of Egypt.
1SAM|12|7|Now therefore stand still that I may plead with you before the LORD concerning all the righteous deeds of the LORD that he performed for you and for your fathers.
1SAM|12|8|When Jacob went into Egypt, and the Egyptians oppressed them, then your fathers cried out to the LORD and the LORD sent Moses and Aaron, who brought your fathers out of Egypt and made them dwell in this place.
1SAM|12|9|But they forgot the LORD their God. And he sold them into the hand of Sisera, commander of the army of Hazor, and into the hand of the Philistines, and into the hand of the king of Moab. And they fought against them.
1SAM|12|10|And they cried out to the LORD and said, 'We have sinned, because we have forsaken the LORD and have served the Baals and the Ashtaroth. But now deliver us out of the hand of our enemies, that we may serve you.'
1SAM|12|11|And the LORD sent Jerubbaal and Barak and Jephthah and Samuel and delivered you out of the hand of your enemies on every side, and you lived in safety.
1SAM|12|12|And when you saw that Nahash the king of the Ammonites came against you, you said to me, 'No, but a king shall reign over us,' when the LORD your God was your king.
1SAM|12|13|And now behold the king whom you have chosen, for whom you have asked; behold, the LORD has set a king over you.
1SAM|12|14|If you will fear the LORD and serve him and obey his voice and not rebel against the commandment of the LORD, and if both you and the king who reigns over you will follow the LORD your God, it will be well.
1SAM|12|15|But if you will not obey the voice of the LORD, but rebel against the commandment of the LORD, then the hand of the LORD will be against you and your king.
1SAM|12|16|Now therefore stand still and see this great thing that the LORD will do before your eyes.
1SAM|12|17|Is it not wheat harvest today? I will call upon the LORD, that he may send thunder and rain. And you shall know and see that your wickedness is great, which you have done in the sight of the LORD, in asking for yourselves a king."
1SAM|12|18|So Samuel called upon the LORD, and the LORD sent thunder and rain that day, and all the people greatly feared the LORD and Samuel.
1SAM|12|19|And all the people said to Samuel, "Pray for your servants to the LORD your God, that we may not die, for we have added to all our sins this evil, to ask for ourselves a king."
1SAM|12|20|And Samuel said to the people, "Do not be afraid; you have done all this evil. Yet do not turn aside from following the LORD, but serve the LORD with all your heart.
1SAM|12|21|And do not turn aside after empty things that cannot profit or deliver, for they are empty.
1SAM|12|22|For the LORD will not forsake his people, for his great name's sake, because it has pleased the LORD to make you a people for himself.
1SAM|12|23|Moreover, as for me, far be it from me that I should sin against the LORD by ceasing to pray for you, and I will instruct you in the good and the right way.
1SAM|12|24|Only fear the LORD and serve him faithfully with all your heart. For consider what great things he has done for you.
1SAM|12|25|But if you still do wickedly, you shall be swept away, both you and your king."
1SAM|13|1|Saul was... years old when he began to reign, and he reigned... and two years over Israel.
1SAM|13|2|Saul chose three thousand men of Israel. Two thousand were with Saul in Michmash and the hill country of Bethel, and a thousand were with Jonathan in Gibeah of Benjamin. The rest of the people he sent home, every man to his tent.
1SAM|13|3|Jonathan defeated the garrison of the Philistines that was at Geba, and the Philistines heard of it. And Saul blew the trumpet throughout all the land, saying, "Let the Hebrews hear."
1SAM|13|4|And all Israel heard it said that Saul had defeated the garrison of the Philistines, and also that Israel had become a stench to the Philistines. And the people were called out to join Saul at Gilgal.
1SAM|13|5|And the Philistines mustered to fight with Israel, thirty thousand chariots and six thousand horsemen and troops like the sand on the seashore in multitude. They came up and encamped in Michmash, to the east of Beth-aven.
1SAM|13|6|When the men of Israel saw that they were in trouble (for the people were hard pressed), the people hid themselves in caves and in holes and in rocks and in tombs and in cisterns,
1SAM|13|7|and some Hebrews crossed the fords of the Jordan to the land of Gad and Gilead. Saul was still at Gilgal, and all the people followed him trembling.
1SAM|13|8|He waited seven days, the time appointed by Samuel. But Samuel did not come to Gilgal, and the people were scattering from him.
1SAM|13|9|So Saul said, "Bring the burnt offering here to me, and the peace offerings." And he offered the burnt offering.
1SAM|13|10|As soon as he had finished offering the burnt offering, behold, Samuel came. And Saul went out to meet him and greet him.
1SAM|13|11|Samuel said, "What have you done?" And Saul said, "When I saw that the people were scattering from me, and that you did not come within the days appointed, and that the Philistines had mustered at Michmash,
1SAM|13|12|I said, 'Now the Philistines will come down against me at Gilgal, and I have not sought the favor of the LORD.' So I forced myself, and offered the burnt offering."
1SAM|13|13|And Samuel said to Saul, "You have done foolishly. You have not kept the command of the LORD your God, with which he commanded you. For then the LORD would have established your kingdom over Israel forever.
1SAM|13|14|But now your kingdom shall not continue. The LORD has sought out a man after his own heart, and the LORD has commanded him to be prince over his people, because you have not kept what the LORD commanded you."
1SAM|13|15|And Samuel arose and went up from Gilgal. The rest of the people went up after Saul to meet the army; they went up from Gilgal to Gibeah of Benjamin. And Saul numbered the people who were present with him, about six hundred men.
1SAM|13|16|And Saul and Jonathan his son and the people who were present with them stayed in Geba of Benjamin, but the Philistines encamped in Michmash.
1SAM|13|17|And raiders came out of the camp of the Philistines in three companies. One company turned toward Ophrah, to the land of Shual;
1SAM|13|18|another company turned toward Beth-horon; and another company turned toward the border that looks down on the valley of Zeboim toward the wilderness.
1SAM|13|19|Now there was no blacksmith to be found throughout all the land of Israel, for the Philistines said, "Lest the Hebrews make themselves swords or spears."
1SAM|13|20|But every one of the Israelites went down to the Philistines to sharpen his plowshare, his mattock, his axe, or his sickle,
1SAM|13|21|and the charge was two-thirds of a shekel for the plowshares and for the mattocks, and a third of a shekel for sharpening the axes and for setting the goads.
1SAM|13|22|So on the day of the battle there was neither sword nor spear found in the hand of any of the people with Saul and Jonathan, but Saul and Jonathan his son had them.
1SAM|13|23|And the garrison of the Philistines went out to the pass of Michmash.
1SAM|14|1|One day Jonathan the son of Saul said to the young man who carried his armor, "Come, let us go over to the Philistine garrison on the other side." But he did not tell his father.
1SAM|14|2|Saul was staying in the outskirts of Gibeah in the pomegranate cave at Migron. The people who were with him were about six hundred men,
1SAM|14|3|including Ahijah the son of Ahitub, Ichabod's brother, son of Phinehas, son of Eli, the priest of the LORD in Shiloh, wearing an ephod. And the people did not know that Jonathan had gone.
1SAM|14|4|Within the passes, by which Jonathan sought to go over to the Philistine garrison, there was a rocky crag on the one side and a rocky crag on the other side. The name of the one was Bozez, and the name of the other Seneh.
1SAM|14|5|The one crag rose on the north in front of Michmash, and the other on the south in front of Geba.
1SAM|14|6|Jonathan said to the young man who carried his armor, "Come, let us go over to the garrison of these uncircumcised. It may be that the LORD will work for us, for nothing can hinder the LORD from saving by many or by few."
1SAM|14|7|And his armor-bearer said to him, "Do all that is in your heart. Do as you wish. Behold, I am with you heart and soul."
1SAM|14|8|Then Jonathan said, "Behold, we will cross over to the men, and we will show ourselves to them.
1SAM|14|9|If they say to us, 'Wait until we come to you,' then we will stand still in our place, and we will not go up to them.
1SAM|14|10|But if they say, 'Come up to us,' then we will go up, for the LORD has given them into our hand. And this shall be the sign to us."
1SAM|14|11|So both of them showed themselves to the garrison of the Philistines. And the Philistines said, "Look, Hebrews are coming out of the holes where they have hidden themselves."
1SAM|14|12|And the men of the garrison hailed Jonathan and his armor-bearer and said, "Come up to us, and we will show you a thing." And Jonathan said to his armor-bearer, "Come up after me, for the LORD has given them into the hand of Israel."
1SAM|14|13|Then Jonathan climbed up on his hands and feet, and his armor-bearer after him. And they fell before Jonathan, and his armor-bearer killed them after him.
1SAM|14|14|And that first strike, which Jonathan and his armor-bearer made, killed about twenty men within as it were half a furrow's length in an acre of land.
1SAM|14|15|And there was a panic in the camp, in the field, and among all the people. The garrison and even the raiders trembled, the earth quaked, and it became a very great panic.
1SAM|14|16|And the watchmen of Saul in Gibeah of Benjamin looked, and behold, the multitude was dispersing here and there.
1SAM|14|17|Then Saul said to the people who were with him, "Count and see who has gone from us." And when they had counted, behold, Jonathan and his armor-bearer were not there.
1SAM|14|18|So Saul said to Ahijah, "Bring the ark of God here." For the ark of God went at that time with the people of Israel.
1SAM|14|19|Now while Saul was talking to the priest, the tumult in the camp of the Philistines increased more and more. So Saul said to the priest, "Withdraw your hand."
1SAM|14|20|Then Saul and all the people who were with him rallied and went into the battle. And behold, every Philistine's sword was against his fellow, and there was very great confusion.
1SAM|14|21|Now the Hebrews who had been with the Philistines before that time and who had gone up with them into the camp, even they also turned to be with the Israelites who were with Saul and Jonathan.
1SAM|14|22|Likewise, when all the men of Israel who had hidden themselves in the hill country of Ephraim heard that the Philistines were fleeing, they too followed hard after them in the battle.
1SAM|14|23|So the LORD saved Israel that day. And the battle passed beyond Beth-aven.
1SAM|14|24|And the men of Israel had been hard pressed that day, so Saul had laid an oath on the people, saying, "Cursed be the man who eats food until it is evening and I am avenged on my enemies." So none of the people had tasted food.
1SAM|14|25|Now when all the people came to the forest, behold, there was honey on the ground.
1SAM|14|26|And when the people entered the forest, behold, the honey was dropping, but no one put his hand to his mouth, for the people feared the oath.
1SAM|14|27|But Jonathan had not heard his father charge the people with the oath, so he put out the tip of the staff that was in his hand and dipped it in the honeycomb and put his hand to his mouth, and his eyes became bright.
1SAM|14|28|Then one of the people said, "Your father strictly charged the people with an oath, saying, 'Cursed be the man who eats food this day.'"And the people were faint.
1SAM|14|29|Then Jonathan said, "My father has troubled the land. See how my eyes have become bright because I tasted a little of this honey.
1SAM|14|30|How much better if the people had eaten freely today of the spoil of their enemies that they found. For now the defeat among the Philistines has not been great."
1SAM|14|31|They struck down the Philistines that day from Michmash to Aijalon. And the people were very faint.
1SAM|14|32|The people pounced on the spoil and took sheep and oxen and calves and slaughtered them on the ground. And the people ate them with the blood.
1SAM|14|33|Then they told Saul, "Behold, the people are sinning against the LORD by eating with the blood." And he said, "You have dealt treacherously; roll a great stone to me here."
1SAM|14|34|And Saul said, "Disperse yourselves among the people and say to them, 'Let every man bring his ox or his sheep and slaughter them here and eat, and do not sin against the LORD by eating with the blood.'"So every one of the people brought his ox with him that night and they slaughtered them there.
1SAM|14|35|And Saul built an altar to the LORD; it was the first altar that he built to the LORD.
1SAM|14|36|Then Saul said, "Let us go down after the Philistines by night and plunder them until the morning light; let us not leave a man of them." And they said, "Do whatever seems good to you." But the priest said, "Let us draw near to God here."
1SAM|14|37|And Saul inquired of God, "Shall I go down after the Philistines? Will you give them into the hand of Israel?" But he did not answer him that day.
1SAM|14|38|And Saul said, "Come here, all you leaders of the people, and know and see how this sin has arisen today.
1SAM|14|39|For as the LORD lives who saves Israel, though it be in Jonathan my son, he shall surely die." But there was not a man among all the people who answered him.
1SAM|14|40|Then he said to all Israel, "You shall be on one side, and I and Jonathan my son will be on the other side." And the people said to Saul, "Do what seems good to you."
1SAM|14|41|Therefore Saul said, "O LORD God of Israel, why have you not answered your servant this day? If this guilt is in me or in Jonathan my son, O LORD, God of Israel, give Urim. But if this guilt is in your people Israel, give Thummim." And Jonathan and Saul were taken, but the people escaped.
1SAM|14|42|Then Saul said, "Cast the lot between me and my son Jonathan." And Jonathan was taken.
1SAM|14|43|Then Saul said to Jonathan, "Tell me what you have done." And Jonathan told him, "I tasted a little honey with the tip of the staff that was in my hand. Here I am; I will die."
1SAM|14|44|And Saul said, "God do so to me and more also; you shall surely die, Jonathan."
1SAM|14|45|Then the people said to Saul, "Shall Jonathan die, who has worked this great salvation in Israel? Far from it! As the LORD lives, there shall not one hair of his head fall to the ground, for he has worked with God this day." So the people ransomed Jonathan, so that he did not die.
1SAM|14|46|Then Saul went up from pursuing the Philistines, and the Philistines went to their own place.
1SAM|14|47|When Saul had taken the kingship over Israel, he fought against all his enemies on every side, against Moab, against the Ammonites, against Edom, against the kings of Zobah, and against the Philistines. Wherever he turned he routed them.
1SAM|14|48|And he did valiantly and struck the Amalekites and delivered Israel out of the hands of those who plundered them.
1SAM|14|49|Now the sons of Saul were Jonathan, Ishvi, and Malchi-shua. And the names of his two daughters were these: the name of the firstborn was Merab, and the name of the younger Michal.
1SAM|14|50|And the name of Saul's wife was Ahinoam the daughter of Ahimaaz. And the name of the commander of his army was Abner the son of Ner, Saul's uncle.
1SAM|14|51|Kish was the father of Saul, and Ner the father of Abner was the son of Abiel.
1SAM|14|52|There was hard fighting against the Philistines all the days of Saul. And when Saul saw any strong man, or any valiant man, he attached him to himself.
1SAM|15|1|And Samuel said to Saul, "The LORD sent me to anoint you king over his people Israel; now therefore listen to the words of the LORD.
1SAM|15|2|Thus says the LORD of hosts, 'I have noted what Amalek did to Israel in opposing them on the way when they came up out of Egypt.
1SAM|15|3|Now go and strike Amalek and devote to destruction all that they have. Do not spare them, but kill both man and woman, child and infant, ox and sheep, camel and donkey.'"
1SAM|15|4|So Saul summoned the people and numbered them in Telaim, two hundred thousand men on foot, and ten thousand men of Judah.
1SAM|15|5|And Saul came to the city of Amalek and lay in wait in the valley.
1SAM|15|6|Then Saul said to the Kenites, "Go, depart; go down from among the Amalekites, lest I destroy you with them. For you showed kindness to all the people of Israel when they came up out of Egypt." So the Kenites departed from among the Amalekites.
1SAM|15|7|And Saul defeated the Amalekites from Havilah as far as Shur, which is east of Egypt.
1SAM|15|8|And he took Agag the king of the Amalekites alive and devoted to destruction all the people with the edge of the sword.
1SAM|15|9|But Saul and the people spared Agag and the best of the sheep and of the oxen and of the fattened calves and the lambs, and all that was good, and would not utterly destroy them. All that was despised and worthless they devoted to destruction.
1SAM|15|10|The word of the LORD came to Samuel:
1SAM|15|11|"I regret that I have made Saul king, for he has turned back from following me and has not performed my commandments." And Samuel was angry, and he cried to the LORD all night.
1SAM|15|12|And Samuel rose early to meet Saul in the morning. And it was told Samuel, "Saul came to Carmel, and behold, he set up a monument for himself and turned and passed on and went down to Gilgal."
1SAM|15|13|And Samuel came to Saul, and Saul said to him, "Blessed be you to the LORD. I have performed the commandment of the LORD."
1SAM|15|14|And Samuel said, "What then is this bleating of the sheep in my ears and the lowing of the oxen that I hear?"
1SAM|15|15|Saul said, "They have brought them from the Amalekites, for the people spared the best of the sheep and of the oxen to sacrifice to the LORD your God, and the rest we have devoted to destruction."
1SAM|15|16|Then Samuel said to Saul, "Stop! I will tell you what the LORD said to me this night." And he said to him, "Speak."
1SAM|15|17|And Samuel said, "Though you are little in your own eyes, are you not the head of the tribes of Israel? The LORD anointed you king over Israel.
1SAM|15|18|And the LORD sent you on a mission and said, 'Go, devote to destruction the sinners, the Amalekites, and fight against them until they are consumed.'
1SAM|15|19|Why then did you not obey the voice of the LORD? Why did you pounce on the spoil and do what was evil in the sight of the LORD?"
1SAM|15|20|And Saul said to Samuel, "I have obeyed the voice of the LORD. I have gone on the mission on which the LORD sent me. I have brought Agag the king of Amalek, and I have devoted the Amalekites to destruction.
1SAM|15|21|But the people took of the spoil, sheep and oxen, the best of the things devoted to destruction, to sacrifice to the LORD your God in Gilgal."
1SAM|15|22|And Samuel said, "Has the LORD as great delight in burnt offerings and sacrifices, as in obeying the voice of the LORD? Behold, to obey is better than sacrifice, and to listen than the fat of rams.
1SAM|15|23|For rebellion is as the sin of divination, and presumption is as iniquity and idolatry. Because you have rejected the word of the LORD, he has also rejected you from being king."
1SAM|15|24|Saul said to Samuel, "I have sinned, for I have transgressed the commandment of the LORD and your words, because I feared the people and obeyed their voice.
1SAM|15|25|Now therefore, please pardon my sin and return with me that I may worship the LORD."
1SAM|15|26|And Samuel said to Saul, "I will not return with you. For you have rejected the word of the LORD, and the LORD has rejected you from being king over Israel."
1SAM|15|27|As Samuel turned to go away, Saul seized the skirt of his robe, and it tore.
1SAM|15|28|And Samuel said to him, "The LORD has torn the kingdom of Israel from you this day and has given it to a neighbor of yours, who is better than you.
1SAM|15|29|And also the Glory of Israel will not lie or have regret, for he is not a man, that he should have regret."
1SAM|15|30|Then he said, "I have sinned; yet honor me now before the elders of my people and before Israel, and return with me, that I may bow before the LORD your God."
1SAM|15|31|So Samuel turned back after Saul, and Saul bowed before the LORD.
1SAM|15|32|Then Samuel said, "Bring here to me Agag the king of the Amalekites." And Agag came to him cheerfully. Agag said, "Surely the bitterness of death is past."
1SAM|15|33|And Samuel said, "As your sword has made women childless, so shall your mother be childless among women." And Samuel hacked Agag to pieces before the LORD in Gilgal.
1SAM|15|34|Then Samuel went to Ramah, and Saul went up to his house in Gibeah of Saul.
1SAM|15|35|And Samuel did not see Saul again until the day of his death, but Samuel grieved over Saul. And the LORD regretted that he had made Saul king over Israel.
1SAM|16|1|The LORD said to Samuel, "How long will you grieve over Saul, since I have rejected him from being king over Israel? Fill your horn with oil, and go. I will send you to Jesse the Bethlehemite, for I have provided for myself a king among his sons."
1SAM|16|2|And Samuel said, "How can I go? If Saul hears it, he will kill me." And the LORD said, "Take a heifer with you and say, 'I have come to sacrifice to the LORD.'
1SAM|16|3|And invite Jesse to the sacrifice, and I will show you what you shall do. And you shall anoint for me him whom I declare to you."
1SAM|16|4|Samuel did what the LORD commanded and came to Bethlehem. The elders of the city came to meet him trembling and said, "Do you come peaceably?"
1SAM|16|5|And he said, "Peaceably; I have come to sacrifice to the LORD. Consecrate yourselves, and come with me to the sacrifice." And he consecrated Jesse and his sons and invited them to the sacrifice.
1SAM|16|6|When they came, he looked on Eliab and thought, "Surely the LORD's anointed is before him."
1SAM|16|7|But the LORD said to Samuel, "Do not look on his appearance or on the height of his stature, because I have rejected him. For the LORD sees not as man sees: man looks on the outward appearance, but the LORD looks on the heart."
1SAM|16|8|Then Jesse called Abinadab and made him pass before Samuel. And he said, "Neither has the LORD chosen this one."
1SAM|16|9|Then Jesse made Shammah pass by. And he said, "Neither has the LORD chosen this one."
1SAM|16|10|And Jesse made seven of his sons pass before Samuel. And Samuel said to Jesse, "The LORD has not chosen these."
1SAM|16|11|Then Samuel said to Jesse, "Are all your sons here?" And he said, "There remains yet the youngest, but behold, he is keeping the sheep." And Samuel said to Jesse, "Send and get him, for we will not sit down till he comes here."
1SAM|16|12|And he sent and brought him in. Now he was ruddy and had beautiful eyes and was handsome. And the LORD said, "Arise, anoint him, for this is he."
1SAM|16|13|Then Samuel took the horn of oil and anointed him in the midst of his brothers. And the Spirit of the LORD rushed upon David from that day forward. And Samuel rose up and went to Ramah.
1SAM|16|14|Now the Spirit of the LORD departed from Saul, and an evil spirit from the LORD tormented him.
1SAM|16|15|And Saul's servants said to him, "Behold now, an evil spirit from God is tormenting you.
1SAM|16|16|Let our lord now command your servants who are before you to seek out a man who is skillful in playing the lyre, and when the evil spirit from God is upon you, he will play it, and you will be well."
1SAM|16|17|So Saul said to his servants, "Provide for me a man who can play well and bring him to me."
1SAM|16|18|One of the young men answered, "Behold, I have seen a son of Jesse the Bethlehemite, who is skillful in playing, a man of valor, a man of war, prudent in speech, and a man of good presence, and the LORD is with him."
1SAM|16|19|Therefore Saul sent messengers to Jesse and said, "Send me David your son, who is with the sheep."
1SAM|16|20|And Jesse took a donkey laden with bread and a skin of wine and a young goat and sent them by David his son to Saul.
1SAM|16|21|And David came to Saul and entered his service. And Saul loved him greatly, and he became his armor-bearer.
1SAM|16|22|And Saul sent to Jesse, saying, "Let David remain in my service, for he has found favor in my sight."
1SAM|16|23|And whenever the evil spirit from God was upon Saul, David took the lyre and played it with his hand. So Saul was refreshed and was well, and the evil spirit departed from him.
1SAM|17|1|Now the Philistines gathered their armies for battle. And they were gathered at Socoh, which belongs to Judah, and encamped between Socoh and Azekah, in Ephes-dammim.
1SAM|17|2|And Saul and the men of Israel were gathered, and encamped in the Valley of Elah, and drew up in line of battle against the Philistines.
1SAM|17|3|And the Philistines stood on the mountain on the one side, and Israel stood on the mountain on the other side, with a valley between them.
1SAM|17|4|And there came out from the camp of the Philistines a champion named Goliath of Gath, whose height was six cubits and a span.
1SAM|17|5|He had a helmet of bronze on his head, and he was armed with a coat of mail, and the weight of the coat was five thousand shekels of bronze.
1SAM|17|6|And he had bronze armor on his legs, and a javelin of bronze slung between his shoulders.
1SAM|17|7|The shaft of his spear was like a weaver's beam, and his spear's head weighed six hundred shekels of iron. And his shield-bearer went before him.
1SAM|17|8|He stood and shouted to the ranks of Israel, "Why have you come out to draw up for battle? Am I not a Philistine, and are you not servants of Saul? Choose a man for yourselves, and let him come down to me.
1SAM|17|9|If he is able to fight with me and kill me, then we will be your servants. But if I prevail against him and kill him, then you shall be our servants and serve us."
1SAM|17|10|And the Philistine said, "I defy the ranks of Israel this day. Give me a man, that we may fight together."
1SAM|17|11|When Saul and all Israel heard these words of the Philistine, they were dismayed and greatly afraid.
1SAM|17|12|Now David was the son of an Ephrathite of Bethlehem in Judah, named Jesse, who had eight sons. In the days of Saul the man was already old and advanced in years.
1SAM|17|13|The three oldest sons of Jesse had followed Saul to the battle. And the names of his three sons who went to the battle were Eliab the firstborn, and next to him Abinadab, and the third Shammah.
1SAM|17|14|David was the youngest. The three eldest followed Saul,
1SAM|17|15|but David went back and forth from Saul to feed his father's sheep at Bethlehem.
1SAM|17|16|For forty days the Philistine came forward and took his stand, morning and evening.
1SAM|17|17|And Jesse said to David his son, "Take for your brothers an ephah of this parched grain, and these ten loaves, and carry them quickly to the camp to your brothers.
1SAM|17|18|Also take these ten cheeses to the commander of their thousand. See if your brothers are well, and bring some token from them."
1SAM|17|19|Now Saul and they and all the men of Israel were in the valley of Elah, fighting with the Philistines.
1SAM|17|20|And David rose early in the morning and left the sheep with a keeper and took the provisions and went, as Jesse had commanded him. And he came to the encampment as the host was going out to the battle line, shouting the war cry.
1SAM|17|21|And Israel and the Philistines drew up for battle, army against army.
1SAM|17|22|And David left the things in charge of the keeper of the baggage and ran to the ranks and went and greeted his brothers.
1SAM|17|23|As he talked with them, behold, the champion, the Philistine of Gath, Goliath by name, came up out of the ranks of the Philistines and spoke the same words as before. And David heard him.
1SAM|17|24|All the men of Israel, when they saw the man, fled from him and were much afraid.
1SAM|17|25|And the men of Israel said, "Have you seen this man who has come up? Surely he has come up to defy Israel. And the king will enrich the man who kills him with great riches and will give him his daughter and make his father's house free in Israel."
1SAM|17|26|And David said to the men who stood by him, "What shall be done for the man who kills this Philistine and takes away the reproach from Israel? For who is this uncircumcised Philistine, that he should defy the armies of the living God?"
1SAM|17|27|And the people answered him in the same way, "So shall it be done to the man who kills him."
1SAM|17|28|Now Eliab his eldest brother heard when he spoke to the men. And Eliab's anger was kindled against David, and he said, "Why have you come down? And with whom have you left those few sheep in the wilderness? I know your presumption and the evil of your heart, for you have come down to see the battle."
1SAM|17|29|And David said, "What have I done now? Was it not but a word?"
1SAM|17|30|And he turned away from him toward another, and spoke in the same way, and the people answered him again as before.
1SAM|17|31|When the words that David spoke were heard, they repeated them before Saul, and he sent for him.
1SAM|17|32|And David said to Saul, "Let no man's heart fail because of him. Your servant will go and fight with this Philistine."
1SAM|17|33|And Saul said to David, "You are not able to go against this Philistine to fight with him, for you are but a youth, and he has been a man of war from his youth."
1SAM|17|34|But David said to Saul, "Your servant used to keep sheep for his father. And when there came a lion, or a bear, and took a lamb from the flock,
1SAM|17|35|I went after him and struck him and delivered it out of his mouth. And if he arose against me, I caught him by his beard and struck him and killed him.
1SAM|17|36|Your servant has struck down both lions and bears, and this uncircumcised Philistine shall be like one of them, for he has defied the armies of the living God."
1SAM|17|37|And David said, "The LORD who delivered me from the paw of the lion and from the paw of the bear will deliver me from the hand of this Philistine." And Saul said to David, "Go, and the LORD be with you!"
1SAM|17|38|Then Saul clothed David with his armor. He put a helmet of bronze on his head and clothed him with a coat of mail,
1SAM|17|39|and David strapped his sword over his armor. And he tried in vain to go, for he had not tested them. Then David said to Saul, "I cannot go with these, for I have not tested them." So David put them off.
1SAM|17|40|Then he took his staff in his hand and chose five smooth stones from the brook and put them in his shepherd's pouch. His sling was in his hand, and he approached the Philistine.
1SAM|17|41|And the Philistine moved forward and came near to David, with his shield-bearer in front of him.
1SAM|17|42|And when the Philistine looked and saw David, he disdained him, for he was but a youth, ruddy and handsome in appearance.
1SAM|17|43|And the Philistine said to David, "Am I a dog, that you come to me with sticks?" And the Philistine cursed David by his gods.
1SAM|17|44|The Philistine said to David, "Come to me, and I will give your flesh to the birds of the air and to the beasts of the field."
1SAM|17|45|Then David said to the Philistine, "You come to me with a sword and with a spear and with a javelin, but I come to you in the name of the LORD of hosts, the God of the armies of Israel, whom you have defied.
1SAM|17|46|This day the LORD will deliver you into my hand, and I will strike you down and cut off your head. And I will give the dead bodies of the host of the Philistines this day to the birds of the air and to the wild beasts of the earth, that all the earth may know that there is a God in Israel,
1SAM|17|47|and that all this assembly may know that the LORD saves not with sword and spear. For the battle is the LORD's, and he will give you into our hand."
1SAM|17|48|When the Philistine arose and came and drew near to meet David, David ran quickly toward the battle line to meet the Philistine.
1SAM|17|49|And David put his hand in his bag and took out a stone and slung it and struck the Philistine on his forehead. The stone sank into his forehead, and he fell on his face to the ground.
1SAM|17|50|So David prevailed over the Philistine with a sling and with a stone, and struck the Philistine and killed him. There was no sword in the hand of David.
1SAM|17|51|Then David ran and stood over the Philistine and took his sword and drew it out of its sheath and killed him and cut off his head with it. When the Philistines saw that their champion was dead, they fled.
1SAM|17|52|And the men of Israel and Judah rose with a shout and pursued the Philistines as far as Gath and the gates of Ekron, so that the wounded Philistines fell on the way from Shaaraim as far as Gath and Ekron.
1SAM|17|53|And the people of Israel came back from chasing the Philistines, and they plundered their camp.
1SAM|17|54|And David took the head of the Philistine and brought it to Jerusalem, but he put his armor in his tent.
1SAM|17|55|As soon as Saul saw David go out against the Philistine, he said to Abner, the commander of the army, "Abner, whose son is this youth?" And Abner said, "As your soul lives, O king, I do not know."
1SAM|17|56|And the king said, "Inquire whose son the boy is."
1SAM|17|57|And as soon as David returned from the striking down of the Philistine, Abner took him, and brought him before Saul with the head of the Philistine in his hand.
1SAM|17|58|And Saul said to him, "Whose son are you, young man?" And David answered, "I am the son of your servant Jesse the Bethlehemite."
1SAM|18|1|As soon as he had finished speaking to Saul, the soul of Jonathan was knit to the soul of David, and Jonathan loved him as his own soul.
1SAM|18|2|And Saul took him that day and would not let him return to his father's house.
1SAM|18|3|Then Jonathan made a covenant with David, because he loved him as his own soul.
1SAM|18|4|And Jonathan stripped himself of the robe that was on him and gave it to David, and his armor, and even his sword and his bow and his belt.
1SAM|18|5|And David went out and was successful wherever Saul sent him, so that Saul set him over the men of war. And this was good in the sight of all the people and also in the sight of Saul's servants.
1SAM|18|6|As they were coming home, when David returned from striking down the Philistine, the women came out of all the cities of Israel, singing and dancing, to meet King Saul, with tambourines, with songs of joy, and with musical instruments.
1SAM|18|7|And the women sang to one another as they celebrated, "Saul has struck down his thousands, and David his ten thousands."
1SAM|18|8|And Saul was very angry, and this saying displeased him. He said, "They have ascribed to David ten thousands, and to me they have ascribed thousands, and what more can he have but the kingdom?"
1SAM|18|9|And Saul eyed David from that day on.
1SAM|18|10|The next day a harmful spirit from God rushed upon Saul, and he raved within his house while David was playing the lyre, as he did day by day. Saul had his spear in his hand.
1SAM|18|11|And Saul hurled the spear, for he thought, "I will pin David to the wall." But David evaded him twice.
1SAM|18|12|Saul was afraid of David because the LORD was with him but had departed from Saul.
1SAM|18|13|So Saul removed him from his presence and made him a commander of a thousand. And he went out and came in before the people.
1SAM|18|14|And David had success in all his undertakings, for the LORD was with him.
1SAM|18|15|And when Saul saw that he had great success, he stood in fearful awe of him.
1SAM|18|16|But all Israel and Judah loved David, for he went out and came in before them.
1SAM|18|17|Then Saul said to David, "Here is my elder daughter Merab. I will give her to you for a wife. Only be valiant for me and fight the LORD's battles." For Saul thought, "Let not my hand be against him, but let the hand of the Philistines be against him."
1SAM|18|18|And David said to Saul, "Who am I, and who are my relatives, my father's clan in Israel, that I should be son-in-law to the king?"
1SAM|18|19|But at the time when Merab, Saul's daughter, should have been given to David, she was given to Adriel the Meholathite for a wife.
1SAM|18|20|Now Saul's daughter Michal loved David. And they told Saul, and the thing pleased him.
1SAM|18|21|Saul thought, "Let me give her to him, that she may be a snare for him and that the hand of the Philistines may be against him." Therefore Saul said to David a second time, "You shall now be my son-in-law."
1SAM|18|22|And Saul commanded his servants, "Speak to David in private and say, 'Behold, the king has delight in you, and all his servants love you. Now then become the king's son-in-law.'"
1SAM|18|23|And Saul's servants spoke those words in the ears of David. And David said, "Does it seem to you a little thing to become the king's son-in-law, since I am a poor man and have no reputation?"
1SAM|18|24|And the servants of Saul told him, "Thus and so did David speak."
1SAM|18|25|Then Saul said, "Thus shall you say to David, 'The king desires no bride-price except a hundred foreskins of the Philistines, that he may be avenged of the king's enemies.'"Now Saul thought to make David fall by the hand of the Philistines.
1SAM|18|26|And when his servants told David these words, it pleased David well to be the king's son-in-law. Before the time had expired,
1SAM|18|27|David arose and went, along with his men, and killed two hundred of the Philistines. And David brought their foreskins, which were given in full number to the king, that he might become the king's son-in-law. And Saul gave him his daughter Michal for a wife.
1SAM|18|28|But when Saul saw and knew that the LORD was with David, and that Michal, Saul's daughter, loved him,
1SAM|18|29|Saul was even more afraid of David. So Saul was David's enemy continually.
1SAM|18|30|Then the princes of the Philistines came out to battle, and as often as they came out David had more success than all the servants of Saul, so that his name was highly esteemed.
1SAM|19|1|And Saul spoke to Jonathan his son and to all his servants, that they should kill David. But Jonathan, Saul's son, delighted much in David.
1SAM|19|2|And Jonathan told David, "Saul my father seeks to kill you. Therefore be on your guard in the morning. Stay in a secret place and hide yourself.
1SAM|19|3|And I will go out and stand beside my father in the field where you are, and I will speak to my father about you. And if I learn anything I will tell you."
1SAM|19|4|And Jonathan spoke well of David to Saul his father and said to him, "Let not the king sin against his servant David, because he has not sinned against you, and because his deeds have brought good to you.
1SAM|19|5|For he took his life in his hand and he struck down the Philistine, and the LORD worked a great salvation for all Israel. You saw it, and rejoiced. Why then will you sin against innocent blood by killing David without cause?"
1SAM|19|6|And Saul listened to the voice of Jonathan. Saul swore, "As the LORD lives, he shall not be put to death."
1SAM|19|7|And Jonathan called David, and Jonathan reported to him all these things. And Jonathan brought David to Saul, and he was in his presence as before.
1SAM|19|8|And there was war again. And David went out and fought with the Philistines and struck them with a great blow, so that they fled before him.
1SAM|19|9|Then a harmful spirit from the LORD came upon Saul, as he sat in his house with his spear in his hand. And David was playing the lyre.
1SAM|19|10|And Saul sought to pin David to the wall with the spear, but he eluded Saul, so that he struck the spear into the wall. And David fled and escaped that night.
1SAM|19|11|Saul sent messengers to David's house to watch him, that he might kill him in the morning. But Michal, David's wife, told him, "If you do not escape with your life tonight, tomorrow you will be killed."
1SAM|19|12|So Michal let David down through the window, and he fled away and escaped.
1SAM|19|13|Michal took an image and laid it on the bed and put a pillow of goats' hair at its head and covered it with the clothes.
1SAM|19|14|And when Saul sent messengers to take David, she said, "He is sick."
1SAM|19|15|Then Saul sent the messengers to see David, saying, "Bring him up to me in the bed, that I may kill him."
1SAM|19|16|And when the messengers came in, behold, the image was in the bed, with the pillow of goats' hair at its head.
1SAM|19|17|Saul said to Michal, "Why have you deceived me thus and let my enemy go, so that he has escaped?" And Michal answered Saul, "He said to me, 'Let me go. Why should I kill you?'"
1SAM|19|18|Now David fled and escaped, and he came to Samuel at Ramah and told him all that Saul had done to him. And he and Samuel went and lived at Naioth.
1SAM|19|19|And it was told Saul, "Behold, David is at Naioth in Ramah."
1SAM|19|20|Then Saul sent messengers to take David, and when they saw the company of the prophets prophesying, and Samuel standing as head over them, the Spirit of God came upon the messengers of Saul, and they also prophesied.
1SAM|19|21|When it was told Saul, he sent other messengers, and they also prophesied. And Saul sent messengers again the third time, and they also prophesied.
1SAM|19|22|Then he himself went to Ramah and came to the great well that is in Secu. And he asked, "Where are Samuel and David?" And one said, "Behold, they are at Naioth in Ramah."
1SAM|19|23|And he went there to Naioth in Ramah. And the Spirit of God came upon him also, and as he went he prophesied until he came to Naioth in Ramah.
1SAM|19|24|And he too stripped off his clothes, and he too prophesied before Samuel and lay naked all that day and all that night. Thus it is said, "Is Saul also among the prophets?"
1SAM|20|1|Then David fled from Naioth in Ramah and came and said before Jonathan, "What have I done? What is my guilt? And what is my sin before your father, that he seeks my life?"
1SAM|20|2|And he said to him, "Far from it! You shall not die. Behold, my father does nothing either great or small without disclosing it to me. And why should my father hide this from me? It is not so."
1SAM|20|3|But David vowed again, saying, "Your father knows well that I have found favor in your eyes, and he thinks, 'Do not let Jonathan know this, lest he be grieved.' But truly, as the LORD lives and as your soul lives, there is but a step between me and death."
1SAM|20|4|Then Jonathan said to David, "Whatever you say, I will do for you."
1SAM|20|5|David said to Jonathan, "Behold, tomorrow is the new moon, and I should not fail to sit at table with the king. But let me go, that I may hide myself in the field till the third day at evening.
1SAM|20|6|If your father misses me at all, then say, 'David earnestly asked leave of me to run to Bethlehem his city, for there is a yearly sacrifice there for all the clan.'
1SAM|20|7|If he says, 'Good!' it will be well with your servant, but if he is angry, then know that harm is determined by him.
1SAM|20|8|Therefore deal kindly with your servant, for you have brought your servant into a covenant of the LORD with you. But if there is guilt in me, kill me yourself, for why should you bring me to your father?"
1SAM|20|9|And Jonathan said, "Far be it from you! If I knew that it was determined by my father that harm should come to you, would I not tell you?"
1SAM|20|10|Then David said to Jonathan, "Who will tell me if your father answers you roughly?"
1SAM|20|11|And Jonathan said to David, "Come, let us go out into the field." So they both went out into the field.
1SAM|20|12|And Jonathan said to David, "The LORD, the God of Israel, be witness! When I have sounded out my father, about this time tomorrow, or the third day, behold, if he is well disposed toward David, shall I not then send and disclose it to you?
1SAM|20|13|But should it please my father to do you harm, the LORD do so to Jonathan and more also if I do not disclose it to you and send you away, that you may go in safety. May the LORD be with you, as he has been with my father.
1SAM|20|14|If I am still alive, show me the steadfast love of the LORD, that I may not die;
1SAM|20|15|and do not cut off your steadfast love from my house forever, when the LORD cuts off every one of the enemies of David from the face of the earth."
1SAM|20|16|And Jonathan made a covenant with the house of David, saying, "May the LORD take vengeance on David's enemies."
1SAM|20|17|And Jonathan made David swear again by his love for him, for he loved him as he loved his own soul.
1SAM|20|18|Then Jonathan said to him, "Tomorrow is the new moon, and you will be missed, because your seat will be empty.
1SAM|20|19|On the third day go down quickly to the place where you hid yourself when the matter was in hand, and remain beside the stone heap.
1SAM|20|20|And I will shoot three arrows to the side of it, as though I shot at a mark.
1SAM|20|21|And behold, I will send the young man, saying, 'Go, find the arrows.' If I say to the young man, 'Look, the arrows are on this side of you, take them,' then you are to come, for, as the LORD lives, it is safe for you and there is no danger.
1SAM|20|22|But if I say to the youth, 'Look, the arrows are beyond you,' then go, for the LORD has sent you away.
1SAM|20|23|And as for the matter of which you and I have spoken, behold, the LORD is between you and me forever."
1SAM|20|24|So David hid himself in the field. And when the new moon came, the king sat down to eat food.
1SAM|20|25|The king sat on his seat, as at other times, on the seat by the wall. Jonathan sat opposite, and Abner sat by Saul's side, but David's place was empty.
1SAM|20|26|Yet Saul did not say anything that day, for he thought, "Something has happened to him. He is not clean; surely he is not clean."
1SAM|20|27|But on the second day, the day after the new moon, David's place was empty. And Saul said to Jonathan his son, "Why has not the son of Jesse come to the meal, either yesterday or today?"
1SAM|20|28|Jonathan answered Saul, "David earnestly asked leave of me to go to Bethlehem.
1SAM|20|29|He said, 'Let me go, for our clan holds a sacrifice in the city, and my brother has commanded me to be there. So now, if I have found favor in your eyes, let me get away and see my brothers.' For this reason he has not come to the king's table."
1SAM|20|30|Then Saul's anger was kindled against Jonathan, and he said to him, "You son of a perverse, rebellious woman, do I not know that you have chosen the son of Jesse to your own shame, and to the shame of your mother's nakedness?
1SAM|20|31|For as long as the son of Jesse lives on the earth, neither you nor your kingdom shall be established. Therefore send and bring him to me, for he shall surely die."
1SAM|20|32|Then Jonathan answered Saul his father, "Why should he be put to death? What has he done?"
1SAM|20|33|But Saul hurled his spear at him to strike him. So Jonathan knew that his father was determined to put David to death.
1SAM|20|34|And Jonathan rose from the table in fierce anger and ate no food the second day of the month, for he was grieved for David, because his father had disgraced him.
1SAM|20|35|In the morning Jonathan went out into the field to the appointment with David, and with him a little boy.
1SAM|20|36|And he said to his boy, "Run and find the arrows that I shoot." As the boy ran, he shot an arrow beyond him.
1SAM|20|37|And when the boy came to the place of the arrow that Jonathan had shot, Jonathan called after the boy and said, "Is not the arrow beyond you?"
1SAM|20|38|And Jonathan called after the boy, "Hurry! Be quick! Do not stay!" So Jonathan's boy gathered up the arrows and came to his master.
1SAM|20|39|But the boy knew nothing. Only Jonathan and David knew the matter.
1SAM|20|40|And Jonathan gave his weapons to his boy and said to him, "Go and carry them to the city."
1SAM|20|41|And as soon as the boy had gone, David rose from beside the stone heap and fell on his face to the ground and bowed three times. And they kissed one another and wept with one another, David weeping the most.
1SAM|20|42|Then Jonathan said to David, "Go in peace, because we have sworn both of us in the name of the LORD, saying, 'The LORD shall be between me and you, and between my offspring and your offspring, forever.'"And he rose and departed, and Jonathan went into the city.
1SAM|21|1|Then David came to Nob to Ahimelech the priest. And Ahimelech came to meet David trembling and said to him, "Why are you alone, and no one with you?"
1SAM|21|2|And David said to Ahimelech the priest, "The king has charged me with a matter and said to me, 'Let no one know anything of the matter about which I send you, and with which I have charged you.' I have made an appointment with the young men for such and such a place.
1SAM|21|3|Now then, what do you have on hand? Give me five loaves of bread, or whatever is here."
1SAM|21|4|And the priest answered David, "I have no common bread on hand, but there is holy bread- if the young men have kept themselves from women."
1SAM|21|5|And David answered the priest, "Truly women have been kept from us as always when I go on an expedition. The vessels of the young men are holy even when it is an ordinary journey. How much more today will their vessels be holy?"
1SAM|21|6|So the priest gave him the holy bread, for there was no bread there but the bread of the Presence, which is removed from before the LORD, to be replaced by hot bread on the day it is taken away.
1SAM|21|7|Now a certain man of the servants of Saul was there that day, detained before the LORD. His name was Doeg the Edomite, the chief of Saul's herdsmen.
1SAM|21|8|Then David said to Ahimelech, "Then have you not here a spear or a sword at hand? For I have brought neither my sword nor my weapons with me, because the king's business required haste."
1SAM|21|9|And the priest said, "The sword of Goliath the Philistine, whom you struck down in the valley of Elah, behold, it is here wrapped in a cloth behind the ephod. If you will take that, take it, for there is none but that here." And David said, "There is none like that; give it to me."
1SAM|21|10|And David rose and fled that day from Saul and went to Achish the king of Gath.
1SAM|21|11|And the servants of Achish said to him, "Is not this David the king of the land? Did they not sing to one another of him in dances, 'Saul has struck down his thousands, and David his ten thousands'?"
1SAM|21|12|And David took these words to heart and was much afraid of Achish the king of Gath.
1SAM|21|13|So he changed his behavior before them and pretended to be insane in their hands and made marks on the doors of the gate and let his spittle run down his beard.
1SAM|21|14|Then Achish said to his servants, "Behold, you see the man is mad. Why then have you brought him to me?
1SAM|21|15|Do I lack madmen, that you have brought this fellow to behave as a madman in my presence? Shall this fellow come into my house?"
1SAM|22|1|David departed from there and escaped to the cave of Adullam. And when his brothers and all his father's house heard it, they went down there to him.
1SAM|22|2|And everyone who was in distress, and everyone who was in debt, and everyone who was bitter in soul, gathered to him. And he became captain over them. And there were with him about four hundred men.
1SAM|22|3|And David went from there to Mizpeh of Moab. And he said to the king of Moab, "Please let my father and my mother stay with you, till I know what God will do for me."
1SAM|22|4|And he left them with the king of Moab, and they stayed with him all the time that David was in the stronghold.
1SAM|22|5|Then the prophet Gad said to David, "Do not remain in the stronghold; depart, and go into the land of Judah." So David departed and went into the forest of Hereth.
1SAM|22|6|Now Saul heard that David was discovered, and the men who were with him. Saul was sitting at Gibeah under the tamarisk tree on the height with his spear in his hand, and all his servants were standing about him.
1SAM|22|7|And Saul said to his servants who stood about him, "Hear now, people of Benjamin; will the son of Jesse give every one of you fields and vineyards, will he make you all commanders of thousands and commanders of hundreds,
1SAM|22|8|that all of you have conspired against me? No one discloses to me when my son makes a covenant with the son of Jesse. None of you is sorry for me or discloses to me that my son has stirred up my servant against me, to lie in wait, as at this day."
1SAM|22|9|Then answered Doeg the Edomite, who stood by the servants of Saul, "I saw the son of Jesse coming to Nob, to Ahimelech the son of Ahitub,
1SAM|22|10|and he inquired of the LORD for him and gave him provisions and gave him the sword of Goliath the Philistine."
1SAM|22|11|Then the king sent to summon Ahimelech the priest, the son of Ahitub, and all his father's house, the priests who were at Nob, and all of them came to the king.
1SAM|22|12|And Saul said, "Hear now, son of Ahitub." And he answered, "Here I am, my lord."
1SAM|22|13|And Saul said to him, "Why have you conspired against me, you and the son of Jesse, in that you have given him bread and a sword and have inquired of God for him, so that he has risen against me, to lie in wait, as at this day?"
1SAM|22|14|Then Ahimelech answered the king, "And who among all your servants is so faithful as David, who is the king's son-in-law, and captain over your bodyguard, and honored in your house?
1SAM|22|15|Is today the first time that I have inquired of God for him? No! Let not the king impute anything to his servant or to all the house of my father, for your servant has known nothing of all this, much or little."
1SAM|22|16|And the king said, "You shall surely die, Ahimelech, you and all your father's house."
1SAM|22|17|And the king said to the guard who stood about him, "Turn and kill the priests of the LORD, because their hand also is with David, and they knew that he fled and did not disclose it to me." But the servants of the king would not put out their hand to strike the priests of the LORD.
1SAM|22|18|Then the king said to Doeg, "You turn and strike the priests." And Doeg the Edomite turned and struck down the priests, and he killed on that day eighty-five persons who wore the linen ephod.
1SAM|22|19|And Nob, the city of the priests, he put to the sword; both man and woman, child and infant, ox, donkey and sheep, he put to the sword.
1SAM|22|20|But one of the sons of Ahimelech the son of Ahitub, named Abiathar, escaped and fled after David.
1SAM|22|21|And Abiathar told David that Saul had killed the priests of the LORD.
1SAM|22|22|And David said to Abiathar, "I knew on that day, when Doeg the Edomite was there, that he would surely tell Saul. I have occasioned the death of all the persons of your father's house.
1SAM|22|23|Stay with me; do not be afraid, for he who seeks my life seeks your life. With me you shall be in safekeeping."
1SAM|23|1|Now they told David, "Behold, the Philistines are fighting against Keilah and are robbing the threshing floors."
1SAM|23|2|Therefore David inquired of the LORD, "Shall I go and attack these Philistines?" And the LORD said to David, "Go and attack the Philistines and save Keilah."
1SAM|23|3|But David's men said to him, "Behold, we are afraid here in Judah; how much more then if we go to Keilah against the armies of the Philistines?"
1SAM|23|4|Then David inquired of the LORD again. And the LORD answered him, "Arise, go down to Keilah, for I will give the Philistines into your hand."
1SAM|23|5|And David and his men went to Keilah and fought with the Philistines and brought away their livestock and struck them with a great blow. So David saved the inhabitants of Keilah.
1SAM|23|6|When Abiathar the son of Ahimelech had fled to David to Keilah, he had come down with an ephod in his hand.
1SAM|23|7|Now it was told Saul that David had come to Keilah. And Saul said, "God has given him into my hand, for he has shut himself in by entering a town that has gates and bars."
1SAM|23|8|And Saul summoned all the people to war, to go down to Keilah, to besiege David and his men.
1SAM|23|9|David knew that Saul was plotting harm against him. And he said to Abiathar the priest, "Bring the ephod here."
1SAM|23|10|Then said David, "O LORD, the God of Israel, your servant has surely heard that Saul seeks to come to Keilah, to destroy the city on my account.
1SAM|23|11|Will the men of Keilah surrender me into his hand? Will Saul come down, as your servant has heard? O LORD, the God of Israel, please tell your servant." And the LORD said, "He will come down."
1SAM|23|12|Then David said, "Will the men of Keilah surrender me and my men into the hand of Saul?" And the LORD said, "They will surrender you."
1SAM|23|13|Then David and his men, who were about six hundred, arose and departed from Keilah, and they went wherever they could go. When Saul was told that David had escaped from Keilah, he gave up the expedition.
1SAM|23|14|And David remained in the strongholds in the wilderness, in the hill country of the Wilderness of Ziph. And Saul sought him every day, but God did not give him into his hand.
1SAM|23|15|David saw that Saul had come out to seek his life. David was in the Wilderness of Ziph at Horesh.
1SAM|23|16|And Jonathan, Saul's son, rose and went to David at Horesh, and strengthened his hand in God.
1SAM|23|17|And he said to him, "Do not fear, for the hand of Saul my father shall not find you. You shall be king over Israel, and I shall be next to you. Saul my father also knows this."
1SAM|23|18|And the two of them made a covenant before the LORD. David remained at Horesh, and Jonathan went home.
1SAM|23|19|Then the Ziphites went up to Saul at Gibeah, saying, "Is not David hiding among us in the strongholds at Horesh, on the hill of Hachilah, which is south of Jeshimon?
1SAM|23|20|Now come down, O king, according to all your heart's desire to come down, and our part shall be to surrender him into the king's hand."
1SAM|23|21|And Saul said, "May you be blessed by the LORD, for you have had compassion on me.
1SAM|23|22|Go, make yet more sure. Know and see the place where his foot is, and who has seen him there, for it is told me that he is very cunning.
1SAM|23|23|See therefore and take note of all the lurking places where he hides, and come back to me with sure information. Then I will go with you. And if he is in the land, I will search him out among all the thousands of Judah."
1SAM|23|24|And they arose and went to Ziph ahead of Saul. Now David and his men were in the wilderness of Maon, in the Arabah to the south of Jeshimon.
1SAM|23|25|And Saul and his men went to seek him. And David was told, so he went down to the rock and lived in the wilderness of Maon. And when Saul heard that, he pursued after David in the wilderness of Maon.
1SAM|23|26|Saul went on one side of the mountain, and David and his men on the other side of the mountain. And David was hurrying to get away from Saul. As Saul and his men were closing in on David and his men to capture them,
1SAM|23|27|a messenger came to Saul, saying, "Hurry and come, for the Philistines have made a raid against the land."
1SAM|23|28|So Saul returned from pursuing after David and went against the Philistines. Therefore that place was called the Rock of Escape.
1SAM|23|29|And David went up from there and lived in the strongholds of Engedi.
1SAM|24|1|When Saul returned from fol- lowing the Philistines, he was told, "Behold, David is in the wilderness of Engedi."
1SAM|24|2|Then Saul took three thousand chosen men out of all Israel and went to seek David and his men in front of the Wildgoats' Rocks.
1SAM|24|3|And he came to the sheepfolds by the way, where there was a cave, and Saul went in to relieve himself. Now David and his men were sitting in the innermost parts of the cave.
1SAM|24|4|And the men of David said to him, "Here is the day of which the LORD said to you, 'Behold, I will give your enemy into your hand, and you shall do to him as it shall seem good to you.'"Then David arose and stealthily cut off a corner of Saul's robe.
1SAM|24|5|And afterward David's heart struck him, because he had cut off a corner of Saul's robe.
1SAM|24|6|He said to his men, "The LORD forbid that I should do this thing to my lord, the LORD's anointed, to put out my hand against him, seeing he is the LORD's anointed."
1SAM|24|7|So David persuaded his men with these words and did not permit them to attack Saul. And Saul rose up and left the cave and went on his way.
1SAM|24|8|Afterward David also arose and went out of the cave, and called after Saul, "My lord the king!" And when Saul looked behind him, David bowed with his face to the earth and paid homage.
1SAM|24|9|And David said to Saul, "Why do you listen to the words of men who say, 'Behold, David seeks your harm'?
1SAM|24|10|Behold, this day your eyes have seen how the LORD gave you today into my hand in the cave. And some told me to kill you, but I spared you. I said, 'I will not put out my hand against my lord, for he is the LORD's anointed.'
1SAM|24|11|See, my father, see the corner of your robe in my hand. For by the fact that I cut off the corner of your robe and did not kill you, you may know and see that there is no wrong or treason in my hands. I have not sinned against you, though you hunt my life to take it.
1SAM|24|12|May the LORD judge between me and you, may the LORD avenge me against you, but my hand shall not be against you.
1SAM|24|13|As the proverb of the ancients says, 'Out of the wicked comes wickedness.' But my hand shall not be against you.
1SAM|24|14|After whom has the king of Israel come out? After whom do you pursue? After a dead dog! After a flea!
1SAM|24|15|May the LORD therefore be judge and give sentence between me and you, and see to it and plead my cause and deliver me from your hand."
1SAM|24|16|As soon as David had finished speaking these words to Saul, Saul said, "Is this your voice, my son David?" And Saul lifted up his voice and wept.
1SAM|24|17|He said to David, "You are more righteous than I, for you have repaid me good, whereas I have repaid you evil.
1SAM|24|18|And you have declared this day how you have dealt well with me, in that you did not kill me when the LORD put me into your hands.
1SAM|24|19|For if a man finds his enemy, will he let him go away safe? So may the LORD reward you with good for what you have done to me this day.
1SAM|24|20|And now, behold, I know that you shall surely be king, and that the kingdom of Israel shall be established in your hand.
1SAM|24|21|Swear to me therefore by the LORD that you will not cut off my offspring after me, and that you will not destroy my name out of my father's house."
1SAM|24|22|And David swore this to Saul. Then Saul went home, but David and his men went up to the stronghold.
1SAM|25|1|Now Samuel died. And all Israel assembled and mourned for him, and they buried him in his house at Ramah. Then David rose and went down to the wilderness of Paran.
1SAM|25|2|And there was a man in Maon whose business was in Carmel. The man was very rich; he had three thousand sheep and a thousand goats. He was shearing his sheep in Carmel.
1SAM|25|3|Now the name of the man was Nabal, and the name of his wife Abigail. The woman was discerning and beautiful, but the man was harsh and badly behaved; he was a Calebite.
1SAM|25|4|David heard in the wilderness that Nabal was shearing his sheep.
1SAM|25|5|So David sent ten young men. And David said to the young men, "Go up to Carmel, and go to Nabal and greet him in my name.
1SAM|25|6|And thus you shall greet him: 'Peace be to you, and peace be to your house, and peace be to all that you have.
1SAM|25|7|I hear that you have shearers. Now your shepherds have been with us, and we did them no harm, and they missed nothing all the time they were in Carmel.
1SAM|25|8|Ask your young men, and they will tell you. Therefore let my young men find favor in your eyes, for we come on a feast day. Please give whatever you have at hand to your servants and to your son David.'"
1SAM|25|9|When David's young men came, they said all this to Nabal in the name of David, and then they waited.
1SAM|25|10|And Nabal answered David's servants, "Who is David? Who is the son of Jesse? There are many servants these days who are breaking away from their masters.
1SAM|25|11|Shall I take my bread and my water and my meat that I have killed for my shearers and give it to men who come from I do not know where?"
1SAM|25|12|So David's young men turned away and came back and told him all this.
1SAM|25|13|And David said to his men, "Every man strap on his sword!" And every man of them strapped on his sword. David also strapped on his sword. And about four hundred men went up after David, while two hundred remained with the baggage.
1SAM|25|14|But one of the young men told Abigail, Nabal's wife, "Behold, David sent messengers out of the wilderness to greet our master, and he railed at them.
1SAM|25|15|Yet the men were very good to us, and we suffered no harm, and we did not miss anything when we were in the fields, as long as we went with them.
1SAM|25|16|They were a wall to us both by night and by day, all the while we were with them keeping the sheep.
1SAM|25|17|Now therefore know this and consider what you should do, for harm is determined against our master and against all his house, and he is such a worthless man that one cannot speak to him."
1SAM|25|18|Then Abigail made haste and took two hundred loaves and two skins of wine and five sheep already prepared and five seahs of parched grain and a hundred clusters of raisins and two hundred cakes of figs, and laid them on donkeys.
1SAM|25|19|And she said to her young men, "Go on before me; behold, I come after you." But she did not tell her husband Nabal.
1SAM|25|20|And as she rode on the donkey and came down under cover of the mountain, behold, David and his men came down toward her, and she met them.
1SAM|25|21|Now David had said, "Surely in vain have I guarded all that this fellow has in the wilderness, so that nothing was missed of all that belonged to him, and he has returned me evil for good.
1SAM|25|22|God do so to the enemies of David and more also, if by morning I leave so much as one male of all who belong to him."
1SAM|25|23|When Abigail saw David, she hurried and got down from the donkey and fell before David on her face and bowed to the ground.
1SAM|25|24|She fell at his feet and said, "On me alone, my lord, be the guilt. Please let your servant speak in your ears, and hear the words of your servant.
1SAM|25|25|Let not my lord regard this worthless fellow, Nabal, for as his name is, so is he. Nabal is his name, and folly is with him. But I your servant did not see the young men of my lord, whom you sent.
1SAM|25|26|Now then, my lord, as the LORD lives, and as your soul lives, because the LORD has restrained you from bloodguilt and from saving with your own hand, now then let your enemies and those who seek to do evil to my lord be as Nabal.
1SAM|25|27|And now let this present that your servant has brought to my lord be given to the young men who follow my lord.
1SAM|25|28|Please forgive the trespass of your servant. For the LORD will certainly make my lord a sure house, because my lord is fighting the battles of the LORD, and evil shall not be found in you so long as you live.
1SAM|25|29|If men rise up to pursue you and to seek your life, the life of my lord shall be bound in the bundle of the living in the care of the LORD your God. And the lives of your enemies he shall sling out as from the hollow of a sling.
1SAM|25|30|And when the LORD has done to my lord according to all the good that he has spoken concerning you and has appointed you prince over Israel,
1SAM|25|31|my lord shall have no cause of grief or pangs of conscience for having shed blood without cause or for my lord taking vengeance himself. And when the LORD has dealt well with my lord, then remember your servant."
1SAM|25|32|And David said to Abigail, "Blessed be the LORD, the God of Israel, who sent you this day to meet me!
1SAM|25|33|Blessed be your discretion, and blessed be you, who have kept me this day from bloodguilt and from avenging myself with my own hand!
1SAM|25|34|For as surely as the LORD the God of Israel lives, who has restrained me from hurting you, unless you had hurried and come to meet me, truly by morning there had not been left to Nabal so much as one male."
1SAM|25|35|Then David received from her hand what she had brought him. And he said to her, "Go up in peace to your house. See, I have obeyed your voice, and I have granted your petition."
1SAM|25|36|And Abigail came to Nabal, and behold, he was holding a feast in his house, like the feast of a king. And Nabal's heart was merry within him, for he was very drunk. So she told him nothing at all until the morning light.
1SAM|25|37|In the morning, when the wine had gone out of Nabal, his wife told him these things, and his heart died within him, and he became as a stone.
1SAM|25|38|And about ten days later the LORD struck Nabal, and he died.
1SAM|25|39|When David heard that Nabal was dead, he said, "Blessed be the LORD who has avenged the insult I received at the hand of Nabal, and has kept back his servant from wrongdoing. The LORD has returned the evil of Nabal on his own head." Then David sent and spoke to Abigail, to take her as his wife.
1SAM|25|40|When the servants of David came to Abigail at Carmel, they said to her, "David has sent us to you to take you to him as his wife."
1SAM|25|41|And she rose and bowed with her face to the ground and said, "Behold, your handmaid is a servant to wash the feet of the servants of my lord."
1SAM|25|42|And Abigail hurried and rose and mounted a donkey, and her five young women attended her. She followed the messengers of David and became his wife.
1SAM|25|43|David also took Ahinoam of Jezreel, and both of them became his wives.
1SAM|25|44|Saul had given Michal his daughter, David's wife, to Palti the son of Laish, who was of Gallim.
1SAM|26|1|Then the Ziphites came to Saul at Gibeah, saying, "Is not David hiding himself on the hill of Hachilah, which is on the east of Jeshimon?"
1SAM|26|2|So Saul arose and went down to the wilderness of Ziph with three thousand chosen men of Israel to seek David in the wilderness of Ziph.
1SAM|26|3|And Saul encamped on the hill of Hachilah, which is beside the road on the east of Jeshimon. But David remained in the wilderness. When he saw that Saul came after him into the wilderness,
1SAM|26|4|David sent out spies and learned that Saul had come.
1SAM|26|5|Then David rose and came to the place where Saul had encamped. And David saw the place where Saul lay, with Abner the son of Ner, the commander of his army. Saul was lying within the encampment, while the army was encamped around him.
1SAM|26|6|Then David said to Ahimelech the Hittite, and to Joab's brother Abishai the son of Zeruiah, "Who will go down with me into the camp to Saul?" And Abishai said, "I will go down with you."
1SAM|26|7|So David and Abishai went to the army by night. And there lay Saul sleeping within the encampment, with his spear stuck in the ground at his head, and Abner and the army lay around him.
1SAM|26|8|Then said Abishai to David, "God has given your enemy into your hand this day. Now please let me pin him to the earth with one stroke of the spear, and I will not strike him twice."
1SAM|26|9|But David said to Abishai, "Do not destroy him, for who can put out his hand against the LORD's anointed and be guiltless?"
1SAM|26|10|And David said, "As the LORD lives, the LORD will strike him, or his day will come to die, or he will go down into battle and perish.
1SAM|26|11|The LORD forbid that I should put out my hand against the LORD's anointed. But take now the spear that is at his head and the jar of water, and let us go."
1SAM|26|12|So David took the spear and the jar of water from Saul's head, and they went away. No man saw it or knew it, nor did any awake, for they were all asleep, because a deep sleep from the LORD had fallen upon them.
1SAM|26|13|Then David went over to the other side and stood far off on the top of the hill, with a great space between them.
1SAM|26|14|And David called to the army, and to Abner the son of Ner, saying, "Will you not answer, Abner?" Then Abner answered, "Who are you who calls to the king?"
1SAM|26|15|And David said to Abner, "Are you not a man? Who is like you in Israel? Why then have you not kept watch over your lord the king? For one of the people came in to destroy the king your lord.
1SAM|26|16|This thing that you have done is not good. As the LORD lives, you deserve to die, because you have not kept watch over your lord, the LORD's anointed. And now see where the king's spear is and the jar of water that was at his head."
1SAM|26|17|Saul recognized David's voice and said, "Is this your voice, my son David?" And David said, "It is my voice, my lord, O king."
1SAM|26|18|And he said, "Why does my lord pursue after his servant? For what have I done? What evil is on my hands?
1SAM|26|19|Now therefore let my lord the king hear the words of his servant. If it is the LORD who has stirred you up against me, may he accept an offering, but if it is men, may they be cursed before the LORD, for they have driven me out this day that I should have no share in the heritage of the LORD, saying, 'Go, serve other gods.'
1SAM|26|20|Now therefore, let not my blood fall to the earth away from the presence of the LORD, for the king of Israel has come out to seek a single flea like one who hunts a partridge in the mountains."
1SAM|26|21|Then Saul said, "I have sinned. Return, my son David, for I will no more do you harm, because my life was precious in your eyes this day. Behold, I have acted foolishly, and have made a great mistake."
1SAM|26|22|And David answered and said, "Here is the spear, O king! Let one of the young men come over and take it.
1SAM|26|23|The LORD rewards every man for his righteousness and his faithfulness, for the LORD gave you into my hand today, and I would not put out my hand against the LORD's anointed.
1SAM|26|24|Behold, as your life was precious this day in my sight, so may my life be precious in the sight of the LORD, and may he deliver me out of all tribulation."
1SAM|26|25|Then Saul said to David, "Blessed be you, my son David! You will do many things and will succeed in them." So David went his way, and Saul returned to his place.
1SAM|27|1|Then David said in his heart, "Now I shall perish one day by the hand of Saul. There is nothing better for me than that I should escape to the land of the Philistines. Then Saul will despair of seeking me any longer within the borders of Israel, and I shall escape out of his hand."
1SAM|27|2|So David arose and went over, he and the six hundred men who were with him, to Achish the son of Maoch, king of Gath.
1SAM|27|3|And David lived with Achish at Gath, he and his men, every man with his household, and David with his two wives, Ahinoam of Jezreel, and Abigail of Carmel, Nabal's widow.
1SAM|27|4|And when it was told Saul that David had fled to Gath, he no longer sought him.
1SAM|27|5|Then David said to Achish, "If I have found favor in your eyes, let a place be given me in one of the country towns, that I may dwell there. For why should your servant dwell in the royal city with you?"
1SAM|27|6|So that day Achish gave him Ziklag. Therefore Ziklag has belonged to the kings of Judah to this day.
1SAM|27|7|And the number of the days that David lived in the country of the Philistines was a year and four months.
1SAM|27|8|Now David and his men went up and made raids against the Geshurites, the Girzites, and the Amalekites, for these were the inhabitants of the land from of old, as far as Shur, to the land of Egypt.
1SAM|27|9|And David would strike the land and would leave neither man nor woman alive, but would take away the sheep, the oxen, the donkeys, the camels, and the garments, and come back to Achish.
1SAM|27|10|When Achish asked, "Where have you made a raid today?" David would say, "Against the Negeb of Judah," or, "Against the Negeb of the Jerahmeelites," or, "Against the Negeb of the Kenites."
1SAM|27|11|And David would leave neither man nor woman alive to bring news to Gath, thinking, "Lest they should tell about us and say, 'So David has done.'"Such was his custom all the while he lived in the country of the Philistines.
1SAM|27|12|And Achish trusted David, thinking, "He has made himself an utter stench to his people Israel; therefore he shall always be my servant."
1SAM|28|1|In those days the Philistines gathered their forces for war, to fight against Israel. And Achish said to David, "Understand that you and your men are to go out with me in the army."
1SAM|28|2|David said to Achish, "Very well, you shall know what your servant can do." And Achish said to David, "Very well, I will make you my bodyguard for life."
1SAM|28|3|Now Samuel had died, and all Israel had mourned for him and buried him in Ramah, his own city. And Saul had put the mediums and the necromancers out of the land.
1SAM|28|4|The Philistines assembled and came and encamped at Shunem. And Saul gathered all Israel, and they encamped at Gilboa.
1SAM|28|5|When Saul saw the army of the Philistines, he was afraid, and his heart trembled greatly.
1SAM|28|6|And when Saul inquired of the LORD, the LORD did not answer him, either by dreams, or by Urim, or by prophets.
1SAM|28|7|Then Saul said to his servants, "Seek out for me a woman who is a medium, that I may go to her and inquire of her." And his servants said to him, "Behold, there is a medium at En-dor."
1SAM|28|8|So Saul disguised himself and put on other garments and went, he and two men with him. And they came to the woman by night. And he said, "Divine for me by a spirit and bring up for me whomever I shall name to you."
1SAM|28|9|The woman said to him, "Surely you know what Saul has done, how he has cut off the mediums and the necromancers from the land. Why then are you laying a trap for my life to bring about my death?"
1SAM|28|10|But Saul swore to her by the LORD, "As the LORD lives, no punishment shall come upon you for this thing."
1SAM|28|11|Then the woman said, "Whom shall I bring up for you?" He said, "Bring up Samuel for me."
1SAM|28|12|When the woman saw Samuel, she cried out with a loud voice. And the woman said to Saul, "Why have you deceived me? You are Saul."
1SAM|28|13|The king said to her, "Do not be afraid. What do you see?" And the woman said to Saul, "I see a god coming up out of the earth."
1SAM|28|14|He said to her, "What is his appearance?" And she said, "An old man is coming up, and he is wrapped in a robe." And Saul knew that it was Samuel, and he bowed with his face to the ground and paid homage.
1SAM|28|15|Then Samuel said to Saul, "Why have you disturbed me by bringing me up?" Saul answered, "I am in great distress, for the Philistines are warring against me, and God has turned away from me and answers me no more, either by prophets or by dreams. Therefore I have summoned you to tell me what I shall do."
1SAM|28|16|And Samuel said, "Why then do you ask me, since the LORD has turned from you and become your enemy?
1SAM|28|17|The LORD has done to you as he spoke by me, for the LORD has torn the kingdom out of your hand and given it to your neighbor, David.
1SAM|28|18|Because you did not obey the voice of the LORD and did not carry out his fierce wrath against Amalek, therefore the LORD has done this thing to you this day.
1SAM|28|19|Moreover, the LORD will give Israel also with you into the hand of the Philistines, and tomorrow you and your sons shall be with me. The LORD will give the army of Israel also into the hand of the Philistines."
1SAM|28|20|Then Saul fell at once full length on the ground, filled with fear because of the words of Samuel. And there was no strength in him, for he had eaten nothing all day and all night.
1SAM|28|21|And the woman came to Saul, and when she saw that he was terrified, she said to him, "Behold, your servant has obeyed you. I have taken my life in my hand and have listened to what you have said to me.
1SAM|28|22|Now therefore, you also obey your servant. Let me set a morsel of bread before you; and eat, that you may have strength when you go on your way."
1SAM|28|23|He refused and said, "I will not eat." But his servants, together with the woman, urged him, and he listened to their words. So he arose from the earth and sat on the bed.
1SAM|28|24|Now the woman had a fattened calf in the house, and she quickly killed it, and she took flour and kneaded it and baked unleavened bread of it,
1SAM|28|25|and she put it before Saul and his servants, and they ate. Then they rose and went away that night.
1SAM|29|1|Now the Philistines had gathered all their forces at Aphek. And the Israelites were encamped by the spring that is in Jezreel.
1SAM|29|2|As the lords of the Philistines were passing on by hundreds and by thousands, and David and his men were passing on in the rear with Achish,
1SAM|29|3|the commanders of the Philistines said, "What are these Hebrews doing here?" And Achish said to the commanders of the Philistines, "Is this not David, the servant of Saul, king of Israel, who has been with me now for days and years, and since he deserted to me I have found no fault in him to this day."
1SAM|29|4|But the commanders of the Philistines were angry with him. And the commanders of the Philistines said to him, "Send the man back, that he may return to the place to which you have assigned him. He shall not go down with us to battle, lest in the battle he become an adversary to us. For how could this fellow reconcile himself to his lord? Would it not be with the heads of the men here?
1SAM|29|5|Is not this David, of whom they sing to one another in dances, 'Saul has struck down his thousands, and David his ten thousands'?"
1SAM|29|6|Then Achish called David and said to him, "As the LORD lives, you have been honest, and to me it seems right that you should march out and in with me in the campaign. For I have found nothing wrong in you from the day of your coming to me to this day. Nevertheless, the lords do not approve of you.
1SAM|29|7|So go back now; and go peaceably, that you may not displease the lords of the Philistines."
1SAM|29|8|And David said to Achish, "But what have I done? What have you found in your servant from the day I entered your service until now, that I may not go and fight against the enemies of my lord the king?"
1SAM|29|9|And Achish answered David and said, "I know that you are as blameless in my sight as an angel of God. Nevertheless, the commanders of the Philistines have said, 'He shall not go up with us to the battle.'
1SAM|29|10|Now then rise early in the morning with the servants of your lord who came with you, and start early in the morning, and depart as soon as you have light."
1SAM|29|11|So David set out with his men early in the morning to return to the land of the Philistines. But the Philistines went up to Jezreel.
1SAM|30|1|Now when David and his men came to Ziklag on the third day, the Amalekites had made a raid against the Negeb and against Ziklag. They had overcome Ziklag and burned it with fire
1SAM|30|2|and taken captive the women and all who were in it, both small and great. They killed no one, but carried them off and went their way.
1SAM|30|3|And when David and his men came to the city, they found it burned with fire, and their wives and sons and daughters taken captive.
1SAM|30|4|Then David and the people who were with him raised their voices and wept until they had no more strength to weep.
1SAM|30|5|David's two wives also had been taken captive, Ahinoam of Jezreel and Abigail the widow of Nabal of Carmel.
1SAM|30|6|And David was greatly distressed, for the people spoke of stoning him, because all the people were bitter in soul, each for his sons and daughters. But David strengthened himself in the LORD his God.
1SAM|30|7|And David said to Abiathar the priest, the son of Ahimelech, "Bring me the ephod." So Abiathar brought the ephod to David.
1SAM|30|8|And David inquired of the LORD, "Shall I pursue after this band? Shall I overtake them?" He answered him, "Pursue, for you shall surely overtake and shall surely rescue."
1SAM|30|9|So David set out, and the six hundred men who were with him, and they came to the brook Besor, where those who were left behind stayed.
1SAM|30|10|But David pursued, he and four hundred men. Two hundred stayed behind, who were too exhausted to cross the brook Besor.
1SAM|30|11|They found an Egyptian in the open country and brought him to David. And they gave him bread and he ate. They gave him water to drink,
1SAM|30|12|and they gave him a piece of a cake of figs and two clusters of raisins. And when he had eaten, his spirit revived, for he had not eaten bread or drunk water for three days and three nights.
1SAM|30|13|And David said to him, "To whom do you belong? And where are you from?" He said, "I am a young man of Egypt, servant to an Amalekite, and my master left me behind because I fell sick three days ago.
1SAM|30|14|We had made a raid against the Negeb of the Cherethites and against that which belongs to Judah and against the Negeb of Caleb, and we burned Ziklag with fire."
1SAM|30|15|And David said to him, "Will you take me down to this band?" And he said, "Swear to me by God that you will not kill me or deliver me into the hands of my master, and I will take you down to this band."
1SAM|30|16|And when he had taken him down, behold, they were spread abroad over all the land, eating and drinking and dancing, because of all the great spoil they had taken from the land of the Philistines and from the land of Judah.
1SAM|30|17|And David struck them down from twilight until the evening of the next day, and not a man of them escaped, except four hundred young men, who mounted camels and fled.
1SAM|30|18|David recovered all that the Amalekites had taken, and David rescued his two wives.
1SAM|30|19|Nothing was missing, whether small or great, sons or daughters, spoil or anything that had been taken. David brought back all.
1SAM|30|20|David also captured all the flocks and herds, and the people drove the livestock before him, and said, "This is David's spoil."
1SAM|30|21|Then David came to the two hundred men who had been too exhausted to follow David, and who had been left at the brook Besor. And they went out to meet David and to meet the people who were with him. And when David came near to the people he greeted them.
1SAM|30|22|Then all the wicked and worthless fellows among the men who had gone with David said, "Because they did not go with us, we will not give them any of the spoil that we have recovered, except that each man may lead away his wife and children, and depart."
1SAM|30|23|But David said, "You shall not do so, my brothers, with what the LORD has given us. He has preserved us and given into our hand the band that came against us.
1SAM|30|24|Who would listen to you in this matter? For as his share is who goes down into the battle, so shall his share be who stays by the baggage. They shall share alike."
1SAM|30|25|And he made it a statute and a rule for Israel from that day forward to this day.
1SAM|30|26|When David came to Ziklag, he sent part of the spoil to his friends, the elders of Judah, saying, "Here is a present for you from the spoil of the enemies of the LORD."
1SAM|30|27|It was for those in Bethel, in Ramoth of the Negeb, in Jattir,
1SAM|30|28|in Aroer, in Siphmoth, in Eshtemoa,
1SAM|30|29|in Racal, in the cities of the Jerahmeelites, in the cities of the Kenites,
1SAM|30|30|in Hormah, in Bor-ashan, in Athach,
1SAM|30|31|in Hebron, for all the places where David and his men had roamed.
1SAM|31|1|Now the Philistines fought against Israel, and the men of Israel fled before the Philistines and fell slain on Mount Gilboa.
1SAM|31|2|And the Philistines overtook Saul and his sons, and the Philistines struck down Jonathan and Abinadab and Malchi-shua, the sons of Saul.
1SAM|31|3|The battle pressed hard against Saul, and the archers found him, and he was badly wounded by the archers.
1SAM|31|4|Then Saul said to his armor-bearer, "Draw your sword, and thrust me through with it, lest these uncircumcised come and thrust me through, and mistreat me." But his armor-bearer would not, for he feared greatly. Therefore Saul took his own sword and fell upon it.
1SAM|31|5|And when his armor-bearer saw that Saul was dead, he also fell upon his sword and died with him.
1SAM|31|6|Thus Saul died, and his three sons, and his armor-bearer, and all his men, on the same day together.
1SAM|31|7|And when the men of Israel who were on the other side of the valley and those beyond the Jordan saw that the men of Israel had fled and that Saul and his sons were dead, they abandoned their cities and fled. And the Philistines came and lived in them.
1SAM|31|8|The next day, when the Philistines came to strip the slain, they found Saul and his three sons fallen on Mount Gilboa.
1SAM|31|9|So they cut off his head and stripped off his armor and sent messengers throughout the land of the Philistines, to carry the good news to the house of their idols and to the people.
1SAM|31|10|They put his armor in the temple of Ashtaroth, and they fastened his body to the wall of Beth-shan.
1SAM|31|11|But when the inhabitants of Jabesh-gilead heard what the Philistines had done to Saul,
1SAM|31|12|all the valiant men arose and went all night and took the body of Saul and the bodies of his sons from the wall of Beth-shan, and they came to Jabesh and burned them there.
1SAM|31|13|And they took their bones and buried them under the tamarisk tree in Jabesh and fasted seven days.
