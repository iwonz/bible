1COR|1|1|Paulus, vocatus apostolus Christi Iesu per voluntatem Dei, et Sosthenes frater
1COR|1|2|ecclesiae Dei, quae est Corinthi, sanctificatis in Christo Iesu, vocatis sanctis cum omnibus, qui invocant nomen Domini nostri Iesu Christi in omni loco ipsorum et nostro:
1COR|1|3|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo.
1COR|1|4|Gratias ago Deo meo semper pro vobis in gratia Dei, quae data est vobis in Christo Iesu,
1COR|1|5|quia in omnibus divites facti estis in illo, in omni verbo et in omni scientia,
1COR|1|6|sicut testimonium Christi confirmatum est in vobis,
1COR|1|7|ita ut nihil vobis desit in ulla donatione, exspectantibus revelationem Domini nostri Iesu Christi;
1COR|1|8|qui et confirmabit vos usque ad finem sine crimine in die Domini nostri Iesu Christi.
1COR|1|9|Fidelis Deus, per quem vocati estis in communionem Filii eius Iesu Christi Domini nostri.
1COR|1|10|Obsecro autem vos, fratres, per nomen Domini nostri Iesu Christi, ut idipsum dicatis omnes, et non sint in vobis schismata, sitis autem perfecti in eodem sensu et in eadem sententia.
1COR|1|11|Significatum est enim mihi de vobis, fratres mei, ab his, qui sunt Chloes, quia contentiones inter vos sunt.
1COR|1|12|Hoc autem dico, quod unusquisque vestrum dicit: " Ego quidem sum Pauli, " Ego autem Apollo ", " Ego vero Cephae ", " Ego autem Christi ".
1COR|1|13|Divisus est Christus? Numquid Paulus crucifixus est pro vobis, aut in nomine Pauli baptizati estis?
1COR|1|14|Gratias ago Deo quod neminem vestrum baptizavi, nisi Crispum et Gaium,
1COR|1|15|ne quis dicat quod in nomine meo baptizati sitis.
1COR|1|16|Baptizavi autem et Stephanae domum; ceterum nescio si quem alium baptizaverim.
1COR|1|17|Non enim misit me Christus baptizare, sed evangelizare; non in sapientia verbi, ut non evacuetur crux Christi.
1COR|1|18|Verbum enim crucis pereuntibus quidem stultitia est; his autem, qui salvi fiunt, id est nobis, virtus Dei est.
1COR|1|19|Scriptum est enim: Perdam sapientiam sapientiumet prudentiam prudentium reprobabo ".
1COR|1|20|Ubi sapiens? Ubi scriba? Ubi conquisitor huius saeculi? Nonne stultam fecit Deus sapientiam huius mundi?
1COR|1|21|Nam quia in Dei sapientia non cognovit mundus per sapientiam Deum, placuit Deo per stultitiam praedicationis salvos facere credentes.
1COR|1|22|Quoniam et Iudaei signa petunt, et Graeci sapientiam quaerunt,
1COR|1|23|nos autem praedicamus Christum crucifixum, Iudaeis quidem scandalum, gentibus autem stultitiam;
1COR|1|24|ipsis autem vocatis, Iudaeis atque Graecis, Christum Dei virtutem et Dei sapientiam;
1COR|1|25|quia quod stultum est Dei, sapientius est hominibus, et, quod infirmum est Dei, fortius est hominibus.
1COR|1|26|Videte enim vocationem vestram, fratres; quia non multi sapientes secundum carnem, non multi potentes, non multi nobiles;
1COR|1|27|sed, quae stulta sunt mundi, elegit Deus, ut confundat sapientes, et infirma mundi elegit Deus, ut confundat fortia,
1COR|1|28|et ignobilia mundi et contemptibilia elegit Deus, quae non sunt, ut ea, quae sunt, destrueret,
1COR|1|29|ut non glorietur omnis caro in conspectu Dei.
1COR|1|30|Ex ipso autem vos estis in Christo Iesu, qui factus est sapientia nobis a Deo et iustitia et sanctificatio et redemptio,
1COR|1|31|ut quemadmodum scriptum est: Qui gloriatur, in Domino glorietur ".
1COR|2|1|Et ego, cum venissem ad vos, fratres, veni non per sublimita tem sermonis aut sapientiae annuntians vobis mysterium Dei.
1COR|2|2|Non enim iudicavi scire me aliquid inter vos nisi Iesum Christum et hunc crucifixum.
1COR|2|3|Et ego in infirmitate et timore et tremore multo fui apud vos,
1COR|2|4|et sermo meus et praedicatio mea non in persuasibilibus sapientiae verbis sed in ostensione Spiritus et virtutis,
1COR|2|5|ut fides vestra non sit in sapientia hominum sed in virtute Dei.
1COR|2|6|Sapientiam autem loquimur inter perfectos, sapientiam vero non huius saeculi neque principum huius saeculi, qui destruuntur,
1COR|2|7|sed loquimur Dei sapientiam in mysterio, quae abscondita est, quam praedestinavit Deus ante saecula in gloriam nostram,
1COR|2|8|quam nemo principum huius saeculi cognovit; si enim cognovissent, numquam Dominum gloriae crucifixissent.
1COR|2|9|Sed sicut scriptum est: " Quod oculus non vidit, nec auris audivit, nec in cor hominis ascendit, quae praeparavit Deus his, qui diligunt illum ".
1COR|2|10|Nobis autem revelavit Deus per Spiritum; Spiritus enim omnia scrutatur, etiam profunda Dei.
1COR|2|11|Quis enim scit hominum, quae sint hominis, nisi spiritus hominis, qui in ipso est? Ita et, quae Dei sunt, nemo cognovit nisi Spiritus Dei.
1COR|2|12|Nos autem non spiritum mundi accepimus, sed Spiritum, qui ex Deo est, ut sciamus, quae a Deo donata sunt nobis;
1COR|2|13|quae et loquimur non in doctis humanae sapientiae sed in doctis Spiritus verbis, spiritalibus spiritalia comparantes.
1COR|2|14|Animalis autem homo non percipit, quae sunt Spiritus Dei, stultitia enim sunt illi, et non potest intellegere, quia spiritaliter examinantur;
1COR|2|15|spiritalis autem iudicat omnia, et ipse a nemine iudicatur.
1COR|2|16|Quis enim cognovit sensum Domini,qui instruat eum?Nos autem sensum Christi habemus.
1COR|3|1|Et ego, fratres, non potui vobis loqui quasi spiritalibus sed qua si carnalibus, tamquam parvulis in Christo.
1COR|3|2|Lac vobis potum dedi, non escam, nondum enim poteratis. Sed ne nunc quidem potestis,
1COR|3|3|adhuc enim estis carnales. Cum enim sit inter vos zelus et contentio, nonne carnales estis et secundum hominem ambulatis?
1COR|3|4|Cum enim quis dicit: " Ego quidem sum Pauli ", alius autem: " Ego Apollo, nonne homines estis?
1COR|3|5|Quid igitur est Apollo? Quid vero Paulus? Ministri, per quos credidistis, et unicuique sicut Dominus dedit.
1COR|3|6|Ego plantavi, Apollo rigavit, sed Deus incrementum dedit;
1COR|3|7|itaque neque qui plantat, est aliquid, neque qui rigat, sed qui incrementum dat, Deus.
1COR|3|8|Qui plantat autem et qui rigat unum sunt; unusquisque autem propriam mercedem accipiet secundum suum laborem.
1COR|3|9|Dei enim sumus adiutores: Dei agri cultura estis, Dei aedificatio estis.
1COR|3|10|Secundum gratiam Dei, quae data est mihi, ut sapiens architectus fundamentum posui; alius autem superaedificat. Unusquisque autem videat quomodo superaedificet;
1COR|3|11|fundamentum enim aliud nemo potest ponere praeter id, quod positum est, qui est Iesus Christus.
1COR|3|12|Si quis autem superaedificat supra fundamentum aurum, argentum, lapides pretiosos, ligna, fenum, stipulam,
1COR|3|13|uniuscuiusque opus manifestum erit; dies enim declarabit: quia in igne revelatur, et uniuscuiusque opus quale sit ignis probabit.
1COR|3|14|Si cuius opus manserit, quod superaedificavit, mercedem accipiet;
1COR|3|15|si cuius opus arserit, detrimentum patietur, ipse autem salvus erit, sic tamen quasi per ignem.
1COR|3|16|Nescitis quia templum Dei estis, et Spiritus Dei habitat in vobis?
1COR|3|17|Si quis autem templum Dei everterit, evertet illum Deus; templum enim Dei sanctum est, quod estis vos.
1COR|3|18|Nemo se seducat; si quis videtur sapiens esse inter vos in hoc saeculo, stultus fiat, ut sit sapiens.
1COR|3|19|Sapientia enim huius mundi stultitia est apud Deum. Scriptum est enim: Qui apprehendit sapientes in astutia eorum ";
1COR|3|20|et iterum: Dominus novit cogitationes sapientium,quoniam vanae sunt ".
1COR|3|21|Itaque nemo glorietur in hominibus. Omnia enim vestra sunt,
1COR|3|22|sive Paulus sive Apollo sive Cephas sive mundus sive vita sive mors sive praesentia sive futura, omnia enim vestra sunt,
1COR|3|23|vos autem Christi, Christus autem Dei.
1COR|4|1|Sic nos existimet homo ut mi nistros Christi et dispensatores mysteriorum Dei.
1COR|4|2|Hic iam quaeritur inter dispensatores, ut fidelis quis inveniatur.
1COR|4|3|Mihi autem pro minimo est, ut a vobis iudicer aut ab humano die. Sed neque meipsum iudico;
1COR|4|4|nihil enim mihi conscius sum, sed non in hoc iustificatus sum. Qui autem iudicat me, Dominus est!
1COR|4|5|Itaque nolite ante tempus quidquam iudicare, quoadusque veniat Dominus, qui et illuminabit abscondita tenebrarum et manifestabit consilia cordium; et tunc laus erit unicuique a Deo.
1COR|4|6|Haec autem, fratres, transfiguravi in me et Apollo propter vos, ut in nobis discatis illud: " Ne supra quae scripta sunt ", ne unus pro alio inflemini adversus alterum.
1COR|4|7|Quis enim te discernit? Quid autem habes, quod non accepisti? Si autem accepisti, quid gloriaris, quasi non acceperis?
1COR|4|8|Iam saturati estis, iam divites facti estis. Sine nobis regnastis; et utinam regnaretis, ut et nos vobiscum regnaremus.
1COR|4|9|Puto enim, Deus nos apostolos novissimos ostendit tamquam morti destinatos, quia spectaculum facti sumus mundo et angelis et hominibus.
1COR|4|10|Nos stulti propter Christum, vos autem prudentes in Christo; nos infirmi, vos autem fortes; vos gloriosi, nos autem ignobiles.
1COR|4|11|Usque in hanc horam et esurimus et sitimus et nudi sumus et colaphis caedimur et instabiles sumus
1COR|4|12|et laboramus operantes manibus nostris; maledicti benedicimus, persecutionem passi sustinemus,
1COR|4|13|blasphemati obsecramus; tamquam purgamenta mundi facti sumus, omnium peripsema, usque adhuc.
1COR|4|14|Non ut confundam vos, haec scribo, sed ut quasi filios meos carissimos moneam;
1COR|4|15|nam si decem milia paedagogorum habeatis in Christo, sed non multos patres, nam in Christo Iesu per evangelium ego vos genui.
1COR|4|16|Rogo ergo vos: imitatorcs mei estote!
1COR|4|17|Ideo misi ad vos Timotheum, qui est filius meus carissimus et fidelis in Domino, qui vos commonefaciat vias meas, quae sunt in Christo, sicut ubique in omni ecclesia doceo.
1COR|4|18|Tamquam non venturus sim ad vos, sic inflati sunt quidam;
1COR|4|19|veniam autem cito ad vos, si Dominus voluerit, et cognoscam non sermonem eorum, qui inflati sunt, sed virtutem;
1COR|4|20|non enim in sermone est regnum Dei sed in virtute.
1COR|4|21|Quid vultis? In virga veniam ad vos an in caritate et spiritu mansuetudinis?
1COR|5|1|Omnino auditur inter vos for nicatio, et talis fornicatio qualis nec inter gentes, ita ut uxorem patris aliquis habeat.
1COR|5|2|Et vos inflati estis et non magis luctum habuistis, ut tollatur de medio vestrum, qui hoc opus fecit?
1COR|5|3|Ego quidem absens corpore, praesens autem spiritu, iam iudicavi ut praesens eum, qui sic operatus est,
1COR|5|4|in nomine Domini nostri Iesu, congregatis vobis et meo spiritu cum virtute Domini nostri Iesu,
1COR|5|5|tradere huiusmodi Satanae in interitum carnis, ut spiritus salvus sit in die Domini.
1COR|5|6|Non bona gloriatio vestra. Nescitis quia modicum fermentum totam massam corrumpit?
1COR|5|7|Expurgate vetus fermentum, ut sitis nova consparsio, sicut estis azymi. Etenim Pascha nostrum immolatus est Christus!
1COR|5|8|Itaque festa celebremus, non in fermento veteri neque in fermento malitiae et nequitiae, sed in azymis sinceritatis et veritatis.
1COR|5|9|Scripsi vobis in epistula: Ne commisceamini fornicariis.
1COR|5|10|Non utique fornicariis huius mundi aut avaris aut rapacibus aut idolis servientibus, alioquin debueratis de hoc mundo exisse!
1COR|5|11|Nunc autem scripsi vobis non commisceri, si is, qui frater nominatur, est fornicator aut avarus aut idolis serviens aut maledicus aut ebriosus aut rapax; cum eiusmodi nec cibum sumere.
1COR|5|12|Quid enim mihi de his, qui foris sunt, iudicare? Nonne de his, qui intus sunt, vos iudicatis?
1COR|5|13|Nam eos, qui foris sunt, Deus iudicabit. Auferte malum ex vobis ipsis!
1COR|6|1|Audet aliquis vestrum habens negotium adversus alterum iu dicari apud iniquos et non apud sanctos?
1COR|6|2|An nescitis quoniam sancti de mundo iudicabunt? Et si in vobis iudicabitur mundus, indigni estis minimis iudiciis?
1COR|6|3|Nescitis quoniam angelos iudicabimus, quanto magis saecularia?
1COR|6|4|Saecularia igitur iudicia si habueritis, contemptibiles, qui sunt in ecclesia, illos constituite ad iudicandum?
1COR|6|5|Ad verecundiam vestram dico! Sic non est inter vos sapiens quisquam, qui possit iudicare inter fratrem suum?
1COR|6|6|Sed frater cum fratre iudicio contendit, et hoc apud infideles?
1COR|6|7|Iam quidem omnino defectio est vobis, quod iudicia habetis inter vosmetipsos! Quare non magis iniuriam accipitis, quare non magis fraudem patimini?
1COR|6|8|Sed vos iniuriam facitis et fraudatis, et hoc fratribus!
1COR|6|9|An nescitis quia iniqui regnum Dei non possidebunt? Nolite errare: neque fornicarii neque idolis servientes neque adulteri neque molles neque masculorum concubitores
1COR|6|10|neque fures neque avari, non ebriosi, non maledici, non rapaces regnum Dei possidebunt.
1COR|6|11|Et haec quidam fuistis. Sed abluti estis, sed sanctificati estis, sed iustificati estis in nomine Domini Iesu Christi et in Spiritu Dei nostri!
1COR|6|12|" Omnia mihi licent! ". Sed non omnia expediunt. " Omnia mihi licent!. Sed ego sub nullius redigar potestate.
1COR|6|13|" Esca ventri, et venter escis! ". Deus autem et hunc et has destruet. Corpus autem non fornicationi sed Domino, et Dominus corpori;
1COR|6|14|Deus vero et Dominum suscitavit et nos suscitabit per virtutem suam.
1COR|6|15|Nescitis quoniam corpora vestra membra Christi sunt? Tollens ergo membra Christi faciam membra meretricis? Absit!
1COR|6|16|An nescitis quoniam, qui adhaeret meretrici, unum corpus est? " Erunt enim, inquit, duo in carne una ".
1COR|6|17|Qui autem adhaeret Domino, unus Spiritus est.
1COR|6|18|Fugite fornicationem! Omne peccatum, quodcumque fecerit homo, extra corpus est; qui autem fornicatur, in corpus suum peccat.
1COR|6|19|An nescitis quoniam corpus vestrum templum est Spiritus Sancti, qui in vobis est, quem habetis a Deo, et non estis vestri?
1COR|6|20|Empti enim estis pretio! Glorificate ergo Deum in corpore vestro.
1COR|7|1|De quibus autem scripsistis, bo num est homini mulierem non non tangere;
1COR|7|2|propter fornicationes autem unusquisque suam uxorem habeat, et unaquaeque suum virum habeat.
1COR|7|3|Uxori vir debitum reddat; similiter autem et uxor viro.
1COR|7|4|Mulier sui corporis potestatem non habet sed vir; similiter autem et vir sui corporis potestatem non habet sed mulier.
1COR|7|5|Nolite fraudare invicem, nisi forte ex consensu ad tempus, ut vacetis orationi et iterum sitis in idipsum, ne tentet vos Satanas propter incontinentiam vestram.
1COR|7|6|Hoc autem dico secundum indulgentiam, non secundum imperium.
1COR|7|7|Volo autem omnes homines esse sicut meipsum; sed unusquisque proprium habet donum ex Deo: alius quidem sic, alius vero sic.
1COR|7|8|Dico autem innuptis et viduis: Bonum est illis si sic maneant, sicut et ego;
1COR|7|9|quod si non se continent, nubant. Melius est enim nubere quam uri.
1COR|7|10|His autem, qui matrimonio iuncti sunt, praecipio, non ego sed Dominus, uxorem a viro non discedere
1COR|7|11|- quod si discesserit, maneat innupta aut viro suo reconcilietur - et virum uxorem non dimittere.
1COR|7|12|Ceteris autem ego dico, non Dominus: Si quis frater uxorem habet infidelem, et haec consentit habitare cum illo, non dimittat illam;
1COR|7|13|et si qua mulier habet virum infidelem, et hic consentit habitare cum illa, non dimittat virum.
1COR|7|14|Sanctificatus est enim vir infidelis in muliere, et sanctificata est mulier infidelis in fratre. Alioquin filii vestri immundi essent; nunc autem sancti sunt.
1COR|7|15|Quod si infidelis discedit, discedat. Non est enim servituti subiectus frater aut soror in eiusmodi; in pace autem vocavit nos Deus.
1COR|7|16|Quid enim scis, mulier, si virum salvum facies? Aut quid scis, vir, si mulierem salvam facies?
1COR|7|17|Nisi unicuique, sicut divisit Dominus, unumquemque, sicut vocavit Deus, ita ambulet; et sic in omnibus ecclesiis doceo.
1COR|7|18|Circumcisus aliquis vocatus est? Non adducat praeputium! In praeputio aliquis vocatus est? Non circumcidatur!
1COR|7|19|Circumcisio nihil est, et praeputium nihil est, sed observatio mandatorum Dei.
1COR|7|20|Unusquisque, in qua vocatione vocatus est, in ea permaneat.
1COR|7|21|Servus vocatus es? Non sit tibi curae; sed et si potes liber fieri, magis utere!
1COR|7|22|Qui enim in Domino vocatus est servus, libertus est Domini; similiter, qui liber vocatus est, servus est Christi!
1COR|7|23|Pretio empti estis! Nolite fieri servi hominum.
1COR|7|24|Unusquisque, in quo vocatus est, fratres, in hoc maneat apud Deum.
1COR|7|25|De virginibus autem praeceptum Domini non habeo; consilium autem do, tamquam misericordiam consecutus a Domino, ut sim fidelis.
1COR|7|26|Existimo ergo hoc bonum esse propter instantem necessitatem, quoniam bonum est homini sic esse.
1COR|7|27|Alligatus es uxori? Noli quaerere solutionem. Solutus es ab uxore? Noli quaerere uxorem.
1COR|7|28|Si autem acceperis uxorem, non peccasti; et si nupserit virgo, non peccavit. Tribulationem tamen carnis habebunt huiusmodi, ego autem vobis parco.
1COR|7|29|Hoc itaque dico, fratres, tempus breviatum est; reliquum est, ut et qui habent uxores, tamquam non habentes sint,
1COR|7|30|et qui flent, tamquam non flentes, et qui gaudent, tamquam non gaudentes, et qui emunt, tamquam non possidentes,
1COR|7|31|et qui utuntur hoc mundo, tamquam non abutentes; praeterit enim figura huius mundi.
1COR|7|32|Volo autem vos sine sollicitudine esse. Qui sine uxore est, sollicitus est, quae Domini sunt, quomodo placeat Domino;
1COR|7|33|qui autem cum uxore est, sollicitus est, quae sunt mundi, quomodo placeat uxori,
1COR|7|34|et divisus est. Et mulier innupta et virgo cogitat, quae Domini sunt, ut sit sancta et corpore et spiritu; quae autem nupta est, cogitat, quae sunt mundi, quomodo placeat viro.
1COR|7|35|Porro hoc ad utilitatem vestram dico, non ut laqueum vobis iniciam, sed ad id quod honestum est, et ut assidue cum Domino sitis sine distractione.
1COR|7|36|Si quis autem turpem se videri existimat super virgine sua, quod sit superadulta, et ita oportet fieri, quod vult, faciat; non peccat: nubant.
1COR|7|37|Qui autem statuit in corde suo firmus, non habens necessitatem, potestatem autem habet suae voluntatis, et hoc iudicavit in corde suo servare virginem suam, bene faciet;
1COR|7|38|igitur et, qui matrimonio iungit virginem suam, bene facit; et, qui non iungit, melius faciet.
1COR|7|39|Mulier alligata est, quanto tempore vir eius vivit; quod si dormierit vir eius, libera est, cui vult nubere, tantum in Domino.
1COR|7|40|Beatior autem erit, si sic permanserit secundum meum consilium; puto autem quod et ego Spiritum Dei habeo.
1COR|8|1|De idolothytis autem, scimus quia omnes scientiam habemus. Scientia inflat, caritas vero aedificat.
1COR|8|2|Si quis se existimat scire aliquid, nondum cognovit, quemadmodum oporteat eum scire;
1COR|8|3|si quis autem diligit Deum, hic cognitus est ab eo.
1COR|8|4|De esu igitur idolothytorum, scimus quia nullum idolum est in mundo, et quod nullus deus nisi Unus.
1COR|8|5|Nam et si sunt, qui dicantur dii sive in caelo sive in terra, si quidem sunt dii multi et domini multi,
1COR|8|6|nobis tamen unus Deus Pater, ex quo omnia et nos in illum, et unus Dominus Iesus Christus, per quem omnia et nos per ipsum.
1COR|8|7|Sed non in omnibus est scientia; quidam autem consuetudine usque nunc idoli quasi idolothytum manducant, et conscientia ipsorum, cum sit infirma, polluitur.
1COR|8|8|Esca autem nos non commendat Deo; neque si non manducaverimus, deficiemus, neque si manducaverimus, abundabimus.
1COR|8|9|Videte autem, ne forte haec licentia vestra offendiculum fiat infirmis.
1COR|8|10|Si enim quis viderit eum, qui habet scientiam, in idolio recumbentem, nonne conscientia eius, cum sit infirma, aedificabitur ad manducandum idolothyta?
1COR|8|11|Peribit enim infirmus in tua scientia, frater, propter quem Christus mortuus est!
1COR|8|12|Sic autem peccantes in fratres et percutientes conscientiam eorum infirmam, in Christum peccatis.
1COR|8|13|Quapropter si esca scandalizat fratrem meum, non manducabo carnem in aeternum, ne fratrem meum scandalizem.
1COR|9|1|Non sum liber? Non sum apo stolus? Nonne Iesum Dominum nostrum vidi? Non opus meum vos estis in Domino?
1COR|9|2|Si aliis non sum apostolus, sed tamen vobis sum; nam signaculum apostolatus mei vos estis in Domino.
1COR|9|3|Mea defensio apud eos, qui me interrogant, haec est.
1COR|9|4|Numquid non habemus potestatem manducandi et bibendi?
1COR|9|5|Numquid non habemus potestatem sororem mulierem circumducendi, sicut et ceteri apostoli et fratres Domini et Cephas?
1COR|9|6|Aut solus ego et Barnabas non habemus potestatem non operandi?
1COR|9|7|Quis militat suis stipendiis umquam? Quis plantat vineam et fructum eius non edit? Aut quis pascit gregem et de lacte gregis non manducat?
1COR|9|8|Numquid secundum hominem haec dico? An et lex haec non dicit?
1COR|9|9|Scriptum est enim in Lege Moysis: " Non alligabis os bovi trituranti ". Numquid de bobus cura est Deo?
1COR|9|10|An propter nos utique dicit? Nam propter nos scripta sunt, quoniam debet in spe, qui arat, arare; et, qui triturat, in spe fructus percipiendi.
1COR|9|11|Si nos vobis spiritalia seminavimus, magnum est, si nos carnalia vestra metamus?
1COR|9|12|Si alii potestatis vestrae participes sunt, non potius nos? Sed non usi sumus hac potestate, sed omnia sustinemus, ne quod offendiculum demus evangelio Christi.
1COR|9|13|Nescitis quoniam, qui sacra operantur, quae de sacrario sunt, edunt; qui altari deserviunt, cum altari participantur?
1COR|9|14|Ita et Dominus ordinavit his, qui evangelium annuntiant, de evangelio vivere.
1COR|9|15|Ego autem nullo horum usus sum. Non scripsi autem haec, ut ita fiant in me; bonum est enim mihi magis mori quam ut gloriam meam quis evacuet.
1COR|9|16|Nam si evangelizavero, non est mihi gloria; necessitas enim mihi incumbit. Vae enim mihi est, si non evangelizavero!
1COR|9|17|Si enim volens hoc ago, mercedem habeo; si autem invitus, dispensatio mihi credita est.
1COR|9|18|Quae est ergo merces mea? Ut evangelium praedicans sine sumptu ponam evangelium, ut non abutar potestate mea in evangelio.
1COR|9|19|Nam cum liber essem ex omnibus, omnium me servum feci, ut plures lucri facerem.
1COR|9|20|Et factus sum Iudaeis tamquam Iudaeus, ut Iudaeos lucrarer; his, qui sub lege sunt, quasi sub lege essem, cum ipse non essem sub lege, ut eos, qui sub lege erant, lucri facerem;
1COR|9|21|his, qui sine lege erant, tamquam sine lege essem, cum sine lege Dei non essem, sed in lege essem Christi, ut lucri facerem eos, qui sine lege erant;
1COR|9|22|factus sum infirmis infirmus, ut infirmos lucri facerem; omnibus omnia factus sum, ut aliquos utique facerem salvos.
1COR|9|23|Omnia autem facio propter evangelium, ut comparticeps eius efficiar.
1COR|9|24|Nescitis quod hi, qui in stadio currunt, omnes quidem currunt, sed unus accipit bravium? Sic currite, ut comprehendatis.
1COR|9|25|Omnis autem, qui in agone contendit, ab omnibus se abstinet; et illi quidem, ut corruptibilem coronam accipiant, nos autem incorruptam.
1COR|9|26|Ego igitur sic curro non quasi in incertum, sic pugno non quasi aerem verberans;
1COR|9|27|sed castigo corpus meum et in servitutem redigo, ne forte, cum aliis praedicaverim, ipse reprobus efficiar.
1COR|10|1|Nolo enim vos ignorare, fra tres, quoniam patres nostri omnes sub nube fuerunt et omnes mare transierunt
1COR|10|2|et omnes in Moyse baptizati sunt in nube et in mari
1COR|10|3|et omnes eandem escam spiritalem manducaverunt
1COR|10|4|et omnes eundem potum spiritalem biberunt; bibebant autem de spiritali, consequente eos, petra; petra autem erat Christus.
1COR|10|5|Sed non in pluribus eorum complacuit sibi Deus, nam prostrati sunt in deserto.
1COR|10|6|Haec autem figurae fuerunt nostrae, ut non simus concupiscentes malorum, sicut et illi concupierunt.
1COR|10|7|Neque idolorum cultores efficiamini, sicut quidam ex ipsis; quemadmodum scriptum est: " Sedit populus manducare et bibere, et surrexerunt ludere.
1COR|10|8|Neque fornicemur, sicut quidam ex ipsis fornicati sunt, et ceciderunt una die viginti tria milia.
1COR|10|9|Neque tentemus Christum, sicut quidam eorum tentaverunt et a serpentibus perierunt.
1COR|10|10|Neque murmuraveritis, sicut quidam eorum murmuraverunt et perierunt ab exterminatore.
1COR|10|11|Haec autem in figura contingebant illis; scripta sunt autem ad correptionem nostram, in quos fines saeculorum devenerunt.
1COR|10|12|Itaque, qui se existimat stare, videat, ne cadat.
1COR|10|13|Tentatio vos non apprehendit nisi humana; fidelis autem Deus, qui non patietur vos tentari super id quod potestis, sed faciet cum tentatione etiam proventum, ut possitis sustinere.
1COR|10|14|Propter quod, carissimi mihi, fugite ab idolorum cultura.
1COR|10|15|Ut prudentibus loquor; vos iudicate, quod dico:
1COR|10|16|Calix benedictionis, cui benedicimus, nonne communicatio sanguinis Christi est? Et panis, quem frangimus, nonne communicatio corporis Christi est?
1COR|10|17|Quoniam unus panis, unum corpus multi sumus, omnes enim de uno pane participamur.
1COR|10|18|Videte Israel secundum carnem: nonne, qui edunt hostias, communicantes sunt altari?
1COR|10|19|Quid ergo dico? Quod idolothytum sit aliquid? Aut quod idolum sit aliquid?
1COR|10|20|Sed, quae immolant, daemoniis immolant et non Deo; nolo autem vos communicantes fieri daemoniis.
1COR|10|21|Non potestis calicem Domini bibere et calicem daemoniorum; non potestis mensae Domini participes esse et mensae daemoniorum.
1COR|10|22|An aemulamur Dominum? Numquid fortiores illo sumus?
1COR|10|23|" Omnia licent! ". Sed non omnia expediunt. " Omnia licent! ". Sed non omnia aedificant.
1COR|10|24|Nemo, quod suum est, quaerat, sed quod alterius.
1COR|10|25|Omne, quod in macello venit, manducate, nihil interrogantes propter conscientiam;
1COR|10|26|Domini enim est terra, et plenitudo eius.
1COR|10|27|Si quis vocat vos infidelium, et vultis ire, omne, quod vobis apponitur, manducate, nihil interrogantes propter conscientiam.
1COR|10|28|Si quis autem vobis dixerit: " Hoc immolaticium est idolis ", nolite manducare, propter illum, qui indicavit, et propter conscientiam;
1COR|10|29|conscientiam autem dico non tuam ipsius sed alterius. Ut quid enim libertas mea iudicatur ab alia conscientia?
1COR|10|30|Si ego cum gratia participo, quid blasphemor pro eo, quod gratias ago?
1COR|10|31|Sive ergo manducatis sive bibitis sive aliud quid facitis, omnia in gloriam Dei facite.
1COR|10|32|Sine offensione estote Iudaeis et Graecis et ecclesiae Dei,
1COR|10|33|sicut et ego per omnia omnibus placeo, non quaerens, quod mihi utile est, sed quod multis, ut salvi fiant.
1COR|11|1|Imitatores mei estote, sicut et ego Christi.
1COR|11|2|Laudo autem vos quod omnia mei memores estis et, sicut tradidi vobis, traditiones meas tenetis.
1COR|11|3|Volo autem vos scire quod omnis viri caput Christus est, caput autem mulieris vir, caput vero Christi Deus.
1COR|11|4|Omnis vir orans aut prophetans velato capite deturpat caput suum;
1COR|11|5|omnis autem mulier orans aut prophetans non velato capite deturpat caput suum; unum est enim atque si decalvetur.
1COR|11|6|Nam si non velatur mulier, et tondeatur! Si vero turpe est mulieri tonderi aut decalvari, veletur.
1COR|11|7|Vir quidem non debet velare caput, quoniam imago et gloria est Dei; mulier autem gloria viri est.
1COR|11|8|Non enim vir ex muliere est, sed mulier ex viro;
1COR|11|9|etenim non est creatus vir propter mulierem, sed mulier propter virum.
1COR|11|10|Ideo debet mulier potestatem habere supra caput propter angelos.
1COR|11|11|Verumtamen neque mulier sine viro, neque vir sine muliere in Domino;
1COR|11|12|nam sicut mulier de viro, ita et vir per mulierem, omnia autem ex Deo.
1COR|11|13|In vobis ipsi iudicate: Decet mulierem non velatam orare Deum?
1COR|11|14|Nec ipsa natura docet vos quod vir quidem, si comam nutriat, ignominia est illi;
1COR|11|15|mulier vero, si comam nutriat, gloria est illi? Quoniam coma pro velamine ei data est.
1COR|11|16|Si quis autem videtur contentiosus esse, nos talem consuetudinem non habemus, neque ecclesiae Dei.
1COR|11|17|Hoc autem praecipio, non laudans quod non in melius sed in deterius convenitis.
1COR|11|18|Primum quidem convenientibus vobis in ecclesia, audio scissuras inter vos esse et ex parte credo.
1COR|11|19|Nam oportet et haereses inter vos esse, ut et, qui probati sunt, manifesti fiant in vobis.
1COR|11|20|Convenientibus ergo vobis in unum, non est dominicam cenam manducare;
1COR|11|21|unusquisque enim suam cenam praesumit in manducando, et alius quidem esurit, alius autem ebrius est.
1COR|11|22|Numquid domos non habetis ad manducandum et bibendum? Aut ecclesiam Dei contemnitis et confunditis eos, qui non habent? Quid dicam vobis? Laudabo vos? In hoc non laudo!
1COR|11|23|Ego enim accepi a Domino, quod et tradidi vobis, quoniam Dominus Iesus, in qua nocte tradebatur, accepit panem
1COR|11|24|et gratias agens fregit et dixit: " Hoc est corpus meum, quod pro vobis est; hoc facite in meam commemorationem ";
1COR|11|25|similiter et calicem, postquam cenatum est, dicens: " Hic calix novum testamentum est in meo sanguine; hoc facite, quotiescumque bibetis, in meam commemorationem ".
1COR|11|26|Quotiescumque enim manducabitis panem hunc et calicem bibetis, mortem Domini annuntiatis, donec veniat.
1COR|11|27|Itaque, quicumque manducaverit panem vel biberit calicem Domini indigne, reus erit corporis et sanguinis Domini.
1COR|11|28|Probet autem seipsum homo, et sic de pane illo edat et de calice bibat;
1COR|11|29|qui enim manducat et bibit, iudicium sibi manducat et bibit non diiudicans corpus.
1COR|11|30|Ideo inter vos multi infirmi et imbecilles et dormiunt multi.
1COR|11|31|Quod si nosmetipsos diiudicaremus, non utique iudicaremur;
1COR|11|32|dum iudicamur autem, a Domino corripimur, ut non cum hoc mundo damnemur
1COR|11|33|Itaque, fratres mei, cum convenitis ad manducandum, invicem exspectate.
1COR|11|34|Si quis esurit, domi manducet, ut non in iudicium conveniatis. Cetera autem, cum venero, disponam.
1COR|12|1|De spiritalibus autem, fra tres, nolo vos ignorare.
1COR|12|2|Scitis quoniam, cum gentes essetis, ad simulacra muta, prout ducebamini, euntes.
1COR|12|3|Ideo notum vobis facio quod nemo in Spiritu Dei loquens dicit: " Anathema Iesus! "; et nemo potest dicere: " Dominus Iesus ", nisi in Spiritu Sancto.
1COR|12|4|Divisiones vero gratiarum sunt, idem autem Spiritus;
1COR|12|5|et divisiones ministrationum sunt, idem autem Dominus;
1COR|12|6|et divisiones operationum sunt, idem vero Deus, qui operatur omnia in omnibus.
1COR|12|7|Unicuique autem datur manifestatio Spiritus ad utilitatem.
1COR|12|8|Alii quidem per Spiritum datur sermo sapientiae, alii autem sermo scientiae secundum eundem Spiritum,
1COR|12|9|alteri fides in eodem Spiritu, alii donationes sanitatum in uno Spiritu,
1COR|12|10|alii operationes virtutum, alii prophetatio, alii discretio spirituum, alii genera linguarum, alii interpretatio linguarum;
1COR|12|11|haec autem omnia operatur unus et idem Spiritus, dividens singulis prout vult.
1COR|12|12|Sicut enim corpus unum est et membra habet multa, omnia autem membra corporis, cum sint multa, unum corpus sunt, ita et Christus;
1COR|12|13|etenim in uno Spiritu omnes nos in unum corpus baptizati sumus, sive Iudaei sive Graeci sive servi sive liberi, et omnes unum Spiritum potati sumus.
1COR|12|14|Nam et corpus non est unum membrum sed multa.
1COR|12|15|Si dixerit pes: "Non sum manus, non sum de corpore ", non ideo non est de corpore;
1COR|12|16|et si dixerit auris: " Non sum oculus, non sum de corpore ", non ideo non est de corpore.
1COR|12|17|Si totum corpus oculus est, ubi auditus? Si totum auditus, ubi odoratus?
1COR|12|18|Nunc autem posuit Deus membra, unumquodque eorum in corpore, sicut voluit.
1COR|12|19|Quod si essent omnia unum membrum, ubi corpus?
1COR|12|20|Nunc autem multa quidem membra, unum autem corpus.
1COR|12|21|Non potest dicere oculus manui: " Non es mihi necessaria! "; aut iterum caput pedibus: " Non estis mihi necessarii! ".
1COR|12|22|Sed multo magis, quae videntur membra corporis infirmiora esse, necessaria sunt;
1COR|12|23|et, quae putamus ignobiliora membra esse corporis, his honorem abundantiorem circumdamus; et, quae inhonesta sunt nostra, abundantiorem honestatem habent,
1COR|12|24|honesta autem nostra nullius egent. Sed Deus temperavit corpus, ei, cui deerat, abundantiorem tribuendo honorem,
1COR|12|25|ut non sit schisma in corpore, sed idipsum pro invicem sollicita sint membra.
1COR|12|26|Et sive patitur unum membrum, compatiuntur omnia membra; sive glorificatur unum membrum, congaudent omnia membra.
1COR|12|27|Vos autem estis corpus Christi et membra ex parte.
1COR|12|28|Et quosdam quidem posuit Deus in ecclesia primum apostolos, secundo prophetas, tertio doctores, deinde virtutes, exinde donationes curationum, opitulationes, gubernationes, genera linguarum.
1COR|12|29|Numquid omnes apostoli? Numquid omnes prophetae? Numquid omnes doctores? Numquid omnes virtutes?
1COR|12|30|Numquid omnes donationes habent curationum? Numquid omnes linguis loquuntur? Numquid omnes interpretantur?
1COR|12|31|Aemulamini autem charismata maiora. Et adhuc excellentiorem viam vobis demonstro.
1COR|13|1|Si linguis hominum loquar et angelorum, caritatem au tem non habeam, factus sum velut aes sonans aut cymbalum tinniens.
1COR|13|2|Et si habuero prophetiam et noverim mysteria omnia et omnem scientiam, et si habuero omnem fidem, ita ut montes transferam, caritatem autem non habuero, nihil sum.
1COR|13|3|Et si distribuero in cibos omnes facultates meas et si tradidero corpus meum, ut glorier, caritatem autem non habuero, nihil mihi prodest.
1COR|13|4|Caritas patiens est, benigna est caritas, non aemulatur, non agit superbe, non inflatur,
1COR|13|5|non est ambitiosa, non quaerit, quae sua sunt, non irritatur, non cogitat malum,
1COR|13|6|non gaudet super iniquitatem, congaudet autem veritati;
1COR|13|7|omnia suffert, omnia credit, omnia sperat, omnia sustinet.
1COR|13|8|Caritas numquam excidit. Sive prophetiae, evacuabuntur; sive linguae, cessabunt; sive scientia, destruetur.
1COR|13|9|Ex parte enim cognoscimus et ex parte prophetamus;
1COR|13|10|cum autem venerit, quod perfectum est, evacuabitur, quod ex parte est.
1COR|13|11|Cum essem parvulus, loquebar ut parvulus, sapiebam ut parvulus, cogitabam ut parvulus; quando factus sum vir, evacuavi, quae erant parvuli.
1COR|13|12|Videmus enim nunc per speculum in aenigmate, tunc autem facie ad faciem; nunc cognosco ex parte, tunc autem cognoscam, sicut et cognitus sum.
1COR|13|13|Nunc autem manet fides, spes, caritas, tria haec; maior autem ex his est caritas.
1COR|14|1|Sectamini caritatem, aemu lamini spiritalia, magis au tem, ut prophetetis.
1COR|14|2|Qui enim loquitur lingua, non hominibus loquitur sed Deo; nemo enim audit, spiritu autem loquitur mysteria.
1COR|14|3|Qui autem prophetat, hominibus loquitur aedificationem et exhortationem et consolationes.
1COR|14|4|Qui loquitur lingua, semetipsum aedificat; qui autem prophetat, ecclesiam aedificat.
1COR|14|5|Volo autem omnes vos loqui linguis, magis autem prophetare; maior autem est qui prophetat, quam qui loquitur linguis, nisi forte interpretetur, ut ecclesia aedificationem accipiat.
1COR|14|6|Nunc autem, fratres, si venero ad vos linguis loquens, quid vobis prodero, nisi vobis loquar aut in revelatione aut in scientia aut in prophetia aut in doctrina?
1COR|14|7|Tamen, quae sine anima sunt vocem dantia, sive tibia sive cithara, nisi distinctionem sonituum dederint, quomodo scietur quod tibia canitur, aut quod citharizatur?
1COR|14|8|Etenim si incertam vocem det tuba, quis parabit se ad bellum?
1COR|14|9|Ita et vos per linguam nisi manifestum sermonem dederitis, quomodo scietur id, quod dicitur? Eritis enim in aera loquentes.
1COR|14|10|Tam multa, ut puta, genera linguarum sunt in mundo, et nihil sine voce est.
1COR|14|11|Si ergo nesciero virtutem vocis, ero ei, qui loquitur, barbarus; et, qui loquitur, mihi barbarus.
1COR|14|12|Sic et vos, quoniam aemulatores estis spirituum, ad aedificationem ecclesiae quaerite, ut abundetis.
1COR|14|13|Et ideo, qui loquitur lingua, oret, ut interpretetur.
1COR|14|14|Nam si orem lingua, spiritus meus orat, mens autem mea sine fructu est.
1COR|14|15|Quid ergo est? Orabo spiritu, orabo et mente; psallam spiritu, psallam et mente.
1COR|14|16|Ceterum si benedixeris in spiritu, qui supplet locum idiotae, quomodo dicet " Amen! " super tuam benedictionem, quoniam quid dicas nescit?
1COR|14|17|Nam tu quidem bene gratias agis, sed alter non aedificatur.
1COR|14|18|Gratias ago Deo, quod omnium vestrum magis linguis loquor;
1COR|14|19|sed in ecclesia volo quinque verba sensu meo loqui, ut et alios instruam, quam decem milia verborum in lingua.
1COR|14|20|Fratres, nolite pueri effici sensibus, sed malitia parvuli estote; sensibus autem perfecti estote.
1COR|14|21|In lege scriptum est: In aliis linguis et in labiis aliorumloquar populo huic,et nec sic exaudient me ",dicit Dominus.
1COR|14|22|Itaque linguae in signum sunt non fidelibus sed infidelibus, prophetia autem non infidelibus sed fidelibus.
1COR|14|23|Si ergo conveniat universa ecclesia in unum, et omnes linguis loquantur, intrent autem idiotae aut infideles, nonne dicent quod insanitis?
1COR|14|24|Si autem omnes prophetent, intret autem quis infidelis vel idiota, convincitur ab omnibus, diiudicatur ab omnibus,
1COR|14|25|occulta cordis eius manifesta fiunt; et ita cadens in faciem adorabit Deum pronuntians: " Vere Deus in vobis est! ".
1COR|14|26|Quid ergo est, fratres? Cum convenitis, unusquisque psalmum habet, doctrinam habet, apocalypsim habet, linguam habet, interpretationem habet: omnia ad aedificationem fiant.
1COR|14|27|Sive lingua quis loquitur, secundum duos aut ut multum tres, et per partes, et unus interpretetur;
1COR|14|28|si autem non fuerit interpres, taceat in ecclesia, sibi autem loquatur et Deo.
1COR|14|29|Prophetae duo aut tres dicant, et ceteri diiudicent;
1COR|14|30|quod si alii revelatum fuerit sedenti, prior taceat.
1COR|14|31|Potestis enim omnes per singulos prophetare, ut omnes discant, et omnes exhortentur;
1COR|14|32|et spiritus prophetarum prophetis subiecti sunt;
1COR|14|33|non enim est dissensionis Deus sed pacis.Sicut in omnibus ecclesiis sanctorum,
1COR|14|34|mulieres in ecclesiis taceant, non enim permittitur eis loqui; sed subditae sint, sicut et Lex dicit.
1COR|14|35|Si quid autem volunt discere, domi viros suos interrogent; turpe est enim mulieri loqui in ecclesia.
1COR|14|36|An a vobis verbum Dei processit aut in vos solos pervenit?
1COR|14|37|Si quis videtur propheta esse aut spiritalis, cognoscat, quae scribo vobis, quia Domini est mandatum.
1COR|14|38|Si quis autem ignorat, ignorabitur.
1COR|14|39|Itaque, fratres mei, aemulamini prophetare et loqui linguis nolite prohibere;
1COR|14|40|omnia autem honeste et secundum ordinem fiant.
1COR|15|1|Notum autem vobis facio, fratres, evangelium, quod evangelizavi vobis, quod et accepistis, in quo et statis,
1COR|15|2|per quod et salvamini, qua ratione evangelizaverim vobis, si tenetis, nisi si frustra credidistis!
1COR|15|3|Tradidi enim vobis in primis, quod et accepi, quoniam Christus mortuus est pro peccatis nostris secundum Scripturas
1COR|15|4|et quia sepultus est et quia suscitatus est tertia die secundum Scripturas
1COR|15|5|et quia visus est Cephae et post haec Duodecim;
1COR|15|6|deinde visus est plus quam quingentis fratribus simul, ex quibus plures manent usque adhuc, quidam autem dormierunt;
1COR|15|7|deinde visus est Iacobo, deinde apostolis omnibus;
1COR|15|8|novissime autem omnium, tamquam abortivo, visus est et mihi.
1COR|15|9|Ego enim sum minimus apostolorum, qui non sum dignus vocari apostolus, quoniam persecutus sum ecclesiam Dei;
1COR|15|10|gratia autem Dei sum id, quod sum, et gratia eius in me vacua non fuit, sed abundantius illis omnibus laboravi; non ego autem, sed gratia Dei mecum.
1COR|15|11|Igitur sive ego sive illi, sic praedicamus, et sic credidistis.
1COR|15|12|Si autem Christus praedicatur quod suscitatus est a mortuis, quomodo quidam dicunt in vobis quoniam resurrectio mortuorum non est?
1COR|15|13|Si autem resurrectio mortuorum non est, neque Christus suscitatus est!
1COR|15|14|Si autem Christus non suscitatus est, inanis est ergo praedicatio nostra, inanis est et fides vestra;
1COR|15|15|invenimur autem et falsi testes Dei, quoniam testimonium diximus adversus Deum quod suscitaverit Christum, quem non suscitavit, si revera mortui non resurgunt.
1COR|15|16|Nam si mortui non resurgunt, neque Christus resurrexit;
1COR|15|17|quod si Christus non resurrexit, stulta est fides vestra; adhuc estis in peccatis vestris.
1COR|15|18|Ergo et, qui dormierunt in Christo, perierunt.
1COR|15|19|Si in hac vita tantum in Christo sperantes sumus, miserabiliores sumus omnibus hominibus.
1COR|15|20|Nunc autem Christus resurrexit a mortuis, primitiae dormientium.
1COR|15|21|Quoniam enim per hominem mors, et per hominem resurrectio mortuorum:
1COR|15|22|sicut enim in Adam omnes moriuntur, ita et in Christo omnes vivificabuntur.
1COR|15|23|Unusquisque autem in suo ordine: primitiae Christus; deinde hi, qui sunt Christi, in adventu eius;
1COR|15|24|deinde finis, cum tradiderit regnum Deo et Patri, cum evacuaverit omnem principatum et omnem potestatem et virtutem.
1COR|15|25|Oportet autem illum regnare, donec ponat omnes inimicos sub pedibus eius.
1COR|15|26|Novissima autem inimica destruetur mors;
1COR|15|27|omnia enim subiecit sub pedibus eius. Cum autem dicat: "Omnia subiecta sunt", sine dubio praeter eum, qui subiecit ei omnia.
1COR|15|28|Cum autem subiecta fuerint illi omnia, tunc ipse Filius subiectus erit illi, qui sibi subiecit omnia, ut sit Deus omnia in omnibus.
1COR|15|29|Alioquin quid facient, qui baptizantur pro mortuis? Si omnino mortui non resurgunt, ut quid et baptizantur pro illis?
1COR|15|30|Ut quid et nos periclitamur omni hora?
1COR|15|31|Cotidie morior, utique per vestram gloriationem, fratres, quam habeo in Christo Iesu Domino nostro!
1COR|15|32|Si secundum hominem ad bestias pugnavi Ephesi, quid mihi prodest? Si mortui non resurgunt, manducemus et bibamus, cras enim moriemur.
1COR|15|33|Noli te seduci: " Corrumpunt mores bonos colloquia mala ".
1COR|15|34|Evigilate iuste et nolite peccare! Ignorantiam enim Dei quidam ha bent; ad reverentiam vobis loquor.
1COR|15|35|Sed dicet aliquis: " Quomodo resurgunt mortui? Quali autem corpore veniunt? ".
1COR|15|36|Insipiens! Tu, quod seminas, non vivificatur, nisi prius moriatur;
1COR|15|37|et, quod seminas, non corpus, quod futurum est, seminas sed nudum granum, ut puta tritici aut alicuius ceterorum.
1COR|15|38|Deus autem dat illi corpus sicut voluit, et unicuique seminum proprium corpus.
1COR|15|39|Non omnis caro eadem caro, sed alia hominum, alia caro pecorum, alia caro volucrum, alia autem piscium.
1COR|15|40|Et corpora caelestia et corpora terrestria, sed alia quidem caelestium gloria, alia autem terrestrium.
1COR|15|41|Alia claritas solis, alia claritas lunae et alia claritas stellarum; stella enim a stella differt in claritate.
1COR|15|42|Sic et resurrectio mortuorum: seminatur in corruptione, resurgit in incorruptione;
1COR|15|43|seminatur in ignobilitate, resurgit in gloria; seminatur in infirmitate, resurgit in virtute;
1COR|15|44|seminatur corpus animale, resurgit corpus spiritale.Si est corpus animale, est et spiritale.
1COR|15|45|Sic et scriptum est: " Factus est primus homo Adam in animam viventem; novissimus Adam in Spiritum vivificantem.
1COR|15|46|Sed non prius, quod spiritale est, sed quod animale est; deinde quod spiritale.
1COR|15|47|Primus homo de terra terrenus, secundus homo de caelo.
1COR|15|48|Qualis terrenus, tales et terreni, et qualis caelestis, tales et caelestes;
1COR|15|49|et sicut portavimus imaginem terreni, portabimus et imaginem caelestis.
1COR|15|50|Hoc autem dico, fratres, quoniam caro et sanguis regnum Dei possidere non possunt, neque corruptio incorruptelam possidebit.
1COR|15|51|Ecce mysterium vobis dico: Non omnes quidem dormiemus, sed omnes immutabimur,
1COR|15|52|in momento, in ictu oculi, in novissima tuba; canet enim, et mortui suscitabuntur incorrupti, et nos immutabimur.
1COR|15|53|Oportet enim corruptibile hoc induere incorruptelam, et mortale induere immortalitatem.
1COR|15|54|Cum autem corruptibile hoc induerit incorruptelam, et mortale hoc induerit immortalitatem, tunc fiet sermo, qui scriptus est: " Absorpta est mors in victoria.
1COR|15|55|Ubi est, mors, victoria tua?Ubi est, mors, stimulus tuus? ".
1COR|15|56|Stimulus autem mortis peccatum est, virtus vero peccati lex.
1COR|15|57|Deo autem gratias, qui dedit nobis victoriam per Dominum nostrum Iesum Christum.
1COR|15|58|Itaque, fratres mei dilecti, stabiles estote, immobiles, abundantes in opere Domini semper, scientes quod labor vester non est inanis in Domino.
1COR|16|1|De collectis autem, quae fiunt in sanctos, sicut ordina vi ecclesiis Galatiae, ita et vos facite.
1COR|16|2|Per primam sabbati unusquisque vestrum apud se ponat recondens, quod ei beneplacuerit, ut non, cum venero, tunc collectae fiant.
1COR|16|3|Cum autem praesens fuero, quos probaveritis, per epistulas hos mittam perferre gratiam vestram in Ierusalem;
1COR|16|4|quod si dignum fuerit, ut et ego eam, mecum ibunt.
1COR|16|5|Veniam autem ad vos, cum Macedoniam pertransiero, nam Macedoniam pertransibo;
1COR|16|6|apud vos autem forsitan manebo vel etiam hiemabo, ut vos me deducatis, quocumque iero.
1COR|16|7|Nolo enim vos modo in transitu videre; spero enim me aliquantum temporis manere apud vos, si Dominus permiserit.
1COR|16|8|Permanebo autem Ephesi usque ad Pentecosten;
1COR|16|9|ostium enim mihi apertum est magnum et efficax, et adversarii multi.
1COR|16|10|Si autem venerit Timotheus, videte, ut sine timore sit apud vos, opus enim Domini operatur, sicut et ego;
1COR|16|11|ne quis ergo illum spernat. Deducite autem illum in pace, ut veniat ad me; exspecto enim illum cum fratribus.
1COR|16|12|De Apollo autem fratre, multum rogavi eum, ut veniret ad vos cum fratribus, et utique non fuit voluntas, ut nunc veniret; veniet autem, cum ei opportunum fuerit.
1COR|16|13|Vigilate, state in fide, viriliter agite, confortamini;
1COR|16|14|omnia vestra in caritate fiant.
1COR|16|15|Obsecro autem vos, fratres: nostis domum Stephanae, quoniam sunt primitiae Achaiae et in ministerium sanctorum ordinaverunt seipsos;
1COR|16|16|ut et vos subditi sitis eiusmodi et omni cooperanti et laboranti.
1COR|16|17|Gaudeo autem in praesentia Stephanae et Fortunati et Achaici, quoniam id quod vobis deerat, ipsi suppleverunt;
1COR|16|18|refecerunt enim et meum spiritum et vestrum. Cognoscite ergo, qui eiusmodi sunt.
1COR|16|19|Salutant vos ecclesiae Asiae. Salutant vos in Domino multum Aquila et Prisca cum domestica sua ecclesia.
1COR|16|20|Salutant vos fratres omnes. Salutate invicem in osculo sancto.
1COR|16|21|Salutatio mea manu Pauli.
1COR|16|22|Si quis non amat Dominum, sit anathema. Marana tha!
1COR|16|23|Gratia Domini Iesu vobiscum.
1COR|16|24|Caritas mea cum omnibus vobis in Christo Iesu.
