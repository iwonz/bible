ECCL|1|1|Слова Екклесиаста, сына Давидова, царя в Иерусалиме.
ECCL|1|2|Суета сует, сказал Екклесиаст, суета сует, – все суета!
ECCL|1|3|Что пользы человеку от всех трудов его, которыми трудится он под солнцем?
ECCL|1|4|Род проходит, и род приходит, а земля пребывает во веки.
ECCL|1|5|Восходит солнце, и заходит солнце, и спешит к месту своему, где оно восходит.
ECCL|1|6|Идет ветер к югу, и переходит к северу, кружится, кружится на ходу своем, и возвращается ветер на круги свои.
ECCL|1|7|Все реки текут в море, но море не переполняется: к тому месту, откуда реки текут, они возвращаются, чтобы опять течь.
ECCL|1|8|Все вещи – в труде: не может человек пересказать всего; не насытится око зрением, не наполнится ухо слушанием.
ECCL|1|9|Что было, то и будет; и что делалось, то и будет делаться, и нет ничего нового под солнцем.
ECCL|1|10|Бывает нечто, о чем говорят: "смотри, вот это новое"; но [это] было уже в веках, бывших прежде нас.
ECCL|1|11|Нет памяти о прежнем; да и о том, что будет, не останется памяти у тех, которые будут после.
ECCL|1|12|Я, Екклесиаст, был царем над Израилем в Иерусалиме;
ECCL|1|13|и предал я сердце мое тому, чтобы исследовать и испытать мудростью все, что делается под небом: это тяжелое занятие дал Бог сынам человеческим, чтобы они упражнялись в нем.
ECCL|1|14|Видел я все дела, какие делаются под солнцем, и вот, все – суета и томление духа!
ECCL|1|15|Кривое не может сделаться прямым, и чего нет, того нельзя считать.
ECCL|1|16|Говорил я с сердцем моим так: вот, я возвеличился и приобрел мудрости больше всех, которые были прежде меня над Иерусалимом, и сердце мое видело много мудрости и знания.
ECCL|1|17|И предал я сердце мое тому, чтобы познать мудрость и познать безумие и глупость: узнал, что и это – томление духа;
ECCL|1|18|потому что во многой мудрости много печали; и кто умножает познания, умножает скорбь.
ECCL|2|1|Сказал я в сердце моем: "дай, испытаю я тебя весельем, и насладись добром"; но и это – суета!
ECCL|2|2|О смехе сказал я: "глупость!", а о веселье: "что оно делает?"
ECCL|2|3|Вздумал я в сердце моем услаждать вином тело мое и, между тем, как сердце мое руководилось мудростью, придержаться и глупости, доколе не увижу, что хорошо для сынов человеческих, что должны были бы они делать под небом в немногие дни жизни своей.
ECCL|2|4|Я предпринял большие дела: построил себе домы, посадил себе виноградники,
ECCL|2|5|устроил себе сады и рощи и насадил в них всякие плодовитые дерева;
ECCL|2|6|сделал себе водоемы для орошения из них рощей, произращающих деревья;
ECCL|2|7|приобрел себе слуг и служанок, и домочадцы были у меня; также крупного и мелкого скота было у меня больше, нежели у всех, бывших прежде меня в Иерусалиме;
ECCL|2|8|собрал себе серебра и золота и драгоценностей от царей и областей; завел у себя певцов и певиц и услаждения сынов человеческих – разные музыкальные орудия.
ECCL|2|9|И сделался я великим и богатым больше всех, бывших прежде меня в Иерусалиме; и мудрость моя пребыла со мною.
ECCL|2|10|Чего бы глаза мои ни пожелали, я не отказывал им, не возбранял сердцу моему никакого веселья, потому что сердце мое радовалось во всех трудах моих, и это было моею долею от всех трудов моих.
ECCL|2|11|И оглянулся я на все дела мои, которые сделали руки мои, и на труд, которым трудился я, делая [их]: и вот, все – суета и томление духа, и нет [от них] пользы под солнцем!
ECCL|2|12|И обратился я, чтобы взглянуть на мудрость и безумие и глупость: ибо что [может сделать] человек после царя [сверх того], что уже сделано?
ECCL|2|13|И увидел я, что преимущество мудрости перед глупостью такое же, как преимущество света перед тьмою:
ECCL|2|14|у мудрого глаза его – в голове его, а глупый ходит во тьме; но узнал я, что одна участь постигает их всех.
ECCL|2|15|И сказал я в сердце моем: "и меня постигнет та же участь, как и глупого: к чему же я сделался очень мудрым?" И сказал я в сердце моем, что и это – суета;
ECCL|2|16|потому что мудрого не будут помнить вечно, как и глупого; в грядущие дни все будет забыто, и увы! мудрый умирает наравне с глупым.
ECCL|2|17|И возненавидел я жизнь, потому что противны стали мне дела, которые делаются под солнцем; ибо все – суета и томление духа!
ECCL|2|18|И возненавидел я весь труд мой, которым трудился под солнцем, потому что должен оставить его человеку, который будет после меня.
ECCL|2|19|И кто знает: мудрый ли будет он, или глупый? А он будет распоряжаться всем трудом моим, которым я трудился и которым показал себя мудрым под солнцем. И это – суета!
ECCL|2|20|И обратился я, чтобы внушить сердцу моему отречься от всего труда, которым я трудился под солнцем,
ECCL|2|21|потому что иной человек трудится мудро, с знанием и успехом, и должен отдать все человеку, не трудившемуся в том, как бы часть его. И это – суета и зло великое!
ECCL|2|22|Ибо что будет иметь человек от всего труда своего и заботы сердца своего, что трудится он под солнцем?
ECCL|2|23|Потому что все дни его – скорби, и его труды – беспокойство; даже и ночью сердце его не знает покоя. И это – суета!
ECCL|2|24|Не во власти человека и то благо, чтобы есть и пить и услаждать душу свою от труда своего. Я увидел, что и это – от руки Божией;
ECCL|2|25|потому что кто может есть и кто может наслаждаться без Него?
ECCL|2|26|Ибо человеку, который добр пред лицем Его, Он дает мудрость и знание и радость; а грешнику дает заботу собирать и копить, чтобы [после] отдать доброму пред лицем Божиим. И это – суета и томление духа!
ECCL|3|1|Всему свое время, и время всякой вещи под небом:
ECCL|3|2|время рождаться, и время умирать; время насаждать, и время вырывать посаженное;
ECCL|3|3|время убивать, и время врачевать; время разрушать, и время строить;
ECCL|3|4|время плакать, и время смеяться; время сетовать, и время плясать;
ECCL|3|5|время разбрасывать камни, и время собирать камни; время обнимать, и время уклоняться от объятий;
ECCL|3|6|время искать, и время терять; время сберегать, и время бросать;
ECCL|3|7|время раздирать, и время сшивать; время молчать, и время говорить;
ECCL|3|8|время любить, и время ненавидеть; время войне, и время миру.
ECCL|3|9|Что пользы работающему от того, над чем он трудится?
ECCL|3|10|Видел я эту заботу, которую дал Бог сынам человеческим, чтобы они упражнялись в том.
ECCL|3|11|Все соделал Он прекрасным в свое время, и вложил мир в сердце их, хотя человек не может постигнуть дел, которые Бог делает, от начала до конца.
ECCL|3|12|Познал я, что нет для них ничего лучшего, как веселиться и делать доброе в жизни своей.
ECCL|3|13|И если какой человек ест и пьет, и видит доброе во всяком труде своем, то это – дар Божий.
ECCL|3|14|Познал я, что все, что делает Бог, пребывает вовек: к тому нечего прибавлять и от того нечего убавить, – и Бог делает так, чтобы благоговели пред лицем Его.
ECCL|3|15|Что было, то и теперь есть, и что будет, то уже было, – и Бог воззовет прошедшее.
ECCL|3|16|Еще видел я под солнцем: место суда, а там беззаконие; место правды, а там неправда.
ECCL|3|17|И сказал я в сердце своем: "праведного и нечестивого будет судить Бог; потому что время для всякой вещи и [суд] над всяким делом там".
ECCL|3|18|Сказал я в сердце своем о сынах человеческих, чтобы испытал их Бог, и чтобы они видели, что они сами по себе животные;
ECCL|3|19|потому что участь сынов человеческих и участь животных – участь одна: как те умирают, так умирают и эти, и одно дыхание у всех, и нет у человека преимущества перед скотом, потому что все – суета!
ECCL|3|20|Все идет в одно место: все произошло из праха и все возвратится в прах.
ECCL|3|21|Кто знает: дух сынов человеческих восходит ли вверх, и дух животных сходит ли вниз, в землю?
ECCL|3|22|Итак увидел я, что нет ничего лучше, как наслаждаться человеку делами своими: потому что это – доля его; ибо кто приведет его посмотреть на то, что будет после него?
ECCL|4|1|И обратился я и увидел всякие угнетения, какие делаются под солнцем: и вот слезы угнетенных, а утешителя у них нет; и в руке угнетающих их – сила, а утешителя у них нет.
ECCL|4|2|И ублажил я мертвых, которые давно умерли, более живых, которые живут доселе;
ECCL|4|3|а блаженнее их обоих тот, кто еще не существовал, кто не видал злых дел, какие делаются под солнцем.
ECCL|4|4|Видел я также, что всякий труд и всякий успех в делах производят взаимную между людьми зависть. И это – суета и томление духа!
ECCL|4|5|Глупый [сидит], сложив свои руки, и съедает плоть свою.
ECCL|4|6|Лучше горсть с покоем, нежели пригоршни с трудом и томлением духа.
ECCL|4|7|И обратился я и увидел еще суету под солнцем;
ECCL|4|8|[человек] одинокий, и другого нет; ни сына, ни брата нет у него; а всем трудам его нет конца, и глаз его не насыщается богатством. "Для кого же я тружусь и лишаю душу мою блага?" И это – суета и недоброе дело!
ECCL|4|9|Двоим лучше, нежели одному; потому что у них есть доброе вознаграждение в труде их:
ECCL|4|10|ибо если упадет один, то другой поднимет товарища своего. Но горе одному, когда упадет, а другого нет, который поднял бы его.
ECCL|4|11|Также, если лежат двое, то тепло им; а одному как согреться?
ECCL|4|12|И если станет преодолевать кто–либо одного, то двое устоят против него: и нитка, втрое скрученная, нескоро порвется.
ECCL|4|13|Лучше бедный, но умный юноша, нежели старый, но неразумный царь, который не умеет принимать советы;
ECCL|4|14|ибо тот из темницы выйдет на царство, хотя родился в царстве своем бедным.
ECCL|4|15|Видел я всех живущих, которые ходят под солнцем, с этим другим юношею, который займет место того.
ECCL|4|16|Не было числа всему народу, который был перед ним, хотя позднейшие не порадуются им. И это – суета и томление духа!
ECCL|4|17|Наблюдай за ногою твоею, когда идешь в дом Божий, и будь готов более к слушанию, нежели к жертвоприношению; ибо они не думают, что худо делают.
ECCL|5|1|Не торопись языком твоим, и сердце твое да не спешит произнести слово пред Богом; потому что Бог на небе, а ты на земле; поэтому слова твои да будут немноги.
ECCL|5|2|Ибо, как сновидения бывают при множестве забот, так голос глупого познается при множестве слов.
ECCL|5|3|Когда даешь обет Богу, то не медли исполнить его, потому что Он не благоволит к глупым: что обещал, исполни.
ECCL|5|4|Лучше тебе не обещать, нежели обещать и не исполнить.
ECCL|5|5|Не дозволяй устам твоим вводить в грех плоть твою, и не говори пред Ангелом [Божиим]: "это – ошибка!" Для чего тебе [делать], чтобы Бог прогневался на слово твое и разрушил дело рук твоих?
ECCL|5|6|Ибо во множестве сновидений, как и во множестве слов, – много суеты; но ты бойся Бога.
ECCL|5|7|Если ты увидишь в какой области притеснение бедному и нарушение суда и правды, то не удивляйся этому: потому что над высоким наблюдает высший, а над ними еще высший;
ECCL|5|8|превосходство же страны в целом есть царь, заботящийся о стране.
ECCL|5|9|Кто любит серебро, тот не насытится серебром, и кто любит богатство, тому нет пользы от того. И это – суета!
ECCL|5|10|Умножается имущество, умножаются и потребляющие его; и какое благо для владеющего им: разве только смотреть своими глазами?
ECCL|5|11|Сладок сон трудящегося, мало ли, много ли он съест; но пресыщение богатого не дает ему уснуть.
ECCL|5|12|Есть мучительный недуг, который видел я под солнцем: богатство, сберегаемое владетелем его во вред ему.
ECCL|5|13|И гибнет богатство это от несчастных случаев: родил он сына, и ничего нет в руках у него.
ECCL|5|14|Как вышел он нагим из утробы матери своей, таким и отходит, каким пришел, и ничего не возьмет от труда своего, что мог бы он понести в руке своей.
ECCL|5|15|И это тяжкий недуг: каким пришел он, таким и отходит. Какая же польза ему, что он трудился на ветер?
ECCL|5|16|А он во все дни свои ел впотьмах, в большом раздражении, в огорчении и досаде.
ECCL|5|17|Вот еще, что я нашел доброго и приятного: есть и пить и наслаждаться добром во всех трудах своих, какими кто трудится под солнцем во все дни жизни своей, которые дал ему Бог; потому что это его доля.
ECCL|5|18|И если какому человеку Бог дал богатство и имущество, и дал ему власть пользоваться от них и брать свою долю и наслаждаться от трудов своих, то это дар Божий.
ECCL|5|19|Недолго будут у него в памяти дни жизни его; потому Бог и вознаграждает его радостью сердца его.
ECCL|6|1|Есть зло, которое видел я под солнцем, и оно часто бывает между людьми:
ECCL|6|2|Бог дает человеку богатство и имущество и славу, и нет для души его недостатка ни в чем, чего не пожелал бы он; но не дает ему Бог пользоваться этим, а пользуется тем чужой человек: это – суета и тяжкий недуг!
ECCL|6|3|Если бы какой человек родил сто [детей], и прожил многие годы, и еще умножились дни жизни его, но душа его не наслаждалась бы добром и не было бы ему и погребения, то я сказал бы: выкидыш счастливее его,
ECCL|6|4|потому что он напрасно пришел и отошел во тьму, и его имя покрыто мраком.
ECCL|6|5|Он даже не видел и не знал солнца: ему покойнее, нежели тому.
ECCL|6|6|А тот, хотя бы прожил две тысячи лет и не наслаждался добром, не все ли пойдет в одно место?
ECCL|6|7|Все труды человека – для рта его, а душа его не насыщается.
ECCL|6|8|Какое же преимущество мудрого перед глупым, какое – бедняка, умеющего ходить перед живущими?
ECCL|6|9|Лучше видеть глазами, нежели бродить душею. И это – также суета и томление духа!
ECCL|6|10|Что существует, тому уже наречено имя, и известно, что это – человек, и что он не может препираться с тем, кто сильнее его.
ECCL|6|11|Много таких вещей, которые умножают суету: что же для человека лучше?
ECCL|6|12|Ибо кто знает, что хорошо для человека в жизни, во все дни суетной жизни его, которые он проводит как тень? И кто скажет человеку, что будет после него под солнцем?
ECCL|7|1|Доброе имя лучше дорогой масти, и день смерти – дня рождения.
ECCL|7|2|Лучше ходить в дом плача об умершем, нежели ходить в дом пира; ибо таков конец всякого человека, и живой приложит [это] к своему сердцу.
ECCL|7|3|Сетование лучше смеха; потому что при печали лица сердце делается лучше.
ECCL|7|4|Сердце мудрых – в доме плача, а сердце глупых – в доме веселья.
ECCL|7|5|Лучше слушать обличения от мудрого, нежели слушать песни глупых;
ECCL|7|6|потому что смех глупых то же, что треск тернового хвороста под котлом. И это – суета!
ECCL|7|7|Притесняя других, мудрый делается глупым, и подарки портят сердце.
ECCL|7|8|Конец дела лучше начала его; терпеливый лучше высокомерного.
ECCL|7|9|Не будь духом твоим поспешен на гнев, потому что гнев гнездится в сердце глупых.
ECCL|7|10|Не говори: "отчего это прежние дни были лучше нынешних?", потому что не от мудрости ты спрашиваешь об этом.
ECCL|7|11|Хороша мудрость с наследством, и особенно для видящих солнце:
ECCL|7|12|потому что под сенью ее [то же, что] под сенью серебра; но превосходство знания в [том, что] мудрость дает жизнь владеющему ею.
ECCL|7|13|Смотри на действование Божие: ибо кто может выпрямить то, что Он сделал кривым?
ECCL|7|14|Во дни благополучия пользуйся благом, а во дни несчастья размышляй: то и другое соделал Бог для того, чтобы человек ничего не мог сказать против Него.
ECCL|7|15|Всего насмотрелся я в суетные дни мои: праведник гибнет в праведности своей; нечестивый живет долго в нечестии своем.
ECCL|7|16|Не будь слишком строг, и не выставляй себя слишком мудрым; зачем тебе губить себя?
ECCL|7|17|Не предавайся греху, и не будь безумен: зачем тебе умирать не в свое время?
ECCL|7|18|Хорошо, если ты будешь держаться одного и не отнимать руки от другого; потому что кто боится Бога, тот избежит всего того.
ECCL|7|19|Мудрость делает мудрого сильнее десяти властителей, которые в городе.
ECCL|7|20|Нет человека праведного на земле, который делал бы добро и не грешил бы;
ECCL|7|21|поэтому не на всякое слово, которое говорят, обращай внимание, чтобы не услышать тебе раба твоего, когда он злословит тебя;
ECCL|7|22|ибо сердце твое знает много случаев, когда и сам ты злословил других.
ECCL|7|23|Все это испытал я мудростью; я сказал: "буду я мудрым"; но мудрость далека от меня.
ECCL|7|24|Далеко то, что было, и глубоко – глубоко: кто постигнет его?
ECCL|7|25|Обратился я сердцем моим к тому, чтобы узнать, исследовать и изыскать мудрость и разум, и познать нечестие глупости, невежества и безумия, –
ECCL|7|26|и нашел я, что горче смерти женщина, потому что она – сеть, и сердце ее – силки, руки ее – оковы; добрый пред Богом спасется от нее, а грешник уловлен будет ею.
ECCL|7|27|Вот это нашел я, сказал Екклесиаст, испытывая одно за другим.
ECCL|7|28|Чего еще искала душа моя, и я не нашел? – Мужчину одного из тысячи я нашел, а женщину между всеми ими не нашел.
ECCL|7|29|Только это я нашел, что Бог сотворил человека правым, а люди пустились во многие помыслы.
ECCL|8|1|Кто – как мудрый, и кто понимает значение вещей? Мудрость человека просветляет лице его, и суровость лица его изменяется.
ECCL|8|2|[Я говорю]: слово царское храни, и [это] ради клятвы пред Богом.
ECCL|8|3|Не спеши уходить от лица его, и не упорствуй в худом деле; потому что он, что захочет, все может сделать.
ECCL|8|4|Где слово царя, там власть; и кто скажет ему: "что ты делаешь?"
ECCL|8|5|Соблюдающий заповедь не испытает никакого зла: сердце мудрого знает и время и устав;
ECCL|8|6|потому что для всякой вещи есть свое время и устав; а человеку великое зло от того,
ECCL|8|7|что он не знает, что будет; и как это будет – кто скажет ему?
ECCL|8|8|Человек не властен над духом, чтобы удержать дух, и нет власти у него над днем смерти, и нет избавления в этой борьбе, и не спасет нечестие нечестивого.
ECCL|8|9|Все это я видел, и обращал сердце мое на всякое дело, какое делается под солнцем. Бывает время, когда человек властвует над человеком во вред ему.
ECCL|8|10|Видел я тогда, что хоронили нечестивых, и приходили и отходили от святого места, и они забываемы были в городе, где они так поступали. И это – суета!
ECCL|8|11|Не скоро совершается суд над худыми делами; от этого и не страшится сердце сынов человеческих делать зло.
ECCL|8|12|Хотя грешник сто раз делает зло и коснеет в нем, но я знаю, что благо будет боящимся Бога, которые благоговеют пред лицем Его;
ECCL|8|13|а нечестивому не будет добра, и, подобно тени, недолго продержится тот, кто не благоговеет пред Богом.
ECCL|8|14|Есть и такая суета на земле: праведников постигает то, чего заслуживали бы дела нечестивых, а с нечестивыми бывает то, чего заслуживали бы дела праведников. И сказал я: и это – суета!
ECCL|8|15|И похвалил я веселье; потому что нет лучшего для человека под солнцем, как есть, пить и веселиться: это сопровождает его в трудах во дни жизни его, которые дал ему Бог под солнцем.
ECCL|8|16|Когда я обратил сердце мое на то, чтобы постигнуть мудрость и обозреть дела, которые делаются на земле, и среди которых [человек] ни днем, ни ночью не знает сна, –
ECCL|8|17|тогда я увидел все дела Божии и [нашел], что человек не может постигнуть дел, которые делаются под солнцем. Сколько бы человек ни трудился в исследовании, он все–таки не постигнет этого; и если бы какой мудрец сказал, что он знает, он не может постигнуть [этого].
ECCL|9|1|На все это я обратил сердце мое для исследования, что праведные и мудрые и деяния их – в руке Божией, и что человек ни любви, ни ненависти не знает во всем том, что перед ним.
ECCL|9|2|Всему и всем – одно: одна участь праведнику и нечестивому, доброму и [злому], чистому и нечистому, приносящему жертву и не приносящему жертвы; как добродетельному, так и грешнику; как клянущемуся, так и боящемуся клятвы.
ECCL|9|3|Это–то и худо во всем, что делается под солнцем, что одна участь всем, и сердце сынов человеческих исполнено зла, и безумие в сердце их, в жизни их; а после того они [отходят] к умершим.
ECCL|9|4|Кто находится между живыми, тому есть еще надежда, так как и псу живому лучше, нежели мертвому льву.
ECCL|9|5|Живые знают, что умрут, а мертвые ничего не знают, и уже нет им воздаяния, потому что и память о них предана забвению,
ECCL|9|6|и любовь их и ненависть их и ревность их уже исчезли, и нет им более части во веки ни в чем, что делается под солнцем.
ECCL|9|7|[Итак] иди, ешь с весельем хлеб твой, и пей в радости сердца вино твое, когда Бог благоволит к делам твоим.
ECCL|9|8|Да будут во всякое время одежды твои светлы, и да не оскудевает елей на голове твоей.
ECCL|9|9|Наслаждайся жизнью с женою, которую любишь, во все дни суетной жизни твоей, и которую дал тебе Бог под солнцем на все суетные дни твои; потому что это – доля твоя в жизни и в трудах твоих, какими ты трудишься под солнцем.
ECCL|9|10|Все, что может рука твоя делать, по силам делай; потому что в могиле, куда ты пойдешь, нет ни работы, ни размышления, ни знания, ни мудрости.
ECCL|9|11|И обратился я, и видел под солнцем, что не проворным достается успешный бег, не храбрым – победа, не мудрым – хлеб, и не у разумных – богатство, и не искусным – благорасположение, но время и случай для всех их.
ECCL|9|12|Ибо человек не знает своего времени. Как рыбы попадаются в пагубную сеть, и как птицы запутываются в силках, так сыны человеческие уловляются в бедственное время, когда оно неожиданно находит на них.
ECCL|9|13|Вот еще какую мудрость видел я под солнцем, и она показалась мне важною:
ECCL|9|14|город небольшой, и людей в нем немного; к нему подступил великий царь и обложил его и произвел против него большие осадные работы;
ECCL|9|15|но в нем нашелся мудрый бедняк, и он спас своею мудростью этот город; и однако же никто не вспоминал об этом бедном человеке.
ECCL|9|16|И сказал я: мудрость лучше силы, и однако же мудрость бедняка пренебрегается, и слов его не слушают.
ECCL|9|17|Слова мудрых, [высказанные] спокойно, выслушиваются [лучше], нежели крик властелина между глупыми.
ECCL|9|18|Мудрость лучше воинских орудий; но один погрешивший погубит много доброго.
ECCL|10|1|Мертвые мухи портят и делают зловонною благовонную масть мироварника: то же делает небольшая глупость уважаемого человека с его мудростью и честью.
ECCL|10|2|Сердце мудрого – на правую сторону, а сердце глупого – на левую.
ECCL|10|3|По какой бы дороге ни шел глупый, у него [всегда] недостает смысла, и всякому он выскажет, что он глуп.
ECCL|10|4|Если гнев начальника вспыхнет на тебя, то не оставляй места твоего; потому что кротость покрывает и большие проступки.
ECCL|10|5|Есть зло, которое видел я под солнцем, это – как бы погрешность, происходящая от властелина;
ECCL|10|6|невежество поставляется на большой высоте, а богатые сидят низко.
ECCL|10|7|Видел я рабов на конях, а князей ходящих, подобно рабам, пешком.
ECCL|10|8|Кто копает яму, тот упадет в нее, и кто разрушает ограду, того ужалит змей.
ECCL|10|9|Кто передвигает камни, тот может надсадить себя, и кто колет дрова, тот может подвергнуться опасности от них.
ECCL|10|10|Если притупится топор, и если лезвие его не будет отточено, то надобно будет напрягать силы; мудрость умеет это исправить.
ECCL|10|11|Если змей ужалит без заговаривания, то не лучше его и злоязычный.
ECCL|10|12|Слова из уст мудрого – благодать, а уста глупого губят его же:
ECCL|10|13|начало слов из уст его – глупость, [а] конец речи из уст его – безумие.
ECCL|10|14|Глупый наговорит много, [хотя] человек не знает, что будет, и кто скажет ему, что будет после него?
ECCL|10|15|Труд глупого утомляет его, потому что не знает [даже] дороги в город.
ECCL|10|16|Горе тебе, земля, когда царь твой отрок, и когда князья твои едят рано!
ECCL|10|17|Благо тебе, земля, когда царь у тебя из благородного рода, и князья твои едят вовремя, для подкрепления, а не для пресыщения!
ECCL|10|18|От лености обвиснет потолок, и когда опустятся руки, то протечет дом.
ECCL|10|19|Пиры устраиваются для удовольствия, и вино веселит жизнь; а за все отвечает серебро.
ECCL|10|20|Даже и в мыслях твоих не злословь царя, и в спальной комнате твоей не злословь богатого; потому что птица небесная может перенести слово [твое], и крылатая – пересказать речь [твою].
ECCL|11|1|Отпускай хлеб твой по водам, потому что по прошествии многих дней опять найдешь его.
ECCL|11|2|Давай часть семи и даже восьми, потому что не знаешь, какая беда будет на земле.
ECCL|11|3|Когда облака будут полны, то они прольют на землю дождь; и если упадет дерево на юг или на север, то оно там и останется, куда упадет.
ECCL|11|4|Кто наблюдает ветер, тому не сеять; и кто смотрит на облака, тому не жать.
ECCL|11|5|Как ты не знаешь путей ветра и того, как [образуются] кости во чреве беременной, так не можешь знать дело Бога, Который делает все.
ECCL|11|6|Утром сей семя твое, и вечером не давай отдыха руке твоей, потому что ты не знаешь, то или другое будет удачнее, или то и другое равно хорошо будет.
ECCL|11|7|Сладок свет, и приятно для глаз видеть солнце.
ECCL|11|8|Если человек проживет [и] много лет, то пусть веселится он в продолжение всех их, и пусть помнит о днях темных, которых будет много: все, что будет, – суета!
ECCL|11|9|Веселись, юноша, в юности твоей, и да вкушает сердце твое радости во дни юности твоей, и ходи по путям сердца твоего и по видению очей твоих; только знай, что за все это Бог приведет тебя на суд.
ECCL|11|10|И удаляй печаль от сердца твоего, и уклоняй злое от тела твоего, потому что детство и юность – суета.
ECCL|12|1|И помни Создателя твоего в дни юности твоей, доколе не пришли тяжелые дни и не наступили годы, о которых ты будешь говорить: "нет мне удовольствия в них!"
ECCL|12|2|доколе не померкли солнце и свет и луна и звезды, и не нашли новые тучи вслед за дождем.
ECCL|12|3|В тот день, когда задрожат стерегущие дом и согнутся мужи силы; и перестанут молоть мелющие, потому что их немного осталось; и помрачатся смотрящие в окно;
ECCL|12|4|и запираться будут двери на улицу; когда замолкнет звук жернова, и будет вставать [человек] по крику петуха и замолкнут дщери пения;
ECCL|12|5|и высоты будут им страшны, и на дороге ужасы; и зацветет миндаль, и отяжелеет кузнечик, и рассыплется каперс. Ибо отходит человек в вечный дом свой, и готовы окружить его по улице плакальщицы; –
ECCL|12|6|доколе не порвалась серебряная цепочка, и не разорвалась золотая повязка, и не разбился кувшин у источника, и не обрушилось колесо над колодезем.
ECCL|12|7|И возвратится прах в землю, чем он и был; а дух возвратился к Богу, Который дал его.
ECCL|12|8|Суета сует, сказал Екклесиаст, все – суета!
ECCL|12|9|Кроме того, что Екклесиаст был мудр, он учил еще народ знанию. Он [все] испытывал, исследовал, [и] составил много притчей.
ECCL|12|10|Старался Екклесиаст приискивать изящные изречения, и слова истины написаны [им] верно.
ECCL|12|11|Слова мудрых – как иглы и как вбитые гвозди, и составители их – от единого пастыря.
ECCL|12|12|А что сверх всего этого, сын мой, того берегись: составлять много книг – конца не будет, и много читать – утомительно для тела.
ECCL|12|13|Выслушаем сущность всего: бойся Бога и заповеди Его соблюдай, потому что в этом все для человека;
ECCL|12|14|ибо всякое дело Бог приведет на суд, и все тайное, хорошо ли оно, или худо.
