ISA|1|1|當 烏西雅 、 約坦 、 亞哈斯 、 希西家 作 猶大 王的時候， 亞摩斯 的兒子 以賽亞 見異象，論到 猶大 和 耶路撒冷 。
ISA|1|2|天哪，要聽！地啊，側耳而聽！ 因為耶和華說： 「我養育兒女，將他們養大， 他們竟悖逆我。
ISA|1|3|牛認識主人， 驢認識主人的槽； 以色列 卻不認識， 我的民卻不明白。」
ISA|1|4|禍哉！犯罪的國民， 擔著罪孽的百姓， 行惡的族類， 敗壞的兒女！ 他們離棄耶和華， 藐視 以色列 的聖者， 背向他，與他疏遠。
ISA|1|5|你們為甚麼屢次悖逆，繼續受責打呢？ 你們已經滿頭疼痛， 全心發昏；
ISA|1|6|從腳掌到頭頂， 沒有一處是完好的， 盡是創傷、瘀青，與流血的傷口， 未曾擠淨，未曾包紮， 也沒有用膏滋潤。
ISA|1|7|你們的土地荒蕪， 城鎮被火燒燬； 你們的田地在你們眼前被陌生人侵吞， 既被陌生人傾覆，就成為荒蕪 。
ISA|1|8|僅存的 錫安 ， 好似葡萄園的草棚， 如瓜田中的茅屋， 又如被圍困的城。
ISA|1|9|若不是萬軍之耶和華為我們留下一些倖存者， 我們早已變成 所多瑪 ，像 蛾摩拉 一樣了。
ISA|1|10|所多瑪 的官長啊， 你們要聽耶和華的言語！ 蛾摩拉 的百姓啊， 要側耳聽我們上帝的教誨！
ISA|1|11|耶和華說： 「你們許多的祭物於我何益呢？ 公綿羊的燔祭和肥畜的油脂， 我已經膩煩了； 公牛、羔羊、公山羊的血， 我都不喜悅。
ISA|1|12|「你們來朝見我， 誰向你們的手要求這些， 使你們踐踏我的院宇呢？
ISA|1|13|不要再獻無謂的供物了， 香是我所憎惡的。 我不能容忍行惡又守嚴肅會： 初一、安息日和召集的大會。
ISA|1|14|你們的初一和節期，我心裏恨惡， 它們成了我的重擔， 擔當這些，令我厭煩。
ISA|1|15|你們舉手禱告，我必遮眼不看， 就算你們多多祈禱，我也不聽； 你們的手沾滿了血。
ISA|1|16|你們要洗滌、自潔， 從我眼前除掉惡行； 要停止作惡，
ISA|1|17|學習行善， 尋求公平， 幫助受欺壓的 ， 替孤兒伸冤， 為寡婦辯護。」
ISA|1|18|耶和華說： 「來吧，我們彼此辯論。 你們的罪雖像硃紅，必變成雪白； 雖紅如丹顏，必白如羊毛。
ISA|1|19|你們若甘心聽從， 必吃地上的美物；
ISA|1|20|若不聽從，反倒悖逆， 必被刀劍吞滅； 這是耶和華親口說的。」
ISA|1|21|忠信的城竟然變為妓女！ 從前充滿了公平， 公義居在其中， 現今卻有兇手居住。
ISA|1|22|你的銀子變為渣滓， 你的酒用水沖淡。
ISA|1|23|你的官長悖逆， 與盜賊為伍， 全都喜愛賄賂， 追求贓物； 他們不為孤兒伸冤， 寡婦的案件也呈不到他們面前。
ISA|1|24|因此，主－萬軍之耶和華、 以色列 的大能者說： 「唉！我要向我的對頭雪恨， 向我的敵人報仇。
ISA|1|25|我必反手對付你， 如鹼煉淨你的渣滓， 除盡你的雜質。
ISA|1|26|我必回復你的審判官，像起初一樣， 回復你的謀士，如起先一般。 然後，你必稱為公義之城， 忠信之邑。」
ISA|1|27|錫安 必因公平得蒙救贖， 其中歸正的人必因公義得蒙救贖。
ISA|1|28|但悖逆的和犯罪的必一同敗亡， 離棄耶和華的必致消滅。
ISA|1|29|那等人必因所喜愛的聖樹抱愧； 你們必因所選擇的園子 蒙羞，
ISA|1|30|因為你們必如葉子枯乾的橡樹， 如無水的園子。
ISA|1|31|有權勢的必如麻線， 他的作為好像火花， 都要一同焚燒，無人撲滅。
ISA|2|1|亞摩斯 的兒子 以賽亞 所見，有關 猶大 和 耶路撒冷 的事。
ISA|2|2|末後的日子，耶和華殿的山必堅立， 超乎諸山，高舉過於萬嶺； 萬國都要流歸這山。
ISA|2|3|必有許多民族前往，說： 「來吧，我們登耶和華的山， 到 雅各 上帝的殿。 他必將他的道教導我們， 我們也要行他的路。」 因為教誨必出於 錫安 ， 耶和華的言語必出於 耶路撒冷 。
ISA|2|4|他必在萬國中施行審判， 為許多民族斷定是非。 他們要將刀打成犁頭， 把槍打成鐮刀； 這國不舉刀攻擊那國， 他們也不再學習戰事。
ISA|2|5|雅各 家啊， 來吧！讓我們在耶和華的光明中行走。
ISA|2|6|你離棄了你的百姓 雅各 家， 因為他們充滿了東方的習俗 ， 又像 非利士 人一樣觀星象， 並與外邦人擊掌。
ISA|2|7|他們的國滿了金銀， 財寶也無窮； 他們的地滿了馬匹， 戰車也無數。
ISA|2|8|他們的地滿了偶像； 他們跪拜自己手所造的， 就是自己手指所做的。
ISA|2|9|有人屈膝， 有人下跪； 所以，不要饒恕他們。
ISA|2|10|當進入磐石，藏在土中， 躲避耶和華的驚嚇和他威嚴的榮光。
ISA|2|11|到那日，眼目高傲的必降卑， 狂妄的人必屈膝； 惟獨耶和華被尊崇。
ISA|2|12|因萬軍之耶和華的一個日子 要臨到所有驕傲狂妄的， 臨到一切自高的， 使他們降為卑；
ISA|2|13|臨到 黎巴嫩 高大的香柏樹、 巴珊 的橡樹，
ISA|2|14|臨到一切高山、 一切峻嶺，
ISA|2|15|臨到一切碉堡、 一切堅固的城牆，
ISA|2|16|臨到 他施 一切的船隻、 一切華麗的船艇。
ISA|2|17|人的驕傲必屈膝， 人的狂妄必降卑； 在那日，惟獨耶和華被尊崇，
ISA|2|18|偶像必全然廢棄。
ISA|2|19|耶和華興起使地大震動的時候， 人就進入石洞和土穴裏， 躲避耶和華的驚嚇和他威嚴的榮光。
ISA|2|20|到那日，人必將造來敬拜的金偶像、銀偶像 拋給田鼠和蝙蝠。
ISA|2|21|耶和華興起使地大震動的時候， 人就進入磐縫和巖隙裏， 躲避耶和華的驚嚇和他威嚴的榮光。
ISA|2|22|你們不要倚靠世人， 他只不過鼻孔裏有氣息， 算得了甚麼呢？
ISA|3|1|看哪，主－萬軍之耶和華要從 耶路撒冷 和 猶大 除掉眾人所倚靠的，所仰賴的， 就是所倚靠的糧，所仰賴的水；
ISA|3|2|除掉勇士和戰士， 審判官和先知， 占卜的和長老，
ISA|3|3|除掉五十夫長和顯要、 謀士和巧匠， 以及擅長法術的人。
ISA|3|4|我必使孩童作他們的領袖， 幼兒管轄他們。
ISA|3|5|百姓要彼此欺壓， 各人欺壓鄰舍； 青年要侮慢老人， 卑賤的要侮慢尊貴的。
ISA|3|6|人在父家拉住自己的兄弟： 「你有外衣，來作我們的官長， 讓這些敗壞的事歸於你的手下吧！」
ISA|3|7|那時，他必揚聲說： 「我不作醫治你們的人； 我家裏沒有糧食，也沒有衣服， 你們不可立我作百姓的官長。」
ISA|3|8|耶路撒冷 敗落， 猶大 傾倒； 因為他們的舌頭和行為與耶和華相悖， 無視於他榮光的眼目。
ISA|3|9|他們的臉色證明自己不正， 他們述說自己像 所多瑪 一樣的罪惡，毫不隱瞞。 他們有禍了！因為作惡自害。
ISA|3|10|你們要對義人說，他是有福的， 因為他必吃自己行為所結的果實。
ISA|3|11|惡人有禍了！他必遭災難！ 因為他要按自己手所做的受報應。
ISA|3|12|至於我的百姓， 統治者剝削你們， 放高利貸的人管轄你們 。 我的百姓啊，引導你的使你走錯， 並毀壞你所行的道路。
ISA|3|13|耶和華興起訴訟， 站著審判萬民。
ISA|3|14|耶和華必審問他國中的長老和領袖： 「你們，你們摧毀葡萄園， 搶奪困苦人，囤積在你們家中。
ISA|3|15|你們為何壓碎我的百姓， 碾磨困苦人的臉呢？」 這是萬軍之主耶和華說的。
ISA|3|16|耶和華說： 因為 錫安 狂傲， 行走挺項，賣弄眼目， 俏步徐行，腳下玎璫，
ISA|3|17|主必使 錫安 頭頂長瘡， 耶和華又暴露其下體。
ISA|3|18|到那日，主必除掉華美的足飾、額帶、月牙圈、
ISA|3|19|耳環、手鐲、面紗、
ISA|3|20|頭巾、足鏈、華帶、香盒、符囊、
ISA|3|21|戒指、鼻環、
ISA|3|22|禮服、外套、披肩、皮包、
ISA|3|23|手鏡、細麻衣、頭飾、紗巾。
ISA|3|24|必有腐爛代替馨香， 繩子代替腰帶， 光禿代替美髮， 麻衣繫腰代替華服， 烙痕代替美貌。
ISA|3|25|你的男丁必倒在刀下， 你的勇士必死在陣上。
ISA|3|26|錫安 的城門必悲傷、哀號； 它必荒涼，坐在地上。
ISA|4|1|在那日，七個女人必拉住一個男人，說：「我們吃自己的食物，穿自己的衣服，但求你允許我們歸你名下，除掉我們的羞恥。」
ISA|4|2|在那日，耶和華的苗必華美尊榮，地的出產必成為倖存的 以色列 民的驕傲和光榮。
ISA|4|3|主以公平的靈和焚燒的靈洗淨 錫安 居民 的污穢，又除淨在 耶路撒冷 流人血的罪。那時，剩在 錫安 、留在 耶路撒冷 的，就是一切住 耶路撒冷 、在生命冊上記名的，必稱為聖。
ISA|4|4|
ISA|4|5|耶和華必在整座 錫安山 ，在會眾之上，白天造雲，黑夜發出煙和火焰的光，因為在一切榮耀之上必有華蓋；
ISA|4|6|這要作為棚子，白天可以遮蔭避暑，暴風雨侵襲時，可作藏身處和避難所。
ISA|5|1|我要為我親愛的唱歌， 我所愛的、他的葡萄園之歌。 我親愛的有葡萄園 在肥沃的山岡上。
ISA|5|2|他刨挖園子，清除石頭， 栽種上等的葡萄樹， 在園中蓋了一座樓， 又鑿出酒池； 指望它結葡萄， 反倒結了野葡萄。
ISA|5|3|耶路撒冷 的居民和 猶大 人哪， 現在，請你們在我與我的葡萄園之間斷定是非。
ISA|5|4|我為我葡萄園所做的之外， 還有甚麼可做的呢？ 我指望它結葡萄， 怎麼倒結了野葡萄呢？
ISA|5|5|現在我告訴你們， 我要向我的葡萄園怎麼做。 我必撤去籬笆，使它被燒燬； 拆毀圍牆，使它被踐踏。
ISA|5|6|我必使它荒廢，不再修剪， 不再鋤草，任荊棘蒺藜生長； 我也必吩咐密雲， 不再降雨在其上。
ISA|5|7|萬軍之耶和華的葡萄園就是 以色列 家； 他所喜愛的樹就是 猶大 人。 他指望公平， 看哪，卻有流血； 指望公義， 看哪，卻有冤聲。
ISA|5|8|禍哉！你們以房接房， 以地連地， 以致不留餘地， 只顧自己獨居境內。
ISA|5|9|我耳聞萬軍之耶和華說： 「許多房屋必然荒廢； 宏偉華麗，無人居住。
ISA|5|10|十畝 的葡萄園只釀出一罷特的酒， 一賀梅珥的穀種只結一伊法糧食。」
ISA|5|11|禍哉！那些清晨早起，追尋烈酒， 因酒狂熱，流連到深夜的人，
ISA|5|12|他們在宴席上 彈琴，鼓瑟，擊鼓，吹笛，飲酒， 卻不留意耶和華的作為， 也不留心他手所做的。
ISA|5|13|所以，我的百姓因無知就被擄去； 尊貴的人甚是飢餓， 平民也極其乾渴。
ISA|5|14|因此，陰間胃口 大開， 張開無限量的口； 令 耶路撒冷 的貴族與平民、狂歡的與作樂的人 都掉落其中。
ISA|5|15|人為之屈膝， 人就降為卑； 高傲的眼目也降為卑。
ISA|5|16|惟有萬軍之耶和華因公平顯為崇高， 神聖的上帝因公義顯為聖。
ISA|5|17|羔羊必來吃草，如同在自己的草場； 在富有人的廢墟，流浪的牲畜也來吃 。
ISA|5|18|禍哉！那些以虛假的繩子牽引罪孽， 以套車的繩索緊拉罪惡的人。
ISA|5|19|他們說： 「任 以色列 的聖者急速前行，快快成就他的作為， 好讓我們看看； 任他的籌算臨近成就， 好使我們知道。」
ISA|5|20|禍哉！那些稱惡為善，稱善為惡， 以暗為光，以光為暗， 以苦為甜，以甜為苦的人。
ISA|5|21|禍哉！那些在自己眼中有智慧， 在自己面前有通達的人。
ISA|5|22|禍哉！那些以飲酒稱雄， 以調烈酒稱霸的人。
ISA|5|23|他們因受賄賂，就稱惡人為義， 將義人的義奪去。
ISA|5|24|火苗怎樣吞滅碎秸， 乾草怎樣落在火焰之中， 照樣，他們的根必然腐朽， 他們的花像灰塵揚起； 因為他們厭棄萬軍之耶和華的教誨， 藐視 以色列 聖者的言語。
ISA|5|25|因此，耶和華的怒氣向他的百姓發作。 他伸手攻擊他們，山嶺就震動； 他們的屍首在街市上好像糞土。 雖然如此，他的怒氣並未轉消， 他的手依然伸出。
ISA|5|26|他必豎立大旗，召集遠方的國民， 把他們從地極叫來。 看哪，他們必急速奔來，
ISA|5|27|其中沒有疲倦的，絆跌的； 沒有打盹的，睡覺的； 腰帶並不放鬆， 鞋帶也不拉斷。
ISA|5|28|他們的箭銳利， 弓也上了弦； 馬蹄如堅石， 車輪像旋風。
ISA|5|29|他們要吼叫，像母獅， 咆哮，像少壯獅子； 他們要咆哮，抓取獵物， 穩穩叼走，無人能救回。
ISA|5|30|那日，他們要向 以色列 人咆哮， 像海浪澎湃； 人若望地，看哪，只有黑暗與禍患， 光明因密雲而變黑暗。
ISA|6|1|當 烏西雅 王崩的那年，我看見主坐在高高的寶座上。他的衣裳下襬遮滿聖殿。
ISA|6|2|上有撒拉弗侍立，各有六個翅膀：兩個翅膀遮臉，兩個翅膀遮腳，兩個翅膀飛翔，
ISA|6|3|彼此呼喊說： 「聖哉！聖哉！聖哉！萬軍之耶和華； 他的榮光遍滿全地！」
ISA|6|4|因呼喊者的聲音，門檻的根基震動，殿裏充滿了煙雲。
ISA|6|5|那時我說：「禍哉！我滅亡了！因為我是嘴唇不潔的人，住在嘴唇不潔的民中，又因我親眼看見大君王－萬軍之耶和華。」
ISA|6|6|有一撒拉弗向我飛來，手裏拿著燒紅的炭，是用火鉗從壇上取下來的，
ISA|6|7|用炭沾我的口，說：「看哪，這炭沾了你的嘴唇，你的罪孽便除掉，你的罪惡就赦免了。」
ISA|6|8|我聽見主的聲音說：「我可以差遣誰呢？誰肯為我們去呢？」我說：「我在這裏，請差遣我！」
ISA|6|9|他說：「你去告訴這百姓說： 『你們聽了又聽，卻不明白； 看了又看，卻不曉得。』
ISA|6|10|要使這百姓心蒙油脂， 耳朵發沉， 眼睛昏花； 恐怕他們眼睛看見， 耳朵聽見， 心裏明白， 回轉過來，就得醫治。」
ISA|6|11|我就說：「主啊，這到幾時為止呢？」他說： 「直到城鎮荒涼，無人居住， 房屋空無一人，土地極其荒蕪；
ISA|6|12|耶和華將人遷到遠方， 國內被撇棄的土地很多。
ISA|6|13|國內剩下的人若還有十分之一， 也必被吞滅。 然而如同大樹與橡樹，雖被砍伐， 殘幹卻仍存留， 聖潔的苗裔是它的殘幹。」
ISA|7|1|烏西雅 的孫子， 約坦 的兒子， 猶大 王 亞哈斯 在位的時候， 亞蘭 王 利汛 和 利瑪利 的兒子 以色列 王 比加 上來攻打 耶路撒冷 ，卻不能攻取。
ISA|7|2|有人告訴 大衛 家說：「 亞蘭 與 以法蓮 已經結盟。」王的心和百姓的心就都顫動，好像林中的樹被風吹動一樣。
ISA|7|3|耶和華對 以賽亞 說：「你和你的兒子 施亞‧雅述 要出去，到 上池 的水溝盡頭，往漂布地的大路上，迎見 亞哈斯 ，
ISA|7|4|對他說：『你要謹慎，要鎮定，不要害怕，不要因 利汛 和 亞蘭 ，以及 利瑪利 的兒子這兩個冒煙火把的頭所發的烈怒而心裏膽怯。
ISA|7|5|因為 亞蘭 、 以法蓮 ，和 利瑪利 的兒子設惡謀要害你，說：
ISA|7|6|我們要上去攻擊 猶大 ，擾亂它，攻破它來歸我們，在其中立 他比勒 的兒子為王。
ISA|7|7|主耶和華如此說： 這事必站立不住， 也不得成就。
ISA|7|8|因為 亞蘭 的首都是 大馬士革 ， 大馬士革 的領袖是 利汛 ； 六十五年之內， 以法蓮 必然國破族亡，
ISA|7|9|以法蓮 的首都是 撒瑪利亞 ； 撒瑪利亞 的領袖是 利瑪利 的兒子。 你們若是不信， 必站立不穩。』」
ISA|7|10|耶和華又吩咐 亞哈斯 ：
ISA|7|11|「你向耶和華－你的上帝求一個預兆：在陰間的深淵，或往上的高處。」
ISA|7|12|但 亞哈斯 說：「我不求；我不試探耶和華。」
ISA|7|13|以賽亞 說：「聽啊， 大衛 家！你們使人厭煩豈算小事，還要使我的上帝厭煩嗎？
ISA|7|14|因此，主自己要給你們一個預兆，看哪，必有童女懷孕生子，給他起名叫 以馬內利 。
ISA|7|15|到他曉得棄惡擇善的時候，他必吃乳酪與蜂蜜。
ISA|7|16|因為在這孩子還不曉得棄惡擇善之先，你所憎惡的那兩個王的土地必被撇棄。
ISA|7|17|耶和華必使 亞述 王臨到你和你的百姓，並你的父家，自從 以法蓮 脫離 猶大 的時候，未曾有過這樣的日子。
ISA|7|18|「那時，耶和華要呼叫，召來 埃及 江河源頭的蒼蠅和 亞述 地的蜂；
ISA|7|19|牠們都必飛來，停在陡峭的谷中、巖石縫裏、一切荊棘叢中和片片草場上。
ISA|7|20|「那時，主必用 大河 外雇來的剃刀，就是 亞述 王，剃去你的頭髮和腳毛，並要剃淨你的鬍鬚。
ISA|7|21|「那時，每一個人要養活一頭母牛犢和兩隻母羊；
ISA|7|22|因為奶量充足，他就有乳酪可吃，國內剩餘的人也都能吃乳酪與蜂蜜。
ISA|7|23|「那時，凡種一千棵葡萄樹、價值一千銀子的地方，必長出荊棘和蒺藜。
ISA|7|24|人到那裏去，必帶弓箭，因為遍地長滿了荊棘和蒺藜。
ISA|7|25|所有鋤頭刨過的山地，你因懼怕荊棘和蒺藜，不敢到那裏去；只能作放牛之處，羊群踐踏之地。」
ISA|8|1|耶和華對我說：「你取一塊大板子，拿人的筆 ，寫上『瑪黑珥‧沙拉勒‧哈施‧罷斯』 。
ISA|8|2|我 要用可靠的證人， 烏利亞 祭司和 耶比利家 的兒子 撒迦利亞 為我作證。」
ISA|8|3|我親近女先知 ；她就懷孕生子，耶和華對我說：「給他起名叫 瑪黑珥‧沙拉勒‧哈施‧罷斯 ；
ISA|8|4|因為在這孩子還不曉得叫爸爸媽媽以前， 大馬士革 的財寶和 撒瑪利亞 的擄物必被 亞述 王掠奪一空。」
ISA|8|5|耶和華又吩咐我：
ISA|8|6|「這百姓既厭棄 西羅亞 緩流的水，喜歡 利汛 以及 利瑪利 的兒子，
ISA|8|7|因此，看哪，主必使 亞述 王和他的威勢如 大河 翻騰洶湧的水上漲，蓋過他們，必上漲超過一切水道，漲過兩岸，
ISA|8|8|必沖入 猶大 ，漲溢氾濫，直到頸項。他展開翅膀，遮蔽你的全地。 以馬內利 啊！」
ISA|8|9|萬民哪，任憑你們行惡 ，終必毀滅； 遠方的眾人哪，當側耳而聽！ 任憑你們束腰，終必毀滅； 你們束起腰來，終必毀滅。
ISA|8|10|任憑你們籌算甚麼，終必無效； 不管你們講定甚麼，總不成立； 因為上帝與我們同在。
ISA|8|11|耶和華以大能的手訓誡我不可行 這百姓所行的道，對我這樣說：
ISA|8|12|「這百姓說同謀背叛的，你們不要說同謀背叛。他們所怕的，你們不要怕，也不要畏懼；
ISA|8|13|但要尊萬軍之耶和華為聖，他才是你們所當怕的，所當畏懼的。
ISA|8|14|他必作為聖所，卻向 以色列 的兩家成為絆腳的石頭，使人跌倒的磐石；作 耶路撒冷 居民的羅網和圈套。
ISA|8|15|許多人在其上絆倒，他們跌倒，甚至跌傷，並且落入陷阱，被抓住了。」
ISA|8|16|你要捲起律法書，在我門徒中間封住教誨。
ISA|8|17|我要等候那轉臉不顧 雅各 家的耶和華，也要仰望他。
ISA|8|18|看哪，我與耶和華所賜給我的兒女成了 以色列 的預兆和奇蹟，這是從住在 錫安山 萬軍之耶和華來的。
ISA|8|19|有人對你們說：「當求問招魂的與行巫術的，他們唧唧喳喳，念念有詞。」然而，百姓不當求問自己的上帝嗎？豈可為活人求問死人呢？
ISA|8|20|當以教誨和律法書為準；人所說的若不與此相符，必沒有黎明。
ISA|8|21|他必經過這地，遇艱難，受飢餓；飢餓的時候，心中焦躁，咒罵自己的君王和上帝。他仰觀上天，
ISA|8|22|俯察下地，看哪，盡是艱難、黑暗和駭人的昏暗。他必被趕入幽暗中去。
ISA|9|1|但那受過痛苦的必不再見幽暗。 從前上帝使 西布倫 地和 拿弗他利 地被藐視，末後卻使這沿海的路， 約旦河 東，外邦人居住的 加利利 地得榮耀。
ISA|9|2|在黑暗中行走的百姓看見了大光； 住在死蔭之地的人有光照耀他們。
ISA|9|3|你使這國民眾多 ， 使他們喜樂大增； 他們在你面前歡喜， 好像收割時的歡喜， 又像人分戰利品那樣的快樂。
ISA|9|4|因為他們所負的重軛 和肩頭上的杖， 並欺壓者的棍， 你都已經折斷， 如同在 米甸 的日子一般。
ISA|9|5|戰士在戰亂中所穿的靴子， 以及那滾在血中的衣服， 都必當作柴火燃燒。
ISA|9|6|因有一嬰孩為我們而生； 有一子賜給我們。 政權必擔在他的肩頭上； 他名稱為「奇妙策士、全能的上帝、永在的父、和平的君」。
ISA|9|7|他的政權與平安必加增無窮。 他必在 大衛 的寶座上治理他的國， 以公平公義使國堅定穩固， 從今直到永遠。 萬軍之耶和華的熱心必成就這事。
ISA|9|8|主向 雅各 家發出言語， 主的話臨到 以色列 家。
ISA|9|9|眾百姓，就是 以法蓮 和 撒瑪利亞 的居民， 都將知道； 他們憑驕傲自大的心說：
ISA|9|10|「磚塊掉落了，我們要鑿石頭重建； 桑樹砍了，我們要改種香柏樹。」
ISA|9|11|因此，耶和華興起 利汛 的敵人 前來攻擊 以色列 ， 要激起它的仇敵，
ISA|9|12|東有 亞蘭 人，西有 非利士 人； 他們張口吞吃 以色列 。 雖然如此，耶和華的怒氣並未轉消； 他的手依然伸出。
ISA|9|13|這百姓還沒有歸向擊打他們的主， 也沒有尋求萬軍之耶和華。
ISA|9|14|耶和華在一日之間 從 以色列 中剪除了頭與尾－ 棕樹枝與蘆葦－
ISA|9|15|長老和顯要就是頭， 以謊言教人的先知就是尾。
ISA|9|16|因為引導這百姓的使他們走入迷途， 被引導的都必被吞滅。
ISA|9|17|所以，主不喜愛 他們的青年， 也不憐憫他們的孤兒和寡婦； 因為他們都是褻瀆的，行惡的， 並且各人的口都說愚妄的話。 雖然如此，耶和華的怒氣並未轉消； 他的手依然伸出。
ISA|9|18|邪惡如火焚燒， 吞滅荊棘和蒺藜， 在稠密的樹林中點燃， 成為煙柱，旋轉上騰。
ISA|9|19|因萬軍之耶和華的烈怒，地都燒遍了； 百姓成為柴火， 無人憐惜弟兄。
ISA|9|20|有人右邊搶奪，猶受飢餓； 左邊吞吃，仍不飽足， 各人吃自己膀臂上的肉。
ISA|9|21|瑪拿西 吞吃 以法蓮 ， 以法蓮 吞吃 瑪拿西 ， 他們又一同攻擊 猶大 。 雖然如此，耶和華的怒氣並未轉消； 他的手依然伸出。
ISA|10|1|禍哉！那些設立不義之律例的， 和記錄奸詐之判詞的，
ISA|10|2|為要扭曲貧寒人的案件， 奪去我民中困苦人的理， 以寡婦當作擄物， 以孤兒當作掠物。
ISA|10|3|到降罰的日子，災禍從遠方臨到， 那時，你們要怎麼辦呢？ 你們要向誰逃奔求救呢？ 你們的財寶要存放何處呢？
ISA|10|4|他們只得屈身在被擄的人之下， 仆倒在被殺的人中間 。 雖然如此，耶和華的怒氣並未轉消； 他的手依然伸出。
ISA|10|5|禍哉！ 亞述 ，我怒氣的棍！ 他們手中的杖是我的惱恨。
ISA|10|6|我要差遣他攻擊褻瀆的國， 吩咐他對付我所惱怒的民， 搶走擄物，奪取掠物， 將他們踐踏，如同街上的泥土一般。
ISA|10|7|然而，這並非他的意念， 他的心不是這樣打算； 他的心要摧毀， 要剪除不少的國家。
ISA|10|8|他說：「我的官長豈不都是君王嗎？
ISA|10|9|迦勒挪 豈不像 迦基米施 嗎？ 哈馬 豈不像 亞珥拔 嗎？ 撒瑪利亞 豈不像 大馬士革 嗎？
ISA|10|10|既然我的手已伸到了這些有偶像的國， 他們所雕刻的偶像 過於 耶路撒冷 和 撒瑪利亞 的偶像，
ISA|10|11|我豈不照樣待 耶路撒冷 和其中的偶像， 如同我待 撒瑪利亞 和其中的偶像嗎？」
ISA|10|12|主在 錫安山 和 耶路撒冷 成就他一切工作的時候，說：「我必懲罰 亞述 王自大的心和他高傲尊貴的眼目。」
ISA|10|13|因為他說： 「我所成就的事是靠我手的能力 和我的智慧， 因為我本有聰明。 我挪移列國的地界， 搶奪他們所積蓄的財寶， 並且像勇士，使坐寶座的降為卑。
ISA|10|14|我的手奪取列國的財寶， 好像人奪取鳥窩； 我得了全地， 好像人拾起被棄的鳥蛋； 沒有振動翅膀的， 沒有張嘴的，也沒有鳴叫的。」
ISA|10|15|斧豈可向用斧砍伐的自誇呢？ 鋸豈可向拉鋸的自大呢？ 這好比棍揮動那舉棍的， 好比杖舉起那不是木頭的人。
ISA|10|16|因此，主－萬軍之耶和華 必使 亞述 王的壯士變為瘦弱， 在他的榮華之下必有火點燃， 如同火在燃燒一般。
ISA|10|17|以色列 的光必變成火， 它的聖者必成為火焰； 一日之間，將 亞述 王的荊棘和蒺藜焚燒淨盡，
ISA|10|18|又毀滅樹林和田園的榮華， 連魂帶體，好像病重的人消逝 一樣。
ISA|10|19|他林中只剩下稀少的樹木， 連孩童也能寫其數目。
ISA|10|20|到那日， 以色列 所剩下的和 雅各 家所逃脫的，必不再倚靠那擊打他們的，卻要誠心仰賴耶和華－ 以色列 的聖者。
ISA|10|21|所剩下的，就是 雅各 家的餘民，必歸回全能的上帝。
ISA|10|22|以色列 啊，你的百姓雖多如海沙，惟有剩下的歸回。滅絕之事已成定局，公義必如水漲溢。
ISA|10|23|因為萬軍之主耶和華在全地必成就所定的滅絕之事。
ISA|10|24|所以，萬軍之主耶和華如此說：「住 錫安 我的百姓啊， 亞述 王雖然用棍擊打你，又如 埃及 舉杖攻擊你，你不要怕他。
ISA|10|25|因為還有一點點時候，我向你們發的憤怒就要結束，我的怒氣要使他們滅亡。
ISA|10|26|萬軍之耶和華要舉起鞭子來攻擊他，好像在 俄立 磐石那裏擊打 米甸 人一樣。他的杖向海伸出，他必把杖舉起，如在 埃及 一般。
ISA|10|27|到那日， 亞述 王的重擔必離開你的肩頭，他的軛必離開你的頸項；那軛必因肥壯而撐斷 。」
ISA|10|28|亞述 王來到 亞葉 ， 經過 米磯崙 ， 在 密抹 安放輜重。
ISA|10|29|他們過了隘口， 要在 迦巴 住宿。 拉瑪 戰兢， 掃羅 的 基比亞 逃命。
ISA|10|30|迦琳 哪，要高聲呼喊！ 注意聽， 萊煞 啊！ 困苦的 亞拿突 啊 ！
ISA|10|31|瑪得米那 躲避， 基柄 的居民逃遁。
ISA|10|32|當那日， 亞述 王要在 挪伯 停留， 揮手攻擊 錫安 的山， 就是 耶路撒冷 的山。
ISA|10|33|看哪，主－萬軍之耶和華 以猛撞削斷樹枝； 巨木必被砍下， 高大的樹必降為低。
ISA|10|34|稠密的樹林，他要用鐵器砍下， 黎巴嫩 必被大能者伐倒 。
ISA|11|1|從 耶西 的殘幹必長出嫩枝， 他的根所抽的枝子必結果實。
ISA|11|2|耶和華的靈必住在他身上， 就是智慧和聰明的靈， 謀略和能力的靈， 知識和敬畏耶和華的靈。
ISA|11|3|他必以敬畏耶和華為樂； 行審判不憑眼見， 斷是非也不憑耳聞；
ISA|11|4|卻要以公義審判貧寒人， 以正直判斷地上的困苦人， 以口中的棍擊打全地， 以嘴裏的氣殺戮惡人。
ISA|11|5|公義必當他的腰帶， 信實必作他脅下的帶子。
ISA|11|6|野狼必與小綿羊同住， 豹子與小山羊同臥； 少壯獅子、牛犢和肥畜同群 ； 孩童要牽引牠們。
ISA|11|7|牛必與熊同食， 牛犢與小熊同臥； 獅子與牛一樣吃草。
ISA|11|8|吃奶的嬰孩在虺蛇的洞口玩耍， 斷奶的幼兒必按手在毒蛇的穴上。
ISA|11|9|在我聖山各處， 牠們都不傷人，不害物； 因為認識耶和華的知識要遍滿全地， 好像水充滿海洋一般。
ISA|11|10|到那日， 耶西 的根立作萬民的大旗；列國的人必尋求他，他安歇之所大有榮耀。
ISA|11|11|當那日，主必再度伸手救回自己百姓中所剩餘的，就是在 亞述 、 埃及 、 巴特羅 、 古實 、 以攔 、 示拿 、 哈馬 ，並眾海島所剩下的。
ISA|11|12|他要向列國豎立大旗， 召集 以色列 被趕散的人， 又從地極四方聚集分散的 猶大 人。
ISA|11|13|以法蓮 的嫉妒必消散， 苦待 猶大 的也被剪除； 以法蓮 必不嫉妒 猶大 ， 猶大 也不苦待 以法蓮 。
ISA|11|14|他們要飛向西方， 撲在 非利士 人的肩頭上， 他們要一同擄掠東方人， 他們的手伸到 以東 和 摩押 ； 亞捫 人也必順服他們。
ISA|11|15|耶和華必使 埃及 的海灣全然毀壞 ， 他舉手在 大河 之上颳起了暴熱的風， 擊打它，使它分成七條溪流， 人穿鞋便可渡過。
ISA|11|16|必有一條大道， 為百姓中從 亞述 逃脫生還的餘民而開， 如當日為 以色列 從 埃及 上來一樣。
ISA|12|1|在那日，你要說： 「耶和華啊，我要稱謝你！ 因為你雖然向我發怒， 你的怒氣卻已轉消； 你又安慰了我。
ISA|12|2|「看哪！上帝是我的拯救； 我要倚靠他，並不懼怕。 因為主耶和華是我的力量， 是我的詩歌， 他也成了我的拯救。」
ISA|12|3|你們必從救恩的泉源歡然取水。
ISA|12|4|在那日，你們要說： 「當稱謝耶和華，求告他的名； 在萬民中傳揚他的作為， 宣告他的名已被尊崇。
ISA|12|5|「你們要向耶和華唱歌， 因他所做的十分宏偉； 但願這事遍傳全地。
ISA|12|6|錫安 的居民哪，當揚聲歡呼， 因為在你們當中的 以色列 聖者最為偉大。」
ISA|13|1|亞摩斯 的兒子 以賽亞 所見，有關 巴比倫 的默示。
ISA|13|2|你們要在荒涼的山上豎立大旗， 向他們揚聲， 揮手招呼他們進入貴族之門。
ISA|13|3|我吩咐我所分別為聖的人， 召喚我的勇士， 就是我那狂喜高傲的人， 為要執行我的怒氣。
ISA|13|4|聽啊，山間有喧鬧的聲音， 好像有許多百姓聚集， 聽啊，多國之民聚集鬧鬨的聲音； 這是萬軍之耶和華召集作戰的軍隊。
ISA|13|5|他們從遠方來， 從天邊來， 耶和華和他惱恨的兵器 要毀滅全地。
ISA|13|6|你們要哀號， 因為耶和華的日子臨近了！ 這日來到，好像毀滅從全能者來到。
ISA|13|7|因此，人的手都變軟弱， 人的心都必惶惶。
ISA|13|8|他們必驚恐， 悲痛和愁苦將他們抓住。 他們陣痛，好像臨產的婦人一樣， 彼此驚奇對看，臉如火焰。
ISA|13|9|看哪！耶和華的日子臨到， 必有殘忍、憤恨、烈怒， 使這地荒蕪， 除滅其中的罪人。
ISA|13|10|天上的星宿都不發光， 太陽一升起就變黑暗， 月亮也不放光。
ISA|13|11|我必因邪惡懲罰世界， 因罪孽懲罰惡人， 我要止息驕傲人的狂妄， 制伏殘暴者的傲慢。
ISA|13|12|我要使人比純金更少， 比 俄斐 的赤金還少。
ISA|13|13|我，萬軍之耶和華狂怒，就是發烈怒的日子， 要令天震動， 地必搖撼，離其本位。
ISA|13|14|人如被追趕的羚羊， 像無人聚集的羊群， 各自歸回本族， 逃到本地。
ISA|13|15|凡被追上的必被刺死， 凡被捉拿的必倒在刀下。
ISA|13|16|他們的嬰孩必在他們眼前被摔死， 他們的房屋被搶劫， 他們的妻子被污辱。
ISA|13|17|看哪，我必激起 瑪代 人攻擊他們， 瑪代 人並不看重銀子， 也不喜愛金子。
ISA|13|18|他們必用弓擊潰青年， 不憐憫婦人所生的； 眼也不顧惜孩子。
ISA|13|19|巴比倫 為列國的榮耀， 為 迦勒底 人所誇耀的華美， 必像上帝所傾覆的 所多瑪 、 蛾摩拉 一樣；
ISA|13|20|國中必永無人煙， 世世代代無人居住； 阿拉伯 人不在那裏支搭帳棚， 牧羊的人也不使羊群躺臥在那裏。
ISA|13|21|曠野的走獸躺臥在那裏， 咆哮的動物擠滿棲身之所； 鴕鳥住在那裏， 山羊鬼魔也在那裏跳舞。
ISA|13|22|土狼必在它的宮殿 呼號， 野狗在華美的殿裏吼叫。 巴比倫 的時辰臨近了， 它的日子必不長久。
ISA|14|1|耶和華要憐憫 雅各 ，再度揀選 以色列 ，將他們安頓在本地。寄居的必與他們聯合，加入 雅各 家。
ISA|14|2|外邦人要將他們帶回本地。 以色列 家必在耶和華的地上得外邦人為僕婢，也要擄掠先前擄掠他們的，轄制先前欺壓他們的。
ISA|14|3|當耶和華使你得享安息，脫離愁苦、煩惱，和被迫做苦工的日子，
ISA|14|4|你必唱這詩歌嘲諷 巴比倫 王說： 「欺壓人的竟然滅亡！ 他的兇暴 竟然止息！
ISA|14|5|耶和華折斷惡人的杖， 打斷統治者的權杖；
ISA|14|6|他們在憤怒中連連攻擊萬民， 在怒氣中轄制列國， 逼迫他們，毫不留情。
ISA|14|7|現在全地得安息，享平靜， 人都出聲歡呼。
ISA|14|8|松樹和 黎巴嫩 的香柏樹 都因你歡樂： 自從你仆倒， 再也無人上來砍伐我們。
ISA|14|9|下面的陰間因你震動， 迎接你的到來； 在世曾為領袖的陰魂為你驚動， 那曾為列國君王的，都從寶座起立。
ISA|14|10|他們都要發言，對你說： 『你也變為軟弱，像我們一樣嗎？ 你也成了我們的樣子嗎？』
ISA|14|11|你的威嚴和琴瑟的聲音都下到陰間。 你下面鋪的是蟲，上面蓋的是蛆。
ISA|14|12|「明亮之星，早晨之子啊， 你竟然從天墜落！ 你這攻敗列國的，竟然被砍倒在地上！
ISA|14|13|你心裏曾說： 『我要升到天上， 我要高舉我的寶座在上帝的眾星之上， 我要坐在會眾聚集的山上，在極北的地方。
ISA|14|14|我要升到高雲之上， 我要與至高者同等。』
ISA|14|15|然而，你必墜落陰間， 到地府極深之處。
ISA|14|16|凡看見你的都要定睛望你， 留意看你，說： 『就是這個人嗎？ 他使大地顫抖， 使列國震動，
ISA|14|17|使世界如同荒野， 使城鎮傾覆； 是他，不釋放被擄的人歸家。』
ISA|14|18|列國的君王各自在自己的墳墓中， 在尊榮裏長眠。
ISA|14|19|惟獨你被拋棄在你的墳墓之外， 有如被厭惡的枝子 ， 被許多用刀刺透殺死的人覆蓋著， 一同墜落地府的石頭那裏， 像被踐踏的屍首。
ISA|14|20|你不得與君王同葬， 因為你毀壞你的國，殺戮你的民。 「惡人的後裔永不留名。
ISA|14|21|為了祖先的罪孽， 要預備他子孫的屠宰場， 免得他們興起，奪得全地， 使城市遍滿地面。」
ISA|14|22|萬軍之耶和華說： 「我必起來攻擊他們， 將 巴比倫 的名號和剩餘的人， 連子帶孫一併剪除； 這是耶和華說的。
ISA|14|23|「我必使 巴比倫 為豪豬佔據， 成為泥沼之地； 我要用滅命的掃帚掃淨它； 這是萬軍之耶和華說的。」
ISA|14|24|萬軍之耶和華起誓說： 「我怎樣思想，必照樣成就； 我怎樣定意，必照樣堅立，
ISA|14|25|要在我的地上擊破 亞述 ， 在我的山上將它踐踏。 它的軛必離開受壓制的人， 它的重擔必離開他們的肩頭。」
ISA|14|26|這是向全地所定的旨意， 向萬國所伸出的手。
ISA|14|27|萬軍之耶和華既然定意，誰能阻撓呢？ 他的手已經伸出，誰能使它縮回呢？
ISA|14|28|亞哈斯 王崩的那年，有默示如下：
ISA|14|29|「全 非利士 啊， 不要因擊打你的杖折斷就喜樂。 因為蛇必生出毒蛇， 牠所生的是會飛的火蛇。
ISA|14|30|貧寒人的長子必有得吃； 貧窮人必安然躺臥。 我必以饑荒滅絕你的根， 牠 必殺盡你所剩餘的人。
ISA|14|31|門哪，哀號吧！ 城啊，呼喊吧！ 全 非利士 都熔化了！ 因為有煙從北方而來， 在它的行伍中沒有掉隊的。」
ISA|14|32|當如何回答外邦的使者呢？ 「耶和華建立了 錫安 ， 在其中他困苦的百姓必有倚靠。」
ISA|15|1|論 摩押 的默示。 一夜之間， 摩押 的 亞珥 變為荒廢， 歸於無有； 一夜之間， 摩押 的 基珥 變為荒廢， 歸於無有。
ISA|15|2|摩押 上到神廟和 底本 的丘壇去哭泣； 它因 尼波 和 米底巴 哀號， 各人頭上光禿，鬍鬚剃淨。
ISA|15|3|他們在街市上腰束麻布， 都在房頂和廣場上哀號， 淚流不停。
ISA|15|4|希實本 和 以利亞利 呼喊， 他們的聲音達到 雅雜 ， 所以 摩押 的士兵高聲喊叫， 他們的心戰兢。
ISA|15|5|我的心 為 摩押 哀號； 它的難民逃到 瑣珥 ， 逃到 伊基拉‧施利施亞 。 他們上 魯希坡 ，隨走隨哭， 在 何羅念 的路上，因毀滅發出哀聲。
ISA|15|6|寧林 的水乾涸， 青草枯乾，嫩草死光， 青綠之物，一無所有。
ISA|15|7|因此， 摩押 人所得的財物和積蓄 都要運過 柳樹河 。
ISA|15|8|哀聲遍傳 摩押 四境， 哀號的聲音達到 以基蓮 ， 哀號的聲音遠及 比珥‧以琳 。
ISA|15|9|底們 的水充滿了血， 然而我還要加添 底們 的災難， 讓獅子追上 摩押 的難民 和那地 剩餘的人。
ISA|16|1|你們當將 羔羊奉送給那地的掌權者， 從 西拉 往曠野，送到 錫安 的山。
ISA|16|2|摩押 的居民 來到 亞嫩 渡口， 如逃遁的飛鳥，被趕離鳥巢 。
ISA|16|3|求你賜謀略，行公平， 使你的影子在正午如黑夜， 掩護逃亡的人，不洩露逃難者的行蹤。
ISA|16|4|願我 摩押 逃亡的人 寄居在你那裏， 你作他們的避難所，躲避滅命者的面。 勒索的人消失， 毀滅的事止息， 欺壓者從國中除滅，
ISA|16|5|在 大衛 帳幕中必有寶座因慈愛堅立， 必有一位君王憑信實坐在其上， 施行審判，尋求公平，迅速行公義。
ISA|16|6|我們聽聞 摩押 的驕傲， 極其驕傲； 它狂妄、驕傲、自大， 它誇大的言詞都是空的。
ISA|16|7|因此， 摩押 人必為 摩押 哀號， 人人都要哀號。 你們要為 吉珥‧哈列設 的葡萄餅哀嘆， 極其憂傷。
ISA|16|8|因為 希實本 的田地 和 西比瑪 的葡萄樹都衰殘了， 列國的君主折斷它的枝幹， 這枝子曾長到 雅謝 ，延伸到曠野， 嫩枝向外伸出，直伸過海；
ISA|16|9|所以，我要為 西比瑪 的葡萄樹哀哭， 像 雅謝 人一樣哀哭。 希實本 、 以利亞利 啊， 我要以眼淚澆灌你， 你因夏天果子和收割的莊稼， 歡呼聲已經止息了。
ISA|16|10|田園中不再有歡喜快樂， 葡萄園裏必無人歌唱，無人歡呼， 在壓酒池中踹酒的不再踹酒了， 我使歡呼的聲音止息了 。
ISA|16|11|因此，我的心腸為 摩押 哀鳴如琴， 我的內心為 吉珥‧哈列設 哀哭。
ISA|16|12|當 摩押 人出現在丘壇，筋疲力盡時，雖然到自己的聖所祈禱，卻仍無濟於事。
ISA|16|13|這是耶和華曾論到 摩押 的話。
ISA|16|14|但現在，耶和華說：「三年之內，按照雇工年數的算法， 摩押 的榮華必變為羞辱，人口雖曾眾多，剩餘的又少又弱。」
ISA|17|1|論 大馬士革 的默示。 看哪， 大馬士革 不再為城市， 變為廢墟。
ISA|17|2|亞羅珥 的城鎮被撇棄 ， 將成為牧羊之處， 羊群在那裏躺臥， 無人使牠們驚嚇。
ISA|17|3|以法蓮 不再有堡壘， 大馬士革 失去其王國， 亞蘭 的百姓所剩無幾， 如 以色列 人的榮美消失一般； 這是萬軍之耶和華說的。
ISA|17|4|到那日， 雅各 的榮美必失色， 它肥胖的身軀漸漸消瘦；
ISA|17|5|像人收割成熟的禾稼， 用手臂割取麥穗， 又像人在 利乏音谷 拾取穗子；
ISA|17|6|其間所剩不多，好像人打橄欖樹， 在最高的樹梢上只剩兩、三顆橄欖， 在多結果子的旁枝上只剩四、五顆； 這是耶和華－ 以色列 的上帝說的。
ISA|17|7|當那日，人必仰望造他們的主，眼目看著 以色列 的聖者。
ISA|17|8|他們必不仰望自己手所築的祭壇，也不理會自己指頭所造的 亞舍拉 和香壇。
ISA|17|9|當那日，他們堅固的城必因 以色列 人的緣故，如同樹林中和山頂上所撇棄的地方 。這樣，地就荒蕪了。
ISA|17|10|因你忘記拯救你的上帝， 忘記那保護你的磐石； 所以，你雖栽上佳美的樹苗， 插上別樣的枝子，
ISA|17|11|栽種的日子，你使它生長， 栽種的早晨，你使它開花， 但在愁苦、極其傷痛的日子， 所收割的都歸無有。
ISA|17|12|唉！萬民鬧鬨，好像海浪澎湃， 列邦喧鬧，如同洪水滔滔，
ISA|17|13|列邦喧鬧，如同大水滔滔； 但上帝一斥責，他們就遠遠躲避， 他們被追趕，如同山上風前的糠秕， 又如暴風前的碎秸；
ISA|17|14|看哪，晚上有驚嚇，未到早晨它就消失無蹤。 這是擄掠我們之人的厄運，是搶奪我們之人的報應。
ISA|18|1|禍哉！ 古實河 的那一邊、翅膀刷刷作響之地，
ISA|18|2|差遣使者在水面上， 坐蒲草船過海。 你們這些疾行的使者， 要到高大光滑的民那裏去； 那民遠近都畏懼， 是強大好征服的國， 土地有河流穿過。
ISA|18|3|世上所有的居民，住在地上的人哪， 山上大旗豎起時，你們要看， 號角吹響時，你們要聽。
ISA|18|4|耶和華對我如此說： 「我要安靜，從我的居所觀看， 如同日光下閃爍的熱氣， 又如收割時 露水蒸發的雲霧。」
ISA|18|5|收割之前，花蕾先謝， 花成了將熟的葡萄； 他必用刀削去嫩枝， 砍掉蔓延的枝條，
ISA|18|6|一起丟給山間的鷙鳥和地上的野獸； 鷙鳥要在其上避暑， 地上一切的野獸都在那裏過冬。
ISA|18|7|到那時，這高大光滑的民， 遠近都畏懼的民、 強大好征服之國、 土地有河流穿過； 他們必被當作 禮物獻給萬軍之耶和華， 獻到 錫安山 － 萬軍之耶和華立他名的地方。
ISA|19|1|論 埃及 的默示。 看哪，耶和華乘駕快雲， 臨到 埃及 ； 埃及 的偶像在他面前戰兢， 埃及 人的心在裏面消溶。
ISA|19|2|我要激起 埃及 人攻擊 埃及 人， 弟兄攻擊弟兄， 鄰舍攻擊鄰舍， 這城攻擊那城， 這國攻擊那國。
ISA|19|3|埃及 人的心神在裏面耗盡， 我要破壞他們的計謀。 他們必求問偶像和念咒的， 求問招魂的與行巫術的人。
ISA|19|4|我要將 埃及 人交在嚴厲的主人手中， 殘暴的君王必管轄他們； 這是主－萬軍之耶和華說的。
ISA|19|5|海水枯竭， 河流乾涸，
ISA|19|6|江河發臭， 埃及 的河水必然減少而枯乾。 蘆葦和蘆荻枯萎，
ISA|19|7|尼羅河 旁的植物 ，在 尼羅河 的沿岸， 並 尼羅河 旁所種的一切 全都枯焦，被風吹去，歸於無有。
ISA|19|8|打魚的哀哭， 所有在 尼羅河 釣魚的都必悲傷， 在水上撒網的也都衰殘。
ISA|19|9|以細緻的麻編織的必羞愧， 織布的必變蒼白 ；
ISA|19|10|織布的心情沮喪 ， 所有的傭工心都愁煩。
ISA|19|11|瑣安 的官長極其愚昧， 法老智慧的謀士籌劃愚謀； 你們怎敢對法老說： 「我是智慧人的子孫， 是古代國王的後裔？」
ISA|19|12|你的智慧人在哪裏？ 萬軍之耶和華向 埃及 所定的旨意， 他們既然知道，就讓他們告訴你吧！
ISA|19|13|瑣安 的官長愚昧， 挪弗 的官長受蒙蔽； 作 埃及 支派棟梁的， 帶領 埃及 走錯了路。
ISA|19|14|耶和華使歪曲的靈滲入 埃及 中間， 讓他們使 埃及 一切所做的都出差錯， 好像醉酒之人嘔吐時東倒西歪一樣。
ISA|19|15|在 埃及 ，無論是頭是尾， 棕樹枝與蘆葦，所做的事都不得成就。
ISA|19|16|到那日， 埃及 必像婦人一樣，因萬軍之耶和華揮手攻擊而戰兢懼怕。
ISA|19|17|猶大 地必使 埃及 驚恐，不論向誰提起，他都懼怕。這是因萬軍之耶和華向 埃及 所定的旨意。
ISA|19|18|當那日， 埃及 地必有五個城市的人說 迦南 的語言，又指著萬軍之耶和華起誓。有一城必稱為「太陽城」 。
ISA|19|19|在那日，在 埃及 地將有獻給耶和華的一座壇，邊界上必有為耶和華立的一根柱子。
ISA|19|20|這都要在 埃及 地為萬軍之耶和華作記號和證據。 埃及 人因受欺壓哀求耶和華，他就差遣一位救主作護衛者，拯救他們，
ISA|19|21|耶和華就被 埃及 所認識。在那日， 埃及 人要認識耶和華，獻牲祭和素祭敬拜他，並向耶和華許願還願。
ISA|19|22|耶和華必擊打 埃及 ，又擊打又醫治， 埃及 人就歸向耶和華。他必應允他們的禱告，醫治他們。
ISA|19|23|在那日，必有從 埃及 通往 亞述 的大道。 亞述 人要進入 埃及 ， 埃及 人也要進入 亞述 ； 埃及 人要與 亞述 人一同敬拜。
ISA|19|24|在那日， 以色列 將與 埃及 、 亞述 三國一起，使地上的人得福。
ISA|19|25|萬軍之耶和華必賜福給他們，說：「 埃及 －我的百姓， 亞述 －我手的工作， 以色列 －我的產業，都有福了！」
ISA|20|1|亞述 元帥 受 亞述 王 撒珥根 派遣往 亞實突 的那年，他攻打 亞實突 ，將城攻取。
ISA|20|2|那時，耶和華吩咐 亞摩斯 的兒子 以賽亞 說：「你去解掉你腰間的麻布，脫下你腳上的鞋。」 以賽亞 就這樣做，赤身赤腳行走。
ISA|20|3|耶和華說：「我僕人 以賽亞 怎樣赤身赤腳行走三年，作為關於 埃及 和 古實 的預兆奇蹟，
ISA|20|4|照樣， 亞述 王必擄去 埃及 人，掠去 古實 人，無論老少，都赤身赤腳，露出下體，使 埃及 蒙羞。
ISA|20|5|以色列 人必驚惶羞愧，因為他們仰望 古實 ，以 埃及 為榮。
ISA|20|6|「那時，沿海一帶的居民必說：『看哪，我們素來所仰望的，就是為躲避 亞述 王所逃往 求救的，不過如此！我們怎能逃脫呢？』」
ISA|21|1|論海邊曠野的默示。 它像 尼革夫 的旋風掃過， 從曠野，從可怕之地而來。
ISA|21|2|有悽慘的異象向我揭示： 「詭詐的在行詭詐，毀滅的在行毀滅。 以攔 哪，前進吧！ 瑪代 啊，圍攻吧！ 我使它一切的嘆息停止了。」
ISA|21|3|為此，我腰部滿是疼痛， 痛苦將我抓住， 好像臨產的婦人一樣的痛。 我疼痛甚至不能聽， 我驚惶甚至不能看 。
ISA|21|4|我心慌亂，驚恐威嚇我。 我所渴望的黃昏，反成為我的恐懼。
ISA|21|5|有人擺設筵席， 鋪上地毯，又吃又喝。 「官長啊，起來， 抹亮盾牌。」
ISA|21|6|主對我如此說： 「你去設立守望者， 讓他報告他所看見的。
ISA|21|7|他會看見一對一對騎著馬的軍隊， 又看見驢隊，駱駝隊， 他要留心聽，仔細地聽。」
ISA|21|8|他如獅子般吼叫 ： 「主啊，我白天常站在暸望樓， 徹夜立在我的暸望臺。」
ISA|21|9|看哪，有一對一對騎著馬的軍隊前來。 他就回應說：「 巴比倫 傾倒了！傾倒了！ 他把 巴比倫 神明的一切雕刻偶像都打碎在地上了。」
ISA|21|10|我被打的禾稼，我禾場上的穀物啊， 我從萬軍之耶和華－ 以色列 的上帝那裏所聽見的，都告訴你們了。
ISA|21|11|論 度瑪 的默示。 有人聲從 西珥 呼喊： 「守望的啊，夜裏如何？ 守望的啊，夜裏如何？」
ISA|21|12|守望者說： 「早晨來到，黑夜將臨。 你們若要問，問吧， 也可以回頭再來。」
ISA|21|13|論 阿拉伯 的默示。 底但 的旅行商隊啊， 你們在 阿拉伯 的樹林中住宿。
ISA|21|14|提瑪 地的居民哪， 提水來迎接口渴的人， 帶餅來迎接難民。
ISA|21|15|他們躲避刀劍和出了鞘的刀， 躲避上了弦的弓與戰爭的重災。
ISA|21|16|主對我這樣說：「一年之內，按照雇工年數的算法， 基達 一切的繁華必歸無有。
ISA|21|17|基達 人中強壯弓箭手剩下的數目甚為稀少，這是耶和華－ 以色列 的上帝說的。」
ISA|22|1|論異象谷的默示。 甚麼事使你們上去， 全都上到屋頂呢？
ISA|22|2|你這四處吶喊、大聲喧嘩的城、 歡樂的邑啊， 你被殺的並非被刀所殺， 也不是因打仗陣亡。
ISA|22|3|你所有的官長一同奔逃， 不用弓箭就被捆綁 ； 你們即使逃往遠方， 也要被找到，一同被捆綁。
ISA|22|4|因此我說： 「不要看我， 讓我痛哭吧！ 不要因我百姓 的毀滅竭力安慰我。」
ISA|22|5|因為這是萬軍之主耶和華使異象谷 混亂、踐踏、煩擾的日子； 城牆被攻破， 哀聲達到山上。
ISA|22|6|以攔 提著箭袋， 有戰車、士兵、騎兵； 吉珥 亮出盾牌，
ISA|22|7|你佳美的山谷遍佈戰車， 騎兵排列在城門前。
ISA|22|8|他除掉 猶大 的防禦。 那時，你指望森林庫裏的兵器。
ISA|22|9|你們看見 大衛城 缺口很多，就匯集 下池 的水；
ISA|22|10|你們數點 耶路撒冷 的房屋，拆毀房屋，用以修補城牆，
ISA|22|11|又在兩道城牆中間挖水池，用以盛舊池的水，卻不仰望成就這事的主，也不顧念從古時定這事的主。
ISA|22|12|當那日，萬軍之主耶和華使人哭泣哀號， 頭上光禿，身披麻布。
ISA|22|13|看哪，人卻歡喜快樂， 宰牛殺羊，吃肉喝酒： 「讓我們吃吃喝喝吧！因為明天要死了。」
ISA|22|14|萬軍之耶和華開啟我的耳朵： 「這罪孽直到你們死，斷不得赦免！」 這是萬軍之主耶和華說的。
ISA|22|15|萬軍之主耶和華如此說：「你到 舍伯那 宮廷總管那裏去，說：
ISA|22|16|『你在這裏憑甚麼？你在這裏靠誰？竟敢在這裏為自己鑿墳墓，在高處為自己鑿墳墓，在巖石中為自己挖安身之所！
ISA|22|17|你這偉大的人，看哪，耶和華必將你用力拋出，將你緊緊纏裹。
ISA|22|18|他必將你捲成一團，好像拋球一樣拋向寬闊之地。你這主人家的羞辱啊，你必死在那裏，你引以為榮的戰車也毀在那裏。
ISA|22|19|我要革除你的官職，你必從原位被逐 。』
ISA|22|20|「到那日，我要召 希勒家 的兒子─我的僕人 以利亞敬 來，
ISA|22|21|將你的外袍給他穿上，將你的腰帶給他繫緊，將你的政權交在他手中。他必作 耶路撒冷 居民和 猶大 家的父。
ISA|22|22|我要將 大衛 家的鑰匙放在他肩頭上。他開了，無人能關；他關了，無人能開。
ISA|22|23|我要使他立穩，像釘子釘在堅固的地方；他必成為他父家榮耀的寶座。
ISA|22|24|他父家所有的榮耀，連兒女帶子孫，有如杯碗、瓶罐的小器皿，都掛在他身上。
ISA|22|25|當那日，萬軍之耶和華說，釘在堅固處的釘子必挪移，被砍斷落地，掛在上面的各樣重擔都被切斷。這是耶和華說的。」
ISA|23|1|論 推羅 的默示。 哀號吧， 他施 的船隻！ 因為 推羅 已成廢墟，沒有房屋存留， 他們從 基提 地來的時候，得到這個消息 。
ISA|23|2|沿海的居民， 西頓 的商家啊， 當靜默無聲。 你差人航海 ，
ISA|23|3|在大水之上， 西曷河 的糧食、 尼羅河 的莊稼是 推羅 的進項， 它就成為列國的商埠。
ISA|23|4|西頓 ，你這海洋中的堡壘啊，應當羞愧， 因為大海說 ： 「我未經歷產痛，也沒有生產， 未曾養育男孩，也沒有撫養女孩。」
ISA|23|5|推羅 的風聲傳到 埃及 時， 他們為這風聲極其疼痛。
ISA|23|6|你們當渡到 他施 去， 哀號吧，沿海的居民！
ISA|23|7|這就是你們那古老歡樂的城市嗎？ 它的腳曾帶人到遠方居住。
ISA|23|8|誰定意 推羅 有這樣的遭遇呢？ 它本是賜冠冕的， 它的商家是王子， 生意人是世上尊貴的人。
ISA|23|9|這是萬軍之耶和華所定的， 為要貶抑一切榮耀的狂傲， 使地上一切尊貴的人被藐視。
ISA|23|10|他施 啊， 你要像 尼羅河 一樣在你的地氾濫， 不再有腰帶的束縛了。
ISA|23|11|耶和華已經向海伸手， 震動列國； 他出令對付 迦南 ， 要拆毀其中的堡壘。
ISA|23|12|他說：「受欺壓的少女 西頓 哪， 你必不再歡樂。 起來！渡到 基提 去， 就是在那裏也不得安歇。
ISA|23|13|看哪， 迦勒底 人之地，這國民如今已不復存在。 亞述 人使它 成為住曠野者的居所。他們建築自己的瞭望樓，拆毀它的宮殿，使它成為荒涼。
ISA|23|14|哀號吧， 他施 的船隻！ 因你們的堡壘已成廢墟。
ISA|23|15|到那時， 推羅 必被忘記七十年，就是一位君王的年數。七十年後， 推羅 的景況必如妓女之歌：
ISA|23|16|「你這被遺忘的妓女啊， 帶著琴周遊城內， 彈得美妙，唱許多歌， 好讓人記得你。」
ISA|23|17|七十年後，耶和華必巡視 推羅 ，使它再度獲利 ，與地面上的世界各國貿易 。
ISA|23|18|它的收益和獲利都要歸耶和華為聖，不再私自屯積存留；因為它的收益必歸給住在耶和華面前的人，使他們吃飽，穿華麗的衣服。
ISA|24|1|看哪，耶和華使地空虛，變為荒蕪， 地面扭曲，居民四散。
ISA|24|2|那時，百姓如何，祭司也如何； 僕人如何，主人也如何； 婢女如何，主母也如何； 買主如何，賣主也如何； 放債的如何，借貸的也如何； 債主如何，欠債的也如何。
ISA|24|3|地必全然空虛，盡都荒蕪， 因為這話是耶和華說的。
ISA|24|4|大地悲哀凋零， 世界敗落衰殘， 地上居高位的人也沒落了。
ISA|24|5|地被其上的居民所污穢， 因為他們犯了律法， 廢了律例，背了永約。
ISA|24|6|所以，詛咒吞滅大地， 住在其上的都有罪； 地上的居民被火焚燒， 剩下的人稀少。
ISA|24|7|新酒悲哀，葡萄樹凋殘， 心中歡樂的都嘆息。
ISA|24|8|擊鼓之樂停止， 狂歡者的喧嘩止住， 彈琴之樂也停止了。
ISA|24|9|人不再飲酒唱歌， 喝烈酒的，必以為苦。
ISA|24|10|荒涼的城拆毀了， 各家關閉，無法進入。
ISA|24|11|有人在街上嚷著要酒喝， 一切的喜樂變為昏暗， 地上的歡樂全都消失。
ISA|24|12|城裏盡是荒涼， 城門全都摧毀。
ISA|24|13|地上的萬民正像打過的橄欖樹， 又如葡萄釀酒以後再去摘取，所剩無幾。
ISA|24|14|他們要高聲歡呼， 從海那邊揚聲讚美耶和華的威嚴。
ISA|24|15|因此，你們要在日出之地榮耀耶和華， 在眾海島榮耀耶和華－ 以色列 上帝的名。
ISA|24|16|我們聽見從地極有人歌唱： 「榮耀歸於公義的那一位！」 我卻說：「我滅亡了！ 我滅亡了，我有禍了！ 詭詐的還在行詭詐， 詭詐的還在大行詭詐。」
ISA|24|17|地上的居民哪， 驚嚇、陷阱、羅網都臨到你；
ISA|24|18|躲過驚嚇之聲的墜入陷阱， 逃離陷阱的又被羅網纏住， 因為天上的窗戶都打開， 地的根基也震動。
ISA|24|19|地必全然破壞，盡都崩裂， 劇烈震動。
ISA|24|20|地要搖搖晃晃，好像醉酒的人， 又如小屋子搖來搖去； 罪過重壓其上， 它就塌陷，不能復起。
ISA|24|21|到那日，耶和華在天上必懲罰天上的軍隊， 在地上必懲罰地上的列王。
ISA|24|22|他們必被聚集， 像囚犯困在牢裏， 他們被關在監獄， 多日之後便受懲罰。
ISA|24|23|那時，月亮要蒙羞，太陽要慚愧， 因為萬軍之耶和華必在 錫安山 ， 在 耶路撒冷 作王， 在他眾長老面前彰顯榮耀。
ISA|25|1|耶和華啊，你是我的上帝， 我要尊崇你，稱頌你的名。 因為你以信實忠信 行遠古所定奇妙的事。
ISA|25|2|你使城市變為廢墟， 使堅固的城荒涼， 使外邦人的城堡不再為城， 永遠不再重建。
ISA|25|3|所以，強大的民必尊敬你， 殘暴之國的城必敬畏你。
ISA|25|4|因為你是貧寒人的保障， 貧窮人急難中的保障， 暴風雨之避難所， 炎熱地之陰涼處。 當殘暴者盛氣凌人的時候， 如暴風直吹牆壁，
ISA|25|5|如乾旱地的熱氣， 你要制止外邦人的喧嚷， 殘暴者的歌要停止， 好像熱氣因雲的陰影而消失。
ISA|25|6|在這山上，萬軍之耶和華必為萬民擺設宴席，有肥甘與美酒，就是滿有骨髓的肥甘與精釀的美酒。
ISA|25|7|在這山上，他必吞滅纏裹萬民的面紗和那遮蓋列國的遮蔽物。
ISA|25|8|他已吞滅死亡直到永遠。主耶和華必擦乾各人臉上的眼淚，在全地除去他百姓的羞辱；這是耶和華說的。
ISA|25|9|到那日，人必說：「看哪，這是我們的上帝，我們向來等候他，他必拯救我們。這是耶和華，我們向來等候他，我們必因他的救恩歡喜快樂。」
ISA|25|10|耶和華的手必按住這山， 摩押 人要被踐踏在他底下，好像乾草被踐踏在糞池 裏。
ISA|25|11|他們要在其中伸展雙手，好像游泳的人伸手游泳。他們的手雖靈巧，耶和華卻使他們的驕傲降為卑下。
ISA|25|12|他使你城牆上堅固的碉堡傾倒，夷為平地，化為塵土。
ISA|26|1|當那日，在 猶大 地，人必唱這歌： 「我們有堅固的城， 耶和華賜救恩為城牆，為城郭。
ISA|26|2|你們要敞開城門， 使守信的公義之民得以進入。
ISA|26|3|堅心倚賴你的，你必保守他十分平安， 因為他倚靠你。
ISA|26|4|你們當倚靠耶和華，直到永遠， 因為耶和華，耶和華是永遠的磐石。
ISA|26|5|他使居住高處的與高處的城市一同降為卑下， 將城拆毀，夷為平地，化為塵土，
ISA|26|6|使它被腳踐踏， 就是被困苦人和貧寒人的腳踐踏。」
ISA|26|7|義人的道是正直的， 正直的主啊，你修平義人的路。
ISA|26|8|耶和華啊，我們在你行審判的路上等候你 ， 我們心裏所渴慕的，就是你的名和你的稱號 。
ISA|26|9|夜間，我的心渴想你， 我裏面的靈切切尋求你。 因為你在地上行審判的時候， 世上的居民就學習公義。
ISA|26|10|惡人雖然領受恩惠， 仍未學到公義。 在正直之地，他行不義， 也不看耶和華的威嚴。
ISA|26|11|耶和華啊，你的手高舉，他們不觀看； 願他們觀看你為百姓發的熱心而羞愧， 願火吞滅你的敵人。
ISA|26|12|耶和華啊，你必賞賜我們平安， 因為我們所做的一切，都是你為我們成就的。
ISA|26|13|耶和華－我們的上帝啊， 在你以外曾有別的主管轄我們， 但我們惟獨稱揚你的名。
ISA|26|14|死去的不能再復活， 陰魂不能再興起； 你懲罰他們，使他們毀滅， 他們的名號 就全然消滅。
ISA|26|15|耶和華啊，你增添國民， 你增添國民，得了榮耀， 又拓展國土的疆界。
ISA|26|16|耶和華啊，他們在急難中尋求你。 你的管教臨到他們身上時， 他們傾吐低聲的禱告。
ISA|26|17|婦人懷孕，臨產疼痛， 在痛苦之中喊叫； 耶和華啊，我們在你面前也是如此。
ISA|26|18|我們曾懷孕，曾疼痛， 所生產的竟像風一樣， 並未帶給地上任何拯救； 世上也未曾有居民生下來 。
ISA|26|19|你的死人要復活， 我的屍首要起來。 睡在塵土裏的啊，要醒起歌唱！ 你的甘露好像晨曦 的甘露， 地要交出陰魂。
ISA|26|20|我的百姓啊，要進入內室， 關上你的門，躲避片刻， 等到憤怒過去。
ISA|26|21|因為，看哪，耶和華從他的居所出來， 要懲罰地上居民的罪孽。 地必露出其中的血， 不再掩蓋被殺的人。
ISA|27|1|到那日，耶和華必用他堅硬銳利的大刀懲罰 力威亞探 ，就是那爬得快的蛇，懲罰 力威亞探 ，就是那彎彎曲曲的蛇，並殺死海裏的大魚。
ISA|27|2|當那日，你們要唱這美好 葡萄園的歌：
ISA|27|3|「我－耶和華看守葡萄園，按時灌溉， 晝夜看守，免得有人損害。
ISA|27|4|我心中不存憤怒。 惟願在戰爭中我有荊棘和蒺藜， 我就起步攻擊他， 把他一同焚燒；
ISA|27|5|或者讓他緊靠我，以我為避難所， 與我和好， 與我和好。」
ISA|27|6|將來 雅各 要扎根， 以色列 要發芽開花， 果實遍滿地面。
ISA|27|7|耶和華擊打 以色列 ， 豈像擊打那些擊打他們的人嗎？ 以色列 被殺戮， 豈像其他人所遭遇的殺戮嗎？
ISA|27|8|你驅趕他們，放逐他們， 與他們相爭。 在颳東風的日子， 他以暴風趕逐他們。
ISA|27|9|所以， 雅各 的罪孽藉此得赦免， 除罪的效果盡在乎此； 他使祭壇的石頭變為粉碎的石灰， 使 亞舍拉 和香壇不再立起。
ISA|27|10|因為堅固的城變為荒涼， 成了被撇棄的居所，像曠野一樣； 牛犢在那裏吃草， 在那裏躺臥，吃盡其中的樹枝。
ISA|27|11|它的枝條一枯乾，就被折斷， 婦女用以點火燃燒。 因為這百姓蒙昧無知， 所以，造他們的必不憐憫他們， 造成他們的也不施恩給他們。
ISA|27|12|到那日， 以色列 人哪，耶和華必像人打樹拾果一般，從 大河 的支流，直到 埃及 的溪谷，將你們一一收集。
ISA|27|13|當那日，號角大響；在 亞述 地將亡的，與被趕散至 埃及 地的，都要前來，在 耶路撒冷 聖山上敬拜耶和華。
ISA|28|1|禍哉！ 以法蓮 酒徒高傲的冠冕， 其榮美竟如花凋殘； 他們在肥沃的山谷頂上， 被酒擊敗。
ISA|28|2|看哪，主有一位大能大力者， 如強烈的冰雹， 如毀滅的暴風雨， 如漲溢的洪水， 他必親手將他們摔落在地。
ISA|28|3|以法蓮 酒徒高傲的冠冕， 必被腳踐踏；
ISA|28|4|那如凋殘之花的榮美， 在肥沃的山谷頂上， 必如夏令前初熟的無花果， 讓看見的人注意， 摘到手裏，隨即吞吃。
ISA|28|5|到那日，萬軍之耶和華 必成為他餘民的榮冠華冕，
ISA|28|6|成為在位審判者的公平之靈， 和城門口制敵的力量。
ISA|28|7|這些人也因酒搖晃， 因烈酒東倒西歪。 祭司和先知因烈酒搖晃， 被酒所困， 因烈酒東倒西歪。 他們錯解默示， 審判時不分是非。
ISA|28|8|筵席上都滿了嘔吐的污穢， 沒有一處乾淨。
ISA|28|9|「他要將知識指教誰呢？ 要向誰闡明信息呢？ 是向那些剛斷奶的， 離開母親胸懷的嗎？
ISA|28|10|因為他咕噥咕噥，咕噥咕噥， 嘮嘮叨叨，嘮嘮叨叨， 這裏一點，那裏一點。」
ISA|28|11|耶和華要藉嘲弄的嘴唇和外邦人的舌頭， 向這百姓說話。
ISA|28|12|他曾對他們說： 「這是安歇之所， 你們要使疲乏的人得安歇， 這是歇息之處。」 他們卻不肯聽。
ISA|28|13|耶和華的話對他們而言是 「咕噥咕噥，咕噥咕噥， 嘮嘮叨叨， 嘮嘮叨叨， 這裏一點，那裏一點」； 以致他們往前行， 卻後仰跌倒，甚至跌傷， 落入陷阱，被抓住了。
ISA|28|14|因此，你們這些傲慢的人， 就是管轄住 耶路撒冷 這百姓的， 要聽耶和華的話。
ISA|28|15|你們曾說： 「我們已與死亡立約， 與陰間結盟， 不可擋的鞭子揮過時， 必不臨到我們； 因我們以謊言為避難所， 靠虛假來藏身」；
ISA|28|16|所以，主耶和華如此說： 「看哪，我在 錫安 放一塊石頭作為根基， 是衡量的石頭， 是寶貴的房角石，穩固的根基； 信靠他的人必不致驚恐。
ISA|28|17|我以公平為準繩， 以公義為鉛垂線； 冰雹必沖去謊言的避難所， 大水必漫過藏身之處。
ISA|28|18|你們與死亡所立的約必廢除， 與陰間所結的盟不得堅立； 不可擋的鞭子揮過時， 你們必被踐踏。
ISA|28|19|每逢它揮來，必將你們擄去； 每早晨它必揮過， 白晝黑夜都是如此。 明白這信息的都必驚恐。」
ISA|28|20|床榻短，人不能伸展； 被子窄，人無從裹身。
ISA|28|21|耶和華必興起，像在 毗拉心山 ， 他必發怒，如在 基遍谷 ； 為要做成他的工，就是非常的工， 成就他的事，就是奇異的事。
ISA|28|22|現在你們不可傲慢， 免得捆綁你們的繩索更結實， 因為我從萬軍之主耶和華那裏聽見， 在全地施行滅絕的事已定。
ISA|28|23|你們當側耳聽我的聲音， 留心聽我的言語。
ISA|28|24|那為撒種而耕地的 會不停地耕地，鬆土，耙地嗎？
ISA|28|25|他剷平了地面， 豈不就種小茴香， 播種大茴香， 按行列種小麥， 在定處種大麥， 在田邊種粗麥嗎？
ISA|28|26|他的上帝教導他， 指導他合宜的方法。
ISA|28|27|原來打小茴香，不用尖利的器具， 軋大茴香，也不是用車輪； 卻要用杖打小茴香， 用棍打大茴香。
ISA|28|28|穀要打， 但不能持續地搗， 用車輪和馬軋， 卻不軋碎它。
ISA|28|29|這也是出於萬軍之耶和華， 他的謀略奇妙， 他的智慧廣大。
ISA|29|1|禍哉！ 亞利伊勒 ， 亞利伊勒 ， 大衛 安營的城， 任憑你年復一年， 節期照常循環，
ISA|29|2|我卻要使 亞利伊勒 遭難； 它必悲傷哀號， 它對我是 亞利伊勒 。
ISA|29|3|我必四圍安營攻擊你， 築臺圍困你， 堆壘攻擊你。
ISA|29|4|你必敗落，從地裏說話， 你的言語細微出於塵埃。 你的聲音必像那招魂者的聲音出於地， 你的言語呢喃出於塵埃。
ISA|29|5|你那成群的陌生人 要像細塵， 暴民要像吹起的糠秕； 這事必頃刻之間忽然臨到。
ISA|29|6|萬軍之耶和華必使雷轟、地震、巨響、旋風、暴風， 並吞滅的火焰臨到它。
ISA|29|7|那時，攻擊 亞利伊勒 列國的軍隊， 與一切攻擊 亞利伊勒 和它城堡， 並帶給它患難的， 必如夢，如夜間的異象；
ISA|29|8|又像飢餓的人在夢中吃飯， 醒了仍覺飢腸轆轆； 或像口渴的人在夢中喝水， 醒了仍覺發昏，心裏想喝。 攻擊 錫安山 列國的軍隊也必如此。
ISA|29|9|你們等候驚奇吧！ 你們沉迷宴樂吧！ 他們醉了，卻非因酒； 東倒西歪，卻非因烈酒。
ISA|29|10|因為耶和華將沉睡的靈澆灌你們， 遮住你們的眼， 眼就是先知， 覆蓋你們的頭， 頭就是先見。
ISA|29|11|所有的默示，在你們看來都如封住的書卷，人將這書卷交給識字的人，說：「請念吧！」他說：「我不能念，因為它封住了。」
ISA|29|12|又將這書卷交給不識字的人，說：「請念吧！」他說：「我不識字。」
ISA|29|13|主說：「因這百姓以口親近我， 用嘴唇尊敬我， 心卻遠離我； 他們敬畏我， 不過是領受前人的命令。
ISA|29|14|所以，看哪，我要在這百姓中行奇妙的事， 就是奇妙又奇妙的事。 他們智慧人的智慧必然消滅， 聰明人的聰明必然消失。」
ISA|29|15|禍哉！那些向耶和華深藏謀略的， 他們在暗中行事，說： 「有誰看見我們呢？ 誰會注意我們呢？」
ISA|29|16|你們把事情顛倒了， 豈可看陶匠如陶土呢？ 受造物豈可論創造者說， 「他並沒有造我」？ 製成物豈可論製作者說， 「他根本不懂」？
ISA|29|17|黎巴嫩 變為田園， 田園看似森林， 不是只需要一些時間嗎？
ISA|29|18|那時，聾子必聽見這書上的話； 盲人的眼必從迷矇黑暗中看見。
ISA|29|19|困苦的人必因耶和華增添歡喜， 人間貧窮的必因 以色列 的聖者快樂。
ISA|29|20|因為殘暴的人歸於無有， 傲慢的人已經滅絕， 一切存心作惡的都被剪除。
ISA|29|21|他們憑一句話定一個人有罪， 為在城門口斷是非的設下羅網， 又用虛無的事屈枉義人。
ISA|29|22|所以，救贖 亞伯拉罕 的耶和華 論到 雅各 家時如此說： 「 雅各 必不再羞愧， 面容也不再變色。
ISA|29|23|當他的兒女看見 我的手在他們當中所成就的事情 ， 他們就必尊我的名為聖， 尊 雅各 的聖者為聖， 他們必敬畏 以色列 的上帝。
ISA|29|24|心中迷糊的必明白， 發怨言的必領受訓誨。」
ISA|30|1|耶和華說： 「禍哉！這悖逆的兒女。 他們同謀，卻不出於我， 結盟，卻不出於我的靈， 以致罪上加罪。
ISA|30|2|他們沒有尋求我的指示，就起身下 埃及 去， 要倚靠法老的庇護堅固自己， 並投在 埃及 的蔭下。
ISA|30|3|但法老的庇護反成為你們的羞辱； 你們投在 埃及 蔭下，反使你們慚愧。
ISA|30|4|他們的領袖已在 瑣安 ， 他們的使臣到了 哈內斯 。
ISA|30|5|他們必因那無益於他們的民蒙羞； 那民並非幫助，也非有益， 只帶來羞恥和凌辱。」
ISA|30|6|論 尼革夫 牲畜的默示。 他們將財物馱在驢背上， 將寶物馱在駱駝的背脊， 經過艱難困苦之地， 就是母獅、公獅、毒蛇、飛蛇之地， 往那無益於他們的民那裏去。
ISA|30|7|埃及 的幫助是徒然的， 因此，我稱它為「毫不中用的 拉哈伯 」 。
ISA|30|8|現在你要去， 在他們面前將這話刻在版上， 寫在書上， 以便流傳後世，直到永永遠遠 。
ISA|30|9|因為他們是悖逆的百姓、說謊的兒女， 是不肯聽從耶和華訓誨的兒女。
ISA|30|10|他們對先見說：「不要再看了」； 對先知說：「不要向我們預言正直的事； 要對我們說好聽的話， 預言虛幻的事。
ISA|30|11|要離開這道，偏離這路， 不要在我們面前再提說 以色列 的聖者。」
ISA|30|12|所以， 以色列 的聖者如此說： 「因你們藐視這話， 倚賴欺壓和詭詐，以此為可靠，
ISA|30|13|因此，這罪孽在你們身上， 好像高牆裏有凸起的裂縫， 頃刻之間忽然坍下來了；
ISA|30|14|它被砸碎，好像把陶匠的瓦器摔碎， 毫不顧惜， 甚至在碎塊中找不到一片 可用以從爐內取火，或從池中舀水。
ISA|30|15|主耶和華－ 以色列 的聖者如此說： 「你們得救在乎歸回安息， 得力在乎平靜安穩。」 你們卻是不肯，
ISA|30|16|你們說：「不然，我們要騎馬奔走」， 所以你們必然奔走。 你們又說：「我們要騎快馬」， 所以追趕你們的，也必飛快。
ISA|30|17|一人叱喝，令千人逃跑， 五人叱喝，你們都逃跑； 以致剩下的如山頂的旗杆， 如山岡上的大旗。
ISA|30|18|耶和華必然等候，要施恩給你們； 必然興起，好憐憫你們。 因為耶和華是公平的上帝； 凡等候他的都是有福的！
ISA|30|19|住在 錫安 、居於 耶路撒冷 的百姓啊，你必不再哭泣。主必因你哀求的聲音施恩給你，他聽見的時候就必應允你。
ISA|30|20|主雖然以艱難給你當餅，以困苦給你當水，你的教師卻不再隱藏，你的眼睛必看見你的教師。
ISA|30|21|你或向左或向右，必聽見後邊有聲音說：「這是正路，要行在其間。」
ISA|30|22|你要玷污那雕刻偶像所包的銀子和鑄造偶像所鍍的金子。你要拋棄它們，如拋棄污穢之物；對偶像說：「去吧！」
ISA|30|23|你撒種在地裏，主必降雨在其上，使地所出的糧食肥美豐盛。那時，你的牲畜必在遼闊的草場吃草。
ISA|30|24|耕地的牛和驢必吃加鹽的飼料，是用鏟子和杈子揚淨的。
ISA|30|25|在大行殺戮的日子，城樓倒塌的時候，高山峻嶺必有川河湧流。
ISA|30|26|當耶和華包紮他百姓的傷口，醫治他所擊打傷痕的日子，月光必像日光，日光必加七倍，像七日的光一樣。
ISA|30|27|看哪，耶和華的名從遠方來， 他的怒氣燒起，濃煙上騰。 他的嘴唇滿有憤恨， 他的舌頭像吞滅的火。
ISA|30|28|他的氣息如漲溢的河水，直漲到頸項， 要用毀滅的篩網篩淨列國， 並在眾民口中安放導錯方向的嚼環。
ISA|30|29|你們必唱歌，像守聖節的夜間一樣；並且心中喜樂，像人吹笛，來到耶和華的山，到 以色列 的磐石那裏。
ISA|30|30|耶和華必使人聽見他威嚴的聲音，又以極大的憤怒、吞滅的火焰、雷雨、暴風和像石塊的冰雹，使人看見他降罰的膀臂。
ISA|30|31|亞述 必因耶和華的聲音驚惶，耶和華必用杖擊打它。
ISA|30|32|耶和華必將定規要打 的杖加在它身上；每打一下，都必配合擊鼓彈琴的節奏。打仗時，耶和華必振臂與它交戰。
ISA|30|33|原來 陀斐特 早已預備好了，是為君王預備的；又深又寬，堆滿了火和木柴；耶和華的氣息猶如一股硫磺使它燃起。
ISA|31|1|禍哉！那些下 埃及 求幫助的， 他們仰賴馬匹，倚靠甚多的戰車， 並倚靠強壯的騎兵， 卻不仰望 以色列 的聖者， 也不求問耶和華。
ISA|31|2|其實，耶和華有智慧， 他降災禍， 並不撤回自己的話， 卻要興起攻擊作惡之家， 攻擊那幫助人作惡的。
ISA|31|3|埃及 人不過是人，並非上帝， 他們的馬不過是血肉，並不是靈。 耶和華一伸手， 那幫助人的必絆跌，受幫助的也必跌倒， 都一同滅亡。
ISA|31|4|耶和華對我如此說， 獅子和少壯獅子為獵物而咆哮， 許多牧人被召來攻擊牠， 牠總不因他們的聲音驚惶， 也不因他們的喧嚷退縮； 萬軍之耶和華也必如此 降臨在 錫安 的大小山岡上爭戰。
ISA|31|5|雀鳥盤旋護衛， 萬軍之耶和華也必照樣保護 耶路撒冷 ； 他必保護拯救， 必逾越而搭救。
ISA|31|6|以色列 人哪，要歸向你們嚴重悖逆的那一位！
ISA|31|7|到那日，你們各人要拋棄親手所造、陷自己於罪中的金偶像和銀偶像。
ISA|31|8|亞述 必倒在刀下，並非人的刀； 有刀要將它吞滅，並非人的刀。 它要逃避這刀， 它的年輕人必做苦工。
ISA|31|9|它的磐石必因驚嚇而消失， 它的領袖必因大旗驚惶； 這是那有火在 錫安 、 有爐在 耶路撒冷 的耶和華說的。
ISA|32|1|看哪，必有一位君王憑公義執政， 必有王子藉公平掌權。
ISA|32|2|必有一人如避風港， 如暴風雨的藏身處； 如乾旱地的溪流， 又如乾燥地巨石的陰影。
ISA|32|3|看的人眼睛不再昏花， 聽的人耳朵必留心聽。
ISA|32|4|性急的人懂得分辨， 口吃的人說話流暢。
ISA|32|5|愚頑人不再稱為君子， 流氓不再稱為紳士。
ISA|32|6|因為愚頑人必說愚妄的話， 他的心作惡 ， 行褻瀆的事， 傳播惡言攻擊耶和華， 使飢餓的人仍然飢餓， 口渴的人無水可喝。
ISA|32|7|流氓的手段邪惡， 他圖謀惡計， 用謊言毀滅困苦人； 貧窮人講求公理時， 他也是如此行。
ISA|32|8|君子卻圖謀高尚的事， 他必因高尚的事站立得穩。
ISA|32|9|安逸的婦女啊，起來聽我的聲音！ 無慮的女子啊，側耳聽我的言語！
ISA|32|10|無慮的女子啊，再過一年，你們必顫慄， 因為無葡萄可摘， 也無果實可收。
ISA|32|11|安逸的婦女啊，要戰兢； 無慮的女子啊，要顫慄， 要脫去衣服，赤著身體， 腰束麻布。
ISA|32|12|你們要為美好的田地 和多結果子的葡萄樹捶胸哀哭。
ISA|32|13|刺草和荊棘要長在我百姓的田地上， 長在歡樂城中一切快樂家園上。
ISA|32|14|宮殿必被撇下， 繁華的城必被拋棄， 堡壘和瞭望樓永為洞穴， 成為野驢的樂土， 羊群的草場。
ISA|32|15|等到聖靈從高處澆灌我們， 曠野將變為田園， 田園看似森林。
ISA|32|16|公平要居住在曠野， 公義要安歇在田園。
ISA|32|17|公義的果實是平安， 公義的效果是平靜和安穩，直到永遠。
ISA|32|18|我的百姓要住在平安的居所， 安穩的住處，寧靜的安歇之地。
ISA|32|19|雖有冰雹擊倒樹林， 城也夷為平地；
ISA|32|20|然而你們在水邊撒種， 牧放牛驢的有福了！
ISA|33|1|禍哉！你這未遭毀滅而毀滅人的人， 人未以詭詐待你而你以詭詐待人的人！ 等你行完了毀滅， 自己必被毀滅； 你行完了詭詐， 人必以詭詐待你。
ISA|33|2|耶和華啊，求你施恩給我們， 我們等候你。 求你每早晨作我們的膀臂， 遭難時作我們的拯救。
ISA|33|3|轟然之聲一發出，萬民就奔逃； 你一興起 ，列國就四散。
ISA|33|4|你們的擄物必被斂盡， 有如螞蚱斂盡禾稼； 人為擄物奔走，宛如蝗蟲蹦跳。
ISA|33|5|耶和華受尊崇，居高處， 使公平和公義充滿 錫安 。
ISA|33|6|他是你這世代安定的力量， 豐盛的救恩、 智慧和知識； 敬畏耶和華是 錫安 的至寶。
ISA|33|7|看哪，他們的英雄在外面哀號 ， 求和的使臣在痛哭。
ISA|33|8|大路荒涼，行人止息； 盟約撕毀，見證 被棄， 人也不受尊重。
ISA|33|9|大地悲哀衰殘， 黎巴嫩 羞愧且枯乾， 沙崙 好像曠野， 巴珊 和 迦密 必凋殘。
ISA|33|10|耶和華說： 「現在我要興起， 要高升， 要受尊崇。
ISA|33|11|你們懷的是糠秕，生的是碎秸； 你們的氣息如火吞滅自己。
ISA|33|12|萬民必像燒著的石灰， 又如斬斷的荊棘，在火裏燃燒。」
ISA|33|13|你們遠方的人，當聽我所做的事； 你們近處的人，當承認我的大能。
ISA|33|14|錫安 的罪人都懼怕， 戰兢抓住不敬虔的人。 我們中間有誰能與吞噬的火同住？ 我們中間有誰能與不滅的火共存呢？
ISA|33|15|那行事公義、說話正直、 憎惡欺壓所得之財、 搖手不受賄賂、 掩耳不聽流血的計謀、 閉眼不看邪惡之事的，
ISA|33|16|這人必居高處， 他的保障是磐石的堡壘， 必有糧食賜給他， 飲水也不致斷絕。
ISA|33|17|你必親眼看見君王的榮美， 看見遼闊之地。
ISA|33|18|你的心必回想那些恐怖的事： 「那數算的人在哪裏？ 秤重的人在哪裏？ 數點城樓的又在哪裏呢？」
ISA|33|19|你必不再看見那兇暴的民， 他們嘴唇說艱澀的言語，難以理解； 舌頭結巴，說無意義的話。
ISA|33|20|你要注視 錫安 ，我們守聖節的城！ 你必親眼看見 耶路撒冷 成為安靜的居所， 成為不挪移的帳幕， 橛子永不拔出， 繩索一根也不折斷。
ISA|33|21|在那裏，威嚴的耶和華對我們是寬闊的江河， 其中必沒有搖槳的小船來往， 也沒有巨大的船舶經過。
ISA|33|22|耶和華是審判我們的， 耶和華為我們設立律法； 耶和華是我們的君王， 他必拯救我們。
ISA|33|23|船上的繩索鬆開， 不能穩住桅杆， 也無法揚起船帆。 那時許多擄物被瓜分， 連瘸腿的也能奪走掠物。
ISA|33|24|城內的居民無人說：「我病了」； 城裏居住的百姓，罪孽都蒙赦免。
ISA|34|1|列國啊，要近前來聽！ 萬民哪，要側耳而聽！ 全地和其上所充滿的， 世界和其中所出的，都應當聽！
ISA|34|2|因為耶和華向列國發怒， 向他們的全軍發烈怒， 要將他們滅盡，任人殺戮。
ISA|34|3|被殺的人必被拋棄， 屍首臭氣上騰， 諸山為他們的血所融化。
ISA|34|4|天上萬象都要朽壞， 天被捲起，有如書卷， 其上的萬象盡都衰殘； 如葡萄樹的葉子凋落， 又如無花果樹枯萎一樣。
ISA|34|5|因為我的刀在天上將要顯現 ； 看哪，這刀臨到 以東 和我所詛咒的民， 要施行審判。
ISA|34|6|耶和華的刀沾滿了血， 是用油脂和羔羊、公山羊的血， 並公綿羊腎上的油脂滋潤的； 因為在 波斯拉 有祭物獻給耶和華， 在 以東 地有大屠殺。
ISA|34|7|野牛與他們一起倒下， 牛犢和壯牛也一同倒下。 他們的地被血染遍， 他們的塵土因油脂肥潤。
ISA|34|8|這是耶和華報仇之日， 為 錫安 伸冤的報應之年。
ISA|34|9|它的河水要變為柏油， 塵埃變為硫磺， 大地成為燃燒的柏油，
ISA|34|10|晝夜總不熄滅， 它的煙永遠上騰， 必世世代代成為荒廢， 永永遠遠無人經過。
ISA|34|11|鵜鶘、豪豬要得它為業， 貓頭鷹、烏鴉要住在其間。 耶和華必將空虛的準繩、 混沌的石垂線，拉在 以東 之上。
ISA|34|12|人必宣稱那裏沒有王國， 它的貴族和所有領袖都歸於無有。
ISA|34|13|以東 的宮殿要長出荊棘， 城堡要生長蒺藜和刺草； 成為野狗的住處， 鴕鳥的居所。
ISA|34|14|野獸要和土狼相遇， 山羊鬼魔要與同伴對唱， 莉莉絲 必在那裏棲身， 為自己尋找安歇之處。
ISA|34|15|箭頭蛇要在那裏做窩， 下蛋，孵蛋，並招聚幼蛇在其保護之下； 鷂鷹也與伴侶聚集在那裏。
ISA|34|16|你們要查考並誦讀耶和華的書； 這些現象必然存在， 沒有一樣動物缺少伴侶。 因為是他，藉著我的口 吩咐， 他的靈將牠們聚集。
ISA|34|17|他為牠們抽籤， 親手用準繩為牠們分地； 直到牠們永遠得地為業， 世世代代住在其間。
ISA|35|1|曠野和乾旱之地必然歡喜， 沙漠也必快樂； 又如玫瑰綻放，
ISA|35|2|朵朵繁茂， 其樂融融，而且歡呼。 黎巴嫩 的榮耀， 並 迦密 與 沙崙 的華美，必賜給它。 人要看見耶和華的榮耀， 看見我們上帝的榮美。
ISA|35|3|你們要使軟弱的手強壯， 使無力的膝蓋穩固；
ISA|35|4|對心裏焦急的人說： 「要剛強，不要懼怕。 看哪，你們的上帝要來施報， 要施行極大的報應， 他必來拯救你們。」
ISA|35|5|那時，盲人的眼必睜開， 聾子的耳必開通。
ISA|35|6|那時，瘸子必跳躍如鹿， 啞巴的舌頭必歡呼。 在曠野有水噴出， 在沙漠有江河湧流。
ISA|35|7|火熱之地要變為水池， 乾渴之地要變為泉源。 野狗躺臥休息之處 必長出青草、蘆葦和蒲草。
ISA|35|8|在那裏必有一條大道， 就是一條路 ，稱為聖路。 污穢的人不得經過， 是專為走路的人 預備的， 愚昧的人也不會迷路。
ISA|35|9|在那裏沒有獅子， 猛獸也不經過； 在那裏牠們未現蹤跡， 只有救贖的民在那裏行走。
ISA|35|10|耶和華救贖的民必歸回， 歌唱來到 錫安 ； 永遠的快樂必歸到他們頭上， 他們必得著歡喜快樂， 憂傷嘆息盡都逃避。
ISA|36|1|希西家 王十四年， 亞述 王 西拿基立 上來攻擊 猶大 的一切堅固的城，將城攻取。
ISA|36|2|亞述 王從 拉吉 差遣將軍 率領大軍前往 耶路撒冷 ，到 希西家 王那裏去。將軍站在 上池 的水溝旁，在往漂布地的大路上。
ISA|36|3|希勒家 的兒子 以利亞敬 宮廷總管、 舍伯那 書記和 亞薩 的兒子 約亞 史官，出來見他。
ISA|36|4|將軍對他們說：「你們去告訴 希西家 ，大王 亞述 王如此說：『你倚靠甚麼，讓你如此自信滿滿？
ISA|36|5|我說 ，你有打仗的計謀和能力，我看不過是空話。你到底倚靠誰，竟敢背叛我呢？
ISA|36|6|看哪，你所倚靠的 埃及 是那斷裂的葦杖，人若倚靠這杖，它就刺進他的手，穿透它。 埃及 王法老向所有倚靠他的人都是這樣。
ISA|36|7|你若對我說：我們倚靠耶和華－我們的上帝， 希西家 豈不是將上帝的丘壇和祭壇廢去，並且吩咐 猶大 和 耶路撒冷 的人說：你們只當在這一個壇前敬拜嗎？
ISA|36|8|現在你與我主 亞述 王打賭，我給你兩千匹馬，看你能否派得出騎士來騎牠們。
ISA|36|9|若不然，怎能使我主臣僕中最小的一個軍官轉臉而逃呢？你難道要倚靠 埃及 的戰車和騎兵嗎？
ISA|36|10|現在我上來攻擊毀滅這地，豈不是出於耶和華嗎？耶和華吩咐我說，你上去攻擊這地，毀滅它吧！』」
ISA|36|11|以利亞敬 、 舍伯那 、 約亞 對將軍說：「求你用 亞蘭 話對僕人說，因為我們聽得懂；不要用 猶大 話對我們說，免得傳到城牆上百姓的耳中。」
ISA|36|12|將軍說：「我主差遣我來，豈是單對你和你的主人說這些話嗎？不也是對這些坐在城牆上，要與你們一同吃自己糞、喝自己尿的人說的嗎？」
ISA|36|13|於是 亞述 將軍站著，用 猶大 話大聲喊著說：「你們當聽大王 亞述 王的話，
ISA|36|14|王如此說：『你們不要被 希西家 欺哄了，因他不能拯救你們。
ISA|36|15|不要聽憑 希西家 說服你們倚靠耶和華，他說，耶和華必要拯救我們，這城必不交在 亞述 王的手中。』
ISA|36|16|你們不要聽 希西家 的話！因 亞述 王如此說：『你們要與我講和，出來投降，各人就可以吃自己葡萄樹和無花果樹的果子，喝自己井裏的水，
ISA|36|17|等我來領你們到一個地方，與你們本地一樣，就是有五穀和新酒之地，有糧食和葡萄園之地。
ISA|36|18|恐怕 希西家 誤導你們說，耶和華必拯救我們。列國的神明有哪一個曾救它本國脫離 亞述 王的手呢？
ISA|36|19|哈馬 和 亞珥拔 的神明在哪裏呢？ 西法瓦音 的神明在哪裏呢？它們曾救 撒瑪利亞 脫離我的手嗎？
ISA|36|20|這些國的神明有誰曾救自己的國家脫離我的手呢？難道耶和華能救 耶路撒冷 脫離我的手嗎？』」
ISA|36|21|百姓靜默不言，一句不答，因為 希西家 王曾吩咐說：「不要回答他。」
ISA|36|22|當下 希勒家 的兒子 以利亞敬 宮廷總管、 舍伯那 書記，和 亞薩 的兒子 約亞 史官都撕裂衣服，來到 希西家 那裏，將 亞述 將軍的話告訴他。
ISA|37|1|希西家 王聽見了，就撕裂衣服，披上麻布，進了耶和華的殿。
ISA|37|2|他差遣 以利亞敬 宮廷總管和 舍伯那 書記，並祭司中年長的，都披上麻布，到 亞摩斯 的兒子 以賽亞 先知那裏去。
ISA|37|3|他們對他說：「 希西家 如此說：『今日是急難、懲罰、凌辱的日子，就如嬰孩快要出生，卻沒有力氣生產。
ISA|37|4|或許耶和華－你的上帝聽見 亞述 將軍的話，就是他主人 亞述 王差他來辱罵永生上帝的話，耶和華－你的上帝就斥責所聽見的這些話。求你為倖存的餘民揚聲禱告。』」
ISA|37|5|希西家 王的臣僕就來到 以賽亞 那裏。
ISA|37|6|以賽亞 對他們說：「要對你們的主人這樣說，耶和華如此說：『你聽見 亞述 王的僕人褻瀆我的話，不要懼怕。
ISA|37|7|看哪，因為我必驚動他的心 ，他要聽見風聲就歸回本地，在那裏我必使他倒在刀下。』」
ISA|37|8|亞述 將軍聽見 亞述 王已拔營離開 拉吉 ，就啟程返回，正遇見 亞述 王去攻打 立拿 。
ISA|37|9|亞述 王聽見有人談論 古實 王 特哈加 說：「他出來要與你爭戰。」 亞述 王一聽見，就差使者去見 希西家 ，說：
ISA|37|10|「你們要對 猶大 王 希西家 如此說：『不要聽你所倚靠的上帝欺哄你說： 耶路撒冷 必不交在 亞述 王的手中。
ISA|37|11|看哪，你總聽說 亞述 諸王向列國所行的是盡行滅絕，難道你能倖免嗎？
ISA|37|12|我祖先所毀滅的，就是 歌散 、 哈蘭 、 利色 和 提‧拉撒 的 伊甸 人；這些國的神明何曾拯救他們呢？
ISA|37|13|哈馬 的王， 亞珥拔 的王， 西法瓦音城 的王， 希拿 和 以瓦 的王，都在哪裏呢？』」
ISA|37|14|希西家 從使者手裏接過書信，看完了，就上耶和華的殿，在耶和華面前展開書信。
ISA|37|15|希西家 向耶和華禱告說：
ISA|37|16|「坐在基路伯之上萬軍之耶和華－ 以色列 的上帝啊，你，惟有你是地上萬國的上帝，你創造了天和地。
ISA|37|17|耶和華啊，求你側耳而聽；耶和華啊，求你睜眼而看，聽 西拿基立 差遣使者辱罵永生上帝的一切話。
ISA|37|18|耶和華啊， 亞述 諸王果然使列國和列國之地變為荒蕪，
ISA|37|19|將列國的神明扔在火裏，因為它們不是神明，是人手所造的，是木頭、石頭，所以被滅絕了。
ISA|37|20|耶和華－我們的上帝啊，現在求你救我們脫離 亞述 王的手，使地上萬國都知道惟有你是耶和華。」
ISA|37|21|亞摩斯 的兒子 以賽亞 就差人去見 希西家 ，說：「耶和華－ 以色列 的上帝如此說，你因 亞述 王 西拿基立 的事向我祈求，
ISA|37|22|所以耶和華論他這樣說： 『少女 錫安 藐視你，嘲笑你； 耶路撒冷 向你搖頭。
ISA|37|23|「『你辱罵誰，褻瀆誰， 揚起聲來，高舉眼目攻擊誰呢？ 你攻擊的是 以色列 的聖者。
ISA|37|24|你藉臣僕辱罵主說： 我率領許多戰車登上高山， 到 黎巴嫩 的頂端； 我要砍伐其中高大的香柏樹 和上好的松樹。 我必上到極高之處， 進入茂盛的森林裏。
ISA|37|25|我已經挖井喝水 我必用腳掌踏乾 埃及 一切的河流。
ISA|37|26|「『你豈沒有聽見 我早先所定、古時所立、現今實現的事嗎？ 就是讓你去毀壞堅固的城鎮，使它們變為廢墟；
ISA|37|27|城裏居民的力量甚小， 他們驚惶羞愧； 像野草，像青菜， 如房頂上的草， 被東風颳散 。
ISA|37|28|「『你站起，你坐下，你出去，你進來， 你向我發烈怒，我都知道。
ISA|37|29|因你向我發烈怒， 你的狂傲上達我耳中， 我要用鉤子鉤住你的鼻子， 將嚼環放在你口裏， 使你從原路轉回去。』
ISA|37|30|「我賜給你的預兆：你們今年要吃野生的，明年也要吃自長的；後年，你們就要耕種收割，栽葡萄園，吃其中的果子。
ISA|37|31|猶大 家所逃脫剩餘的，仍要往下扎根，向上結果。
ISA|37|32|必有剩餘的民從 耶路撒冷 而出；有逃脫的人從 錫安山 而來。萬軍之耶和華的熱心必成就這事。
ISA|37|33|「所以耶和華論 亞述 王如此說：他必不得來到這城，也不在這裏射箭，不得拿盾牌到城前，也不能建土堆攻城。
ISA|37|34|他從哪條路來，必從那條路回去，必不得來到這城。這是耶和華說的。
ISA|37|35|因我為自己的緣故，又為我僕人 大衛 的緣故，必保護拯救這城。」
ISA|37|36|耶和華的使者出去，在 亞述 營中殺了十八萬五千人。清早有人起來，看哪，都是死屍。
ISA|37|37|亞述 王 西拿基立 就拔營回去，住在 尼尼微 。
ISA|37|38|一日，他在他的神明 尼斯洛 廟裏叩拜，他兒子 亞得米勒 和 沙利色 用刀殺了他，然後逃到 亞拉臘 地；他兒子 以撒．哈頓 接續他作王。
ISA|38|1|那些日子， 希西家 病得要死， 亞摩斯 的兒子 以賽亞 先知來見他，對他說：「耶和華如此說：『你當留遺囑給你的家，因為你必死，不能活了。』」
ISA|38|2|希西家 就轉臉朝牆，向耶和華禱告，
ISA|38|3|說：「耶和華啊，求你記念我在你面前怎樣存完全的心，按誠實行事，又做你眼中看為善的事。」 希西家 就痛哭。
ISA|38|4|耶和華的話臨到 以賽亞 說：
ISA|38|5|「你去告訴 希西家 說，耶和華－你祖先 大衛 的上帝如此說：『我聽見了你的禱告，看見了你的眼淚。看哪，我必加添你十五年的壽數；
ISA|38|6|我要救你和這城脫離 亞述 王的手，也要保護這城。』
ISA|38|7|「耶和華必成就他所說的這話。這是耶和華給你的預兆：
ISA|38|8|看哪，我要使 亞哈斯 日晷上隨太陽前進的影子，往後退十度。」於是，在日晷上照下來的日影果然往後退了十度。
ISA|38|9|猶大 王 希西家 患病痊癒後的詩：
ISA|38|10|我說，在如日中天的時候我就走了， 將剩餘的年歲交給陰間的門。
ISA|38|11|我說，我必不得見耶和華，不得在活人之地見耶和華， 也不再看見世人，就是短暫世界 中的居民。
ISA|38|12|我的住處好像牧人的帳棚， 遭人掀起，離我而去； 我將性命捲起， 像織布的捲布一樣。 他從織布機頭那裏將我剪斷， 你使我命喪於旦夕。
ISA|38|13|我令自己安靜 直到天亮； 他像獅子折斷我所有的骨頭， 你使我命喪於旦夕。
ISA|38|14|我像燕子呢喃， 像白鶴鳴叫， 又如鴿子哀鳴； 我因仰望，眼睛困倦。 主啊，我受欺壓， 求你為我作保。
ISA|38|15|我還有甚麼可說的呢？ 他應許我的 ，他已成就了。 我因心裏的苦楚， 在一生的年日必謙卑而行 。
ISA|38|16|主啊，人得存活是在乎此， 我的靈存活也全在乎此 ； 求你使我痊癒，仍然存活。
ISA|38|17|看哪，我受大苦是為使我得平安； 你愛我，救我的性命脫離敗壞的地府， 將我一切的罪扔在你背後。
ISA|38|18|原來，陰間不能稱謝你， 死亡不能頌揚你， 下到地府的人也不能盼望你的信實。
ISA|38|19|只有活人，活人必稱謝你， 像我今日稱謝你一樣。 為父的，必使兒女知道你的信實。
ISA|38|20|耶和華肯救我， 所以，我們要一生一世 在耶和華殿中 彈奏我弦樂的歌。
ISA|38|21|以賽亞 說：「拿一塊無花果餅來，貼在瘡上，王必痊癒。」
ISA|38|22|希西家 說：「我能上耶和華的殿，有甚麼預兆呢？」
ISA|39|1|那時， 巴拉但 的兒子， 巴比倫 王 米羅達‧巴拉但 聽見 希西家 病得痊癒，就送書信和禮物給他。
ISA|39|2|希西家 歡喜見使者，就將自己寶庫裏的金子、銀子、香料、貴重的膏油和他軍械庫裏一切的兵器，以及他所有的財寶，都給他們看；在他家中和全國之內， 希西家 沒有一樣不給他們看的。
ISA|39|3|於是 以賽亞 先知到 希西家 王那裏去，對他說：「這些人說了些甚麼？他們從哪裏來見你？」 希西家 說：「他們從遠方的 巴比倫 來見我。」
ISA|39|4|以賽亞 說：「他們在你家裏看見了甚麼？」 希西家 說：「凡我家中所有的，他們都看見了；我財寶中沒有一樣東西不給他們看的。」
ISA|39|5|以賽亞 對 希西家 說：「你要聽萬軍之耶和華的話，
ISA|39|6|耶和華說：『看哪，日子將到，凡你家裏所有的，並你祖先積蓄到如今的一切，都要被擄到 巴比倫 去，不留下一樣；
ISA|39|7|從你本身所生的孩子，其中必有被擄到 巴比倫 王宮當太監的。』」
ISA|39|8|希西家 對 以賽亞 說：「你所說耶和華的話甚好。」因為他想：「在我有生之年必有太平和安穩。」
ISA|40|1|你們的上帝說： 「要安慰，安慰我的百姓。
ISA|40|2|要對 耶路撒冷 說安慰的話， 向它宣告， 它的戰爭已結束， 它的罪孽已赦免； 它為自己一切的罪， 已從耶和華手中加倍受罰。」
ISA|40|3|有聲音呼喊著： 「要在曠野為耶和華預備道路， 在沙漠為我們的上帝修直大道。
ISA|40|4|一切山窪都要填滿， 大小山岡都要削平； 陡峭的要變為平坦， 崎嶇的必成為平原。
ISA|40|5|耶和華的榮耀必然顯現， 凡有血肉之軀的都一同看見， 因為這是耶和華親口說的。」
ISA|40|6|有聲音說：「你喊叫吧！」 我 說：「我喊叫甚麼呢？」 凡有血肉之軀的盡都如草， 他的一切榮美像野地的花。
ISA|40|7|耶和華吹一口氣， 草就枯乾，花也凋謝。 百姓誠然是草；
ISA|40|8|草必枯乾，花必凋謝， 惟有我們上帝的話永遠立定。
ISA|40|9|報好信息的 錫安 哪， 要登高山； 報好信息的 耶路撒冷 啊， 要極力揚聲。 揚聲不要懼怕， 對 猶大 的城鎮說： 「看哪，你們的上帝！」
ISA|40|10|看哪，主耶和華必以大能臨到， 他的膀臂必為他掌權； 看哪，他的賞賜在他那裏， 他的報應在他面前。
ISA|40|11|他要像牧人牧養自己的羊群， 用膀臂聚集羔羊，抱在胸懷， 慢慢引導那乳養小羊的。
ISA|40|12|誰曾用手心量諸水， 用手虎口量蒼天， 用升斗盛大地的塵土， 用秤稱山嶺， 用天平稱岡陵呢？
ISA|40|13|誰曾測度耶和華的靈， 或作他的謀士指教他呢？
ISA|40|14|他與誰商議， 誰教導他， 以公平的路指示他， 將知識傳授與他， 又將通達的道指教他呢？
ISA|40|15|看哪，列國都像水桶裏的一滴， 又如天平上的微塵； 看哪，他舉起眾海島，好像舉起極微小之物。
ISA|40|16|黎巴嫩 不夠當柴燒， 其中的走獸也不夠作燔祭。
ISA|40|17|列國在他面前如同不存在， 在他看來微不足道，只是虛空。
ISA|40|18|你們究竟將誰比上帝， 用甚麼形像與他相較呢？
ISA|40|19|至於偶像，匠人鑄造它， 銀匠用金子包裹它， 又為它鑄造銀鏈。
ISA|40|20|沒有能力捐獻的人， 就挑選不易朽壞的木頭， 為自己尋找巧匠， 豎立不會倒的偶像。
ISA|40|21|你們豈不知道嗎？ 豈未曾聽見嗎？ 難道沒有人從起頭就告訴你們嗎？ 自從地的根基立定， 你們豈不明白嗎？
ISA|40|22|上帝坐在地的穹窿之上， 地上的居民有如蚱蜢。 他鋪張穹蒼如幔子， 展開諸天如可住的帳棚。
ISA|40|23|他使君王歸於虛無， 使地上的審判官成為虛空。
ISA|40|24|他們剛栽上， 剛種好， 根也剛扎在地裏， 經他一吹，就都枯乾； 旋風將他們吹去，像碎秸一樣。
ISA|40|25|那聖者說：「你們將誰與我相比， 與我相等呢？」
ISA|40|26|你們要向上舉目， 看是誰創造這萬象， 按數目領出它們， 一一稱其名， 以他的權能 和他的大能大力， 使它們一個都不缺。
ISA|40|27|雅各 啊，你為何說， 以色列 啊，你為何言， 「我的道路向耶和華隱藏， 我的冤屈上帝並不查問」？
ISA|40|28|你豈不曾知道嗎？ 你豈未曾聽見嗎？ 永在的上帝耶和華，創造地極的主， 他不疲乏，也不困倦； 他的智慧無法測度。
ISA|40|29|疲乏的，他賜能力； 軟弱的，他加力量。
ISA|40|30|就是年輕人也要疲乏困倦， 強壯的也必全然跌倒。
ISA|40|31|但那等候耶和華的必重新得力。 他們必如鷹展翅上騰； 他們奔跑卻不困倦， 行走卻不疲乏。
ISA|41|1|眾海島啊，在我面前靜默； 萬民要重新得力， 讓他們近前來陳述， 我們可以彼此辯論。
ISA|41|2|誰從東方興起一人， 憑公義召他來到腳前？ 誰將列國交給他， 使他管轄列王， 把他們如灰塵交與他的刀， 如風吹的碎秸交與他的弓？
ISA|41|3|他追趕君王， 安然走過， 快速地腳不落地 。
ISA|41|4|誰做成這事， 從起初宣召歷代呢？ 就是我－耶和華！ 我是首先的， 也與末後的同在。
ISA|41|5|眾海島看見就都害怕， 地極也都戰兢， 他們近前來；
ISA|41|6|各人互相幫助， 對弟兄說：「壯膽吧！」
ISA|41|7|木匠鼓勵銀匠， 用鎚子打光的鼓勵打砧的， 對銲工說：「銲得好！」 又用釘子釘穩，免得它倒下。
ISA|41|8|惟你 以色列 ，我的僕人， 雅各 ，我所揀選的， 我朋友 亞伯拉罕 的後裔，
ISA|41|9|你是我從地極領來， 從地角召來的， 我對你說：「你是我的僕人； 我揀選你，並不棄絕你。」
ISA|41|10|你不要害怕，因為我與你同在； 不要驚惶，因為我是你的上帝。 我必堅固你，幫助你， 用我公義的右手扶持你。
ISA|41|11|看哪，凡向你發怒的都抱愧蒙羞， 與你相爭的必如無有，並要滅亡。
ISA|41|12|與你爭鬥的，你要尋找他們，卻遍尋不著； 與你爭戰的必如無有，成為虛無。
ISA|41|13|因為我耶和華－你的上帝 必攙扶你的右手， 對你說：「不要害怕！ 我必幫助你。」
ISA|41|14|蟲子 雅各 ， 以色列 人哪， 不要害怕！ 我必幫助你； 救贖你的是 以色列 的聖者。 這是耶和華說的。
ISA|41|15|看哪，我使你成為 全新的打穀機，齒輪銳利； 你要把山嶺打得粉碎， 使岡陵如同糠秕。
ISA|41|16|你要簸揚它們，風要將它們吹去； 旋風要颳散它們。 你卻要以耶和華為喜樂， 因 以色列 的聖者誇耀。
ISA|41|17|困苦貧窮人尋找水，卻尋不著； 他們因口渴，舌頭乾燥。 我－耶和華必應允他們， 我─ 以色列 的上帝必不離棄他們。
ISA|41|18|我要在光禿的高地開江河， 在谷中開泉源； 我要使沙漠變為水池， 使乾地變為湧泉。
ISA|41|19|我要在曠野栽植香柏樹、 皂莢樹、番石榴樹，和野橄欖樹。 在沙漠一同栽上松樹、杉樹， 和黃楊樹，
ISA|41|20|好叫人看見，知道， 思想，明白； 這是耶和華親手做的， 是 以色列 的聖者所造的。
ISA|41|21|耶和華說： 「你們要呈上你們的案件。」 雅各 的君王說： 「你們要提出你們的理由。」
ISA|41|22|讓它們近前來，告訴我們將來要發生甚麼事！ 你們要說明先前發生的事，好讓我們思索； 或者告訴我們將來的事，使我們得知事情的結局。
ISA|41|23|你們要指明未來的事， 使我們知道你們是神明！ 你們或降福，或降禍， 好使我們驚奇，一同觀看。
ISA|41|24|看哪，你們屬乎虛無， 你們的作為也屬虛空； 那選擇你們的是可憎惡的。
ISA|41|25|我從北方興起一人， 他從日出之地而來， 是求告我名的； 他必踩踏 掌權者，如踩踏泥土， 又如陶匠踹泥一般。
ISA|41|26|有誰從起初宣佈這事，使我們知道呢？ 有誰從先前指明，使我們說「他是對的」呢？ 沒有人宣佈， 沒有人指明， 也沒有人聽見你們的話。
ISA|41|27|我首先對 錫安 說，看哪，他們在此！ 我要將一位報好信息的賜給 耶路撒冷 。
ISA|41|28|然而我觀看，並無一人； 我詢問的時候， 他們中間也沒有謀士可回答。
ISA|41|29|看哪，他們盡是麻煩 ， 所做的工都屬虛無； 所鑄的偶像是風，是虛空。
ISA|42|1|看哪，我的僕人， 我所扶持、所揀選、心所喜悅的！ 我已將我的靈賜給他， 他必將公理傳給萬邦。
ISA|42|2|他不喧嚷，不揚聲， 也不使街上聽見他的聲音。
ISA|42|3|壓傷的蘆葦，他不折斷； 將殘的燈火，他不吹滅。 他憑信實將公理傳開。
ISA|42|4|他不灰心，也不喪膽， 直到他在地上設立公理； 眾海島都等候他的訓誨。
ISA|42|5|那創造諸天，鋪張穹蒼， 鋪開地與地的出產， 賜氣息給地上眾人， 賜生命給行走其上之人的 上帝耶和華如此說：
ISA|42|6|「我－耶和華憑公義召你， 要攙扶你的手，保護你， 要藉著你與百姓立約， 使你成為萬邦之光，
ISA|42|7|開盲人的眼， 領囚犯出監獄， 領坐在黑暗中的出地牢。
ISA|42|8|我是耶和華，這是我的名； 我必不將我的榮耀歸給別神 ， 也不將我所得的頌讚歸給雕刻的偶像。
ISA|42|9|看哪，先前的事已經成就， 現在我要指明新事， 告訴你們尚未發生的事。
ISA|42|10|航海的人和海中一切所有的， 眾海島和其中的居民， 都當向耶和華唱新歌， 從地極讚美他。
ISA|42|11|曠野和其中的城鎮， 並 基達 人居住的村莊都當揚聲 ； 西拉 的居民當歡呼， 在山頂上大聲呼喊。
ISA|42|12|願他們將榮耀歸給耶和華， 在海島中傳揚頌讚他的話。
ISA|42|13|耶和華必如勇士出征， 如戰士激起憤恨， 他要喊叫，大聲吶喊， 擊敗他的敵人。
ISA|42|14|我許久閉口不言，沉默不語； 現在我要像臨產的婦人，大聲喊叫， 呼吸急促而喘氣。
ISA|42|15|我要使大小山岡變為荒蕪， 使其上的花草都枯乾； 我要使江河變為沙洲， 使水池盡都乾涸。
ISA|42|16|我要引導盲人行他們所不認識的道， 引領他們走他們未曾走過的路； 我在他們面前使黑暗變為光明， 使彎曲變為平直。 這些事我都要做， 並不離棄他們。
ISA|42|17|但那倚靠雕刻的偶像， 對鑄造的偶像說： 「你是我們的神明」； 這種人要退後，大大蒙羞。
ISA|42|18|你們這耳聾的，聽吧！ 你們這眼瞎的，看吧， 使你們得以看見！
ISA|42|19|誰比我的僕人眼瞎呢？ 誰比我所差遣的使者耳聾呢？ 誰瞎眼像那獻身給我的人？ 誰瞎眼 像耶和華的僕人呢？
ISA|42|20|看見許多事卻不領會， 耳朵開通卻聽不見。
ISA|42|21|耶和華因自己的公義， 樂意使律法為大為尊。
ISA|42|22|但這百姓是被搶被奪的， 全都陷在洞穴中，關在監牢裏； 他們成了掠物，無人拯救， 成了擄物，無人索還。
ISA|42|23|你們中間誰肯側耳聽這話， 誰肯留心聽，以防將來呢？
ISA|42|24|誰將 雅各 交出作為擄物， 將 以色列 交給搶奪者呢？ 豈不是耶和華 ─我們所得罪的那位嗎？ 他們不肯遵行他的道， 也不聽從他的訓誨。
ISA|42|25|所以，他將猛烈的怒氣和戰爭的威力 傾倒在 以色列 身上； 在他周圍如火燃起，他竟然不知， 燒著了，他也不在意。
ISA|43|1|雅各 啊，創造你的耶和華， 以色列 啊，造成你的那位， 現在如此說： 「你不要害怕，因為我救贖了你； 我曾提你的名召你，你是屬我的。
ISA|43|2|你從水中經過，我必與你同在， 你渡過江河，水必不漫過你； 你在火中行走，也不被燒傷， 火焰必不燒著你身。
ISA|43|3|因為我是耶和華－你的上帝， 是 以色列 的聖者－你的救主； 我使 埃及 作你的贖價， 使 古實 和 西巴 代替你。
ISA|43|4|因我看你為寶貝為尊貴； 又因我愛你， 所以使人代替你， 使萬民替換你的生命。
ISA|43|5|你不要害怕，因我與你同在； 我必領你的後裔從東方來， 又從西方召集你。
ISA|43|6|我要對北方說，交出來！ 對南方說，不可扣留！ 要將我的兒子從遠方帶來， 將我的女兒從地極領回，
ISA|43|7|就是凡稱為我名下的人， 是我為自己的榮耀創造的， 是我所塑造，所做成的。」
ISA|43|8|你要將有眼卻瞎、 有耳卻聾的民都帶出來！
ISA|43|9|任憑萬國聚集， 任憑萬民會合。 他們當中誰能說明， 並將先前的事指示我們呢？ 讓他們帶來見證，顯明他們有理， 看是否聽見的人會說：「果然是真的。」
ISA|43|10|你們是我的見證， 是我所揀選的僕人， 為了要使你們知道，且信服我， 又明白我就是耶和華。 在我以前沒有任何被造的真神， 在我以後也必沒有。 這是耶和華說的。
ISA|43|11|我，惟有我是耶和華； 除我以外沒有救主。
ISA|43|12|我曾指示，我曾拯救，我曾說明， 並沒有外族的神明 在你們中間。 你們是我的見證， 我是上帝。 這是耶和華說的。
ISA|43|13|自有日子以來，我就是上帝， 誰也不能救人脫離我的手。 我要行事，誰能逆轉呢？
ISA|43|14|耶和華─你們的救贖主、 以色列 的聖者如此說： 「因你們的緣故， 我已派遣人到 巴比倫 去； 要使 迦勒底 人都如難民， 坐自己素來宴樂的船下來。
ISA|43|15|我是耶和華－你們的聖者， 是創造 以色列 的，是你們的君王。」
ISA|43|16|那在滄海中開道， 在大水中開路， 使戰車、馬匹、軍兵、勇士一同出來， 使他們仆倒，不再起來， 使他們滅沒，好像熄滅之燈火的耶和華如此說：
ISA|43|17|
ISA|43|18|「你們不要追念從前的事， 也不要思想古時的事。
ISA|43|19|看哪，我要行一件新事， 如今就要顯明，你們豈不知道嗎？ 我必在曠野開道路， 在沙漠開江河 。
ISA|43|20|野地的走獸要尊敬我， 野狗和鴕鳥也必尊敬我。 因我使曠野有水， 使沙漠有河， 好賜給我的百姓、我的選民喝。
ISA|43|21|這百姓是我為自己造的， 為要述說我的美德。」
ISA|43|22|「 雅各 啊，你並沒有求告我； 以色列 啊，你倒厭煩我。
ISA|43|23|你並沒有將你的羊帶來獻給我做燔祭， 也沒有用牲祭尊敬我； 我未曾因素祭使你操勞， 也沒有因乳香使你厭煩。
ISA|43|24|你沒有用銀子為我買香菖蒲， 也沒有用祭物的油脂使我飽足； 倒使我因你的罪惡操勞， 使我因你的罪孽厭煩。
ISA|43|25|我，惟有我為自己的緣故塗去你的過犯， 我也不再記得你的罪惡。
ISA|43|26|你儘管提醒我，讓我們來辯論； 儘管陳述，自顯為義。
ISA|43|27|你的始祖犯罪， 你的師傅違背我；
ISA|43|28|因此，我要凌辱聖所的領袖 ， 使 雅各 遭毀滅， 使 以色列 受辱罵。」
ISA|44|1|「我的僕人 雅各 ， 我所揀選的 以色列 啊， 現在你當聽。
ISA|44|2|那位造你，使你在母腹中成形， 並要幫助你的耶和華如此說： 我的僕人 雅各 ， 我所揀選的 耶書崙 哪， 不要害怕！
ISA|44|3|因為我要把水澆灌乾渴的地方， 使水湧流在乾旱之地。 我要將我的靈澆灌你的後裔， 使我的福臨到你的子孫。
ISA|44|4|他們要在草叢中生長 ， 如溪水旁的柳樹。
ISA|44|5|這個要說：『我是屬耶和華的』， 那個要以 雅各 的名自稱， 又有一個在手上寫著：『歸耶和華』， 並自稱為 以色列 。」
ISA|44|6|耶和華－ 以色列 的君王， 以色列 的救贖主－萬軍之耶和華如此說： 「我是首先的，也是末後的； 除我以外再沒有上帝。
ISA|44|7|自從古時我設立了人， 誰能像我宣告，指明，又為自己陳說呢？ 讓他指明未來的事和必成的事吧！
ISA|44|8|你們不要恐懼，也不要害怕。 我豈不是從上古就告訴並指示你們了嗎？ 你們是我的見證人！ 除我以外，豈有上帝呢？ 誠然沒有磐石，就我所知，一個也沒有！」
ISA|44|9|製造偶像的人盡都虛空，他們所喜悅的全無益處；偶像的見證人毫無所見，毫無所知，以致他們羞愧。
ISA|44|10|誰製造神像，鑄造偶像？這些都是無益的。
ISA|44|11|看哪，他的同夥都必羞愧。工匠不過是人，任他們聚集，任他們站立吧！他們都必懼怕，一同羞愧。
ISA|44|12|鐵匠用工具在火炭上工作 ，用鎚打出形狀，用他有力的膀臂來錘。他因飢餓而無力氣；因未喝水而疲倦。
ISA|44|13|木匠拉線，用筆劃出樣子，用鉋子鉋成形狀，又用圓規劃了模樣。他仿照人的體態，做出美妙的人形，放在廟裏。
ISA|44|14|他砍伐香柏樹，又取杉樹和橡樹，在樹林中讓它茁壯；或栽種松樹，得雨水滋潤長大。
ISA|44|15|這樹，人可用以生火；他拿一些來取暖，又搧火烤餅，而且做神像供跪拜，做雕刻的偶像向它叩拜。
ISA|44|16|他將一半的木頭燒在火中，用它烤肉來吃；吃飽了，就自己取暖說：「啊哈，我暖和了，我看到火了！」
ISA|44|17|然後又用剩下的一半做了一個神明，就是雕刻的偶像，向這偶像俯伏叩拜，向它禱告說：「求你拯救我，因你是我的神明。」
ISA|44|18|他們既無知，又不思想；因為耶和華蒙蔽他們的眼，使他們看不見，塞住他們的心，使他們不明白。
ISA|44|19|沒有一個心裏醒悟，有知識，有聰明，能說：「我曾拿一部分用火燃燒，在炭火上烤餅，也烤肉來吃。這剩下的，我豈要做可憎之像嗎？我豈可向木頭叩拜呢？」
ISA|44|20|他以灰塵為食，心裏迷糊，以致偏邪，不能自救，也不能說：「我右手中豈不是有虛謊嗎？」
ISA|44|21|雅各 啊，要思念這些事； 以色列 啊，你是我的僕人。 我造了你，你是我的僕人， 以色列 啊，我必不忘記你 。
ISA|44|22|我塗去你的過犯，像厚雲消散； 塗去你的罪惡，如薄霧消失。 你當歸向我，因我救贖了你。
ISA|44|23|諸天哪，應當歌唱， 因為耶和華成就這事。 地的深處啊，應當歡呼； 眾山哪，要出聲歌唱； 樹林和其中所有的樹木啊，你們都當歌唱！ 因為耶和華救贖了 雅各 ， 並要因 以色列 榮耀自己。
ISA|44|24|從你在母腹中就造了你，你的救贖主－耶和華如此說： 「我－耶和華創造萬物， 獨自鋪張諸天，親自展開大地 ；
ISA|44|25|我使虛謊的預兆失效， 愚弄占卜的人， 使智慧人退後， 使他的知識變為愚拙；
ISA|44|26|卻使我僕人的話站得住， 成就我使者的籌算。 我論 耶路撒冷 說：『必有人居住』； 論 猶大 的城鎮說：『必被建造， 我必重建其中的廢墟。』
ISA|44|27|我對深淵說：『乾了吧！ 我要使你的江河乾涸』；
ISA|44|28|論 居魯士 說：『他是我的牧人， 他要成就我所喜悅的， 下令建造 耶路撒冷 ， 發命令立穩聖殿的根基。』」
ISA|45|1|耶和華對所膏的 居魯士 如此說， 他的右手我曾攙扶， 使列國降服在他面前， 列王的腰帶我曾鬆開， 使城門在他面前敞開， 不得關閉：
ISA|45|2|「我要在你前面行， 修平崎嶇之地。 我必打破銅門， 砍斷鐵閂。
ISA|45|3|我要將暗中的寶物和隱藏的財富賜給你， 使你知道提名召你的 就是我－耶和華， 以色列 的上帝。
ISA|45|4|因我的僕人 雅各 ， 我所揀選的 以色列 ， 我提名召你； 你雖不認識我， 我也加給你名號。
ISA|45|5|我是耶和華，再沒有別的了； 除了我以外再沒有上帝。 你雖不認識我， 我必給你束腰。
ISA|45|6|從日出之地到日落之處使人都知道 除我以外，沒有別的。 我是耶和華，再沒有別的了。
ISA|45|7|我造光，又造暗； 施平安，又降災禍； 做成這一切的是我－耶和華。
ISA|45|8|「諸天哪，要如雨傾盆而降， 雲要降下公義， 地要裂開，救恩湧出 ， 使公義也一同滋長； 這都是我－耶和華造的。」
ISA|45|9|「那與造他的主爭論的人有禍了！ 他不過是地上瓦塊中的一片 。 泥土豈可對塑造它的說：『你做的是甚麼？ 你所做的物怎麼沒有把手呢？ 』
ISA|45|10|有人對父親說， 『你生的是甚麼』， 對母親 說， 『你生產的是甚麼』； 這人有禍了！」
ISA|45|11|耶和華－ 以色列 的聖者， 就是造 以色列 的如此說： 「難道我孩子的未來，你們能質問我， 我手的工作，你們可以吩咐我嗎？
ISA|45|12|我造大地，又創造人在地上。 我親手鋪張諸天， 天上萬象也是我所任命的。
ISA|45|13|我憑公義興起 居魯士 ， 又要修直他一切的道路。 他必建造我的城， 釋放我被擄的民， 不為工價，也不為獎賞。」 這是萬軍之耶和華說的。
ISA|45|14|耶和華如此說： 「 埃及 的出產和 古實 的貨物必歸你； 身量高大的 西巴 人，他們必過來歸你，為你所有。 他們必帶著鎖鏈過來跟隨你， 向你下拜，祈求你說： 『上帝真是在你中間，再沒有別的， 沒有別的上帝。』」
ISA|45|15|救主－ 以色列 的上帝啊， 你誠然是隱藏自己的上帝。
ISA|45|16|製造偶像的都要抱愧蒙羞， 他們要一同歸於慚愧。
ISA|45|17|惟有 以色列 必蒙耶和華拯救， 得永遠的救恩。 你們必不蒙羞，也不抱愧， 直到永世無盡。
ISA|45|18|耶和華如此說， 他創造諸天，他是上帝； 他造了地，形成它，堅固它， 並非創造它為荒涼， 而是要給人居住： 「我是耶和華，再沒有別的。
ISA|45|19|我不在隱密黑暗之地說話， 也沒有對 雅各 的後裔說， 『你們尋求我是徒然的』， 我－耶和華所講的是公義， 所說的是正直。」
ISA|45|20|「你們從列國逃脫的人， 要一同聚集前來。 那些抬著雕刻的木偶、 祈求不能救人之神明的， 毫無知識。
ISA|45|21|你們要近前來說明， 讓他們彼此商議。 誰從古時指明這事？ 誰從上古述說它？ 不是我－耶和華嗎？ 除了我以外，再沒有上帝； 我是公義的上帝，又是救主； 除了我以外，再沒有別的了。
ISA|45|22|「地的四極都當轉向我， 就必得救； 因為我是上帝，再沒有別的。
ISA|45|23|我指著自己起誓， 公義從我的口發出，這話並不返回： 『萬膝必向我跪拜， 萬口必憑我起誓。』
ISA|45|24|人論我說 ， 「公義、能力，惟獨在乎耶和華。 人必歸向他， 凡向他發怒的都必蒙羞。
ISA|45|25|以色列 的後裔必因耶和華得稱為義， 並要彼此誇耀。」
ISA|46|1|彼勒 叩拜， 尼波 屈身； 巴比倫 的偶像馱在走獸和牲畜背上。 你們所抬的成了重馱， 使牲畜疲乏。
ISA|46|2|這些神明一同屈身叩拜， 不能救自己 ， 反倒遭人擄去。
ISA|46|3|雅各 家， 以色列 家所有的餘民哪， 你們自從生下就蒙我抱， 自出母胎便由我來背， 你們都要聽從我。
ISA|46|4|直到你們年老，我不改變； 直到你們髮白，我仍扶持。 我已造你，就必背你； 我必抱你，也必拯救。
ISA|46|5|你們將誰與我相比，與我相等， 將誰與我相較，使我們相似呢？
ISA|46|6|他們從錢囊中倒出金子， 用天平秤出銀子， 雇銀匠造成神像， 他們又俯伏，又叩拜。
ISA|46|7|他們抬起神像，扛在肩上， 安置在定處，使它站立， 不離本位； 人呼求它，它卻不回答， 也無法救人脫離災難。
ISA|46|8|你們當記得這事，立定心意 。 叛逆的人哪，要留心思想。
ISA|46|9|要追念上古的事， 因為我是上帝，並無別的； 我是上帝，沒有能與我相比的。
ISA|46|10|我從起初就指明末後的事， 從古時便言明未成的事， 說：「我的籌算必立定； 凡我所喜悅的，我必成就。」
ISA|46|11|我召鷙鳥從東方來， 召那成就我籌算的人從遠方來。 我已說出，就必成就； 我已謀定，也必做成。
ISA|46|12|你們這些心中頑固、 遠離公義的人，要聽從我。
ISA|46|13|我使我的公義臨近，它已不遠。 我的救恩必不遲延。 我要為 以色列 －我的榮耀 在 錫安 施行救恩。
ISA|47|1|少女 巴比倫 哪， 下來坐在塵埃； 迦勒底 啊， 沒有寶座，要坐在地上； 你不再稱為柔弱嬌嫩。
ISA|47|2|要用磨磨麵， 揭去面紗， 脫去長裙， 露腿渡河。
ISA|47|3|你的下體必被露出； 你的羞辱必被看見。 我要報復， 誰也不寬容 。
ISA|47|4|我們的救贖主是 以色列 的聖者， 他的名為萬軍之耶和華。
ISA|47|5|迦勒底 啊， 你要靜坐，進入黑暗中， 因你不再稱為萬國之后。
ISA|47|6|我向我的百姓發怒， 使我的產業受凌辱， 將他們交在你手中； 然而你毫不憐憫他們， 連老年人你也加極重的軛。
ISA|47|7|你說：「我必永遠為后。」 你不將這事放在心上， 也不思想事情的結局。
ISA|47|8|你這專好宴樂、以為地位穩固的， 現在當聽這話。 你心中說： 「惟有我，除我以外再沒有別的。 我必不致寡居， 也不經歷喪子之痛。」
ISA|47|9|哪知，喪子、寡居這兩件事 一日之間忽然臨到你； 你雖多行邪術、廣施魔咒， 這兩件事必全然臨到你身上。
ISA|47|10|你倚靠自己的惡行，說： 「無人看見我。」 你的智慧聰明使你走偏， 你心裏說： 「惟有我，除我以外再沒有別的了。」
ISA|47|11|但災禍臨到你， 你不知如何驅除； 災害落在你身上， 你也無法除掉， 你所不知道的毀滅必忽然臨到你身上。
ISA|47|12|儘管使用從幼年就施行的魔符和眾多的邪術吧！ 或許有些幫助， 或許可以致勝。
ISA|47|13|你籌劃太多，以致疲倦。 讓那些觀天象，看星宿， 在初一說預言的都起來， 救你脫離所要臨到你的事！
ISA|47|14|看哪，他們要像碎秸被火焚燒， 無法救自己脫離火焰的魔掌； 沒有炭火可以取暖 ， 你也不能坐在火旁。
ISA|47|15|你所操勞的事都像這樣； 從你幼年以來與你交易的都各奔己路， 沒有一人來救你。
ISA|48|1|雅各 家，稱為 以色列 名下， 從 猶大 的源頭而出的啊， 你們指著耶和華的名起誓， 提說 以色列 的上帝， 卻不憑誠信，也不憑公義； 你們自稱為聖城之民， 倚靠名為萬軍之耶和華－ 以色列 的上帝； 現在，當聽我言：
ISA|48|2|
ISA|48|3|「先前的事，我自古已說明， 已從我口而出， 是我所指示的； 我瞬間行事，事便成就。
ISA|48|4|因為我知道你是頑梗的； 你的頸項是鐵的， 你的額頭是銅的。
ISA|48|5|所以，我自古就給你說明， 在事未成以先指示你， 免得你說：『這些事是我的偶像所行的， 是我雕刻的偶像和鑄造的神像所命定的。』
ISA|48|6|「你既已聽見，現在要察看這一切； 你們不是要說明嗎？ 從今以後，我要指示你新事， 就是你所不知道的隱密事。
ISA|48|7|這事是現今造的，並非自古就有， 在今日以先，你未曾聽見； 免得你說：『看哪，這事我早已知道了。』
ISA|48|8|誠然你未曾聽見，也未曾知道； 你的耳朵從來未曾開通。 我原知道你行事極其詭詐， 你自從出母胎以來， 就稱為悖逆的。
ISA|48|9|「我為我的名暫且忍怒， 為了我的榮耀向你容忍， 不將你剪除。
ISA|48|10|看哪，我熬煉你，卻不像熬煉銀子； 你在苦難的火爐中，我試煉 你。
ISA|48|11|我為自己的緣故必做這事， 我豈能被褻瀆？ 我必不將我的榮耀歸給別神 。
ISA|48|12|雅各 －我所選召的 以色列 啊， 當聽從我： 我是耶和華， 「我是首先的，也是末後的。
ISA|48|13|我親手立了地的根基， 以右手鋪張諸天； 我一召喚，天地就都立定。
ISA|48|14|你們都當聚集而聽， 偶像 之中誰曾說明這些事？ 耶和華愛他，他必向 巴比倫 成就耶和華的旨意， 耶和華的膀臂也要加在 迦勒底 人身上 。
ISA|48|15|我，惟有我曾說過， 我選召他，領他來， 他的道路必亨通。
ISA|48|16|你們要接近我來聽這話， 我從起初就未曾在隱密之處說話， 萬事之始，我就在那裏。」 現在，主耶和華差遣了我， 帶著他的靈而來 。
ISA|48|17|耶和華－你的救贖主， 以色列 的聖者如此說： 「我是耶和華－你的上帝， 我教導你，使你得益處， 指引你當走的路。
ISA|48|18|甚願你聽從我的命令， 你的平安就會如河水， 你的公義如海浪，
ISA|48|19|你的後裔必多如海沙， 你腹中所生的必多如沙粒。 他的名絕不從我面前剪除， 也不滅絕。」
ISA|48|20|你們要從 巴比倫 出來， 從 迦勒底 人中逃脫， 以歡呼的聲音宣告， 將這事傳揚到地極，說： 耶和華救贖了他的僕人 雅各 ！
ISA|48|21|他引導他們經過沙漠， 他們卻未嘗乾渴； 他為他們使水從磐石流出， 磐石裂開，水就湧出。
ISA|48|22|耶和華說： 「惡人必不得平安！」
ISA|49|1|眾海島啊，當聽從我！ 遠方的眾民哪，要留心聽！ 自出母胎，耶和華就選召我； 自出母腹，他就稱呼我的名。
ISA|49|2|他使我的口如快刀， 把我藏在他手蔭之下； 又使我成為磨利的箭， 把我藏在他箭袋之中；
ISA|49|3|對我說：「你是我的僕人 以色列 ； 我必因你得榮耀。」
ISA|49|4|我卻說：「我勞碌是徒然， 我盡力是虛無虛空。 耶和華誠然以公平待我， 我的賞賜在我的上帝那裏。」
ISA|49|5|現在耶和華說話，他從我出母胎，就造我作他的僕人， 要使 雅各 歸向他， 使 以色列 聚集在他那裏。 耶和華看我為尊貴， 我的上帝是我的力量。
ISA|49|6|他說：「你作我的僕人， 使 雅各 眾支派復興， 使 以色列 中蒙保存的人歸回； 然而此事尚小， 我還要使你作萬邦之光， 使你施行我的救恩，直到地極。」
ISA|49|7|救贖主－ 以色列 的聖者耶和華 對那被人藐視、本國憎惡、 統治者奴役的如此說： 「君王看見就站起來， 領袖也要下拜； 這都是因信實的耶和華， 因揀選你的 以色列 的聖者。」
ISA|49|8|耶和華如此說： 「在悅納的時候，我應允了你； 在拯救的日子，我幫助了你。 我要保護你， 要藉著你與百姓立約， 為了復興遍地， 使人承受荒蕪之地為業；
ISA|49|9|對那被捆綁的人說：『出來吧！』 對在黑暗裏的人說：『顯現吧！』 他們在路上必得飲食， 在光禿的高地必有食物。
ISA|49|10|他們不飢不渴， 炎熱和烈日必不傷害他們； 因為憐憫他們的必引導他們， 領他們到水泉旁邊。
ISA|49|11|我必在眾山開闢路徑， 大道也要填高。
ISA|49|12|看哪，他們從遠方來； 有些從北方來，有些從西方來， 有些從 色弗尼 地來。」
ISA|49|13|諸天哪，應當歡呼！ 大地啊，應當快樂！ 眾山哪，應當揚聲歌唱！ 因為耶和華已經安慰他的百姓， 他要憐憫他的困苦之民。
ISA|49|14|錫安 說：「耶和華離棄了我， 主忘記了我。」
ISA|49|15|婦人焉能忘記她吃奶的嬰孩， 不憐憫她所生的兒子？ 即或有忘記的， 我卻不忘記你。
ISA|49|16|看哪，我將你銘刻在我掌上， 你的城牆常在我眼前。
ISA|49|17|建立你的勝過毀壞你的， 使你荒廢的必都離你而去。
ISA|49|18|你舉目向四圍觀看， 他們都聚集來到你這裏。 我指著我的永生起誓， 你定要以他們為妝飾佩戴， 帶著他們，像新娘一樣。 這是耶和華說的。
ISA|49|19|至於你荒廢淒涼之處， 並你被毀壞之地， 如今居民必嫌太窄， 吞滅你的必離你遙遠。
ISA|49|20|你要再聽見喪失子女後所生的兒女說： 「這地方我居住太窄， 請你給我地方居住。」
ISA|49|21|那時你心裏必說：「我既喪子不育， 被擄，飄流在外 ， 誰給我生了這些？ 誰將他們養大呢？ 看哪，我被撇下獨自一人時， 他們都在哪裏呢？」
ISA|49|22|主耶和華如此說： 「看哪，我必向列國舉手， 向萬民豎立大旗； 他們必將你的兒子抱在懷中帶來， 將你的女兒背在肩上扛來。
ISA|49|23|列王必作你的養父， 王后必作你的乳母。 他們必以臉伏地，向你下拜， 並舔你腳上的塵土。 你就知道我是耶和華， 等候我的必不致羞愧。」
ISA|49|24|勇士搶去的豈能奪回？ 被殘暴者擄掠的豈能得解救呢？
ISA|49|25|但耶和華如此說： 「就是勇士所擄掠的，也可以奪回； 殘暴者所搶的，也可以得解救。 與你相爭的，我必與他相爭， 我也要拯救你的兒女。
ISA|49|26|我必使那欺壓你的吃自己的肉， 飲自己的血，如喝甜酒喝醉一樣。 凡有血肉之軀的都必知道我－耶和華是你的救主， 是你的救贖主，是 雅各 的大能者。」
ISA|50|1|耶和華如此說： 「我休了你們的母親， 她的休書在哪裏呢？ 我將你們賣給了我哪一個債主呢？ 看哪，你們被賣是因你們的罪孽； 你們的母親被休，是因你們的過犯。
ISA|50|2|我來的時候，為何沒有人呢？ 我呼喚的時候，為何無人回應呢？ 我的膀臂豈是過短、不能救贖嗎？ 我豈無拯救之力嗎？ 看哪，我一斥責，海就乾了； 我使江河變為曠野， 其中的魚因無水腥臭，乾渴而死。
ISA|50|3|我使諸天以黑暗為衣， 以麻布為遮蓋。」
ISA|50|4|主耶和華賜我受教者的舌頭， 使我知道怎樣用言語扶助疲乏的人。 主每天早晨喚醒，喚醒我的耳朵， 使我能聽，像受教者一樣。
ISA|50|5|主耶和華開啟我的耳朵， 我並未違背，也未退後。
ISA|50|6|人打我的背，我任他打； 人拔我兩頰的鬍鬚，我由他拔； 人侮辱我，向我吐唾沫，我並不掩面。
ISA|50|7|主耶和華必幫助我， 所以我不抱愧。 我硬著臉面好像堅石， 也知道我必不致蒙羞。
ISA|50|8|稱我為義的與我相近； 誰與我爭論， 讓我們來對質； 誰與我作對， 讓他近前來吧！
ISA|50|9|看哪，主耶和華必幫助我， 誰能定我有罪呢？ 看哪，他們都要像衣服漸漸破舊， 被蛀蟲蛀光。
ISA|50|10|你們當中有誰是敬畏耶和華， 聽從他僕人的話語， 卻行在黑暗中，沒有亮光的， 當倚靠耶和華的名， 仰賴自己的上帝。
ISA|50|11|看哪，你們當中所有點火、以火把圍繞自己的人， 當行走在你們的火焰 裏， 並你們所點的火把中。 這是我親手為你們定的： 你們必躺臥在悲慘之中。
ISA|51|1|追求公義、 尋求耶和華的人哪， 當聽從我！ 你們要追想自己是從哪塊磐石鑿出， 從哪個巖穴挖掘而來；
ISA|51|2|要追想你們的祖宗 亞伯拉罕 和生你們的 撒拉 ； 因為我選召 亞伯拉罕 時，他只有一個人， 但我賜福給他， 使他增多。
ISA|51|3|耶和華已經安慰 錫安 ， 安慰了 錫安 一切的廢墟， 使曠野如 伊甸 ， 使沙漠像耶和華的園子； 其中必有歡喜、快樂、感謝， 和歌唱的聲音。
ISA|51|4|我的民哪，要留心聽我， 我的國啊，要向我側耳； 因為訓誨必從我而出， 我必使我的公理成為萬民之光。
ISA|51|5|我的公義臨近， 我的救恩發出。 我的膀臂要審判萬民， 眾海島都要等候我，倚賴我的膀臂。
ISA|51|6|你們要向天舉目， 觀看下面的地； 天必像煙雲消散， 地必如衣服漸漸破舊； 其上的居民也要如此 死亡。 惟有我的救恩永遠長存， 我的公義也不廢掉。
ISA|51|7|知道公義、將我的訓誨存在心中的人哪， 當聽從我！ 不要怕人的辱罵， 也不要因人的毀謗驚惶。
ISA|51|8|因為他們必像衣服被蛀蟲蛀； 像羊毛被蟲子咬。 惟有我的公義永遠長存， 我的救恩直到萬代。
ISA|51|9|耶和華的膀臂啊，興起，興起！ 以能力為衣穿上， 像古時的年日，像上古的世代一樣興起！ 從前砍碎 拉哈伯 、 刺透大魚的，不是你嗎？
ISA|51|10|使海與深淵的水乾涸， 在海的深處開路， 使救贖的民走過的，不是你嗎？
ISA|51|11|耶和華救贖的民必歸回， 歌唱來到 錫安 ； 永恆的喜樂必歸到他們頭上。 他們必得著歡喜快樂， 憂傷嘆息盡都逃避。
ISA|51|12|我，惟有我是安慰你們的。 你是誰，竟怕那必死的人， 怕那生命如草的世人，
ISA|51|13|卻忘記鋪張諸天、立定地基、 造你的耶和華？ 你因欺壓者圖謀毀滅所發的暴怒， 終日害怕， 其實那欺壓者的暴怒在哪裏呢？
ISA|51|14|被擄的即將得釋放， 不至於死而下入地府， 也不致缺乏食物。
ISA|51|15|我是耶和華－你的上帝， 我攪動大海，使海中的波浪澎湃， 萬軍之耶和華是我的名。
ISA|51|16|我已將我的話放在你口中， 用我的手影遮蔽你， 為要安定諸天，立定地基， 並對 錫安 說：「你是我的百姓。」
ISA|51|17|耶路撒冷 啊，興起，興起！ 站起來！ 你從耶和華手中喝了他憤怒的杯， 那使人東倒西歪的杯，直到喝盡。
ISA|51|18|她所生育的孩子中，沒有一個攙她的； 她所撫養的孩子中，沒有一個扶她的。
ISA|51|19|這雙重的災難臨到你， 有誰憐憫你呢？ 破壞和毀滅，饑荒和戰爭臨到， 我如何能安慰你呢 ？
ISA|51|20|你的孩子發昏， 在各街頭躺臥， 如同網羅裏的羚羊， 滿了耶和華的憤怒， 滿了你上帝的斥責。
ISA|51|21|因此，你這困苦卻非因酒而醉的， 當聽這話，
ISA|51|22|你的主，耶和華， 就是為他百姓辯護的上帝如此說： 「看哪，我已從你手中接過 那使人東倒西歪的杯， 就是我憤怒的杯， 你必不再喝。
ISA|51|23|我必將這杯遞在苦待你的人 手中。 他們曾對你說：『你屈身， 任我們踐踏過去吧！』 你就以背為地， 又如街道，任人走過。
ISA|52|1|錫安 哪，興起！興起！ 穿上你的能力！ 聖城 耶路撒冷 啊，穿上你華美的衣服！ 因為從今以後， 未受割禮、不潔淨的必不再進入你中間。
ISA|52|2|耶路撒冷 啊，抖去塵埃， 起來坐在王位上！ 被擄的 錫安 哪， 解開你頸上的鎖鏈！
ISA|52|3|耶和華如此說：「你們白白地被賣，也必不用銀子贖回。」
ISA|52|4|主耶和華如此說：「先前我的百姓下到 埃及 ，在那裏寄居，末後又有 亞述 人欺壓他們。」
ISA|52|5|我的百姓既是白白地被擄，如今我在這裏做甚麼呢？這是耶和華說的。轄制他們的人歡呼 ，我的名終日不斷受褻瀆，這是耶和華說的。
ISA|52|6|因此，我的百姓必認識我的名；在那日，他們必知道說這話的就是我。看哪，是我！」
ISA|52|7|在山上報佳音，傳平安， 報好信息，傳揚救恩， 那人的腳蹤何等佳美啊！ 他對 錫安 說：「你的上帝作王了！」
ISA|52|8|聽啊，你守望之人的聲音， 他們揚聲一同歡唱； 因為他們必親眼看見耶和華返回 錫安 。
ISA|52|9|耶路撒冷 的廢墟啊， 要出聲一同歡唱； 因為耶和華安慰了他的百姓， 救贖了 耶路撒冷 。
ISA|52|10|耶和華在萬國眼前露出聖臂， 地的四極都要看見我們上帝的救恩。
ISA|52|11|離開吧！離開吧！ 你們要從 巴比倫 出來。 你們扛抬耶和華器皿的人哪， 不要沾不潔淨的東西， 離去時務要保持潔淨。
ISA|52|12|你們出來必不致匆忙， 也不致奔逃； 因為耶和華要在你們前頭行， 以色列 的上帝必作你們的後盾。
ISA|52|13|看哪，我的僕人行事必有智慧， 他必被高升，高舉， 升到至高之處。
ISA|52|14|許多人因他 驚奇 ─他的面貌比別人憔悴， 他的外表比世人枯槁─
ISA|52|15|同樣，他也必使許多國家驚奇 ， 君王要向他閉口。 未曾傳給他們的，他們必看見； 未曾聽見過的事，他們要明白。
ISA|53|1|我們所傳的有誰信呢？ 耶和華的膀臂向誰顯露呢？
ISA|53|2|他在耶和華面前生長如嫩芽， 像根出於乾地。 他無佳形美容使我們注視他， 也無美貌使我們仰慕他。
ISA|53|3|他被藐視，被人厭棄； 多受痛苦，常經憂患。 他被藐視， 好像被人掩面不看的一樣， 我們也不尊重他。
ISA|53|4|他誠然擔當我們的憂患， 背負我們的痛苦； 我們卻以為他受責罰， 是被上帝擊打苦待。
ISA|53|5|他為我們的過犯受害， 為我們的罪孽被壓傷。 因他受的懲罰，我們得平安； 因他受的鞭傷，我們得醫治。
ISA|53|6|我們都如羊走迷， 各人偏行己路； 耶和華使我們眾人的罪孽都歸在他身上。
ISA|53|7|他被欺壓受苦， 卻不開口； 他像羔羊被牽去宰殺， 又像羊在剪毛的人手下無聲， 他也是這樣不開口。
ISA|53|8|因受欺壓和審判，他被奪去， 誰能想到他的世代呢？ 因為他從活人之地被剪除， 為我百姓 的罪過他被帶到死裏 。
ISA|53|9|他雖然未行殘暴， 口中也沒有詭詐， 人還使他與惡人同穴， 與財主同墓 。
ISA|53|10|耶和華的旨意要壓傷他， 使他受苦。 當他的生命作為贖罪祭時 ， 他必看見後裔，他的年日必然長久。 耶和華所喜悅的事，必在他手中亨通。
ISA|53|11|因自己的勞苦，他必看見光 就心滿意足。 因自己的認識，我的義僕使許多人得稱為義， 他要擔當他們的罪孽。
ISA|53|12|因此，我要使他與位大的同份， 與強盛的均分擄物。 因為他傾倒自己的生命，以致於死， 也列在罪犯之中。 他卻擔當多人的罪， 為他們的過犯代求 。
ISA|54|1|你這不懷孕、不生育的，要歡呼； 你這未曾經過產難的，要歡呼，揚聲呼喊； 因為被遺棄的婦人， 比有丈夫的人兒女更多； 這是耶和華說的。
ISA|54|2|要擴張你帳幕之地， 伸展你居所的幔子，不要縮回； 要放長你的繩子， 堅固你的橛子。
ISA|54|3|因為你要向左向右開展， 你的後裔必得列國為業， 又使荒廢的城鎮有人居住。
ISA|54|4|不要懼怕，因你必不致蒙羞； 不要抱愧，因你必不致受辱。 你必忘記年輕時的羞愧， 不再記得守寡的恥辱。
ISA|54|5|因為造你的是你的丈夫， 萬軍之耶和華是他的名； 救贖你的是 以色列 的聖者， 他必稱為全地之上帝。
ISA|54|6|耶和華召你， 如同召回心中憂傷遭遺棄的婦人， 就是年輕時所娶被遺棄的妻子； 這是你的上帝說的。
ISA|54|7|我離棄你不過片時， 卻要大施憐憫將你尋回。
ISA|54|8|我因漲溢的怒氣， 一時向你轉臉， 但我要以永遠的慈愛憐憫你； 這是耶和華－你的救贖主說的。
ISA|54|9|這事於我有如 挪亞 的洪水； 我怎樣起誓不再使 挪亞 的洪水淹沒全地， 也照樣起誓不再向你發怒， 且不斥責你。
ISA|54|10|大山可以挪開， 小山可以遷移， 但我的慈愛必不離開你， 我平安的約也不遷移； 這是憐憫你的耶和華說的。
ISA|54|11|你這受困苦、被暴風捲走、不得憐憫的城， 看哪，我必以灰泥來做你的石頭， 以藍寶石立你的根基，
ISA|54|12|又以紅寶石造你的女牆， 以晶瑩的珠玉造你的城門， 以珍貴的寶石造你四圍的邊界。
ISA|54|13|你的兒女都要領受耶和華的教導， 你的兒女必大享平安。
ISA|54|14|你必因公義得堅立， 必遠離欺壓，毫不懼怕； 你必遠離驚嚇，驚嚇必不臨近你。
ISA|54|15|若有人攻擊你，這非出於我； 凡攻擊你的，必因你仆倒。
ISA|54|16|看哪，我造了那吹炭火、打造合用兵器的鐵匠； 我也造了那殘害人、行毀滅的人。
ISA|54|17|凡為攻擊你而造的兵器必無效用； 在審判時興起用口舌攻擊你的， 你必駁倒他。 這是耶和華僕人的產業， 是他們從我所得的義； 這是耶和華說的。
ISA|55|1|來！你們所有乾渴的，都當來到水邊； 沒有銀錢的也可以來。 你們都來，買了吃； 不用銀錢，不付代價， 就可買酒和奶。
ISA|55|2|你們為何花錢買那不是食物的東西， 用勞碌得來的買那無法使人飽足的呢？ 你們要留意聽從我的話，就能吃那美物， 得享肥甘，心中喜樂。
ISA|55|3|當側耳而聽，來到我這裏； 要聽，就必存活。 我要與你們立永約， 就是應許給 大衛 那可靠的慈愛。
ISA|55|4|看哪，我已立他作萬民的見證， 立他作萬民的君王和發令者。
ISA|55|5|看哪，你要召集素不認識的國民， 素不認識的國民要奔向你； 這都因耶和華─你的上帝， 因 以色列 的聖者已經榮耀了你。
ISA|55|6|當趁耶和華可尋找的時候尋找他， 在他接近的時候求告他。
ISA|55|7|惡人當離棄自己的道路， 不義的人應除掉自己的意念。 歸向耶和華，耶和華就必憐憫他； 當歸向我們的上帝，因為他必廣行赦免。
ISA|55|8|我的意念非同你們的意念， 我的道路非同你們的道路。 這是耶和華說的。
ISA|55|9|天怎樣高過地， 照樣，我的道路高過你們的道路， 我的意念高過你們的意念。
ISA|55|10|雨雪從天而降，並不返回， 卻要滋潤土地，使地面發芽結實， 使撒種的有種，使要吃的有糧。
ISA|55|11|我口所出的話也必如此， 絕不徒然返回， 卻要成就我的旨意， 達成我差它的目的。
ISA|55|12|你們必歡歡喜喜出來， 平平安安蒙引導。 大山小山必在你們面前歡呼， 田野的樹木也都拍掌。
ISA|55|13|松樹長出，代替荊棘； 番石榴長出，代替蒺藜。 這要為耶和華留名， 作為永不磨滅的證據。
ISA|56|1|耶和華如此說： 「你們當守公平，行公義； 因我的救恩臨近， 我的公義將要顯現。
ISA|56|2|謹守安息日不予干犯， 禁止己手不作惡， 如此行、如此持守的人有福了！」
ISA|56|3|與耶和華聯合的外邦人不要說： 「耶和華將我和他的子民分別出來。」 太監也不要說：「看哪，我是枯樹。」
ISA|56|4|因為耶和華如此說： 「那些謹守我的安息日， 選擇我旨意， 持守我約的太監，
ISA|56|5|我必使他們在我殿中，在我牆內， 有紀念碑，有名號， 勝過有兒有女； 我必賜他們永遠的名，不能剪除。
ISA|56|6|「那些與耶和華聯合， 事奉他，愛他名， 作他僕人的外邦人， 凡謹守安息日不予干犯， 又持守我約的人，
ISA|56|7|我必領他們到我的聖山， 使他們在我的禱告的殿中喜樂。 他們的燔祭和祭物， 在我壇上必蒙悅納， 因我的殿必稱為萬民禱告的殿。
ISA|56|8|我還要召集更多的人 歸併到這些被召集的人中。 這是召集被趕散的 以色列 人的 主耶和華說的。」
ISA|56|9|野地的走獸，你們都來吞吃吧！ 林中的野獸，你們也來吞吃！
ISA|56|10|以色列 的守望者都瞎了眼， 沒有知識； 都是啞狗，不會吠叫， 只知做夢，躺臥，貪睡，
ISA|56|11|這些狗貪食，不知飽足。 這些牧人不知明辨， 他們都偏行己路， 人人追求自己的利益。
ISA|56|12|他們說：「來吧！我去拿酒， 讓我們暢飲烈酒吧！ 明天必和今天一樣， 甚至更好！」
ISA|57|1|義人死亡， 無人放在心上； 虔誠的人被接去， 無人理解； 義人被接去，以免禍患。
ISA|57|2|行為正直的人進入平安， 得以在床上安歇 。
ISA|57|3|到這裏來吧！ 你們這些巫婆的兒子， 姦夫和妓女的後代；
ISA|57|4|你們向誰戲笑？ 向誰張口吐舌呢？ 你們豈不是叛逆所生的兒女， 虛謊所生的後代嗎？
ISA|57|5|你們在橡樹 中間，在各青翠的樹下慾火攻心； 在山谷間，在巖隙下殺了兒女；
ISA|57|6|去拜谷中光滑的石頭有你們的份， 這些就是你們的命運。 你向它們獻澆酒祭，獻供物， 這事我豈能容忍嗎？
ISA|57|7|你在高而又高的山上安設床舖， 上那裏去獻祭。
ISA|57|8|你在門後，在門框後， 立起你的牌來； 你離棄了我，赤露己身， 又爬上自己所鋪寬闊的床鋪， 與它們立約； 你喜愛它們的床，看著它們的赤體 。
ISA|57|9|你帶了油到 摩洛 那裏， 加上許多香水。 你派遣使者往遠方去， 甚至降到陰間，
ISA|57|10|因路途遙遠，你就疲倦， 卻不說，這是枉然， 以為能找到復興之力， 所以不覺疲憊。
ISA|57|11|你怕誰，因誰恐懼， 竟說謊，不記得我， 不將這事放在心上。 是否因我許久閉口不言， 你就不怕我了呢？
ISA|57|12|我可以宣告你的公義和你的作為， 但它們與你無益。
ISA|57|13|你哀求的時候， 讓你所搜集的神像 拯救你吧！ 風要把它們全都颳散， 吹一口氣就都吹走。 但那投靠我的必得地產， 承受我的聖山為業。
ISA|57|14|耶和華說： 「你們要修築，修築，要預備道路， 除掉我百姓路中的絆腳石。」
ISA|57|15|那至高無上、永遠長存、 名為聖者的如此說： 「我住在至高至聖的所在， 卻與心靈痛悔的謙卑人同住； 要使謙卑的人心靈甦醒， 使痛悔的人內心復甦。
ISA|57|16|我必不長久控訴，也不永遠懷怒， 因為我雖使靈性發昏，我也造了人的氣息。
ISA|57|17|我因人貪婪的罪孽，發怒擊打他； 我轉臉向他發怒， 他卻仍隨意背道而行。
ISA|57|18|我看見他的行為， 要醫治他，引導他 ， 使他和與他一同哀傷的人都得安慰。
ISA|57|19|我要醫治他， 他要結出嘴唇的果實。 平安，平安，歸給遠處和近處的人！ 這是耶和華說的。」
ISA|57|20|但是惡人好像翻騰的海， 不得平靜； 其中的水常湧出污穢和淤泥。
ISA|57|21|我的上帝說：「惡人必不得平安！」
ISA|58|1|你要大聲喊叫，不要停止； 要揚聲，好像吹角； 向我的百姓宣告他們的過犯， 向 雅各 家陳述他們的罪惡。
ISA|58|2|他們天天尋求我， 樂意明白我的道， 好像行義的國家， 未離棄它的上帝的典章； 他們向我求問公義的判詞， 喜悅親近上帝。
ISA|58|3|「我們禁食，你為何不看呢？ 我們刻苦己心，你為何不理會呢？」 看哪，你們禁食的時候仍追求私利， 剝削為你們做苦工的人。
ISA|58|4|看哪，你們禁食，卻起紛爭興訟， 以兇惡的拳頭打人。 你們今日這種禁食 無法使你們的聲音聽聞於高處。
ISA|58|5|這豈是我所要的禁食， 為人所用以刻苦己心的日子嗎？ 我難道只是叫人如蘆葦般低頭， 鋪上麻布和灰燼嗎？ 你能稱此為禁食， 為耶和華所悅納的日子嗎？
ISA|58|6|我所要的禁食，豈不是要你鬆開兇惡的繩， 解開軛上的索， 使被欺壓的得自由， 折斷一切的軛嗎？
ISA|58|7|豈不是要你把食物分給飢餓的人， 將流浪的窮人接到家中， 見赤身的給他衣服遮體， 而不隱藏自己避開你的骨肉嗎？
ISA|58|8|這樣，必有光如晨光破曉照耀你， 你也要快快得到醫治； 你的公義在你前面行， 耶和華的榮光必作你的後盾。
ISA|58|9|那時你求告，耶和華必應允； 你呼求，他必說：「我在這裏。」 你若從你中間除掉重軛 和指摘人的指頭，並發惡言的事，
ISA|58|10|向飢餓的人施憐憫， 使困苦的人得滿足； 你在黑暗中就必得著光明， 你的幽暗必變如正午。
ISA|58|11|耶和華必時常引導你， 在乾旱之地使你心滿意足， 又使你骨頭強壯。 你必如有水澆灌的園子， 又像水流不絕的泉源。
ISA|58|12|你們中間必有人起來修造久已荒廢之處， 立起代代相承的根基。 你必稱為修補裂痕的， 和重修路徑給人居住的。
ISA|58|13|你若禁止自己的腳踐踏安息日， 不在我的聖日做自己高興的事， 稱安息日為「可喜樂的」， 稱耶和華的聖日為「可尊重的」， 尊敬這日， 不走自己的道路， 不求自己的喜悅， 也不隨意說話；
ISA|58|14|那麼，你就會以耶和華為樂。 耶和華要使你乘駕於地的高處， 又要以你祖先 雅各 的產業養育你； 這是耶和華親口說的。
ISA|59|1|看哪，耶和華的膀臂並非過短，不能拯救， 耳朵並非發沉，不能聽見，
ISA|59|2|但你們的罪孽使你們與上帝隔絕， 你們的罪惡使他轉臉不聽你們。
ISA|59|3|因你們的手掌被血沾染， 你們的指頭被罪玷污， 你們的嘴唇說謊言， 你們的舌頭出惡語。
ISA|59|4|無人按公義控訴， 也無人憑誠實辯白； 卻倚靠虛妄，口說謊言， 懷毒害，生罪孽。
ISA|59|5|他們孵毒蛇蛋， 結蜘蛛網。 凡吃這蛋的必死， 蛋一打破，就孵出蛇來。
ISA|59|6|所結的網不能當衣服， 無法掩蓋自己所作所為。 他們的行為全是邪惡， 手所做的盡都殘暴。
ISA|59|7|他們的腳奔跑行惡， 急速流無辜者的血； 他們的思想全是惡念， 走過的路盡是破壞與毀滅。
ISA|59|8|平安的路，他們不知道， 所行的事無一公平。 他們為自己修築彎曲的路， 凡走這路的都不得平安。
ISA|59|9|因此，公平離我們甚遠， 公義追不上我們。 我們指望光亮，看哪，卻只有黑暗， 指望光明，卻行在幽暗中。
ISA|59|10|我們用手摸牆，好像盲人， 四處摸索，如同失明的人； 中午時我們絆倒，如在黃昏一樣， 在強壯的人中，我們好像死人一般。
ISA|59|11|我們全都咆哮如熊， 哀鳴如鴿子； 指望公平，卻得不著； 指望救恩，它卻遠離。
ISA|59|12|我們的過犯在你面前增加， 罪惡作證控告我們； 過犯與我們同在。 至於我們的罪孽，我們都知道：
ISA|59|13|就是悖逆，否認耶和華， 轉去不跟從我們的上帝， 口說欺壓和叛逆的話， 心懷謊言，隨即說出；
ISA|59|14|公平轉而退後， 公義站在遠處， 誠實仆倒在廣場上， 正直不得進入；
ISA|59|15|誠實少見， 離棄邪惡的人反成掠物。 那時，耶和華見沒有公平， 就不喜悅。
ISA|59|16|他見無人， 竟無一人代求，甚為詫異， 就用自己的膀臂拯救他， 以公義扶持他。
ISA|59|17|他穿上公義為鎧甲， 戴上救恩為頭盔， 穿上報復為衣服， 披戴熱心為外袍。
ISA|59|18|他必按人的行為報應， 惱怒他的敵人， 報復他的仇敵， 向眾海島施行報應。
ISA|59|19|在日落之處，人必敬畏耶和華的名； 在日出之地，人必敬畏他的榮耀。 他必如湍急的河流沖來， 耶和華的靈催逼他自己。
ISA|59|20|必有一位救贖主來到 錫安 ， 來到 雅各 族中離棄過犯的人那裏； 這是耶和華說的。
ISA|59|21|耶和華說：「這就是我與他們所立的約：我加給你的靈，傳給你的話，必不離你的口，也不離你後裔與你後裔之後裔的口，從今直到永遠；這是耶和華說的。」
ISA|60|1|興起，發光！因為你的光已來到！ 耶和華的榮光發出照耀著你。
ISA|60|2|看哪，黑暗籠罩大地， 幽暗遮蓋萬民， 耶和華卻要升起照耀你， 他的榮光要顯在你身上。
ISA|60|3|列國要來就你的光， 列王要來就你發出的光輝。
ISA|60|4|你舉目向四圍觀看， 眾人都聚集到你這裏。 你的兒子從遠方來， 你的女兒也被抱著帶來。
ISA|60|5|那時，你看見就有光榮， 你的心興奮歡暢 ； 因為大海那邊的財富必歸你， 列國的財寶也來歸你。
ISA|60|6|成群的駱駝， 並 米甸 和 以法 的獨峰駝遮滿你； 示巴 的眾人都必來到， 要奉上黃金和乳香， 又要傳揚讚美耶和華的話。
ISA|60|7|基達 的羊群都聚集到你這裏， 尼拜約 的公羊供你使用， 獻在我壇上蒙悅納； 我必榮耀我那榮耀的殿。
ISA|60|8|那些飛來如雲、 又像鴿子飛向窗戶的是誰呢？
ISA|60|9|眾海島必等候我 ， 他施 的船隻領先， 將你的兒女，連同他們的金銀從遠方帶來， 這都因 以色列 的聖者、耶和華－你上帝的名， 因為他已經榮耀了你。
ISA|60|10|外邦人要建造你的城牆， 他們的君王必服事你。 我曾發怒擊打你， 如今卻施恩憐憫你。
ISA|60|11|你的城門必時常開放， 晝夜不關， 使人將列國的財物帶來歸你， 他們的君王也被牽引而來。
ISA|60|12|不事奉你的那邦、那國要滅亡， 那些國家必全然荒廢。
ISA|60|13|黎巴嫩 的榮耀， 就是松樹、杉樹、黃楊樹， 都必一同歸你， 用以裝飾我聖所坐落之處； 我也要使我腳所踏之地得榮耀。
ISA|60|14|壓制你的，他的子孫必來向你屈身； 藐視你的，都要在你腳前下拜。 人要稱你為「耶和華的城」， 為「 以色列 聖者的 錫安 」。
ISA|60|15|你雖曾被拋棄，被恨惡， 甚至無人經過， 我卻使你有永遠的榮華， 成為世世代代的喜樂。
ISA|60|16|你要吃列國的奶， 吃列王的乳。 你就知道我－耶和華是你的救主， 是你的救贖主，是 雅各 的大能者。
ISA|60|17|我要賞賜金子代替銅， 賞賜銀子代替鐵， 銅代替木頭， 鐵代替石頭。 我要以和平為你的官長， 以公義為你的監督。
ISA|60|18|你的地不再聽聞殘暴的事， 境內不再聽見破壞與毀滅。 你必稱你的牆為「拯救」， 稱你的門為「讚美」。
ISA|60|19|白晝太陽不再作你的光， 月亮 也不再發光照耀你； 耶和華卻要作你永遠的光， 你的上帝要成為你的榮耀。
ISA|60|20|你的太陽不再落下， 月亮也不消失； 因為耶和華必作你永遠的光。 你悲哀的日子定要結束。
ISA|60|21|你的居民全是義人， 永遠得地為業； 他們是我栽的苗，是我手的工作， 為了彰顯我的榮耀。
ISA|60|22|稀少的要成為大族， 弱小的要變為強國。 我－耶和華到了時候必速速成就這事。
ISA|61|1|主耶和華的靈在我身上， 因為耶和華用膏膏我， 叫我報好信息給貧窮的人， 差遣我醫好傷心的人， 報告被擄的得釋放， 被捆綁的得自由；
ISA|61|2|宣告耶和華的恩年 和我們的上帝報仇的日子； 安慰所有悲哀的人，
ISA|61|3|為 錫安 悲哀的人，賜華冠代替灰燼， 喜樂的油代替悲哀， 讚美為衣代替憂傷的靈； 稱他們為「公義樹」， 是耶和華所栽植的，為要彰顯他的榮耀。
ISA|61|4|他們必修造久已荒涼的廢墟， 建立先前淒涼之處， 重修歷代荒涼之城。
ISA|61|5|那時，陌生人要伺候、牧放你們的羊群； 外邦人必為你們耕種田地， 修整你們的葡萄園。
ISA|61|6|但你們要稱為「耶和華的祭司」， 稱作「我們上帝的僕人」。 你們必享用列國的財物， 必承受他們的財富 。
ISA|61|7|因為他們所受雙倍的羞辱， 凌辱被稱為他們的命運， 因此，他們在境內必得雙倍的產業， 永遠之樂必歸給他們。
ISA|61|8|因為我－耶和華喜愛公平， 恨惡搶奪與惡行 ； 我要憑誠實施行報償， 與我的百姓立永約。
ISA|61|9|他們的後裔必在列國中為人所知， 他們的子孫在萬民中為人所識； 凡看見他們的必承認他們是耶和華所賜福的後裔。
ISA|61|10|我因耶和華大大歡喜， 我的心因上帝喜樂； 因他以拯救為衣給我穿上， 以公義為外袍給我披上， 好像新郎戴上華冠， 又如新娘佩戴首飾。
ISA|61|11|地怎樣使芽長出， 園子怎樣使所栽種的生長， 主耶和華也必照樣 使公義和讚美在萬國中發出。
ISA|62|1|我因 錫安 必不靜默， 為 耶路撒冷 必不安寧， 直到它的公義如光輝發出， 它的救恩如火把燃燒。
ISA|62|2|列國要看見你的公義， 列王要看見你的榮耀。 你必得新的名字， 是耶和華親口起的。
ISA|62|3|你在耶和華的手中成為華冠， 在你上帝的掌上成為冠冕。
ISA|62|4|你不再稱為「被撇棄的」， 你的地也不再稱為「荒蕪的」； 你要稱為「我所喜悅的」， 你的地要稱為「有歸屬的」。 因為耶和華喜悅你， 你的地必歸屬於他。
ISA|62|5|年輕人怎樣娶童女， 你的百姓也要照樣娶你； 新郎怎樣因新娘而喜樂， 你的上帝也要如此以你為樂。
ISA|62|6|耶路撒冷 啊， 我在你城牆上設立守望者， 他們晝夜不停地呼喊。 呼求耶和華的啊，你們不要歇息，
ISA|62|7|也不要使他歇息， 直等他建立 耶路撒冷 ， 使 耶路撒冷 在地上為人所讚美。
ISA|62|8|耶和華指著自己的右手和大能的膀臂起誓說： 「我必不再將你的五穀給仇敵作食物， 外邦人也必不再喝你勞碌得來的新酒。
ISA|62|9|惟有那收割的要吃，並讚美耶和華； 那儲藏葡萄的要在我聖所院內喝。」
ISA|62|10|你們當從門經過，經過， 預備百姓的路。 你們要修築，修築大道， 清除石頭， 為萬民豎立大旗。
ISA|62|11|看哪，耶和華曾宣告到地極， 你們要對 錫安 說： 「看哪，你的拯救者已來到。 看哪，他的賞賜在他那裏， 他的報償在他面前。」
ISA|62|12|人稱他們為「聖民」，為「耶和華救贖的民」， 你也必稱為「受眷顧的」，為「不被撇棄的城」。
ISA|63|1|這從 以東 的 波斯拉 來， 穿紅衣服， 裝扮華美， 能力廣大， 大步向前邁進的是誰呢？ 就是我， 憑公義說話， 以大能施行拯救的。
ISA|63|2|你為何以紅色裝扮？ 你的衣服為何像踹醡酒池的人呢？
ISA|63|3|我獨自踹醡酒池， 萬民中並無一人與我同在。 我發怒，將他們踹下， 發烈怒將他們踐踏。 他們的血濺在我的衣服上， 玷污了我一切的衣裳。
ISA|63|4|因為報仇之日在我心中， 救贖我民之年已經來到。
ISA|63|5|我仰望，見無人幫助； 我詫異，竟無人扶持。 因此，我的膀臂為我施行拯救； 我的烈怒將我扶持。
ISA|63|6|我發怒，踹下眾民； 發烈怒，使他們喝醉， 又將他們的血倒在地上。
ISA|63|7|我要照耶和華一切所賜給我們的， 並他憑憐憫與豐盛的慈愛 所賜給 以色列 家的大恩， 述說他的慈愛和美德。
ISA|63|8|他說：「他們誠然是我的百姓， 未行虛假的子民。」 這樣，他就作了他們的救主。
ISA|63|9|他們在一切苦難當中， 他也同受苦難， 並且他面前的使者拯救他們 。 他以慈愛和憐憫救贖他們， 在古時的日子時常抱他們，背他們。
ISA|63|10|他們竟然悖逆，使他的聖靈憂傷。 他就轉變，成為他們的仇敵， 親自攻擊他們。
ISA|63|11|那時，他的百姓想起古時 摩西 的日子： 「那將百姓和牧養群羊的人 從海裏領上來的在哪裏呢？ 那將聖靈降在他們中間，
ISA|63|12|以榮耀的膀臂在 摩西 右邊行動， 在百姓面前將水分開， 為要建立自己永遠的名，
ISA|63|13|又帶領他們經過深處的在哪裏呢？」 他們如馬行走曠野，不致絆跌；
ISA|63|14|又如牲畜下到山谷， 耶和華的靈使他們得安息； 照樣，你也引導你的百姓， 為要建立自己榮耀的名。
ISA|63|15|求你從天上， 從你神聖榮耀的居所垂顧觀看。 你的熱心和你大能的作為在哪裏呢？ 你內心的關懷和你的憐憫向我們停止了。
ISA|63|16|亞伯拉罕 雖然不承認我們， 以色列 也不承認我們， 你卻是我們的父。 耶和華啊，你是我們的父； 自古以來，你的名是「我們的救贖主」。
ISA|63|17|耶和華啊，你為何使我們偏離你的道， 使我們心裏剛硬、不敬畏你呢？ 求你為你的僕人， 為你產業的支派而回轉。
ISA|63|18|你的聖民暫時得你的聖所， 但我們的敵人踐踏了它。
ISA|63|19|我們就成了你未曾治理的人， 成了未曾稱為你名下的人。
ISA|64|1|願你破天而降， 願山在你面前震動，
ISA|64|2|好像火燒乾柴， 又如火將水燒開， 使你敵人知道你的名， 列國必在你面前發顫！
ISA|64|3|你曾做我們不能逆料可畏的事； 那時你降臨，山嶺在你面前震動。
ISA|64|4|自古以來，人未曾聽見，未曾耳聞，未曾眼見， 除你以外，還有上帝能為等候他的人行事。
ISA|64|5|你迎見那歡喜行義、記念你道的人； 看哪，你曾發怒，因我們犯了罪； 這景況已久，我們還能得救嗎？
ISA|64|6|我們都如不潔淨的人， 所行的義都像污穢的衣服。 我們如葉子漸漸枯乾， 罪孽像風把我們吹走。
ISA|64|7|無人求告你的名， 無人奮力抓住你。 你轉臉不顧我們， 你使我們因罪孽而融化 。
ISA|64|8|但耶和華啊，現在你仍是我們的父！ 我們是泥，你是陶匠； 我們都是你親手所造的。
ISA|64|9|耶和華啊，求你不要大發震怒， 也不要永遠記得罪孽； 看哪，求你垂顧我們， 因我們都是你的百姓。
ISA|64|10|你的聖城已變為曠野； 錫安 變為曠野， 耶路撒冷 成為廢墟。
ISA|64|11|我們那神聖華美的殿， 就是我們祖先讚美你的地方，已被火焚燒； 我們所羨慕的美地盡都荒蕪。
ISA|64|12|耶和華啊，有這些事，你還能忍受嗎？ 你還靜默，使我們大受苦難嗎？
ISA|65|1|沒有求問我的，我要讓他們找到； 沒有尋找我的，我要讓他們尋見； 我對沒有呼求我名的國 說： 「我在這裏！我在這裏！」
ISA|65|2|我整天向那悖逆的百姓招手， 他們隨自己的意念行不善之道。
ISA|65|3|這百姓時常當面惹我發怒， 在園中獻祭， 在磚上燒香，
ISA|65|4|在墳墓間停留， 在隱密處過夜， 吃豬肉， 器皿中有不潔淨之肉熬的湯；
ISA|65|5|且對人說：「你站開吧！ 不要挨近我，因為我對你來說太神聖了 。」 這些人惹我鼻中冒煙， 如終日燃燒的火。
ISA|65|6|看哪，這些都寫在我面前。 我必不靜默，卻要施行報應， 將你們和你們祖先的罪孽 全都報應在後人身上； 因為他們在山上燒香， 在岡上褻瀆我， 我要按他們先前所行的，報應在他們身上 ； 這是耶和華說的。
ISA|65|7|
ISA|65|8|耶和華如此說： 「人在葡萄中尋得新酒時會說： 『不要毀壞它，因為它還有用處』； 同樣，我必因我僕人的緣故， 不將他們全然毀滅。
ISA|65|9|我必從 雅各 中領出後裔， 從 猶大 中領出那要繼承我眾山的； 我的選民要繼承它， 我的僕人要在那裏居住。
ISA|65|10|沙崙 必成為羊群的圈， 亞割谷 成為牛群躺臥之處， 都為尋求我的民所得。
ISA|65|11|但你們這些離棄耶和華， 就是忘記我的聖山、 為『幸運之神』擺設筵席、 為『命運之神』裝滿調和酒的，
ISA|65|12|我命定你們歸於刀下， 你們都要屈身被殺； 因為我呼喚，你們不回應； 我說話，你們不聽從； 反倒做我眼中看為惡的事， 選擇我所不喜悅的事。」
ISA|65|13|所以，主耶和華如此說： 「看哪，我的僕人必得吃，你們卻飢餓； 看哪，我的僕人必得喝，你們卻乾渴； 看哪，我的僕人必歡喜，你們卻蒙羞。
ISA|65|14|看哪，我的僕人因心中喜樂而歡呼， 你們卻因心裏悲痛而哀哭， 因靈裏憂傷而哀號。
ISA|65|15|你們必留下自己的名 給我選民指著賭咒： 主耶和華必殺你們， 另起別名稱呼他的僕人。
ISA|65|16|在地上為自己求福的， 必憑真實的上帝求福； 在地上起誓的， 必指著真實的上帝起誓。 因為從前的患難已被遺忘， 從我眼前消逝。」
ISA|65|17|「看哪，我造新天新地！ 從前的事不再被記念，也不被人放在心上；
ISA|65|18|當因我所造的歡喜快樂，直到永遠； 看哪，因為我造 耶路撒冷 為人所喜， 造其中的居民為人所樂。
ISA|65|19|我必因 耶路撒冷 歡喜， 因我的百姓快樂， 那裏不再聽見哭泣和哀號的聲音。
ISA|65|20|那裏沒有數日夭折的嬰孩， 也沒有壽數不滿的老人； 因為百歲死的仍算孩童， 未達百歲而亡的 算是被詛咒的。
ISA|65|21|他們建造房屋，居住其中， 栽葡萄園，吃園中的果子；
ISA|65|22|並非造了給別人居住， 也非栽種給別人享用； 因為我百姓的日子必長久如樹木， 我的選民必享受親手勞碌得來的。
ISA|65|23|他們必不徒然勞碌， 所生產的，也不遭災害， 因為他們和他們的子孫 都是蒙耶和華賜福的後裔。
ISA|65|24|他們尚未求告，我就應允； 正說話的時候，我就垂聽。
ISA|65|25|野狼必與羔羊同食， 獅子必吃草，與牛一樣， 蛇必以塵土為食物； 在我聖山的遍處， 牠們都不傷人，也不害物； 這是耶和華說的。」
ISA|66|1|耶和華如此說： 「天是我的座位； 地是我的腳凳。 你們能為我造怎樣的殿宇呢？ 哪裏是我安歇的地方呢？
ISA|66|2|這一切是我手所造的， 這一切就都存在了。 我所看顧的是困苦、靈裏痛悔、 因我言語而戰兢的人。 這是耶和華說的。
ISA|66|3|「至於那些宰牛，殺人， 獻羔羊，打斷狗頸項， 獻豬血為供物， 燒乳香，稱頌偶像的， 他們選擇自己的道路， 心裏喜愛可憎惡的事；
ISA|66|4|我也必選擇苦待他們， 使他們所懼怕的臨到他們； 因為我呼喚，無人回應； 我說話，他們不聽從； 反倒做我眼中看為惡的事， 選擇我所不喜悅的事。」
ISA|66|5|你們因耶和華言語而戰兢的人哪，當聽他的話： 「你們的弟兄，就是恨惡你們， 因我名趕出你們的，曾說： 『願耶和華彰顯榮耀 ， 好讓我們看見你們的喜樂。』 但蒙羞的終究是他們！
ISA|66|6|「有喧嘩的聲音出自城中！ 有聲音來自殿裏！ 是耶和華向仇敵施行報應的聲音！
ISA|66|7|「 錫安 未曾陣痛就生產， 疼痛尚未來到，就生出男孩。
ISA|66|8|國豈能一日而生？ 民豈能一時而產？ 但 錫安 一陣痛就生下兒女， 這樣的事有誰聽見， 有誰看見呢？
ISA|66|9|耶和華說：我使人臨產， 豈不讓她 生產呢？ 你的上帝說：我使人生產， 難道還讓她關閉 不生嗎？
ISA|66|10|「你們所有愛慕 耶路撒冷 的啊， 要與她一同歡喜，為她高興； 你們所有為她悲哀的啊， 都要與她一同樂上加樂；
ISA|66|11|使你們在她安慰的懷中吃奶得飽， 盡情吸取她豐盛的榮耀，滿心喜樂。」
ISA|66|12|耶和華如此說： 「看哪，我要使平安臨到她，好像江河； 使列國的榮耀及於她，如同漲溢的溪流。 你們要盡情吸吮； 你們必被抱在身旁 ，搖弄在膝上。
ISA|66|13|我要安慰你們，如同母親安慰兒女； 你們也必在 耶路撒冷 得安慰。
ISA|66|14|你們看見，心裏就喜樂， 你們的骨頭必如草生長； 耶和華的手在他僕人身上彰顯， 他卻要向他的仇敵發怒。」
ISA|66|15|看哪，耶和華必在火中降臨， 他的戰車宛如暴風， 以烈怒施行報應， 以火焰施行責罰；
ISA|66|16|耶和華必以火與刀審判凡有血肉之軀的， 被耶和華所殺的很多。
ISA|66|17|那些潔淨自己獻給偶像，進入園內，跟隨其中一個人去吃豬肉和鼠肉，並可憎之物的，他們必一同滅絕。這是耶和華說的。
ISA|66|18|我知道他們的行為和他們的意念。聚集萬國萬族 的時候到了 ，他們要來瞻仰我的榮耀；
ISA|66|19|我要在他們中間顯神蹟，差遣他們當中的倖存者到列國去，就是到 他施 、 普勒 、以善射聞名的 路德 、 土巴 、 雅完 ，和未曾聽見我名聲，未曾看見我榮耀的遙遠海島那裏去；他們必在列國中傳揚我的榮耀。
ISA|66|20|他們要將你們的弟兄從列國中帶回，或騎馬，或坐車，或乘蓬車，或騎騾子，或騎獨峰駝，到我的聖山 耶路撒冷 ，作為供物獻給耶和華。這是耶和華說的。正如 以色列 人用潔淨的器皿盛供物奉到耶和華的殿中，
ISA|66|21|我也必從他們中間立人作祭司，作 利未 人。這是耶和華說的。
ISA|66|22|「我所造的新天新地在我面前長存， 你們的後裔和你們的名號也必照樣長存。 這是耶和華說的。
ISA|66|23|每逢初一、安息日， 凡有血肉之軀的必前來，在我面前下拜； 這是耶和華說的。
ISA|66|24|「他們要出去觀看那些違背我的人的屍首， 他們的蟲是不死的， 他們的火是不滅的， 凡有血肉之軀的都必憎惡他們。」
