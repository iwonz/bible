2CHR|1|1|И утвердился Соломон, сын Давидов, в царстве своем; и Господь Бог его [был] с ним, и вознес его высоко.
2CHR|1|2|И приказал Соломон [собраться] всему Израилю: тысяченачальникам и стоначальникам, и судьям, и всем начальствующим во всем Израиле – главам поколений.
2CHR|1|3|И пошли Соломон и все собрание с ним на высоту, что в Гаваоне, ибо там была Божия скиния собрания, которую устроил Моисей, раб Господень, в пустыне.
2CHR|1|4|Ковчег Божий принес Давид из Кириаф–Иарима на место, которое приготовил для него Давид, устроив для него скинию в Иерусалиме.
2CHR|1|5|А медный жертвенник, который сделал Веселеил, сын Урия, сына Орова, [оставался] там, пред скиниею Господнею, и взыскал его Соломон с собранием.
2CHR|1|6|И там пред лицем Господа, на медном жертвеннике, который пред скиниею собрания, вознес Соломон тысячу всесожжений.
2CHR|1|7|В ту ночь явился Бог Соломону и сказал ему: проси, что Мне дать тебе.
2CHR|1|8|И сказал Соломон Богу: Ты сотворил Давиду, отцу моему, великую милость и поставил меня царем вместо него.
2CHR|1|9|Да исполнится же, Господи Боже, слово Твое к Давиду, отцу моему. Так как Ты воцарил меня над народом многочисленным, как прах земной,
2CHR|1|10|то ныне дай мне премудрость и знание, чтобы я [умел] выходить пред народом сим и входить, ибо кто может управлять сим народом Твоим великим?
2CHR|1|11|И сказал Бог Соломону: за то, что это было на сердце твоем, и ты не просил богатства, имения и славы и души неприятелей твоих, и также не просил ты многих дней, а просил себе премудрости и знания, чтобы управлять народом Моим, над которым Я воцарил тебя,
2CHR|1|12|премудрость и знание дается тебе, а богатство и имение и славу Я дам тебе такие, подобных которым не бывало у царей прежде тебя и не будет после тебя.
2CHR|1|13|И пришел Соломон с высоты, что в Гаваоне, от скинии собрания, в Иерусалим и царствовал над Израилем.
2CHR|1|14|И набрал Соломон колесниц и всадников; и было у него тысяча четыреста колесниц и двенадцать тысяч всадников; и он разместил их в колесничных городах и при царе в Иерусалиме.
2CHR|1|15|И сделал царь серебро и золото в Иерусалиме равноценным [простому] камню, а кедры, по множеству их, сделал равноценными сикоморам, которые на низких местах.
2CHR|1|16|Коней Соломону приводили из Египта и из Кувы; купцы царские из Кувы получали их за деньги.
2CHR|1|17|Колесница получаема и доставляема была из Египта за шестьсот [сиклей] серебра, а конь за сто пятьдесят. Таким же образом они руками своими доставляли [это] всем царям Хеттейским и царям Арамейским.
2CHR|1|18|И положил Соломон построить дом имени Господню и дом царский для себя.
2CHR|2|1|И отчислил Соломон семьдесят тысяч носильщиков и восемьдесят тысяч каменосеков в горах, и надзирателей над ними три тысячи шестьсот.
2CHR|2|2|И послал Соломон к Хираму, царю Тирскому, сказать: как поступал ты с Давидом, отцом моим, и присылал ему кедры на построение дома для его жительства, [так поступи и со мною].
2CHR|2|3|Вот я строю дом имени Господа Бога моего, для посвящения Ему, чтобы возжигать пред Ним благовонное курение, представлять постоянно хлебы предложения и [возносить там] всесожжения утром и вечером в субботы, и в новомесячия, и в праздники Господа Бога нашего, что навсегда заповедано Израилю.
2CHR|2|4|И дом, который я строю, велик, потому что велик Бог наш, выше всех богов.
2CHR|2|5|И достанет ли у кого силы построить Ему дом, когда небо и небеса небес не вмещают Его? И кто я, чтобы мог построить Ему дом? Разве [только] для курения пред лицем Его.
2CHR|2|6|Итак пришли мне человека, умеющего делать [изделия] из золота, и из серебра, и из меди, и из железа, и из [пряжи] пурпурового, багряного и яхонтового [цвета], и знающего вырезывать резную работу, вместе с художниками, какие есть у меня в Иудее и в Иерусалиме, которых приготовил Давид, отец мой.
2CHR|2|7|И пришли мне кедровых дерев, и кипарису и певгового дерева с Ливана, ибо я знаю, что рабы твои умеют рубить дерева Ливанские. И вот рабы мои пойдут с рабами твоими,
2CHR|2|8|чтобы мне приготовить множество дерев, потому что дом, который я строю, великий и чудный.
2CHR|2|9|И вот древосекам, рубящим дерева, рабам твоим, я даю в пищу: пшеницы двадцать тысяч коров, и ячменю двадцать тысяч коров, и вина двадцать тысяч батов, и оливкового масла двадцать тысяч батов.
2CHR|2|10|И отвечал Хирам, царь Тирский, письмом, которое прислал к Соломону: по любви к народу Своему, Господь поставил тебя царем над ним.
2CHR|2|11|И [еще] сказал Хирам: благословен Господь Бог Израилев, создавший небо и землю, давший царю Давиду сына мудрого, имеющего смысл и разум, который намерен строить дом Господу и дом царский для себя.
2CHR|2|12|Итак я посылаю [тебе] человека умного, имеющего знания, Хирам–Авия,
2CHR|2|13|сына [одной] женщины из дочерей Дановых, – а отец его Тирянин, – умеющего делать [изделия] из золота и из серебра, из меди, из железа, из камней и из дерев, из [пряжи] пурпурового, яхонтового [цвета], и из виссона, и из багряницы, и вырезывать всякую резьбу, и исполнять все, что будет поручено ему вместе с художниками твоими и с художниками господина моего Давида, отца твоего.
2CHR|2|14|А пшеницу и ячмень, оливковое масло и вино, о которых говорил ты, господин мой, пошли рабам твоим.
2CHR|2|15|Мы же нарубим дерев с Ливана, сколько нужно тебе, и пригоним их в плотах по морю в Яфу, а ты отвезешь их в Иерусалим.
2CHR|2|16|И исчислил Соломон всех пришельцев, бывших [тогда] в земле Израилевой, после исчисления их, сделанного Давидом, отцом его, – и нашлось их сто пятьдесят три тысячи шестьсот.
2CHR|2|17|И сделал он из них семьдесят тысяч носильщиков и восемьдесят тысяч каменосеков на горах и три тысячи шестьсот надзирателей, чтобы они побуждали народ к работе.
2CHR|3|1|И начал Соломон строить дом Господень в Иерусалиме на горе Мориа, которая указана была Давиду, отцу его, на месте, которое приготовил Давид, на гумне Орны Иевусеянина.
2CHR|3|2|Начал же он строить во второй [день] второго месяца, в четвертый год царствования своего.
2CHR|3|3|И вот основание, [положенное] Соломоном при строении дома Божия: длина [его] шестьдесят локтей, по прежней мере, а ширина двадцать локтей;
2CHR|3|4|и притвор, который пред домом, длиною по ширине дома в двадцать локтей, а вышиною во сто двадцать. И обложил его внутри чистым золотом.
2CHR|3|5|Дом же главный обшил деревом кипарисовым и обложил его лучшим золотом, и выделал на нем пальмы и цепочки.
2CHR|3|6|И обложил дом дорогими камнями для красоты; золото же [было] золото Парваимское.
2CHR|3|7|И покрыл дом, бревна, пороги и стены его и двери его золотом, и вырезал на стенах херувимов.
2CHR|3|8|И сделал Святое Святых: длина его по широте дома в двадцать локтей, и ширина его в двадцать локтей; и покрыл его лучшим золотом на шестьсот талантов.
2CHR|3|9|В гвоздях весу до пятидесяти сиклей золота. Горницы также покрыл золотом.
2CHR|3|10|И сделал он во Святом Святых двух херувимов резной работы и покрыл их золотом.
2CHR|3|11|Крылья херувимов длиною [были] в двадцать локтей. Одно крыло в пять локтей касалось стены дома, а другое крыло в пять же локтей сходилось с крылом другого херувима;
2CHR|3|12|[равно] и крыло другого херувима в пять локтей касалось стены дома, а другое крыло в пять локтей сходилось с крылом другого херувима.
2CHR|3|13|Крылья сих херувимов [были] распростерты на двадцать локтей; и они стояли на ногах своих, лицами своими к храму.
2CHR|3|14|И сделал завесу из яхонтовой, пурпуровой и багряной [ткани] и из виссона и изобразил на ней херувимов.
2CHR|3|15|И сделал пред храмом два столба, длиною по тридцати пяти локтей, и капитель на верху каждого в пять локтей.
2CHR|3|16|И сделал цепочки, [как] во святилище, и положил на верху столбов, и сделал сто гранатовых яблок и положил на цепочки.
2CHR|3|17|И поставил столбы пред храмом, один по правую сторону, другой по левую, и дал имя правому Иахин, а левому имя Воаз.
2CHR|4|1|И сделал медный жертвенник: двадцать локтей длина его и двадцать локтей ширина его и десять локтей вышина его.
2CHR|4|2|И сделал море литое, – от края его до края его десять локтей, – все круглое, вышиною в пять локтей; и снурок в тридцать локтей обнимал его кругом;
2CHR|4|3|и [литые] подобия волов стояли под ним кругом со всех сторон; на десять локтей окружали море кругом два ряда волов, вылитых одним литьем с ним.
2CHR|4|4|Стояло оно на двенадцати волах: три глядели к северу и три глядели к западу, и три глядели к югу, и три глядели к востоку, – и море на них сверху; зады же их были обращены внутрь под него.
2CHR|4|5|Толщиною оно [было] в ладонь; и края его, сделанные, как края чаши, [походили] на распустившуюся лилию. Оно вмещало до трех тысяч батов.
2CHR|4|6|И сделал десять омывальниц, и поставил пять по правую сторону и пять по левую, чтоб омывать в них, – приготовляемое ко всесожжению омывали в них; море же – для священников, чтоб они омывались в нем.
2CHR|4|7|И сделал десять золотых светильников, как им быть надлежало, и поставил в храме, пять по правую сторону и пять по левую.
2CHR|4|8|И сделал десять столов и поставил в храме, пять по правую сторону и пять по левую, и сделал сто золотых чаш.
2CHR|4|9|И сделал священнический двор и большой двор и двери к двору, и вереи их обложил медью.
2CHR|4|10|Море поставил на правой стороне, к юго–востоку.
2CHR|4|11|И сделал Хирам тазы, и лопатки, и чаши. И кончил Хирам работу, которую производил для царя Соломона в доме Божием:
2CHR|4|12|два столба и две опояски венцов на верху столбов, и две сетки для покрытия двух опоясок венцов, которые на главе столбов,
2CHR|4|13|и четыреста гранатовых яблок на двух сетках, два ряда гранатовых яблок для каждой сетки, для покрытия двух опоясок венцов, которые на столбах.
2CHR|4|14|И подставы сделал он, и омывальницы сделал на подставах;
2CHR|4|15|одно море, и двенадцать волов под ним,
2CHR|4|16|и тазы, и лопатки, и вилки, и весь прибор их сделал Хирам–Авий царю Соломону для дома Господня из полированной меди.
2CHR|4|17|В окрестности Иордана выливал их царь, в глинистой земле, между Сокхофом и Цередою.
2CHR|4|18|И сделал Соломон все вещи сии в великом множестве, так что не знали веса меди.
2CHR|4|19|Также сделал Соломон все вещи для дома Божия и золотой жертвенник, и столы, на которых хлебы предложения,
2CHR|4|20|и светильники и лампады их, чтобы возжигать их по уставу пред давиром, из чистого золота;
2CHR|4|21|и цветы, и лампады, и щипцы из золота, из самого чистого золота,
2CHR|4|22|и ножи, и кропильницы, и чаши, и лотки из золота самого чистого, и двери храма, – двери его внутренние во Святое Святых, и двери храма во святилище, – из золота.
2CHR|5|1|И окончилась вся работа, которую производил Соломон для дома Господня. И принес Соломон посвященное Давидом, отцом его, и серебро и золото и все вещи отдал в сокровищницы дома Божия.
2CHR|5|2|Тогда собрал Соломон старейшин Израилевых и всех глав колен, начальников поколений сынов Израилевых, в Иерусалим, для перенесения ковчега завета Господня из города Давидова, то есть [с] Сиона.
2CHR|5|3|И собрались к царю все Израильтяне на праздник, в седьмой месяц.
2CHR|5|4|И пришли все старейшины Израилевы. Левиты взяли ковчег
2CHR|5|5|и понесли ковчег и скинию собрания и все вещи священные, которые в скинии, – понесли их священники и левиты.
2CHR|5|6|Царь же Соломон и все общество Израилево, собравшееся к нему пред ковчегом, приносили жертвы из овец и волов, которых невозможно исчислить и определить, по причине множества.
2CHR|5|7|И принесли священники ковчег завета Господня на место его, в давир храма – во Святое Святых, под крылья херувимов.
2CHR|5|8|И херувимы распростирали крылья над местом ковчега, и покрывали херувимы ковчег и шесты его сверху.
2CHR|5|9|И выдвинулись шесты, так что головки шестов ковчега видны были пред давиром, но не выказывались наружу, и они там до сего дня.
2CHR|5|10|Не было в ковчеге ничего кроме двух скрижалей, которые положил Моисей на Хориве, когда Господь заключил [завет] с сынами Израилевыми, по исходе их из Египта.
2CHR|5|11|Когда священники вышли из святилища, ибо все священники, находившиеся там, освятились без различия отделов;
2CHR|5|12|и левиты певцы, – все они, [то есть] Асаф, Еман, Идифун и сыновья их, и братья их, – одетые в виссон, с кимвалами и с псалтирями и цитрами стояли на восточной стороне жертвенника, и с ними сто двадцать священников, трубивших трубами,
2CHR|5|13|и были, как один, трубящие и поющие, издавая один голос к восхвалению и славословию Господа; и когда загремел звук труб и кимвалов и музыкальных орудий, и восхваляли Господа, ибо Он благ, ибо вовек милость Его; тогда дом, дом Господень, наполнило облако,
2CHR|5|14|и не могли священники стоять на служении по причине облака, потому что слава Господня наполнила дом Божий.
2CHR|6|1|Тогда сказал Соломон: Господь сказал, что Он благоволит обитать во мгле,
2CHR|6|2|а я построил дом в жилище Тебе, место для вечного Твоего пребывания.
2CHR|6|3|И обратился царь лицем своим и благословил все собрание Израильтян, – все собрание Израильтян стояло, –
2CHR|6|4|и сказал: благословен Господь Бог Израилев, Который, что сказал устами Своими Давиду, отцу моему, исполнил [ныне] рукою Своею! Он говорил:
2CHR|6|5|"с того дня, как Я вывел народ Мой из земли Египетской, Я не избрал города ни в одном из колен Израилевых для построения дома, в котором пребывало бы имя Мое, и не избрал человека, который был бы правителем народа Моего Израиля,
2CHR|6|6|но избрал Иерусалим, чтобы там пребывало имя Мое, и избрал Давида, чтоб он был над народом Моим Израилем".
2CHR|6|7|И было на сердце у Давида, отца моего, построить дом имени Господа, Бога Израилева.
2CHR|6|8|Но Господь сказал Давиду, отцу моему: "у тебя есть на сердце построить храм имени Моему; хорошо, что это на сердце у тебя.
2CHR|6|9|Однако не ты построишь храм, а сын твой, который произойдет из чресл твоих, – он построит храм имени Моему".
2CHR|6|10|И исполнил Господь слово Свое, которое изрек: я вступил на место Давида, отца моего, и воссел на престоле Израилевом, как сказал Господь, и построил дом имени Господа Бога Израилева.
2CHR|6|11|И я поставил там ковчег, в котором завет Господа, заключенный Им с сынами Израилевыми.
2CHR|6|12|И стал [Соломон] у жертвенника Господня впереди всего собрания Израильтян, и воздвиг руки свои, –
2CHR|6|13|ибо Соломон сделал медный амвон длиною в пять локтей и шириною в пять локтей, а вышиною в три локтя, и поставил его среди двора; и стал на нем, и преклонил колени впереди всего собрания Израильтян, и воздвиг руки свои к небу, –
2CHR|6|14|и сказал: Господи Боже Израилев! Нет Бога, подобного Тебе, ни на небе, ни на земле. Ты хранишь завет и милость к рабам Твоим, ходящим пред Тобою всем сердцем своим:
2CHR|6|15|Ты исполнил рабу Твоему Давиду, отцу моему, что Ты говорил ему; что изрек Ты устами Твоими, то в день сей исполнил рукою Твоею.
2CHR|6|16|И ныне, Господи Боже Израилев! исполни рабу Твоему Давиду, отцу моему, то, что Ты сказал ему, говоря: не прекратится у тебя [муж], сидящий пред лицем Моим на престоле Израилевом, если только сыновья твои будут наблюдать за путями своими, ходя по закону Моему так, как ты ходил предо Мною.
2CHR|6|17|И ныне, Господи Боже Израилев! да будет верно слово Твое, которое Ты изрек рабу Твоему Давиду.
2CHR|6|18|Поистине, Богу ли жить с человеками на земле? Если небо и небеса небес не вмещают Тебя, тем менее храм сей, который построил я.
2CHR|6|19|Но призри на молитву раба Твоего и на прошение его, Господи Боже мой! услышь воззвание и молитву, которою раб Твой молится пред Тобою.
2CHR|6|20|Да будут очи Твои отверсты на храм сей днем и ночью, на место, где Ты обещал положить имя Твое, чтобы слышать молитву, которою раб Твой будет молиться на месте сем.
2CHR|6|21|Услышь моления раба Твоего и народа Твоего Израиля, какими они будут молиться на месте сем; услышь с места обитания Твоего, с небес, услышь и помилуй!
2CHR|6|22|Когда кто согрешит против ближнего своего, и потребуют от него клятвы, чтоб он поклялся, и будет совершаться клятва пред жертвенником Твоим в храме сем,
2CHR|6|23|тогда Ты услышь с неба и соверши суд над рабами Твоими, воздай виновному, возложив поступок его на голову его, и оправдай правого, воздав ему по правде его.
2CHR|6|24|Когда поражен будет народ Твой Израиль неприятелем за то, что согрешил пред Тобою, и они обратятся [к Тебе], и исповедают имя Твое, и будут просить и молиться пред Тобою в храме сем,
2CHR|6|25|тогда Ты услышь с неба, и прости грех народа Твоего Израиля, и возврати их в землю, которую Ты дал им и отцам их.
2CHR|6|26|Когда заключится небо и не будет дождя за то, что они согрешили пред Тобою, и будут молиться на месте сем, и исповедают имя Твое, и обратятся от греха своего, потому что Ты смирил их,
2CHR|6|27|тогда Ты услышь с неба и прости грех рабов Твоих и народа Твоего Израиля, указав им добрый путь, по которому идти им, и пошли дождь на землю Твою, которую Ты дал народу Твоему в наследие.
2CHR|6|28|Голод ли будет на земле, будет ли язва моровая, будет ли ветер палящий или ржа, саранча или червь, будут ли теснить его неприятели его на земле владений его, [будет ли] какое бедствие, какая болезнь,
2CHR|6|29|всякую молитву, всякое прошение, какое будет от какого–либо человека или от всего народа Твоего Израиля, когда они почувствуют каждый бедствие свое и горе свое и прострут руки свои к храму сему,
2CHR|6|30|Ты услышь с неба – места обитания Твоего, и прости, и воздай каждому по всем путям его, как Ты знаешь сердце его, – ибо Ты один знаешь сердце сынов человеческих, –
2CHR|6|31|чтобы они боялись Тебя и ходили путями Твоими во все дни, доколе живут на земле, которую Ты дал отцам нашим.
2CHR|6|32|Даже и иноплеменник, который не от народа Твоего Израиля, когда он придет из земли далекой ради имени Твоего великого и руки Твоей могущественной и мышцы Твоей простертой, и придет и будет молиться у храма сего,
2CHR|6|33|Ты услышь с неба, с места обитания Твоего, и сделай все, о чем будет взывать к Тебе иноплеменник, чтобы все народы земли узнали имя Твое, и чтобы боялись Тебя, как народ Твой Израиль, и знали, что Твоим именем называется дом сей, который построил я.
2CHR|6|34|Когда выйдет народ Твой на войну против неприятелей своих путем, которым Ты пошлешь его, и будет молиться Тебе, обратившись к городу сему, который избрал Ты, и к храму, который я построил имени Твоему,
2CHR|6|35|тогда услышь с неба молитву их и прошение их и сделай, что потребно для них.
2CHR|6|36|Когда они согрешат пред Тобою, – ибо нет человека, который не согрешил бы, – и Ты прогневаешься на них, и предашь их врагу, и отведут их пленившие их в землю далекую или близкую,
2CHR|6|37|и когда они в земле, в которую будут пленены, войдут в себя и обратятся и будут молиться Тебе в земле пленения своего, говоря: мы согрешили, сделали беззаконие, мы виновны,
2CHR|6|38|и обратятся к Тебе всем сердцем своим и всею душею своею в земле пленения своего, куда отведут их в плен, и будут молиться, обратившись к земле своей, которую Ты дал отцам их, и к городу, который избрал Ты, и к храму, который я построил имени Твоему, –
2CHR|6|39|тогда услышь с неба, с места обитания Твоего, молитву их и прошение их, и сделай, что потребно для них, и прости народу Твоему, в чем он согрешил пред Тобою.
2CHR|6|40|Боже мой! да будут очи Твои отверсты и уши Твои внимательны к молитве на месте сем.
2CHR|6|41|И ныне, Господи Боже, стань на [место] покоя Твоего, Ты и ковчег могущества Твоего. Священники Твои, Господи Боже, да облекутся во спасение, и преподобные Твои да насладятся благами.
2CHR|6|42|Господи Боже! не отврати лица помазанника Твоего, помяни милости к Давиду, рабу Твоему.
2CHR|7|1|Когда окончил Соломон молитву, сошел огонь с неба и поглотил всесожжение и жертвы, и слава Господня наполнила дом.
2CHR|7|2|И не могли священники войти в дом Господень, потому что слава Господня наполнила дом Господень.
2CHR|7|3|И все сыны Израилевы, видя, как сошел огонь и слава Господня на дом, пали лицем на землю, на помост, и поклонились, и славословили Господа, ибо Он благ, ибо вовек милость Его.
2CHR|7|4|Царь же и весь народ стали приносить жертвы пред лицем Господа.
2CHR|7|5|И принес царь Соломон в жертву двадцать две тысячи волов и сто двадцать тысяч овец: так освятили дом Божий царь и весь народ.
2CHR|7|6|Священники стояли в служении своем, и левиты с музыкальными орудиями Господа, которые сделал царь Давид для прославления Господа, ибо вечна милость Его, так как Давид славословил чрез них; священники же трубили перед ним, и весь Израиль стоял.
2CHR|7|7|Освятил Соломон и внутреннюю часть двора, которая пред домом Господним: ибо принес там всесожжения и тук мирных жертв, так как жертвенник медный, сделанный Соломоном, не мог вмещать всесожжения и хлебного приношения, и туков.
2CHR|7|8|И сделал Соломон в то время семидневный праздник, и весь Израиль с ним – собрание весьма большое, [сошедшееся] от входа в Емаф до реки Египетской;
2CHR|7|9|а в день восьмой сделали попразднство, ибо освящение жертвенника совершали семь дней и праздник семь дней.
2CHR|7|10|И в двадцать третий день седьмого месяца [царь] отпустил народ в шатры их, радующийся и веселящийся в сердце о благе, какое сделал Господь Давиду и Соломону и Израилю, народу Своему.
2CHR|7|11|И окончил Соломон дом Господень и дом царский; и все, что предположил Соломон в сердце своем сделать в доме Господнем и в доме своем, совершил он успешно.
2CHR|7|12|И явился Господь Соломону ночью и сказал ему: Я услышал молитву твою и избрал Себе место сие в дом жертвоприношения.
2CHR|7|13|Если Я заключу небо и не будет дождя, и если повелю саранче поядать землю, или пошлю моровую язву на народ Мой,
2CHR|7|14|и смирится народ Мой, который именуется именем Моим, и будут молиться, и взыщут лица Моего, и обратятся от худых путей своих, то Я услышу с неба и прощу грехи их и исцелю землю их.
2CHR|7|15|Ныне очи Мои будут отверсты и уши Мои внимательны к молитве на месте сем.
2CHR|7|16|И ныне Я избрал и освятил дом сей, чтобы имя Мое было там во веки; и очи Мои и сердце Мое будут там во все дни.
2CHR|7|17|И если ты будешь ходить пред лицем Моим, как ходил Давид, отец твой, и будешь делать все, что Я повелел тебе, и будешь хранить уставы Мои и законы Мои,
2CHR|7|18|то утвержу престол царства твоего, как Я обещал Давиду, отцу твоему, говоря: не прекратится у тебя [муж], владеющий Израилем.
2CHR|7|19|Если же вы отступите и оставите уставы Мои и заповеди Мои, которые Я дал вам, и пойдете и станете служить богам иным и поклоняться им,
2CHR|7|20|то Я истреблю [Израиля] с лица земли Моей, которую Я дал им, и храм сей, который Я освятил имени Моему, отвергну от лица Моего и сделаю его притчею и посмешищем у всех народов.
2CHR|7|21|И о храме сем высоком всякий, проходящий мимо него, ужаснется и скажет: за что поступил так Господь с землею сею и с храмом сим?
2CHR|7|22|И скажут: за то, что они оставили Господа, Бога отцов своих, Который вывел их из земли Египетской, и прилепились к богам иным, и поклонялись им, и служили им, – за то Он навел на них все это бедствие.
2CHR|8|1|По окончании двадцати лет, в которые Соломон строил дом Господень и свой дом,
2CHR|8|2|Соломон обстроил и города, которые дал Соломону Хирам, и поселил в них сынов Израилевых.
2CHR|8|3|И пошел Соломон на Емаф–Сува и взял его.
2CHR|8|4|И построил он Фадмор в пустыне, и все города для запасов, какие основал в Емафе.
2CHR|8|5|Он обстроил Вефорон верхний и Вефорон нижний, города укрепленные, со стенами, воротами и запорами,
2CHR|8|6|и Ваалаф и все города для запасов, которые были у Соломона, и все города для колесниц, и города для конных, и все, что хотел Соломон построить в Иерусалиме и на Ливане и во всей земле владения своего.
2CHR|8|7|Весь народ, оставшийся от Хеттеев, и Аморреев, и Ферезеев, и Евеев и Иевусеев, которые были не из сынов Израилевых, –
2CHR|8|8|детей их, оставшихся после них на земле, которых не истребили сыны Израилевы, – сделал Соломон оброчными до сего дня.
2CHR|8|9|Сынов же Израилевых не делал Соломон работниками по делам своим, но они были воинами, и начальниками телохранителей его, и вождями колесниц его и всадников его.
2CHR|8|10|И было главных приставников у царя Соломона, управлявших народом, двести пятьдесят.
2CHR|8|11|А дочь Фараонову перевел Соломон из города Давидова в дом, который построил для нее, потому что, говорил он, не должна жить женщина у меня в доме Давида, царя Израилева, ибо свят он, так как вошел в него ковчег Господень.
2CHR|8|12|Тогда стал возносить Соломон всесожжения Господу на жертвеннике Господнем, который он устроил пред притвором,
2CHR|8|13|чтобы по уставу каждого дня приносить всесожжения, по заповеди Моисеевой, в субботы, и в новомесячия, и в праздники три раза в год: в праздник опресноков, и в праздник седмиц, и в праздник кущей.
2CHR|8|14|И установил он, по распоряжению Давида, отца своего, череды священников по службе их и левитов по стражам их, чтобы они славословили и служили при священниках по уставу каждого дня, и привратников по чередам их, к каждым воротам, потому что таково было завещание Давида, человека Божия.
2CHR|8|15|И не отступали от повелений царя о священниках и левитах ни в чем, ни в отношении сокровищ.
2CHR|8|16|Так устроено было все дело Соломоново от дня основания дома Господня до совершенного окончания его – дома Господня.
2CHR|8|17|Тогда пошел Соломон в Ецион–Гавер и в Елаф, который на берегу моря, в земле Идумейской.
2CHR|8|18|И прислал ему Хирам чрез слуг своих корабли и рабов, знающих море, и отправились они с слугами Соломоновыми в Офир, и добыли оттуда четыреста пятьдесят талантов золота, и привезли царю Соломону.
2CHR|9|1|Царица Савская, услышав о славе Соломона, пришла испытать Соломона загадками в Иерусалим, с весьма большим богатством, и с верблюдами, навьюченными благовониями и множеством золота и драгоценных камней. И пришла к Соломону и беседовала с ним обо всем, что было на сердце у нее.
2CHR|9|2|И объяснил ей Соломон все слова ее, и не нашлось ничего незнакомого Соломону, чего он не объяснил бы ей.
2CHR|9|3|И увидела царица Савская мудрость Соломона и дом, который он построил,
2CHR|9|4|и пищу за столом его, и жилище рабов его, и чинность служащих ему и одежду их, и виночерпиев его и одежду их, и ход, которым он ходил в дом Господень, – и была она вне себя.
2CHR|9|5|И сказала царю: верно то, что я слышала в земле моей о делах твоих и о мудрости твоей,
2CHR|9|6|но я не верила словам о них, доколе не пришла и не увидела глазами своими. И вот, мне и вполовину не сказано о множестве мудрости твоей: ты превосходишь молву, какую я слышала.
2CHR|9|7|Блаженны люди твои, и блаженны сии слуги твои, всегда предстоящие пред тобою и слышащие мудрость твою!
2CHR|9|8|Да будет благословен Господь Бог твой, Который благоволил посадить тебя на престол Свой в царя у Господа Бога твоего. По любви Бога твоего к Израилю, чтоб утвердить его на веки, Он поставил тебя царем над ним – творить суд и правду.
2CHR|9|9|И подарила она царю сто двадцать талантов золота и великое множество благовоний и драгоценных камней; и не бывало таких благовоний, какие подарила царица Савская царю Соломону.
2CHR|9|10|И слуги Хирамовы и слуги Соломоновы, которые привезли золото из Офира, привезли и красного дерева и драгоценных камней.
2CHR|9|11|И сделал царь из этого красного дерева лестницы к дому Господню и к дому царскому, и цитры и псалтири для певцов. И не видано было подобного сему прежде в земле Иудейской.
2CHR|9|12|Царь же Соломон дал царице Савской все, чего она желала и чего она просила, кроме таких вещей, какие она привезла царю. И она отправилась обратно в землю свою, она и слуги ее.
2CHR|9|13|Весу в золоте, которое приходило к Соломону в один год, [было] шестьсот шестьдесят шесть талантов золота.
2CHR|9|14|Сверх того, послы и купцы приносили, и все цари Аравийские и начальники областные приносили золото и серебро Соломону.
2CHR|9|15|И сделал царь Соломон двести больших щитов из кованого золота, – по шестисот [сиклей] кованого золота пошло на каждый щит, –
2CHR|9|16|и триста щитов меньших из кованого золота, – по триста [сиклей] золота пошло на каждый щит; и поставил их царь в доме из Ливанского дерева.
2CHR|9|17|И сделал царь большой престол из слоновой кости и обложил его чистым золотом,
2CHR|9|18|и шесть ступеней к престолу и золотое подножие, к престолу приделанное, и локотники по обе стороны у места сидения, и двух львов, стоящих возле локотников,
2CHR|9|19|и [еще] двенадцать львов, стоящих там на шести ступенях, по обе стороны. Не бывало такого [престола] ни в одном царстве.
2CHR|9|20|И все сосуды для питья у царя Соломона [были] из золота, и все сосуды в доме из Ливанского дерева [были] из золота отборного; серебро во дни Соломона вменялось ни во что,
2CHR|9|21|ибо корабли царя ходили в Фарсис с слугами Хирама, и в три года раз возвращались корабли из Фарсиса и привозили золото и серебро, слоновую кость и обезьян и павлинов.
2CHR|9|22|И превзошел царь Соломон всех царей земли богатством и мудростью.
2CHR|9|23|И все цари земли искали видеть Соломона, чтобы послушать мудрости его, которую вложил Бог в сердце его.
2CHR|9|24|И каждый из них подносил от себя в дар сосуды серебряные и сосуды золотые и одежды, оружие и благовония, коней и лошаков, из года в год.
2CHR|9|25|И было у Соломона четыре тысячи стойл для коней и колесниц и двенадцать тысяч всадников; и он разместил их в городах колесничных и при царе – в Иерусалиме;
2CHR|9|26|и господствовал он над всеми царями, от реки [Евфрата] до земли Филистимской и до пределов Египта.
2CHR|9|27|И сделал царь серебро в Иерусалиме равноценным [простому] камню, а кедры, по их множеству, сделал равноценными сикоморам, которые на низких местах.
2CHR|9|28|Коней приводили Соломону из Египта и из всех земель.
2CHR|9|29|Прочие деяния Соломоновы, первые и последние, описаны в записях Нафана пророка и в пророчестве Ахии Силомлянина и в видениях прозорливца Иоиля о Иеровоаме, сыне Наватовом.
2CHR|9|30|Царствовал же Соломон в Иерусалиме над всем Израилем сорок лет.
2CHR|9|31|И почил Соломон с отцами своими, и похоронили его в городе Давида, отца его. И воцарился Ровоам, сын его, вместо него.
2CHR|10|1|И пошел Ровоам в Сихем, потому что в Сихем сошлись все Израильтяне, чтобы поставить его царем.
2CHR|10|2|Когда услышал [о сем] Иеровоам, сын Наватов, – он находился в Египте, куда убежал от царя Соломона, – то возвратился Иеровоам из Египта.
2CHR|10|3|И послали и звали его; и пришел Иеровоам и весь Израиль, и говорили Ровоаму так:
2CHR|10|4|отец твой наложил на нас тяжкое иго; но ты облегчи жестокую работу отца твоего и тяжкое иго, которое он наложил на нас, и мы будем служить тебе.
2CHR|10|5|И сказал им [Ровоам]: через три дня придите опять ко мне. И разошелся народ.
2CHR|10|6|И советовался царь Ровоам со старейшинами, которые предстояли пред лицем Соломона, отца его, при жизни его, и говорил: как вы посоветуете отвечать народу сему?
2CHR|10|7|Они сказали ему: если ты будешь добр к народу сему и угодишь им и будешь говорить с ними ласково, то они будут тебе рабами на все дни.
2CHR|10|8|Но он оставил совет старейшин, который они давали ему, и стал советоваться с людьми молодыми, которые выросли вместе с ним, предстоящими пред лицем его;
2CHR|10|9|и сказал им: что вы посоветуете мне отвечать народу сему, говорившему мне так: облегчи иго, которое наложил на нас отец твой?
2CHR|10|10|И говорили ему молодые люди, выросшие вместе с ним, и сказали: так скажи народу, говорившему тебе: отец твой наложил на нас тяжкое иго, а ты облегчи нас, – так скажи им: мизинец мой толще чресл отца моего.
2CHR|10|11|Отец мой наложил на вас тяжкое иго, а я увеличу иго ваше; отец мой наказывал вас бичами, а я [буду бить вас] скорпионами.
2CHR|10|12|И пришел Иеровоам и весь народ к Ровоаму на третий день, как приказал царь, сказав: придите ко мне опять чрез три дня.
2CHR|10|13|Тогда царь отвечал им сурово, ибо оставил царь Ровоам совет старейшин, и говорил им по совету молодых людей так:
2CHR|10|14|отец мой наложил на вас тяжкое иго, а я увеличу его; отец мой наказывал вас бичами, а я [буду бить вас] скорпионами.
2CHR|10|15|И не послушал царь народа, потому что так устроено было от Бога, чтоб исполнить Господу слово Свое, которое изрек Он чрез Ахию Силомлянина Иеровоаму, сыну Наватову.
2CHR|10|16|Когда весь Израиль увидел, что не слушает его царь, то отвечал народ царю, говоря: какая нам часть в Давиде? Нет нам доли в сыне Иессеевом; по шатрам своим, Израиль! Теперь знай свой дом, Давид. И разошлись все Израильтяне по шатрам своим.
2CHR|10|17|Только над сынами Израилевыми, жившими в городах Иудиных, остался царем Ровоам.
2CHR|10|18|И послал царь Ровоам Адонирама, начальника над собиранием даней, и забросали его сыны Израилевы каменьями, и он умер. Царь же Ровоам поспешил сесть на колесницу, чтобы убежать в Иерусалим.
2CHR|10|19|Так отложились Израильтяне от дома Давидова до сего дня.
2CHR|11|1|И прибыл Ровоам в Иерусалим и созвал из дома Иудина и Вениаминова сто восемьдесят тысяч отборных воинов, чтобы воевать с Израилем и возвратить царство Ровоаму.
2CHR|11|2|И было слово Господне к Самею, человеку Божию, и сказано:
2CHR|11|3|скажи Ровоаму, сыну Соломонову, царю Иудейскому, и всему Израилю в [колене] Иудином и Вениаминовом:
2CHR|11|4|так говорит Господь: не ходите и не начинайте войны с братьями вашими; возвратитесь каждый в дом свой, ибо Мною сделано это. Они послушались слов Господних и возвратились из похода против Иеровоама.
2CHR|11|5|Ровоам жил в Иерусалиме; он обнес города в Иудее стенами.
2CHR|11|6|Он укрепил Вифлеем и Ефам, и Фекою,
2CHR|11|7|и Вефцур, и Сохо, и Одоллам,
2CHR|11|8|и Геф, и Марешу, и Зиф,
2CHR|11|9|и Адораим, и Лахис, и Азеку,
2CHR|11|10|и Цору, и Аиалон, и Хеврон, находившиеся в колене Иудином и Вениаминовом.
2CHR|11|11|И утвердил он крепости сии, и устроил в них начальников и хранилища для хлеба и деревянного масла и вина.
2CHR|11|12|И [дал] в каждый город щиты и копья и утвердил их весьма сильно. И оставались за ним Иуда и Вениамин.
2CHR|11|13|И священники и левиты, какие [были] по всей земле Израильской, собрались к нему из всех пределов,
2CHR|11|14|ибо оставили левиты свои городские предместья и свои владения и пришли в Иудею и в Иерусалим, так как оставил их Иеровоам и сыновья его от священства Господня
2CHR|11|15|и поставил у себя жрецов к высотам, и к козлам, и к тельцам, которых он сделал.
2CHR|11|16|А за ними и из всех колен Израилевых расположившие сердце свое, чтобы взыскать Господа Бога Израилева, приходили в Иерусалим, дабы приносить жертвы Господу Богу отцов своих.
2CHR|11|17|И укрепили они царство Иудино и поддерживали Ровоама, сына Соломонова, три года, потому что ходили путем Давида и Соломона в сии три года.
2CHR|11|18|И взял себе Ровоам в жену Махалафу, дочь Иеромофа, сына Давидова, и Авихаиль, дочь Елиава, сына Иессеева,
2CHR|11|19|и она родила ему сыновей: Иеуса и Шемарию и Загама.
2CHR|11|20|После нее он взял Мааху, дочь Авессалома, и она родила ему Авию и Аттая, и Зизу и Шеломифа.
2CHR|11|21|И любил Ровоам Мааху, дочь Авессалома, более всех жен и наложниц своих, ибо он имел восемнадцать жен и шестьдесят наложниц и родил двадцать восемь сыновей и шестьдесят дочерей.
2CHR|11|22|И поставил Ровоам Авию, сына Маахи, главою [и] князем над братьями его, потому что [хотел] воцарить его.
2CHR|11|23|И действовал благоразумно, и разослал всех сыновей своих по всем землям Иуды и Вениамина во все укрепленные города, и дал им содержание большое и приискал много жен.
2CHR|12|1|Когда царство Ровоама утвердилось, и он сделался силен, тогда он оставил закон Господень, и весь Израиль с ним.
2CHR|12|2|На пятом году царствования Ровоама, Сусаким, царь Египетский, пошел на Иерусалим, – потому что они отступили от Господа, –
2CHR|12|3|с тысячью и двумя стами колесниц и шестьюдесятью тысячами всадников; и не было числа народу, который пришел с ним из Египта, Ливиянам, Сукхитам и Ефиоплянам;
2CHR|12|4|и взял укрепленные города в Иудее и пришел к Иерусалиму.
2CHR|12|5|Тогда Самей пророк пришел к Ровоаму и князьям Иудеи, которые собрались в Иерусалим, [спасаясь] от Сусакима, и сказал им: так говорит Господь: вы оставили Меня, за то и Я оставляю вас в руки Сусакиму.
2CHR|12|6|И смирились князья Израилевы и царь и сказали: праведен Господь!
2CHR|12|7|Когда увидел Господь, что они смирились, тогда было слово Господне к Самею, и сказано: они смирились; не истреблю их и вскоре дам им избавление, и не прольется гнев Мой на Иерусалим рукою Сусакима;
2CHR|12|8|однакоже они будут слугами его, чтобы знали, каково служить Мне и служить царствам земным.
2CHR|12|9|И пришел Сусаким, царь Египетский, в Иерусалим и взял сокровища дома Господня и сокровища дома царского; все взял он, взял и щиты золотые, которые сделал Соломон.
2CHR|12|10|И сделал царь Ровоам, вместо их, щиты медные, и отдал их на руки начальникам телохранителей, охранявших вход дома царского.
2CHR|12|11|Когда выходил царь в дом Господень, приходили телохранители и несли их, и потом опять относили их в палату телохранителей.
2CHR|12|12|И когда он смирился, тогда отвратился от него гнев Господа и не погубил его до конца; притом и в Иудее было нечто доброе.
2CHR|12|13|И утвердился царь Ровоам в Иерусалиме и царствовал. Сорок один год было Ровоаму, когда он воцарился, и семнадцать лет царствовал в Иерусалиме, в городе, который из всех колен Израилевых избрал Господь, чтобы там пребывало имя Его. Имя матери его Наама, Аммонитянка.
2CHR|12|14|И делал он зло, потому что не расположил сердца своего к тому, чтобы взыскать Господа.
2CHR|12|15|Деяния Ровоамовы, первые и последние, описаны в записях Самея пророка и Адды прозорливца при родословиях. И были войны у Ровоама с Иеровоамом во все дни.
2CHR|12|16|И почил Ровоам с отцами своими и погребен в городе Давидовом. И воцарился Авия, сын его, вместо него.
2CHR|13|1|В восемнадцатый год царствования Иеровоама воцарился Авия над Иудою.
2CHR|13|2|Три года он царствовал в Иерусалиме; имя матери его Михаия, дочь Уриилова, из Гивы. И была война у Авии с Иеровоамом.
2CHR|13|3|И вывел Авия на войну войско, состоявшее из людей храбрых, из четырехсот тысяч человек отборных; а Иеровоам выступил против него на войну с восемью стами тысяч человек, [также] отборных, храбрых.
2CHR|13|4|И стал Авия на вершине горы Цемараимской, одной из гор Ефремовых, и говорил: послушайте меня, Иеровоам и все Израильтяне!
2CHR|13|5|Не знаете ли вы, что Господь Бог Израилев дал царство Давиду над Израилем навек, ему и сыновьям его, по завету соли?
2CHR|13|6|Но восстал Иеровоам, сын Наватов, раб Соломона, сына Давидова, и возмутился против господина своего.
2CHR|13|7|И собрались вокруг него люди пустые, люди развращенные, и укрепились против Ровоама, сына Соломонова; Ровоам же был молод и слаб сердцем и не устоял против них.
2CHR|13|8|И ныне вы думаете устоять против царства Господня в руке сынов Давидовых, [потому что] вас великое множество, и у вас золотые тельцы, которых Иеровоам сделал вам богами.
2CHR|13|9|Не вы ли изгнали священников Господних, сынов Аарона, и левитов, и поставили у себя священников, какие у народов [других] земель? Всякий, кто приходит для посвящения своего с тельцом и с семью овнами, делается [у вас] священником лжебогов.
2CHR|13|10|А у нас – Господь Бог наш; мы не оставляли Его, и Господу служат священники, сыны Аароновы, и левиты при [своем] деле.
2CHR|13|11|И сожигают они Господу всесожжения каждое утро и каждый вечер, и благовонное курение, и полагают рядами хлебы на столе чистом, и [зажигают] золотой светильник и лампады его, чтобы горели каждый вечер, потому что мы соблюдаем установление Господа Бога нашего, а вы оставили Его.
2CHR|13|12|И вот, у нас во главе Бог, и священники Его, и трубы громогласные, чтобы греметь против вас. Сыны Израилевы! не воюйте с Господом Богом отцов ваших, ибо не получите успеха.
2CHR|13|13|Между тем Иеровоам послал отряд в засаду с тыла им, так что [сам] [он] был впереди Иудеев, а засада позади их.
2CHR|13|14|И оглянулись Иудеи, и вот, им битва спереди и сзади; и возопили они к Господу, а священники затрубили трубами.
2CHR|13|15|И воскликнули Иудеи. И когда воскликнули Иудеи, Бог поразил Иеровоама и всех Израильтян пред лицем Авии и Иуды.
2CHR|13|16|И побежали сыны Израилевы от Иудеев, и предал их Бог в руки им.
2CHR|13|17|И произвели у них Авия и народ его поражение сильное; и пало убитых у Израиля пятьсот тысяч человек отборных.
2CHR|13|18|И смирились тогда сыны Израилевы, и были сильны сыны Иудины, потому что уповали на Господа Бога отцов своих.
2CHR|13|19|И преследовал Авия Иеровоама и взял у него города: Вефиль и зависящие от него города, и Иешану и зависящие от нее города, и Ефрон и зависящие от него города.
2CHR|13|20|И не входил уже в силу Иеровоам во дни Авии. И поразил его Господь, и он умер.
2CHR|13|21|Авия же усилился; и взял себе четырнадцать жен и родил двадцать два сына и шестнадцать дочерей.
2CHR|13|22|Прочие деяния Авии и его поступки и слова описаны в сказании пророка Адды.
2CHR|13|23|И почил Авия с отцами своими, и похоронили его в городе Давидовом. И воцарился Аса, сын его, вместо него. Во дни его покоилась земля десять лет.
2CHR|14|1|И делал Аса доброе и угодное в очах Господа Бога своего:
2CHR|14|2|и отверг он жертвенники [богов] чужих и высоты, и разбил статуи, и вырубил [посвященные] дерева;
2CHR|14|3|и повелел Иудеям взыскать Господа Бога отцов своих, и исполнять закон [Его] и заповеди;
2CHR|14|4|и отменил он во всех городах Иудиных высоты и статуи солнца. И спокойно было при нем царство.
2CHR|14|5|И построил он укрепленные города в Иудее, ибо спокойна была земля, и не было у него войны в те годы, так как Господь дал покой ему.
2CHR|14|6|И сказал он Иудеям: построим города сии и обнесем их стенами с башнями, с воротами и запорами. Земля еще наша, потому что мы взыскали Господа Бога нашего: мы взыскали Его, – и Он дал нам покой со всех сторон. И стали строить, и имели успех.
2CHR|14|7|И было у Асы военной силы: вооруженных щитом и копьем из [колена] Иудина триста тысяч, и из [колена] Вениаминова вооруженных щитом и стрелявших из лука двести восемьдесят тысяч, людей храбрых.
2CHR|14|8|И вышел на них Зарай Ефиоплянин с войском в тысячу тысяч и с тремя стами колесниц и дошел до Мареши.
2CHR|14|9|И выступил Аса против него, и построились к сражению на долине Цефата у Мареши.
2CHR|14|10|И воззвал Аса к Господу Богу своему, и сказал: Господи! не в Твоей ли силе помочь сильному или бессильному? помоги же нам, Господи Боже наш: ибо мы на Тебя уповаем и во имя Твое вышли мы против множества сего. Господи! Ты Бог наш: да не превозможет Тебя человек.
2CHR|14|11|И поразил Господь Ефиоплян пред лицем Асы и пред лицем Иуды, и побежали Ефиопляне.
2CHR|14|12|И преследовал их Аса и народ, бывший с ним, до Герара, и пали Ефиопляне, так что у них никого [не осталось] в живых, потому что они поражены были пред Господом и пред воинством Его. И набрали добычи великое множество.
2CHR|14|13|И разрушили все города вокруг Герара, потому что напал на них ужас от Господа; и разграбили все города и вынесли из них весьма много добычи.
2CHR|14|14|Также и пастушеские шалаши разорили и угнали множество стад мелкого скота и верблюдов и возвратились в Иерусалим.
2CHR|15|1|Тогда на Азарию, сына Одедова, сошел Дух Божий,
2CHR|15|2|и вышел он навстречу Асе и сказал ему: послушайте меня, Аса и весь Иуда и Вениамин: Господь с вами, когда вы с Ним; и если будете искать Его, Он будет найден вами; если же оставите Его, Он оставит вас.
2CHR|15|3|Многие дни Израиль [будет] без Бога истинного, и без священника учащего, и без закона;
2CHR|15|4|но когда он обратится в тесноте своей к Господу Богу Израилеву и взыщет Его, Он даст им найти Себя.
2CHR|15|5|В те времена не будет мира ни выходящему, ни входящему, ибо великие волнения будут у всех жителей земель;
2CHR|15|6|народ будет сражаться с народом, и город с городом, потому что Бог приведет их в смятение всякими бедствиями.
2CHR|15|7|Но вы укрепитесь, и пусть не ослабевают руки ваши, потому что есть возмездие за дела ваши.
2CHR|15|8|Когда услышал Аса слова сии и пророчество, [сына] Одеда пророка, то ободрился и изверг мерзости [языческие] из всей земли Иудиной и Вениаминовой и из городов, которые он взял на горе Ефремовой, и обновил жертвенник Господень, который пред притвором Господним.
2CHR|15|9|И собрал всего Иуду и Вениамина и живущих с ними переселенцев от Ефрема и Манассии и Симеона; ибо многие от Израиля перешли к нему, когда увидели, что Господь, Бог его, с ним.
2CHR|15|10|И собрались в Иерусалим в третий месяц, в пятнадцатый год царствования Асы;
2CHR|15|11|и принесли в день тот жертву Господу из добычи, которую привели, из крупного скота семьсот и из мелкого семь тысяч;
2CHR|15|12|и вступили в завет, чтобы взыскать Господа Бога отцов своих от всего сердца своего и от всей души своей;
2CHR|15|13|а всякий, кто не станет искать Господа Бога Израилева, должен умереть, малый ли он или большой, мужчина ли или женщина.
2CHR|15|14|И клялись Господу громогласно и с восклицанием и при [звуке] труб и рогов.
2CHR|15|15|И радовались все Иудеи сей клятве, потому что от всего сердца своего клялись и со всем усердием взыскали Его, и Он дал им найти Себя. И дал им Господь покой со всех сторон.
2CHR|15|16|И Мааху, мать свою, царь Аса лишил царского достоинства за то, что она сделала истукан для дубравы. И ниспроверг Аса истукан ее, и изрубил в куски, и сжег на долине Кедрона.
2CHR|15|17|Хотя высоты не были отменены у Израиля, но сердце Асы было вполне предано [Господу] во все дни его.
2CHR|15|18|И внес он посвященное отцом его и свое посвящение в дом Божий, серебро и золото и сосуды.
2CHR|15|19|И не было войны до тридцать пятого года царствования Асы.
2CHR|16|1|В тридцать шестой год царствования Асы, пошел Вааса, царь Израильский, на Иудею и начал строить Раму, чтобы не позволить [никому] ни уходить от Асы, царя Иудейского, ни приходить [к нему].
2CHR|16|2|И вынес Аса серебро и золото из сокровищниц дома Господня и дома царского и послал к Венададу, царю Сирийскому, жившему в Дамаске, говоря:
2CHR|16|3|союз да будет между мною и тобою, как был между отцом моим и отцом твоим; вот, я посылаю тебе серебра и золота: пойди, расторгни союз твой с Ваасою, царем Израильским, чтоб он отступил от меня.
2CHR|16|4|И послушался Венадад царя Асы и послал военачальников, которые [были] у него, против городов Израильских, и они опустошили Ийон и Дан и Авелмаим и все запасы в городах Неффалимовых.
2CHR|16|5|И когда услышал [о сем] Вааса, то перестал строить Раму и прекратил работу свою.
2CHR|16|6|Аса же царь собрал всех Иудеев, и они вывезли [из] Рамы камни и дерева, которые употреблял Вааса для строения, – и выстроил из них Геву и Мицфу.
2CHR|16|7|В то время пришел Ананий прозорливец к Асе, царю Иудейскому, и сказал ему: так как ты понадеялся на царя Сирийского и не уповал на Господа Бога твоего, потому и спаслось войско царя Сирийского от руки твоей.
2CHR|16|8|Не были ли Ефиопляне и Ливияне с силою большею и с колесницами и всадниками весьма многочисленными? Но как ты уповал на Господа, то Он предал их в руку твою,
2CHR|16|9|ибо очи Господа обозревают всю землю, чтобы поддерживать тех, [чье] сердце вполне предано Ему. Безрассудно ты поступил теперь. За то отныне будут у тебя войны.
2CHR|16|10|И разгневался Аса на прозорливца, и заключил его в темницу, так как за это был в раздражении на него; притеснял Аса и [некоторых] из народа в то время.
2CHR|16|11|И вот, деяния Асы, первые и последние, описаны в книге царей Иудейских и Израильских.
2CHR|16|12|И сделался Аса болен ногами на тридцать девятом году царствования своего, и болезнь его поднялась до верхних частей тела; но он в болезни своей взыскал не Господа, а врачей.
2CHR|16|13|И почил Аса с отцами своими, и умер на сорок первом году царствования своего.
2CHR|16|14|И похоронили его в гробнице, которую он устроил для себя в городе Давидовом; и положили его на одре, который наполнили благовониями и разными искусственными мастями, и сожгли их для него великое множество.
2CHR|17|1|И воцарился Иосафат, сын его, вместо него; и укрепился он против Израильтян.
2CHR|17|2|И поставил он войско во все укрепленные города Иудеи и расставил охранное войско по земле Иудейской и по городам Ефремовым, которыми овладел Аса, отец его.
2CHR|17|3|И был Господь с Иосафатом, потому что он ходил первыми путями Давида, отца своего, и не взыскал Ваалов,
2CHR|17|4|но взыскал он Бога отца своего и поступал по заповедям Его, а не по деяниям Израильтян.
2CHR|17|5|И утвердил Господь царство в руке его, и давали все Иудеи дары Иосафату, и было у него много богатства и славы.
2CHR|17|6|И возвысилось сердце его на путях Господних; притом и высоты отменил он и дубравы в Иудее.
2CHR|17|7|И в третий год царствования своего он послал князей своих Бенхаила и Овадию, и Захарию и Нафанаила и Михея, чтоб учили по городам Иудиным народ,
2CHR|17|8|и с ними левитов: Шемаию и Нефанию, и Зевадию и Азаила, и Шемирамофа и Ионафана, и Адонию и Товию и Тов–Адонию, и с ними Елишаму и Иорама, священников.
2CHR|17|9|И они учили в Иудее, имея с собою книгу закона Господня; и обходили все города Иудеи и учили народ.
2CHR|17|10|И был страх Господень на всех царствах земель, которые вокруг Иудеи, и не воевали с Иосафатом.
2CHR|17|11|А от Филистимлян приносили Иосафату дары и в дань серебро; также Аравитяне пригоняли к нему мелкий скот: овнов семь тысяч семьсот и козлов семь тысяч семьсот.
2CHR|17|12|И возвышался Иосафат все более и более и построил в Иудее крепости и города для запасов.
2CHR|17|13|Много было у него запасов в городах Иудейских, а в Иерусалиме людей военных, храбрых.
2CHR|17|14|И вот список их по поколениям их: у Иуды начальники тысяч: Адна начальник, и у него отличных воинов триста тысяч;
2CHR|17|15|за ним Иоханан начальник, и у него двести восемьдесят тысяч;
2CHR|17|16|за ним Амасия, сын Зихри, посвятивший себя Господу, и у него двести тысяч воинов отличных.
2CHR|17|17|У Вениамина: отличный воин Елиада, и у него вооруженных луком и щитом двести тысяч;
2CHR|17|18|за ним Иегозавад, и у него сто восемьдесят тысяч вооруженных воинов.
2CHR|17|19|Вот служившие царю, сверх тех, которых расставил царь в укрепленных городах по всей Иудее.
2CHR|18|1|И было у Иосафата много богатства и славы; и породнился он с Ахавом.
2CHR|18|2|И пошел чрез несколько лет к Ахаву в Самарию; и заколол для него Ахав множество скота мелкого и крупного, и для людей, бывших с ним, и склонял его идти на Рамоф Галаадский.
2CHR|18|3|И говорил Ахав, царь Израильский, Иосафату, царю Иудейскому: пойдешь ли со мною в Рамоф Галаадский? Тот сказал ему: как ты, так и я, как твой народ, так и мой народ: [иду] с тобою на войну!
2CHR|18|4|И сказал Иосафат царю Израильскому: вопроси сегодня, что скажет Господь.
2CHR|18|5|И собрал царь Израильский пророков четыреста человек и сказал им: идти ли нам на Рамоф Галаадский войною, или удержаться? Они сказали: иди, и Бог предаст [его] в руку царя.
2CHR|18|6|И сказал Иосафат: нет ли здесь еще пророка Господня? спросим и у него.
2CHR|18|7|И сказал царь Израильский Иосафату: есть еще один человек, чрез которого можно вопросить Господа; но я не люблю его, потому что он не пророчествует обо мне доброго, а постоянно пророчествует худое; это Михей, сын Иемвлая. И сказал Иосафат: не говори так, царь.
2CHR|18|8|И позвал царь Израильский одного евнуха, и сказал: сходи поскорее за Михеем, сыном Иемвлая.
2CHR|18|9|Царь же Израильский и Иосафат, царь Иудейский, сидели каждый на своем престоле, одетые в [царские] одежды; сидели на площади у ворот Самарии, и все пророки пророчествовали пред ними.
2CHR|18|10|И сделал себе Седекия, сын Хенааны, железные рога и сказал: так говорит Господь: сими избодешь Сириян до истребления их.
2CHR|18|11|И все пророки пророчествовали то же, говоря: иди на Рамоф Галаадский; будет успех тебе, и предаст [его] Господь в руку царя.
2CHR|18|12|Посланный, который пошел позвать Михея, говорил ему: вот, пророки единогласно предрекают доброе царю; пусть бы и твое слово было такое же, как каждого из них: изреки и ты доброе.
2CHR|18|13|И сказал Михей: жив Господь, – что скажет мне Бог мой, то изреку я.
2CHR|18|14|И пришел он к царю, и сказал ему царь: Михей, идти ли нам войной на Рамоф Галаадский, или удержаться? И сказал тот: идите, будет вам успех, и они преданы будут в руки ваши.
2CHR|18|15|И сказал ему царь: сколько раз мне заклинать тебя, чтобы ты не говорил мне ничего, кроме истины, во имя Господне?
2CHR|18|16|Тогда [Михей] сказал: я видел всех сынов Израиля, рассеянных по горам, как овец, у которых нет пастыря, – и сказал Господь: нет у них начальника, пусть возвратятся каждый в дом свой с миром.
2CHR|18|17|И сказал царь Израильский Иосафату: не говорил ли я тебе, что он не пророчествует о мне доброго, а только худое?
2CHR|18|18|И сказал [Михей]: так выслушайте слово Господне: я видел Господа, седящего на престоле Своем, и все воинство небесное стояло по правую и по левую руку Его.
2CHR|18|19|И сказал Господь: кто увлек бы Ахава, царя Израильского, чтобы он пошел и пал в Рамофе Галаадском? И один говорил так, другой говорил иначе.
2CHR|18|20|И выступил один дух, и стал пред лицем Господа, и сказал: я увлеку его. И сказал ему Господь: чем?
2CHR|18|21|Тот сказал: я выйду, и буду духом лжи в устах всех пророков его. И сказал Он: ты увлечешь его, и успеешь; пойди и сделай так.
2CHR|18|22|И теперь, вот попустил Господь духу лжи [войти] в уста сих пророков твоих, но Господь изрек о тебе недоброе.
2CHR|18|23|И подошел Седекия, сын Хенааны, и ударил Михея по щеке, и сказал: по какой это дороге отошел от меня Дух Господень, чтобы говорить в тебе?
2CHR|18|24|И сказал Михей: вот, ты увидишь [это] в тот день, когда будешь бегать из комнаты в комнату, чтобы укрыться.
2CHR|18|25|И сказал царь Израильский: возьмите Михея и отведите его к Амону градоначальнику и к Иоасу, сыну царя,
2CHR|18|26|и скажите: так говорит царь: посадите этого в темницу и кормите его хлебом и водою скудно, доколе я не возвращусь в мире.
2CHR|18|27|И сказал Михей: если ты возвратишься в мире, то не Господь говорил чрез меня. И сказал: слушайте [это], все люди!
2CHR|18|28|И пошел царь Израильский и Иосафат, царь Иудейский, к Рамофу Галаадскому.
2CHR|18|29|И сказал царь Израильский Иосафату: я переоденусь и вступлю в сражение, а ты надень свои [царские] одежды. И переоделся царь Израильский, и вступили в сражение.
2CHR|18|30|И царь Сирийский повелел начальникам колесниц, бывших у него, сказав: не сражайтесь ни с малым, ни с великим, а только с одним царем Израильским.
2CHR|18|31|И когда увидели Иосафата начальники колесниц, то подумали: это царь Израильский, – и окружили его, чтобы сразиться с ним. Но Иосафат закричал, и Господь помог ему, и отвел их Бог от него.
2CHR|18|32|И когда увидели начальники колесниц, что [это] не был царь Израильский, то поворотили от него.
2CHR|18|33|Между тем один человек случайно натянул лук свой, и ранил царя Израильского сквозь швы лат. И сказал он вознице: повороти назад, и вези меня от войска, ибо я ранен.
2CHR|18|34|Но сражение в тот день усилилось; и царь Израильский стоял на колеснице напротив Сириян до вечера и умер на закате солнца.
2CHR|19|1|И возвращался Иосафат, царь Иудейский, в мире в дом свой в Иерусалим.
2CHR|19|2|И выступил навстречу ему Ииуй, сын Анании, прозорливец, и сказал царю Иосафату: [следовало] ли тебе помогать нечестивцу и любить ненавидящих Господа? За это на тебя гнев от лица Господня.
2CHR|19|3|Впрочем и доброе найдено в тебе, потому что ты истребил кумиры в земле [Иудейской] и расположил сердце свое к тому, чтобы взыскать Бога.
2CHR|19|4|И жил Иосафат в Иерусалиме. И опять стал он обходить народ [свой] от Вирсавии до горы Ефремовой, и обращал их к Господу, Богу отцов их.
2CHR|19|5|И поставил судей на земле по всем укрепленным городам Иудеи в каждом городе,
2CHR|19|6|и сказал судьям: смотрите, что вы делаете, вы творите не суд человеческий, но суд Господа; и [Он] с вами в деле суда.
2CHR|19|7|Итак да будет страх Господень на вас: действуйте осмотрительно, ибо нет у Господа Бога нашего неправды, ни лицеприятия, ни мздоимства.
2CHR|19|8|И в Иерусалиме приставил Иосафат [некоторых] из левитов и священников и глав поколений у Израиля – к суду Господню и к тяжбам. И возвратились в Иерусалим.
2CHR|19|9|И дал им повеление, говоря: так действуйте в страхе Господнем, с верностью и с чистым сердцем:
2CHR|19|10|во всяком деле спорном, какое поступит к вам от братьев ваших, живущих в городах своих, о кровопролитии ли, или о законе, заповеди, уставах и обрядах, наставляйте их, чтобы они не провинились пред Господом, и не было бы гнева [Его] на вас и на братьев ваших; так действуйте, – и вы не погрешите.
2CHR|19|11|И вот Амария первосвященник, над вами во всяком деле Господнем, а Зевадия, сын Исмаилов, князь дома Иудина, во всяком деле царя, и надзиратели левиты пред вами. Будьте тверды и действуйте, и будет Господь с добрым.
2CHR|20|1|После сего Моавитяне и Аммонитяне, а с ними некоторые из страны Маонитской, пошли войною на Иосафата.
2CHR|20|2|И пришли, и донесли Иосафату, говоря: идет на тебя множество великое из–за моря, от Сирии, и вот они в Хацацон–Фамаре, то есть в Енгедди.
2CHR|20|3|И убоялся Иосафат, и обратил лице свое взыскать Господа, и объявил пост по всей Иудее.
2CHR|20|4|И собрались Иудеи просить [помощи] у Господа; из всех городов Иудиных пришли они умолять Господа.
2CHR|20|5|И стал Иосафат в собрании Иудеев и Иерусалимлян в доме Господнем, пред новым двором,
2CHR|20|6|и сказал: Господи Боже отцов наших! Не Ты ли Бог на небе? И Ты владычествуешь над всеми царствами народов, и в Твоей руке сила и крепость, и никто не устоит против Тебя!
2CHR|20|7|Не Ты ли, Боже наш, изгнал жителей земли сей пред лицем народа Твоего Израиля и отдал ее семени Авраама, друга Твоего, навек?
2CHR|20|8|И они поселились на ней и построили Тебе на ней святилище во имя Твое, говоря:
2CHR|20|9|если придет на нас бедствие: меч наказующий, или язва, или голод, то мы станем пред домом сим и пред лицем Твоим, ибо имя Твое в доме сем; и воззовем к Тебе в тесноте нашей, и Ты услышишь и спасешь.
2CHR|20|10|И ныне вот Аммонитяне и Моавитяне и [обитатели] горы Сеира, чрез земли которых Ты не позволил пройти Израильтянам, когда они шли из земли Египетской, а потому они миновали их и не истребили их, –
2CHR|20|11|вот они платят нам [тем], что пришли выгнать нас из наследственного владения Твоего, которое Ты отдал нам.
2CHR|20|12|Боже наш! Ты суди их. Ибо нет в нас силы против множества сего великого, пришедшего на нас, и мы не знаем, что делать, но к Тебе очи наши!
2CHR|20|13|И все Иудеи стояли пред лицем Господним, и малые дети их, жены их и сыновья их.
2CHR|20|14|Тогда на Иозиила, сына Захарии, сына Ванеи, сына Иеиела, сына Матфании, левита из сынов Асафовых, сошел Дух Господень среди собрания
2CHR|20|15|и сказал он: слушайте, все Иудеи и жители Иерусалима и царь Иосафат! Так говорит Господь к вам: не бойтесь и не ужасайтесь множества сего великого, ибо не ваша война, а Божия.
2CHR|20|16|Завтра выступите против них: вот они всходят на возвышенность Циц, и вы найдете их на конце долины, пред пустынею Иеруилом.
2CHR|20|17|Не вам сражаться на сей раз; вы станьте, стойте и смотрите на спасение Господне, [посылаемое] вам. Иуда и Иерусалим! не бойтесь и не ужасайтесь. Завтра выступите навстречу им, и Господь будет с вами.
2CHR|20|18|И преклонился Иосафат лицем до земли, и все Иудеи и жители Иерусалима пали пред Господом, чтобы поклониться Господу.
2CHR|20|19|И встали левиты из сынов Каафовых и из сынов Кореевых – хвалить Господа Бога Израилева, голосом весьма громким.
2CHR|20|20|И встали они рано утром, и выступили к пустыне Фекойской; и когда они выступили, стал Иосафат и сказал: послушайте меня, Иудеи и жители Иерусалима! Верьте Господу Богу вашему, и будьте тверды; верьте пророкам Его, и будет успех вам.
2CHR|20|21|И совещался он с народом, и поставил певцов Господу, чтобы они в благолепии святыни, выступая впереди вооруженных, славословили и говорили: славьте Господа, ибо вовек милость Его!
2CHR|20|22|И в то время, [как] они стали восклицать и славословить, Господь возбудил несогласие между Аммонитянами, Моавитянами и [обитателями] горы Сеира, пришедшими на Иудею, и были они поражены:
2CHR|20|23|ибо восстали Аммонитяне и Моавитяне на обитателей горы Сеира, побивая и истребляя [их], а когда покончили с жителями Сеира, тогда стали истреблять друг друга.
2CHR|20|24|И когда Иудеи пришли на возвышенность к пустыне и взглянули на то многолюдство, и вот – трупы, лежащие на земле, и нет уцелевшего.
2CHR|20|25|И пришел Иосафат и народ его забирать добычу, и нашли у них во множестве и имущество, и одежды, и драгоценные вещи, и набрали себе столько, что не [могли] нести. И три дня они забирали добычу; так велика [была] она!
2CHR|20|26|А в четвертый день собрались на долину благословения, так как там они благословили Господа. Посему и называют то место долиною благословения до сего дня.
2CHR|20|27|И пошли назад все Иудеи и Иерусалимляне и Иосафат во главе их, чтобы возвратиться в Иерусалим с веселием, потому что дал им Господь торжество над врагами их.
2CHR|20|28|И пришли в Иерусалим с псалтирями, и цитрами, и трубами, к дому Господню.
2CHR|20|29|И был страх Божий на всех царствах земных, когда они услышали, что [Сам] Господь воевал против врагов Израиля.
2CHR|20|30|И спокойно стало царство Иосафатово, и дал ему Бог его покой со всех сторон.
2CHR|20|31|Так царствовал Иосафат над Иудеею: тридцати пяти лет он [был], когда воцарился, и двадцать пять лет царствовал в Иерусалиме. Имя матери его Азува, дочь Салаила.
2CHR|20|32|И ходил он путем отца своего Асы и не уклонился от него, делая угодное в очах Господних.
2CHR|20|33|Только высоты не были отменены, и народ еще не обратил твердо сердца своего к Богу отцов своих.
2CHR|20|34|Прочие деяния Иосафата, первые и последние, описаны в записях Ииуя, сына Ананиева, которые внесены в книгу царей Израилевых.
2CHR|20|35|Но после того вступил Иосафат, царь Иудейский в общение с Охозиею, царем Израильским, который поступал беззаконно,
2CHR|20|36|и соединился с ним, чтобы построить корабли для отправления в Фарсис; и построили они корабли в Ецион–Гавере.
2CHR|20|37|И изрек [тогда] Елиезер, сын Додавы из Мареши, пророчество на Иосафата, говоря: так как ты вступил в общение с Охозиею, то разрушил Господь дело твое. – И разбились корабли, и не могли идти в Фарсис.
2CHR|21|1|И почил Иосафат с отцами своими, и похоронен с отцами своими в городе Давидовом. И воцарился Иорам, сын его, вместо него.
2CHR|21|2|И у него [были] братья, сыновья Иосафата: Азария и Иехиил, и Захария и Азария, и Михаил и Сафатия: все сии сыновья Иосафата, царя Израилева.
2CHR|21|3|И дал им отец их большие подарки серебром и золотом и драгоценностями, вместе с укрепленными городами в Иудее; царство же отдал Иораму, потому что он первенец.
2CHR|21|4|И вступил Иорам на царство отца своего и утвердился, и умертвил всех братьев своих мечом и также [некоторых] из князей Израилевых.
2CHR|21|5|Тридцати двух лет [был] Иорам, когда воцарился, и восемь лет царствовал в Иерусалиме;
2CHR|21|6|и ходил он путем царей Израильских, как поступал дом Ахавов, потому что дочь Ахава была женою его, – и делал он неугодное в очах Господних.
2CHR|21|7|Однакоже не хотел Господь погубить дома Давидова ради завета, который заключил с Давидом, и потому что обещал дать ему светильник и сыновьям его на все времена.
2CHR|21|8|Во дни его вышел Едом из–под власти Иуды, и поставили над собою царя.
2CHR|21|9|И пошел Иорам с военачальниками своими, и все колесницы с ним; и встав ночью, поразил Идумеян, которые окружили его, и начальствующих над колесницами.
2CHR|21|10|Однако вышел Едом из–под власти Иуды до сего дня. В то же время вышла и Ливна из–под власти его, потому что он оставил Господа Бога отцов своих.
2CHR|21|11|Также высоты устроил он на горах Иудейских, и ввел в блужение жителей Иерусалима и соблазнил Иудею.
2CHR|21|12|И пришло к нему письмо от Илии пророка, в котором было сказано: так говорит Господь Бог Давида, отца твоего: за то, что ты не пошел путями Иосафата, отца твоего, и путями Асы, царя Иудейского,
2CHR|21|13|а пошел путем царей Израильских и ввел в блужение Иудею и жителей Иерусалима, как вводил в блужение дом Ахавов, еще же и братьев твоих, дом отца твоего, которые лучше тебя, ты умертвил,
2CHR|21|14|[за то], вот Господь поразит поражением великим народ твой и сыновей твоих, и жен твоих, и все имущество твое,
2CHR|21|15|тебя же [самого] – болезнью сильною, болезнью внутренностей твоих до того, что будут выпадать внутренности твои от болезни со дня на день.
2CHR|21|16|И возбудил Господь против Иорама дух Филистимлян и Аравитян, сопредельных Ефиоплянам;
2CHR|21|17|и они пошли на Иудею и ворвались в нее, и захватили все имущество, находившееся в доме царя, также и сыновей его и жен его; и не осталось у него сына, кроме Охозии, меньшего из сыновей его.
2CHR|21|18|А после всего этого поразил Господь внутренности его болезнью неизлечимою.
2CHR|21|19|Так было со дня на день, а к концу второго года выпали внутренности его от болезни его, и он умер в жестоких страданиях; и не сожег для него народ его [благовоний], как делал то для отцов его.
2CHR|21|20|Тридцати двух [лет] был он, когда воцарился, и восемь лет царствовал в Иерусалиме, и отошел неоплаканный, и похоронили его в городе Давидовом, но не в царских гробницах.
2CHR|22|1|И поставили царем жители Иерусалима Охозию, меньшего сына его, вместо него, так как всех старших избило полчище, приходившее с Аравитянами к стану, – и воцарился Охозия, сын Иорама, царя Иудейского.
2CHR|22|2|Двадцати двух лет [был] Охозия, когда воцарился, и один год царствовал в Иерусалиме; имя матери его Гофолия, дочь Амврия.
2CHR|22|3|Он также ходил путями дома Ахавова, потому что мать его была советницею ему на беззаконные дела.
2CHR|22|4|И делал он неугодное в очах Господних, подобно дому Ахавову, потому что он был ему советником, по смерти отца его, на погибель ему.
2CHR|22|5|Также следуя их совету, он пошел с Иорамом, сыном Ахавовым, царем Израильским, на войну против Азаила, царя Сирийского, в Рамоф Галаадский. И ранили Сирияне Иорама,
2CHR|22|6|и возвратился он в Изреель лечиться от ран, которые причинили ему в Раме, когда он воевал с Азаилом, царем Сирийским. И Охозия, сын Иорама, царь Иудейский, пришел посетить Иорама, сына Ахавова, в Изреель, потому что тот был болен.
2CHR|22|7|И от Бога было это на погибель Охозии, что он пришел к Иораму: ибо, по приходе своем, он вышел с Иорамом против Ииуя, сына Намессиева, которого помазал Господь на истребление дома Ахавова.
2CHR|22|8|Когда совершал Ииуй суд над домом Ахава, тогда он нашел князей Иудийских и сыновей братьев Охозии, служивших Охозии, и умертвил их.
2CHR|22|9|И [велел] он искать Охозию, и взяли его, когда он скрывался в Самарии, и привели его к Ииую, и умертвили его, и похоронили его, ибо говорили: он сын Иосафата, который взыскал Господа от всего сердца своего. И не [осталось] в доме Охозии, [кто] мог бы царствовать.
2CHR|22|10|Ибо Гофолия, мать Охозии, увидев, что умер сын ее, встала и истребила все царское племя дома Иудина.
2CHR|22|11|Но Иосавеф, дочь царя, взяла Иоаса, сына Охозии, и похитила его из среды царских сыновей умерщвляемых, и поместила его и кормилицу его в спальной комнате; и таким образом Иосавеф, дочь царя Иорама, жена Иодая священника, сестра Охозии, скрыла Иоаса от Гофолии, и она не умертвила его.
2CHR|22|12|И был он у них в доме Божием скрываем шесть лет; Гофолия же царствовала над землею.
2CHR|23|1|Но в седьмой год ободрился Иодай и принял в союз с собою начальников сотен: Азарию, сына Иерохамова, и Исмаила, сына Иегохананова, и Азарию, сына Оведова, и Маасею, сына Адаии, и Елишафата, сына Зихри.
2CHR|23|2|И они прошли по Иудее и собрали левитов из всех городов Иудеи и глав поколений Израилевых, и пришли в Иерусалим.
2CHR|23|3|И заключило все собрание союз в доме Божием с царем. И сказал им [Иодай]: вот сын царя должен быть царем, как изрек Господь о сыновьях Давидовых.
2CHR|23|4|Вот что вы сделайте: треть вас, приходящих в субботу, из священников и левитов, [будет] привратниками у порогов,
2CHR|23|5|и треть при доме царском, и треть у ворот Иесод, а весь народ на дворах дома Господня.
2CHR|23|6|И [никто] пусть не входит в дом Господень, кроме священников и служащих из левитов. Они могут войти, потому что освящены; весь же народ пусть стоит на страже Господней.
2CHR|23|7|И пусть левиты окружат царя со всех сторон, всякий с оружием своим в руке своей, и кто будет входить в храм, да будет умерщвлен. И будьте вы при царе, когда он будет входить и выходить.
2CHR|23|8|И сделали левиты и все Иудеи, что приказал Иодай священник; и взяли каждый людей своих, приходящих в субботу с отходящими в субботу, потому что не отпустил священник Иодай [сменившихся] черед.
2CHR|23|9|И роздал Иодай священник начальникам сотен копья и малые и большие щиты царя Давида, которые [были] в доме Божием;
2CHR|23|10|и поставил весь народ, каждого с оружием его в руке его, от правой стороны храма до левой стороны храма, у жертвенника и у дома, вокруг царя.
2CHR|23|11|И вывели сына царя, и возложили на него венец и украшения, и поставили его царем; и помазали его Иодай и сыновья его и сказали: да живет царь!
2CHR|23|12|И услышала Гофолия голос народа, бегущего и провозглашающего о царе, и вышла к народу в дом Господень,
2CHR|23|13|и увидела: и вот царь стоит на возвышении своем при входе, и князья и трубы подле царя, и весь народ земли веселится, и трубят трубами, и певцы с орудиями музыкальными и искусные в славословии. И разодрала Гофолия одежды свои и закричала: заговор! заговор!
2CHR|23|14|И вызвал Иодай священник начальников сотен, начальствующих над войском, и сказал им: выведите ее вон, и, кто последует за нею, да будет умерщвлен мечом. Потому что священник сказал: не умертвите ее в доме Господнем.
2CHR|23|15|И дали ей место, и когда она пришла ко входу конских ворот царского дома, там умертвили ее.
2CHR|23|16|И заключил Иодай завет между собою и между всем народом и царем, чтобы быть [им] народом Господним.
2CHR|23|17|И пошел весь народ в капище Ваала, и разрушили его, и жертвенники его и истуканов его сокрушили; и Матфана, жреца Ваалова, умертвили пред жертвенниками.
2CHR|23|18|И поручил Иодай дела дома Господня священникам и левитам, как распределил Давид в доме Господнем, для возношения всесожжений Господу, как написано в законе Моисеевом, с радостью и пением, по уставу Давидову.
2CHR|23|19|И поставил он привратников у ворот дома Господня, чтобы не [мог] входить нечистый почему–нибудь.
2CHR|23|20|И взял начальников сотен, и вельмож, и начальствующих в народе, и весь народ земли, и проводил царя из дома Господня, и прошли чрез верхние ворота в дом царский, и посадили царя на царский престол.
2CHR|23|21|И веселился весь народ земли, и город успокоился. А Гофолию умертвили мечом.
2CHR|24|1|Семи лет [был] Иоас, когда воцарился, и сорок лет царствовал в Иерусалиме; имя матери его Цивья из Вирсавии.
2CHR|24|2|И делал Иоас угодное в очах Господних во все дни Иодая священника.
2CHR|24|3|И взял ему Иодай двух жен, и он имел [от них] сыновей и дочерей.
2CHR|24|4|И после сего пришло на сердце Иоасу обновить дом Господень,
2CHR|24|5|и собрал он священников и левитов и сказал им: пойдите по городам Иудеи и собирайте со всех Израильтян серебро для поддержания дома Бога вашего из года в год, и поспешите в этом деле. Но не поспешили левиты.
2CHR|24|6|И призвал царь Иодая, главу [их], и сказал ему: почему ты не требуешь от левитов, чтобы они доставляли с Иудеи и Иерусалима дань, [установленную] Моисеем, рабом Господним, и собранием Израильтян для скинии собрания?
2CHR|24|7|Ибо нечестивая Гофолия и сыновья ее разорили дом Божий и все посвященное для дома Господня употребили для Ваалов.
2CHR|24|8|И приказал царь, и сделали один ящик, и поставили его у входа в дом Господень извне.
2CHR|24|9|И провозгласили по Иудее и Иерусалиму, чтобы приносили Господу дань, [наложенную] Моисеем, рабом Божиим, на Израильтян в пустыне.
2CHR|24|10|И обрадовались все начальствующие и весь народ, и приносили и клали в ящик дотоле, доколе он не наполнился.
2CHR|24|11|В то время, когда приносили ящик к царским чиновникам чрез левитов, и когда они видели, что серебра много, приходил писец царя и поверенный первосвященника, и высыпали из ящика, и относили его и ставили его на свое место. Так делали они изо дня в день, и собрали множество серебра.
2CHR|24|12|И отдавали его царь и Иодай производителям работ по дому Господню, и они нанимали каменотесов и плотников для подновления дома Господня, также кузнецов и медников для укрепления дома Господня.
2CHR|24|13|И работали производители работ, и совершилось исправление руками их, и привели дом Божий в надлежащее состояние его, и укрепили его.
2CHR|24|14|И кончив [все], они представили царю и Иодаю остаток серебра. И сделали из него сосуды для дома Господня, сосуды служебные и [для] всесожжений, чаши и [другие] сосуды золотые и серебряные. И приносили всесожжения в доме Господнем постоянно во все дни Иодая.
2CHR|24|15|И состарился Иодай и, насытившись днями [жизни], умер: сто тридцать лет [было] ему, когда он умер.
2CHR|24|16|И похоронили его в городе Давидовом с царями, потому что он делал доброе в Израиле и для Бога, и для дома Его.
2CHR|24|17|Но по смерти Иодая пришли князья Иудейские и поклонились царю; тогда царь стал слушаться их.
2CHR|24|18|И оставили дом Господа Бога отцов своих и стали служить деревам [посвященным] и идолам, – и был гнев [Господень] на Иуду и Иерусалим за сию вину их.
2CHR|24|19|И он посылал к ним пророков для обращения их к Господу, и они увещевали их, но те не слушали.
2CHR|24|20|И Дух Божий облек Захарию, сына Иодая священника, и он стал на возвышении пред народом и сказал им: так говорит Господь: для чего вы преступаете повеления Господни? не будет успеха вам; и как вы оставили Господа, то и Он оставит вас.
2CHR|24|21|И сговорились против него, и побили его камнями, по приказанию царя, на дворе дома Господня.
2CHR|24|22|И не вспомнил царь Иоас благодеяния, какое сделал ему Иодай, отец его, и убил сына его. И он умирая говорил: да видит Господь и да взыщет!
2CHR|24|23|И по истечении года выступило против него войско Сирийское, и вошли в Иудею и в Иерусалим, и истребили из народа всех князей народа, и всю добычу, [взятую] у них, отослали к царю в Дамаск.
2CHR|24|24|Хотя в небольшом числе людей приходило войско Сирийское, но Господь предал в руку их весьма многочисленную силу за то, что оставили Господа Бога отцов своих. И над Иоасом совершили они суд,
2CHR|24|25|и когда они ушли от него, оставив его в тяжкой болезни, то составили против него заговор рабы его, за кровь сына Иодая священника, и убили его на постели его, и он умер. И похоронили его в городе Давидовом, но не похоронили его в царских гробницах.
2CHR|24|26|Заговорщиками же против него были: Завад, сын Шимеафы Аммонитянки, и Иегозавад, сын Шимрифы Моавитянки.
2CHR|24|27|О сыновьях его и о множестве пророчеств против него и об устроении дома Божия написано в книге царей. И воцарился Амасия, сын его, вместо него.
2CHR|25|1|Двадцати пяти лет воцарился Амасия и двадцать девять лет царствовал в Иерусалиме; имя матери его Иегоаддань из Иерусалима.
2CHR|25|2|И делал он угодное в очах Господних, но не от полного сердца.
2CHR|25|3|Когда утвердилось за ним царство, тогда он умертвил рабов своих, убивших царя, отца его.
2CHR|25|4|Но детей их не умертвил, так как написано в законе, в книге Моисеевой, где заповедал Господь, говоря: не должны быть умерщвляемы отцы за детей, и дети не должны быть умерщвляемы за отцов, но каждый за свое преступление должен умереть.
2CHR|25|5|И собрал Амасия Иудеев и поставил их по поколениям под власть тысяченачальников и стоначальников, всех Иудеев и Вениаминян, и пересчитал их от двадцати лет и выше, и нашел их триста тысяч человек отборных, ходящих на войну, держащих копье и щит.
2CHR|25|6|И [еще] нанял из Израильтян сто тысяч храбрых воинов за сто талантов серебра.
2CHR|25|7|Но человек Божий пришел к нему и сказал: царь! пусть не идет с тобою войско Израильское, потому что нет Господа с Израильтянами, со всеми сынами Ефрема.
2CHR|25|8|Но иди ты [один], делай дело, мужественно подвизайся на войне. [Иначе] повергнет тебя Бог пред лицем врага, ибо есть сила у Бога поддержать и повергнуть.
2CHR|25|9|И сказал Амасия человеку Божию: что же делать со ста талантами, которые я отдал войску Израильскому? И сказал человек Божий: может Господь дать тебе более сего.
2CHR|25|10|И отделил их Амасия, – войско, пришедшее к нему из [земли] Ефремовой, – чтоб они шли в свое место. И возгорелся сильно гнев их на Иудею, и они пошли назад в свое место, в пылу гнева.
2CHR|25|11|А Амасия отважился и повел народ свой, и пошел на долину Соляную и побил сынов Сеира десять тысяч;
2CHR|25|12|и десять тысяч живых взяли сыны Иудины в плен, и привели их на вершину скалы, и низринули их с вершины скалы, и все они разбились совершенно.
2CHR|25|13|Войско же, которое Амасия отослал обратно, чтоб оно не ходило с ним на войну, рассыпалось по городам Иудеи от Самарии до Вефорона и перебило в них три тысячи, и награбило множество добычи.
2CHR|25|14|Амасия, придя после поражения Идумеян, принес богов сынов Сеира и поставил их у себя богами, и пред ними кланялся и им кадил.
2CHR|25|15|И воспылал гнев Господа на Амасию, и послал Он к нему пророка, и тот сказал ему: зачем ты прибегаешь к богам народа сего, которые не избавили народа своего от руки твоей?
2CHR|25|16|Когда он говорил ему, [царь] отвечал: разве советником царским поставили тебя? перестань, чтобы не убили тебя. И перестал пророк, сказав: знаю, что решил Бог погубить тебя, потому что ты сделал сие и не слушаешь совета моего.
2CHR|25|17|И посоветовался Амасия, царь Иудейский, и послал к Иоасу, сыну Иоахаза, сына Ииуева, царю Израильскому, сказать: выходи, повидаемся лично.
2CHR|25|18|И послал Иоас, царь Израильский, к Амасии, царю Иудейскому, сказать: терн, который на Ливане, послал к кедру, который на Ливане же, сказать: отдай дочь свою в жену сыну моему. Но прошли звери дикие, которые на Ливане, и истоптали этот терн.
2CHR|25|19|Ты говоришь: вот я побил Идумеян, – и вознеслось сердце твое до тщеславия. Сиди лучше у себя дома. К чему тебе затевать опасное дело? Падешь ты и Иудея с тобою.
2CHR|25|20|Но не послушался Амасия, так как от Бога [было] это, дабы предать их в руку [Иоаса] за то, что стали прибегать к богам Идумейским.
2CHR|25|21|И выступил Иоас, царь Израильский, и увиделись лично, он и Амасия, царь Иудейский, в Вефсамисе Иудейском.
2CHR|25|22|И были разбиты Иудеи Израильтянами, и разбежались каждый в шатер свой.
2CHR|25|23|И Амасию, царя Иудейского, сына Иоаса, сына Иоахазова, захватил Иоас, царь Израильский, в Вефсамисе и привел его в Иерусалим, и разрушил стену Иерусалимскую от ворот Ефремовых до ворот угольных, на четыреста локтей;
2CHR|25|24|и [взял] все золото и серебро, и все сосуды, находившиеся в доме Божием у Овед–Едома, и сокровища дома царского, и заложников, и возвратился в Самарию.
2CHR|25|25|И жил Амасия, сын Иоасов, царь Иудейский, по смерти Иоаса, сына Иоахазова, царя Израильского, пятнадцать лет.
2CHR|25|26|Прочие дела Амасии, первые и последние, описаны в книге царей Иудейских и Израильских.
2CHR|25|27|И после того времени, как Амасия отступил от Господа, составили против него заговор в Иерусалиме, и он убежал в Лахис. И послали за ним в Лахис, и умертвили его там.
2CHR|25|28|И привезли его на конях, и похоронили его с отцами его в городе Иудином.
2CHR|26|1|И взял весь народ Иудейский Озию, которому [было] шестнадцать лет, и поставили его царем на место отца его Амасии.
2CHR|26|2|Он обстроил Елаф и возвратил его Иудее, после того как почил царь с отцами своими.
2CHR|26|3|Шестнадцати лет [был] Озия, когда воцарился, и пятьдесят два года царствовал в Иерусалиме; имя матери его Иехолия из Иерусалима.
2CHR|26|4|И делал он угодное в очах Господних точно так, как делал Амасия, отец его;
2CHR|26|5|и прибегал он к Богу во дни Захарии, поучавшего страху Божию; и в те дни, когда он прибегал к Господу, споспешествовал ему Бог.
2CHR|26|6|И он вышел и сразился с Филистимлянами, и разрушил стены Гефа и стены Иавнеи и стены Азота; и построил города в [области] Азотской и у Филистимлян.
2CHR|26|7|И помогал ему Бог против Филистимлян и против Аравитян, живущих в Гур–Ваале, и [против] Меунитян;
2CHR|26|8|и давали Аммонитяне дань Озии, и дошло имя его до пределов Египта, потому что он был весьма силен.
2CHR|26|9|И построил Озия башни в Иерусалиме над воротами угольными и над воротами долины и на углу, и укрепил их.
2CHR|26|10|И построил башни в пустыне, и иссек много водоемов, потому что имел много скота, и на низменности и на равнине, и земледельцев и садовников на горах и на Кармиле, ибо он любил земледелие.
2CHR|26|11|Было у Озии и войско, выходившее на войну отрядами, по счету в списке их, составленном рукою Иеиела писца и Маасеи надзирателя, под предводительством Ханании, [одного] из главных сановников царских.
2CHR|26|12|Все число глав поколений, из храбрых воинов, [было] две тысячи шестьсот,
2CHR|26|13|и под рукою их военной силы триста семь тысяч пятьсот, вступавших в сражение с воинским мужеством, на помощь царю против неприятеля.
2CHR|26|14|И заготовил для них Озия, для всего войска, щиты и копья, и шлемы и латы, и луки и пращные камни.
2CHR|26|15|И сделал он в Иерусалиме искусно придуманные машины, чтоб они находились на башнях и на углах для метания стрел и больших камней. И пронеслось имя его далеко, потому что он дивно оградил себя и сделался силен.
2CHR|26|16|Но когда он сделался силен, возгордилось сердце его на погибель [его], и он сделался преступником пред Господом Богом своим, ибо вошел в храм Господень, чтобы воскурить [фимиам] на алтаре кадильном.
2CHR|26|17|И пошел за ним Азария священник, и с ним восемьдесят священников Господних, людей отличных,
2CHR|26|18|и воспротивились Озии царю и сказали ему: не тебе, Озия, кадить Господу; это [дело] священников, сынов Аароновых, посвященных для каждения; выйди из святилища, ибо ты поступил беззаконно, и не [будет] тебе это в честь у Господа Бога.
2CHR|26|19|И разгневался Озия, – а в руке у него кадильница для каждения; и когда разгневался он на священников, проказа явилась на челе его, пред лицем священников, в доме Господнем, у алтаря кадильного.
2CHR|26|20|И взглянул на него Азария первосвященник и все священники; и вот у него проказа на челе его. И понуждали его выйти оттуда, да и сам он спешил удалиться, так как поразил его Господь.
2CHR|26|21|И был царь Озия прокаженным до дня смерти своей, и жил в отдельном доме и отлучен был от дома Господня. А Иоафам, сын его, начальствовал над домом царским и управлял народом земли.
2CHR|26|22|Прочие деяния Озии, первые и последние, описал Исаия, сын Амоса, пророк.
2CHR|26|23|И почил Озия с отцами своими, и похоронили его с отцами его на поле царских гробниц, ибо говорили: он прокаженный. И воцарился Иоафам, сын его, вместо него.
2CHR|27|1|Двадцати пяти лет [был] Иоафам, когда воцарился, и шестнадцать лет царствовал в Иерусалиме; имя матери его Иеруша, дочь Садока.
2CHR|27|2|И делал он угодное в очах Господних точно так, как делал Озия, отец его, только он не входил в храм Господень, и народ продолжал еще грешить.
2CHR|27|3|Он построил верхние ворота дома Господня, и многое построил на стене Офела;
2CHR|27|4|и города построил на горе Иудейской, и в лесах построил дворцы и башни.
2CHR|27|5|Он воевал с царем Аммонитян и одолел их, и дали ему Аммонитяне в тот год сто талантов серебра и десять тысяч коров пшеницы и ячменя десять тысяч. Это давали ему Аммонитяне и на другой год, и на третий.
2CHR|27|6|Так силен был Иоафам потому, что устроял пути свои пред лицем Господа Бога своего.
2CHR|27|7|Прочие деяния Иоафама и все войны его и поведение его описаны в книге царей Израильских и Иудейских:
2CHR|27|8|двадцати пяти лет был он, когда воцарился, и шестнадцать лет царствовал в Иерусалиме.
2CHR|27|9|И почил Иоафам с отцами своими, и похоронили его в городе Давидовом. И воцарился Ахаз, сын его, вместо него.
2CHR|28|1|Двадцати лет был Ахаз, когда воцарился, и шестнадцать лет царствовал в Иерусалиме; и он не делал угодного в очах Господних, как [делал] Давид, отец его:
2CHR|28|2|он шел путями царей Израильских, и даже сделал литые статуи Ваалов;
2CHR|28|3|и он совершал курения на долине сынов Еннома, и проводил сыновей своих через огонь, подражая мерзостям народов, которых изгнал Господь пред лицем сынов Израилевых;
2CHR|28|4|и приносил жертвы и курения на высотах и на холмах и под всяким ветвистым деревом.
2CHR|28|5|И предал его Господь Бог его в руку царя Сириян, и они поразили его и взяли у него множество пленных и отвели в Дамаск. Также и в руку царя Израильского был предан он, и тот произвел у него великое поражение.
2CHR|28|6|И избил Факей, сын Ремалиин, Иудеев сто двадцать тысяч в один день, людей воинственных, потому что они оставили Господа Бога отцов своих.
2CHR|28|7|Зихрий же, силач из Ефремлян, убил Маасею, сына царя, и Азрикама, начальствующего над дворцом, и Елкану, второго по царе.
2CHR|28|8|И взяли сыны Израилевы в плен у братьев своих, [Иудеев], двести тысяч жен, сыновей и дочерей; также и множество добычи награбили у них, и отправили добычу в Самарию.
2CHR|28|9|Там был пророк Господень, имя его Одед. Он вышел пред лице войска, шедшего в Самарию, и сказал им: вот Господь Бог отцов ваших, во гневе на Иудеев, предал их в руку вашу, и вы избили их с такою яростью, которая достигла до небес.
2CHR|28|10|И теперь вы думаете поработить сынов Иуды и Иерусалима в рабы и рабыни себе. А разве на самих вас нет вины пред Господом Богом вашим?
2CHR|28|11|Итак послушайте меня, и возвратите пленных, которых вы захватили из братьев ваших, ибо пламень гнева Господня на вас.
2CHR|28|12|И встали некоторые из начальников сынов Ефремовых: Азария, сын Иегоханана, Берехия, сын Мешиллемофа, и Езекия, сын Шаллума, и Амаса, сын Хадлая, против шедших с войны,
2CHR|28|13|и сказали им: не вводите сюда пленных, потому что грех был бы нам пред Господом. Неужели вы думаете прибавить к грехам нашим и к преступлениям нашим? велика вина наша, и пламень гнева [Господня] над Израилем.
2CHR|28|14|И оставили вооруженные пленных и добычу у военачальников и всего собрания.
2CHR|28|15|И встали мужи, упомянутые по именам, и взяли пленных, и всех нагих из них одели из добычи, – и одели их, и обули их, и накормили их, и напоили их, и помазали их елеем, и посадили на ослов всех слабых из них, и отправили их в Иерихон, город пальм, к братьям их, и возвратились в Самарию.
2CHR|28|16|В то время послал царь Ахаз к царям Ассирийским, чтоб они помогли ему,
2CHR|28|17|ибо Идумеяне и еще приходили, и [многих] побили в Иудее, и взяли в плен;
2CHR|28|18|и Филистимляне рассыпались по городам низменного края и юга Иудеи и взяли Вефсамис и Аиалон, и Гедероф и Сохо и зависящие от него города, и Фимну и зависящие от нее города, и Гимзо и зависящие от него города, и поселились там.
2CHR|28|19|Так унизил Господь Иудею за Ахаза, царя Иудейского, потому что он развратил Иудею и тяжко грешил пред Господом.
2CHR|28|20|И пришел к нему Феглафелласар, царь Ассирийский, но был в тягость ему, вместо того, чтобы помочь ему,
2CHR|28|21|потому что Ахаз взял [сокровища] из дома Господня и дома царского и у князей и отдал царю Ассирийскому, но не в помощь себе.
2CHR|28|22|И в тесное для себя время он продолжал беззаконно поступать пред Господом, он – царь Ахаз.
2CHR|28|23|И приносил он жертвы богам Дамасским, [думая, что] они поражали его, и говорил: боги царей Сирийских помогают им; принесу я жертву им, и они помогут мне. Но они были на падение ему и всему Израилю.
2CHR|28|24|И собрал Ахаз сосуды дома Божия, и сокрушил сосуды дома Божия, и запер двери дома Господня, и устроил себе жертвенники по всем углам в Иерусалиме,
2CHR|28|25|и по всем городам Иудиным устроил высоты для каждения богам иным, и раздражал Господа Бога отцов своих.
2CHR|28|26|Прочие дела его и все поступки его, первые и последние, описаны в книге царей Иудейских и Израильских.
2CHR|28|27|И почил Ахаз с отцами своими, и похоронили его в городе, в Иерусалиме, но не внесли его в гробницы царей Израилевых. И воцарился Езекия, сын его, вместо него.
2CHR|29|1|Езекия воцарился двадцати пяти лет, и двадцать девять лет царствовал в Иерусалиме; имя матери его Авия, дочь Захарии.
2CHR|29|2|И делал он угодное в очах Господних точно так, как делал Давид, отец его.
2CHR|29|3|В первый же год царствования своего, в первый месяц, он отворил двери дома Господня и возобновил их,
2CHR|29|4|и велел прийти священникам и левитам, и собрал их на площади восточной,
2CHR|29|5|и сказал им: послушайте меня, левиты! Ныне освятитесь [сами] и освятите дом Господа Бога отцов ваших, и выбросьте нечистоту из святилища.
2CHR|29|6|Ибо отцы наши поступали беззаконно, и делали неугодное в очах Господа Бога нашего, и оставили Его, и отвратили они лица свои от жилища Господня, и оборотились спиною,
2CHR|29|7|и заперли двери притвора, и погасили светильники, и не сожигали курения, и не возносили всесожжений во святилище Бога Израилева.
2CHR|29|8|И был гнев Господа на Иудею и на Иерусалим, и Он отдал их на позор, на опустошение и на посмеяние, как вы видите глазами вашими.
2CHR|29|9|И вот, пали отцы наши от меча, а сыновья наши и дочери наши и жены наши за это в плену доныне.
2CHR|29|10|Теперь у меня на сердце – заключить завет с Господом Богом Израилевым, да отвратит от нас пламень гнева Своего.
2CHR|29|11|Дети мои! не будьте небрежны, ибо вас избрал Господь предстоять лицу Его, служить Ему и быть у Него служителями и возжигателями курений.
2CHR|29|12|И встали левиты: Махаф, сын Амасая, и Иоель, сын Азарии, из сыновей Каафовых; и из сыновей Мерариных: Кис, сын Авдия, и Азария, сын Иегаллелела; и из племени Гирсонова: Иоах, сын Зиммы, и Еден, сын Иоаха;
2CHR|29|13|и из сыновей Елицафановых: Шимри и Иеиел; и из сыновей Асафовых: Захария и Матфания;
2CHR|29|14|и из сыновей Емановых: Иехиел и Шимей; и из сыновей Идифуновых: Шемаия и Уззиел.
2CHR|29|15|Они собрали братьев своих и освятились, и пошли по приказанию царя очищать дом Господень по словам Господа.
2CHR|29|16|И вошли священники внутрь дома Господня для очищения, и вынесли все нечистое, что нашли в храме Господнем, на двор дома Господня, а левиты взяли это, чтобы вынести вон к потоку Кедрону.
2CHR|29|17|И начали освящать в первый [день] первого месяца, и в восьмой день [того же] месяца вошли в притвор Господень; и освящали дом Господень восемь дней, и в шестнадцатый день первого месяца кончили.
2CHR|29|18|И пришли в дом к царю Езекии и сказали: мы очистили дом Господень, и жертвенник для всесожжения, и все сосуды его, и стол [для хлебов] предложения, и все сосуды его;
2CHR|29|19|и все сосуды, которые забросил царь Ахаз во время царствования своего, в беззаконии своем, мы приготовили и освятили, и вот они пред жертвенником Господним.
2CHR|29|20|И встал царь Езекия рано утром и собрал начальников города, и пошел в дом Господень.
2CHR|29|21|И привели семь тельцов и семь овнов, и семь агнцев и семь козлов на жертву о грехе за царство и за святилище и за Иудею; и приказал он сынам Аароновым, священникам, вознести всесожжение на жертвенник Господень.
2CHR|29|22|И закололи тельцов, и взяли священники кровь, и окропили жертвенник, и закололи овнов, и окропили кровью жертвенник; и закололи агнцев, и окропили кровью жертвенник.
2CHR|29|23|И привели козлов за грех пред лице царя и собрания, и они возложили руки свои на них.
2CHR|29|24|И закололи их священники, и очистили кровью их жертвенник для заглаждения грехов всего Израиля, ибо за всего Израиля приказал царь [принести] всесожжение и жертву о грехе.
2CHR|29|25|И поставил он левитов в доме Господнем с кимвалами, псалтирями и цитрами, по уставу Давида и Гада, прозорливца царева, и Нафана пророка, так как от Господа [был] устав этот чрез пророков Его.
2CHR|29|26|И стали левиты с [музыкальными] орудиями Давидовыми и священники с трубами.
2CHR|29|27|И приказал Езекия вознести всесожжение на жертвенник. И в то время, как началось всесожжение, началось пение Господу, при [звуке] труб и орудий Давида, царя Израилева.
2CHR|29|28|И все собрание молилось, и певцы пели, и трубили трубы, доколе не окончилось всесожжение.
2CHR|29|29|По окончании же всесожжения царь и все находившиеся при нем преклонились и поклонились.
2CHR|29|30|И сказал царь Езекия и князья левитам, чтоб они славили Господа словами Давида и Асафа прозорливца, и они славили с радостью и преклонялись и поклонялись.
2CHR|29|31|И продолжал Езекия и сказал: теперь вы посвятили себя Господу; приступайте и приносите жертвы и благодарственные приношения в дом Господень. И понесло [все] собрание жертвы и благодарственные приношения, и всякий, кто расположен был сердцем, – всесожжения.
2CHR|29|32|И было число всесожжений, которые привели собравшиеся: семьдесят волов, сто овнов, двести агнцев – все это для всесожжения Господу.
2CHR|29|33|[Других] священных жертв [было]: шестьсот из крупного скота и три тысячи из мелкого скота.
2CHR|29|34|Но священников было мало, и они не могли сдирать кож со всех всесожжений, и помогали им братья их левиты, до окончания дела и доколе освятились [прочие] священники, ибо левиты были более тщательны в освящении себя, нежели священники.
2CHR|29|35|Притом же всесожжений [было] множество с туками мирных жертв и с возлияниями при всесожжении. Так восстановлено служение в доме Господнем.
2CHR|29|36|И радовался Езекия и весь народ о том, что Бог [так] расположил народ, ибо это сделалось неожиданно.
2CHR|30|1|И послал Езекия по всей [земле] Израильской и Иудее, и письма писал к Ефрему и Манассии, чтобы пришли в дом Господень, в Иерусалим, для совершения пасхи Господу Богу Израилеву.
2CHR|30|2|И положили на совете царь и князья его и все собрание в Иерусалиме – совершить пасху во второй месяц,
2CHR|30|3|ибо не могли совершить ее в свое время, потому что священники [еще] не освятились в достаточном числе и народ не собрался в Иерусалим.
2CHR|30|4|И понравилось это царю и всему собранию.
2CHR|30|5|И определили объявить по всему Израилю, от Вирсавии до Дана, чтобы шли в Иерусалим для совершения пасхи Господу Богу Израилеву, потому что давно не совершали [ее], как предписано.
2CHR|30|6|И пошли гонцы с письмами от царя и от князей его по всей [земле] Израильской и Иудее, и по повелению царя говорили: дети Израиля! обратитесь к Господу Богу Авраама, Исаака и Израиля, и Он обратится к остатку, уцелевшему у вас от руки царей Ассирийских.
2CHR|30|7|И не будьте таковы, как отцы ваши и братья ваши, которые беззаконно поступали пред Господом Богом отцов своих; и Он предал их на опустошение, как вы видите.
2CHR|30|8|Ныне не будьте жестоковыйны, как отцы ваши, покоритесь Господу и приходите во святилище Его, которое Он освятил навек; и служите Господу Богу вашему, и Он отвратит от вас пламень гнева Своего.
2CHR|30|9|Когда вы обратитесь к Господу, тогда братья ваши и дети ваши [будут] в милости у пленивших их и возвратятся в землю сию, ибо благ и милосерд Господь Бог ваш и не отвратит лица от вас, если вы обратитесь к Нему.
2CHR|30|10|И ходили гонцы из города в город по земле Ефремовой и Манассииной и до Завулоновой, но над ними смеялись и издевались.
2CHR|30|11|Однако некоторые из [колена] Асирова, Манассиина и Завулонова смирились и пришли в Иерусалим.
2CHR|30|12|И над Иудеею была рука Божия, даровавшая им единое сердце, чтоб исполнить повеление царя и князей, по слову Господню.
2CHR|30|13|И собралось в Иерусалим множество народа для совершения праздника опресноков, во второй месяц, – собрание весьма многочисленное.
2CHR|30|14|И встали и ниспровергли жертвенники, которые были в Иерусалиме; и все, на чем совершаемо было курение [идолам], разрушили и бросили в поток Кедрон;
2CHR|30|15|и закололи пасхального агнца в четырнадцатый [день] второго месяца. Священники и левиты устыдившись освятились и принесли всесожжения в дом Господень,
2CHR|30|16|и стали на своем месте по уставу своему, по закону Моисея, человека Божия. Священники кропили кровью [принимая ее] из рук левитов.
2CHR|30|17|Так как много [было] в собрании таких, которые не освятились, то вместо нечистых левиты закололи пасхального агнца, для посвящения Господу.
2CHR|30|18|Многие из народа, большею частью из колена Ефремова и Манассиина, Иссахарова и Завулонова, не очистились; однакоже они ели пасху, не по уставу.
2CHR|30|19|Но Езекия помолился за них, говоря: Господь благий да простит каждого, кто расположил сердце свое к тому, чтобы взыскать Господа Бога, Бога отцов своих, хотя и без очищения священного!
2CHR|30|20|И услышал Господь Езекию и простил народ.
2CHR|30|21|И совершили сыны Израилевы, находившиеся в Иерусалиме, праздник опресноков в семь дней, с великим веселием; каждый день левиты и священники славили Господа на орудиях, [устроенных] для славословия Господа.
2CHR|30|22|И говорил Езекия по сердцу всем левитам, имевшим доброе разумение [в служении] Господу. И ели праздничное семь дней, принося жертвы мирные и славя Господа Бога отцов своих.
2CHR|30|23|И решило все собрание праздновать другие семь дней, и провели эти семь дней в веселии,
2CHR|30|24|потому что Езекия, царь Иудейский, выставил для собравшихся тысячу тельцов и десять тысяч мелкого скота, и вельможи выставили для собравшихся тысячу тельцов и десять тысяч мелкого скота; и священников освятилось [уже] много.
2CHR|30|25|И веселились все собравшиеся из Иудеи, и священники и левиты, и все собрание, пришедшее от Израиля, и пришельцы, пришедшие из земли Израильской и обитавшие в Иудее.
2CHR|30|26|И было веселие великое в Иерусалиме, потому что со дней Соломона, сына Давидова, царя Израилева, [не бывало] подобного сему в Иерусалиме.
2CHR|30|27|И встали священники и левиты, и благословили народ; и услышан был голос их, и взошла молитва их в святое жилище Его на небеса.
2CHR|31|1|И по окончании всего этого, пошли все Израильтяне, [там] находившиеся, в города Иудейские и разбили статуи, срубили [посвященные] дерева, и разрушили высоты и жертвенники во всей Иудее и в [земле] Вениаминовой, Ефремовой и Манассииной, до конца. И [потом] возвратились все сыны Израилевы, каждый во владение свое, в города свои.
2CHR|31|2|И поставил Езекия череды священников и левитов, по их распределению, каждого при деле своем, священническом или левитском, при всесожжении и при жертвах мирных, для службы, для хваления и славословия, у ворот дома Господня.
2CHR|31|3|И [определил] царь часть из имущества своего на всесожжения: на всесожжения утренние и вечерние, и на всесожжения в субботы и в новомесячия, и в праздники, как написано в законе Господнем.
2CHR|31|4|И повелел он народу, живущему в Иерусалиме, давать определенное содержание священникам и левитам, чтоб они были ревностны в законе Господнем.
2CHR|31|5|Когда обнародовано было это повеление, тогда нанесли сыны Израилевы множество начатков хлеба, вина, и масла, и меду, и всяких произведений полевых; и десятин из всего нанесли множество.
2CHR|31|6|И Израильтяне и Иудеи, живущие по городам Иудейским, также представили десятины из крупного и мелкого скота и десятины из пожертвований, посвященных Господу Богу их; и наложили груды, груды.
2CHR|31|7|В третий месяц начали класть груды, и в седьмой месяц кончили.
2CHR|31|8|И пришли Езекия и вельможи, и увидели груды, и благодарили Господа и народ Его Израиля.
2CHR|31|9|И спросил Езекия священников и левитов об этих грудах.
2CHR|31|10|И отвечал ему Азария первосвященник из дома Садокова и сказал: с того времени, как начали носить приношения в дом Господень, мы ели досыта, и многое осталось, потому что Господь благословил народ Свой. Из оставшегося [составилось] такое множество.
2CHR|31|11|И приказал Езекия приготовить комнаты при доме Господнем. И приготовили.
2CHR|31|12|И перенесли [туда] приношения, и десятины, и пожертвования, со [всею] точностью. И [был] начальником при них Хонания левит, и Симей, брат его, вторым.
2CHR|31|13|А Иехиил и Азазия, и Нахаф и Асаил, и Иеримоф и Иозавад, и Елиел и Исмахия, и Махаф и Бенания [были] смотрителями под рукою Хонании и Симея, брата его, по распоряжению царя Езекии и Азарии, начальника при доме Божием.
2CHR|31|14|Коре, сын Имны, левит, привратник на восточной стороне, [был] при добровольных приношениях Богу, для выдачи принесенного Господу и важнейших из вещей посвященных.
2CHR|31|15|И под его [ведением находились] Еден, и Миниамин, и Иешуа, и Шемаия, и Амария и Шехания в городах священнических, чтобы верно раздавать братьям своим части, как большому, так и малому,
2CHR|31|16|сверх списка их, [всем] мужеского пола от трех лет и выше, всем ходящим в дом Господа для дел ежедневных, для служения их, по должностям их и по отделам их,
2CHR|31|17|и внесенным в список священникам, по поколениям их, и левитам от двадцати лет и выше, по должностям их, по отделам их,
2CHR|31|18|и внесенным в список, со всеми малолетними их, с женами их и с сыновьями их и с дочерями их, – всему обществу, ибо они со [всею] верностью посвятили себя на священную службу.
2CHR|31|19|И для сынов Аароновых, священников в селениях вокруг городов их, при каждом городе [поставлены были] мужи поименованные, чтобы раздавать участки всем мужеского пола у священников и всем внесенным в список у левитов.
2CHR|31|20|Вот что сделал Езекия во всей Иудее, – и он делал доброе, и справедливое, и истинное пред лицем Господа Бога своего.
2CHR|31|21|И во всем, что он предпринимал на служение дому Божию и для соблюдения закона и заповедей, помышляя о Боге своем, он действовал от всего сердца своего и имел успех.
2CHR|32|1|После таких дел и верности, пришел Сеннахирим, царь Ассирийский, и вступил в Иудею, и осадил укрепленные города, и думал отторгнуть их себе.
2CHR|32|2|Когда Езекия увидел, что пришел Сеннахирим с намерением воевать против Иерусалима,
2CHR|32|3|тогда решил с князьями своими и с военными людьми своими засыпать источники воды, которые вне города, и те помогли ему.
2CHR|32|4|И собралось множество народа, и засыпали все источники и поток, протекавший по стране, говоря: да не найдут цари Ассирийские, придя [сюда], много воды.
2CHR|32|5|И ободрился он, и восстановил всю обрушившуюся стену, и поднял ее до башни, и извне [построил] другую стену, и укрепил Милло в городе Давидовом, и наготовил множество оружия и щитов.
2CHR|32|6|И поставил военачальников над народом, и собрал их к себе на площадь у городских ворот, и говорил к сердцу их, и сказал:
2CHR|32|7|будьте тверды и мужественны, не бойтесь и не страшитесь царя Ассирийского и всего множества, которое с ним, потому что с нами более, нежели с ним;
2CHR|32|8|с ним мышца плотская, а с нами Господь Бог наш, чтобы помогать нам и сражаться на бранях наших. И подкрепился народ словами Езекии, царя Иудейского.
2CHR|32|9|После сего послал Сеннахирим, царь Ассирийский, рабов своих в Иерусалим, – сам он [стоял] против Лахиса, и вся сила его с ним, – к Езекии, царю Иудейскому, и ко всем Иудеям, которые в Иерусалиме, сказать:
2CHR|32|10|так говорит Сеннахирим, царь Ассирийский: на что вы надеетесь и сидите в крепости в Иерусалиме?
2CHR|32|11|Не обольщает ли вас Езекия, чтобы предать вас смерти от голода и жажды, говоря: Господь Бог наш спасет нас от руки царя Ассирийского?
2CHR|32|12|Не этот ли Езекия разрушил высоты Его и жертвенники Его, и сказал Иудее и Иерусалиму: пред жертвенником единым поклоняйтесь и на нем совершайте курения?
2CHR|32|13|Разве вы не знаете, что сделал я и отцы мои со всеми народами земель? Могли ли боги народов земных спасти землю свою от руки моей?
2CHR|32|14|Кто из всех богов народов, истребленных отцами моими, мог спасти народ свой от руки моей? [Как же] возможет ваш Бог спасти вас от руки моей?
2CHR|32|15|И ныне пусть не обольщает вас Езекия и не отклоняет вас таким образом; не верьте ему: если не в силах был ни один бог ни одного народа и царства спасти народ свой от руки моей и от руки отцов моих, то и ваш Бог не спасет вас от руки моей.
2CHR|32|16|И еще [многое] говорили рабы его против Господа Бога и против Езекии, раба Его.
2CHR|32|17|И письма писал он, [в которых] поносил Господа Бога Израилева и говорил против Него такие слова: как боги народов земных не спасли народов своих от руки моей, так Бог Езекии не спасет народа Своего от руки моей.
2CHR|32|18|И кричали громким голосом на Иудейском языке к народу Иерусалимскому, который [был] на стене, чтоб устрашить его и напугать его, и взять город.
2CHR|32|19|И говорили о Боге Иерусалима, как о богах народов земли, – изделии рук человеческих.
2CHR|32|20|И помолился царь Езекия и Исаия, сын Амосов, пророк, и возопили к небу.
2CHR|32|21|И послал Господь Ангела, и он истребил всех храбрых и главноначальствующего и начальствующих в войске царя Ассирийского. И возвратился он со стыдом в землю свою; и когда пришел в дом бога своего, – исшедшие из чресл его поразили его там мечом.
2CHR|32|22|Так спас Господь Езекию и жителей Иерусалима от руки Сеннахирима, царя Ассирийского, и от руки всех и оберегал их отовсюду.
2CHR|32|23|Тогда многие приносили дары Господу в Иерусалим и дорогие вещи Езекии, царю Иудейскому. И он возвеличился после сего в глазах всех народов.
2CHR|32|24|В те дни заболел Езекия смертельно. И помолился Господу, и Он услышал его и дал ему знамение.
2CHR|32|25|Но не воздал Езекия за оказанные ему благодеяния, ибо возгордилось сердце его. И был на него гнев [Божий] и на Иудею, и на Иерусалим.
2CHR|32|26|Но как смирился Езекия в гордости сердца своего, – сам и жители Иерусалима, то не пришел на них гнев Господень во дни Езекии.
2CHR|32|27|И было у Езекии богатства и славы весьма много, и хранилище он сделал у себя для серебра и золота, и камней драгоценных, и для ароматов и щитов, и для всяких драгоценных сосудов;
2CHR|32|28|и кладовые для произведений [земли], для хлеба, вина и масла, и стойла для всякого рода скота, и дворы для стад.
2CHR|32|29|И города построил себе. И стад мелкого и крупного скота [было] [у него] множество, потому что дал ему Бог весьма большое имущество.
2CHR|32|30|Он же, Езекия, запер верхний проток вод Геона и провел их вниз к западной стороне города Давидова. И действовал успешно Езекия во всяком деле своем.
2CHR|32|31|Только при послах царей Вавилонских, которые присылали к нему спросить о знамении, бывшем на земле, оставил его Бог, чтоб испытать его и открыть все, что у него на сердце.
2CHR|32|32|Прочие деяния Езекии и добродетели его описаны в видении Исаии, сына Амосова, пророка, и в книге царей Иудейских и Израильских.
2CHR|32|33|И почил Езекия с отцами своими, и похоронили его над гробницами сыновей Давидовых, и почесть воздали ему по смерти его все Иудеи и жители Иерусалима. И воцарился Манассия, сын его, вместо него.
2CHR|33|1|Двенадцати лет [был] Манассия, когда воцарился, и пятьдесят пять лет царствовал в Иерусалиме,
2CHR|33|2|и делал он неугодное в очах Господних, подражая мерзостям народов, которых прогнал Господь от лица сынов Израилевых,
2CHR|33|3|и снова построил высоты, которые разрушил Езекия, отец его, и поставил жертвенники Ваалам, и устроил дубравы, и поклонялся всему воинству небесному, и служил ему,
2CHR|33|4|и соорудил жертвенники в доме Господнем, о котором сказал Господь: в Иерусалиме будет имя Мое вечно;
2CHR|33|5|и соорудил жертвенники всему воинству небесному на обоих дворах дома Господня.
2CHR|33|6|Он же проводил сыновей своих чрез огонь в долине сына Енномова, и гадал, и ворожил, и чародействовал, и учредил вызывателей мертвецов и волшебников; много делал он неугодного в очах Господа, к прогневлению Его.
2CHR|33|7|И поставил резного идола, которого сделал, в доме Божием, о котором говорил Бог Давиду и Соломону, сыну его: в доме сем и в Иерусалиме, который Я избрал из всех колен Израилевых, Я положу имя Мое навек;
2CHR|33|8|и не дам впредь выступить ноге Израиля из земли сей, которую Я укрепил за отцами их, если только они будут стараться исполнять все, что Я заповедал им, по всему закону и уставам и повелениям, [данным] рукою Моисея.
2CHR|33|9|Но Манассия довел Иудею и жителей Иерусалима до того, что они поступали хуже тех народов, которых истребил Господь от лица сынов Израилевых.
2CHR|33|10|И говорил Господь к Манассии и к народу его, но они не слушали.
2CHR|33|11|И привел Господь на них военачальников царя Ассирийского, и заковали они Манассию в кандалы и оковали его цепями, и отвели его в Вавилон.
2CHR|33|12|И в тесноте своей он стал умолять лице Господа Бога своего и глубоко смирился пред Богом отцов своих.
2CHR|33|13|И помолился Ему, и [Бог] преклонился к нему и услышал моление его, и возвратил его в Иерусалим на царство его. И узнал Манассия, что Господь есть Бог.
2CHR|33|14|И после того построил внешнюю стену города Давидова, на западной стороне Геона, по лощине и до входа в Рыбные ворота, и провел ее вокруг Офела и высоко поднял ее. И поставил военачальников по всем укрепленным городам в Иудее,
2CHR|33|15|и низверг чужеземных богов и идола из дома Господня, и все капища, которые соорудил на горе дома Господня и в Иерусалиме, и выбросил их за город.
2CHR|33|16|И восстановил жертвенник Господень и принес на нем жертвы мирные и хвалебные, и сказал Иудеям, чтобы они служили Господу Богу Израилеву.
2CHR|33|17|Но народ еще приносил жертвы на высотах, хотя и Господу Богу своему.
2CHR|33|18|Прочие дела Манассии, и молитва его к Богу своему, и слова прозорливцев, говоривших к нему именем Господа Бога Израилева, находятся в записях царей Израилевых.
2CHR|33|19|И молитва его, и то, что [Бог] преклонился к нему, и все грехи его и беззакония его, и места, на которых он построил высоты и поставил изображения Астарты и истуканов, прежде нежели смирился, описаны в записях Хозая.
2CHR|33|20|И почил Манассия с отцами своими, и похоронили его в доме его. И воцарился Амон, сын его, вместо него.
2CHR|33|21|Двадцати двух лет был Амон, когда воцарился, и два года царствовал в Иерусалиме.
2CHR|33|22|И делал неугодное в очах Господних так, как делал Манассия, отец его; и всем истуканам, которых сделал Манассия, отец его, приносил Амон жертвы и служил им.
2CHR|33|23|И не смирился пред лицем Господним, как смирился Манассия, отец его; напротив, Амон умножил [свои] грехи.
2CHR|33|24|И составили против него заговор слуги его, и умертвили его в доме его.
2CHR|33|25|Но народ земли перебил всех, бывших в заговоре против царя Амона, и воцарил народ земли Иосию, сына его, вместо него.
2CHR|34|1|Восемь лет было Иосии, когда он воцарился, и тридцать один год царствовал в Иерусалиме,
2CHR|34|2|и делал он угодное в очах Господних, и ходил путями Давида, отца своего, и не уклонялся ни направо, ни налево.
2CHR|34|3|В восьмой год царствования своего, будучи еще отроком, он начал прибегать к Богу Давида, отца своего, а в двенадцатый год начал очищать Иудею и Иерусалим от высот и [посвященных] дерев и от резных и литых кумиров.
2CHR|34|4|И разрушили пред лицем его жертвенники Ваалов и статуи, возвышавшиеся над ними; и [посвященные] дерева он срубил, и резные и литые кумиры изломал и разбил в прах, и рассыпал на гробах тех, которые приносили им жертвы,
2CHR|34|5|и кости жрецов сжег на жертвенниках их, и очистил Иудею и Иерусалим,
2CHR|34|6|и в городах Манассии, и Ефрема, и Симеона, [даже] до колена Неффалимова, и в опустошенных окрестностях их
2CHR|34|7|он разрушил жертвенники и [посвященные] дерева, и кумиры разбил в прах, и все статуи сокрушил по всей земле Израильской, и возвратился в Иерусалим.
2CHR|34|8|В восемнадцатый год царствования своего, по очищении земли и дома [Божия], он послал Шафана, сына Ацалии, и Маасею градоначальника, и Иоаха, сына Иоахазова, дееписателя, возобновить дом Господа Бога своего.
2CHR|34|9|И пришли они к Хелкии первосвященнику, и отдали серебро, принесенное в дом Божий, которое левиты, стоящие на страже у порога, собрали из рук Манассии и Ефрема и всех прочих Израильтян, и от всего Иуды и Вениамина, и от жителей Иерусалима,
2CHR|34|10|и отдали в руки производителям работ, приставленным к дому Господню, чтоб они раздавали его работникам, которые работали в доме Господнем, при исправлении и возобновлении дома.
2CHR|34|11|И они раздавали плотникам и строителям на покупку тесаных камней и дерев для связей и для покрытия зданий, которые разорили цари Иудейские.
2CHR|34|12|Люди сии действовали честно при работе, и для надзора над ними поставлены были Иахаф и Овадия, левиты из сыновей Мерариных, и Захария и Мешуллам из сыновей Каафовых, и все левиты, умеющие играть на музыкальных орудиях.
2CHR|34|13|Они же [были] приставниками над носильщиками и наблюдали над всеми работниками при каждой работе; из левитов же [были и] писцы, и надзиратели, и привратники.
2CHR|34|14|Когда вынимали они серебро, принесенное в дом Господень, тогда Хелкия священник нашел книгу закона Господня, [данную] рукою Моисея.
2CHR|34|15|И начал Хелкия, и сказал Шафану писцу: книгу закона нашел я в доме Господнем. И подал Хелкия ту книгу Шафану.
2CHR|34|16|И понес Шафан книгу к царю, и принес при этом царю известие: все, что поручено рабам твоим, они делают;
2CHR|34|17|и высыпали серебро, найденное в доме Господнем, и передали его в руки приставникам и в руки производителям работ.
2CHR|34|18|И [также] донес Шафан писец царю, говоря: книгу дал мне Хелкия священник. И читал ее Шафан перед царем.
2CHR|34|19|Когда услышал царь слова закона, то разодрал одежды свои.
2CHR|34|20|И дал царь повеление Хелкии и Ахикаму, сыну Шафанову, и Авдону, сыну Михея, и Шафану писцу, и Асаии, слуге царскому, говоря:
2CHR|34|21|пойдите, вопросите Господа за меня и за оставшихся у Израиля и за Иуду о словах сей найденной книги, потому что велик гнев Господа, который воспылал на нас за то, что не соблюдали отцы наши слова Господня, чтобы поступать по всему написанному в книге сей.
2CHR|34|22|И пошел Хелкия и те, которые от царя, к Олдане пророчице, жене Шаллума, сына Тавкегафа, сына Хасры, хранителя одежд, – а жила она во второй части Иерусалима, – и говорили с нею об этом.
2CHR|34|23|И она сказала им: так говорит Господь Бог Израилев: скажите тому человеку, который послал вас ко мне:
2CHR|34|24|так говорит Господь: вот Я наведу бедствие на место сие и на жителей его все проклятия, написанные в книге, которую читали пред лицем царя Иудейского,
2CHR|34|25|за то, что они оставили Меня и кадили богам другим, чтобы прогневлять Меня всеми делами рук своих. И гнев Мой возгорится над местом сим и не угаснет.
2CHR|34|26|А царю Иудейскому, пославшему вас вопросить Господа, так скажите: так говорит Господь Бог Израилев о словах, которые ты слышал:
2CHR|34|27|так как смягчилось сердце твое, и ты смирился пред Богом, услышав слова Его о месте сем и о жителях его, – и ты смирился предо Мною, и разодрал одежды свои, и плакал предо Мною, то и Я услышал [тебя], говорит Господь.
2CHR|34|28|Вот Я приложу тебя к отцам твоим, и положен будешь в гробницу твою в мире, и не увидят глаза твои всего того бедствия, которое Я наведу на место сие и на жителей его. И принесли царю ответ.
2CHR|34|29|И послал царь, и собрал всех старейшин Иудеи и Иерусалима,
2CHR|34|30|и пошел царь в дом Господень, и [с ним] все Иудеи и жители Иерусалима, и священники и левиты, и весь народ, от большого до малого; и он прочитал вслух их все слова книги завета, найденной в доме Господнем.
2CHR|34|31|И стал царь на месте своем, и заключил завет пред лицем Господа последовать Господу и соблюдать заповеди Его и откровения Его, и уставы Его, от всего сердца своего и от всей души своей, чтобы выполнить слова завета, написанные в книге сей.
2CHR|34|32|И велел царь подтвердить [это] всем находившимся в Иерусалиме и в земле Вениаминовой; и стали поступать жители Иерусалима по завету Бога, Бога отцов своих.
2CHR|34|33|И изверг Иосия все мерзости из всех земель, которые у сынов Израилевых, и повелел всем, находившимся в [земле] Израилевой служить Господу Богу своему. И во все дни [жизни] его они не отступали от Господа Бога отцов своих.
2CHR|35|1|И совершил Иосия в Иерусалиме пасху Господу, и закололи пасхального агнца в четырнадцатый [день] первого месяца.
2CHR|35|2|И поставил он священников на местах их, и ободрял их на служение в доме Господнем,
2CHR|35|3|и сказал левитам, наставникам всех Израильтян, посвященным Господу: поставьте ковчег святый в храме, который построил Соломон, сын Давидов, царь Израилев; нет вам нужды носить [его] на раменах; служите теперь Господу Богу нашему и народу Его Израилю;
2CHR|35|4|станьте по поколениям вашим, по чередам вашим, как предписано Давидом, царем Израилевым, и как предписано Соломоном, сыном его,
2CHR|35|5|и стойте во святилище, по распределениям поколений у братьев ваших, сынов народа, и по разделению поколений у левитов,
2CHR|35|6|и заколите пасхального агнца, и освятитесь, и приготовьте его для братьев ваших, поступая согласно со словом Господним чрез Моисея.
2CHR|35|7|И дал Иосия в дар сынам народа, всем, находившимся там, из мелкого скота агнцев и козлов молодых, все для жертвы пасхальной, числом тридцать тысяч и три тысячи волов. Это из имущества царя.
2CHR|35|8|И князья его по усердию давали в дар народу, священникам и левитам: Хелкия и Захария и Иехиил, начальствующие в доме Божием, дали священникам для жертвы пасхальной две тысячи шестьсот [овец, агнцев и козлов] и триста волов;
2CHR|35|9|и Хонания, и Шемаия, и Нафанаил, братья его, и Хашавия, и Иеиел, и Иозавад, начальники левитов, подарили левитам для жертвы пасхальной [овец] пять тысяч и пятьсот волов.
2CHR|35|10|Так устроено было служение. И стали священники на место свое и левиты по чередам своим, по повелению царскому;
2CHR|35|11|и закололи пасхального агнца. И кропили священники [кровью], принимая ее из рук левитов, а левиты снимали кожу;
2CHR|35|12|и распределили [назначенное] для всесожжения, чтобы раздать то по отделениям поколений у сынов народа, для принесения Господу, как написано в книге Моисеевой. То же [сделали] и с волами.
2CHR|35|13|И испекли пасхального агнца на огне, по уставу; и священные жертвы сварили в котлах, горшках и кастрюлях, и поспешно роздали всему народу,
2CHR|35|14|а после приготовили для себя и для священников, ибо священники, сыны Аароновы, [заняты были] приношением всесожжения и туков до ночи; потому–то и готовили левиты для себя и для священников, сынов Аароновых.
2CHR|35|15|И певцы, сыновья Асафовы, [оставались] на местах своих, по установлению Давида и Асафа, и Емана и Идифуна, прозорливца царского, и привратники у каждых ворот: не для чего [было] им отходить от служения своего, так как братья их левиты готовили для них.
2CHR|35|16|Так устроено было все служение Господу в тот день, чтобы совершить пасху и принести всесожжения на жертвеннике Господнем, по повелению царя Иосии.
2CHR|35|17|И совершали сыны Израилевы, находившиеся [там], пасху в то время и праздник опресноков в течение семи дней.
2CHR|35|18|И не была совершаема такая пасха у Израиля от дней Самуила пророка; и из всех царей Израилевых ни один не совершал такой пасхи, какую совершил Иосия, и священники, и левиты, и все Иудеи, и Израильтяне, [там] находившиеся, и жители Иерусалима.
2CHR|35|19|В восемнадцатый год царствования Иосии совершена сия пасха.
2CHR|35|20|После всего того, что сделал Иосия в доме [Божием], пошел Нехао, царь Египетский, на войну к Кархемису на Евфрате; и Иосия вышел навстречу ему.
2CHR|35|21|И послал к нему [Нехао] послов сказать: что мне и тебе, царь Иудейский? Не против тебя теперь [иду я,] но туда, где у меня война. И Бог повелел мне поспешать; не противься Богу, Который со мною, чтоб Он не погубил тебя.
2CHR|35|22|Но Иосия не отстранился от него, а приготовился, чтобы сразиться с ним, и не послушал слов Нехао от лица Божия и выступил на сражение на равнину Мегиддо.
2CHR|35|23|И выстрелили стрельцы в царя Иосию, и сказал царь слугам своим: уведите меня, потому что я тяжело ранен.
2CHR|35|24|И свели его слуги его с колесницы, и посадили его в другую повозку, которая [была] у него, и отвезли его в Иерусалим. И умер он, и похоронен в гробницах отцов своих. И вся Иудея и Иерусалим оплакали Иосию.
2CHR|35|25|Оплакал Иосию и Иеремия в песне плачевной; и говорили все певцы и певицы об Иосии в плачевных песнях своих, [известных] до сего дня, и передали их в употребление у Израиля; и вот они вписаны в [книгу] плачевных песней.
2CHR|35|26|Прочие деяния Иосии и добродетели его, согласные с предписанным в законе Господнем,
2CHR|35|27|и деяния его, первые и последние, описаны в книге царей Израильских и Иудейских.
2CHR|36|1|И взял народ земли Иоахаза, сына Иосиина, и воцарили его, вместо отца его, в Иерусалиме.
2CHR|36|2|Двадцати трех лет был Иоахаз, когда воцарился, и три месяца царствовал в Иерусалиме.
2CHR|36|3|И низложил его царь Египетский в Иерусалиме, наложил на землю пени сто талантов серебра и талант золота.
2CHR|36|4|И воцарил царь Египетский над Иудеею и Иерусалимом Елиакима, брата его, и переменил имя его на Иоакима, а Иоахаза, брата его, взял Нехао и отвел его в Египет.
2CHR|36|5|Двадцати пяти лет [был] Иоаким, когда воцарился, и одиннадцать лет царствовал в Иерусалиме. И делал он неугодное в очах Господа Бога своего.
2CHR|36|6|Против него вышел Навуходоносор, царь Вавилонский, и оковал его оковами, чтоб отвести его в Вавилон.
2CHR|36|7|И часть сосудов дома Господня перенес Навуходоносор в Вавилон и положил их в капище своем в Вавилоне.
2CHR|36|8|Прочие дела Иоакима и мерзости его, какие он делал и какие найдены в нем, описаны в книге царей Израильских и Иудейских. И воцарился Иехония, сын его, вместо него.
2CHR|36|9|Восемнадцати лет [был] Иехония, когда воцарился, и три месяца и десять дней царствовал в Иерусалиме, и делал он неугодное в очах Господних.
2CHR|36|10|По прошествии года послал царь Навуходоносор и велел взять его в Вавилон вместе с драгоценными сосудами дома Господня, и воцарил над Иудеею и Иерусалимом Седекию, брата его.
2CHR|36|11|Двадцати одного года [был] Седекия, когда воцарился, и одиннадцать лет царствовал в Иерусалиме,
2CHR|36|12|и делал он неугодное в очах Господа Бога своего. Он не смирился пред Иеремиею пророком, [пророчествовавшим] от уст Господних,
2CHR|36|13|и отложился от царя Навуходоносора, взявшего клятву с него [именем] Бога, – и сделал упругою шею свою и ожесточил сердце свое до того, что не обратился к Господу Богу Израилеву.
2CHR|36|14|Да и все начальствующие над священниками и над народом много грешили, подражая всем мерзостям язычников, и сквернили дом Господа, который Он освятил в Иерусалиме.
2CHR|36|15|И посылал к ним Господь Бог отцов их, посланников Своих от раннего утра, потому что Он жалел Свой народ и Свое жилище.
2CHR|36|16|Но они издевались над посланными от Бога и пренебрегали словами Его, и ругались над пророками Его, доколе не сошел гнев Господа на народ Его, так что не было [ему] спасения.
2CHR|36|17|И Он навел на них царя Халдейского, – и тот умертвил юношей их мечом в доме святыни их и не пощадил ни юноши, ни девицы, ни старца, ни седовласого: все предал [Бог] в руку его.
2CHR|36|18|И все сосуды дома Божия, большие и малые, и сокровища дома Господня, и сокровища царя и князей его, все принес он в Вавилон.
2CHR|36|19|И сожгли дом Божий, и разрушили стену Иерусалима, и все чертоги его сожгли огнем, и все драгоценности его истребили.
2CHR|36|20|И переселил он оставшихся от меча в Вавилон, и были они рабами его и сыновей его, до воцарения царя Персидского,
2CHR|36|21|доколе, во исполнение слова Господня, [сказанного] устами Иеремии, земля не отпраздновала суббот своих. Во все дни запустения она субботствовала до исполнения семидесяти лет.
2CHR|36|22|А в первый год Кира, царя Персидского, во исполнение слова Господня, [сказанного] устами Иеремии, возбудил Господь дух Кира, царя Персидского, и он велел объявить по всему царству своему, словесно и письменно, и сказать:
2CHR|36|23|так говорит Кир, царь Персидский: все царства земли дал мне Господь Бог небесный, и Он повелел мне построить Ему дом в Иерусалиме, что в Иудее. Кто есть из вас – из всего народа Его, [да будет] Господь Бог его с ним, и пусть он туда идет.
2CHR|36|24|МОЛИТВА МАНАССИИ, ЦАРЯ ИУДЕЙСКОГО, КОГДА ОН СОДЕРЖАЛСЯ В ПЛЕНУ В ВАВИЛОНЕ Господи Вседержителю, Боже отцев наших, Авраама и Исаака и Иакова, и семени их праведного [а], сотворивший небо и землю со всем благолепием их, связавший море словом повеления Твоего, заключивший бездну и запечатавший ее страшным и славным именем Твоим, которого все боятся, и трепещут от лица силы Твоея, потому что никто не может устоять пред великолепием славы Твоея, и нестерпим гнев [б] прещения Твоего на грешников [в]! Но безмерна и неисследима милость обетования Твоего [г], ибо Ты Господь вышний, благий, долготерпеливый и многомилостивый и кающийся о злобах человеческих. Ты, Господи, по множеству Твоей благости, обещал покаяние [д] и отпущение согрешившим Тебе, и множеством щедрот Твоих определил покаяние грешникам во спасение. Итак Ты, Господи, Боже праведных, не положил покаяния праведным [е] Аврааму и Исааку и Иакову, не согрешившим Тебе, но положил покаяние мне грешнику, потому что я согрешил паче числа песка морского. Многочисленны беззакония мои, Господи, многочисленны беззакония мои, и я недостоин взирать и смотреть на высоту небесную от множества неправд моих. Я согбен многими железными узами [з], так что не могу поднять головы моей, и нет мне отдохновения, потому что прогневал Тебя и сделал пред Тобою злое [и]: не исполнил воли Твоей, не сохранил повелений Твоих, поставил мерзости и умножил соблазны. И ныне преклоняю колени сердца моего, умоляя Тебя о благости [к]. Согрешил я, Господи, согрешил, и беззакония мои я знаю, но прошу, молясь Тебе: отпусти мне, Господи, отпусти мне, и не погуби меня с беззакониями моими и не оссуди меня в преисподнюю. Ибо Ты Бог, Бог кающихся, и на мне яви всю благость Твою, спасши меня недостойного по великой милости Твоей, и буду прославлять Тебя во все дни жизни моей [л], потому что Тебя славят все силы небесные, и Твоя слава во веки веков. Аминь.
