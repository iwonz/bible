LAM|1|1|唉！先前人口稠密的城市， 现在为何独坐！ 先前在列国中为大的， 现在竟如寡妇！ 先前在各省中为王后的， 现在竟成为服苦役的人！
LAM|1|2|她 夜间痛哭，泪流满颊， 在所有亲爱的人中，找不到一个安慰她的。 她的朋友都以诡诈待她， 成为她的仇敌。
LAM|1|3|犹大 被掳， 遭遇苦难，多服劳役。 她住在列国中，得不着安息； 追逼她的在狭窄之地追上她。
LAM|1|4|锡安 的道路因无人前来过节就哀伤， 她的城门荒凉， 祭司叹息， 少女悲伤； 她自己充满痛苦。
LAM|1|5|她的敌人作主， 她的仇敌亨通； 耶和华因她过犯多而使她受苦， 她的孩童在敌人面前去作俘虏。
LAM|1|6|锡安 的威荣全都失去。 她的领袖如找不着草场的鹿， 在追赶的人面前无力行走。
LAM|1|7|耶路撒冷 在困苦窘迫之时， 就追想古时一切的荣华。 她的百姓落在敌人手中，无人帮助； 敌人看见，就因她的毁灭嗤笑。
LAM|1|8|耶路撒冷 犯了大罪， 因此成为不洁净； 素来尊敬她的，见她裸露就都藐视她， 她自己也叹息退后。
LAM|1|9|她的污秽是在下摆上； 她未曾思想自己的结局， 她的败落令人惊诧， 无人安慰她。 “耶和华啊，求你看顾我的苦难， 因为仇敌强大。”
LAM|1|10|敌人伸手夺取她的一切贵重物品； 她眼见列国侵入她的圣所， 你曾吩咐他们不可进入你的集会。
LAM|1|11|她的百姓都叹息，寻求食物； 他们用贵重物品换取粮食，要救性命。 “耶和华啊，求你观看， 留意我多么卑微。”
LAM|1|12|所有过路的人哪，愿这事不要发生在你们身上 。 你们要留意观看， 有像这样临到我的痛苦没有？ 耶和华在他发烈怒的日子使我受苦。
LAM|1|13|他从高处降火进入我的骨头， 克制了我； 他张开网，绊我的脚， 使我退后， 又令我终日凄凉发昏。
LAM|1|14|他用手绑我罪过的轭， 卷绕着加在我颈项上； 他使我力量衰败。 主将我交在我不能抵挡的人手中。
LAM|1|15|主弃绝我们当中所有的勇士， 聚集会众攻击我， 要压碎我的年轻人。 主踹下少女 犹大 ， 在醡酒池中。
LAM|1|16|我因这些事哭泣， 眼泪汪汪； 因为那安慰我、使我重新得力的， 离我甚远。 我的儿女孤苦， 因为仇敌得胜了。
LAM|1|17|锡安 伸出双手，却无人安慰。 论到 雅各 ，耶和华已经出令， 使四围的人作他的仇敌； 耶路撒冷 在他们中间成为不洁净。
LAM|1|18|耶和华是公义的！ 我违背了他的命令。 万民哪，请听， 来看我的痛苦； 我的少女和壮丁都被掳去。
LAM|1|19|我招呼我所亲爱的， 他们却欺骗了我。 我的祭司和长老寻找食物，要救性命的时候， 就在城中断了气。
LAM|1|20|耶和华啊，求你观看， 因为我在急难中； 我的心肠烦乱， 我心在我里面翻转， 因我大大背逆。 在外，刀剑使人丧亡； 在家，犹如死亡。
LAM|1|21|有人听见我叹息 ， 却无人安慰我！ 我所有的仇敌听见我的患难就喜乐， 因这是你所做的。 你使你所宣告的日子来临， 愿他们像我一样。
LAM|1|22|愿他们的恶行都呈现在你面前； 你怎样因我一切的罪过待我， 求你也照样待他们； 因我叹息甚多，心中发昏。
LAM|2|1|唉！主竟发怒，使黑云遮蔽 锡安 ！ 他将 以色列 的华美从天扔在地上， 在他发怒的日子并不顾念自己的脚凳。
LAM|2|2|主吞灭 雅各 一切的住处，并不顾惜。 他发怒倾覆 犹大 的堡垒， 将它们夷为平地， 凌辱这国与她的领袖。
LAM|2|3|他发烈怒，砍断 以色列 一切的角， 在仇敌面前收回右手。 他将 雅各 烧毁，如火焰四围吞灭。
LAM|2|4|他张弓好像仇敌， 他站立举起右手， 如同敌人杀戮我们眼目所喜爱的。 他在 锡安 的帐棚 倾倒愤怒，如火一般。
LAM|2|5|主如仇敌吞灭 以色列 ， 吞灭它一切的宫殿， 毁坏境内的堡垒； 在 犹大 加添悲伤和哭号。
LAM|2|6|他摧毁自己的帐幕如摧毁园子， 毁坏自己的会幕。 耶和华使节庆和安息日在 锡安 尽被遗忘， 又在极其愤怒中厌弃君王与祭司。
LAM|2|7|耶和华撇弃自己的祭坛， 憎恶自己的圣所， 把宫殿的墙交给仇敌。 他们在耶和华的殿中喧嚷， 如在节庆之日一样。
LAM|2|8|耶和华定意拆毁 锡安 的城墙； 他拉了准绳， 不将手收回，定要毁灭。 他使城郭和城墙都悲哀， 一同衰败。
LAM|2|9|锡安 的门陷入地里， 主毁坏，折断她的门闩。 她的君王和官长都置身列国中，没有律法； 她的先知也不再从耶和华领受异象。
LAM|2|10|锡安 的长老坐在地上，默默无声； 他们扬起尘土落在头上，腰束麻布； 耶路撒冷 的少女垂头至地。
LAM|2|11|我的眼睛流泪，以致失明； 我的心肠烦乱，肝胆落地， 都因我的百姓 遭毁灭， 又因孩童和吃奶的在城内的广场上昏厥。
LAM|2|12|他们如受伤的人在城内广场上昏厥， 在母亲的怀里将要丧命时， 就对母亲说：“饼和酒在哪里呢？”
LAM|2|13|耶路撒冷 啊，我可用什么向你证明 呢？ 我可用什么与你相比呢？ 少女 锡安 哪，我拿什么和你比较，好安慰你呢？ 因你的裂伤大如海； 谁能医治你呢？
LAM|2|14|你的先知为你看见虚假和粉饰的异象， 并未揭露你的罪孽， 使你被掳的归回； 却传给你虚假与误导人的默示。
LAM|2|15|凡过路的都向你拍掌。 他们向 耶路撒冷 嗤笑，摇头： “这就是人称为全美的、 称为全地所喜悦的城吗？”
LAM|2|16|你所有的仇敌 张口来攻击你； 他们嗤笑，切齿，说： “我们把她吞灭了， 这是我们所盼望的日子！ 我们终于等到了，亲眼看见了！”
LAM|2|17|耶和华成就了他所定的， 应验了他古时所命定的。 他倾覆，并不顾惜， 他使仇敌向你夸耀， 使你敌人的角高举。
LAM|2|18|他们的心哀求主。 锡安 的城墙啊， 愿你日夜泪流如河，不让自己休息， 你眼中的瞳人也不歇息。
LAM|2|19|夜间每逢时辰开始，要起来呼喊， 在主面前倾心吐意如水。 你的孩童在街头上挨饿昏厥， 你要为他们的性命向主举手。
LAM|2|20|耶和华啊，求你观看， 留意你向谁这样行。 妇人岂可吃自己所生、所抚育的婴孩吗？ 祭司和先知岂可在主的圣所中被杀吗？
LAM|2|21|年轻人和老年人躺卧在街上， 我的少女和壮丁都倒在刀下。 你在发怒的日子杀了他们， 你杀戮，并不顾惜。
LAM|2|22|你从四围招聚使我惊吓的人， 像在节庆的日子一样。 耶和华发怒的日子， 无人逃脱，无人生还。 我所抚育养大的， 仇敌都杀尽了。
LAM|3|1|因耶和华愤怒的杖， 我是遭遇困苦的人。
LAM|3|2|他驱赶我走入黑暗， 没有光明。
LAM|3|3|他反手攻击我， 终日不停。
LAM|3|4|他使我皮肉枯干， 折断我的骨头。
LAM|3|5|他筑垒攻击我， 以苦楚和艰难围困我；
LAM|3|6|使我住在幽暗之处， 像死了许久的人一样。
LAM|3|7|他围住我，使我无法脱身； 他使我的铜链沉重。
LAM|3|8|尽管我哀号求救， 他仍拦阻我的祷告。
LAM|3|9|他用凿过的石头挡住我的道路， 使我的路径弯曲。
LAM|3|10|他向我如埋伏的熊， 如在隐密处的狮子。
LAM|3|11|他使我转离正路， 把我撕碎 ，使我凄凉。
LAM|3|12|他拉弓，命我站立， 作为箭靶；
LAM|3|13|把箭袋中的箭 射入我的肺腑。
LAM|3|14|我成了全体百姓的笑柄， 成了他们终日的歌曲。
LAM|3|15|他使我受尽苦楚， 饱食茵蔯；
LAM|3|16|用沙石磨断我的牙， 以灰尘覆盖我。
LAM|3|17|你使我远离平安， 我忘了何为福乐。
LAM|3|18|于是我说：“我的力量衰败， 在耶和华那里我毫无指望！”
LAM|3|19|求你记得我的困苦和流离， 它如茵蔯和苦胆一般；
LAM|3|20|我心想念这些， 就在我里面忧闷 。
LAM|3|21|但我的心回转过来， 因此就有指望；
LAM|3|22|因耶和华的慈爱，我们不致灭绝 ， 因他的怜悯永不断绝，
LAM|3|23|每早晨，这些都是新的； 你的信实极其广大！
LAM|3|24|我心里说：“耶和华是我的福分， 因此，我要仰望他。”
LAM|3|25|凡等候耶和华，心里寻求他的， 耶和华必施恩给他。
LAM|3|26|人仰望耶和华， 安静等候他的救恩， 这是好的。
LAM|3|27|人在年轻时负轭， 这是好的。
LAM|3|28|他当安静独坐， 因为这是耶和华加在他身上的。
LAM|3|29|让他脸伏于地 吧！ 或者还会有指望。
LAM|3|30|让人打他耳光， 使他饱受凌辱吧！
LAM|3|31|主必不永远撇弃，
LAM|3|32|他虽使人忧愁， 还要照他丰盛的慈爱施怜悯；
LAM|3|33|他并不存心要人受苦， 令世人忧愁。
LAM|3|34|把世上所有的囚犯 踹在脚下，
LAM|3|35|在至高者面前 扭曲人的公正，
LAM|3|36|在人的诉讼上 颠倒是非， 这都是主看不中的。
LAM|3|37|若非主发命令， 谁能说了就成呢？
LAM|3|38|是祸，是福， 不都出于至高者的口吗？
LAM|3|39|人都有自己的罪， 活人有什么好发怨言的呢？
LAM|3|40|让我们省察，检讨自己的行为， 归向耶和华吧！
LAM|3|41|让我们献上我们的心， 向天上的上帝举手！
LAM|3|42|我们犯罪悖逆， 你并未赦免。
LAM|3|43|你浑身是怒气，追赶我们； 你施行杀戮，并不顾惜。
LAM|3|44|你以密云围着自己， 祷告不能穿透。
LAM|3|45|你使我们在万民中 成为污物和垃圾。
LAM|3|46|我们所有的仇敌 张口来攻击我们；
LAM|3|47|惊吓和陷阱临到我们， 残害和毁灭也临到我们。
LAM|3|48|因我百姓 遭毁灭， 我的眼睛泪流成河。
LAM|3|49|我的眼睛流泪不停， 流泪不止，
LAM|3|50|直等到耶和华垂顾， 从天上观看。
LAM|3|51|为我城中的百姓 ， 我眼所见的使我心痛。
LAM|3|52|无故与我为敌的追逼我， 像追捕雀鸟一样。
LAM|3|53|他们要在坑中了结我的性命， 丢石头在我身上。
LAM|3|54|众水淹没我的头， 我说：“我没命了！”
LAM|3|55|耶和华啊， 在极深的地府里，我求告你的名。
LAM|3|56|我的声音你听见了， 求你不要掩耳不听 我的呼声，我的求救。
LAM|3|57|我求告你的时候， 你临近我，说：“不要惧怕！”
LAM|3|58|主啊，你为我伸冤， 你救赎了我的命。
LAM|3|59|耶和华啊，你已看见我的委屈， 求你为我主持正义。
LAM|3|60|他们要报复，谋害我， 你都看见了。
LAM|3|61|耶和华啊，你听见他们的辱骂， 他们害我的一切计谋，
LAM|3|62|那些起来攻击我的人嘴唇所说的话 和他们终日攻击我的计谋。
LAM|3|63|求你留意！ 他们无论坐下或起来， 我都是他们的笑柄。
LAM|3|64|耶和华啊，求你照他们手所做的 向他们施行报应。
LAM|3|65|求你使他们心里刚硬， 使你的诅咒临到他们。
LAM|3|66|求你发怒追赶他们， 从耶和华的地上 除灭他们。
LAM|4|1|唉！黄金竟然无光！ 纯金竟然变色！ 圣所的石头散落在街上。
LAM|4|2|锡安 宝贝的孩子虽然好比精金， 现在竟当作陶匠手所做的瓦瓶！
LAM|4|3|野狗尚且哺乳其子， 我百姓 的妇人反倒残忍， 如旷野的鸵鸟一般；
LAM|4|4|吃奶孩子的舌头因干渴贴住上膛， 孩童求饼，却无人擘给他们。
LAM|4|5|素来吃美好食物的， 如今遭遗弃在街上； 素来穿着朱红衣裳长大的， 如今却拥抱粪堆。
LAM|4|6|我百姓的罪孽比 所多玛 的罪还大； 所多玛 虽无人伸手攻击， 转眼之间就被倾覆。
LAM|4|7|锡安 的拿细耳人 比雪纯净， 比奶更白； 他们的身体比宝石更红， 身躯之美如蓝宝石一般。
LAM|4|8|但如今他们的面貌比煤炭更黑， 在街上无人认识； 他们的皮肤紧贴骨头， 枯干形同槁木。
LAM|4|9|被刀剑刺杀的 胜过因饥饿而死 的； 饥饿者由于缺乏田里的出产 就消瘦而亡 。
LAM|4|10|当我百姓遭毁灭的时候， 慈心的妇人亲手烹煮自己的儿女为食物。
LAM|4|11|耶和华发尽他的愤怒， 倾倒他的烈怒， 用火焚烧 锡安 ， 烧毁 锡安 的根基。
LAM|4|12|地上的君王和世上的居民都不信 敌人和仇敌竟能进入 耶路撒冷 的城门。
LAM|4|13|这都因她先知的罪恶和祭司的罪孽， 他们在城中流了义人的血。
LAM|4|14|他们如盲人在街上徘徊， 又被血玷污， 以致人不敢摸他们的衣服。
LAM|4|15|人向他们喊着： “你这不洁净的，走开！ 走开！走开！不要摸我！” 他们逃走流浪的时候， 列国中有人说： “他们不可再寄居此地。”
LAM|4|16|耶和华亲自赶散他们， 不再眷顾他们； 不看重祭司，也不厚待长老。
LAM|4|17|我们的眼目徒然仰望帮助，以致失明， 我们从了望台所守望的，竟是一个不能救人的国！
LAM|4|18|仇敌追逐我们的脚踪， 使我们不敢在自己的街上行走。 我们的结局临近， 日子已满， 我们的结局已经来到。
LAM|4|19|追赶我们的比空中的鹰更快； 他们在山上追逼我们， 在旷野埋伏，等候我们。
LAM|4|20|耶和华的受膏者是我们鼻中的气， 被抓到他们的坑里， 论到他，我们曾说： “我们必在他荫下， 在列国中存活。”
LAM|4|21|住 乌斯 地的 以东 啊，尽管欢喜快乐， 苦杯必传到你那里； 你要喝醉，裸露自己。
LAM|4|22|锡安 哪，你罪孽的惩罚已经结束， 耶和华必不再使你被掳去。 以东 啊，耶和华必惩罚你的罪孽， 揭露你的罪恶。
LAM|5|1|耶和华啊，求你顾念我们所遭遇的， 留意看我们所受的凌辱。
LAM|5|2|我们的产业归陌生人， 我们的房屋归外邦人。
LAM|5|3|我们是无父的孤儿， 我们的母亲如同寡妇。
LAM|5|4|我们出银钱才得水喝， 我们的柴也是用钱买来的。
LAM|5|5|我们被追赶，迫及颈项， 疲乏却不得歇息。
LAM|5|6|我们束手投降 埃及 和 亚述 ， 为要得粮吃饱。
LAM|5|7|我们的祖先犯罪，而今他们不在了， 我们却担当他们的罪孽。
LAM|5|8|奴仆辖制我们， 无人救我们脱离他们的手。
LAM|5|9|因旷野有刀剑， 我们冒生命的危险才能得粮食。
LAM|5|10|因饥荒的干热， 我们的皮肤热如火炉。
LAM|5|11|他们在 锡安 玷污妇人， 在 犹大 城镇污辱少女。
LAM|5|12|他们吊起领袖的手， 使长老脸上无光。
LAM|5|13|年轻人扛磨石， 孩童背木柴而跌倒。
LAM|5|14|城门口不再有老年人， 年轻人也不再奏乐。
LAM|5|15|我们心中的快乐止息， 跳舞转为悲哀。
LAM|5|16|冠冕从我们的头上掉落； 我们有祸了，因为犯了罪。
LAM|5|17|因这些事我们心里发昏， 眼睛昏花。
LAM|5|18|锡安山 荒凉， 狐狸行在其上。
LAM|5|19|耶和华啊，你治理直到永远， 你的宝座万代长存。
LAM|5|20|你为何全然忘记我们？ 为何长久离弃我们？
LAM|5|21|耶和华啊，求你使我们回转归向你， 我们就得以回转。 求你更新我们的年日，像古时一样，
LAM|5|22|难道你全然弃绝了我们， 向我们大发烈怒？
