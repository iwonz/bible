2PET|1|1|Simon Peter, a servant and an apostle of Jesus Christ, to them that have obtained like precious faith with us through the righteousness of God and our Saviour Jesus Christ:
2PET|1|2|Grace and peace be multiplied unto you through the knowledge of God, and of Jesus our Lord,
2PET|1|3|According as his divine power hath given unto us all things that pertain unto life and godliness, through the knowledge of him that hath called us to glory and virtue:
2PET|1|4|Whereby are given unto us exceeding great and precious promises: that by these ye might be partakers of the divine nature, having escaped the corruption that is in the world through lust.
2PET|1|5|And beside this, giving all diligence, add to your faith virtue; and to virtue knowledge;
2PET|1|6|And to knowledge temperance; and to temperance patience; and to patience godliness;
2PET|1|7|And to godliness brotherly kindness; and to brotherly kindness charity.
2PET|1|8|For if these things be in you, and abound, they make you that ye shall neither be barren nor unfruitful in the knowledge of our Lord Jesus Christ.
2PET|1|9|But he that lacketh these things is blind, and cannot see afar off, and hath forgotten that he was purged from his old sins.
2PET|1|10|Wherefore the rather, brethren, give diligence to make your calling and election sure: for if ye do these things, ye shall never fall:
2PET|1|11|For so an entrance shall be ministered unto you abundantly into the everlasting kingdom of our Lord and Saviour Jesus Christ.
2PET|1|12|Wherefore I will not be negligent to put you always in remembrance of these things, though ye know them, and be established in the present truth.
2PET|1|13|Yea, I think it meet, as long as I am in this tabernacle, to stir you up by putting you in remembrance;
2PET|1|14|Knowing that shortly I must put off this my tabernacle, even as our Lord Jesus Christ hath shewed me.
2PET|1|15|Moreover I will endeavour that ye may be able after my decease to have these things always in remembrance.
2PET|1|16|For we have not followed cunningly devised fables, when we made known unto you the power and coming of our Lord Jesus Christ, but were eyewitnesses of his majesty.
2PET|1|17|For he received from God the Father honour and glory, when there came such a voice to him from the excellent glory, This is my beloved Son, in whom I am well pleased.
2PET|1|18|And this voice which came from heaven we heard, when we were with him in the holy mount.
2PET|1|19|We have also a more sure word of prophecy; whereunto ye do well that ye take heed, as unto a light that shineth in a dark place, until the day dawn, and the day star arise in your hearts:
2PET|1|20|Knowing this first, that no prophecy of the scripture is of any private interpretation.
2PET|1|21|For the prophecy came not in old time by the will of man: but holy men of God spake as they were moved by the Holy Ghost.
2PET|2|1|But there were false prophets also among the people, even as there shall be false teachers among you, who privily shall bring in damnable heresies, even denying the Lord that bought them, and bring upon themselves swift destruction.
2PET|2|2|And many shall follow their pernicious ways; by reason of whom the way of truth shall be evil spoken of.
2PET|2|3|And through covetousness shall they with feigned words make merchandise of you: whose judgment now of a long time lingereth not, and their damnation slumbereth not.
2PET|2|4|For if God spared not the angels that sinned, but cast them down to hell, and delivered them into chains of darkness, to be reserved unto judgment;
2PET|2|5|And spared not the old world, but saved Noah the eighth person, a preacher of righteousness, bringing in the flood upon the world of the ungodly;
2PET|2|6|And turning the cities of Sodom and Gomorrha into ashes condemned them with an overthrow, making them an ensample unto those that after should live ungodly;
2PET|2|7|And delivered just Lot, vexed with the filthy conversation of the wicked:
2PET|2|8|(For that righteous man dwelling among them, in seeing and hearing, vexed his righteous soul from day to day with their unlawful deeds;)
2PET|2|9|The Lord knoweth how to deliver the godly out of temptations, and to reserve the unjust unto the day of judgment to be punished:
2PET|2|10|But chiefly them that walk after the flesh in the lust of uncleanness, and despise government. Presumptuous are they, selfwilled, they are not afraid to speak evil of dignities.
2PET|2|11|Whereas angels, which are greater in power and might, bring not railing accusation against them before the Lord.
2PET|2|12|But these, as natural brute beasts, made to be taken and destroyed, speak evil of the things that they understand not; and shall utterly perish in their own corruption;
2PET|2|13|And shall receive the reward of unrighteousness, as they that count it pleasure to riot in the day time. Spots they are and blemishes, sporting themselves with their own deceivings while they feast with you;
2PET|2|14|Having eyes full of adultery, and that cannot cease from sin; beguiling unstable souls: an heart they have exercised with covetous practices; cursed children:
2PET|2|15|Which have forsaken the right way, and are gone astray, following the way of Balaam the son of Bosor, who loved the wages of unrighteousness;
2PET|2|16|But was rebuked for his iniquity: the dumb ass speaking with man's voice forbad the madness of the prophet.
2PET|2|17|These are wells without water, clouds that are carried with a tempest; to whom the mist of darkness is reserved for ever.
2PET|2|18|For when they speak great swelling words of vanity, they allure through the lusts of the flesh, through much wantonness, those that were clean escaped from them who live in error.
2PET|2|19|While they promise them liberty, they themselves are the servants of corruption: for of whom a man is overcome, of the same is he brought in bondage.
2PET|2|20|For if after they have escaped the pollutions of the world through the knowledge of the Lord and Saviour Jesus Christ, they are again entangled therein, and overcome, the latter end is worse with them than the beginning.
2PET|2|21|For it had been better for them not to have known the way of righteousness, than, after they have known it, to turn from the holy commandment delivered unto them.
2PET|2|22|But it is happened unto them according to the true proverb, The dog is turned to his own vomit again; and the sow that was washed to her wallowing in the mire.
2PET|3|1|This second epistle, beloved, I now write unto you; in both which I stir up your pure minds by way of remembrance:
2PET|3|2|That ye may be mindful of the words which were spoken before by the holy prophets, and of the commandment of us the apostles of the Lord and Saviour:
2PET|3|3|Knowing this first, that there shall come in the last days scoffers, walking after their own lusts,
2PET|3|4|And saying, Where is the promise of his coming? for since the fathers fell asleep, all things continue as they were from the beginning of the creation.
2PET|3|5|For this they willingly are ignorant of, that by the word of God the heavens were of old, and the earth standing out of the water and in the water:
2PET|3|6|Whereby the world that then was, being overflowed with water, perished:
2PET|3|7|But the heavens and the earth, which are now, by the same word are kept in store, reserved unto fire against the day of judgment and perdition of ungodly men.
2PET|3|8|But, beloved, be not ignorant of this one thing, that one day is with the Lord as a thousand years, and a thousand years as one day.
2PET|3|9|The Lord is not slack concerning his promise, as some men count slackness; but is longsuffering to us-ward, not willing that any should perish, but that all should come to repentance.
2PET|3|10|But the day of the Lord will come as a thief in the night; in the which the heavens shall pass away with a great noise, and the elements shall melt with fervent heat, the earth also and the works that are therein shall be burned up.
2PET|3|11|Seeing then that all these things shall be dissolved, what manner of persons ought ye to be in all holy conversation and godliness,
2PET|3|12|Looking for and hasting unto the coming of the day of God, wherein the heavens being on fire shall be dissolved, and the elements shall melt with fervent heat?
2PET|3|13|Nevertheless we, according to his promise, look for new heavens and a new earth, wherein dwelleth righteousness.
2PET|3|14|Wherefore, beloved, seeing that ye look for such things, be diligent that ye may be found of him in peace, without spot, and blameless.
2PET|3|15|And account that the longsuffering of our Lord is salvation; even as our beloved brother Paul also according to the wisdom given unto him hath written unto you;
2PET|3|16|As also in all his epistles, speaking in them of these things; in which are some things hard to be understood, which they that are unlearned and unstable wrest, as they do also the other scriptures, unto their own destruction.
2PET|3|17|Ye therefore, beloved, seeing ye know these things before, beware lest ye also, being led away with the error of the wicked, fall from your own stedfastness.
2PET|3|18|But grow in grace, and in the knowledge of our Lord and Saviour Jesus Christ. To him be glory both now and for ever. Amen.
