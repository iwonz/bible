JONAH|1|1|耶和華的話臨到 亞米太 的兒子 約拿 ，說：
JONAH|1|2|「起來，到 尼尼微 大城去，向其中的居民宣告，因為他們的惡已達到我面前。」
JONAH|1|3|約拿 卻起身，逃往 他施 去躲避耶和華。他下到 約帕 ，遇見一條船要往 他施 去。 約拿 付了船費，就上船，與船上的人同往 他施 ，為要躲避耶和華。
JONAH|1|4|耶和華在海上颳起大風，海就狂風大作，船幾乎破裂。
JONAH|1|5|水手都懼怕，各人哀求自己的神明。他們把船上的貨物拋進海裏，為要減輕載重。 約拿 卻下到艙底，躺臥沉睡。
JONAH|1|6|船長到他那裏，對他說：「你怎麼還在沉睡呢？起來，求告你的神明，或者神明顧念我們，使我們不致滅亡。」
JONAH|1|7|船上的人彼此說：「來吧，我們來抽籤，看看這災難臨到我們是因誰的緣故。」於是他們就抽籤，抽出 約拿 來。
JONAH|1|8|他們對 約拿 說：「請你告訴我們，這災難臨到我們是因誰的緣故呢？你做甚麼行業？你從哪裏來？你是哪一國的人？屬哪一族？」
JONAH|1|9|他說：「我是 希伯來 人，我敬畏耶和華，天上的上帝，他創造了滄海和陸地。」
JONAH|1|10|那些人就大大懼怕，對他說：「你做的是甚麼事呢？」原來他們已經知道他在躲避耶和華，因為他告訴了他們。
JONAH|1|11|海浪越來越洶湧，他們就問他說：「我們當向你做甚麼，才能使海浪平靜呢？」
JONAH|1|12|他對他們說：「你們把我抬起來，拋進海裏，海就會平靜了；我知道你們遭遇這大風浪是因我的緣故。」
JONAH|1|13|然而那些人竭力划槳，想要把船靠回陸地，卻是不能；因風浪愈來愈大，撲向他們。
JONAH|1|14|於是他們求告耶和華說：「耶和華啊，求求你不要因這人的性命使我們滅亡，不要使流無辜人血的罪歸給我們；因為你－耶和華隨自己的旨意行事。」
JONAH|1|15|他們把 約拿 抬起來，拋進海裏，海的狂浪就平息了。
JONAH|1|16|那些人就大大懼怕耶和華，向耶和華獻祭許願。
JONAH|1|17|耶和華安排一條大魚吞下 約拿 ， 約拿 在魚腹中三日三夜。
JONAH|2|1|約拿 在魚腹中向耶和華－他的上帝禱告，
JONAH|2|2|說： 「我在患難中求告耶和華， 他就應允我； 我從陰間的深處呼求， 你就俯聽我的聲音。
JONAH|2|3|你將我投下深淵， 直到海心； 大水環繞我， 你的波浪洪濤漫過我身。
JONAH|2|4|我說：『我從你眼前被驅逐， 然而我仍要仰望你的聖殿。』
JONAH|2|5|眾水環繞我，幾乎淹沒我； 深淵圍住我； 海草纏繞我的頭。
JONAH|2|6|我下沉到山的根基， 地的門閂將我永遠關住。 耶和華－我的上帝啊， 你卻將我的性命從地府裏救出來。
JONAH|2|7|我心靈發昏時， 就想起耶和華。 我的禱告進入你的聖殿， 達到你面前。
JONAH|2|8|那信奉虛無神明 的人， 丟棄自己的慈愛；
JONAH|2|9|但我要以感謝的聲音向你獻祭。 我所許的願，我必償還。 救恩出於耶和華。」
JONAH|2|10|耶和華吩咐那魚，魚就把 約拿 吐在陸地上。
JONAH|3|1|耶和華的話第二次臨到 約拿 ，說：
JONAH|3|2|「起來，到 尼尼微 大城去，把我告訴你的信息向其中的居民宣告。」
JONAH|3|3|約拿 就照耶和華的話起來，到 尼尼微 去。 尼尼微 是一座極大的城，約有三天的路程。
JONAH|3|4|約拿 進城，走了一天，宣告說：「再過四十天， 尼尼微 要傾覆了！」
JONAH|3|5|尼尼微 人就信服上帝，宣告禁食，從最大的到最小的都穿上麻衣。
JONAH|3|6|這消息傳到 尼尼微 王那裏，他就從寶座起來，脫下朝服，披上麻布，坐在灰中。
JONAH|3|7|他叫人通告 尼尼微 全城，說：「王和大臣有令，人、畜、牛、羊都不可嘗任何東西，不可吃，也不可喝水。
JONAH|3|8|人與牲畜都要披上麻布，切切求告上帝。各人要回轉離開惡道，離棄自己掌中的殘暴。
JONAH|3|9|誰知道上帝也許會回心轉意，不發烈怒，使我們不致滅亡。」
JONAH|3|10|上帝察看他們的行為，見他們離開惡道，上帝就改變心意，原先所說要降與他們的災難，他不降了。
JONAH|4|1|這事令 約拿 大大不悅，甚至發怒。
JONAH|4|2|他就向耶和華禱告，說：「耶和華啊，這不就是我仍在本國的時候所說的嗎？我知道你是有恩惠，有憐憫的上帝，不輕易發怒，有豐盛的慈愛，並且會改變心意，不降那災難。我就是因為這樣，才急速逃往 他施 去的呀！
JONAH|4|3|耶和華啊，現在求你取走我的性命吧！因為我死了比活著更好。」
JONAH|4|4|耶和華說：「你這樣發怒，對嗎？」
JONAH|4|5|約拿 出城，坐在城的東邊，在那裏為自己搭了一座棚。他坐在棚子的蔭下，要看看城裏會發生甚麼事。
JONAH|4|6|耶和華上帝安排了一棵蓖麻，使它生長高過 約拿 ，影子遮蓋他的頭，使他免受苦難； 約拿 因這棵蓖麻大大歡喜。
JONAH|4|7|次日黎明，上帝卻安排一條蟲來咬這蓖麻，以致枯乾。
JONAH|4|8|太陽出來的時候，上帝安排炎熱的東風，太陽曝曬 約拿 的頭，使他發昏，他就為自己求死，說：「我死了比活著更好！」
JONAH|4|9|上帝對 約拿 說：「你因這棵蓖麻這樣發怒，對嗎？」他說：「我發怒以至於死，都是對的！」
JONAH|4|10|耶和華說：「這棵蓖麻你沒有為它操勞，也不是你使它長大的；它一夜生長，一夜枯死，你尚且愛惜；
JONAH|4|11|何況這 尼尼微 大城，其中不能分辨左右手的就有十二萬多人，還有許多牲畜，我豈能不愛惜呢？」
