1CHR|1|1|亞當 ， 塞特 ， 以挪士 ，
1CHR|1|2|該南 ， 瑪勒列 ， 雅列 ，
1CHR|1|3|以諾 ， 瑪土撒拉 ， 拉麥 ，
1CHR|1|4|挪亞 ， 閃 ， 含 ， 雅弗 。
1CHR|1|5|雅弗 的兒子是 歌篾 、 瑪各 、 瑪代 、 雅完 、 土巴 、 米設 和 提拉 。
1CHR|1|6|歌篾 的兒子是 亞實基拿 、 低法 和 陀迦瑪 。
1CHR|1|7|雅完 的兒子是 以利沙 、 他施 、 基提 和 羅單 人 。
1CHR|1|8|含 的兒子是 古實 、 麥西 、 弗 和 迦南 。
1CHR|1|9|古實 的兒子是 西巴 、 哈腓拉 、 撒弗他 、 拉瑪 和 撒弗提迦 。 拉瑪 的兒子是 示巴 和 底但 。
1CHR|1|10|古實 又生 寧錄 ，他是地上第一個勇士。
1CHR|1|11|麥西 生 路低 人、 亞拿米 人、 利哈比 人、 拿弗土希 人、
1CHR|1|12|帕斯魯細 人、 迦斯路希 人和 迦斐託 人； 非利士 人是從 迦斐託 人 出來的。
1CHR|1|13|迦南 生了長子 西頓 ，又生 赫
1CHR|1|14|和 耶布斯 人、 亞摩利 人、 革迦撒 人、
1CHR|1|15|希未 人、 亞基 人、 西尼 人、
1CHR|1|16|亞瓦底 人、 洗瑪利 人和 哈馬 人。
1CHR|1|17|閃 的兒子是 以攔 、 亞述 、 亞法撒 、 路德 、 亞蘭 、 烏斯 、 戶勒 、 基帖 和 米設 。
1CHR|1|18|亞法撒 生 沙拉 ； 沙拉 生 希伯 。
1CHR|1|19|希伯 生了兩個兒子：一個名叫 法勒 ，因為那時人分地居住； 法勒 的兄弟名叫 約坍 。
1CHR|1|20|約坍 生 亞摩答 、 沙列 、 哈薩瑪非 、 耶拉 、
1CHR|1|21|哈多蘭 、 烏薩 、 德拉 、
1CHR|1|22|以巴錄 、 亞比瑪利 、 示巴 、
1CHR|1|23|阿斐 、 哈腓拉 和 約巴 。這些都是 約坍 的兒子。
1CHR|1|24|閃 ， 亞法撒 ， 沙拉 ，
1CHR|1|25|希伯 ， 法勒 ， 拉吳 ，
1CHR|1|26|西鹿 ， 拿鶴 ， 他拉 ，
1CHR|1|27|亞伯蘭 ， 亞伯蘭 就是 亞伯拉罕 。
1CHR|1|28|亞伯拉罕 的兒子是 以撒 和 以實瑪利 。
1CHR|1|29|以實瑪利 的後代如下： 以實瑪利 的長子是 尼拜約 ，又有 基達 、 亞德別 、 米比衫 、
1CHR|1|30|米施瑪 、 度瑪 、 瑪撒 、 哈大 、 提瑪 、
1CHR|1|31|伊突 、 拿非施 和 基底瑪 。這些都是 以實瑪利 的兒子。
1CHR|1|32|亞伯拉罕 的妾 基土拉 所生的兒子，就是 心蘭 、 約珊 、 米但 、 米甸 、 伊施巴 和 書亞 。 約珊 的兒子是 示巴 和 底但 。
1CHR|1|33|米甸 的兒子是 以法 、 以弗 、 哈諾 、 亞比大 和 以勒大 。這些都是 基土拉 的子孫。
1CHR|1|34|亞伯拉罕 生 以撒 ； 以撒 的兒子是 以掃 和 以色列 。
1CHR|1|35|以掃 的兒子是 以利法 、 流珥 、 耶烏施 、 雅蘭 和 可拉 。
1CHR|1|36|以利法 的兒子是 提幔 、 阿抹 、 洗玻 、 迦坦 、 基納斯 、 亭納 和 亞瑪力 。
1CHR|1|37|流珥 的兒子是 拿哈 、 謝拉 、 沙瑪 和 米撒 。
1CHR|1|38|西珥 的兒子是 羅坍 、 朔巴 、 祭便 、 亞拿 、 底順 、 以察 和 底珊 。
1CHR|1|39|羅坍 的兒子是 何利 和 荷幔 ； 羅坍 的妹妹是 亭納 。
1CHR|1|40|朔巴 的兒子是 亞勒文 、 瑪拿轄 、 以巴錄 、 示非 和 阿南 。 祭便 的兒子是 愛亞 和 亞拿 。
1CHR|1|41|亞拿 的兒子是 底順 。 底順 的兒子是 哈默蘭 、 伊是班 、 益蘭 和 基蘭 。
1CHR|1|42|以察 的兒子是 辟罕 、 撒番 ，和 亞干 。 底珊 的兒子是 烏斯 和 亞蘭 。
1CHR|1|43|以色列 人未有君王治理之前，這些是在 以東 地作王的。有 比珥 的兒子 比拉 ，他的城名叫 亭哈巴 。
1CHR|1|44|比拉 死了， 波斯拉 人 謝拉 的兒子 約巴 接續他作王。
1CHR|1|45|約巴 死了， 提幔 人之地的 戶珊 接續他作王。
1CHR|1|46|戶珊 死了， 比達 的兒子 哈達 接續他作王， 哈達 曾在 摩押 地擊敗 米甸 人，他的城名叫 亞未得 。
1CHR|1|47|哈達 死了， 瑪士利加 人 桑拉 接續他作王。
1CHR|1|48|桑拉 死了， 大河 邊的 利河伯 人 掃羅 接續他作王。
1CHR|1|49|掃羅 死了， 亞革波 的兒子 巴勒‧哈南 接續他作王。
1CHR|1|50|巴勒‧哈南 死了， 哈達 接續他作王，他的城名叫 巴伊 。他的妻子名叫 米希她別 ，是 米‧薩合 的孫女， 瑪特列 的女兒。
1CHR|1|51|哈達 死了。 以東 的族長有： 亭納 族長、 亞勒瓦 族長、 耶帖 族長、
1CHR|1|52|阿何利巴瑪 族長、 以拉 族長、 比嫩 族長、
1CHR|1|53|基納斯 族長、 提幔 族長、 米比薩 族長、
1CHR|1|54|瑪基疊 族長、 以蘭 族長。這些都是 以東 的族長。
1CHR|2|1|以色列 的兒子是 呂便 、 西緬 、 利未 、 猶大 、 以薩迦 、 西布倫 、
1CHR|2|2|但 、 約瑟 、 便雅憫 、 拿弗他利 、 迦得 和 亞設 。
1CHR|2|3|猶大 的兒子是 珥 、 俄南 和 示拉 ，這三人是 迦南 女子 拔．書亞 所生的。 猶大 的長子 珥 在耶和華眼中看為惡，耶和華就殺死了他。
1CHR|2|4|猶大 的媳婦 她瑪 為 猶大 生了 法勒斯 和 謝拉 。 猶大 共有五個兒子。
1CHR|2|5|法勒斯 的兒子是 希斯崙 和 哈母勒 。
1CHR|2|6|謝拉 的兒子是 心利 、 以探 、 希幔 、 甲各 和 大拉 ，共五人。
1CHR|2|7|迦米 的兒子是 亞迦 ，他在當滅的物上犯了罪，連累了 以色列 人。
1CHR|2|8|以探 的兒子是 亞撒利雅 。
1CHR|2|9|希斯崙 所生的兒子是 耶拉篾 、 蘭 和 基路拜 。
1CHR|2|10|蘭 生 亞米拿達 ； 亞米拿達 生 拿順 ， 拿順 是 猶大 人的領袖。
1CHR|2|11|拿順 生 撒門 ； 撒門 生 波阿斯 ；
1CHR|2|12|波阿斯 生 俄備得 ； 俄備得 生 耶西 ；
1CHR|2|13|耶西 生長子 以利押 ，次子 亞比拿達 ，三子 示米亞 ，
1CHR|2|14|四子 拿坦業 ，五子 拉代 ，
1CHR|2|15|六子 阿鮮 ，七子 大衛 。
1CHR|2|16|他們的姊妹是 洗魯雅 和 亞比該 。 洗魯雅 的兒子是 亞比篩 、 約押 和 亞撒黑 ，共三人。
1CHR|2|17|亞比該 生 亞瑪撒 ； 亞瑪撒 的父親是 以實瑪利 人 益帖 。
1CHR|2|18|希斯崙 的兒子 迦勒 娶 阿蘇巴 和 耶略 為妻， 阿蘇巴 的兒子是 耶設 、 朔罷 和 押墩 。
1CHR|2|19|阿蘇巴 死了， 迦勒 又娶 以法她 ，生了 戶珥 。
1CHR|2|20|戶珥 生 烏利 ； 烏利 生 比撒列 。
1CHR|2|21|後來， 希斯崙 六十歲時娶了 基列 的父親 瑪吉 的女兒，與她同房； 瑪吉 的女兒為他生了 西割 ；
1CHR|2|22|西割 生 睚珥 。 睚珥 在 基列 地有二十三座城。
1CHR|2|23|後來 基述 和 亞蘭 奪了 哈倭特．睚珥 ，以及 基納 和所屬的鄉鎮 ，共六十個。這些城鎮的人全都是 基列 的父親 瑪吉 的子孫。
1CHR|2|24|希斯崙 在 迦勒‧以法他 死後，他的妻子 亞比雅 為他生了 提哥亞 的父親 亞施戶 。
1CHR|2|25|希斯崙 的長子 耶拉篾 的兒子有長子 蘭 、 布拿 、 阿連 、 阿鮮 和 亞希雅 。
1CHR|2|26|耶拉篾 又娶一妻名叫 亞她拉 ，是 阿南 的母親。
1CHR|2|27|耶拉篾 的長子 蘭 的兒子有 瑪斯 、 雅憫 和 以結 。
1CHR|2|28|阿南 的兒子是 沙買 和 雅大 。 沙買 的兒子是 拿答 和 亞比述 。
1CHR|2|29|亞比述 的妻子名叫 亞比孩 ，為他生了 亞辦 和 摩利 。
1CHR|2|30|拿答 的兒子是 西列 和 亞遍 ； 西列 死了，沒有兒子。
1CHR|2|31|亞遍 的兒子是 以示 ； 以示 的兒子是 示珊 ； 示珊 的兒子是 亞來 。
1CHR|2|32|沙買 的兄弟 雅大 的兒子是 益帖 和 約拿單 ； 益帖 死了，沒有兒子。
1CHR|2|33|約拿單 的兒子是 比勒 和 撒薩 。這些都是 耶拉篾 的子孫。
1CHR|2|34|示珊 沒有兒子，只有女兒。 示珊 有一個僕人名叫 耶哈 ，是 埃及 人。
1CHR|2|35|示珊 把女兒嫁給僕人 耶哈 ，她為他生了 亞太 。
1CHR|2|36|亞太 生 拿單 ； 拿單 生 撒拔 ；
1CHR|2|37|撒拔 生 以弗拉 ； 以弗拉 生 俄備得 ；
1CHR|2|38|俄備得 生 耶戶 ； 耶戶 生 亞撒利雅 ；
1CHR|2|39|亞撒利雅 生 希利斯 ； 希利斯 生 以利亞薩 ；
1CHR|2|40|以利亞薩 生 西斯買 ； 西斯買 生 沙龍 ；
1CHR|2|41|沙龍 生 耶加米雅 ； 耶加米雅 生 以利沙瑪 。
1CHR|2|42|耶拉篾 的兄弟 迦勒 的眾兒子：長子是 米沙 ， 米沙 是 西弗 的父親，還有 希伯倫 的父親 瑪利沙 的眾兒子。
1CHR|2|43|希伯倫 的兒子是 可拉 、 他普亞 、 利肯 和 示瑪 。
1CHR|2|44|示瑪 生 拉含 ，是 約干 之祖。 利肯 生 沙買 。
1CHR|2|45|沙買 的兒子是 瑪雲 ； 瑪雲 是 伯‧夙 的父親。
1CHR|2|46|迦勒 的妾 以法 生 哈蘭 、 摩撒 和 迦謝 ； 哈蘭 生 迦卸 。
1CHR|2|47|雅代 的兒子是 利健 、 約坦 、 基珊 、 毗力 、 以法 和 沙亞弗 。
1CHR|2|48|迦勒 的妾 瑪迦 生 示別 和 特哈拿 ，
1CHR|2|49|又生 麥瑪拿 的父親 沙亞弗 ，又生 抹比拿 和 基比亞 的父親 示法 。 迦勒 的女兒是 押撒 。
1CHR|2|50|這些都是 迦勒 的子孫。 以法她 的長子 戶珥 的子孫： 基列‧耶琳 之祖 朔巴 ，
1CHR|2|51|伯利恆 之祖 薩瑪 ， 伯‧迦得 之祖 哈勒 。
1CHR|2|52|基列‧耶琳 之祖 朔巴 的子孫是 哈羅以 和一半的 米努哈 人 。
1CHR|2|53|基列‧耶琳 的宗族有 以帖 人、 布特 人、 舒瑪 人、 密來 人，又從這些宗族生出 瑣拉 人和 以實陶 人。
1CHR|2|54|薩瑪 的子孫有 伯利恆 人、 尼陀法 人、 亞他綠‧伯‧約押 人、一半的 瑪拿哈 人、 瑣利 人。
1CHR|2|55|住 雅比斯 的文士的宗族有 特拉 人、 示米押 人和 蘇甲 人。這些都是 利甲 家之祖 哈末 所生的 基尼 人。
1CHR|3|1|大衛 在 希伯崙 所生的兒子如下：長子 暗嫩 是 耶斯列 人 亞希暖 生的。次子 但以利 是 迦密 人 亞比該 生的。
1CHR|3|2|三子 押沙龍 是 基述 王 達買 的女兒 瑪迦 生的。四子 亞多尼雅 是 哈及 生的。
1CHR|3|3|五子 示法提雅 是 亞比她 生的。六子 以特念 是 大衛 的妻子 以格拉 生的。
1CHR|3|4|這六人都是 大衛 在 希伯崙 生的。 大衛 在 希伯崙 作王七年六個月，在 耶路撒冷 作王三十三年。
1CHR|3|5|大衛 在 耶路撒冷 所生的兒子是 示米亞 、 朔罷 、 拿單 和 所羅門 。這四人是 亞米利 的女兒 拔‧書亞 生的。
1CHR|3|6|還有 益轄 、 以利沙瑪 、 以利法列 、
1CHR|3|7|挪迦 、 尼斐 、 雅非亞 、
1CHR|3|8|以利沙瑪 、 以利雅大 、 以利法列 ，共九人。
1CHR|3|9|這些全都是 大衛 的兒子，妃嬪的兒子不在其內； 她瑪 是他們的妹妹。
1CHR|3|10|所羅門 的後裔如下： 羅波安 ，他的兒子 亞比雅 ，他的兒子 亞撒 ，他的兒子 約沙法 ，
1CHR|3|11|他的兒子 約蘭 ，他的兒子 亞哈謝 ，他的兒子 約阿施 ，
1CHR|3|12|他的兒子 亞瑪謝 ，他的兒子 亞撒利雅 ，他的兒子 約坦 ；
1CHR|3|13|他的兒子 亞哈斯 ，他的兒子 希西家 ，他的兒子 瑪拿西 ，
1CHR|3|14|他的兒子 亞們 ，他的兒子 約西亞 ，
1CHR|3|15|他的長子 約哈難 ，次子 約雅敬 ，三子 西底家 ，四子 沙龍 。
1CHR|3|16|約雅敬 的後裔：他的兒子 耶哥尼雅 ，他的兒子 西底家 。
1CHR|3|17|被擄的 耶哥尼雅 的後裔如下：他的兒子 撒拉鐵 、
1CHR|3|18|瑪基蘭 、 毗大雅 、 示拿薩 、 耶加米 、 何沙瑪 和 尼大比雅 。
1CHR|3|19|毗大雅 的兒子是 所羅巴伯 和 示每 。 所羅巴伯 的兒子是 米書蘭 和 哈拿尼雅 ， 示羅密 是他們的妹妹；
1CHR|3|20|還有 哈舒巴 、 阿黑 、 比利家 、 哈撒底 、 于沙‧希悉 ，共五人。
1CHR|3|21|哈拿尼雅 的兒子是 毗拉提 和 耶篩亞 。還有 利法雅 的眾兒子， 亞珥難 的眾兒子， 俄巴底亞 的眾兒子， 示迦尼 的眾兒子。
1CHR|3|22|示迦尼 的後裔： 示瑪雅 ， 示瑪雅 的兒子 哈突 、 以甲 、 巴利亞 、 尼利雅 、 沙法 ，共六人。
1CHR|3|23|尼利雅 的兒子是 以利約乃 、 希西家 、 亞斯利干 ，共三人。
1CHR|3|24|以利約乃 的兒子是 何大雅 、 以利亞實 、 毗萊雅 、 阿谷 、 約哈難 、 第萊雅 、 阿拿尼 ，共七人。
1CHR|4|1|猶大 的兒子是 法勒斯 、 希斯崙 、 迦米 、 戶珥 和 朔巴 。
1CHR|4|2|朔巴 的兒子 利亞雅 生 雅哈 ； 雅哈 生 亞戶買 和 拉哈 。這些是 瑣拉 人的宗族。
1CHR|4|3|以坦 之祖 是 耶斯列 、 伊施瑪 和 伊得巴 ；他們的妹妹名叫 哈悉勒玻尼 。
1CHR|4|4|基多 之祖是 毗努伊勒 。 戶沙 之祖是 以謝珥 。這些都是 伯利恆 之祖， 以法她 的長子 戶珥 的後裔。
1CHR|4|5|提哥亞 的父親 亞施戶 有兩個妻子， 希拉 和 拿拉 。
1CHR|4|6|拿拉 為 亞施戶 生 亞戶撒 、 希弗 、 提米尼 和 哈轄斯他利 。這些都是 拿拉 的兒子。
1CHR|4|7|希拉 生的是 洗列 、 瑣轄 和 伊提南 。
1CHR|4|8|哥斯 生 亞諾 、 瑣比巴 和 哈崙 的兒子 亞哈黑 的宗族。
1CHR|4|9|雅比斯 比他眾兄弟更尊貴，他母親給他起名叫 雅比斯 ，意思說：「我生他甚是痛苦。」
1CHR|4|10|雅比斯 求告 以色列 的上帝說：「甚願你賜福與我，擴張我的疆界，你的手常與我同在，保佑我不遭患難，不受艱苦。」上帝就應允他所求的。
1CHR|4|11|書哈 的兄弟 基綠 生 米黑 ， 米黑 是 伊施屯 的父親。
1CHR|4|12|伊施屯 生 伯拉巴 、 巴西亞 和 珥．拿轄 之祖 提欣拿 。這些都是 利迦 人。
1CHR|4|13|基納斯 的兒子是 俄陀聶 和 西萊雅 。 俄陀聶 的兒子是 哈塔 。
1CHR|4|14|憫挪太 生 俄弗拉 ； 西萊雅 生 革‧夏納欣 之祖 約押 。他們都是工匠。
1CHR|4|15|耶孚尼 的兒子 迦勒 的後裔： 以路 、 以拉 和 拿安 。 以拉 的兒子是 基納斯 。
1CHR|4|16|耶哈利勒 的兒子是 西弗 、 西法 、 提利 和 亞撒列 。
1CHR|4|17|以斯拉 的兒子是 益帖 、 米列 、 以弗 和 雅倫 。 米列 所娶法老的女兒 比提雅 的後裔如下：她懷了 米利暗 、 沙買 ，和 以實提摩 之祖 益巴 。 米列 的 猶大 妻子生 基多 之祖 雅列 ， 梭哥 之祖 希伯 ，和 撒挪亞 之祖 耶古鐵 。
1CHR|4|18|
1CHR|4|19|拿含 的妹妹， 荷第雅 的妻子所生的是 達利亞 ， 迦米 人 基伊拉 和 瑪迦 人 以實提摩 的祖先。
1CHR|4|20|示門 的兒子是 暗嫩 、 林拿 、 便‧哈南 和 提倫 。 以示 的兒子是 梭黑 和 便‧梭黑 。
1CHR|4|21|猶大 的兒子 示拉 的後裔： 利迦 之祖 珥 ， 瑪利沙 之祖 拉大 ，和住在 伯‧亞實比 織細麻布的各宗族。
1CHR|4|22|還有 約敬 、 哥西巴 人、 約阿施 ，和那在 摩押 娶妻，回到 利恆 的 薩拉 。這都是古時的記載。
1CHR|4|23|這些人都是陶匠，是 尼他應 和 基底拉 的居民。他們住在王那裏，為王做工。
1CHR|4|24|西緬 的後裔如下： 尼母利 、 雅憫 、 雅立 、 謝拉 和 掃羅 ；
1CHR|4|25|他的兒子 沙龍 ，他的兒子 米比衫 ，他的兒子 米施瑪 ；
1CHR|4|26|米施瑪 的後裔：他的兒子 哈母利 ，他的兒子 撒刻 ，他的兒子 示每 。
1CHR|4|27|示每 有十六個兒子和六個女兒，但他兄弟的兒女不多，他們各家族也不如 猶大 族那樣人丁興旺。
1CHR|4|28|西緬 人住在 別是巴 、 摩拉大 、 哈薩‧書亞 、
1CHR|4|29|辟拉 、 以森 、 陀臘 、
1CHR|4|30|彼土利 、 何珥瑪 、 洗革拉 、
1CHR|4|31|伯‧瑪加博 、 哈薩‧蘇撒 、 伯‧比利 和 沙拉音 ，這些城鎮直到 大衛 作王的時候都是屬 西緬 人的；
1CHR|4|32|還有所屬的村莊 以坦 、 亞因 、 臨門 、 陀健 、 亞珊 ，共五個城鎮；
1CHR|4|33|連同環繞這些城鎮的一切鄉村，直到 巴力 。這是他們的住處，他們都有家譜。
1CHR|4|34|還有 米所巴 、 雅米勒 、 亞瑪謝 的兒子 約沙 、
1CHR|4|35|約珥 ，和 亞薛 的曾孫， 西萊雅 的孫子， 約示比 的兒子 耶戶 。
1CHR|4|36|還有 以利約乃 、 雅哥巴 、 約朔海 、 亞帥雅 、 亞底業 、 耶西篾 、 比拿雅 、
1CHR|4|37|細撒 ； 細撒 是 示非 的兒子， 示非 是 亞龍 的兒子， 亞龍 是 耶大雅 的兒子， 耶大雅 是 申利 的兒子， 申利 是 示瑪雅 的兒子。
1CHR|4|38|以上所記的人名都是作族長的，他們父系的家屬大量增加。
1CHR|4|39|他們往平原東邊 基多口 去，尋找牧放羊群的草場，
1CHR|4|40|找到了肥沃優美的草場，又寬闊又平靜安寧之地；從前住那裏的是 含 族的人。
1CHR|4|41|以上紀錄上有名的人，在 猶大 王 希西家 的日子，來攻擊 含 族人的帳棚和那裏所有的 米烏尼 人，把他們滅盡，就住在他們的地方，直到今日，因為那裏有草場可以牧放羊群。
1CHR|4|42|這些 西緬 人中有五百人上 西珥山 ，率領他們的是 以示 的兒子 毗拉提 、 尼利雅 、 利法雅 和 烏薛 。
1CHR|4|43|他們殺了 亞瑪力 剩下的殘存之民，就住在那裏，直到今日。
1CHR|5|1|以色列 的長子 呂便 的後裔。 呂便 玷污了父親的床，他長子的名分就歸了 以色列 的兒子 約瑟 的後裔；因此，家譜就不按出生順序登錄。
1CHR|5|2|雖然 猶大 比他兄弟強盛，君王也從他而出，然而長子的名分卻歸 約瑟 。
1CHR|5|3|以色列 長子 呂便 的後裔如下： 哈諾 、 法路 、 希斯倫 和 迦米 。
1CHR|5|4|約珥 的後裔：他的兒子 示瑪雅 ，他的兒子 歌革 ，他的兒子 示每 ，
1CHR|5|5|他的兒子 米迦 ，他的兒子 利亞雅 ，他的兒子 巴力 ，
1CHR|5|6|他的兒子 備拉 ；這 備拉 作 呂便 支派的領袖，被 亞述 王 提革拉‧毗列色 擄去。
1CHR|5|7|他的弟兄照著宗族，按著家譜作族長的是 耶利 、 撒迦利雅 、
1CHR|5|8|比拉 ； 比拉 是 亞撒 的兒子， 亞撒 是 示瑪 的兒子， 示瑪 是 約珥 的兒子； 約珥 住在 亞羅珥 ，直到 尼波 和 巴力‧免 。
1CHR|5|9|他也住在東邊，直到 幼發拉底河 這邊的曠野邊界，因為他們在 基列 地牲畜增多。
1CHR|5|10|掃羅 年間，他們與 夏甲 人爭戰， 夏甲 人倒在他們手下，他們就在 基列 東邊的全地，住在 夏甲 人的帳棚裏。
1CHR|5|11|迦得 的後裔在 呂便 對面，住在 巴珊 地，延伸到 撒迦 ：
1CHR|5|12|有作族長的 約珥 ，有作副族長的 沙番 ，還有 雅乃 和住在 巴珊 的 沙法 。
1CHR|5|13|按著家族，他們的弟兄是 米迦勒 、 米書蘭 、 示巴 、 約賴 、 雅干 、 細亞 和 希伯 ，共七人。
1CHR|5|14|這些都是 亞比孩 的兒子； 亞比孩 是 戶利 的兒子， 戶利 是 耶羅亞 的兒子， 耶羅亞 是 基列 的兒子， 基列 是 米迦勒 的兒子， 米迦勒 是 耶示篩 的兒子， 耶示篩 是 耶哈多 的兒子， 耶哈多 是 布斯 的兒子；
1CHR|5|15|古尼 的孫子， 押比疊 的兒子 亞希 是他們的族長。
1CHR|5|16|他們住在 基列 、 巴珊 和所屬的鄉鎮，以及 沙崙 一切的郊野，直到四圍的交界。
1CHR|5|17|這些人在 猶大 王 約坦 和 以色列 王 耶羅波安 年間，都載入家譜。
1CHR|5|18|呂便 人、 迦得 人和 瑪拿西 半支派的人，能拿盾牌和刀劍、拉弓、出征善戰的勇士共有四萬四千七百六十名。
1CHR|5|19|他們與 夏甲 人、 伊突 人、 拿非施 人、 挪答 人打仗。
1CHR|5|20|他們在打仗的時候得了上帝的幫助， 夏甲 人和所有跟隨 夏甲 人的人都交在他們手中；因為他們在陣上呼求上帝，倚賴他，他就應允他們。
1CHR|5|21|他們擄掠了 夏甲 人的牲畜，有五萬匹駱駝，二十五萬隻羊，二千匹驢，又有十萬人；
1CHR|5|22|被殺仆倒的很多，因為這戰爭是出乎上帝。他們就住在 夏甲 人的地上，直到被擄的時候。
1CHR|5|23|瑪拿西 半支派的人住在那地，從 巴珊 延到 巴力‧黑門 、 示尼珥 和 黑門山 ，他們人數增多 。
1CHR|5|24|他們的族長如下： 以弗 、 以示 、 以利業 、 亞斯列 、 耶利米 、 何達威雅 和 雅疊 ；他們都是大能的勇士，有名的人，是作族長的。
1CHR|5|25|但他們得罪了他們列祖的上帝，隨從當地百姓的神明而行淫，這百姓就是上帝在他們面前所除滅的。
1CHR|5|26|因此， 以色列 的上帝激發 亞述 王 普勒 ，就是 亞述 王 提革拉‧毗列色 的心，他擄掠了 呂便 人、 迦得 人、 瑪拿西 半支派的人，把他們帶到 哈臘 、 哈博 、 哈拉 與 歌散河 邊，直到今日。
1CHR|6|1|利未 的後裔： 革順 、 哥轄 和 米拉利 。
1CHR|6|2|哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 和 烏薛 。
1CHR|6|3|暗蘭 的兒女是 亞倫 、 摩西 和 米利暗 。 亞倫 的兒子是 拿答 、 亞比戶 、 以利亞撒 和 以他瑪 。
1CHR|6|4|以利亞撒 生 非尼哈 ； 非尼哈 生 亞比書 ；
1CHR|6|5|亞比書 生 布基 ； 布基 生 烏西 ；
1CHR|6|6|烏西 生 西拉希雅 ； 西拉希雅 生 米拉約 ；
1CHR|6|7|米拉約 生 亞瑪利雅 ； 亞瑪利雅 生 亞希突 ；
1CHR|6|8|亞希突 生 撒督 ； 撒督 生 亞希瑪斯 ；
1CHR|6|9|亞希瑪斯 生 亞撒利雅 ； 亞撒利雅 生 約哈難 ；
1CHR|6|10|約哈難 生 亞撒利雅 ， 亞撒利雅 在 所羅門 建造的 耶路撒冷 殿中擔任祭司的職分；
1CHR|6|11|亞撒利雅 生 亞瑪利雅 ； 亞瑪利雅 生 亞希突 ；
1CHR|6|12|亞希突 生 撒督 ； 撒督 生 沙龍 ；
1CHR|6|13|沙龍 生 希勒家 ； 希勒家 生 亞撒利雅 ；
1CHR|6|14|亞撒利雅 生 西萊雅 ； 西萊雅 生 約薩答 。
1CHR|6|15|當耶和華藉 尼布甲尼撒 的手擄掠 猶大 和 耶路撒冷 的時候， 約薩答 也被擄去。
1CHR|6|16|利未 的後裔： 革順 、 哥轄 和 米拉利 。
1CHR|6|17|革順 的兒子名叫 立尼 和 示每 。
1CHR|6|18|哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 和 烏薛 。
1CHR|6|19|米拉利 的兒子是 抹利 和 母示 。這是按著父系所分 利未 人的宗族。
1CHR|6|20|屬 革順 的：他的兒子 立尼 ，他的兒子 雅哈 ，他的兒子 薪瑪 ，
1CHR|6|21|他的兒子 約亞 ，他的兒子 易多 ，他的兒子 謝拉 ，他的兒子 耶特賴 。
1CHR|6|22|哥轄 的後裔：他的兒子 亞米拿達 ，他的兒子 可拉 ，他的兒子 亞惜 ，
1CHR|6|23|他的兒子 以利加拿 ，他的兒子 以比雅撒 ，他的兒子 亞惜 ，
1CHR|6|24|他的兒子 他哈 ，他的兒子 烏列 ，他的兒子 烏西雅 ，他的兒子 少羅 。
1CHR|6|25|以利加拿 的兒子是 亞瑪賽 、 亞希摩 、
1CHR|6|26|以利加拿 。 以利加拿 的後裔：他的兒子 瑣菲 ，他的兒子 拿哈 ，
1CHR|6|27|他的兒子 以利押 ，他的兒子 耶羅罕 ，他的兒子 以利加拿 ，他的兒子 撒母耳 。
1CHR|6|28|撒母耳 的兒子是長子 約珥 和次子 亞比亞 。
1CHR|6|29|米拉利 的後裔： 抹利 ，他的兒子 立尼 ，他的兒子 示每 ，他的兒子 烏撒 ，
1CHR|6|30|他的兒子 示米亞 ，他的兒子 哈基雅 ，他的兒子 亞帥雅 。
1CHR|6|31|這些是約櫃安設之後， 大衛 派在耶和華殿中管理歌唱事奉的人。
1CHR|6|32|他們在會幕前負責歌唱的事奉，及至 所羅門 在 耶路撒冷 建造了耶和華的殿，他們就按著班次供職。
1CHR|6|33|供職的人和他們的子孫如下： 哥轄 的子孫中有歌唱的 希幔 ； 希幔 是 約珥 的兒子， 約珥 是 撒母耳 的兒子，
1CHR|6|34|撒母耳 是 以利加拿 的兒子， 以利加拿 是 耶羅罕 的兒子， 耶羅罕 是 以利業 的兒子， 以利業 是 陀亞 的兒子，
1CHR|6|35|陀亞 是 蘇弗 的兒子， 蘇弗 是 以利加拿 的兒子， 以利加拿 是 瑪哈 的兒子， 瑪哈 是 亞瑪賽 的兒子，
1CHR|6|36|亞瑪賽 是 以利加拿 的兒子， 以利加拿 是 約珥 的兒子， 約珥 是 亞撒利雅 的兒子， 亞撒利雅 是 西番雅 的兒子，
1CHR|6|37|西番雅 是 他哈 的兒子， 他哈 是 亞惜 的兒子， 亞惜 是 以比雅撒 的兒子， 以比雅撒 是 可拉 的兒子，
1CHR|6|38|可拉 是 以斯哈 的兒子， 以斯哈 是 哥轄 的兒子， 哥轄 是 利未 的兒子， 利未 是 以色列 的兒子。
1CHR|6|39|希幔 的弟兄 亞薩 在 希幔 的右邊供職； 亞薩 是 比利家 的兒子， 比利家 是 示米亞 的兒子，
1CHR|6|40|示米亞 是 米迦勒 的兒子， 米迦勒 是 巴西雅 的兒子， 巴西雅 是 瑪基雅 的兒子，
1CHR|6|41|瑪基雅 是 伊特尼 的兒子， 伊特尼 是 謝拉 的兒子， 謝拉 是 亞大雅 的兒子，
1CHR|6|42|亞大雅 是 以探 的兒子， 以探 是 薪瑪 的兒子， 薪瑪 是 示每 的兒子，
1CHR|6|43|示每 是 雅哈 的兒子， 雅哈 是 革順 的兒子， 革順 是 利未 的兒子。
1CHR|6|44|他們的弟兄 米拉利 的子孫，在他們左邊供職的有 以探 ； 以探 是 基示 的兒子， 基示 是 亞伯底 的兒子， 亞伯底 是 瑪鹿 的兒子，
1CHR|6|45|瑪鹿 是 哈沙比雅 的兒子， 哈沙比雅 是 亞瑪謝 的兒子， 亞瑪謝 是 希勒家 的兒子，
1CHR|6|46|希勒家 是 暗西 的兒子， 暗西 是 巴尼 的兒子， 巴尼 是 沙麥 的兒子，
1CHR|6|47|沙麥 是 末力 的兒子， 末力 是 母示 的兒子， 母示 是 米拉利 的兒子， 米拉利 是 利未 的兒子。
1CHR|6|48|他們的弟兄 利未 人也被派辦理上帝殿中帳幕的一切事務。
1CHR|6|49|亞倫 和他的子孫在燔祭壇和香壇上獻祭燒香，辦理至聖所一切的事，為 以色列 贖罪，正如上帝僕人 摩西 所吩咐的一切。
1CHR|6|50|亞倫 的後裔如下：他的兒子 以利亞撒 ，他的兒子 非尼哈 ，他的兒子 亞比書 ，
1CHR|6|51|他的兒子 布基 ，他的兒子 烏西 ，他的兒子 西拉希雅 ，
1CHR|6|52|他的兒子 米拉約 ，他的兒子 亞瑪利雅 ，他的兒子 亞希突 ，
1CHR|6|53|他的兒子 撒督 ，他的兒子 亞希瑪斯 。
1CHR|6|54|他們的住處按著境內的營寨如下： 亞倫 的子孫 哥轄 族先抽籤得地，
1CHR|6|55|得了 猶大 地的 希伯崙 和四圍的郊野；
1CHR|6|56|只是這城的田地和所屬的村莊都為 耶孚尼 的兒子 迦勒 所得。
1CHR|6|57|亞倫 的子孫所得逃城如下： 希伯崙 、 立拿 與其郊野、 雅提珥 、 以實提莫 與其郊野、
1CHR|6|58|希崙 與其郊野、 底璧 與其郊野、
1CHR|6|59|亞珊 與其郊野、 伯‧示麥 與其郊野。
1CHR|6|60|他們也從 便雅憫 支派中得了 迦巴 與其郊野、 阿勒篾 與其郊野、 亞拿突 與其郊野。他們宗族所得的城共十三座。
1CHR|6|61|哥轄 族其餘的人抽籤，按支派的宗族，從半個支派，就是 瑪拿西 半支派中得了十座城。
1CHR|6|62|革順 族按著宗族，從 以薩迦 支派、 亞設 支派、 拿弗他利 支派、 巴珊 內的 瑪拿西 支派中，得了十三座城。
1CHR|6|63|米拉利 族按著宗族抽籤，從 呂便 支派、 迦得 支派、 西布倫 支派中，得了十二座城。
1CHR|6|64|以色列 人把這些城與其郊野給了 利未 人。
1CHR|6|65|以色列 人用抽籤的方式，從 猶大 人、 西緬 人、 便雅憫 人三支派中，把以上提到名字的城給了他們。
1CHR|6|66|哥轄 子孫中有幾個宗族從 以法蓮 支派中也得了城鎮作為他們的區域。
1CHR|6|67|他們在 以法蓮 山區所得的逃城： 示劍 與其郊野、 基色 與其郊野、
1CHR|6|68|約緬 與其郊野、 伯‧和崙 與其郊野、
1CHR|6|69|亞雅崙 與其郊野、 迦特‧臨門 與其郊野。
1CHR|6|70|哥轄 其餘的子孫從 瑪拿西 半支派中得了 亞乃 與其郊野、 比連 與其郊野。
1CHR|6|71|革順 子孫從 瑪拿西 半支派中得了 巴珊 的 哥蘭 與其郊野、 亞斯她錄 與其郊野；
1CHR|6|72|從 以薩迦 支派中得了 基低斯 與其郊野、 大比拉 與其郊野、
1CHR|6|73|拉末 與其郊野、 亞年 與其郊野；
1CHR|6|74|從 亞設 支派中得了 瑪沙 與其郊野、 押頓 與其郊野、
1CHR|6|75|戶割 與其郊野、 利合 與其郊野；
1CHR|6|76|從 拿弗他利 支派中得了 加利利 的 基低斯 與其郊野、 哈們 與其郊野、 基列亭 與其郊野。
1CHR|6|77|米拉利 其餘的子孫從 西布倫 支派中得了 臨摩挪 與其郊野、 他泊 與其郊野；
1CHR|6|78|又在 耶利哥 的 約旦河 東，從 呂便 支派中得了曠野的 比悉 與其郊野、 雅雜 與其郊野，
1CHR|6|79|基底莫 與其郊野、 米法押 與其郊野；
1CHR|6|80|又從 迦得 支派中得了 基列 的 拉末 與其郊野、 瑪哈念 與其郊野、
1CHR|6|81|希實本 與其郊野、 雅謝 與其郊野。
1CHR|7|1|以薩迦 的後裔： 陀拉 、 普瓦 、 雅述 和 伸崙 ，共四人。
1CHR|7|2|陀拉 的後裔： 烏西 、 利法雅 、 耶勒 、 雅買 、 易伯散 和 示母利 ，都是 陀拉 的族長，在他們世代中是大能的勇士。到 大衛 年間，他們的人數共有二萬二千六百名。
1CHR|7|3|烏西 的後裔： 伊斯拉希 ， 伊斯拉希 的兒子 米迦勒 、 俄巴底亞 、 約珥 和 伊示雅 ，共五人，全都是族長。
1CHR|7|4|他們所率領的，按著家譜，照著父家，可作戰的軍隊共有三萬六千人，因為他們的妻子和兒子眾多。
1CHR|7|5|他們的弟兄在 以薩迦 各族中的大能勇士，登記在家譜中的全部共有八萬七千人。
1CHR|7|6|便雅憫 ： 比拉 、 比結 和 耶疊 ，共三人。
1CHR|7|7|比拉 的兒子： 以斯本 、 烏西 、 烏薛 、 耶利末 和 以利 ，共五人，都是族長，是大能的勇士。登記在家譜中的人共有二萬二千零三十四人。
1CHR|7|8|比結 的兒子： 細米拉 、 約阿施 、 以利以謝 、 以利約乃 、 暗利 、 耶列末 、 亞比雅 、 亞拿突 和 亞拉篾 ；這些全都是 比結 的兒子。
1CHR|7|9|登記在家譜中，按家譜的族長，大能的勇士，共有二萬零二百人。
1CHR|7|10|耶疊 的後裔： 比勒罕 ， 比勒罕 的兒子 耶烏施 、 便雅憫 、 以笏 、 基拿拿 、 細坦 、 他施 和 亞希沙哈 。
1CHR|7|11|這些全都是 耶疊 的後裔，都是族長，是大能的勇士，能上陣打仗的共有一萬七千二百人。
1CHR|7|12|還有 以珥 的兒子 書品 和 戶品 ，以及 亞黑 的兒子 戶伸 。
1CHR|7|13|拿弗他利 的後裔： 雅薛 、 沽尼 、 耶色 和 沙龍 ，都是 辟拉 的子孫。
1CHR|7|14|瑪拿西 的兒子 亞斯烈 是他的妾 亞蘭 女子所生的；她又生了 瑪吉 ，是 基列 的父親。
1CHR|7|15|瑪吉 為 戶品 和 書品 各娶了一妻，他的姊妹名叫 瑪迦 。第二個名叫 西羅非哈 ； 西羅非哈 只有女兒。
1CHR|7|16|瑪吉 的妻子 瑪迦 生了一個兒子， 瑪迦 給他起名叫 毗利施 。 毗利施 的弟弟名叫 示利施 ； 示利施 的兒子是 烏蘭 和 利金 。
1CHR|7|17|烏蘭 的兒子是 比但 。這些都是 基列 的子孫； 基列 是 瑪吉 的兒子， 瑪吉 是 瑪拿西 的兒子。
1CHR|7|18|基列 的妹妹 哈摩利吉 生了 伊施荷 、 亞比以謝 和 瑪拉 。
1CHR|7|19|示米大 的兒子是 亞現 、 示劍 、 利克希 和 阿尼安 。
1CHR|7|20|以法蓮 的後裔： 書提拉 ，他的兒子 比列 ，他的兒子 他哈 ，他的兒子 以拉大 ，他的兒子 他哈 ，
1CHR|7|21|他的兒子 撒拔 ，他的兒子 書提拉 。 以法蓮 又生 以謝 和 以列 ；這二人因為下去奪取 迦特 人的牲畜，被本地的 迦特 人殺了。
1CHR|7|22|他們的父親 以法蓮 為他們悲哀了多日，他的兄弟都來安慰他。
1CHR|7|23|以法蓮 與妻子同房，妻子懷孕生了一子， 以法蓮 因為家裏遭禍，就給這兒子起名叫 比利亞 。
1CHR|7|24|他的女兒名叫 舍伊拉 ， 舍伊拉 建築了 上伯‧和崙 、 下伯‧和崙 和 烏羨‧舍伊拉 。
1CHR|7|25|他的兒子 利法 和 利悉 ，他的兒子 他拉 ，他的兒子 他罕 ，
1CHR|7|26|他的兒子 拉但 ，他的兒子 亞米忽 ，他的兒子 以利沙瑪 ，
1CHR|7|27|他的兒子 嫩 ，他的兒子 約書亞 。
1CHR|7|28|以法蓮 人的地業和住處是 伯特利 和所屬的鄉鎮，東邊 拿蘭 ，西邊 基色 和所屬的鄉鎮， 示劍 和所屬的鄉鎮，直到 艾雅 和所屬的鄉鎮；
1CHR|7|29|還有靠近 瑪拿西 人的邊界， 伯‧善 和所屬的鄉鎮， 他納 和所屬的鄉鎮， 米吉多 和所屬的鄉鎮， 多珥 和所屬的鄉鎮。 以色列 兒子 約瑟 的子孫住在這些地方。
1CHR|7|30|亞設 的後裔： 音拿 、 亦施瓦 、 亦施韋 和 比利亞 ，還有他們的妹妹 西拉 。
1CHR|7|31|比利亞 的兒子是 希別 和 瑪結 ； 瑪結 是 比撒威 的父親。
1CHR|7|32|希別 生 雅弗勒 、 朔默 、 何坦 和他們的妹妹 書雅 。
1CHR|7|33|雅弗勒 的兒子是 巴薩 、 賓哈 和 亞施法 ；這些都是 雅弗勒 的兒子。
1CHR|7|34|朔默 的兒子是 亞希 、 羅迦 、 耶戶巴 和 亞蘭 。
1CHR|7|35|朔默 的兄弟 希連 的兒子是 瑣法 、 音那 、 示利斯 和 亞抹 。
1CHR|7|36|瑣法 的兒子是 書亞 、 哈尼弗 、 書阿勒 、 比利 、 音拉 、
1CHR|7|37|比悉 、 河得 、 珊瑪 、 施沙 、 益蘭 和 比拉 。
1CHR|7|38|益帖 的兒子是 耶孚尼 、 毗斯巴 和 亞拉 。
1CHR|7|39|烏拉 的兒子是 亞拉 、 漢尼業 和 利寫 。
1CHR|7|40|這些全都是 亞設 的子孫，都是族長，是精壯大能的勇士，也是領袖中的領袖。登記在家譜中，能上陣打仗的共有二萬六千人。
1CHR|8|1|便雅憫 生長子 比拉 ，次子 亞實別 ，三子 亞哈拉 ，
1CHR|8|2|四子 挪哈 ，五子 拉法 。
1CHR|8|3|比拉 的兒子是 亞大 、 基拉 、 亞比忽 、
1CHR|8|4|亞比書 、 乃幔 、 亞何亞 、
1CHR|8|5|基拉 、 示孚汛 和 戶蘭 。
1CHR|8|6|以忽 的後裔如下，他們是 迦巴 居民的族長，曾被擄到 瑪拿轄 ：
1CHR|8|7|乃幔 、 亞希亞 、 基拉 ；他擄了他們，又生了 烏撒 和 亞希忽 。
1CHR|8|8|沙哈連 休了兩個妻子 戶伸 和 巴拉 之後，在 摩押 地生了兒子。
1CHR|8|9|他與妻子 賀得 生了 約巴 、 洗比雅 、 米沙 、 瑪拉干 、
1CHR|8|10|耶烏斯 、 沙迦 和 米瑪 ；這些是他的兒子，都是族長。
1CHR|8|11|戶伸 為他生了 亞比突 和 以利巴力 。
1CHR|8|12|以利巴力 的兒子是 希伯 、 米珊 和 沙麥 ； 沙麥 建立 阿挪 、 羅德 和所屬的鄉鎮。
1CHR|8|13|比利亞 和 示瑪 是 亞雅崙 居民的族長，他們驅逐了 迦特 的居民。
1CHR|8|14|亞希約 、 沙煞 、 耶列末 、
1CHR|8|15|西巴第雅 、 亞拉得 、 亞得 、
1CHR|8|16|米迦勒 、 伊施巴 和 約哈 都是 比利亞 的兒子。
1CHR|8|17|西巴第雅 、 米書蘭 、 希西基 、 希伯 、
1CHR|8|18|伊施米萊 、 伊斯利亞 和 約巴 都是 以利巴力 的兒子。
1CHR|8|19|雅金 、 細基利 、 撒底 、
1CHR|8|20|以利乃 、 洗勒太 、 以利業 、
1CHR|8|21|亞大雅 、 比拉雅 和 申拉 都是 示每 的兒子。
1CHR|8|22|伊施班 、 希伯 、 以利業 、
1CHR|8|23|亞伯頓 、 細基利 、 哈難 、
1CHR|8|24|哈拿尼雅 、 以攔 、 安陀提雅 、
1CHR|8|25|伊弗底雅 、 毗努伊勒 都是 沙煞 的兒子。
1CHR|8|26|珊示萊 、 示哈利 、 亞他利雅 、
1CHR|8|27|雅利西 、 以利亞 和 細基利 都是 耶羅罕 的兒子。
1CHR|8|28|這些人按照他們的家譜都是族長，是領袖，都住在 耶路撒冷 。
1CHR|8|29|在 基遍 住的有 基遍 的父親 耶利 ，他的妻子名叫 瑪迦 ；
1CHR|8|30|他的長子是 亞伯頓 ，還有 蘇珥 、 基士 、 巴力 、 拿答 、
1CHR|8|31|基多 、 亞希約 和 撒迦 。
1CHR|8|32|米基羅 生 示米暗 。這些人在他們弟兄的對面，和他們的弟兄同住在 耶路撒冷 。
1CHR|8|33|尼珥 生 基士 ； 基士 生 掃羅 ； 掃羅 生 約拿單 、 麥基‧舒亞 、 亞比拿達 和 伊施巴力 。
1CHR|8|34|約拿單 的兒子是 米力‧巴力 ； 米力‧巴力 生 米迦 。
1CHR|8|35|米迦 的兒子是 毗敦 、 米勒 、 他利亞 和 亞哈斯 ；
1CHR|8|36|亞哈斯 生 耶何阿達 ； 耶何阿達 生 亞拉篾 、 亞斯瑪威 和 心利 ； 心利 生 摩撒 ；
1CHR|8|37|摩撒 生 比尼亞 ； 比尼亞 的兒子是 拉法 ， 拉法 的兒子是 以利亞薩 ， 以利亞薩 的兒子是 亞悉 。
1CHR|8|38|亞悉 有六個兒子，他們的名字是 亞斯利干 、 波基路 、 以實瑪利 、 示亞利雅 、 俄巴底雅 和 哈難 ；這些全都是 亞悉 的兒子。
1CHR|8|39|亞悉 兄弟 以設 的兒子：長子是 烏蘭 ，次子是 耶烏施 ，三子是 以利法列 。
1CHR|8|40|烏蘭 的兒子都是大能的勇士，是弓箭手，他們有許多的子孫，共一百五十名，都是 便雅憫 人。
1CHR|9|1|以色列 眾人按家譜登記，看哪，都寫在《以色列諸王記》上。 猶大 人因背叛被擄到 巴比倫 。
1CHR|9|2|從 巴比倫 先回來，住在自己地業城鎮中的有 以色列 人、祭司、 利未 人和殿役。
1CHR|9|3|住在 耶路撒冷 的有 猶大 人、 便雅憫 人、 以法蓮 人和 瑪拿西 人：
1CHR|9|4|猶大 兒子 法勒斯 的子孫中有 烏太 ， 烏太 是 亞米忽 的兒子， 亞米忽 是 暗利 的兒子， 暗利 是 音利 的兒子， 音利 是 巴尼 的兒子；
1CHR|9|5|示羅 人中有長子 亞帥雅 和他的眾兒子；
1CHR|9|6|謝拉 的子孫中有 耶烏利 和他的弟兄，共六百九十人；
1CHR|9|7|便雅憫 人中有 哈西努亞 的曾孫， 何達威雅 的孫子， 米書蘭 的兒子 撒路 ；
1CHR|9|8|又有 耶羅罕 的兒子 伊比內雅 ； 米基立 的孫子， 烏西 的兒子 以拉 ； 伊比尼雅 的曾孫， 流珥 的孫子， 示法提雅 的兒子 米書蘭 ；
1CHR|9|9|和他們的弟兄，按著家譜登記，共有九百五十六名；這些人都是族長。
1CHR|9|10|祭司中有 耶大雅 、 耶何雅立 、 雅斤 ，
1CHR|9|11|還有管理上帝殿的 亞撒利雅 ， 亞撒利雅 是 希勒家 的兒子， 希勒家 是 米書蘭 的兒子， 米書蘭 是 撒督 的兒子， 撒督 是 米拉約 的兒子， 米拉約 是 亞希突 的兒子。
1CHR|9|12|還有 瑪基雅 的曾孫， 巴施戶珥 的孫子， 耶羅罕 的兒子 亞大雅 ；又有 瑪賽 ， 瑪賽 是 亞第業 的兒子， 亞第業 是 雅希細拉 的兒子， 雅希細拉 是 米書蘭 的兒子， 米書蘭 是 米實利密 的兒子， 米實利密 是 音麥 的兒子。
1CHR|9|13|他們和他們的弟兄都是族長，共有一千七百六十人，都善於做上帝殿的事工。
1CHR|9|14|利未 人 米拉利 的子孫中有 哈沙比雅 的曾孫， 押利甘 的孫子， 哈述 的兒子 示瑪雅 ；
1CHR|9|15|有 拔巴甲 、 黑勒施 、 加拉 和 亞薩 的曾孫， 細基利 的孫子， 米迦 的兒子 瑪探雅 ；
1CHR|9|16|又有 耶杜頓 的曾孫， 加拉 的孫子， 示瑪雅 的兒子 俄巴底 ，還有 以利加拿 的孫子， 亞撒 的兒子 比利家 。他們都住在 尼陀法 人的村莊。
1CHR|9|17|守衛是 沙龍 、 亞谷 、 達們 、 亞希幔 和他們的弟兄； 沙龍 是領袖。
1CHR|9|18|從前這些人看守朝東的王門，如今是 利未 人營中的守衛。
1CHR|9|19|可拉 的曾孫， 以比雅撒 的孫子， 可利 的兒子 沙龍 ，和他父家的弟兄 可拉 人管理事務，看守會幕的門。他們的祖宗曾管理耶和華的軍營，把守營的入口。
1CHR|9|20|從前 以利亞撒 的兒子 非尼哈 管理他們，耶和華也與他同在。
1CHR|9|21|米施利米雅 的兒子 撒迦利雅 是看守會幕門口的。
1CHR|9|22|被選作門口守衛的總共有二百一十二名。他們在自己的村莊，按著家譜登記，是 大衛 和 撒母耳 先見所派擔當這受託之職任的。
1CHR|9|23|他們和他們的子孫看守耶和華殿的門，就是會幕的門口。
1CHR|9|24|在東西南北，四方 都有守衛。
1CHR|9|25|他們的弟兄住在村莊，每七日來與他們換班。
1CHR|9|26|這些守衛的四個領袖都是 利未 人，各有受託的職任，看守上帝殿的房間和寶庫。
1CHR|9|27|他們住在上帝殿的四圍，受託看守聖殿，負責每日早晨開門。
1CHR|9|28|利未 人中有人管理所使用的器皿，拿出拿入都按數目點算。
1CHR|9|29|又有人管理器具和聖所一切的器皿，以及細麵、酒、油、乳香和香料。
1CHR|9|30|祭司的子孫中有人用香料做膏油。
1CHR|9|31|利未 人 瑪他提雅 是 可拉 族 沙龍 的長子，他受託做烤餅。
1CHR|9|32|他們弟兄 哥轄 子孫中，有人負責每安息日排列供餅。
1CHR|9|33|歌唱的有 利未 人的族長，住在殿的房間，晝夜供職，不做別樣的工。
1CHR|9|34|以上都是 利未 人的族長，按各世系作領袖，他們都住在 耶路撒冷 。
1CHR|9|35|在 基遍 住的有 基遍 的父親 耶利 ，他的妻子名叫 瑪迦 ；
1CHR|9|36|他的長子是 亞伯頓 ，還有 蘇珥 、 基士 、 巴力 、 尼珥 、 拿答 、
1CHR|9|37|基多 、 亞希約 、 撒迦利雅 和 米基羅 。
1CHR|9|38|米基羅 生 示米暗 。這些人在他們弟兄的對面，和他們的弟兄同住在 耶路撒冷 。
1CHR|9|39|尼珥 生 基士 ； 基士 生 掃羅 ； 掃羅 生 約拿單 、 麥基‧舒亞 、 亞比拿達 和 伊施巴力 。
1CHR|9|40|約拿單 的兒子是 米力‧巴力 ； 米力‧巴力 生 米迦 。
1CHR|9|41|米迦 的兒子是 毗敦 、 米勒 、 他利亞 和 亞哈斯 。
1CHR|9|42|亞哈斯 生 雅拉 ； 雅拉 生 亞拉篾 、 亞斯瑪威 和 心利 ； 心利 生 摩撒 ；
1CHR|9|43|摩撒 生 比尼亞 ； 比尼亞 的兒子是 利法雅 ， 利法雅 的兒子是 以利亞薩 ， 以利亞薩 的兒子是 亞悉 。
1CHR|9|44|亞悉 有六個兒子，他們的名字是 亞斯利干 、 波基路 、 以實瑪利 、 示亞利雅 、 俄巴底雅 和 哈難 ；這些都是 亞悉 的兒子。
1CHR|10|1|非利士 人攻打 以色列 。 以色列 人在 非利士 人面前逃跑，很多人 在 基利波山 被殺仆倒。
1CHR|10|2|非利士 人緊追 掃羅 和他的兒子，殺了 掃羅 的兒子 約拿單 、 亞比拿達 、 麥基‧舒亞 。
1CHR|10|3|攻擊 掃羅 的戰事激烈， 掃羅 被弓箭手射中，被他們射傷。
1CHR|10|4|掃羅 吩咐拿他兵器的人說：「你拔出刀來，把我刺死，免得那些未受割禮的人來凌辱我。」但拿兵器的人非常懼怕，不肯刺他。於是 掃羅 拿起刀來，伏在刀上。
1CHR|10|5|拿兵器的人見 掃羅 已死，也伏在刀上死了。
1CHR|10|6|這樣， 掃羅 和他三個兒子，以及他的全家都一起陣亡了。
1CHR|10|7|住平原的 以色列 眾人見 以色列 軍兵 逃跑， 掃羅 和他兒子都死了，就棄城逃跑。 非利士 人前來，佔據了他們的城。
1CHR|10|8|次日， 非利士 人來剝那些被殺之人的衣服，看見 掃羅 和他兒子仆倒在 基利波山 。
1CHR|10|9|他們剝了他的軍裝，拿著他的首級和盔甲，派人到 非利士 人之地的四境，報信給他們的偶像和百姓。
1CHR|10|10|他們將 掃羅 的盔甲放在他們神明的廟裏，把他的首級釘在 大袞 廟中。
1CHR|10|11|基列 的 雅比 居民聽見 非利士 人向 掃羅 所行的一切事，
1CHR|10|12|他們中間所有的勇士就起身，把 掃羅 和他兒子的屍身送到 雅比 ，把他們的屍骨葬在 雅比 的橡樹下，禁食七日。
1CHR|10|13|這樣， 掃羅 為了他的不忠死了；因為他干犯耶和華，沒有遵守耶和華的話，又因他求問招魂的婦人，
1CHR|10|14|不求問耶和華，所以耶和華使他被殺，把王國給了 耶西 的兒子 大衛 。
1CHR|11|1|以色列 眾人聚集到 希伯崙 見 大衛 ，說：「看哪，我們是你的骨肉。
1CHR|11|2|從前 掃羅 作王的時候，率領 以色列 人出入的是你；耶和華－你的上帝也曾對你說：『你必牧養我的百姓 以色列 ，你必作我百姓 以色列 的君王。』」
1CHR|11|3|於是 以色列 的眾長老都來到 希伯崙 見王。 大衛 在 希伯崙 ，在耶和華面前與他們立約，他們就膏 大衛 作 以色列 的王，正如耶和華藉 撒母耳 所說的話。
1CHR|11|4|大衛 和 以色列 眾人到了 耶路撒冷 ，就是 耶布斯 ；那時 耶布斯 人住在那裏。
1CHR|11|5|耶布斯 人對 大衛 說：「你必不能進到這裏。」然而 大衛 攻取了 錫安 的堡壘，就是 大衛 的城。
1CHR|11|6|大衛 說：「誰先攻打 耶布斯 人，必作領袖，作元帥。」 洗魯雅 的兒子 約押 先上去，就作了領袖。
1CHR|11|7|大衛 住在堡壘裏，所以那堡壘叫作 大衛城 。
1CHR|11|8|大衛 又從 米羅 起，四圍建築城牆，其餘的由 約押 修建。
1CHR|11|9|大衛 日見強大，萬軍之耶和華與他同在。
1CHR|11|10|以下是跟隨 大衛 勇士的領袖；他們奮勇幫助他得到國度，並照著耶和華吩咐 以色列 的話，與 以色列 眾人一同立他作王。
1CHR|11|11|大衛 勇士的名單如下： 哈革摩尼 的兒子 雅朔班 ，他是軍官的統領 ，曾一次舉槍殺了三百人。
1CHR|11|12|其次是 亞何亞 人 朵多 的兒子 以利亞撒 ，他是三個勇士裏的一個。
1CHR|11|13|他從前與 大衛 在 巴斯‧大憫 ， 非利士 人聚集要打仗。那裏有一塊長滿大麥的田。百姓在 非利士 人面前逃跑，
1CHR|11|14|他們 卻站在那塊田的中間，防守那田，擊敗了 非利士 人。耶和華大獲全勝。
1CHR|11|15|三十個領袖中的三個人下到磐石那裏，進了 亞杜蘭洞 見 大衛 ； 非利士 的軍隊在 利乏音谷 安營。
1CHR|11|16|那時 大衛 在山寨， 非利士 人的駐軍在 伯利恆 。
1CHR|11|17|大衛 渴想著說：「但願有人從 伯利恆 城門旁的井裏打水來給我喝！」
1CHR|11|18|這三個勇士就闖過 非利士 人的軍營，從 伯利恆 城門旁的井裏打水，拿來給 大衛 喝。 大衛 卻不肯喝，將水澆在耶和華面前，
1CHR|11|19|說：「我的上帝啊，我絕不做這事！這些人冒死去打水，這水是他們用生命換來的，我怎能喝他們的血呢？」 大衛 不肯喝這水。這是三個勇士所做的事。
1CHR|11|20|約押 的兄弟 亞比篩 是這三個 勇士的領袖；他曾舉槍殺了三百人，就在三個勇士中得了名。
1CHR|11|21|他在這三個勇士裏比其他兩個更有名望，所以作他們的領袖，只是不及前三個勇士。
1CHR|11|22|耶何耶大 的兒子 比拿雅 是來自 甲薛 的勇士，曾行了大事。他殺了 摩押 人 亞利伊勒 的兩個兒子，又在下雪的時候下到坑裏去，殺了一隻獅子。
1CHR|11|23|他又殺了一個身高五肘的 埃及 人； 埃及 人手裏拿著槍，槍桿粗如織布機的軸。 比拿雅 只拿著棍子下到他那裏去，從 埃及 人手裏奪過槍來，用那槍殺死了他。
1CHR|11|24|這些是 耶何耶大 的兒子 比拿雅 所做的事，就在三個勇士裏得了名。
1CHR|11|25|看哪，他比那三十個勇士更有名望，只是不及前三個勇士。 大衛 立他作護衛長。
1CHR|11|26|軍中的勇士有 約押 的兄弟 亞撒黑 ， 伯利恆 人 朵多 的兒子 伊勒哈難 ，
1CHR|11|27|哈律 人 沙瑪 ， 比倫 人 希利斯 ，
1CHR|11|28|提哥亞 人 益吉 的兒子 以拉 ， 亞拿突 人 亞比以謝 ，
1CHR|11|29|戶沙 人 西比該 ， 亞何亞 人 以來 ，
1CHR|11|30|尼陀法 人 瑪哈萊 ， 尼陀法 人 巴拿 的兒子 希立 ，
1CHR|11|31|便雅憫 族 基比亞 人 利拜 的兒子 以太 ， 比拉頓 人 比拿雅 ，
1CHR|11|32|迦實溪 人 戶萊 ， 亞拉巴 人 亞比 ，
1CHR|11|33|巴路米 人 押斯瑪弗 ， 沙本 人 以利雅哈巴 ，
1CHR|11|34|基孫 人 哈深 的眾兒子， 哈拉 人 沙基 的兒子 約拿單 ，
1CHR|11|35|哈拉 人 沙甲 的兒子 亞希暗 ， 吾珥 的兒子 以利法勒 ，
1CHR|11|36|米基拉 人 希弗 ， 比倫 人 亞希雅 ，
1CHR|11|37|迦密 人 希斯羅 ， 伊斯拜 的兒子 拿萊 ，
1CHR|11|38|拿單 的兄弟 約珥 ， 哈基利 的兒子 彌伯哈 ，
1CHR|11|39|亞捫 人 洗勒 ， 比錄 人 拿哈萊 ，他是給 洗魯雅 的兒子 約押 拿兵器的，
1CHR|11|40|以帖 人 以拉 ， 以帖 人 迦立 ，
1CHR|11|41|赫 人 烏利亞 ， 亞萊 的兒子 撒拔 ，
1CHR|11|42|呂便 人 示撒 的兒子 亞第拿 ，是 呂便 支派中的一個領袖，率領三十人，
1CHR|11|43|瑪迦 的兒子 哈難 ， 彌特尼 人 約沙法 ，
1CHR|11|44|亞施他拉 人 烏西亞 ， 亞羅珥 人 何坦 的兒子 沙瑪 和 耶利 ，
1CHR|11|45|提洗 人 申利 的兒子 耶疊 和他的兄弟 約哈 ，
1CHR|11|46|瑪哈未 人 以利業 ， 伊利拿安 的兒子 耶利拜 和 約沙未雅 ， 摩押 人 伊特瑪 、
1CHR|11|47|以利業 、 俄備得 ，以及 米瑣八 人 雅西業 。
1CHR|12|1|以下是 大衛 因 基士 的兒子 掃羅 的緣故被放逐到 洗革拉 的時候，到他那裏幫助他打仗的勇士；
1CHR|12|2|他們是弓箭手，能左右甩石，開弓射箭，都是 便雅憫 人 掃羅 同族的弟兄：
1CHR|12|3|為首的是 亞希以謝 ，其次是 約阿施 ，都是 基比亞 人 示瑪 的兒子。還有 亞斯瑪威 的兒子 耶薛 和 毗力 ， 比拉迦 ， 亞拿突 人 耶戶 ，
1CHR|12|4|基遍 人 以實買雅 ，他在三十人中是勇士，管理這三十人，又有 耶利米 ， 雅哈悉 ， 約哈難 ， 基底拉 人 約撒拔 ，
1CHR|12|5|伊利烏賽 ， 耶利末 ， 比亞利雅 ， 示瑪利雅 ， 哈律弗 人 示法提雅 ，
1CHR|12|6|可拉 人 以利加拿 、 耶西亞 、 亞薩列 、 約以謝 、 雅朔班 ，
1CHR|12|7|基多 人 耶羅罕 的兒子 猶拉 和 西巴第雅 。
1CHR|12|8|迦得 人中有人到曠野的山寨投奔 大衛 ，都是大能的勇士，能拿盾牌和槍的戰士。他們的面貌好像獅子，敏捷如山上的鹿。
1CHR|12|9|第一 以薛 ，第二 俄巴底雅 ，第三 以利押 ，
1CHR|12|10|第四 彌施瑪拿 ，第五 耶利米 ，
1CHR|12|11|第六 亞太 ，第七 以利業 ，
1CHR|12|12|第八 約哈難 ，第九 以利薩巴 ，
1CHR|12|13|第十 耶利米 ，第十一 末巴奈 。
1CHR|12|14|這些都是 迦得 人中的軍官，小的能抵一百人，大的能抵一千人 。
1CHR|12|15|正月， 約旦河 水漲過兩岸的時候，他們過河，使所有住河谷的人東奔西逃。
1CHR|12|16|便雅憫 人和 猶大 人中有人來到山寨 大衛 那裏。
1CHR|12|17|大衛 出去迎接他們，回答他們說：「你們若和平地來幫助我，我的心就與你們契合；但你們若把我這雙手無辜的人賣給敵人，願我們列祖的上帝察看責罰。」
1CHR|12|18|那時軍官 的領袖 亞瑪撒 受靈的感動說： 「 大衛 啊，我們歸向你！ 耶西 的兒子啊，我們幫助你！ 願你平平安安， 願幫助你的也都平安！ 因為你的上帝幫助你。」 大衛 就收留他們，派他們作軍官。
1CHR|12|19|大衛 從前與 非利士 人同去，要與 掃羅 爭戰，有些 瑪拿西 人來投奔 大衛 。其實他們並沒有幫助 非利士 人，因為 非利士 人的領袖商議，打發他回去，說：「恐怕 大衛 拿我們的首級去向他的主人 掃羅 投誠。」
1CHR|12|20|大衛 往 洗革拉 去的時候，有 瑪拿西 人的千夫長 押拿 、 約撒拔 、 耶疊 、 米迦勒 、 約撒拔 、 以利戶 、 洗勒太 都來投奔他。
1CHR|12|21|他們幫助 大衛 攻擊敵軍；因為他們都是大能的勇士，又作軍官。
1CHR|12|22|那時天天有人來幫助 大衛 ，以致成了強大的軍隊，如上帝的軍隊一樣。
1CHR|12|23|以下是來到 希伯崙 見 大衛 ，要照耶和華的話把 掃羅 的國位歸給 大衛 的武裝士兵的數目：
1CHR|12|24|猶大 人，拿盾牌和槍的武裝戰士有六千八百人。
1CHR|12|25|西緬 人中，能上陣的大能勇士有七千一百人。
1CHR|12|26|利未 人中，有四千六百人。
1CHR|12|27|耶何耶大 是 亞倫 家的領袖，跟從他的有三千七百人。
1CHR|12|28|還有大能的青年勇士 撒督 ，同他本族的二十二個軍官。
1CHR|12|29|便雅憫 人中， 掃羅 同族的弟兄也有三千人；直到現在他們大部分仍然效忠 掃羅 家。
1CHR|12|30|以法蓮 人中，在本族中著名的大能勇士有二萬零八百人。
1CHR|12|31|瑪拿西 半支派，冊上有名來擁立 大衛 作王的，有一萬八千人。
1CHR|12|32|以薩迦 人中，通達時務，知道 以色列 所當行，同族弟兄也都聽從他們命令的族長有二百人。
1CHR|12|33|西布倫 中，能上陣用各樣作戰的兵器、不生二心幫助打仗的有五萬人。
1CHR|12|34|拿弗他利 中，有一千個軍官；跟從他們、拿盾牌和槍的有三萬七千人。
1CHR|12|35|但 人中，能擺陣的有二萬八千六百人。
1CHR|12|36|亞設 中，能上陣打仗的有四萬人。
1CHR|12|37|約旦河 東的 呂便 人、 迦得 人、 瑪拿西 半支派，拿各樣兵器打仗的有十二萬人。
1CHR|12|38|以上都是能列隊上陣的戰士，他們都全心來到 希伯崙 ，要擁立 大衛 作全 以色列 的王。 以色列 其餘的人也都一心要擁立 大衛 作王。
1CHR|12|39|他們在那裏三日，與 大衛 一同吃喝，因為他們同族的弟兄已經為他們預備好了。
1CHR|12|40|他們附近的人，以及 以薩迦 、 西布倫 、 拿弗他利 人，都將食物，許多麵餅、無花果餅、乾葡萄、酒、油，用驢、駱駝、騾子、牛馱來，又帶了許多的牛和羊來，因為在 以色列 中充滿了歡樂。
1CHR|13|1|大衛 與千夫長、百夫長，以及所有的領袖商議。
1CHR|13|2|大衛 對 以色列 全會眾說：「你們若以為好，見這事是出於耶和華－我們的上帝，我們就派人到遠近各處去見仍留在 以色列 各地我們的弟兄，以及住在有郊野之城的祭司和 利未 人，使他們都到我們這裏來聚集。
1CHR|13|3|我們要把上帝的約櫃接到這裏來；因為在 掃羅 年間，我們沒有去尋求約櫃 。」
1CHR|13|4|全會眾都說可以這麼做，因這事在眾百姓眼中都看為好。
1CHR|13|5|於是， 大衛 把 以色列 眾人從 埃及 的 西曷河 直到 哈馬口 都召集了來，要從 基列‧耶琳 將上帝的約櫃接來。
1CHR|13|6|大衛 率領 以色列 眾人上到 巴拉 ，就是屬 猶大 的 基列‧耶琳 ，要將耶和華上帝的約櫃從那裏接上來，他坐在二基路伯之上，這約櫃是以他的名來命名的。
1CHR|13|7|他們將上帝的約櫃從 亞比拿達 的家裏抬出來，放在新車上，由 烏撒 和 亞希約 趕車。
1CHR|13|8|大衛 和 以色列 眾人在上帝面前隨著詩歌、琴、瑟、鼓、鈸、號，極力跳舞。
1CHR|13|9|到了 基頓 的禾場，因為牛失前蹄 ， 烏撒 就伸手扶住約櫃。
1CHR|13|10|耶和華的怒氣向 烏撒 發作，因他伸手扶住約櫃而擊殺他，他就死在那裏，在上帝面前。
1CHR|13|11|大衛 因耶和華突然衝出撞死 烏撒 就生氣，稱那地方為 毗列斯‧烏撒 ，直到今日。
1CHR|13|12|那日， 大衛 懼怕上帝，說：「我怎能將上帝的約櫃接到我這裏來呢？」
1CHR|13|13|於是 大衛 不將約櫃接進 大衛城 他自己的地方，卻轉送到 迦特 人 俄別‧以東 的家中。
1CHR|13|14|上帝的約櫃停在 俄別‧以東 家中三個月，耶和華賜福給 俄別‧以東 的家和他一切所有的。
1CHR|14|1|推羅 王 希蘭 派使者把香柏木運到 大衛 那裏，又派石匠和木匠給 大衛 建造宮殿。
1CHR|14|2|大衛 知道耶和華堅立他作 以色列 王，又為自己百姓 以色列 的緣故，使他的國興盛。
1CHR|14|3|大衛 在 耶路撒冷 又立后妃，又生兒女。
1CHR|14|4|在 耶路撒冷 所生的孩子名字是 沙母亞 、 朔罷 、 拿單 、 所羅門 、
1CHR|14|5|益轄 、 以利書亞 、 以法列 、
1CHR|14|6|挪迦 、 尼斐 、 雅非亞 、
1CHR|14|7|以利沙瑪 、 比利雅大 、 以利法列 。
1CHR|14|8|非利士 人聽見 大衛 受膏作全 以色列 的王， 非利士 眾人就上來尋索 大衛 。 大衛 聽見了，就出去迎敵。
1CHR|14|9|非利士 人來了，侵犯 利乏音谷 。
1CHR|14|10|大衛 求問上帝說：「我可以上去攻打 非利士 人嗎？你將他們交在我手裏嗎？」耶和華對他說：「你可以上去，我必將他們交在你手裏。」
1CHR|14|11|非利士 人上到 巴力‧毗拉心 ， 大衛 在那裏擊敗他們。 大衛 說：「上帝藉我的手沖破敵人，如水沖破一樣。」因此那地方稱為 巴力‧毗拉心 。
1CHR|14|12|非利士 人把神像拋棄在那裏， 大衛 吩咐人用火焚燒了。
1CHR|14|13|非利士 人又侵犯 利乏音谷 。
1CHR|14|14|大衛 再求問上帝。上帝對他說：「不要從他們後頭追上去，要繞道離開他們，從桑樹林對面攻打他們。
1CHR|14|15|你聽見桑樹梢上有腳步的聲音，那時你就要出戰，因為上帝已經出去，在你前頭攻打 非利士 人的軍隊了。」
1CHR|14|16|大衛 就遵照上帝所吩咐的去做，攻打 非利士 人的軍隊，從 基遍 直到 基色 。
1CHR|14|17|於是 大衛 的名傳揚到萬邦，耶和華使萬國都懼怕他。
1CHR|15|1|大衛 在 大衛城 為自己建造宮殿，又為上帝的約櫃預備地方，支搭帳幕。
1CHR|15|2|那時 大衛 說：「除了 利未 人之外，無人可抬上帝的約櫃，因為耶和華揀選他們抬上帝的約櫃，永遠事奉他。」
1CHR|15|3|大衛 召集 以色列 眾人到 耶路撒冷 ，要將耶和華的約櫃接到他所預備的地方。
1CHR|15|4|大衛 又召集 亞倫 的子孫和 利未 人：
1CHR|15|5|哥轄 子孫中有領袖 烏列 和他的弟兄一百二十人，
1CHR|15|6|米拉利 子孫中有領袖 亞帥雅 和他的弟兄二百二十人，
1CHR|15|7|革順 子孫中有領袖 約珥 和他的弟兄一百三十人，
1CHR|15|8|以利撒反 子孫中有領袖 示瑪雅 和他的弟兄二百人，
1CHR|15|9|希伯倫 子孫中有領袖 以利業 和他的弟兄八十人，
1CHR|15|10|烏薛 子孫中有領袖 亞米拿達 和他的弟兄一百一十二人。
1CHR|15|11|大衛 召來 撒督 和 亞比亞他 二位祭司，以及 利未 人 烏列 、 亞帥雅 、 約珥 、 示瑪雅 、 以利業 、 亞米拿達 ，
1CHR|15|12|對他們說：「你們是 利未 人的族長，你們和你們的弟兄應當使自己分別為聖，好將耶和華－ 以色列 上帝的約櫃接到我所預備的地方。
1CHR|15|13|因為你們上一次沒有抬這約櫃，並且我們沒有按規矩求問耶和華－我們的上帝，所以他衝出來攻擊我們。」
1CHR|15|14|於是祭司和 利未 人使自己分別為聖，將耶和華－ 以色列 上帝的約櫃接上來。
1CHR|15|15|利未 子孫用槓，把上帝的約櫃抬在肩上，正如 摩西 按照耶和華的話所吩咐的。
1CHR|15|16|大衛 吩咐 利未 人的領袖派他們歌唱的弟兄用琴瑟和鈸的樂器奏樂，歡歡喜喜地大聲歌頌。
1CHR|15|17|於是 利未 人派 約珥 的兒子 希幔 和他弟兄中 比利家 的兒子 亞薩 ，以及他們同族弟兄 米拉利 子孫裏 古沙雅 的兒子 以探 。
1CHR|15|18|其次還有跟隨他們的弟兄 撒迦利雅 、 便‧雅薛 、 示米拉末 、 耶歇 、 烏尼 、 以利押 、 比拿雅 、 瑪西雅 、 瑪他提雅 、 以利斐利戶 、 彌克尼雅 ，以及門口的守衛 俄別‧以東 和 耶利 。
1CHR|15|19|歌唱的 希幔 、 亞薩 和 以探 ，敲銅鈸，聲音響亮；
1CHR|15|20|撒迦利雅 、 雅薛 、 示米拉末 、 耶歇 、 烏尼 、 以利押 、 瑪西雅 、 比拿雅 鼓瑟，調用女音；
1CHR|15|21|瑪他提雅 、 以利斐利戶 、 彌克尼雅 、 俄別‧以東 、 耶利 、 亞撒西雅 用琴指揮，調用第八。
1CHR|15|22|基拿尼雅 是 利未 人聖詠團的領袖，又教導人唱歌，因為他精通此事。
1CHR|15|23|比利家 和 以利加拿 是約櫃的守衛。
1CHR|15|24|示巴尼 、 約沙法 、 拿坦業 、 亞瑪賽 、 撒迦利雅 、 比拿亞 、 以利以謝 眾祭司在上帝的約櫃前吹號。 俄別‧以東 和 耶希亞 也是約櫃的守衛。
1CHR|15|25|於是， 大衛 和 以色列 的長老，以及千夫長都去，歡歡喜喜地將耶和華的約櫃從 俄別‧以東 家中接上來。
1CHR|15|26|上帝賜恩給抬耶和華約櫃的 利未 人，他們就獻上七頭公牛，七隻公羊。
1CHR|15|27|大衛 和所有抬約櫃的 利未 人，以及聖詠團的領袖 基拿尼雅 和歌唱的人，都穿著細麻布外袍； 大衛 另外穿著細麻布以弗得。
1CHR|15|28|這樣， 以色列 眾人歡呼、吹角、吹號、敲鈸、鼓瑟、彈琴，聲音響亮，將耶和華的約櫃接上來。
1CHR|15|29|耶和華的約櫃進 大衛城 的時候， 掃羅 的女兒 米甲 從窗戶裏往外觀看，見 大衛 王踴躍跳舞，心裏就輕視他。
1CHR|16|1|眾人將上帝的約櫃請進去，安放在 大衛 為它搭的帳幕中，就在上帝面前獻燔祭和平安祭。
1CHR|16|2|大衛 獻完了燔祭和平安祭，就奉耶和華的名祝福百姓，
1CHR|16|3|並且分給每一個 以色列 人，無論男女，每人一個餅，一個棗子餅 ，一個葡萄餅。
1CHR|16|4|大衛 派幾個 利未 人在耶和華的約櫃前事奉，頌揚，稱謝，讚美耶和華－ 以色列 的上帝：
1CHR|16|5|為首的是 亞薩 ，其次是 撒迦利雅 、 耶利 、 示米拉末 、 耶歇 、 瑪他提雅 、 以利押 、 比拿雅 、 俄別‧以東 、 耶利 ；他們鼓瑟彈琴， 亞薩 敲鈸，聲音響亮；
1CHR|16|6|比拿雅 和 雅哈悉 二位祭司常在上帝的約櫃前吹號。
1CHR|16|7|那日， 大衛 初次指派 亞薩 和他的弟兄稱謝耶和華。
1CHR|16|8|你們要稱謝耶和華，求告他的名， 在萬民中傳揚他的作為！
1CHR|16|9|要向他唱詩，向他歌頌， 述說他一切奇妙的作為！
1CHR|16|10|要誇耀他的聖名！ 願尋求耶和華的人心中歡喜！
1CHR|16|11|要尋求耶和華與他的能力， 時常尋求他的面。
1CHR|16|12|他僕人 以色列 的後裔， 他所揀選 雅各 的子孫哪， 要記念他奇妙的作為和他的奇事， 並他口中的判語。
1CHR|16|13|
1CHR|16|14|他是耶和華－我們的上帝， 全地都有他的判斷。
1CHR|16|15|要記念他的約，直到永遠； 記念他吩咐的話，直到千代，
1CHR|16|16|就是他與 亞伯拉罕 所立的約， 向 以撒 所起的誓。
1CHR|16|17|他將這約向 雅各 定為律例， 向 以色列 定為永遠的約，
1CHR|16|18|說：「我必將 迦南 地賜給你， 作你們應得的產業。」
1CHR|16|19|當時，你們人丁有限， 數目稀少，在那地寄居。
1CHR|16|20|他們從這邦遊到那邦， 從這國去到另一民族。
1CHR|16|21|他不容人欺負他們， 為他們的緣故責備君王：
1CHR|16|22|「不可傷害我的受膏者， 也不可惡待我的先知。」
1CHR|16|23|全地都要向耶和華歌唱！ 天天傳揚他的救恩！
1CHR|16|24|在列國中述說他的榮耀！ 在萬民中述說他的奇事！
1CHR|16|25|因耶和華本為大，當受極大的讚美； 他在萬神之上，當受敬畏。
1CHR|16|26|因萬民的神明都屬虛無； 惟獨耶和華創造諸天。
1CHR|16|27|有尊榮和威嚴在他面前， 有能力和喜樂在他自己的地方。
1CHR|16|28|民中的萬族啊，要將榮耀、能力歸給耶和華， 都歸給耶和華！
1CHR|16|29|要將耶和華的名所當得的榮耀歸給他， 拿供物來獻在他面前； 當敬拜神聖榮耀的耶和華 。
1CHR|16|30|全地都要在他面前戰抖！ 世界堅定，不得動搖。
1CHR|16|31|願天歡喜，願地快樂！ 願人在列國中說： 「耶和華作王了！」
1CHR|16|32|願海和其中所充滿的澎湃！ 願田和其中所有的都歡樂！
1CHR|16|33|那時，林中的樹木都要在耶和華面前歡呼， 因為他來要審判全地。
1CHR|16|34|你們要稱謝耶和華，因他本為善， 他的慈愛永遠長存！
1CHR|16|35|你們要說： 「拯救我們的上帝啊，求你拯救我們， 聚集我們，救我們脫離列國， 我們好頌揚你的聖名， 以讚美你為誇勝。
1CHR|16|36|耶和華－ 以色列 的上帝是應當稱頌的， 從亙古直到永遠。」 全體百姓都說：「阿們！」並且讚美耶和華。
1CHR|16|37|大衛 把 亞薩 和他的弟兄留在耶和華的約櫃那裏，經常在約櫃前事奉，天天盡本分供職，
1CHR|16|38|又有 俄別‧以東 和他的弟兄六十八人； 耶杜頓 的兒子 俄別‧以東 ，以及 何薩 作門口的守衛。
1CHR|16|39|還有 撒督 祭司和他弟兄眾祭司在 基遍 的丘壇、耶和華的帳幕前，
1CHR|16|40|在燔祭壇上，每日早晚，照著寫在耶和華律法書上所吩咐 以色列 的，經常獻燔祭給耶和華。
1CHR|16|41|與他們一同的還有 希幔 、 耶杜頓 ，和其餘被選、名字錄在冊上的，為要稱謝耶和華，因他的慈愛永遠長存。
1CHR|16|42|希幔 、 耶杜頓 同他們吹號、敲鈸，聲音響亮，並用其他樂器配合，歌頌上帝。 耶杜頓 的子孫作門口的守衛。
1CHR|16|43|於是眾百姓各自回家， 大衛 也回去為家人祝福。
1CHR|17|1|大衛 住在自己宮中，對 拿單 先知說：「看哪，我住在香柏木的宮中，耶和華的約櫃卻在幔子裏。」
1CHR|17|2|拿單 對 大衛 說：「你可以完全照你的心意去做，因為上帝與你同在。」
1CHR|17|3|當夜上帝的話臨到 拿單 ，說：
1CHR|17|4|「你去對我僕人 大衛 說：『耶和華如此說：你不可建造殿宇給我居住。
1CHR|17|5|自從我領 以色列 人上來，直到今日，我未曾住過殿宇；我從這會幕到那會幕，從這帳幕到那帳幕 。
1CHR|17|6|凡我同 以色列 人所走的地方，我何曾向 以色列 的一個士師，就是我吩咐牧養我百姓的，說過這話：你們為何不給我建造香柏木的殿宇呢？』
1CHR|17|7|現在，你要對我僕人 大衛 這樣說：『萬軍之耶和華如此說：我從羊圈中將你召來，叫你不再牧放羊群，立你作我百姓 以色列 的君王。
1CHR|17|8|你無論往哪裏去，我都與你同在，剪除你所有的仇敵。我必使你得大名，好像世上偉人的名一樣。
1CHR|17|9|我必為我百姓 以色列 選定一個地方，栽植他們，使他們住自己的地方，不再受攪擾；兇惡之子也不再像從前那樣擾亂他們，
1CHR|17|10|並不像我命令士師治理我百姓 以色列 的日子。我必制伏你所有的仇敵，並且我應許你 ，耶和華必為你建立家室。
1CHR|17|11|當你壽數滿足歸你祖先的時候，我必使你的後裔，你自己的兒子接續你；我也必堅定他的國。
1CHR|17|12|他必為我建造殿宇，我必堅定他的王位，直到永遠。
1CHR|17|13|我要作他的父，他要作我的子；我必不使我的慈愛離開他，像離開在你以前的那位一樣。
1CHR|17|14|我要永遠堅立他在我的家和我的國裏；他的王位也必堅定，直到永遠。』」
1CHR|17|15|拿單 就按這一切話，照這一切異象告訴 大衛 。
1CHR|17|16|於是 大衛 王進去，坐在耶和華面前，說：「耶和華上帝啊，我是誰，我的家算甚麼，你竟帶領我到這地步呢？
1CHR|17|17|上帝啊，這在你眼中還看為小，你又說到你僕人的家將來的情況。耶和華上帝啊，你看顧我好像看顧尊貴的人。
1CHR|17|18|你加於僕人的尊榮， 大衛 還有甚麼可以對你說呢？你是知道你僕人的。
1CHR|17|19|耶和華啊，因你僕人的緣故，也照著你的心意，你行這一切大事，為了顯明這一切偉大的事。
1CHR|17|20|耶和華啊，照我們耳中一切所聽見的，沒有可比你的，除你以外再沒有上帝。
1CHR|17|21|世上有何國能比你的百姓 以色列 呢？上帝親自去救贖世上的一國 ，作自己的子民，又行大而可畏的事，顯出你的大名，在你從 埃及 贖出來的子民面前驅逐了列國。
1CHR|17|22|你使你的百姓 以色列 作你的子民，直到永遠；你－耶和華也作他們的上帝。
1CHR|17|23|現在，耶和華啊，你所應許僕人和僕人家的話，求你堅定，直到永遠；求你照你所說的而行。
1CHR|17|24|願你的名永遠堅立，被尊為大，人要說：『萬軍之耶和華－ 以色列 的上帝，是 以色列 的上帝。』這樣，你僕人 大衛 的家必在你面前堅立。
1CHR|17|25|我的上帝啊，因你啟示你的僕人，要為他建立家室，所以僕人大膽在你面前祈禱。
1CHR|17|26|現在，耶和華啊，惟有你是上帝！你應許將這福氣賜給僕人。
1CHR|17|27|現在，你喜悅賜福給僕人的家，可以永存在你面前。耶和華啊，因你已經賜福，還要賜福到永遠。」
1CHR|18|1|此後， 大衛 攻打 非利士 人，制伏了他們，從 非利士 人手中奪取了 迦特 和所屬的鄉鎮。
1CHR|18|2|他又攻打 摩押 ， 摩押 人就臣服 大衛 ，向他進貢。
1CHR|18|3|瑣巴 王 哈大底謝 往 幼發拉底河 去，要鞏固自己的國權。 大衛 攻打他，直到 哈馬 ，
1CHR|18|4|奪了他的戰車一千，俘擄了騎兵七千人，步兵二萬人。 大衛 把所有戰馬的蹄筋砍斷，只留下一百輛戰車。
1CHR|18|5|大馬士革 的 亞蘭 人來幫助 瑣巴 王 哈大底謝 ， 大衛 殺了 亞蘭 人二萬二千。
1CHR|18|6|於是 大衛 在 大馬士革 的 亞蘭 地設立軍營 ， 亞蘭 人就臣服 大衛 ，向他進貢。 大衛 無論往哪裏去，耶和華都使他得勝。
1CHR|18|7|大衛 奪了 哈大底謝 臣僕擁有的金盾牌，帶到 耶路撒冷 。
1CHR|18|8|大衛 又從 哈大底謝 的 提巴 和 均 二城奪取了許多的銅；後來 所羅門 用這些銅製造銅海、銅柱和銅器。
1CHR|18|9|哈馬 王 陀烏 聽見 大衛 擊敗 瑣巴 王 哈大底謝 的全軍，
1CHR|18|10|就派他兒子 哈多蘭 到 大衛 王那裏，向他請安，為他祝福，因他與 哈大底謝 爭戰，並且擊敗了他；原來 哈大底謝 與 陀烏 常常爭戰。 哈多蘭 帶了金銀銅的各樣器皿來。
1CHR|18|11|大衛 王把這些器皿，以及從各國奪來的金銀，就是從 以東 、 摩押 、 亞捫 人、 非利士 人、 亞瑪力 所奪來的，都分別為聖獻給耶和華。
1CHR|18|12|洗魯雅 的兒子 亞比篩 在 鹽谷 擊殺了一萬八千 以東 人。
1CHR|18|13|大衛 在 以東 設立軍營， 以東 人就都臣服他。 大衛 無論往哪裏去，耶和華都使他得勝。
1CHR|18|14|大衛 作全 以色列 的王，又向眾百姓秉公行義。
1CHR|18|15|洗魯雅 的兒子 約押 作元帥； 亞希律 的兒子 約沙法 作史官；
1CHR|18|16|亞希突 的兒子 撒督 和 亞比亞他 的兒子 亞希米勒 作祭司； 沙威沙 作書記；
1CHR|18|17|耶何耶大 的兒子 比拿雅 管轄 基利提 人和 比利提 人。 大衛 的眾兒子都在王的左右作領袖。
1CHR|19|1|此後， 亞捫 人的王 拿轄 死了，他兒子接續他作王。
1CHR|19|2|大衛 說：「 哈嫩 的父親 拿轄 怎樣向我施恩，我也要怎樣向 哈嫩 施恩。」於是 大衛 派使者為他的父親安慰他。 大衛 的臣僕到了 亞捫 人的境內來見 哈嫩 ，要安慰他。
1CHR|19|3|但 亞捫 人的領袖對 哈嫩 說：「 大衛 派人來安慰你，你看他是要尊敬你父親嗎？他的臣僕來見你，不是為了要窺探偵察，而傾覆這地嗎？」
1CHR|19|4|哈嫩 就抓住 大衛 的臣僕，剃去他們的鬍鬚，又割斷他們下半截的衣服，露出臀部，然後放了他們。
1CHR|19|5|他們走了，有人把臣僕所遭遇的事告訴 大衛 ，他就派人去迎接他們，因為這些人覺得很羞恥。王說：「可以住在 耶利哥 ，等到鬍鬚長出來再回來。」
1CHR|19|6|亞捫 人看到 大衛 憎惡他們， 哈嫩 和 亞捫 人就派人拿一千他連得銀子，從 美索不達米亞 、 亞蘭‧瑪迦 、 瑣巴 雇用戰車和騎兵。
1CHR|19|7|他們雇了三萬二千輛戰車，以及 瑪迦 王和他的軍兵；這些部隊來安營在 米底巴 前。 亞捫 人也從他們的城裏出來，聚集預備作戰。
1CHR|19|8|大衛 聽見了，就派 約押 和所有勇猛的軍隊出去。
1CHR|19|9|亞捫 人出來，在城門前擺陣，前來的諸王另在郊野擺陣。
1CHR|19|10|約押 看見戰陣對著他前後擺列，就把從 以色列 所有精兵中挑選出來的，擺陣迎戰 亞蘭 人。
1CHR|19|11|他把其餘的兵交在他兄弟 亞比篩 手裏，他們就擺陣迎戰 亞捫 人。
1CHR|19|12|約押 說：「 亞蘭 人若強過我，你就來幫助我； 亞捫 人若強過你，我就去幫助你。
1CHR|19|13|你要剛強，我們要為自己的百姓，為我們上帝的城鎮奮勇。願耶和華照他所看為好的去做！」
1CHR|19|14|於是， 約押 和跟隨他的士兵前進攻打 亞蘭 人； 亞蘭 人在他面前逃跑。
1CHR|19|15|亞捫 人見 亞蘭 人逃跑，他們也在 約押 的兄弟 亞比篩 面前逃跑進城。 約押 就回 耶路撒冷 去了。
1CHR|19|16|亞蘭 人見自己被 以色列 打敗，就派使者把 大河 那邊的 亞蘭 人調來，由 哈大底謝 的將軍 朔法 在他們前面率領。
1CHR|19|17|有人告訴 大衛 ，他就聚集 以色列 眾人過 約旦河 ，來到 亞蘭 人那裏，迎著他們擺陣。 大衛 擺陣攻擊 亞蘭 人， 亞蘭 人就與他打仗。
1CHR|19|18|亞蘭 人在 以色列 人面前逃跑。 大衛 殺了 亞蘭 七千輛戰車的士兵，四萬步兵，又殺死 亞蘭 的將軍 朔法 。
1CHR|19|19|哈大底謝 的臣僕見自己被 以色列 打敗，就與 大衛 講和，臣服他。於是 亞蘭 人不願再幫助 亞捫 人了。
1CHR|20|1|到了年初，諸王出征的時候， 約押 率領軍兵蹂躪 亞捫 人的地，前來圍攻 拉巴 ； 大衛 仍住在 耶路撒冷 。 約押 攻打 拉巴 ，把它毀壞。
1CHR|20|2|大衛 奪了 米勒公 所戴的冠冕，其上的金子重一他連得，又嵌著寶石。這冠冕就戴在 大衛 頭上。 大衛 又從城裏奪了許多財物，
1CHR|20|3|把城裏的百姓拉出來，放在鋸下，或鐵耙下，或斧 的下面； 大衛 待 亞捫 各城的居民都是如此。於是， 大衛 和全軍都回 耶路撒冷 去了。
1CHR|20|4|後來， 以色列 人在 基色 與 非利士 人打仗。 戶沙 人 西比該 殺了巨人族的後裔 細派 ， 非利士 人就被制伏了。
1CHR|20|5|他們又與 非利士 人打仗。 睚珥 的兒子 伊勒哈難 殺了 迦特 人 歌利亞 的兄弟 拉哈米 ；這人的槍桿粗如織布機的軸。
1CHR|20|6|又有一次，他們在 迦特 打仗。那裏有一個身材高大的人，手指腳趾都是六根，共有二十四根；他也是巨人族的後裔。
1CHR|20|7|他向 以色列 罵陣， 大衛 的哥哥 示米亞 的兒子 約拿單 就殺了他。
1CHR|20|8|這些人是 迦特 巨人族的後裔，都仆倒在 大衛 和他僕人的手下。
1CHR|21|1|撒但起來攻擊 以色列 ，激起 大衛 數點以色列人。
1CHR|21|2|大衛 對 約押 和百姓的領袖說：「去，數點 以色列 人，從 別是巴 直到 但 ，回來告訴我，我好知道他們的數目。」
1CHR|21|3|約押 說：「願耶和華使他的百姓比現在加增百倍。我主我王啊，他們不都是我主的僕人嗎？我主為何吩咐行這事，為何使 以色列 陷入罪裏呢？」
1CHR|21|4|但王堅持他對 約押 的命令。 約押 就出去，來回走遍 以色列 ，然後回到 耶路撒冷 。
1CHR|21|5|約押 向 大衛 報告百姓的總數：全 以色列 拿刀的有一百一十萬人； 猶大 拿刀的有四十七萬人。
1CHR|21|6|惟有 利未 人和 便雅憫 人沒有算在其中，因為 約押 厭惡王的這命令。
1CHR|21|7|這件事在上帝眼中看為惡，上帝就降災給 以色列 。
1CHR|21|8|大衛 對上帝說：「我做這事大大有罪了。現在求你除掉僕人的罪孽，因為我所做的非常愚昧。」
1CHR|21|9|耶和華吩咐 迦得 ， 大衛 的先見，說：
1CHR|21|10|「你去告訴 大衛 說：『耶和華如此說：我列出三樣災禍給你，隨你選擇一樣，我好降與你。』」
1CHR|21|11|於是， 迦得 來到 大衛 那裏，對他說：「耶和華如此說：『你可以隨意選擇：
1CHR|21|12|三年的饑荒，或敗在敵人面前，被敵人的刀追殺三個月，或在國中三日有耶和華的刀，就是瘟疫，讓耶和華的使者在 以色列 全境施行毀滅呢？』現在你要想一想，我怎樣去回覆那差我來的。」
1CHR|21|13|大衛 對 迦得 說：「我很為難。我寧願落在耶和華的手裏，因為他有豐盛的憐憫；我不願落在人的手裏。」
1CHR|21|14|於是，耶和華降瘟疫給 以色列 ， 以色列 中死了七萬人。
1CHR|21|15|上帝派遣使者去毀滅 耶路撒冷 ，剛要毀滅的時候，耶和華看見就改變心意，不降這災了。他吩咐那滅城的天使說：「夠了，住手吧！」耶和華的使者正站在 耶布斯 人 阿珥楠 的禾場那裏。
1CHR|21|16|大衛 舉目，看見耶和華的使者站在天和地之間，手裏有拔出來的刀，伸在 耶路撒冷 以上。 大衛 和長老都披上麻布，臉伏於地。
1CHR|21|17|大衛 向上帝說：「吩咐數點百姓的不是我嗎？是我犯了罪，行了大惡，但這群羊做了甚麼呢？耶和華－我的上帝啊，願你的手攻擊我和我的父家，不要降瘟疫給你的百姓。」
1CHR|21|18|耶和華的使者吩咐 迦得 去告訴 大衛 ，叫他上去，在 耶布斯 人 阿珥楠 的禾場上為耶和華立一座壇。
1CHR|21|19|大衛 就照著 迦得 奉耶和華名所說的話上去。
1CHR|21|20|阿珥楠 回頭看見天使，跟他在一起的四個兒子都藏起來了， 阿珥楠 繼續打麥子。
1CHR|21|21|大衛 到了 阿珥楠 那裏， 阿珥楠 觀看，看見 大衛 ，就從禾場上出去，臉伏於地，向他下拜。
1CHR|21|22|大衛 對 阿珥楠 說：「你把這禾場的地方給我，照著十足的價錢賣給我，我好在其上為耶和華築一座壇，使瘟疫在百姓中停止。」
1CHR|21|23|阿珥楠 對 大衛 說：「請用這禾場吧，願我主我王照你眼中看為好的去做。看，我提供牛作燔祭，打糧的器具作柴，麥子作素祭，這一切我全都提供。」
1CHR|21|24|大衛 王對 阿珥楠 說：「不，我一定要按十足的價錢買；因我不能用你的東西獻給耶和華，也不能用白得之物獻為燔祭。」
1CHR|21|25|於是 大衛 為那個地方付了六百舍客勒重的金子給 阿珥楠 。
1CHR|21|26|大衛 在那裏為耶和華築了一座壇，獻燔祭和平安祭，求告耶和華。耶和華就應允他，使火從天降在燔祭壇上。
1CHR|21|27|耶和華吩咐使者，他就收刀入鞘。
1CHR|21|28|那時， 大衛 見耶和華在 耶布斯 人 阿珥楠 的禾場上應允了他，就在那裏獻祭。
1CHR|21|29|摩西 在曠野所造之耶和華的帳幕和燔祭壇，當時都在 基遍 的丘壇，
1CHR|21|30|只是 大衛 不能前去求問上帝，因為他懼怕耶和華使者的刀。
1CHR|22|1|大衛 說：「這是耶和華上帝的殿，這是 以色列 獻燔祭的壇。」
1CHR|22|2|大衛 吩咐人召集住 以色列 地的寄居者，又派石匠鑿石頭，要建造上帝的殿。
1CHR|22|3|大衛 預備許多鐵，要做門上的釘子和鉤子，又預備許多銅，多得無法可秤；
1CHR|22|4|還有無數的香柏木，因為 西頓 人和 推羅 人給 大衛 運了許多香柏木來。
1CHR|22|5|大衛 說：「我兒子 所羅門 還年幼脆弱，要為耶和華建造的殿宇必須高大輝煌，使名聲榮耀傳遍萬國，所以我要為殿預備。」於是， 大衛 在未死之前預備了許多材料。
1CHR|22|6|大衛 召了他兒子 所羅門 來，吩咐他為耶和華－ 以色列 的上帝建造殿宇。
1CHR|22|7|大衛 對 所羅門 說：「我兒啊，我心裏本想為耶和華－我上帝的名建造殿宇，
1CHR|22|8|可是耶和華的話臨到我說：『你流了許多的血，打了多次大仗；你不可為我的名建造殿宇，因為你在我面前使許多血流在地上。
1CHR|22|9|看哪，你要生一個兒子，他必成為安寧的人；我必使他得享安寧，不被四圍仇敵擾亂。他的名字要叫 所羅門 ，在他的日子，我必使 以色列 平安康泰。
1CHR|22|10|他必為我的名建造殿宇。他要作我的子，我要作他的父。我必堅定他國度的王位，使他治理 以色列 ，直到永遠。』
1CHR|22|11|我兒啊，現今願耶和華與你同在，使你亨通，建造耶和華－你上帝的殿，正如他指著你所說的。
1CHR|22|12|但願耶和華賜你聰明智慧，好按著他吩咐你的去治理 以色列 ，遵行耶和華－你上帝的律法。
1CHR|22|13|那時候，你若謹守遵行耶和華藉 摩西 吩咐 以色列 的律例典章，就得亨通。你當剛強壯膽，不要懼怕，也不要驚惶。
1CHR|22|14|看哪，我辛苦地為耶和華的殿預備了十萬他連得金子，一百萬他連得銀子，銅和鐵多得無法可秤；我也預備了木頭、石頭，你還可以增添。
1CHR|22|15|你有許多工匠，就是石匠、木匠，和一切能做各樣工的巧匠，
1CHR|22|16|以及無數的金銀銅鐵。你當起來做工，願耶和華與你同在。」
1CHR|22|17|大衛 又吩咐 以色列 的眾官長幫助他兒子 所羅門 ：
1CHR|22|18|「耶和華－你們的上帝不是與你們同在嗎？他不是使你們四圍都平安嗎？因他已將這地的居民交在我手中，這地已在耶和華與他百姓面前制伏了。
1CHR|22|19|現在你們應當立定心意，尋求耶和華－你們的上帝。你們當起來建造耶和華上帝的聖所，好將耶和華的約櫃和上帝神聖的器皿都搬進為耶和華的名建造的殿裏。」
1CHR|23|1|大衛 年紀老邁，日子滿足，就立他兒子 所羅門 作 以色列 的王。
1CHR|23|2|大衛 召集 以色列 的眾領袖、祭司和 利未 人。
1CHR|23|3|利未 人三十歲以上的都被數點，他們男丁的數目共有三萬八千；
1CHR|23|4|其中有二萬四千人管理耶和華殿的事務，有六千人作官長和審判官，
1CHR|23|5|有四千人作門口的守衛，又有四千人頌讚耶和華，用 大衛 造的樂器來頌讚。
1CHR|23|6|大衛 把 利未 人 革順 、 哥轄 、 米拉利 的子孫分了班次。
1CHR|23|7|屬 革順 的有 拉但 和 示每 。
1CHR|23|8|拉但 的長子是 耶歇 ，還有 西坦 和 約珥 ，共三人。
1CHR|23|9|示每 的兒子是 示羅密 、 哈薛 、 哈蘭 三人。這是 拉但 族的族長。
1CHR|23|10|示每 的兒子是 雅哈 、 細拿 、 耶烏施 、 比利亞 ，這四人是 示每 的兒子。
1CHR|23|11|雅哈 是長子， 細撒 是次子。但 耶烏施 和 比利亞 的子孫不多，所以算為一族。
1CHR|23|12|哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 、 烏薛 ，共四人。
1CHR|23|13|暗蘭 的兒子是 亞倫 和 摩西 。 亞倫 被分別出來，把至聖之物分別為聖，使他和他的子孫在耶和華面前燒香、事奉他，奉他的名祝福，直到永遠。
1CHR|23|14|至於神人 摩西 ，他的子孫記名在 利未 支派下。
1CHR|23|15|摩西 的兒子是 革舜 和 以利以謝 。
1CHR|23|16|革舜 的兒子，長子是 細布業 ；
1CHR|23|17|以利以謝 的兒子，長子是 利哈比雅 。 以利以謝 沒有別的兒子，但 利哈比雅 的子孫很多。
1CHR|23|18|以斯哈 的兒子，長子是 示羅密 。
1CHR|23|19|希伯倫 的兒子，長子是 耶利雅 ，次子是 亞瑪利亞 ，三子是 雅哈悉 ，四子是 耶加面 。
1CHR|23|20|烏薛 的兒子，長子是 米迦 ，次子是 耶西雅 。
1CHR|23|21|米拉利 的兒子是 抹利 和 母示 。 抹利 的兒子是 以利亞撒 和 基士 。
1CHR|23|22|以利亞撒 死了，沒有兒子，只有女兒，他們本族 基士 的幾個兒子娶了她們為妻。
1CHR|23|23|母示 的兒子是 末力 、 以得 、 耶列末 ，共三人。
1CHR|23|24|以上是 利未 子孫作族長的，按著父系、照著男丁的數目，二十歲以上登記的，都辦理耶和華殿的事務。
1CHR|23|25|大衛 說：「耶和華－ 以色列 的上帝已經使他的百姓得享安寧，他永遠住在 耶路撒冷 。
1CHR|23|26|因此， 利未 人不必再抬帳幕和其中所使用的一切器皿了。」
1CHR|23|27|照著 大衛 臨終的話， 利未 人二十歲以上的都被數點。
1CHR|23|28|他們的職務是作 亞倫 子孫的幫手，在耶和華的殿事奉，照管院子和屋子，潔淨一切聖物，辦理上帝殿的事務。
1CHR|23|29|他們負責預備供餅、素祭的細麵和無酵薄餅，或用盤烤，或用油調和的祭物，確認其數量和大小。
1CHR|23|30|每日早晚、安息日、初一，以及節期，按數照例，經常獻燔祭給耶和華的時候，他們站立稱謝讚美耶和華。
1CHR|23|31|
1CHR|23|32|他們照管會幕和聖所，服事他們的弟兄 亞倫 的子孫，辦理耶和華殿的事務。
1CHR|24|1|亞倫 子孫的班次如下： 亞倫 的兒子是 拿答 、 亞比戶 、 以利亞撒 、 以他瑪 。
1CHR|24|2|拿答 和 亞比戶 死在他們父親之先，沒有留下兒子；因此， 以利亞撒 和 以他瑪 擔任祭司的職分。
1CHR|24|3|大衛 和 以利亞撒 的子孫 撒督 ，以及 以他瑪 的子孫 亞希米勒 ，把他們按照任務分成班次，
1CHR|24|4|發現 以利亞撒 子孫中作領袖的，比 以他瑪 子孫中作領袖的更多，就分班如下： 以利亞撒 的子孫中有十六個族長， 以他瑪 的子孫中有八個族長。
1CHR|24|5|他們抽籤分配，彼此一樣。在聖所和上帝面前作領袖的有 以利亞撒 的子孫，也有 以他瑪 的子孫。
1CHR|24|6|作書記的 利未 人 拿坦業 的兒子 示瑪雅 在王和領袖，與 撒督 祭司、 亞比亞他 的兒子 亞希米勒 ，以及祭司和 利未 人的族長面前記錄他們的名字；在 以利亞撒 的子孫中取一族，在 以他瑪 的子孫中也取一族。
1CHR|24|7|抽籤的時候，第一籤抽到的是 耶何雅立 ，第二是 耶大雅 ，
1CHR|24|8|第三是 哈琳 ，第四是 梭琳 ，
1CHR|24|9|第五是 瑪基雅 ，第六是 米雅民 ，
1CHR|24|10|第七是 哈歌斯 ，第八是 亞比雅 ，
1CHR|24|11|第九是 耶書亞 ，第十是 示迦尼 ，
1CHR|24|12|第十一是 以利亞實 ，第十二是 雅金 ，
1CHR|24|13|第十三是 胡巴 ，第十四是 耶是比押 ，
1CHR|24|14|第十五是 璧迦 ，第十六是 音麥 ，
1CHR|24|15|第十七是 希悉 ，第十八是 哈闢悉 ，
1CHR|24|16|第十九是 毗他希雅 ，第二十是 以西結 ，
1CHR|24|17|第二十一是 雅斤 ，第二十二是 迦末 ，
1CHR|24|18|第二十三是 第來雅 ，第二十四是 瑪西亞 。
1CHR|24|19|這就是他們事奉的班次，要照耶和華－ 以色列 的上帝藉他們祖宗 亞倫 所吩咐的條例，進入耶和華的殿辦理事務。
1CHR|24|20|利未 其餘的子孫如下： 暗蘭 的子孫中有 書巴業 ； 書巴業 的子孫中有 耶希底亞 。
1CHR|24|21|屬 利哈比雅 ， 利哈比雅 的兒子中有長子 伊示雅 。
1CHR|24|22|屬 以斯哈 人的有 示羅摩 ； 示羅摩 的子孫中有 雅哈 。
1CHR|24|23|希伯倫 的兒子中有長子 耶利雅 ，次子 亞瑪利亞 ，三子 雅哈悉 ，四子 耶加面 。
1CHR|24|24|烏薛 的子孫中有 米迦 ； 米迦 的子孫中有 沙密 。
1CHR|24|25|米迦 的兄弟是 伊示雅 ； 伊示雅 的子孫中有 撒迦利雅 。
1CHR|24|26|米拉利 的兒子是 抹利 和 母示 ； 雅西雅 的子孫中有 比挪 ；
1CHR|24|27|米拉利 的子孫中有屬 雅西雅 的 比挪 、 朔含 、 撒刻 、 伊比利 。
1CHR|24|28|屬 抹利 的有 以利亞撒 ； 以利亞撒 沒有兒子。
1CHR|24|29|屬 基士 ， 基士 的子孫中有 耶拉篾 。
1CHR|24|30|母示 的兒子是 末力 、 以得 、 耶利末 。按著宗族，這些都是 利未 的子孫。
1CHR|24|31|他們在 大衛 王和 撒督 ，以及 亞希米勒 與祭司和 利未 人的族長面前也抽籤，正如他們弟兄 亞倫 的子孫一樣。各族的族長與最年輕的兄弟都一樣。
1CHR|25|1|大衛 和事奉團隊的眾領袖分派 亞薩 、 希幔 ，以及 耶杜頓 的子孫唱歌 ，以彈琴、鼓瑟、敲鈸伴奏。他們供職的人數如下：
1CHR|25|2|亞薩 的兒子 撒刻 、 約瑟 、 尼探雅 、 亞薩利拉 ， 亞薩 的兒子都在 亞薩 的指導下，遵王的指示唱歌。
1CHR|25|3|屬 耶杜頓 ， 耶杜頓 的兒子 基大利 、 西利 、 耶篩亞 、 示每 、 哈沙比雅 、 瑪他提雅 共六人，都在他們父親 耶杜頓 的指導下唱歌，以彈琴伴奏，稱謝，頌讚耶和華。
1CHR|25|4|屬 希幔 ， 希幔 的兒子是 布基雅 、 瑪探雅 、 烏薛 、 細布業 、 耶利末 、 哈拿尼雅 、 哈拿尼 、 以利亞他 、 基大利提 、 羅幔提‧以謝 、 約施比加沙 、 瑪羅提 、 何提 、 瑪哈秀 。
1CHR|25|5|這些都是 希幔 的兒子； 希幔 奉上帝之命作王的先見，吹角頌讚。上帝賜給 希幔 十四個兒子，三個女兒，
1CHR|25|6|他們都在父親的指導下，在耶和華的殿唱歌，以敲鈸、彈琴、鼓瑟伴奏，遵從王的指示，在上帝的殿裏事奉。 亞薩 、 耶杜頓 、 希幔 ，
1CHR|25|7|他們和他們的弟兄學習頌讚耶和華，精通者的數目共有二百八十八人。
1CHR|25|8|這些人無論大小，為師的、為徒的，都一同抽籤分了班次。
1CHR|25|9|抽籤的時候，第一籤抽到的是 亞薩 的兒子 約瑟 。第二是 基大利 ；他和他兄弟，以及兒子共十二人。
1CHR|25|10|第三是 撒刻 ，他兒子和他兄弟共十二人。
1CHR|25|11|第四是 伊洗利 ，他兒子和他兄弟共十二人。
1CHR|25|12|第五是 尼探雅 ，他兒子和他兄弟共十二人。
1CHR|25|13|第六是 布基雅 ，他兒子和他兄弟共十二人。
1CHR|25|14|第七是 耶薩利拉 ，他兒子和他兄弟共十二人。
1CHR|25|15|第八是 耶篩亞 ，他兒子和他兄弟共十二人。
1CHR|25|16|第九是 瑪探雅 ，他兒子和他兄弟共十二人。
1CHR|25|17|第十是 示每 ，他兒子和他兄弟共十二人。
1CHR|25|18|第十一是 亞薩烈 ，他兒子和他兄弟共十二人。
1CHR|25|19|第十二是 哈沙比雅 ，他兒子和他兄弟共十二人。
1CHR|25|20|第十三是 書巴業 ，他兒子和他兄弟共十二人。
1CHR|25|21|第十四是 瑪他提雅 ，他兒子和他兄弟共十二人。
1CHR|25|22|第十五是 耶列末 ，他兒子和他兄弟共十二人。
1CHR|25|23|第十六是 哈拿尼雅 ，他兒子和他兄弟共十二人。
1CHR|25|24|第十七是 約施比加沙 ，他兒子和他兄弟共十二人。
1CHR|25|25|第十八是 哈拿尼 ，他兒子和他兄弟共十二人。
1CHR|25|26|第十九是 瑪羅提 ，他兒子和他兄弟共十二人。
1CHR|25|27|第二十是 以利亞他 ，他兒子和他兄弟共十二人。
1CHR|25|28|第二十一是 何提 ，他兒子和他兄弟共十二人。
1CHR|25|29|第二十二是 基大利提 ，他兒子和他兄弟共十二人。
1CHR|25|30|第二十三是 瑪哈秀 ，他兒子和他兄弟共十二人。
1CHR|25|31|第二十四是 羅幔提‧以謝 ，他兒子和他兄弟共十二人。
1CHR|26|1|門口守衛的班次如下： 可拉 族 以比雅撒 的子孫中，有 可利 的兒子 米施利米雅 。
1CHR|26|2|米施利米雅 的長子是 撒迦利亞 ，次子是 耶疊 ，三子是 西巴第雅 ，四子是 耶提聶 ，
1CHR|26|3|五子是 以攔 ，六子是 約哈難 ，七子是 以利約乃 。
1CHR|26|4|俄別‧以東 的長子是 示瑪雅 ，次子是 約薩拔 ，三子是 約亞 ，四子是 沙甲 ，五子是 拿坦業 ，
1CHR|26|5|六子是 亞米利 ，七子是 以薩迦 ，八子是 毗烏利太 ，因為上帝賜福給 俄別‧以東 。
1CHR|26|6|他的兒子 示瑪雅 生了幾個兒子，都是大能的勇士，管理父親的家。
1CHR|26|7|示瑪雅 的兒子是 俄得尼 、 利法益 、 俄備得 、 以利薩巴 。 以利薩巴 的兄弟 以利戶 和 西瑪迦 是能人。
1CHR|26|8|這些都是 俄別‧以東 的子孫，他們和他們的兒子，以及兄弟，都是善於辦事的能人。屬 俄別‧以東 的共六十二人。
1CHR|26|9|米施利米雅 的兒子和兄弟都是能人，共十八人。
1CHR|26|10|米拉利 子孫中的 何薩 有幾個兒子：為首的是 申利 ；他原不是長子，是他父親立他為首的，
1CHR|26|11|次子是 希勒家 ，三子是 底巴利雅 ，四子是 撒迦利亞 。 何薩 的兒子和兄弟共十三人。
1CHR|26|12|這些是門口守衛的班次，各隨他們的班長，與他們的兄弟一同在耶和華殿裏按班供職。
1CHR|26|13|他們無論大小，都按著父系抽籤，分守各門。
1CHR|26|14|抽到東門的是 示利米雅 ；他的兒子 撒迦利亞 是精明的謀士，抽到北門。
1CHR|26|15|俄別‧以東 守南門，他的兒子守倉庫。
1CHR|26|16|書聘 與 何薩 守西門，在靠近 沙利基 門、通往上去的街道上，守衛與守衛相對。
1CHR|26|17|東門有六個 利未 人 ，北門每日有四人，南門每日有四人，庫房有兩人輪流替換。
1CHR|26|18|至於走廊，在西面街道上有四人，在走廊上有兩人。
1CHR|26|19|以上是 可拉 子孫和 米拉利 子孫門口守衛的班次。
1CHR|26|20|利未 人中有 亞希雅 管理上帝殿的庫房和聖物的庫房。
1CHR|26|21|拉但 子孫中， 革順 族屬 拉但 、作族長的是 革順 族屬 拉但 的 耶希伊利 。
1CHR|26|22|耶希伊利 的兒子 西坦 和他兄弟 約珥 管理耶和華殿的庫房。
1CHR|26|23|暗蘭 人、 以斯哈 人、 希伯倫 人、 烏薛 人也有職務。
1CHR|26|24|摩西 的孫子， 革舜 的兒子 細布業 管理庫房。
1CHR|26|25|還有他的弟兄： 以利以謝 ， 以利以謝 的兒子 利哈比雅 ， 利哈比雅 的兒子 耶篩亞 ， 耶篩亞 的兒子 約蘭 ， 約蘭 的兒子 細基利 ， 細基利 的兒子 示羅密 。
1CHR|26|26|這 示羅密 和他的兄弟管理一切庫房的聖物，就是 大衛 王和眾族長、千夫長、百夫長，以及軍官所分別為聖之物。
1CHR|26|27|他們把打仗時奪取的一些財物分別為聖，用來修造耶和華的殿。
1CHR|26|28|凡 撒母耳 先見、 基士 的兒子 掃羅 、 尼珥 的兒子 押尼珥 、 洗魯雅 的兒子 約押 分別為聖的，一切分別為聖之物都歸 示羅密 和他的兄弟掌管。
1CHR|26|29|以斯哈 人有 基拿尼雅 和他眾兒子作官長和審判官，管理 以色列 對外的事務。
1CHR|26|30|希伯倫 人有 哈沙比雅 和他弟兄一千七百人，都是能人，在 約旦河 西監督 以色列 人，辦理耶和華的一切工作和王的事務。
1CHR|26|31|希伯倫 人中有 耶利雅 作族長。 大衛 作王第四十年在各族各家從事尋訪，在 基列 的 雅謝 ，從這族中發現大能的勇士。
1CHR|26|32|耶利雅 的弟兄有二千七百人，都是能人，又是族長； 大衛 王派他們在 呂便 人、 迦得 人、 瑪拿西 半支派中管理上帝和王的一切事務。
1CHR|27|1|以色列 人的族長、千夫長、百夫長和官長都分配班次，每班二萬四千人，整年按月輪流出入，按班次服事王。
1CHR|27|2|正月第一班的班長是 撒巴第業 的兒子 雅朔班 ；他班內有二萬四千人。
1CHR|27|3|他是 法勒斯 的後裔，統管正月軍隊所有的官長。
1CHR|27|4|二月的班長是 亞何亞 人 朵代 ，他的班有總長 密基羅 ；他班內有二萬四千人。
1CHR|27|5|三月第三班的班長是 耶何耶大 祭司長的兒子 比拿雅 ；他班內有二萬四千人。
1CHR|27|6|這 比拿雅 是那三十人中的勇士，管理那三十人；他班內又有他兒子 暗米薩拔 。
1CHR|27|7|四月第四班的班長是 約押 的兄弟 亞撒黑 。接續他的是他兒子 西巴第雅 ；他班內有二萬四千人。
1CHR|27|8|五月第五班的班長是 伊斯拉 人 珊合 ；他班內有二萬四千人。
1CHR|27|9|六月第六班的班長是 提哥亞 人 益吉 的兒子 以拉 ；他班內有二萬四千人。
1CHR|27|10|七月第七班的班長是 以法蓮 族 比倫 人 希利斯 ；他班內有二萬四千人。
1CHR|27|11|八月第八班的班長是 謝拉 族 戶沙 人 西比該 ；他班內有二萬四千人。
1CHR|27|12|九月第九班的班長是 便雅憫 族 亞拿突 人 亞比以謝 ；他班內有二萬四千人。
1CHR|27|13|十月第十班的班長是 謝拉 族 尼陀法 人 瑪哈萊 ；他班內有二萬四千人。
1CHR|27|14|十一月第十一班的班長是 以法蓮 族 比拉頓 人 比拿雅 ；他班內有二萬四千人。
1CHR|27|15|十二月第十二班的班長是 俄陀聶 族 尼陀法 人 黑玳 ；他班內有二萬四千人。
1CHR|27|16|管理 以色列 眾支派的如下：管 呂便 人的是 細基利 的兒子 以利以謝 ；管 西緬 人的是 瑪迦 的兒子 示法提雅 ；
1CHR|27|17|管 利未 的是 基摩利 的兒子 哈沙比雅 ；管 亞倫 子孫的是 撒督 ；
1CHR|27|18|管 猶大 的是 大衛 的一個哥哥 以利戶 ；管 以薩迦 的是 米迦勒 的兒子 暗利 ；
1CHR|27|19|管 西布倫 的是 俄巴第雅 的兒子 伊施瑪雅 ；管 拿弗他利 的是 亞斯列 的兒子 耶利摩 ；
1CHR|27|20|管 以法蓮 的是 阿撒細雅 的兒子 何細亞 ；管 瑪拿西 半支派的是 毗大雅 的兒子 約珥 ；
1CHR|27|21|管 基列 地 瑪拿西 半支派的是 撒迦利亞 的兒子 易多 ；管 便雅憫 的是 押尼珥 的兒子 雅西業 ；
1CHR|27|22|管 但 的是 耶羅罕 的兒子 亞薩列 。以上是 以色列 眾支派的領袖。
1CHR|27|23|以色列 人二十歲以下的， 大衛 沒有記其數目；因耶和華曾應許，必加增 以色列 人如天上的星那樣多。
1CHR|27|24|洗魯雅 的兒子 約押 開始數點，卻還沒有數完。為了這事，烈怒臨到 以色列 ，數點的數目也沒有寫在《大衛王記》上。
1CHR|27|25|管理王的庫房的是 亞疊 的兒子 押斯馬威 。管理田野、城鎮、村莊、堡壘之倉庫的是 烏西雅 的兒子 約拿單 。
1CHR|27|26|管理耕田種地的是 基綠 的兒子 以斯利 。
1CHR|27|27|管理葡萄園的是 拉瑪 人 示每 。管理葡萄園酒窖的是 實弗米 人 撒巴底 。
1CHR|27|28|管理 謝非拉 橄欖樹和桑樹的是 基第利 人 巴勒‧哈南 。管理油庫的是 約阿施 。
1CHR|27|29|管理 沙崙 牧放牛群的是 沙崙 人 施提萊 。管理山谷牧養牛群的是 亞第萊 的兒子 沙法 。
1CHR|27|30|管理駱駝群的是 以實瑪利 人 阿比勒 。管理驢群的是 米崙 人 耶希底亞 。管理羊群的是 夏甲 人 雅悉 。
1CHR|27|31|這些都是為 大衛 王管理產業的領袖。
1CHR|27|32|大衛 的叔父 約拿單 作謀士；這人有智慧，又作書記。 哈摩尼 的兒子 耶歇 陪伴王的眾兒子。
1CHR|27|33|亞希多弗 作王的謀士。 亞基 人 戶篩 作王的顧問。
1CHR|27|34|亞希多弗 之後，有 比拿雅 的兒子 耶何耶大 ，以及 亞比亞他 接續他。 約押 作王的元帥。
1CHR|28|1|大衛 召集 以色列 所有的領袖，各支派的領袖、輪班服事王的官長、千夫長、百夫長、掌管王和王子一切產業牲畜的、宮廷官員、勇士，和所有大能的勇士，都到 耶路撒冷 來。
1CHR|28|2|大衛 王站起來，說：「我的弟兄，我的百姓啊，請聽我說！我心裏本想建造殿宇，安放耶和華的約櫃，作為我們上帝的腳凳，並且我已經預備了建造的材料。
1CHR|28|3|只是上帝對我說：『你不可為我的名建造殿宇，因你是戰士，流了人的血。』
1CHR|28|4|然而，耶和華－ 以色列 的上帝在我父的全家揀選我作 以色列 的王，直到永遠。因他揀選 猶大 為領袖，在 猶大 家中揀選我父家，在我父的眾兒子裏喜悅我，立我作全 以色列 的王。
1CHR|28|5|耶和華賜我許多兒子，在我兒子中揀選我兒子 所羅門 坐耶和華國度的王位，治理 以色列 。
1CHR|28|6|耶和華對我說：『你兒子 所羅門 必建造我的殿和院宇，因為我揀選他作我的子，我也必作他的父。
1CHR|28|7|他若恆久遵行我的誡命典章如今日一樣，我就必堅定他的國，直到永遠。』
1CHR|28|8|現今在 以色列 眾人眼前，在耶和華的會中，在我們上帝的垂聽下，你們務要遵行並尋求耶和華－你們上帝的一切誡命，如此你們就可以承受這美地，並留給你們的子孫，永遠為業。
1CHR|28|9|「我兒 所羅門 哪，你當認識耶和華－你父的上帝，全心樂意地事奉他，因為耶和華鑒察眾人的心，知道一切心思意念。你若尋求他，他必使你尋見；你若離棄他，他必永遠丟棄你。
1CHR|28|10|現在你當謹慎，因耶和華揀選你建造殿宇作為聖所。你當剛強去做。」
1CHR|28|11|大衛 指示他兒子 所羅門 有關殿的走廊、屋子、庫房、樓房、內殿和櫃蓋 之處的樣式，
1CHR|28|12|被靈感動所得的一切樣式：耶和華殿的院子、周圍一切的房屋、上帝殿的庫房和聖物庫房；
1CHR|28|13|祭司和 利未 人的班次，耶和華殿裏各樣事奉的工作，耶和華殿裏一切事奉用的器皿，
1CHR|28|14|以及各樣事奉所用金器的重量，和各樣事奉所用銀器的重量，
1CHR|28|15|金燈臺和金燈的重量，按每一個燈臺和燈的重量；銀燈臺和銀燈的重量，按每一個燈臺和燈的重量，都按照每一個燈臺的用途；
1CHR|28|16|每張供餅桌子的金子重量，和銀桌子的銀子重量，
1CHR|28|17|純金的肉叉子、盤子，和壺的重量，金碗，按每個金碗的重量，和銀碗，按每個銀碗的重量，
1CHR|28|18|純金香壇的重量，金基路伯座車的樣式，基路伯張開翅膀，遮蓋耶和華的約櫃。
1CHR|28|19|大衛 說：「這一切，所有工作的樣式，是耶和華用手寫的文件使我明白的。」
1CHR|28|20|大衛 又對他兒子 所羅門 說：「你當剛強壯膽去做！不要懼怕，也不要驚惶，因為耶和華上帝，我的上帝與你同在。他必不撇下你，也不丟棄你，直到耶和華殿的工作都完畢。
1CHR|28|21|看哪，有祭司和 利未 人的班次，為要辦理上帝殿各樣的事務，又有擅長做各樣事務的人，樂意在各樣工作上幫助你，並且領袖和眾百姓也都聽從你的一切命令。」
1CHR|29|1|大衛 王對全會眾說：「我兒子 所羅門 是上帝特選的，還年幼脆弱，但這工程浩大，因這殿不是為人，而是為耶和華上帝建造的。
1CHR|29|2|我為我上帝的殿已經盡力，預備金子做金器，銀子做銀器，銅做銅器，鐵做鐵器，木做木器，還有紅瑪瑙、可鑲嵌的寶石、彩石、各樣的寶石和許多大理石。
1CHR|29|3|此外，因我愛慕我上帝的殿，在預備建造聖殿的一切材料之外，又將我自己積蓄的金銀獻給我上帝的殿，
1CHR|29|4|就是三千他連得 俄斐 金子、七千他連得純銀，用來貼殿的牆；
1CHR|29|5|金子做金器，銀子做銀器，並藉工匠的手做一切的工。今日有誰願意將自己獻給耶和華呢？」
1CHR|29|6|於是，眾族長和 以色列 各支派的領袖、千夫長、百夫長，以及監管王工作的官長，都樂意奉獻。
1CHR|29|7|他們為上帝殿的工程獻上五千他連得又一萬達利克 金子，一萬他連得銀子，一萬八千他連得銅，十萬他連得鐵。
1CHR|29|8|凡有寶石的都送入耶和華殿的庫房，由 革順 人 耶歇 的手管理。
1CHR|29|9|因這些人全心樂意獻給耶和華，百姓就歡喜， 大衛 王也大大歡喜。
1CHR|29|10|大衛 在全會眾眼前稱頌耶和華； 大衛 說：「耶和華－ 以色列 的上帝，我們的父，你是應當稱頌的，直到永永遠遠！
1CHR|29|11|耶和華啊，尊大、能力、榮耀、勝利、威嚴都是你的；天上地下的一切都是你的；耶和華啊，國度是你的，並且你為至高，為萬有之首。
1CHR|29|12|豐富尊榮都從你而來，你也治理萬物。在你手裏有大能大力，你的手使人尊大強盛。
1CHR|29|13|我們的上帝啊，現在我們稱謝你，讚美你榮耀之名！
1CHR|29|14|「我算甚麼，我的百姓算甚麼，竟然能夠如此樂意奉獻？因為萬物都從你而來，我們把從你的手得來的獻給你。
1CHR|29|15|我們在你面前是客旅，是寄居的，與我們的列祖一樣。我們在世的日子如影子，沒有盼望。
1CHR|29|16|耶和華－我們的上帝啊，我們預備這許多材料，要為你的聖名建造殿宇，都是從你的手而來，都是屬你的。
1CHR|29|17|我的上帝啊，我知道你察驗人心，喜悅正直；我以正直的心樂意獻上這一切。現在我歡喜見你的百姓在此樂意奉獻給你。
1CHR|29|18|耶和華－我們列祖 亞伯拉罕 、 以撒 、 以色列 的上帝啊，求你使你的百姓心中常存這樣的心思意念，堅定他們的心歸向你，
1CHR|29|19|又求你賜我兒子 所羅門 全心遵守你的命令、法度、律例，成就這一切的事，用我所預備的建造殿宇。」
1CHR|29|20|大衛 對全會眾說：「你們應當稱頌耶和華－你們的上帝。」於是全會眾稱頌耶和華－他們列祖的上帝，低頭向耶和華和王下拜。
1CHR|29|21|次日，他們向耶和華獻平安祭和燔祭，獻一千頭公牛，一千隻公綿羊，一千隻羔羊，以及同獻的澆酒祭，並為 以色列 眾人獻許多的祭。
1CHR|29|22|那日，他們在耶和華面前吃喝，大大歡樂。 他們再次立 大衛 的兒子 所羅門 作王，膏他歸耶和華作君王，又膏 撒督 作祭司。
1CHR|29|23|於是 所羅門 坐在耶和華所賜的王位上，接續他父親 大衛 作王；他萬事亨通，全 以色列 都聽從他。
1CHR|29|24|眾領袖和勇士，以及 大衛 王的眾兒子，都順服 所羅門 王。
1CHR|29|25|耶和華使 所羅門 在 以色列 眾人眼前非常尊大，賜他君王的威嚴，勝過他以前任何一位 以色列 王。
1CHR|29|26|耶西 的兒子 大衛 作全 以色列 的王。
1CHR|29|27|他作 以色列 王的時期共四十年：在 希伯崙 作王七年，在 耶路撒冷 作王三十三年。
1CHR|29|28|他死的時候年紀老邁，日子滿足，享盡榮華富貴。他的兒子 所羅門 接續他作王。
1CHR|29|29|大衛 王自始至終的事蹟，看哪，都寫在 撒母耳 先見的書上、 拿單 先知的書上和 迦得 先見的書上，
1CHR|29|30|包括他治國的一切和他英勇的事蹟，以及他和 以色列 與世上列國所經歷的事。
