EXOD|1|1|haec sunt nomina filiorum Israhel qui ingressi sunt Aegyptum cum Iacob singuli cum domibus suis introierunt
EXOD|1|2|Ruben Symeon Levi Iuda
EXOD|1|3|Isachar Zabulon et Beniamin
EXOD|1|4|Dan et Nepthalim Gad et Aser
EXOD|1|5|erant igitur omnes animae eorum qui egressi sunt de femore Iacob septuaginta Ioseph autem in Aegypto erat
EXOD|1|6|quo mortuo et universis fratribus eius omnique cognatione illa
EXOD|1|7|filii Israhel creverunt et quasi germinantes multiplicati sunt ac roborati nimis impleverunt terram
EXOD|1|8|surrexit interea rex novus super Aegyptum qui ignorabat Ioseph
EXOD|1|9|et ait ad populum suum ecce populus filiorum Israhel multus et fortior nobis
EXOD|1|10|venite sapienter opprimamus eum ne forte multiplicetur et si ingruerit contra nos bellum addatur inimicis nostris expugnatisque nobis egrediatur e terra
EXOD|1|11|praeposuit itaque eis magistros operum ut adfligerent eos oneribus aedificaveruntque urbes tabernaculorum Pharaoni Phiton et Ramesses
EXOD|1|12|quantoque opprimebant eos tanto magis multiplicabantur et crescebant
EXOD|1|13|oderantque filios Israhel Aegyptii et adfligebant inludentes eis
EXOD|1|14|atque ad amaritudinem perducebant vitam eorum operibus duris luti et lateris omnique famulatu quo in terrae operibus premebantur
EXOD|1|15|dixit autem rex Aegypti obsetricibus Hebraeorum quarum una vocabatur Sephra altera Phua
EXOD|1|16|praecipiens eis quando obsetricabitis Hebraeas et partus tempus advenerit si masculus fuerit interficite illum si femina reservate
EXOD|1|17|timuerunt autem obsetrices Deum et non fecerunt iuxta praeceptum regis Aegypti sed conservabant mares
EXOD|1|18|quibus ad se accersitis rex ait quidnam est hoc quod facere voluistis ut pueros servaretis
EXOD|1|19|quae responderunt non sunt hebraeae sicut aegyptiae mulieres ipsae enim obsetricandi habent scientiam et priusquam veniamus ad eas pariunt
EXOD|1|20|bene ergo fecit Deus obsetricibus et crevit populus confortatusque est nimis
EXOD|1|21|et quia timuerant obsetrices Deum aedificavit illis domos
EXOD|1|22|praecepit autem Pharao omni populo suo dicens quicquid masculini sexus natum fuerit in flumen proicite quicquid feminei reservate
EXOD|2|1|egressus est post haec vir de domo Levi accepta uxore stirpis suae
EXOD|2|2|quae concepit et peperit filium et videns eum elegantem abscondit tribus mensibus
EXOD|2|3|cumque iam celare non posset sumpsit fiscellam scirpeam et linivit eam bitumine ac pice posuitque intus infantulum et exposuit eum in carecto ripae fluminis
EXOD|2|4|stante procul sorore eius et considerante eventum rei
EXOD|2|5|ecce autem descendebat filia Pharaonis ut lavaretur in flumine et puellae eius gradiebantur per crepidinem alvei quae cum vidisset fiscellam in papyrione misit unam e famulis suis et adlatam
EXOD|2|6|aperiens cernensque in ea parvulum vagientem miserta eius ait de infantibus Hebraeorum est
EXOD|2|7|cui soror pueri vis inquit ut vadam et vocem tibi hebraeam mulierem quae nutrire possit infantulum
EXOD|2|8|respondit vade perrexit puella et vocavit matrem eius
EXOD|2|9|ad quam locuta filia Pharaonis accipe ait puerum istum et nutri mihi ego tibi dabo mercedem tuam suscepit mulier et nutrivit puerum adultumque tradidit filiae Pharaonis
EXOD|2|10|quem illa adoptavit in locum filii vocavitque nomen eius Mosi dicens quia de aqua tuli eum
EXOD|2|11|in diebus illis postquam creverat Moses egressus ad fratres suos vidit adflictionem eorum et virum aegyptium percutientem quendam de Hebraeis fratribus suis
EXOD|2|12|cumque circumspexisset huc atque illuc et nullum adesse vidisset percussum Aegyptium abscondit sabulo
EXOD|2|13|et egressus die altero conspexit duos Hebraeos rixantes dixitque ei qui faciebat iniuriam quare percutis proximum tuum
EXOD|2|14|qui respondit quis constituit te principem et iudicem super nos num occidere me tu dicis sicut occidisti Aegyptium timuit Moses et ait quomodo palam factum est verbum istud
EXOD|2|15|audivitque Pharao sermonem hunc et quaerebat occidere Mosen qui fugiens de conspectu eius moratus est in terra Madian et sedit iuxta puteum
EXOD|2|16|erant sacerdoti Madian septem filiae quae venerunt ad hauriendas aquas et impletis canalibus adaquare cupiebant greges patris sui
EXOD|2|17|supervenere pastores et eiecerunt eas surrexitque Moses et defensis puellis adaquavit oves earum
EXOD|2|18|quae cum revertissent ad Raguhel patrem suum dixit ad eas cur velocius venistis solito
EXOD|2|19|responderunt vir aegyptius liberavit nos de manu pastorum insuper et hausit aquam nobiscum potumque dedit ovibus
EXOD|2|20|at ille ubi est inquit quare dimisistis hominem vocate eum ut comedat panem
EXOD|2|21|iuravit ergo Moses quod habitaret cum eo accepitque Sefforam filiam eius
EXOD|2|22|quae peperit filium quem vocavit Gersam dicens advena fui in terra aliena
EXOD|2|23|post multum temporis mortuus est rex Aegypti et ingemescentes filii Israhel propter opera vociferati sunt ascenditque clamor eorum ad Deum ab operibus
EXOD|2|24|et audivit gemitum eorum ac recordatus foederis quod pepigerat cum Abraham et Isaac et Iacob
EXOD|2|25|respexit filios Israhel et cognovit eos
EXOD|3|1|Moses autem pascebat oves Iethro cognati sui sacerdotis Madian cumque minasset gregem ad interiora deserti venit ad montem Dei Horeb
EXOD|3|2|apparuitque ei Dominus in flamma ignis de medio rubi et videbat quod rubus arderet et non conbureretur
EXOD|3|3|dixit ergo Moses vadam et videbo visionem hanc magnam quare non conburatur rubus
EXOD|3|4|cernens autem Dominus quod pergeret ad videndum vocavit eum de medio rubi et ait Moses Moses qui respondit adsum
EXOD|3|5|at ille ne adpropies inquit huc solve calciamentum de pedibus tuis locus enim in quo stas terra sancta est
EXOD|3|6|et ait ego sum Deus patris tui Deus Abraham Deus Isaac Deus Iacob abscondit Moses faciem suam non enim audebat aspicere contra Deum
EXOD|3|7|cui ait Dominus vidi adflictionem populi mei in Aegypto et clamorem eius audivi propter duritiam eorum qui praesunt operibus
EXOD|3|8|et sciens dolorem eius descendi ut liberarem eum de manibus Aegyptiorum et educerem de terra illa in terram bonam et spatiosam in terram quae fluit lacte et melle ad loca Chananei et Hetthei et Amorrei Ferezei et Evei et Iebusei
EXOD|3|9|clamor ergo filiorum Israhel venit ad me vidique adflictionem eorum qua ab Aegyptiis opprimuntur
EXOD|3|10|sed veni mittam te ad Pharaonem ut educas populum meum filios Israhel de Aegypto
EXOD|3|11|dixit Moses ad Deum quis ego sum ut vadam ad Pharaonem et educam filios Israhel de Aegypto
EXOD|3|12|qui dixit ei ero tecum et hoc habebis signum quod miserim te cum eduxeris populum de Aegypto immolabis Deo super montem istum
EXOD|3|13|ait Moses ad Deum ecce ego vadam ad filios Israhel et dicam eis Deus patrum vestrorum misit me ad vos si dixerint mihi quod est nomen eius quid dicam eis
EXOD|3|14|dixit Deus ad Mosen ego sum qui sum ait sic dices filiis Israhel qui est misit me ad vos
EXOD|3|15|dixitque iterum Deus ad Mosen haec dices filiis Israhel Dominus Deus patrum vestrorum Deus Abraham Deus Isaac et Deus Iacob misit me ad vos hoc nomen mihi est in aeternum et hoc memoriale meum in generationem et generatione
EXOD|3|16|vade congrega seniores Israhel et dices ad eos Dominus Deus patrum vestrorum apparuit mihi Deus Abraham et Deus Isaac et Deus Iacob dicens visitans visitavi vos et omnia quae acciderunt vobis in Aegypto
EXOD|3|17|et dixi ut educam vos de adflictione Aegypti in terram Chananei et Hetthei et Amorrei Ferezei et Evei et Iebusei ad terram fluentem lacte et melle
EXOD|3|18|et audient vocem tuam ingredierisque tu et seniores Israhel ad regem Aegypti et dices ad eum Dominus Deus Hebraeorum vocavit nos ibimus viam trium dierum per solitudinem ut immolemus Domino Deo nostro
EXOD|3|19|sed ego scio quod non dimittet vos rex Aegypti ut eatis nisi per manum validam
EXOD|3|20|extendam enim manum meam et percutiam Aegyptum in cunctis mirabilibus meis quae facturus sum in medio eorum post haec dimittet vos
EXOD|3|21|daboque gratiam populo huic coram Aegyptiis et cum egrediemini non exibitis vacui
EXOD|3|22|sed postulabit mulier a vicina sua et ab hospita vasa argentea et aurea ac vestes ponetisque eas super filios et filias vestras et spoliabitis Aegyptum
EXOD|4|1|respondens Moses ait non credent mihi neque audient vocem meam sed dicent non apparuit tibi Dominus
EXOD|4|2|dixit ergo ad eum quid est hoc quod tenes in manu tua respondit virga
EXOD|4|3|ait proice eam in terram proiecit et versa est in colubrum ita ut fugeret Moses
EXOD|4|4|dixitque Dominus extende manum tuam et adprehende caudam eius extendit et tenuit versaque est in virgam
EXOD|4|5|ut credant inquit quod apparuerit tibi Dominus Deus patrum tuorum Deus Abraham Deus Isaac Deus Iacob
EXOD|4|6|dixitque Dominus rursum mitte manum in sinum tuum quam cum misisset in sinum protulit leprosam instar nivis
EXOD|4|7|retrahe ait manum in sinum tuum retraxit et protulit iterum et erat similis carni reliquae
EXOD|4|8|si non crediderint inquit tibi neque audierint sermonem signi prioris credent verbo signi sequentis
EXOD|4|9|quod si nec duobus quidem his signis crediderint neque audierint vocem tuam sume aquam fluminis et effunde eam super aridam et quicquid hauseris de fluvio vertetur in sanguinem
EXOD|4|10|ait Moses obsecro Domine non sum eloquens ab heri et nudius tertius et ex quo locutus es ad servum tuum inpeditioris et tardioris linguae sum
EXOD|4|11|dixit Dominus ad eum quis fecit os hominis aut quis fabricatus est mutum et surdum videntem et caecum nonne ego
EXOD|4|12|perge igitur et ego ero in ore tuo doceboque te quid loquaris
EXOD|4|13|at ille obsecro inquit Domine mitte quem missurus es
EXOD|4|14|iratus Dominus in Mosen ait Aaron frater tuus Levites scio quod eloquens sit ecce ipse egreditur in occursum tuum vidensque te laetabitur corde
EXOD|4|15|loquere ad eum et pone verba mea in ore eius ego ero in ore tuo et in ore illius et ostendam vobis quid agere debeatis
EXOD|4|16|ipse loquetur pro te ad populum et erit os tuum tu autem eris ei in his quae ad Deum pertinent
EXOD|4|17|virgam quoque hanc sume in manu tua in qua facturus es signa
EXOD|4|18|abiit Moses et reversus est ad Iethro cognatum suum dixitque ei vadam et revertar ad fratres meos in Aegyptum ut videam si adhuc vivunt cui ait Iethro vade in pace
EXOD|4|19|dixit ergo Dominus ad Mosen in Madian vade revertere in Aegyptum mortui sunt omnes qui quaerebant animam tuam
EXOD|4|20|tulit Moses uxorem et filios suos et inposuit eos super asinum reversusque est in Aegyptum portans virgam Dei in manu sua
EXOD|4|21|dixitque ei Dominus revertenti in Aegyptum vide ut omnia ostenta quae posui in manu tua facias coram Pharaone ego indurabo cor eius et non dimittet populum
EXOD|4|22|dicesque ad eum haec dicit Dominus filius meus primogenitus meus Israhel
EXOD|4|23|dixi tibi dimitte filium meum ut serviat mihi et noluisti dimittere eum ecce ego interficiam filium tuum primogenitum
EXOD|4|24|cumque esset in itinere in diversorio occurrit ei Dominus et volebat occidere eum
EXOD|4|25|tulit ilico Seffora acutissimam petram et circumcidit praeputium filii sui tetigitque pedes eius et ait sponsus sanguinum tu mihi es
EXOD|4|26|et dimisit eum postquam dixerat sponsus sanguinum ob circumcisionem
EXOD|4|27|dixit autem Dominus ad Aaron vade in occursum Mosi in deserto qui perrexit ei obviam in montem Dei et osculatus est eum
EXOD|4|28|narravitque Moses Aaron omnia verba Domini quibus miserat eum et signa quae mandaverat
EXOD|4|29|veneruntque simul et congregaverunt cunctos seniores filiorum Israhel
EXOD|4|30|locutusque est Aaron omnia verba quae dixerat Dominus ad Mosen et fecit signa coram populo
EXOD|4|31|et credidit populus audieruntque quod visitasset Dominus filios Israhel et quod respexisset adflictionem eorum et proni adoraverunt
EXOD|5|1|post haec ingressi sunt Moses et Aaron et dixerunt Pharaoni haec dicit Dominus Deus Israhel dimitte populum meum ut sacrificet mihi in deserto
EXOD|5|2|at ille respondit quis est Dominus ut audiam vocem eius et dimittam Israhel nescio Dominum et Israhel non dimittam
EXOD|5|3|dixerunt Deus Hebraeorum vocavit nos ut eamus viam trium dierum in solitudinem et sacrificemus Domino Deo nostro ne forte accidat nobis pestis aut gladius
EXOD|5|4|ait ad eos rex Aegypti quare Moses et Aaron sollicitatis populum ab operibus suis ite ad onera vestra
EXOD|5|5|dixitque Pharao multus est populus terrae videtis quod turba succreverit quanto magis si dederitis eis requiem ab operibus
EXOD|5|6|praecepit ergo in die illo praefectis operum et exactoribus populi dicens
EXOD|5|7|nequaquam ultra dabitis paleas populo ad conficiendos lateres sicut prius sed ipsi vadant et colligant stipulam
EXOD|5|8|et mensuram laterum quos prius faciebant inponetis super eos nec minuetis quicquam vacant enim et idcirco vociferantur dicentes eamus et sacrificemus Deo nostro
EXOD|5|9|opprimantur operibus et expleant ea ut non adquiescant verbis mendacibus
EXOD|5|10|igitur egressi praefecti operum et exactores ad populum dixerunt sic dicit Pharao non do vobis paleas
EXOD|5|11|ite et colligite sicubi invenire potueritis nec minuetur quicquam de opere vestro
EXOD|5|12|dispersusque est populus per omnem terram Aegypti ad colligendas paleas
EXOD|5|13|praefecti quoque operum instabant dicentes conplete opus vestrum cotidie ut prius facere solebatis quando dabantur vobis paleae
EXOD|5|14|flagellatique sunt qui praeerant operibus filiorum Israhel ab exactoribus Pharaonis dicentibus quare non impletis mensuram laterum sicut prius nec heri nec hodie
EXOD|5|15|veneruntque praepositi filiorum Israhel et vociferati sunt ad Pharaonem dicentes cur ita agis contra servos tuos
EXOD|5|16|paleae non dantur nobis et lateres similiter imperantur en famuli tui flagellis caedimur et iniuste agitur contra populum tuum
EXOD|5|17|qui ait vacatis otio et idcirco dicitis eamus et sacrificemus Domino
EXOD|5|18|ite ergo et operamini paleae non dabuntur vobis et reddetis consuetum numerum laterum
EXOD|5|19|videbantque se praepositi filiorum Israhel in malo eo quod diceretur eis non minuetur quicquam de lateribus per singulos dies
EXOD|5|20|occurreruntque Mosi et Aaron qui stabant ex adverso egredientes a Pharaone
EXOD|5|21|et dixerunt ad eos videat Dominus et iudicet quoniam fetere fecistis odorem nostrum coram Pharao et servis eius et praebuistis ei gladium ut occideret nos
EXOD|5|22|reversusque Moses ad Dominum ait Domine cur adflixisti populum istum quare misisti me
EXOD|5|23|ex eo enim quo ingressus sum ad Pharaonem ut loquerer nomine tuo adflixit populum tuum et non liberasti eos
EXOD|6|1|dixit Dominus ad Mosen nunc videbis quae facturus sum Pharaoni per manum enim fortem dimittet eos et in manu robusta eiciet illos de terra sua
EXOD|6|2|locutusque est Dominus ad Mosen dicens ego Dominus
EXOD|6|3|qui apparui Abraham Isaac et Iacob in Deo omnipotente et nomen meum Adonai non indicavi eis
EXOD|6|4|pepigique cum eis foedus ut darem illis terram Chanaan terram peregrinationis eorum in qua fuerunt advenae
EXOD|6|5|ego audivi gemitum filiorum Israhel quo Aegyptii oppresserunt eos et recordatus sum pacti mei
EXOD|6|6|ideo dic filiis Israhel ego Dominus qui educam vos de ergastulo Aegyptiorum et eruam de servitute ac redimam in brachio excelso et iudiciis magnis
EXOD|6|7|et adsumam vos mihi in populum et ero vester Deus scietisque quod ego sim Dominus Deus vester qui eduxerim vos de ergastulo Aegyptiorum
EXOD|6|8|et induxerim in terram super quam levavi manum meam ut darem eam Abraham Isaac et Iacob daboque illam vobis possidendam ego Dominus
EXOD|6|9|narravit ergo Moses omnia filiis Israhel qui non adquieverunt ei propter angustiam spiritus et opus durissimum
EXOD|6|10|locutusque est Dominus ad Mosen dicens
EXOD|6|11|ingredere et loquere ad Pharao regem Aegypti ut dimittat filios Israhel de terra sua
EXOD|6|12|respondit Moses coram Domino ecce filii Israhel non me audiunt et quomodo audiet me Pharao praesertim cum sim incircumcisus labiis
EXOD|6|13|locutus est Dominus ad Mosen et Aaron et dedit mandatum ad filios Israhel et ad Pharao regem Aegypti ut educerent filios Israhel de terra Aegypti
EXOD|6|14|isti sunt principes domorum per familias suas filii Ruben primogeniti Israhelis Enoch et Phallu Aesrom et Charmi
EXOD|6|15|hae cognationes Ruben filii Symeon Iamuhel et Iamin et Aod Iachin et Soer et Saul filius Chananitidis hae progenies Symeon
EXOD|6|16|et haec nomina filiorum Levi per cognationes suas Gerson et Caath et Merari anni autem vitae Levi fuerunt centum triginta septem
EXOD|6|17|filii Gerson Lobeni et Semei per cognationes suas
EXOD|6|18|filii Caath Amram et Isuar et Hebron et Ozihel annique vitae Caath centum triginta tres
EXOD|6|19|filii Merari Mooli et Musi hae cognationes Levi per familias suas
EXOD|6|20|accepit autem Amram uxorem Iocabed patruelem suam quae peperit ei Aaron et Mosen fueruntque anni vitae Amram centum triginta septem
EXOD|6|21|filii quoque Isuar Core et Napheg et Zechri
EXOD|6|22|filii quoque Ozihel Misahel et Elsaphan et Sethri
EXOD|6|23|accepit autem Aaron uxorem Elisabe filiam Aminadab sororem Naasson quae peperit ei Nadab et Abiu et Eleazar et Ithamar
EXOD|6|24|filii quoque Core Asir et Helcana et Abiasab hae sunt cognationes Coritarum
EXOD|6|25|at vero Eleazar filius Aaron accepit uxorem de filiabus Phutihel quae peperit ei Finees hii sunt principes familiarum leviticarum per cognationes suas
EXOD|6|26|iste est Aaron et Moses quibus praecepit Dominus ut educerent filios Israhel de terra Aegypti per turmas suas
EXOD|6|27|hii sunt qui loquuntur ad Pharao regem Aegypti ut educant filios Israhel de Aegypto iste Moses et Aaron
EXOD|6|28|in die qua locutus est Dominus ad Mosen in terra Aegypti
EXOD|6|29|et locutus est Dominus ad Mosen dicens ego Dominus loquere ad Pharao regem Aegypti omnia quae ego loquor tibi
EXOD|6|30|et ait Moses coram Domino en incircumcisus labiis sum quomodo audiet me Pharao
EXOD|7|1|dixitque Dominus ad Mosen ecce constitui te Deum Pharaonis Aaron frater tuus erit propheta tuus
EXOD|7|2|tu loqueris omnia quae mando tibi ille loquetur ad Pharaonem ut dimittat filios Israhel de terra sua
EXOD|7|3|sed ego indurabo cor eius et multiplicabo signa et ostenta mea in terra Aegypti
EXOD|7|4|et non audiet vos inmittamque manum meam super Aegyptum et educam exercitum et populum meum filios Israhel de terra Aegypti per iudicia maxima
EXOD|7|5|et scient Aegyptii quod ego sim Dominus qui extenderim manum meam super Aegyptum et eduxerim filios Israhel de medio eorum
EXOD|7|6|fecit itaque Moses et Aaron sicut praeceperat Dominus ita egerunt
EXOD|7|7|erat autem Moses octoginta annorum et Aaron octoginta trium quando locuti sunt ad Pharaonem
EXOD|7|8|dixitque Dominus ad Mosen et Aaron
EXOD|7|9|cum dixerit vobis Pharao ostendite signa dices ad Aaron tolle virgam tuam et proice eam coram Pharao ac vertatur in colubrum
EXOD|7|10|ingressi itaque Moses et Aaron ad Pharaonem fecerunt sicut praeceperat Dominus tulitque Aaron virgam coram Pharao et servis eius quae versa est in colubrum
EXOD|7|11|vocavit autem Pharao sapientes et maleficos et fecerunt etiam ipsi per incantationes aegyptias et arcana quaedam similiter
EXOD|7|12|proieceruntque singuli virgas suas quae versae sunt in dracones sed devoravit virga Aaron virgas eorum
EXOD|7|13|induratumque est cor Pharaonis et non audivit eos sicut praeceperat Dominus
EXOD|7|14|dixit autem Dominus ad Mosen ingravatum est cor Pharaonis non vult dimittere populum
EXOD|7|15|vade ad eum mane ecce egredietur ad aquas et stabis in occursum eius super ripam fluminis et virgam quae conversa est in draconem tolles in manu tua
EXOD|7|16|dicesque ad eum Dominus Deus Hebraeorum misit me ad te dicens dimitte populum meum ut mihi sacrificet in deserto et usque ad praesens audire noluisti
EXOD|7|17|haec igitur dicit Dominus in hoc scies quod Dominus sim ecce percutiam virga quae in manu mea est aquam fluminis et vertetur in sanguinem
EXOD|7|18|pisces quoque qui sunt in fluvio morientur et conputrescent aquae et adfligentur Aegyptii bibentes aquam fluminis
EXOD|7|19|dixit quoque Dominus ad Mosen dic ad Aaron tolle virgam tuam et extende manum tuam super aquas Aegypti et super fluvios eorum et rivos ac paludes et omnes lacus aquarum ut vertantur in sanguinem et sit cruor in omni terra Aegypti tam in ligneis vasis quam in saxeis
EXOD|7|20|feceruntque ita Moses et Aaron sicut praeceperat Dominus et elevans virgam percussit aquam fluminis coram Pharao et servis eius quae versa est in sanguinem
EXOD|7|21|et pisces qui erant in flumine mortui sunt conputruitque fluvius et non poterant Aegyptii bibere aquam fluminis et fuit sanguis in tota terra Aegypti
EXOD|7|22|feceruntque similiter malefici Aegyptiorum incantationibus suis et induratum est cor Pharaonis nec audivit eos sicut praeceperat Dominus
EXOD|7|23|avertitque se et ingressus est domum suam nec adposuit cor etiam hac vice
EXOD|7|24|foderunt autem omnes Aegyptii per circuitum fluminis aquam ut biberent non enim poterant bibere de aqua fluminis
EXOD|7|25|impletique sunt septem dies postquam percussit Dominus fluvium
EXOD|8|1|dixitque Dominus ad Mosen ingredere ad Pharao et dices ad eum haec dicit Dominus dimitte populum meum ut sacrificet mihi
EXOD|8|2|sin autem nolueris dimittere ecce ego percutiam omnes terminos tuos ranis
EXOD|8|3|et ebulliet fluvius ranas quae ascendent et ingredientur domum tuam et cubiculum lectuli tui et super stratum tuum et in domos servorum tuorum et in populum tuum et in furnos tuos et in reliquias ciborum tuorum
EXOD|8|4|et ad te et ad populum tuum et ad omnes servos tuos intrabunt ranae
EXOD|8|5|dixitque Dominus ad Mosen dic Aaron extende manum tuam super fluvios et super rivos ac paludes et educ ranas super terram Aegypti
EXOD|8|6|extendit Aaron manum super aquas Aegypti et ascenderunt ranae operueruntque terram Aegypti
EXOD|8|7|fecerunt autem et malefici per incantationes suas similiter eduxeruntque ranas super terram Aegypti
EXOD|8|8|vocavit autem Pharao Mosen et Aaron et dixit orate Dominum ut auferat ranas a me et a populo meo et dimittam populum ut sacrificet Domino
EXOD|8|9|dixitque Moses Pharaoni constitue mihi quando deprecer pro te et pro servis tuis et pro populo tuo ut abigantur ranae a te et a domo tua et tantum in flumine remaneant
EXOD|8|10|qui respondit cras at ille iuxta verbum inquit tuum ut scias quoniam non est sicut Dominus Deus noster
EXOD|8|11|et recedent ranae a te et a domo tua et a servis tuis et a populo tuo tantum in flumine remanebunt
EXOD|8|12|egressique sunt Moses et Aaron a Pharaone et clamavit Moses ad Dominum pro sponsione ranarum quam condixerat Pharaoni
EXOD|8|13|fecitque Dominus iuxta verbum Mosi et mortuae sunt ranae de domibus et de villis et de agris
EXOD|8|14|congregaveruntque eas in inmensos aggeres et conputruit terra
EXOD|8|15|videns autem Pharao quod data esset requies ingravavit cor suum et non audivit eos sicut praeceperat Dominus
EXOD|8|16|dixitque Dominus ad Mosen loquere ad Aaron extende virgam tuam et percute pulverem terrae et sint scinifes in universa terra Aegypti
EXOD|8|17|feceruntque ita et extendit Aaron manu virgam tenens percussitque pulverem terrae et facti sunt scinifes in hominibus et in iumentis omnis pulvis terrae versus est in scinifes per totam terram Aegypti
EXOD|8|18|feceruntque similiter malefici incantationibus suis ut educerent scinifes et non potuerunt erantque scinifes tam in hominibus quam in iumentis
EXOD|8|19|et dixerunt malefici ad Pharao digitus Dei est induratumque est cor Pharaonis et non audivit eos sicut praeceperat Dominus
EXOD|8|20|dixit quoque Dominus ad Mosen consurge diluculo et sta coram Pharaone egreditur enim ad aquas et dices ad eum haec dicit Dominus dimitte populum meum ut sacrificet mihi
EXOD|8|21|quod si non dimiseris eum ecce ego inmittam in te et in servos tuos et in populum tuum et in domos tuas omne genus muscarum et implebuntur domus Aegyptiorum muscis diversi generis et in universa terra in qua fuerint
EXOD|8|22|faciamque mirabilem in die illa terram Gessen in qua populus meus est ut non sint ibi muscae et scias quoniam ego Dominus in medio terrae
EXOD|8|23|ponamque divisionem inter populum meum et populum tuum cras erit signum istud
EXOD|8|24|fecitque Dominus ita et venit musca gravissima in domos Pharaonis et servorum eius et in omnem terram Aegypti corruptaque est terra ab huiuscemodi muscis
EXOD|8|25|vocavit Pharao Mosen et Aaron et ait eis ite sacrificate Deo vestro in terra
EXOD|8|26|et ait Moses non potest ita fieri abominationes enim Aegyptiorum immolabimus Domino Deo nostro quod si mactaverimus ea quae colunt Aegyptii coram eis lapidibus nos obruent
EXOD|8|27|via trium dierum pergemus in solitudine et sacrificabimus Domino Deo nostro sicut praeceperit nobis
EXOD|8|28|dixitque Pharao ego dimittam vos ut sacrificetis Domino Deo vestro in deserto verumtamen longius ne abeatis rogate pro me
EXOD|8|29|et ait Moses egressus a te orabo Dominum et recedet musca a Pharaone et a servis et a populo eius cras verumtamen noli ultra fallere ut non dimittas populum sacrificare Domino
EXOD|8|30|egressusque Moses a Pharao oravit Dominum
EXOD|8|31|qui fecit iuxta verbum illius et abstulit muscas a Pharao et a servis et a populo eius non superfuit ne una quidem
EXOD|8|32|et ingravatum est cor Pharaonis ita ut ne hac quidem vice dimitteret populum
EXOD|9|1|dixit autem Dominus ad Mosen ingredere ad Pharaonem et loquere ad eum haec dicit Dominus Deus Hebraeorum dimitte populum meum ut sacrificet mihi
EXOD|9|2|quod si adhuc rennuis et retines eos
EXOD|9|3|ecce manus mea erit super agros tuos et super equos et asinos et camelos et boves et oves pestis valde gravis
EXOD|9|4|et faciet Dominus mirabile inter possessiones Israhel et possessiones Aegyptiorum ut nihil omnino intereat ex his quae pertinent ad filios Israhel
EXOD|9|5|constituitque Dominus tempus dicens cras faciet Dominus verbum istud in terra
EXOD|9|6|fecit ergo Dominus verbum hoc altero die mortuaque sunt omnia animantia Aegyptiorum de animalibus vero filiorum Israhel nihil omnino periit
EXOD|9|7|et misit Pharao ad videndum nec erat quicquam mortuum de his quae possidebat Israhel ingravatumque est cor Pharaonis et non dimisit populum
EXOD|9|8|et dixit Dominus ad Mosen et Aaron tollite plenas manus cineris de camino et spargat illud Moses in caelum coram Pharao
EXOD|9|9|sitque pulvis super omnem terram Aegypti erunt enim in hominibus et in iumentis vulnera et vesicae turgentes in universa terra Aegypti
EXOD|9|10|tuleruntque cinerem de camino et steterunt contra Pharao et sparsit illud Moses in caelum factaque sunt vulnera vesicarum turgentium in hominibus et in iumentis
EXOD|9|11|nec poterant malefici stare coram Mosen propter vulnera quae in illis erant et in omni terra Aegypti
EXOD|9|12|induravitque Dominus cor Pharaonis et non audivit eos sicut locutus est Dominus ad Mosen
EXOD|9|13|dixit quoque Dominus ad Mosen mane consurge et sta coram Pharao et dices ad eum haec dicit Dominus Deus Hebraeorum dimitte populum meum ut sacrificet mihi
EXOD|9|14|quia in hac vice mittam omnes plagas meas super cor tuum super servos tuos et super populum tuum ut scias quod non sit similis mei in omni terra
EXOD|9|15|nunc enim extendens manum percutiam te et populum tuum peste peribisque de terra
EXOD|9|16|idcirco autem posui te ut ostendam in te fortitudinem meam et narretur nomen meum in omni terra
EXOD|9|17|adhuc retines populum meum et non vis eum dimittere
EXOD|9|18|en pluam hac ipsa hora cras grandinem multam nimis qualis non fuit in Aegypto a die qua fundata est usque in praesens tempus
EXOD|9|19|mitte ergo iam nunc et congrega iumenta tua et omnia quae habes in agro homines enim et iumenta et universa quae inventa fuerint foris nec congregata de agris cecideritque super ea grando morientur
EXOD|9|20|qui timuit verbum Domini de servis Pharao fecit confugere servos suos et iumenta in domos
EXOD|9|21|qui autem neglexit sermonem Domini dimisit servos suos et iumenta in agris
EXOD|9|22|et dixit Dominus ad Mosen extende manum tuam in caelum ut fiat grando in universa terra Aegypti super homines et super iumenta et super omnem herbam agri in terra Aegypti
EXOD|9|23|extenditque Moses virgam in caelum et Dominus dedit tonitrua et grandinem ac discurrentia fulgura super terram pluitque Dominus grandinem super terram Aegypti
EXOD|9|24|et grando et ignis inmixta pariter ferebantur tantaeque fuit magnitudinis quanta ante numquam apparuit in universa terra Aegypti ex quo gens illa condita est
EXOD|9|25|et percussit grando in omni terra Aegypti cuncta quae fuerunt in agris ab homine usque ad iumentum cunctam herbam agri percussit grando et omne lignum regionis confregit
EXOD|9|26|tantum in terra Gessen ubi erant filii Israhel grando non cecidit
EXOD|9|27|misitque Pharao et vocavit Mosen et Aaron dicens ad eos peccavi etiam nunc Dominus iustus ego et populus meus impii
EXOD|9|28|orate Dominum et desinant tonitrua Dei et grando ut dimittam vos et nequaquam hic ultra maneatis
EXOD|9|29|ait Moses cum egressus fuero de urbe extendam palmas meas ad Dominum et cessabunt tonitrua et grando non erit ut scias quia Domini est terra
EXOD|9|30|novi autem quod et tu et servi tui necdum timeatis Dominum Deum
EXOD|9|31|linum ergo et hordeum laesum est eo quod hordeum esset virens et linum iam folliculos germinaret
EXOD|9|32|triticum autem et far non sunt laesa quia serotina erant
EXOD|9|33|egressusque Moses a Pharaone et ex urbe tetendit manus ad Dominum et cessaverunt tonitrua et grando nec ultra stillavit pluvia super terram
EXOD|9|34|videns autem Pharao quod cessasset pluvia et grando et tonitrua auxit peccatum
EXOD|9|35|et ingravatum est cor eius et servorum illius et induratum nimis nec dimisit filios Israhel sicut praeceperat Dominus per manum Mosi
EXOD|10|1|et dixit Dominus ad Mosen ingredere ad Pharao ego enim induravi cor eius et servorum illius ut faciam signa mea haec in eo
EXOD|10|2|et narres in auribus filii tui et nepotum tuorum quotiens contriverim Aegyptios et signa mea fecerim in eis et sciatis quia ego Dominus
EXOD|10|3|introierunt ergo Moses et Aaron ad Pharaonem et dixerunt ad eum haec dicit Dominus Deus Hebraeorum usquequo non vis subici mihi dimitte populum meum ut sacrificet mihi
EXOD|10|4|sin autem resistis et non vis dimittere eum ecce ego inducam cras lucustam in fines tuos
EXOD|10|5|quae operiat superficiem terrae nec quicquam eius appareat sed comedatur quod residuum fuit grandini conrodet enim omnia ligna quae germinant in agris
EXOD|10|6|et implebunt domos tuas et servorum tuorum et omnium Aegyptiorum quantam non viderunt patres tui et avi ex quo orti sunt super terram usque in praesentem diem avertitque se et egressus est a Pharaone
EXOD|10|7|dixerunt autem servi Pharaonis ad eum usquequo patiemur hoc scandalum dimitte homines ut sacrificent Domino Deo suo nonne vides quod perierit Aegyptus
EXOD|10|8|revocaveruntque Mosen et Aaron ad Pharaonem qui dixit eis ite sacrificate Domino Deo vestro quinam sunt qui ituri sunt
EXOD|10|9|ait Moses cum parvulis nostris et senibus pergemus cum filiis et filiabus cum ovibus et armentis est enim sollemnitas Domini nostri
EXOD|10|10|et respondit sic Dominus sit vobiscum quomodo ego dimittam vos et parvulos vestros cui dubium est quod pessime cogitetis
EXOD|10|11|non fiet ita sed ite tantum viri et sacrificate Domino hoc enim et ipsi petistis statimque eiecti sunt de conspectu Pharaonis
EXOD|10|12|dixit autem Dominus ad Mosen extende manum tuam super terram Aegypti ad lucustam ut ascendat super eam et devoret omnem herbam quae residua fuit grandini
EXOD|10|13|extendit Moses virgam super terram Aegypti et Dominus induxit ventum urentem tota illa die ac nocte et mane facto ventus urens levavit lucustas
EXOD|10|14|quae ascenderunt super universam terram Aegypti et sederunt in cunctis finibus Aegyptiorum innumerabiles quales ante illud tempus non fuerant nec postea futurae sunt
EXOD|10|15|operueruntque universam superficiem terrae vastantes omnia devorata est igitur herba terrae et quicquid pomorum in arboribus fuit quae grando dimiserat nihilque omnino virens relictum est in lignis et in herbis terrae in cuncta Aegypto
EXOD|10|16|quam ob rem festinus Pharao vocavit Mosen et Aaron et dixit eis peccavi in Dominum Deum vestrum et in vos
EXOD|10|17|sed nunc dimittite peccatum mihi etiam hac vice et rogate Dominum Deum vestrum ut auferat a me mortem istam
EXOD|10|18|egressusque est de conspectu Pharaonis et oravit Dominum
EXOD|10|19|qui flare fecit ventum ab occidente vehementissimum et arreptam lucustam proiecit in mare Rubrum non remansit ne una quidem in cunctis finibus Aegypti
EXOD|10|20|et induravit Dominus cor Pharaonis nec dimisit filios Israhel
EXOD|10|21|dixit autem Dominus ad Mosen extende manum tuam in caelum et sint tenebrae super terram Aegypti tam densae ut palpari queant
EXOD|10|22|extendit Moses manum in caelum et factae sunt tenebrae horribiles in universa terra Aegypti tribus diebus
EXOD|10|23|nemo vidit fratrem suum nec movit se de loco in quo erat ubicumque autem habitabant filii Israhel lux erat
EXOD|10|24|vocavitque Pharao Mosen et Aaron et dixit eis ite sacrificate Domino oves tantum vestrae et armenta remaneant parvuli vestri eant vobiscum
EXOD|10|25|ait Moses hostias quoque et holocausta dabis nobis quae offeramus Domino Deo nostro
EXOD|10|26|cuncti greges pergent nobiscum non remanebit ex eis ungula quae necessaria sunt in cultum Domini Dei nostri praesertim cum ignoremus quid debeat immolari donec ad ipsum locum perveniamus
EXOD|10|27|induravit autem Dominus cor Pharaonis et noluit dimittere eos
EXOD|10|28|dixitque Pharao ad eum recede a me cave ne ultra videas faciem meam quocumque die apparueris mihi morieris
EXOD|10|29|respondit Moses ita fiat ut locutus es non videbo ultra faciem tuam
EXOD|11|1|et dixit Dominus ad Mosen adhuc una plaga tangam Pharaonem et Aegyptum et post haec dimittet vos et exire conpellet
EXOD|11|2|dices ergo omni plebi ut postulet vir ab amico suo et mulier a vicina sua vasa argentea et aurea
EXOD|11|3|dabit autem Dominus gratiam populo coram Aegyptiis fuitque Moses vir magnus valde in terra Aegypti coram servis Pharao et omni populo
EXOD|11|4|et ait haec dicit Dominus media nocte egrediar in Aegyptum
EXOD|11|5|et morietur omne primogenitum in terra Aegyptiorum a primogenito Pharaonis qui sedet in solio eius usque ad primogenitum ancillae quae est ad molam et omnia primogenita iumentorum
EXOD|11|6|eritque clamor magnus in universa terra Aegypti qualis nec ante fuit nec postea futurus est
EXOD|11|7|apud omnes autem filios Israhel non muttiet canis ab homine usque ad pecus ut sciatis quanto miraculo dividat Dominus Aegyptios et Israhel
EXOD|11|8|descendentque omnes servi tui isti ad me et adorabunt me dicentes egredere tu et omnis populus qui subiectus est tibi post haec egrediemur
EXOD|11|9|et exivit a Pharaone iratus nimis dixit autem Dominus ad Mosen non audiet vos Pharao ut multa signa fiant in terra Aegypti
EXOD|11|10|Moses autem et Aaron fecerunt omnia ostenta quae scripta sunt coram Pharaone et induravit Dominus cor Pharaonis nec dimisit filios Israhel de terra sua
EXOD|12|1|dixit quoque Dominus ad Mosen et Aaron in terra Aegypti
EXOD|12|2|mensis iste vobis principium mensuum primus erit in mensibus anni
EXOD|12|3|loquimini ad universum coetum filiorum Israhel et dicite eis decima die mensis huius tollat unusquisque agnum per familias et domos suas
EXOD|12|4|sin autem minor est numerus ut sufficere possit ad vescendum agnum adsumet vicinum suum qui iunctus est domui eius iuxta numerum animarum quae sufficere possunt ad esum agni
EXOD|12|5|erit autem agnus absque macula masculus anniculus iuxta quem ritum tolletis et hedum
EXOD|12|6|et servabitis eum usque ad quartamdecimam diem mensis huius immolabitque eum universa multitudo filiorum Israhel ad vesperam
EXOD|12|7|et sument de sanguine ac ponent super utrumque postem et in superliminaribus domorum in quibus comedent illum
EXOD|12|8|et edent carnes nocte illa assas igni et azymos panes cum lactucis agrestibus
EXOD|12|9|non comedetis ex eo crudum quid nec coctum aqua sed assum tantum igni caput cum pedibus eius et intestinis vorabitis
EXOD|12|10|nec remanebit ex eo quicquam usque mane si quid residui fuerit igne conburetis
EXOD|12|11|sic autem comedetis illum renes vestros accingetis calciamenta habebitis in pedibus tenentes baculos in manibus et comedetis festinantes est enim phase id est transitus Domini
EXOD|12|12|et transibo per terram Aegypti nocte illa percutiamque omne primogenitum in terra Aegypti ab homine usque ad pecus et in cunctis diis Aegypti faciam iudicia ego Dominus
EXOD|12|13|erit autem sanguis vobis in signum in aedibus in quibus eritis et videbo sanguinem ac transibo vos nec erit in vobis plaga disperdens quando percussero terram Aegypti
EXOD|12|14|habebitis autem hanc diem in monumentum et celebrabitis eam sollemnem Domino in generationibus vestris cultu sempiterno
EXOD|12|15|septem diebus azyma comedetis in die primo non erit fermentum in domibus vestris quicumque comederit fermentatum peribit anima illa de Israhel a primo die usque ad diem septimum
EXOD|12|16|dies prima erit sancta atque sollemnis et dies septima eadem festivitate venerabilis nihil operis facietis in eis exceptis his quae ad vescendum pertinent
EXOD|12|17|et observabitis azyma in eadem enim ipsa die educam exercitum vestrum de terra Aegypti et custodietis diem istum in generationes vestras ritu perpetuo
EXOD|12|18|primo mense quartadecima die mensis ad vesperam comedetis azyma usque ad diem vicesimam primam eiusdem mensis ad vesperam
EXOD|12|19|septem diebus fermentum non invenietur in domibus vestris qui comederit fermentatum peribit anima eius de coetu Israhel tam de advenis quam de indigenis terrae
EXOD|12|20|omne fermentatum non comedetis in cunctis habitaculis vestris edetis azyma
EXOD|12|21|vocavit autem Moses omnes seniores filiorum Israhel et dixit ad eos ite tollentes animal per familias vestras immolate phase
EXOD|12|22|fasciculumque hysopi tinguite sanguine qui est in limine et aspergite ex eo superliminare et utrumque postem nullus vestrum egrediatur ostium domus suae usque mane
EXOD|12|23|transibit enim Dominus percutiens Aegyptios cumque viderit sanguinem in superliminari et in utroque poste transcendet ostium et non sinet percussorem ingredi domos vestras et laedere
EXOD|12|24|custodi verbum istud legitimum tibi et filiis tuis usque in aeternum
EXOD|12|25|cumque introieritis terram quam Dominus daturus est vobis ut pollicitus est observabitis caerimonias istas
EXOD|12|26|et cum dixerint vobis filii vestri quae est ista religio
EXOD|12|27|dicetis eis victima transitus Domini est quando transivit super domos filiorum Israhel in Aegypto percutiens Aegyptios et domos nostras liberans incurvatusque populus adoravit
EXOD|12|28|et egressi filii Israhel fecerunt sicut praeceperat Dominus Mosi et Aaron
EXOD|12|29|factum est autem in noctis medio percussit Dominus omne primogenitum in terra Aegypti a primogenito Pharaonis qui sedebat in solio eius usque ad primogenitum captivae quae erat in carcere et omne primogenitum iumentorum
EXOD|12|30|surrexitque Pharao nocte et omnes servi eius cunctaque Aegyptus et ortus est clamor magnus in Aegypto neque enim erat domus in qua non iaceret mortuus
EXOD|12|31|vocatisque Mosen et Aaron nocte ait surgite egredimini a populo meo et vos et filii Israhel ite immolate Domino sicut dicitis
EXOD|12|32|oves vestras et armenta adsumite ut petieratis et abeuntes benedicite mihi
EXOD|12|33|urguebantque Aegyptii populum de terra exire velociter dicentes omnes moriemur
EXOD|12|34|tulit igitur populus conspersam farinam antequam fermentaretur et ligans in palliis posuit super umeros suos
EXOD|12|35|feceruntque filii Israhel sicut praeceperat Moses et petierunt ab Aegyptiis vasa argentea et aurea vestemque plurimam
EXOD|12|36|dedit autem Dominus gratiam populo coram Aegyptiis ut commodarent eis et spoliaverunt Aegyptios
EXOD|12|37|profectique sunt filii Israhel de Ramesse in Soccoth sescenta ferme milia peditum virorum absque parvulis
EXOD|12|38|sed et vulgus promiscuum innumerabile ascendit cum eis oves et armenta et animantia diversi generis multa nimis
EXOD|12|39|coxeruntque farinam quam dudum conspersam de Aegypto tulerant et fecerunt subcinericios panes azymos neque enim poterant fermentari cogentibus exire Aegyptiis et nullam facere sinentibus moram nec pulmenti quicquam occurrerant praeparare
EXOD|12|40|habitatio autem filiorum Israhel qua manserant in Aegypto fuit quadringentorum triginta annorum
EXOD|12|41|quibus expletis eadem die egressus est omnis exercitus Domini de terra Aegypti
EXOD|12|42|nox est ista observabilis Domini quando eduxit eos de terra Aegypti hanc observare debent omnes filii Israhel in generationibus suis
EXOD|12|43|dixitque Dominus ad Mosen et Aaron haec est religio phase omnis alienigena non comedet ex eo
EXOD|12|44|omnis autem servus empticius circumcidetur et sic comedet
EXOD|12|45|advena et mercennarius non edent ex eo
EXOD|12|46|in una domo comedetur nec efferetis de carnibus eius foras nec os illius confringetis
EXOD|12|47|omnis coetus filiorum Israhel faciet illud
EXOD|12|48|quod si quis peregrinorum in vestram voluerit transire coloniam et facere phase Domini circumcidetur prius omne masculinum eius et tunc rite celebrabit eritque sicut indigena terrae si quis autem circumcisus non fuerit non vescetur ex eo
EXOD|12|49|eadem lex erit indigenae et colono qui peregrinatur apud vos
EXOD|12|50|fecerunt omnes filii Israhel sicut praeceperat Dominus Mosi et Aaron
EXOD|12|51|et in eadem die eduxit Dominus filios Israhel de terra Aegypti per turmas suas
EXOD|13|1|locutusque est Dominus ad Mosen dicens
EXOD|13|2|sanctifica mihi omne primogenitum quod aperit vulvam in filiis Israhel tam de hominibus quam de iumentis mea sunt enim omnia
EXOD|13|3|et ait Moses ad populum mementote diei huius in qua egressi estis de Aegypto et de domo servitutis quoniam in manu forti eduxit vos Dominus de loco isto ut non comedatis fermentatum panem
EXOD|13|4|hodie egredimini mense novarum frugum
EXOD|13|5|cumque te introduxerit Dominus in terram Chananei et Hetthei et Amorrei et Evei et Iebusei quam iuravit patribus tuis ut daret tibi terram fluentem lacte et melle celebrabis hunc morem sacrorum mense isto
EXOD|13|6|septem diebus vesceris azymis et in die septimo erit sollemnitas Domini
EXOD|13|7|azyma comedetis septem diebus non apparebit apud te aliquid fermentatum nec in cunctis finibus tuis
EXOD|13|8|narrabisque filio tuo in die illo dicens hoc est quod fecit Dominus mihi quando egressus sum de Aegypto
EXOD|13|9|et erit quasi signum in manu tua et quasi monumentum ante oculos tuos et ut lex Domini semper in ore tuo in manu enim forti eduxit te Dominus de Aegypto
EXOD|13|10|custodies huiuscemodi cultum statuto tempore a diebus in dies
EXOD|13|11|cumque introduxerit te in terram Chananei sicut iuravit tibi et patribus tuis et dederit eam tibi
EXOD|13|12|separabis omne quod aperit vulvam Domino et quod primitivum est in pecoribus tuis quicquid habueris masculini sexus consecrabis Domino
EXOD|13|13|primogenitum asini mutabis ove quod si non redemeris interficies omne autem primogenitum hominis de filiis tuis pretio redimes
EXOD|13|14|cumque interrogaverit te filius tuus cras dicens quid est hoc respondebis ei in manu forti eduxit nos Dominus de Aegypto de domo servitutis
EXOD|13|15|nam cum induratus esset Pharao et nollet nos dimittere occidit Dominus omne primogenitum in terra Aegypti a primogenito hominis usque ad primogenitum iumentorum idcirco immolo Domino omne quod aperit vulvam masculini sexus et omnia primogenita filiorum meorum redimo
EXOD|13|16|erit igitur quasi signum in manu tua et quasi adpensum quid ob recordationem inter oculos tuos eo quod in manu forti eduxerit nos Dominus de Aegypto
EXOD|13|17|igitur cum emisisset Pharao populum non eos duxit Dominus per viam terrae Philisthim quae vicina est reputans ne forte paeniteret eum si vidisset adversum se bella consurgere et reverteretur in Aegyptum
EXOD|13|18|sed circumduxit per viam deserti quae est iuxta mare Rubrum et armati ascenderunt filii Israhel de terra Aegypti
EXOD|13|19|tulit quoque Moses ossa Ioseph secum eo quod adiurasset filios Israhel dicens visitabit vos Deus efferte ossa mea hinc vobiscum
EXOD|13|20|profectique de Soccoth castrametati sunt in Etham in extremis finibus solitudinis
EXOD|13|21|Dominus autem praecedebat eos ad ostendendam viam per diem in columna nubis et per noctem in columna ignis ut dux esset itineris utroque tempore
EXOD|13|22|numquam defuit columna nubis per diem nec columna ignis per noctem coram populo
EXOD|14|1|locutus est autem Dominus ad Mosen dicens
EXOD|14|2|loquere filiis Israhel reversi castrametentur e regione Phiahiroth quae est inter Magdolum et mare contra Beelsephon in conspectu eius castra ponetis super mare
EXOD|14|3|dicturusque est Pharao super filiis Israhel coartati sunt in terra conclusit eos desertum
EXOD|14|4|et indurabo cor eius ac persequetur vos et glorificabor in Pharao et in omni exercitu eius scientque Aegyptii quia ego sum Dominus feceruntque ita
EXOD|14|5|et nuntiatum est regi Aegyptiorum quod fugisset populus inmutatumque est cor Pharaonis et servorum eius super populo et dixerunt quid voluimus facere ut dimitteremus Israhel ne serviret nobis
EXOD|14|6|iunxit ergo currum et omnem populum suum adsumpsit secum
EXOD|14|7|tulitque sescentos currus electos quicquid in Aegypto curruum fuit et duces totius exercitus
EXOD|14|8|induravitque Dominus cor Pharaonis regis Aegypti et persecutus est filios Israhel at illi egressi erant in manu excelsa
EXOD|14|9|cumque persequerentur Aegyptii vestigia praecedentium reppererunt eos in castris super mare omnis equitatus et currus Pharaonis et universus exercitus erant in Ahiroth contra Beelsephon
EXOD|14|10|cumque adpropinquasset Pharao levantes filii Israhel oculos viderunt Aegyptios post se et timuerunt valde clamaveruntque ad Dominum
EXOD|14|11|et dixerunt ad Mosen forsitan non erant sepulchra in Aegypto ideo tulisti nos ut moreremur in solitudine quid hoc facere voluisti ut educeres nos ex Aegypto
EXOD|14|12|nonne iste est sermo quem loquebamur ad te in Aegypto dicentes recede a nobis ut serviamus Aegyptiis multo enim melius est servire eis quam mori in solitudine
EXOD|14|13|et ait Moses ad populum nolite timere state et videte magnalia Domini quae facturus est hodie Aegyptios enim quos nunc videtis nequaquam ultra videbitis usque in sempiternum
EXOD|14|14|Dominus pugnabit pro vobis et vos tacebitis
EXOD|14|15|dixitque Dominus ad Mosen quid clamas ad me loquere filiis Israhel ut proficiscantur
EXOD|14|16|tu autem eleva virgam tuam et extende manum super mare et divide illud ut gradiantur filii Israhel in medio mari per siccum
EXOD|14|17|ego autem indurabo cor Aegyptiorum ut persequantur vos et glorificabor in Pharaone et in omni exercitu eius in curribus et in equitibus illius
EXOD|14|18|et scient Aegyptii quia ego sum Dominus cum glorificatus fuero in Pharaone et in curribus atque in equitibus eius
EXOD|14|19|tollensque se angelus Dei qui praecedebat castra Israhel abiit post eos et cum eo pariter columna nubis priora dimittens post tergum
EXOD|14|20|stetit inter castra Aegyptiorum et castra Israhel et erat nubes tenebrosa et inluminans noctem ut ad se invicem toto noctis tempore accedere non valerent
EXOD|14|21|cumque extendisset Moses manum super mare abstulit illud Dominus flante vento vehementi et urente tota nocte et vertit in siccum divisaque est aqua
EXOD|14|22|et ingressi sunt filii Israhel per medium maris sicci erat enim aqua quasi murus a dextra eorum et leva
EXOD|14|23|persequentesque Aegyptii ingressi sunt post eos omnis equitatus Pharaonis currus eius et equites per medium maris
EXOD|14|24|iamque advenerat vigilia matutina et ecce respiciens Dominus super castra Aegyptiorum per columnam ignis et nubis interfecit exercitum eorum
EXOD|14|25|et subvertit rotas curruum ferebanturque in profundum dixerunt ergo Aegyptii fugiamus Israhelem Dominus enim pugnat pro eis contra nos
EXOD|14|26|et ait Dominus ad Mosen extende manum tuam super mare ut revertantur aquae ad Aegyptios super currus et equites eorum
EXOD|14|27|cumque extendisset Moses manum contra mare reversum est primo diluculo ad priorem locum fugientibusque Aegyptiis occurrerunt aquae et involvit eos Dominus in mediis fluctibus
EXOD|14|28|reversaeque sunt aquae et operuerunt currus et equites cuncti exercitus Pharaonis qui sequentes ingressi fuerant mare ne unus quidem superfuit ex eis
EXOD|14|29|filii autem Israhel perrexerunt per medium sicci maris et aquae eis erant quasi pro muro a dextris et a sinistris
EXOD|14|30|liberavitque Dominus in die illo Israhel de manu Aegyptiorum
EXOD|14|31|et viderunt Aegyptios mortuos super litus maris et manum magnam quam exercuerat Dominus contra eos timuitque populus Dominum et crediderunt Domino et Mosi servo eius
EXOD|15|1|tunc cecinit Moses et filii Israhel carmen hoc Domino et dixerunt cantemus Domino gloriose enim magnificatus est equum et ascensorem deiecit in mare
EXOD|15|2|fortitudo mea et laus mea Dominus et factus est mihi in salutem iste Deus meus et glorificabo eum Deus patris mei et exaltabo eum
EXOD|15|3|Dominus quasi vir pugnator Omnipotens nomen eius
EXOD|15|4|currus Pharaonis et exercitum eius proiecit in mare electi principes eius submersi sunt in mari Rubro
EXOD|15|5|abyssi operuerunt eos descenderunt in profundum quasi lapis
EXOD|15|6|dextera tua Domine magnifice in fortitudine dextera tua Domine percussit inimicum
EXOD|15|7|et in multitudine gloriae tuae deposuisti adversarios meos misisti iram tuam quae devoravit eos ut stipulam
EXOD|15|8|et in spiritu furoris tui congregatae sunt aquae stetit unda fluens congregatae sunt abyssi in medio mari
EXOD|15|9|dixit inimicus persequar et conprehendam dividam spolia implebitur anima mea evaginabo gladium meum interficiet eos manus mea
EXOD|15|10|flavit spiritus tuus et operuit eos mare submersi sunt quasi plumbum in aquis vehementibus
EXOD|15|11|quis similis tui in fortibus Domine quis similis tui magnificus in sanctitate terribilis atque laudabilis et faciens mirabilia
EXOD|15|12|extendisti manum tuam et devoravit eos terra
EXOD|15|13|dux fuisti in misericordia tua populo quem redemisti et portasti eum in fortitudine tua ad habitaculum sanctum tuum
EXOD|15|14|adtenderunt populi et irati sunt dolores obtinuerunt habitatores Philisthim
EXOD|15|15|tunc conturbati sunt principes Edom robustos Moab obtinuit tremor obriguerunt omnes habitatores Chanaan
EXOD|15|16|inruat super eos formido et pavor in magnitudine brachii tui fiant inmobiles quasi lapis donec pertranseat populus tuus Domine donec pertranseat populus tuus iste quem possedisti
EXOD|15|17|introduces eos et plantabis in monte hereditatis tuae firmissimo habitaculo tuo quod operatus es Domine sanctuarium Domine quod firmaverunt manus tuae
EXOD|15|18|Dominus regnabit in aeternum et ultra
EXOD|15|19|ingressus est enim equus Pharao cum curribus et equitibus eius in mare et reduxit super eos Dominus aquas maris filii autem Israhel ambulaverunt per siccum in medio eius
EXOD|15|20|sumpsit ergo Maria prophetis soror Aaron tympanum in manu egressaeque sunt omnes mulieres post eam cum tympanis et choris
EXOD|15|21|quibus praecinebat dicens cantemus Domino gloriose enim magnificatus est equum et ascensorem eius deiecit in mare
EXOD|15|22|tulit autem Moses Israhel de mari Rubro et egressi sunt in desertum Sur ambulaveruntque tribus diebus per solitudinem et non inveniebant aquam
EXOD|15|23|et venerunt in Marath nec poterant bibere aquas de Mara eo quod essent amarae unde et congruum loco nomen inposuit vocans illud Mara id est amaritudinem
EXOD|15|24|et murmuravit populus contra Mosen dicens quid bibemus
EXOD|15|25|at ille clamavit ad Dominum qui ostendit ei lignum quod cum misisset in aquas in dulcedinem versae sunt ibi constituit ei praecepta atque iudicia et ibi temptavit eum
EXOD|15|26|dicens si audieris vocem Domini Dei tui et quod rectum est coram eo feceris et oboedieris mandatis eius custodierisque omnia praecepta illius cunctum languorem quem posui in Aegypto non inducam super te ego enim Dominus sanator tuus
EXOD|15|27|venerunt autem in Helim ubi erant duodecim fontes aquarum et septuaginta palmae et castrametati sunt iuxta aquas
EXOD|16|1|profectique sunt de Helim et venit omnis multitudo filiorum Israhel in desertum Sin quod est inter Helim et Sinai quintodecimo die mensis secundi postquam egressi sunt de terra Aegypti
EXOD|16|2|et murmuravit omnis congregatio filiorum Israhel contra Mosen et contra Aaron in solitudine
EXOD|16|3|dixeruntque ad eos filii Israhel utinam mortui essemus per manum Domini in terra Aegypti quando sedebamus super ollas carnium et comedebamus panes in saturitate cur eduxistis nos in desertum istud ut occideretis omnem multitudinem fame
EXOD|16|4|dixit autem Dominus ad Mosen ecce ego pluam vobis panes de caelo egrediatur populus et colligat quae sufficiunt per singulos dies ut temptem eum utrum ambulet in lege mea an non
EXOD|16|5|die autem sexta parent quod inferant et sit duplum quam colligere solebant per singulos dies
EXOD|16|6|dixeruntque Moses et Aaron ad omnes filios Israhel vespere scietis quod Dominus eduxerit vos de terra Aegypti
EXOD|16|7|et mane videbitis gloriam Domini audivit enim murmur vestrum contra Dominum nos vero quid sumus quia mussitatis contra nos
EXOD|16|8|et ait Moses dabit Dominus vobis vespere carnes edere et mane panes in saturitate eo quod audierit murmurationes vestras quibus murmurati estis contra eum nos enim quid sumus nec contra nos est murmur vestrum sed contra Dominum
EXOD|16|9|dixitque Moses ad Aaron dic universae congregationi filiorum Israhel accedite coram Domino audivit enim murmur vestrum
EXOD|16|10|cumque loqueretur Aaron ad omnem coetum filiorum Israhel respexerunt ad solitudinem et ecce gloria Domini apparuit in nube
EXOD|16|11|locutus est autem Dominus ad Mosen dicens
EXOD|16|12|audivi murmurationes filiorum Israhel loquere ad eos vespere comedetis carnes et mane saturabimini panibus scietisque quod sim Dominus Deus vester
EXOD|16|13|factum est ergo vespere et ascendens coturnix operuit castra mane quoque ros iacuit per circuitum castrorum
EXOD|16|14|cumque operuisset superficiem terrae apparuit in solitudine minutum et quasi pilo tunsum in similitudinem pruinae super terram
EXOD|16|15|quod cum vidissent filii Israhel dixerunt ad invicem man hu quod significat quid est hoc ignorabant enim quid esset quibus ait Moses iste est panis quem dedit Dominus vobis ad vescendum
EXOD|16|16|hic est sermo quem praecepit Dominus colligat ex eo unusquisque quantum sufficiat ad vescendum gomor per singula capita iuxta numerum animarum vestrarum quae habitant in tabernaculo sic tolletis
EXOD|16|17|feceruntque ita filii Israhel et collegerunt alius plus alius minus
EXOD|16|18|et mensi sunt ad mensuram gomor nec qui plus collegerat habuit amplius nec qui minus paraverat repperit minus sed singuli iuxta id quod edere poterant congregarunt
EXOD|16|19|dixitque Moses ad eos nullus relinquat ex eo in mane
EXOD|16|20|qui non audierunt eum sed dimiserunt quidam ex eis usque mane et scatere coepit vermibus atque conputruit et iratus est contra eos Moses
EXOD|16|21|colligebant autem mane singuli quantum sufficere poterat ad vescendum cumque incaluisset sol liquefiebat
EXOD|16|22|in die vero sexta collegerunt cibos duplices id est duo gomor per singulos homines venerunt autem omnes principes multitudinis et narraverunt Mosi
EXOD|16|23|qui ait eis hoc est quod locutus est Dominus requies sabbati sanctificata erit Domino cras quodcumque operandum est facite et quae coquenda sunt coquite quicquid autem reliquum fuerit reponite usque in mane
EXOD|16|24|feceruntque ita ut praeceperat Moses et non conputruit neque vermis inventus est in eo
EXOD|16|25|dixitque Moses comedite illud hodie quia sabbatum est Domino non invenietur hodie in agro
EXOD|16|26|sex diebus colligite in die autem septimo sabbatum est Domino idcirco non invenietur
EXOD|16|27|venit septima dies et egressi de populo ut colligerent non invenerunt
EXOD|16|28|dixit autem Dominus ad Mosen usquequo non vultis custodire mandata mea et legem meam
EXOD|16|29|videte quod Dominus dederit vobis sabbatum et propter hoc tribuerit vobis die sexto cibos duplices maneat unusquisque apud semet ipsum nullus egrediatur de loco suo die septimo
EXOD|16|30|et sabbatizavit populus die septimo
EXOD|16|31|appellavitque domus Israhel nomen eius man quod erat quasi semen coriandri album gustusque eius quasi similae cum melle
EXOD|16|32|dixit autem Moses iste est sermo quem praecepit Dominus imple gomor ex eo et custodiatur in futuras retro generationes ut noverint panem quo alui vos in solitudine quando educti estis de terra Aegypti
EXOD|16|33|dixitque Moses ad Aaron sume vas unum et mitte ibi man quantum potest capere gomor et repone coram Domino ad servandum in generationes vestras
EXOD|16|34|sicut praecepit Dominus Mosi posuitque illud Aaron in tabernaculo reservandum
EXOD|16|35|filii autem Israhel comederunt man quadraginta annis donec venirent in terram habitabilem hoc cibo aliti sunt usquequo tangerent fines terrae Chanaan
EXOD|16|36|gomor autem decima pars est oephi
EXOD|17|1|igitur profecta omnis multitudo filiorum Israhel de deserto Sin per mansiones suas iuxta sermonem Domini castrametata est in Raphidim ubi non erat aqua ad bibendum populo
EXOD|17|2|qui iurgatus contra Mosen ait da nobis aquam ut bibamus quibus respondit Moses quid iurgamini contra me cur temptatis Dominum
EXOD|17|3|sitivit ergo populus ibi pro aquae penuria et murmuravit contra Mosen dicens cur nos exire fecisti de Aegypto ut occideres et nos et liberos nostros ac iumenta siti
EXOD|17|4|clamavit autem Moses ad Dominum dicens quid faciam populo huic adhuc pauxillum et lapidabunt me
EXOD|17|5|ait Dominus ad Mosen antecede populum et sume tecum de senibus Israhel et virgam qua percussisti fluvium tolle in manu tua et vade
EXOD|17|6|en ego stabo coram te ibi super petram Horeb percutiesque petram et exibit ex ea aqua ut bibat populus fecit Moses ita coram senibus Israhel
EXOD|17|7|et vocavit nomen loci illius Temptatio propter iurgium filiorum Israhel et quia temptaverunt Dominum dicentes estne Dominus in nobis an non
EXOD|17|8|venit autem Amalech et pugnabat contra Israhel in Raphidim
EXOD|17|9|dixitque Moses ad Iosue elige viros et egressus pugna contra Amalech cras ego stabo in vertice collis habens virgam Dei in manu mea
EXOD|17|10|fecit Iosue ut locutus ei erat Moses et pugnavit contra Amalech Moses autem et Aaron et Hur ascenderunt super verticem collis
EXOD|17|11|cumque levaret Moses manus vincebat Israhel sin autem paululum remisisset superabat Amalech
EXOD|17|12|manus autem Mosi erant graves sumentes igitur lapidem posuerunt subter eum in quo sedit Aaron autem et Hur sustentabant manus eius ex utraque parte et factum est ut manus ipsius non lassarentur usque ad occasum solis
EXOD|17|13|fugavitque Iosue Amalech et populum eius in ore gladii
EXOD|17|14|dixit autem Dominus ad Mosen scribe hoc ob monumentum in libro et trade auribus Iosue delebo enim memoriam Amalech sub caelo
EXOD|17|15|aedificavitque Moses altare et vocavit nomen eius Dominus exaltatio mea dicens
EXOD|17|16|quia manus solii Domini et bellum Dei erit contra Amalech a generatione in generationem
EXOD|18|1|cumque audisset Iethro sacerdos Madian cognatus Mosi omnia quae fecerat Deus Mosi et Israhel populo suo eo quod eduxisset Dominus Israhel de Aegypto
EXOD|18|2|tulit Sefforam uxorem Mosi quam remiserat
EXOD|18|3|et duos filios eius quorum unus vocabatur Gersan dicente patre advena fui in terra aliena
EXOD|18|4|alter vero Eliezer Deus enim ait patris mei adiutor meus et eruit me de gladio Pharaonis
EXOD|18|5|venit ergo Iethro cognatus Mosi et filii eius et uxor ad Mosen in desertum ubi erat castrametatus iuxta montem Dei
EXOD|18|6|et mandavit Mosi dicens ego cognatus tuus Iethro venio ad te et uxor tua et duo filii tui cum ea
EXOD|18|7|qui egressus in occursum cognati sui adoravit et osculatus est eum salutaveruntque se mutuo verbis pacificis cumque intrasset tabernaculum
EXOD|18|8|narravit Moses cognato suo cuncta quae fecerat Deus Pharaoni et Aegyptiis propter Israhel universum laborem qui accidisset eis in itinere quo liberarat eos Dominus
EXOD|18|9|laetatusque est Iethro super omnibus bonis quae fecerat Dominus Israheli eo quod eruisset eum de manu Aegyptiorum
EXOD|18|10|et ait benedictus Dominus qui liberavit vos de manu Aegyptiorum et de manu Pharaonis qui eruit populum suum de manu Aegypti
EXOD|18|11|nunc cognovi quia magnus Dominus super omnes deos eo quod superbe egerint contra illos
EXOD|18|12|obtulit ergo Iethro cognatus Mosi holocausta et hostias Deo veneruntque Aaron et omnes senes Israhel ut comederent panem cum eo coram Domino
EXOD|18|13|altero autem die sedit Moses ut iudicaret populum qui adsistebat Mosi de mane usque ad vesperam
EXOD|18|14|quod cum vidisset cognatus eius omnia scilicet quae agebat in populo ait quid est hoc quod facis in plebe cur solus sedes et omnis populus praestolatur de mane usque ad vesperam
EXOD|18|15|cui respondit Moses venit ad me populus quaerens sententiam Dei
EXOD|18|16|cumque acciderit eis aliqua disceptatio veniunt ad me ut iudicem inter eos et ostendam praecepta Dei et leges eius
EXOD|18|17|at ille non bonam inquit rem facis
EXOD|18|18|stulto labore consumeris et tu et populus iste qui tecum est ultra vires tuas est negotium solus illud non poteris sustinere
EXOD|18|19|sed audi verba mea atque consilia et erit Deus tecum esto tu populo in his quae ad Deum pertinent ut referas quae dicuntur ad eum
EXOD|18|20|ostendasque populo caerimonias et ritum colendi viamque per quam ingredi debeant et opus quod facere
EXOD|18|21|provide autem de omni plebe viros potentes et timentes Deum in quibus sit veritas et qui oderint avaritiam et constitue ex eis tribunos et centuriones et quinquagenarios et decanos
EXOD|18|22|qui iudicent populum omni tempore quicquid autem maius fuerit referant ad te et ipsi minora tantummodo iudicent leviusque tibi sit partito in alios onere
EXOD|18|23|si hoc feceris implebis imperium Dei et praecepta eius poteris sustentare et omnis hic populus revertetur cum pace ad loca sua
EXOD|18|24|quibus auditis Moses fecit omnia quae ille suggesserat
EXOD|18|25|et electis viris strenuis de cuncto Israhel constituit eos principes populi tribunos et centuriones et quinquagenarios et decanos
EXOD|18|26|qui iudicabant plebem omni tempore quicquid autem gravius erat referebant ad eum faciliora tantummodo iudicantes
EXOD|18|27|dimisitque cognatum qui reversus abiit in terram suam
EXOD|19|1|mense tertio egressionis Israhel de terra Aegypti in die hac venerunt in solitudinem Sinai
EXOD|19|2|nam profecti de Raphidim et pervenientes usque in desertum Sinai castrametati sunt in eodem loco ibique Israhel fixit tentoria e regione montis
EXOD|19|3|Moses autem ascendit ad Deum vocavitque eum Dominus de monte et ait haec dices domui Iacob et adnuntiabis filiis Israhel
EXOD|19|4|vos ipsi vidistis quae fecerim Aegyptiis quomodo portaverim vos super alas aquilarum et adsumpserim mihi
EXOD|19|5|si ergo audieritis vocem meam et custodieritis pactum meum eritis mihi in peculium de cunctis populis mea est enim omnis terra
EXOD|19|6|et vos eritis mihi regnum sacerdotale et gens sancta haec sunt verba quae loqueris ad filios Israhel
EXOD|19|7|venit Moses et convocatis maioribus natu populi exposuit omnes sermones quos mandaverat Dominus
EXOD|19|8|responditque universus populus simul cuncta quae locutus est Dominus faciemus cumque rettulisset Moses verba populi ad Dominum
EXOD|19|9|ait ei Dominus iam nunc veniam ad te in caligine nubis ut audiat me populus loquentem ad te et credat tibi in perpetuum nuntiavit ergo Moses verba populi ad Dominum
EXOD|19|10|qui dixit ei vade ad populum et sanctifica illos hodie et cras laventque vestimenta sua
EXOD|19|11|et sint parati in diem tertium die enim tertio descendet Dominus coram omni plebe super montem Sinai
EXOD|19|12|constituesque terminos populo per circuitum et dices cavete ne ascendatis in montem nec tangatis fines illius omnis qui tetigerit montem morte morietur
EXOD|19|13|manus non tanget eum sed lapidibus opprimetur aut confodietur iaculis sive iumentum fuerit sive homo non vivet cum coeperit clangere bucina tunc ascendant in montem
EXOD|19|14|descenditque Moses de monte ad populum et sanctificavit eum cumque lavissent vestimenta sua
EXOD|19|15|ait ad eos estote parati in diem tertium ne adpropinquetis uxoribus vestris
EXOD|19|16|iam advenerat tertius dies et mane inclaruerat et ecce coeperunt audiri tonitrua ac micare fulgura et nubes densissima operire montem clangorque bucinae vehementius perstrepebat timuit populus qui erat in castris
EXOD|19|17|cumque eduxisset eos Moses in occursum Dei de loco castrorum steterunt ad radices montis
EXOD|19|18|totus autem mons Sinai fumabat eo quod descendisset Dominus super eum in igne et ascenderet fumus ex eo quasi de fornace eratque mons omnis terribilis
EXOD|19|19|et sonitus bucinae paulatim crescebat in maius et prolixius tendebatur Moses loquebatur et Dominus respondebat ei
EXOD|19|20|descenditque Dominus super montem Sinai in ipso montis vertice et vocavit Mosen in cacumen eius quo cum ascendisset
EXOD|19|21|dixit ad eum descende et contestare populum ne forte velint transcendere terminos ad videndum Dominum et pereat ex eis plurima multitudo
EXOD|19|22|sacerdotes quoque qui accedunt ad Dominum sanctificentur ne percutiat eos
EXOD|19|23|dixitque Moses ad Dominum non poterit vulgus ascendere in montem Sinai tu enim testificatus es et iussisti dicens pone terminos circa montem et sanctifica illum
EXOD|19|24|cui ait Dominus vade descende ascendesque tu et Aaron tecum sacerdotes autem et populus ne transeant terminos nec ascendant ad Dominum ne forte interficiat illos
EXOD|19|25|descendit Moses ad populum et omnia narravit eis
EXOD|20|1|locutus quoque est Dominus cunctos sermones hos
EXOD|20|2|ego sum Dominus Deus tuus qui eduxi te de terra Aegypti de domo servitutis
EXOD|20|3|non habebis deos alienos coram me
EXOD|20|4|non facies tibi sculptile neque omnem similitudinem quae est in caelo desuper et quae in terra deorsum nec eorum quae sunt in aquis sub terra
EXOD|20|5|non adorabis ea neque coles ego sum Dominus Deus tuus fortis zelotes visitans iniquitatem patrum in filiis in tertiam et quartam generationem eorum qui oderunt me
EXOD|20|6|et faciens misericordiam in milia his qui diligunt me et custodiunt praecepta mea
EXOD|20|7|non adsumes nomen Domini Dei tui in vanum nec enim habebit insontem Dominus eum qui adsumpserit nomen Domini Dei sui frustra
EXOD|20|8|memento ut diem sabbati sanctifices
EXOD|20|9|sex diebus operaberis et facies omnia opera tua
EXOD|20|10|septimo autem die sabbati Domini Dei tui non facies omne opus tu et filius tuus et filia tua servus tuus et ancilla tua iumentum tuum et advena qui est intra portas tuas
EXOD|20|11|sex enim diebus fecit Dominus caelum et terram et mare et omnia quae in eis sunt et requievit in die septimo idcirco benedixit Dominus diei sabbati et sanctificavit eum
EXOD|20|12|honora patrem tuum et matrem tuam ut sis longevus super terram quam Dominus Deus tuus dabit tibi
EXOD|20|13|non occides
EXOD|20|14|non moechaberis
EXOD|20|15|non furtum facies
EXOD|20|16|non loqueris contra proximum tuum falsum testimonium
EXOD|20|17|non concupisces domum proximi tui nec desiderabis uxorem eius non servum non ancillam non bovem non asinum nec omnia quae illius sunt
EXOD|20|18|cunctus autem populus videbat voces et lampadas et sonitum bucinae montemque fumantem et perterriti ac pavore concussi steterunt procul
EXOD|20|19|dicentes Mosi loquere tu nobis et audiemus non loquatur nobis Dominus ne forte moriamur
EXOD|20|20|et ait Moses ad populum nolite timere ut enim probaret vos venit Deus et ut terror illius esset in vobis et non peccaretis
EXOD|20|21|stetitque populus de longe Moses autem accessit ad caliginem in qua erat Deus
EXOD|20|22|dixit praeterea Dominus ad Mosen haec dices filiis Israhel vos vidistis quod de caelo locutus sum vobis
EXOD|20|23|non facietis mecum deos argenteos nec deos aureos facietis vobis
EXOD|20|24|altare de terra facietis mihi et offeretis super eo holocausta et pacifica vestra oves vestras et boves in omni loco in quo memoria fuerit nominis mei veniam ad te et benedicam tibi
EXOD|20|25|quod si altare lapideum feceris mihi non aedificabis illud de sectis lapidibus si enim levaveris cultrum tuum super eo polluetur
EXOD|20|26|non ascendes per gradus ad altare meum ne reveletur turpitudo tua
EXOD|21|1|haec sunt iudicia quae propones eis
EXOD|21|2|si emeris servum hebraeum sex annis serviet tibi in septimo egredietur liber gratis
EXOD|21|3|cum quali veste intraverit cum tali exeat si habens uxorem et uxor egredietur simul
EXOD|21|4|sin autem dominus dederit illi uxorem et peperit filios et filias mulier et liberi eius erunt domini sui ipse vero exibit cum vestitu suo
EXOD|21|5|quod si dixerit servus diligo dominum meum et uxorem ac liberos non egrediar liber
EXOD|21|6|offeret eum dominus diis et adplicabitur ad ostium et postes perforabitque aurem eius subula et erit ei servus in saeculum
EXOD|21|7|si quis vendiderit filiam suam in famulam non egredietur sicut ancillae exire consuerunt
EXOD|21|8|si displicuerit oculis domini sui cui tradita fuerit dimittet eam populo autem alieno vendendi non habet potestatem si spreverit eam
EXOD|21|9|sin autem filio suo desponderit eam iuxta morem filiarum faciet illi
EXOD|21|10|quod si alteram ei acceperit providebit puellae nuptias et vestimenta et pretium pudicitiae non negabit
EXOD|21|11|si tria ista non fecerit egredietur gratis absque pecunia
EXOD|21|12|qui percusserit hominem volens occidere morte moriatur
EXOD|21|13|qui autem non est insidiatus sed Deus illum tradidit in manu eius constituam tibi locum quo fugere debeat
EXOD|21|14|si quis de industria occiderit proximum suum et per insidias ab altari meo evelles eum ut moriatur
EXOD|21|15|qui percusserit patrem suum et matrem morte moriatur
EXOD|21|16|qui furatus fuerit hominem et vendiderit eum convictus noxae morte moriatur
EXOD|21|17|qui maledixerit patri suo et matri morte moriatur
EXOD|21|18|si rixati fuerint viri et percusserit alter proximum suum lapide vel pugno et ille mortuus non fuerit sed iacuerit in lectulo
EXOD|21|19|si surrexerit et ambulaverit foris super baculum suum innocens erit qui percussit ita tamen ut operas eius et inpensas in medicos restituat
EXOD|21|20|qui percusserit servum suum vel ancillam virga et mortui fuerint in manibus eius criminis reus erit
EXOD|21|21|sin autem uno die supervixerit vel duobus non subiacebit poenae quia pecunia illius est
EXOD|21|22|si rixati fuerint viri et percusserit quis mulierem praegnantem et abortivum quidem fecerit sed ipsa vixerit subiacebit damno quantum expetierit maritus mulieris et arbitri iudicarint
EXOD|21|23|sin autem mors eius fuerit subsecuta reddet animam pro anima
EXOD|21|24|oculum pro oculo dentem pro dente manum pro manu pedem pro pede
EXOD|21|25|adustionem pro adustione vulnus pro vulnere livorem pro livore
EXOD|21|26|si percusserit quispiam oculum servi sui aut ancillae et luscos eos fecerit dimittet liberos pro oculo quem eruit
EXOD|21|27|dentem quoque si excusserit servo vel ancillae suae similiter dimittet eos liberos
EXOD|21|28|si bos cornu petierit virum aut mulierem et mortui fuerint lapidibus obruetur et non comedentur carnes eius dominusque bovis innocens erit
EXOD|21|29|quod si bos cornipeta fuerit ab heri et nudius tertius et contestati sunt dominum eius nec reclusit eum occideritque virum aut mulierem et bos lapidibus obruetur et dominum illius occident
EXOD|21|30|quod si pretium ei fuerit inpositum dabit pro anima sua quicquid fuerit postulatus
EXOD|21|31|filium quoque et filiam si cornu percusserit simili sententiae subiacebit
EXOD|21|32|si servum ancillamque invaserit triginta siclos argenti dabit domino bos vero lapidibus opprimetur
EXOD|21|33|si quis aperuerit cisternam et foderit et non operuerit eam cecideritque bos vel asinus in eam
EXOD|21|34|dominus cisternae reddet pretium iumentorum quod autem mortuum est ipsius erit
EXOD|21|35|si bos alienus bovem alterius vulnerarit et ille mortuus fuerit vendent bovem vivum et divident pretium cadaver autem mortui inter se dispertient
EXOD|21|36|sin autem sciebat quod bos cornipeta esset ab heri et nudius tertius et non custodivit eum dominus suus reddet bovem pro bove et cadaver integrum accipiet
EXOD|22|1|si quis furatus fuerit bovem aut ovem et occiderit vel vendiderit quinque boves pro uno bove restituet et quattuor oves pro una ove
EXOD|22|2|si effringens fur domum sive suffodiens fuerit inventus et accepto vulnere mortuus fuerit percussor non erit reus sanguinis
EXOD|22|3|quod si orto sole hoc fecerit homicidium perpetravit et ipse morietur si non habuerit quod pro furto reddat venundabitur
EXOD|22|4|si inventum fuerit apud eum quod furatus est vivens sive bos sive asinus sive ovis duplum restituet
EXOD|22|5|si laeserit quispiam agrum vel vineam et dimiserit iumentum suum ut depascatur aliena quicquid optimum habuerit in agro suo vel in vinea pro damni aestimatione restituet
EXOD|22|6|si egressus ignis invenerit spinas et conprehenderit acervos frugum sive stantes segetes in agris reddet damnum qui ignem succenderit
EXOD|22|7|si quis commendaverit amico pecuniam aut vas in custodiam et ab eo qui susceperat furto ablata fuerint si invenitur fur duplum reddet
EXOD|22|8|si latet dominus domus adplicabitur ad deos et iurabit quod non extenderit manum in rem proximi sui
EXOD|22|9|ad perpetrandam fraudem tam in bove quam in asino et ove ac vestimento et quicquid damnum inferre potest ad deos utriusque causa perveniet et si illi iudicaverint duplum restituet proximo suo
EXOD|22|10|si quis commendaverit proximo suo asinum bovem ovem et omne iumentum ad custodiam et mortuum fuerit aut debilitatum vel captum ab hostibus nullusque hoc viderit
EXOD|22|11|iusiurandum erit in medio quod non extenderit manum ad rem proximi sui suscipietque dominus iuramentum et ille reddere non cogetur
EXOD|22|12|quod si furto ablatum fuerit restituet damnum domino
EXOD|22|13|si comestum a bestia deferet ad eum quod occisum est et non restituet
EXOD|22|14|qui a proximo suo quicquam horum mutuo postularit et debilitatum aut mortuum fuerit domino non praesente reddere conpelletur
EXOD|22|15|quod si inpraesentiarum fuit dominus non restituet maxime si conductum venerat pro mercede operis sui
EXOD|22|16|si seduxerit quis virginem necdum desponsatam et dormierit cum ea dotabit eam et habebit uxorem
EXOD|22|17|si pater virginis dare noluerit reddet pecuniam iuxta modum dotis quam virgines accipere consuerunt
EXOD|22|18|maleficos non patieris vivere
EXOD|22|19|qui coierit cum iumento morte moriatur
EXOD|22|20|qui immolat diis occidetur praeter Domino soli
EXOD|22|21|advenam non contristabis neque adfliges eum advenae enim et ipsi fuistis in terra Aegypti
EXOD|22|22|viduae et pupillo non nocebitis
EXOD|22|23|si laeseritis eos vociferabuntur ad me et ego audiam clamorem eorum
EXOD|22|24|et indignabitur furor meus percutiamque vos gladio et erunt uxores vestrae viduae et filii vestri pupilli
EXOD|22|25|si pecuniam mutuam dederis populo meo pauperi qui habitat tecum non urgues eum quasi exactor nec usuris opprimes
EXOD|22|26|si pignus a proximo tuo acceperis vestimentum ante solis occasum redde ei
EXOD|22|27|ipsum enim est solum quo operitur indumentum carnis eius nec habet aliud in quo dormiat si clamaverit ad me exaudiam eum quia misericors sum
EXOD|22|28|diis non detrahes et principi populi tui non maledices
EXOD|22|29|decimas tuas et primitias non tardabis offerre primogenitum filiorum tuorum dabis mihi
EXOD|22|30|de bubus quoque et ovibus similiter facies septem diebus sit cum matre sua die octavo reddes illum mihi
EXOD|22|31|viri sancti eritis mihi carnem quae a bestiis fuerit praegustata non comedetis sed proicietis canibus
EXOD|23|1|non suscipies vocem mendacii nec iunges manum tuam ut pro impio dicas falsum testimonium
EXOD|23|2|non sequeris turbam ad faciendum malum nec in iudicio plurimorum adquiesces sententiae ut a vero devies
EXOD|23|3|pauperis quoque non misereberis in negotio
EXOD|23|4|si occurreris bovi inimici tui aut asino erranti reduc ad eum
EXOD|23|5|si videris asinum odientis te iacere sub onere non pertransibis sed sublevabis cum eo
EXOD|23|6|non declinabis in iudicio pauperis
EXOD|23|7|mendacium fugies insontem et iustum non occides quia aversor impium
EXOD|23|8|nec accipias munera quae excaecant etiam prudentes et subvertunt verba iustorum
EXOD|23|9|peregrino molestus non eris scitis enim advenarum animas quia et ipsi peregrini fuistis in terra Aegypti
EXOD|23|10|sex annis seminabis terram tuam et congregabis fruges eius
EXOD|23|11|anno autem septimo dimittes eam et requiescere facies ut comedant pauperes populi tui et quicquid reliqui fuerit edant bestiae agri ita facies in vinea et in oliveto tuo
EXOD|23|12|sex diebus operaberis septima die cessabis ut requiescat bos et asinus tuus et refrigeretur filius ancillae tuae et advena
EXOD|23|13|omnia quae dixi vobis custodite et per nomen externorum deorum non iurabitis neque audietur ex ore vestro
EXOD|23|14|tribus vicibus per singulos annos mihi festa celebrabitis
EXOD|23|15|sollemnitatem azymorum custodies septem diebus comedes azyma sicut praecepi tibi tempore mensis novorum quando egressus es de Aegypto non apparebis in conspectu meo vacuus
EXOD|23|16|et sollemnitatem messis primitivorum operis tui quaecumque serueris in agro sollemnitatem quoque in exitu anni quando congregaveris omnes fruges tuas de agro
EXOD|23|17|ter in anno apparebit omne masculinum tuum coram Domino Deo
EXOD|23|18|non immolabis super fermento sanguinem victimae meae nec remanebit adeps sollemnitatis meae usque mane
EXOD|23|19|primitias frugum terrae tuae deferes in domum Domini Dei tui nec coques hedum in lacte matris suae
EXOD|23|20|ecce ego mittam angelum meum qui praecedat te et custodiat in via et introducat ad locum quem paravi
EXOD|23|21|observa eum et audi vocem eius nec contemnendum putes quia non dimittet cum peccaveritis et est nomen meum in illo
EXOD|23|22|quod si audieris vocem eius et feceris omnia quae loquor inimicus ero inimicis tuis et adfligam adfligentes te
EXOD|23|23|praecedetque te angelus meus et introducet te ad Amorreum et Hettheum et Ferezeum Chananeumque et Eveum et Iebuseum quos ego contribo
EXOD|23|24|non adorabis deos eorum nec coles eos non facies opera eorum sed destrues eos et confringes statuas eorum
EXOD|23|25|servietisque Domino Deo vestro ut benedicam panibus tuis et aquis et auferam infirmitatem de medio tui
EXOD|23|26|non erit infecunda nec sterilis in terra tua numerum dierum tuorum implebo
EXOD|23|27|terrorem meum mittam in praecursum tuum et occidam omnem populum ad quem ingredieris cunctorumque inimicorum tuorum coram te terga vertam
EXOD|23|28|emittens crabrones prius qui fugabunt Eveum et Chananeum et Hettheum antequam introeas
EXOD|23|29|non eiciam eos a facie tua anno uno ne terra in solitudinem redigatur et crescant contra te bestiae
EXOD|23|30|paulatim expellam eos de conspectu tuo donec augearis et possideas terram
EXOD|23|31|ponam autem terminos tuos a mari Rubro usque ad mare Palestinorum et a deserto usque ad Fluvium tradam manibus vestris habitatores terrae et eiciam eos de conspectu vestro
EXOD|23|32|non inibis cum eis foedus nec cum diis eorum
EXOD|23|33|non habitent in terra tua ne forte peccare te faciant in me si servieris diis eorum quod tibi certo erit in scandalum
EXOD|24|1|Mosi quoque dixit ascende ad Dominum tu et Aaron Nadab et Abiu et septuaginta senes ex Israhel et adorabitis procul
EXOD|24|2|solusque Moses ascendet ad Dominum et illi non adpropinquabunt nec populus ascendet cum eo
EXOD|24|3|venit ergo Moses et narravit plebi omnia verba Domini atque iudicia responditque cunctus populus una voce omnia verba Domini quae locutus est faciemus
EXOD|24|4|scripsit autem Moses universos sermones Domini et mane consurgens aedificavit altare ad radices montis et duodecim titulos per duodecim tribus Israhel
EXOD|24|5|misitque iuvenes de filiis Israhel et obtulerunt holocausta immolaveruntque victimas pacificas Domino vitulos
EXOD|24|6|tulit itaque Moses dimidiam partem sanguinis et misit in crateras partem autem residuam fudit super altare
EXOD|24|7|adsumensque volumen foederis legit audiente populo qui dixerunt omnia quae locutus est Dominus faciemus et erimus oboedientes
EXOD|24|8|ille vero sumptum sanguinem respersit in populum et ait hic est sanguis foederis quod pepigit Dominus vobiscum super cunctis sermonibus his
EXOD|24|9|ascenderuntque Moses et Aaron Nadab et Abiu et septuaginta de senioribus Israhel
EXOD|24|10|et viderunt Deum Israhel sub pedibus eius quasi opus lapidis sapphirini et quasi caelum cum serenum est
EXOD|24|11|nec super eos qui procul recesserant de filiis Israhel misit manum suam videruntque Deum et comederunt ac biberunt
EXOD|24|12|dixit autem Dominus ad Mosen ascende ad me in montem et esto ibi daboque tibi tabulas lapideas et legem ac mandata quae scripsi ut doceas eos
EXOD|24|13|surrexerunt Moses et Iosue minister eius ascendensque Moses in montem Dei
EXOD|24|14|senioribus ait expectate hic donec revertamur ad vos habetis Aaron et Hur vobiscum si quid natum fuerit quaestionis referetis ad eos
EXOD|24|15|cumque ascendisset Moses operuit nubes montem
EXOD|24|16|et habitavit gloria Domini super Sinai tegens illum nube sex diebus septimo autem die vocavit eum de medio caliginis
EXOD|24|17|erat autem species gloriae Domini quasi ignis ardens super verticem montis in conspectu filiorum Israhel
EXOD|24|18|ingressusque Moses medium nebulae ascendit in montem et fuit ibi quadraginta diebus et quadraginta noctibus
EXOD|25|1|locutusque est Dominus ad Mosen dicens
EXOD|25|2|loquere filiis Israhel ut tollant mihi primitias ab omni homine qui offert ultroneus accipietis eas
EXOD|25|3|haec sunt autem quae accipere debetis aurum et argentum et aes
EXOD|25|4|hyacinthum et purpuram coccumque bis tinctum et byssum pilos caprarum
EXOD|25|5|et pelles arietum rubricatas pelles ianthinas et ligna setthim
EXOD|25|6|oleum ad luminaria concinnanda aromata in unguentum et thymiama boni odoris
EXOD|25|7|lapides onychinos et gemmas ad ornandum ephod ac rationale
EXOD|25|8|facientque mihi sanctuarium et habitabo in medio eorum
EXOD|25|9|iuxta omnem similitudinem tabernaculi quod ostendam tibi et omnium vasorum in cultum eius sicque facietis illud
EXOD|25|10|arcam de lignis setthim conpingite cuius longitudo habeat duos semis cubitos latitudo cubitum et dimidium altitudo cubitum similiter ac semissem
EXOD|25|11|et deaurabis eam auro mundissimo intus et foris faciesque supra coronam auream per circuitum
EXOD|25|12|et quattuor circulos aureos quos pones per quattuor arcae angulos duo circuli sint in latere uno et duo in altero
EXOD|25|13|facies quoque vectes de lignis setthim et operies eos auro
EXOD|25|14|inducesque per circulos qui sunt in arcae lateribus ut portetur in eis
EXOD|25|15|qui semper erunt in circulis nec umquam extrahentur ab eis
EXOD|25|16|ponesque in arcam testificationem quam dabo tibi
EXOD|25|17|facies et propitiatorium de auro mundissimo duos cubitos et dimidium tenebit longitudo eius cubitum ac semissem latitudo
EXOD|25|18|duos quoque cherubin aureos et productiles facies ex utraque parte oraculi
EXOD|25|19|cherub unus sit in latere uno et alter in altero
EXOD|25|20|utrumque latus propitiatorii tegant expandentes alas et operientes oraculum respiciantque se mutuo versis vultibus in propitiatorium quo operienda est arca
EXOD|25|21|in qua pones testimonium quod dabo tibi
EXOD|25|22|inde praecipiam et loquar ad te supra propitiatorio scilicet ac medio duorum cherubin qui erunt super arcam testimonii cuncta quae mandabo per te filiis Israhel
EXOD|25|23|facies et mensam de lignis setthim habentem duos cubitos longitudinis et in latitudine cubitum et in altitudine cubitum ac semissem
EXOD|25|24|et inaurabis eam auro purissimo faciesque illi labium aureum per circuitum
EXOD|25|25|et ipsi labio coronam interrasilem altam quattuor digitis et super illam alteram coronam aureolam
EXOD|25|26|quattuor quoque circulos aureos praeparabis et pones eos in quattuor angulis eiusdem mensae per singulos pedes
EXOD|25|27|subter coronam erunt circuli aurei ut mittantur vectes per eos et possit mensa portari
EXOD|25|28|ipsosque vectes facies de lignis setthim et circumdabis auro ad subvehendam mensam
EXOD|25|29|parabis et acetabula ac fialas turibula et cyatos in quibus offerenda sunt libamina ex auro purissimo
EXOD|25|30|et pones super mensam panes propositionis in conspectu meo semper
EXOD|25|31|facies et candelabrum ductile de auro mundissimo hastile eius et calamos scyphos et spherulas ac lilia ex ipso procedentia
EXOD|25|32|sex calami egredientur de lateribus tres ex uno latere et tres ex altero
EXOD|25|33|tres scyphi quasi in nucis modum per calamos singulos spherulaque simul et lilium et tres similiter scyphi instar nucis in calamo altero spherulaque et lilium hoc erit opus sex calamorum qui producendi sunt de hastili
EXOD|25|34|in ipso autem candelabro erunt quattuor scyphi in nucis modum spherulaeque per singulos et lilia
EXOD|25|35|spherula sub duobus calamis per tria loca qui simul sex fiunt procedentes de hastili uno
EXOD|25|36|et spherae igitur et calami ex ipso erunt universa ductilia de auro purissimo
EXOD|25|37|facies et lucernas septem et pones eas super candelabrum ut luceant ex adverso
EXOD|25|38|emunctoria quoque et ubi quae emuncta sunt extinguantur fient de auro purissimo
EXOD|25|39|omne pondus candelabri cum universis vasis suis habebit talentum auri mundissimi
EXOD|25|40|inspice et fac secundum exemplar quod tibi in monte monstratum est
EXOD|26|1|tabernaculum vero ita fiet decem cortinas de bysso retorta et hyacintho ac purpura coccoque bis tincto variatas opere plumario facies
EXOD|26|2|longitudo cortinae unius habebit viginti octo cubitos latitudo quattuor cubitorum erit unius mensurae fient universa tentoria
EXOD|26|3|quinque cortinae sibi iungentur mutuo et aliae quinque nexu simili coherebunt
EXOD|26|4|ansulas hyacinthinas in lateribus ac summitatibus facies cortinarum ut possint invicem copulari
EXOD|26|5|quinquagenas ansulas cortina habebit in utraque parte ita insertas ut ansa contra ansam veniat et altera alteri possit aptari
EXOD|26|6|facies et quinquaginta circulos aureos quibus cortinarum vela iungenda sunt ut unum tabernaculum fiat
EXOD|26|7|facies et saga cilicina undecim ad operiendum tectum tabernaculi
EXOD|26|8|longitudo sagi unius habebit triginta cubitos et latitudo quattuor aequa erit mensura sagorum omnium
EXOD|26|9|e quibus quinque iunges seorsum et sex sibi mutuo copulabis ita ut sextum sagum in fronte tecti duplices
EXOD|26|10|facies et quinquaginta ansas in ora sagi unius ut coniungi cum altero queat et quinquaginta ansas in ora sagi alterius ut cum altero copuletur
EXOD|26|11|quinquaginta fibulas aeneas quibus iungantur ansae et unum ex omnibus operimentum fiat
EXOD|26|12|quod autem superfuerit in sagis quae parantur tecto id est unum sagum quod amplius est ex medietate eius operies posteriora tabernaculi
EXOD|26|13|et cubitus ex una parte pendebit et alter ex altera qui plus est in sagorum longitudine utrumque latus tabernaculi protegens
EXOD|26|14|facies et operimentum aliud tecto de pellibus arietum rubricatis et super hoc rursum aliud operimentum de ianthinis pellibus
EXOD|26|15|facies et tabulas stantes tabernaculi de lignis setthim
EXOD|26|16|quae singulae denos cubitos in longitudine habeant et in latitudine singulos ac semissem
EXOD|26|17|in lateribus tabulae duae incastraturae fient quibus tabula alteri tabulae conectatur atque in hunc modum cunctae tabulae parabuntur
EXOD|26|18|quarum viginti erunt in latere meridiano quod vergit ad austrum
EXOD|26|19|quibus quadraginta bases argenteas fundes ut binae bases singulis tabulis per duos angulos subiciantur
EXOD|26|20|in latere quoque secundo tabernaculi quod vergit ad aquilonem viginti tabulae erunt
EXOD|26|21|quadraginta habentes bases argenteas binae bases singulis tabulis subponentur
EXOD|26|22|ad occidentalem vero plagam tabernaculi facies sex tabulas
EXOD|26|23|et rursum alias duas quae in angulis erigantur post tergum tabernaculi
EXOD|26|24|eruntque coniunctae a deorsum usque sursum et una omnes conpago retinebit duabus quoque tabulis quae in angulis ponendae sunt similis iunctura servabitur
EXOD|26|25|et erunt simul tabulae octo bases earum argenteae sedecim duabus basibus per unam tabulam supputatis
EXOD|26|26|facies et vectes de lignis setthim quinque ad continendas tabulas in uno latere tabernaculi
EXOD|26|27|et quinque alios in altero et eiusdem numeri ad occidentalem plagam
EXOD|26|28|qui mittentur per medias tabulas a summo usque ad summum
EXOD|26|29|ipsasque tabulas deaurabis et fundes eis anulos aureos per quos vectes tabulata contineant quos operies lamminis aureis
EXOD|26|30|et eriges tabernaculum iuxta exemplum quod tibi in monte monstratum est
EXOD|26|31|facies et velum de hyacintho et purpura coccoque bis tincto et bysso retorta opere plumario et pulchra varietate contextum
EXOD|26|32|quod adpendes ante quattuor columnas de lignis setthim quae ipsae quidem deauratae erunt et habebunt capita aurea sed bases argenteas
EXOD|26|33|inseretur autem velum per circulos intra quod pones arcam testimonii et quo sanctuarium et sanctuarii sanctuaria dividentur
EXOD|26|34|pones et propitiatorium super arcam testimonii in sancta sanctorum
EXOD|26|35|mensamque extra velum et contra mensam candelabrum in latere tabernaculi meridiano mensa enim stabit in parte aquilonis
EXOD|26|36|facies et tentorium in introitu tabernaculi de hyacintho et purpura coccoque bis tincto et bysso retorta opere plumarii
EXOD|26|37|et quinque columnas deaurabis lignorum setthim ante quas ducetur tentorium quarum erunt capita aurea et bases aeneae
EXOD|27|1|facies et altare de lignis setthim quod habebit quinque cubitos in longitudine et totidem in latitudine id est quadrum et tres cubitos in altitudine
EXOD|27|2|cornua autem per quattuor angulos ex ipso erunt et operies illud aere
EXOD|27|3|faciesque in usus eius lebetas ad suscipiendos cineres et forcipes atque fuscinulas et ignium receptacula omnia vasa ex aere fabricabis
EXOD|27|4|craticulamque in modum retis aeneam per cuius quattuor angulos erunt quattuor anuli aenei
EXOD|27|5|quos pones subter arulam altaris eritque craticula usque ad altaris medium
EXOD|27|6|facies et vectes altaris de lignis setthim duos quos operies lamminis aeneis
EXOD|27|7|et induces per circulos eruntque ex utroque latere altaris ad portandum
EXOD|27|8|non solidum sed inane et cavum intrinsecus facies illud sicut tibi in monte monstratum est
EXOD|27|9|facies et atrium tabernaculi in cuius plaga australi contra meridiem erunt tentoria de bysso retorta centum cubitos unum latus tenebit in longitudine
EXOD|27|10|et columnas viginti cum basibus totidem aeneis quae capita cum celaturis suis habebunt argentea
EXOD|27|11|similiter in latere aquilonis per longum erunt tentoria centum cubitorum columnae viginti et bases aeneae eiusdem numeri et capita earum cum celaturis suis argentea
EXOD|27|12|in latitudine vero atrii quod respicit ad occidentem erunt tentoria per quinquaginta cubitos et columnae decem basesque totidem
EXOD|27|13|in ea quoque atrii latitudine quae respicit ad orientem quinquaginta cubiti erunt
EXOD|27|14|in quibus quindecim cubitorum tentoria lateri uno deputabuntur columnaeque tres et bases totidem
EXOD|27|15|et in latere altero erunt tentoria cubitos obtinentia quindecim columnas tres et bases totidem
EXOD|27|16|in introitu vero atrii fiet tentorium cubitorum viginti ex hyacintho et purpura coccoque bis tincto et bysso retorta opere plumarii columnas habebit quattuor cum basibus totidem
EXOD|27|17|omnes columnae atrii per circuitum vestitae erunt argenti lamminis capitibus argenteis et basibus aeneis
EXOD|27|18|in longitudine occupabit atrium cubitos centum in latitudine quinquaginta altitudo quinque cubitorum erit fietque de bysso retorta et habebit bases aeneas
EXOD|27|19|cuncta vasa tabernaculi in omnes usus et caerimonias tam paxillos eius quam atrii ex aere facies
EXOD|27|20|praecipe filiis Israhel ut adferant tibi oleum de arboribus olivarum purissimum piloque contusum ut ardeat lucerna semper
EXOD|27|21|in tabernaculo testimonii extra velum quod oppansum est testimonio et conlocabunt eam Aaron et filii eius ut usque mane luceat coram Domino perpetuus erit cultus per successiones eorum a filiis Israhel
EXOD|28|1|adplica quoque ad te Aaron fratrem tuum cum filiis suis de medio filiorum Israhel ut sacerdotio fungantur mihi Aaron Nadab et Abiu Eleazar et Ithamar
EXOD|28|2|faciesque vestem sanctam fratri tuo in gloriam et decorem
EXOD|28|3|et loqueris cunctis sapientibus corde quos replevi spiritu prudentiae ut faciant vestes Aaron in quibus sanctificatus ministret mihi
EXOD|28|4|haec autem erunt vestimenta quae facient rationale et superumerale tunicam et lineam strictam cidarim et balteum facient vestimenta sancta Aaron fratri tuo et filiis eius ut sacerdotio fungantur mihi
EXOD|28|5|accipientque aurum et hyacinthum et purpuram coccumque bis tinctum et byssum
EXOD|28|6|facient autem superumerale de auro et hyacintho ac purpura coccoque bis tincto et bysso retorta opere polymito
EXOD|28|7|duas oras iunctas habebit in utroque latere summitatum ut in unum redeant
EXOD|28|8|ipsaque textura et cuncta operis varietas erit ex auro et hyacintho et purpura coccoque bis tincto et bysso retorta
EXOD|28|9|sumesque duos lapides onychinos et sculpes in eis nomina filiorum Israhel
EXOD|28|10|sex nomina in lapide uno et sex reliqua in altero iuxta ordinem nativitatis eorum
EXOD|28|11|opere sculptoris et celatura gemmarii sculpes eos nominibus filiorum Israhel inclusos auro atque circumdatos
EXOD|28|12|et pones in utroque latere superumeralis memoriale filiis Israhel portabitque Aaron nomina eorum coram Domino super utrumque umerum ob recordationem
EXOD|28|13|facies et uncinos ex auro
EXOD|28|14|et duas catenulas auri purissimi sibi invicem coherentes quas inseres uncinis
EXOD|28|15|rationale quoque iudicii facies opere polymito iuxta texturam superumeralis ex auro hyacintho et purpura coccoque bis tincto et bysso retorta
EXOD|28|16|quadrangulum erit et duplex mensuram palmi habebit tam in longitudine quam in latitudine
EXOD|28|17|ponesque in eo quattuor ordines lapidum in primo versu erit lapis sardius et topazius et zmaragdus
EXOD|28|18|in secundo carbunculus sapphyrus et iaspis
EXOD|28|19|in tertio ligyrius achates et amethistus
EXOD|28|20|in quarto chrysolitus onychinus et berillus inclusi auro erunt per ordines suos
EXOD|28|21|habebuntque nomina filiorum Israhel duodecim nominibus celabuntur singuli lapides nominibus singulorum per duodecim tribus
EXOD|28|22|facies in rationali catenas sibi invicem coherentes ex auro purissimo
EXOD|28|23|et duos anulos aureos quos pones in utraque rationalis summitate
EXOD|28|24|catenasque aureas iunges anulis qui sunt in marginibus eius
EXOD|28|25|et ipsarum catenarum extrema duobus copulabis uncinis in utroque latere superumeralis quod rationale respicit
EXOD|28|26|facies et duos anulos aureos quos pones in summitatibus rationalis et in oris quae e regione sunt superumeralis et posteriora eius aspiciunt
EXOD|28|27|nec non et alios duos anulos aureos qui ponendi sunt in utroque latere superumeralis deorsum quod respicit contra faciem iuncturae inferioris ut aptari possit cum superumerali
EXOD|28|28|et stringatur rationale anulis suis cum anulis superumeralis vitta hyacinthina ut maneat iunctura fabrefacta et a se invicem rationale et superumerale nequeant separari
EXOD|28|29|portabitque Aaron nomina filiorum Israhel in rationali iudicii super pectus suum quando ingreditur sanctuarium memoriale coram Domino in aeternum
EXOD|28|30|pones autem in rationali iudicii doctrinam et veritatem quae erunt in pectore Aaron quando ingreditur coram Domino et gestabit iudicium filiorum Israhel in pectore suo in conspectu Domini semper
EXOD|28|31|facies et tunicam superumeralis totam hyacinthinam
EXOD|28|32|in cuius medio supra erit capitium et ora per gyrum eius textilis sicut fieri solet in extremis vestium partibus ne facile rumpatur
EXOD|28|33|deorsum vero ad pedes eiusdem tunicae per circuitum quasi mala punica facies ex hyacintho et purpura et cocco bis tincto mixtis in medio tintinabulis
EXOD|28|34|ita ut tintinabulum sit aureum et malum rursumque tintinabulum aliud aureum et malum punicum
EXOD|28|35|et vestietur ea Aaron in officio ministerii ut audiatur sonitus quando ingreditur et egreditur sanctuarium in conspectu Domini et non moriatur
EXOD|28|36|facies et lamminam de auro purissimo in qua sculpes opere celatoris Sanctum Domino
EXOD|28|37|ligabisque eam vitta hyacinthina et erit super tiaram
EXOD|28|38|inminens fronti pontificis portabitque Aaron iniquitates eorum quae obtulerint et sanctificaverint filii Israhel in cunctis muneribus et donariis suis erit autem lammina semper in fronte eius ut placatus eis sit Dominus
EXOD|28|39|stringesque tunicam bysso et tiaram byssinam facies et balteum opere plumarii
EXOD|28|40|porro filiis Aaron tunicas lineas parabis et balteos ac tiaras in gloriam et decorem
EXOD|28|41|vestiesque his omnibus Aaron fratrem tuum et filios eius cum eo et cunctorum consecrabis manus sanctificabisque illos ut sacerdotio fungantur mihi
EXOD|28|42|facies et feminalia linea ut operiant carnem turpitudinis suae a renibus usque ad femina
EXOD|28|43|et utentur eis Aaron et filii eius quando ingredientur tabernaculum testimonii vel quando adpropinquant ad altare ut ministrent in sanctuario ne iniquitatis rei moriantur legitimum sempiternum erit Aaron et semini eius post eum
EXOD|29|1|sed et hoc facies ut mihi in sacerdotio consecrentur tolle vitulum de armento et arietes duos inmaculatos
EXOD|29|2|panesque azymos et crustula absque fermento quae conspersa sint oleo lagana quoque azyma oleo lita de simila triticea cuncta facies
EXOD|29|3|et posita in canistro offeres vitulum autem et duos arietes
EXOD|29|4|et Aaron ac filios eius adplicabis ad ostium tabernaculi testimonii cumque laveris patrem cum filiis aqua
EXOD|29|5|indues Aaron vestimentis suis id est linea et tunica et superumerali et rationali quod constringes balteo
EXOD|29|6|et pones tiaram in capite eius et lamminam sanctam super tiaram
EXOD|29|7|et oleum unctionis fundes super caput eius atque hoc ritu consecrabitur
EXOD|29|8|filios quoque illius adplicabis et indues tunicis lineis cingesque balteo
EXOD|29|9|Aaron scilicet et liberos eius et inpones eis mitras eruntque sacerdotes mei in religione perpetua postquam initiaveris manus eorum
EXOD|29|10|adplicabis et vitulum coram tabernaculo testimonii inponentque Aaron et filii eius manus super caput illius
EXOD|29|11|et mactabis eum in conspectu Domini iuxta ostium tabernaculi testimonii
EXOD|29|12|sumptumque de sanguine vituli pones super cornua altaris digito tuo reliquum autem sanguinem fundes iuxta basim eius
EXOD|29|13|sumes et adipem totum qui operit intestina et reticulum iecoris ac duos renes et adipem qui super eos est et offeres incensum super altare
EXOD|29|14|carnes vero vituli et corium et fimum conbures foris extra castra eo quod pro peccato sit
EXOD|29|15|unum quoque arietum sumes super cuius caput ponent Aaron et filii eius manus
EXOD|29|16|quem cum mactaveris tolles de sanguine eius et fundes circa altare
EXOD|29|17|ipsum autem arietem secabis in frusta lotaque intestina eius ac pedes pones super concisas carnes et super caput illius
EXOD|29|18|et offeres totum arietem in incensum super altare oblatio est Domini odor suavissimus victimae Dei
EXOD|29|19|tolles quoque arietem alterum super cuius caput Aaron et filii eius ponent manus
EXOD|29|20|quem cum immolaveris sumes de sanguine ipsius et pones super extremum dextrae auriculae Aaron et filiorum eius et super pollices manus eorum et pedis dextri fundesque sanguinem super altare per circuitum
EXOD|29|21|cumque tuleris de sanguine qui est super altare et de oleo unctionis asperges Aaron et vestes eius filios et vestimenta eorum consecratisque et ipsis et vestibus
EXOD|29|22|tolles adipem de ariete et caudam et arvinam quae operit vitalia ac reticulum iecoris et duos renes atque adipem qui super eos est armumque dextrum eo quod sit aries consecrationum
EXOD|29|23|tortam panis unius crustulum conspersum oleo laganum de canistro azymorum quod positum est in conspectu Domini
EXOD|29|24|ponesque omnia super manus Aaron et filiorum eius et sanctificabis eos elevans coram Domino
EXOD|29|25|suscipiesque universa de manibus eorum et incendes super altare in holocaustum odorem suavissimum in conspectu Domini quia oblatio eius est
EXOD|29|26|sumes quoque pectusculum de ariete quo initiatus est Aaron sanctificabisque illud elatum coram Domino et cedet in partem tuam
EXOD|29|27|sanctificabis et pectusculum consecratum et armum quem de ariete separasti
EXOD|29|28|quo initiatus est Aaron et filii eius cedentque in partem Aaron et filiorum eius iure perpetuo a filiis Israhel quia primitiva sunt et initia de victimis eorum pacificis quae offerunt Domino
EXOD|29|29|vestem autem sanctam qua utitur Aaron habebunt filii eius post eum ut unguantur in ea et consecrentur manus eorum
EXOD|29|30|septem diebus utetur illa qui pontifex pro eo fuerit constitutus de filiis eius et qui ingredietur tabernaculum testimonii ut ministret in sanctuario
EXOD|29|31|arietem autem consecrationum tolles et coques carnes eius in loco sancto
EXOD|29|32|quibus vescetur Aaron et filii eius panes quoque qui sunt in canistro in vestibulo tabernaculi testimonii comedent
EXOD|29|33|ut sit placabile sacrificium et sanctificentur offerentium manus alienigena non vescetur ex eis quia sancti sunt
EXOD|29|34|quod si remanserit de carnibus consecratis sive de panibus usque mane conbures reliquias igni non comedentur quia sanctificata sunt
EXOD|29|35|omnia quae praecepi tibi facies super Aaron et filiis eius septem diebus consecrabis manus eorum
EXOD|29|36|et vitulum pro peccato offeres per singulos dies ad expiandum mundabisque altare cum immolaris expiationis hostiam et ungues illud in sanctificationem
EXOD|29|37|septem diebus expiabis altare et sanctificabis et erit sanctum sanctorum omnis qui tetigerit illud sanctificabitur
EXOD|29|38|hoc est quod facies in altari agnos anniculos duos per singulos dies iugiter
EXOD|29|39|unum agnum mane et alterum vespere
EXOD|29|40|decimam partem similae conspersae oleo tunso quod habeat mensuram quartam partem hin et vinum ad libandum eiusdem mensurae in agno uno
EXOD|29|41|alterum vero agnum offeres ad vesperam iuxta ritum matutinae oblationis et iuxta ea quae diximus in odorem suavitatis
EXOD|29|42|sacrificium Domino oblatione perpetua in generationes vestras ad ostium tabernaculi testimonii coram Domino ubi constituam ut loquar ad te
EXOD|29|43|ibique praecipiam filiis Israhel et sanctificabitur altare in gloria mea
EXOD|29|44|sanctificabo et tabernaculum testimonii cum altari et Aaron cum filiis eius ut sacerdotio fungantur mihi
EXOD|29|45|et habitabo in medio filiorum Israhel eroque eis Deus
EXOD|29|46|et scient quia ego Dominus Deus eorum qui eduxi eos de terra Aegypti ut manerem inter illos ego Dominus Deus ipsorum
EXOD|30|1|facies quoque altare in adolendum thymiama de lignis setthim
EXOD|30|2|habens cubitum longitudinis et alterum latitudinis id est quadrangulum et duos cubitos in altitudine cornua ex ipso procedent
EXOD|30|3|vestiesque illud auro purissimo tam craticulam eius quam parietes per circuitum et cornua faciesque ei coronam aureolam per gyrum
EXOD|30|4|et duos anulos aureos sub corona per singula latera ut mittantur in eos vectes et altare portetur
EXOD|30|5|ipsos quoque vectes facies de lignis setthim et inaurabis
EXOD|30|6|ponesque altare contra velum quod ante arcam pendet testimonii coram propitiatorio quo tegitur testimonium ubi loquar tibi
EXOD|30|7|et adolebit incensum super eo Aaron suave fraglans mane quando conponet lucernas incendet illud
EXOD|30|8|et quando conlocat eas ad vesperum uret thymiama sempiternum coram Domino in generationes vestras
EXOD|30|9|non offeretis super eo thymiama conpositionis alterius nec oblationem et victimam nec liba libabitis
EXOD|30|10|et deprecabitur Aaron super cornua eius semel per annum in sanguine quod oblatum est pro peccato et placabit super eo in generationibus vestris sanctum sanctorum erit Domino
EXOD|30|11|locutusque est Dominus ad Mosen dicens
EXOD|30|12|quando tuleris summam filiorum Israhel iuxta numerum dabunt singuli pretium pro animabus suis Domino et non erit plaga in eis cum fuerint recensiti
EXOD|30|13|hoc autem dabit omnis qui transit ad nomen dimidium sicli iuxta mensuram templi siclus viginti obolos habet media pars sicli offeretur Domino
EXOD|30|14|qui habetur in numero a viginti annis et supra dabit pretium
EXOD|30|15|dives non addet ad medium sicli et pauper nihil minuet
EXOD|30|16|susceptamque pecuniam quae conlata est a filiis Israhel trades in usus tabernaculi testimonii ut sit monumentum eorum coram Domino et propitietur animabus illorum
EXOD|30|17|locutusque est Dominus ad Mosen dicens
EXOD|30|18|facies et labium aeneum cum basi sua ad lavandum ponesque illud inter tabernaculum testimonii et altare et missa aqua
EXOD|30|19|lavabunt in eo Aaron et filii eius manus suas ac pedes
EXOD|30|20|quando ingressuri sunt tabernaculum testimonii et quando accessuri ad altare ut offerant in eo thymiama Domino
EXOD|30|21|ne forte moriantur legitimum sempiternum erit ipsi et semini eius per successiones
EXOD|30|22|locutusque est Dominus ad Mosen
EXOD|30|23|dicens sume tibi aromata prima et zmyrnae electae quingentos siclos et cinnamomi medium id est ducentos quinquaginta calami similiter ducentos quinquaginta
EXOD|30|24|cassiae autem quingentos siclos in pondere sanctuarii olei de olivetis mensuram hin
EXOD|30|25|faciesque unctionis oleum sanctum unguentum conpositum opere unguentarii
EXOD|30|26|et ungues ex eo tabernaculum testimonii et arcam testamenti
EXOD|30|27|mensamque cum vasis suis candelabrum et utensilia eius altaria thymiamatis
EXOD|30|28|et holocausti et universam supellectilem quae ad cultum eorum pertinent
EXOD|30|29|sanctificabisque omnia et erunt sancta sanctorum qui tetigerit ea sanctificabitur
EXOD|30|30|Aaron et filios eius ungues sanctificabisque eos ut sacerdotio fungantur mihi
EXOD|30|31|filiis quoque Israhel dices hoc oleum unctionis sanctum erit mihi in generationes vestras
EXOD|30|32|caro hominis non unguetur ex eo et iuxta conpositionem eius non facietis aliud quia sanctificatum est et sanctum erit vobis
EXOD|30|33|homo quicumque tale conposuerit et dederit ex eo alieno exterminabitur de populo suo
EXOD|30|34|dixitque Dominus ad Mosen sume tibi aromata stacten et onycha galbanen boni odoris et tus lucidissimum aequalis ponderis erunt omnia
EXOD|30|35|faciesque thymiama conpositum opere unguentarii mixtum diligenter et purum et sanctificatione dignissimum
EXOD|30|36|cumque in tenuissimum pulverem universa contuderis pones ex eo coram testimonio tabernaculi in quo loco apparebo tibi sanctum sanctorum erit vobis thymiama
EXOD|30|37|talem conpositionem non facietis in usus vestros quia sanctum est Domino
EXOD|30|38|homo quicumque fecerit simile ut odore illius perfruatur peribit de populis suis
EXOD|31|1|locutusque est Dominus ad Mosen dicens
EXOD|31|2|ecce vocavi ex nomine Beselehel filium Uri filii Hur de tribu Iuda
EXOD|31|3|et implevi eum spiritu Dei sapientia intellegentia et scientia in omni opere
EXOD|31|4|ad excogitandum fabre quicquid fieri potest ex auro et argento et aere
EXOD|31|5|marmore et gemmis et diversitate lignorum
EXOD|31|6|dedique ei socium Hooliab filium Achisamech de tribu Dan et in corde omnis eruditi posui sapientiam ut faciant cuncta quae praecepi tibi
EXOD|31|7|tabernaculum foederis et arcam testimonii et propitiatorium quod super eam est et cuncta vasa tabernaculi
EXOD|31|8|mensamque et vasa eius candelabrum purissimum cum vasis suis et altaria thymiamatis
EXOD|31|9|et holocausti et omnia vasa eorum labium cum basi sua
EXOD|31|10|vestes sanctas in ministerio Aaron sacerdoti et filiis eius ut fungantur officio suo in sacris
EXOD|31|11|oleum unctionis et thymiama aromatum in sanctuario omnia quae praecepi tibi facient
EXOD|31|12|et locutus est Dominus ad Mosen dicens
EXOD|31|13|loquere filiis Israhel et dices ad eos videte ut sabbatum meum custodiatis quia signum est inter me et vos in generationibus vestris ut sciatis quia ego Dominus qui sanctifico vos
EXOD|31|14|custodite sabbatum sanctum est enim vobis qui polluerit illud morte morietur qui fecerit in eo opus peribit anima illius de medio populi sui
EXOD|31|15|sex diebus facietis opus in die septimo sabbatum est requies sancta Domino omnis qui fecerit opus in hac die morietur
EXOD|31|16|custodiant filii Israhel sabbatum et celebrent illud in generationibus suis pactum est sempiternum
EXOD|31|17|inter me et filios Israhel signumque perpetuum sex enim diebus fecit Dominus caelum et terram et in septimo ab opere cessavit
EXOD|31|18|dedit quoque Mosi conpletis huiuscemodi sermonibus in monte Sinai duas tabulas testimonii lapideas scriptas digito Dei
EXOD|32|1|videns autem populus quod moram faceret descendendi de monte Moses congregatus adversus Aaron ait surge fac nobis deos qui nos praecedant Mosi enim huic viro qui nos eduxit de terra Aegypti ignoramus quid acciderit
EXOD|32|2|dixitque ad eos Aaron tollite inaures aureas de uxorum filiorumque et filiarum vestrarum auribus et adferte ad me
EXOD|32|3|fecit populus quae iusserat deferens inaures ad Aaron
EXOD|32|4|quas cum ille accepisset formavit opere fusorio et fecit ex eis vitulum conflatilem dixeruntque hii sunt dii tui Israhel qui te eduxerunt de terra Aegypti
EXOD|32|5|quod cum vidisset Aaron aedificavit altare coram eo et praeconis voce clamavit dicens cras sollemnitas Domini est
EXOD|32|6|surgentesque mane obtulerunt holocausta et hostias pacificas et sedit populus comedere ac bibere et surrexerunt ludere
EXOD|32|7|locutus est autem Dominus ad Mosen vade descende peccavit populus tuus quem eduxisti de terra Aegypti
EXOD|32|8|recesserunt cito de via quam ostendisti eis feceruntque sibi vitulum conflatilem et adoraverunt atque immolantes ei hostias dixerunt isti sunt dii tui Israhel qui te eduxerunt de terra Aegypti
EXOD|32|9|rursumque ait Dominus ad Mosen cerno quod populus iste durae cervicis sit
EXOD|32|10|dimitte me ut irascatur furor meus contra eos et deleam eos faciamque te in gentem magnam
EXOD|32|11|Moses autem orabat Dominum Deum suum dicens cur Domine irascitur furor tuus contra populum tuum quem eduxisti de terra Aegypti in fortitudine magna et in manu robusta
EXOD|32|12|ne quaeso dicant Aegyptii callide eduxit eos ut interficeret in montibus et deleret e terra quiescat ira tua et esto placabilis super nequitia populi tui
EXOD|32|13|recordare Abraham Isaac et Israhel servorum tuorum quibus iurasti per temet ipsum dicens multiplicabo semen vestrum sicut stellas caeli et universam terram hanc de qua locutus sum dabo semini vestro et possidebitis eam semper
EXOD|32|14|placatusque est Dominus ne faceret malum quod locutus fuerat adversus populum suum
EXOD|32|15|et reversus est Moses de monte portans duas tabulas testimonii manu scriptas ex utraque parte
EXOD|32|16|et factas opere Dei scriptura quoque Dei erat sculpta in tabulis
EXOD|32|17|audiens autem Iosue tumultum populi vociferantis dixit ad Mosen ululatus pugnae auditur in castris
EXOD|32|18|qui respondit non est clamor adhortantium ad pugnam neque vociferatio conpellentium ad fugam sed vocem cantantium ego audio
EXOD|32|19|cumque adpropinquasset ad castra vidit vitulum et choros iratusque valde proiecit de manu tabulas et confregit eas ad radices montis
EXOD|32|20|arripiensque vitulum quem fecerant conbusit et contrivit usque ad pulverem quem sparsit in aqua et dedit ex eo potum filiis Israhel
EXOD|32|21|dixitque ad Aaron quid tibi fecit hic populus ut induceres super eum peccatum maximum
EXOD|32|22|cui ille respondit ne indignetur dominus meus tu enim nosti populum istum quod pronus sit ad malum
EXOD|32|23|dixerunt mihi fac nobis deos qui praecedant nos huic enim Mosi qui nos eduxit de terra Aegypti nescimus quid acciderit
EXOD|32|24|quibus ego dixi quis vestrum habet aurum tulerunt et dederunt mihi et proieci illud in ignem egressusque est hic vitulus
EXOD|32|25|videns ergo Moses populum quod esset nudatus spoliaverat enim eum Aaron propter ignominiam sordis et inter hostes nudum constituerat
EXOD|32|26|et stans in porta castrorum ait si quis est Domini iungatur mihi congregatique sunt ad eum omnes filii Levi
EXOD|32|27|quibus ait haec dicit Dominus Deus Israhel ponat vir gladium super femur suum ite et redite de porta usque ad portam per medium castrorum et occidat unusquisque fratrem et amicum et proximum suum
EXOD|32|28|fecerunt filii Levi iuxta sermonem Mosi cecideruntque in die illo quasi tria milia hominum
EXOD|32|29|et ait Moses consecrastis manus vestras hodie Domino unusquisque in filio et fratre suo ut detur vobis benedictio
EXOD|32|30|facto autem die altero locutus est Moses ad populum peccastis peccatum maximum ascendam ad Dominum si quo modo eum quivero deprecari pro scelere vestro
EXOD|32|31|reversusque ad Dominum ait obsecro peccavit populus iste peccatum magnum feceruntque sibi deos aureos aut dimitte eis hanc noxam
EXOD|32|32|aut si non facis dele me de libro tuo quem scripsisti
EXOD|32|33|cui respondit Dominus qui peccaverit mihi delebo eum de libro meo
EXOD|32|34|tu autem vade et duc populum istum quo locutus sum tibi angelus meus praecedet te ego autem in die ultionis visitabo et hoc peccatum eorum
EXOD|32|35|percussit ergo Dominus populum pro reatu vituli quem fecit Aaron
EXOD|33|1|locutusque est Dominus ad Mosen vade ascende de loco isto tu et populus tuus quem eduxisti de terra Aegypti in terram quam iuravi Abraham Isaac et Iacob dicens semini tuo dabo eam
EXOD|33|2|et mittam praecursorem tui angelum ut eiciam Chananeum et Amorreum et Hettheum et Ferezeum et Eveum et Iebuseum
EXOD|33|3|et intres in terram fluentem lacte et melle non enim ascendam tecum quia populus durae cervicis est ne forte disperdam te in via
EXOD|33|4|audiens populus sermonem hunc pessimum luxit et nullus ex more indutus est cultu suo
EXOD|33|5|dixitque Dominus ad Mosen loquere filiis Israhel populus durae cervicis es semel ascendam in medio tui et delebo te iam nunc depone ornatum tuum ut sciam quid faciam tibi
EXOD|33|6|deposuerunt ergo filii Israhel ornatum suum a monte Horeb
EXOD|33|7|Moses quoque tollens tabernaculum tetendit extra castra procul vocavitque nomen eius tabernaculum foederis et omnis populus qui habebat aliquam quaestionem egrediebatur ad tabernaculum foederis extra castra
EXOD|33|8|cumque egrederetur Moses ad tabernaculum surgebat universa plebs et stabat unusquisque in ostio papilionis sui aspiciebantque tergum Mosi donec ingrederetur tentorium
EXOD|33|9|ingresso autem illo tabernaculum foederis descendebat columna nubis et stabat ad ostium loquebaturque cum Mosi
EXOD|33|10|cernentibus universis quod columna nubis staret ad ostium tabernaculi stabantque ipsi et adorabant per fores tabernaculorum suorum
EXOD|33|11|loquebatur autem Dominus ad Mosen facie ad faciem sicut loqui solet homo ad amicum suum cumque ille reverteretur in castra minister eius Iosue filius Nun puer non recedebat de tabernaculo
EXOD|33|12|dixit autem Moses ad Dominum praecipis ut educam populum istum et non indicas mihi quem missurus es mecum praesertim cum dixeris novi te ex nomine et invenisti gratiam coram me
EXOD|33|13|si ergo inveni gratiam in conspectu tuo ostende mihi viam tuam ut sciam te et inveniam gratiam ante oculos tuos respice populum tuum gentem hanc
EXOD|33|14|dixitque Dominus facies mea praecedet te et requiem dabo tibi
EXOD|33|15|et ait Moses si non tu ipse praecedes ne educas nos de loco isto
EXOD|33|16|in quo enim scire poterimus ego et populus tuus invenisse nos gratiam in conspectu tuo nisi ambulaveris nobiscum ut glorificemur ab omnibus populis qui habitant super terram
EXOD|33|17|dixit autem Dominus ad Mosen et verbum istud quod locutus es faciam invenisti enim gratiam coram me et te ipsum novi ex nomine
EXOD|33|18|qui ait ostende mihi gloriam tuam
EXOD|33|19|respondit ego ostendam omne bonum tibi et vocabo in nomine Domini coram te et miserebor cui voluero et clemens ero in quem mihi placuerit
EXOD|33|20|rursumque ait non poteris videre faciem meam non enim videbit me homo et vivet
EXOD|33|21|et iterum ecce inquit est locus apud me stabis super petram
EXOD|33|22|cumque transibit gloria mea ponam te in foramine petrae et protegam dextera mea donec transeam
EXOD|33|23|tollamque manum meam et videbis posteriora mea faciem autem meam videre non poteris
EXOD|34|1|ac deinceps praecide ait tibi duas tabulas lapideas instar priorum et scribam super eas verba quae habuerunt tabulae quas fregisti
EXOD|34|2|esto paratus mane ut ascendas statim in montem Sinai stabisque mecum super verticem montis
EXOD|34|3|nullus ascendat tecum nec videatur quispiam per totum montem boves quoque et oves non pascantur e contra
EXOD|34|4|excidit ergo duas tabulas lapideas quales ante fuerant et de nocte consurgens ascendit in montem Sinai sicut ei praeceperat Dominus portans secum tabulas
EXOD|34|5|cumque descendisset Dominus per nubem stetit Moses cum eo invocans nomen Domini
EXOD|34|6|quo transeunte coram eo ait Dominator Domine Deus misericors et clemens patiens et multae miserationis ac verus
EXOD|34|7|qui custodis misericordiam in milia qui aufers iniquitatem et scelera atque peccata nullusque apud te per se innocens est qui reddis iniquitatem patrum in filiis ac nepotibus in tertiam et quartam progeniem
EXOD|34|8|festinusque Moses curvatus est pronus in terram et adorans
EXOD|34|9|ait si inveni gratiam in conspectu tuo Domine obsecro ut gradiaris nobiscum populus enim durae cervicis est et auferas iniquitates nostras atque peccata nosque possideas
EXOD|34|10|respondit Dominus ego inibo pactum videntibus cunctis signa faciam quae numquam sunt visa super terram nec in ullis gentibus ut cernat populus in cuius es medio opus Domini terribile quod facturus sum
EXOD|34|11|observa cuncta quae hodie mando tibi ego ipse eiciam ante faciem tuam Amorreum et Chananeum et Hettheum Ferezeum quoque et Eveum et Iebuseum
EXOD|34|12|cave ne umquam cum habitatoribus terrae illius iungas amicitias quae tibi sint in ruinam
EXOD|34|13|sed aras eorum destrue confringe statuas lucosque succide
EXOD|34|14|noli adorare deum alienum Dominus Zelotes nomen eius Deus est aemulator
EXOD|34|15|ne ineas pactum cum hominibus illarum regionum ne cum fornicati fuerint cum diis suis et adoraverint simulacra eorum vocet te quispiam ut comedas de immolatis
EXOD|34|16|nec uxorem de filiabus eorum accipies filiis tuis ne postquam ipsae fuerint fornicatae fornicari faciant et filios tuos in deos suos
EXOD|34|17|deos conflatiles non facies tibi
EXOD|34|18|sollemnitatem azymorum custodies septem diebus vesceris azymis sicut praecepi tibi in tempore mensis novorum mense enim verni temporis egressus es de Aegypto
EXOD|34|19|omne quod aperit vulvam generis masculini meum erit de cunctis animantibus tam de bubus quam de ovibus meum erit
EXOD|34|20|primogenitum asini redimes ove sin autem nec pretium pro eo dederis occidetur primogenitum filiorum tuorum redimes nec apparebis in conspectu meo vacuus
EXOD|34|21|sex diebus operaberis die septimo cessabis arare et metere
EXOD|34|22|sollemnitatem ebdomadarum facies tibi in primitiis frugum messis tuae triticeae et sollemnitatem quando redeunte anni tempore cuncta conduntur
EXOD|34|23|tribus temporibus anni apparebit omne masculinum tuum in conspectu omnipotentis Domini Dei Israhel
EXOD|34|24|cum enim tulero gentes a facie tua et dilatavero terminos tuos nullus insidiabitur terrae tuae ascendente te et apparente in conspectu Domini Dei tui ter in anno
EXOD|34|25|non immolabis super fermento sanguinem hostiae meae neque residebit mane de victima sollemnitatis phase
EXOD|34|26|primitias frugum terrae tuae offeres in domum Domini Dei tui non coques hedum in lacte matris suae
EXOD|34|27|dixitque Dominus ad Mosen scribe tibi verba haec quibus et tecum et cum Israhel pepigi foedus
EXOD|34|28|fecit ergo ibi cum Domino quadraginta dies et quadraginta noctes panem non comedit et aquam non bibit et scripsit in tabulis verba foederis decem
EXOD|34|29|cumque descenderet Moses de monte Sinai tenebat duas tabulas testimonii et ignorabat quod cornuta esset facies sua ex consortio sermonis Dei
EXOD|34|30|videntes autem Aaron et filii Israhel cornutam Mosi faciem timuerunt prope accedere
EXOD|34|31|vocatique ab eo reversi sunt tam Aaron quam principes synagogae et postquam locutus est
EXOD|34|32|venerunt ad eum etiam omnes filii Israhel quibus praecepit cuncta quae audierat a Domino in monte Sinai
EXOD|34|33|impletisque sermonibus posuit velamen super faciem suam
EXOD|34|34|quod ingressus ad Dominum et loquens cum eo auferebat donec exiret et tunc loquebatur ad filios Israhel omnia quae sibi fuerant imperata
EXOD|34|35|qui videbant faciem egredientis Mosi esse cornutam sed operiebat rursus ille faciem suam si quando loquebatur ad eos
EXOD|35|1|igitur congregata omni turba filiorum Israhel dixit ad eos haec sunt quae iussit Dominus fieri
EXOD|35|2|sex diebus facietis opus septimus dies erit vobis sanctus sabbatum et requies Domini qui fecerit opus in eo occidetur
EXOD|35|3|non succendetis ignem in omnibus habitaculis vestris per diem sabbati
EXOD|35|4|et ait Moses ad omnem catervam filiorum Israhel iste est sermo quem praecepit Dominus dicens
EXOD|35|5|separate apud vos primitias Domino omnis voluntarius et proni animi offerat eas Domino aurum et argentum et aes
EXOD|35|6|hyacinthum purpuram coccumque bis tinctum et byssum pilos caprarum
EXOD|35|7|et pelles arietum rubricatas et ianthinas
EXOD|35|8|ligna setthim
EXOD|35|9|et oleum ad luminaria concinnanda et ut conficiatur unguentum et thymiama suavissimum
EXOD|35|10|lapides onychinos et gemmas ad ornatum superumeralis et rationalis
EXOD|35|11|quisquis vestrum est sapiens veniat et faciat quod Dominus imperavit
EXOD|35|12|tabernaculum scilicet et tectum eius atque operimentum anulos et tabulata cum vectibus paxillos et bases
EXOD|35|13|arcam et vectes propitiatorium et velum quod ante illud oppanditur
EXOD|35|14|mensam cum vectibus et vasis et propositionis panibus
EXOD|35|15|candelabrum ad luminaria sustentanda vasa illius et lucernas et oleum ad nutrimenta ignium
EXOD|35|16|altare thymiamatis et vectes oleum unctionis et thymiama ex aromatibus tentorium ad ostium tabernaculi
EXOD|35|17|altare holocausti et craticulam eius aeneam cum vectibus et vasis suis labrum et basim eius
EXOD|35|18|cortinas atrii cum columnis et basibus tentorium in foribus vestibuli
EXOD|35|19|paxillos tabernaculi et atrii cum funiculis suis
EXOD|35|20|vestimenta quorum usus est in ministerio sanctuarii vestes Aaron pontificis ac filiorum eius ut sacerdotio fungantur mihi
EXOD|35|21|egressaque omnis multitudo filiorum Israhel de conspectu Mosi
EXOD|35|22|obtulit mente promptissima atque devota primitias Domino ad faciendum opus tabernaculi testimonii quicquid in cultum et ad vestes sanctas necessarium erat
EXOD|35|23|viri cum mulieribus praebuerunt armillas et inaures anulos et dextralia omne vas aureum in donaria Domini separatum est
EXOD|35|24|si quis habuit hyacinthum purpuram coccumque bis tinctum byssum et pilos caprarum pelles arietum rubricatas et ianthinas
EXOD|35|25|argenti et aeris metalla obtulerunt Domino lignaque setthim in varios usus
EXOD|35|26|sed et mulieres doctae dederunt quae neverant hyacinthum purpuram et vermiculum ac byssum
EXOD|35|27|et pilos caprarum sponte propria cuncta tribuentes
EXOD|35|28|principes vero obtulerunt lapides onychinos et gemmas ad superumerale et rationale
EXOD|35|29|aromataque et oleum ad luminaria concinnanda et ad praeparandum unguentum ac thymiama odoris suavissimi conponendum
EXOD|35|30|omnes viri et mulieres mente devota obtulerunt donaria ut fierent opera quae iusserat Dominus per manum Mosi cuncti filii Israhel voluntaria Domino dedicaverunt
EXOD|35|31|dixitque Moses ad filios Israhel ecce vocavit Dominus ex nomine Beselehel filium Uri filii Hur de tribu Iuda
EXOD|35|32|implevitque eum spiritu Dei sapientiae et intellegentiae et scientiae omni doctrina
EXOD|35|33|ad excogitandum et faciendum opus in auro et argento et aere sculpendisque lapidibus et opere carpentario quicquid fabre adinveniri potest
EXOD|35|34|dedit in corde eius Hooliab quoque filium Achisamech de tribu Dan
EXOD|35|35|ambos erudivit sapientia ut faciant opera abietarii polymitarii ac plumarii de hyacintho et purpura coccoque bis tincto et bysso et texant omnia ac nova quaeque repperiant
EXOD|36|1|fecit ergo Beselehel et Hooliab et omnis vir sapiens quibus dedit Dominus sapientiam et intellectum ut scirent fabre operari quae in usus sanctuarii necessaria sunt et quae praecepit Dominus
EXOD|36|2|cumque vocasset eos Moses et omnem eruditum virum cui dederat Deus sapientiam et qui sponte sua obtulerant se ad faciendum opus
EXOD|36|3|tradidit eis universa donaria filiorum Israhel qui cum instarent operi cotidie mane vota populus offerebat
EXOD|36|4|unde artifices venire conpulsi
EXOD|36|5|dixerunt Mosi plus offert populus quam necessarium est
EXOD|36|6|iussit ergo Moses praeconis voce cantari nec vir nec mulier quicquam ultra offerat in opere sanctuarii sicque cessatum est a muneribus offerendis
EXOD|36|7|eo quod oblata sufficerent et superabundarent
EXOD|36|8|feceruntque omnes corde sapientes ad explendum opus tabernaculi cortinas decem de bysso retorta et hyacintho et purpura coccoque bis tincto opere vario et arte polymita
EXOD|36|9|quarum una habebat in longitudine viginti octo cubitos et in latitudine quattuor una mensura erat omnium cortinarum
EXOD|36|10|coniunxitque cortinas quinque alteram alteri et alias quinque sibi invicem copulavit
EXOD|36|11|fecit et ansas hyacinthinas in ora cortinae unius ex utroque latere et in ora cortinae alterius similiter
EXOD|36|12|ut contra se invicem venirent ansae et mutuo iungerentur
EXOD|36|13|unde et quinquaginta fudit circulos aureos qui morderent cortinarum ansas et fieret unum tabernaculum
EXOD|36|14|fecit et saga undecim de pilis caprarum ad operiendum tectum tabernaculi
EXOD|36|15|unum sagum habebat in longitudine cubitos triginta et in latitudine cubitos quattuor unius mensurae erant omnia saga
EXOD|36|16|quorum quinque iunxit seorsum et sex alia separatim
EXOD|36|17|fecitque ansas quinquaginta in ora sagi unius et quinquaginta in ora sagi alterius ut sibi invicem iungerentur
EXOD|36|18|et fibulas aeneas quinquaginta quibus necteretur tectum et unum pallium ex omnibus sagis fieret
EXOD|36|19|fecit et opertorium tabernaculi de pellibus arietum rubricatis aliudque desuper velamentum de pellibus ianthinis
EXOD|36|20|fecit et tabulas tabernaculi de lignis setthim stantes
EXOD|36|21|decem cubitorum erat longitudo tabulae unius et unum ac semis cubitum latitudo retinebat
EXOD|36|22|binae incastraturae erant per singulas tabulas ut altera alteri iungeretur sic fecit in omnibus tabulis tabernaculi
EXOD|36|23|e quibus viginti ad plagam meridianam erant contra austrum
EXOD|36|24|cum quadraginta basibus argenteis duae bases sub una tabula ponebantur ex utraque angulorum parte ubi incastraturae laterum in angulis terminantur
EXOD|36|25|ad plagam quoque tabernaculi quae respicit ad aquilonem fecit viginti tabulas
EXOD|36|26|cum quadraginta argenteis basibus duas bases per singulas tabulas
EXOD|36|27|contra occidentem vero id est ad eam partem tabernaculi quae mare respicit fecit sex tabulas
EXOD|36|28|et duas alias per singulos angulos tabernaculi retro
EXOD|36|29|quae iunctae erant deorsum usque sursum et in unam conpagem pariter ferebantur ita fecit ex utraque parte per angulos
EXOD|36|30|ut octo essent simul tabulae et haberent bases argenteas sedecim binas scilicet bases sub singulis tabulis
EXOD|36|31|fecit et vectes de lignis setthim quinque ad continendas tabulas unius lateris tabernaculi
EXOD|36|32|et quinque alios ad alterius lateris tabulas coaptandas et extra hos quinque alios vectes ad occidentalem plagam tabernaculi contra mare
EXOD|36|33|fecit quoque vectem alium qui per medias tabulas ab angulo usque ad angulum perveniret
EXOD|36|34|ipsa autem tabulata deauravit et circulos eorum fecit aureos per quos vectes induci possint quos et ipsos aureis lamminis operuit
EXOD|36|35|fecit et velum de hyacintho purpura vermiculo ac bysso retorta opere polymitario varium atque distinctum
EXOD|36|36|et quattuor columnas de lignis setthim quas cum capitibus deauravit fusis basibus earum argenteis
EXOD|36|37|fecit et tentorium in introitu tabernaculi ex hyacintho purpura vermiculo byssoque retorta opere plumarii
EXOD|36|38|et columnas quinque cum capitibus suis quas operuit auro basesque earum fudit aeneas
EXOD|37|1|fecit autem Beselehel et arcam de lignis setthim habentem duos semis cubitos in longitudinem et cubitum ac semissem in latitudinem altitudo quoque uno cubito fuit et dimidio vestivitque eam auro purissimo intus ac foris
EXOD|37|2|et fecit illi coronam auream per gyrum
EXOD|37|3|conflans quattuor anulos aureos per quattuor angulos eius duos anulos in latere uno et duos in altero
EXOD|37|4|vectes quoque fecit de lignis setthim quos vestivit auro
EXOD|37|5|et quos misit in anulos qui erant in lateribus arcae ad portandum eam
EXOD|37|6|fecit et propitiatorium id est oraculum de auro mundissimo duorum cubitorum et dimidio in longitudine et cubito ac semisse in latitudine
EXOD|37|7|duos etiam cherubin ex auro ductili quos posuit ex utraque parte propitiatorii
EXOD|37|8|cherub unum in summitate huius partis et cherub alterum in summitate partis alterius duos cherubin in singulis summitatibus propitiatorii
EXOD|37|9|extendentes alas et tegentes propitiatorium seque mutuo et illud respectantes
EXOD|37|10|fecit et mensam de lignis setthim in longitudine duorum cubitorum et in latitudine unius cubiti quae habebat in altitudine cubitum ac semissem
EXOD|37|11|circumdeditque eam auro mundissimo et fecit illi labium aureum per gyrum
EXOD|37|12|ipsique labio coronam interrasilem quattuor digitorum et super eandem alteram coronam auream
EXOD|37|13|fudit et quattuor circulos aureos quos posuit in quattuor angulis per singulos pedes mensae
EXOD|37|14|contra coronam misitque in eos vectes ut possit mensa portari
EXOD|37|15|ipsos quoque vectes fecit de lignis setthim et circumdedit eos auro
EXOD|37|16|et vasa ad diversos usus mensae acetabula fialas cyatos et turibula ex auro puro in quibus offerenda sunt liba
EXOD|37|17|fecit et candelabrum ductile de auro mundissimo de cuius vecte calami scyphi spherulae ac lilia procedebant
EXOD|37|18|sex in utroque latere tres calami ex parte una et tres ex altera
EXOD|37|19|tres scyphi in nucis modum per calamos singulos spherulaeque simul et lilia et tres scyphi instar nucis in calamo altero spherulaeque simul et lilia aequum erat opus sex calamorum qui procedebant de stipite candelabri
EXOD|37|20|in ipso autem vecte erant quattuor scyphi in nucis modum spherulaeque per singulos et lilia
EXOD|37|21|et spherae sub duobus calamis per loca tria qui simul sex fiunt calami procedentes de vecte uno
EXOD|37|22|et spherae igitur et calami ex ipso erant universa ductilia de auro purissimo
EXOD|37|23|fecit et lucernas septem cum emunctoriis suis et vasa ubi quae emuncta sunt extinguuntur de auro mundissimo
EXOD|37|24|talentum auri adpendebat candelabrum cum omnibus vasis suis
EXOD|37|25|fecit et altare thymiamatis de lignis setthim habens per quadrum singulos cubitos et in altitudine duos e cuius angulis procedebant cornua
EXOD|37|26|vestivitque illud auro purissimo cum craticula ac parietibus et cornibus
EXOD|37|27|fecitque ei coronam aureolam per gyrum et duos anulos aureos sub corona per singula latera ut mittantur in eos vectes et possit altare portari
EXOD|37|28|ipsos autem vectes fecit de lignis setthim et operuit lamminis aureis
EXOD|37|29|conposuit et oleum ad sanctificationis unguentum et thymiama de aromatibus mundissimis opere pigmentarii
EXOD|38|1|fecit et altare holocausti de lignis setthim quinque cubitorum per quadrum et trium in altitudine
EXOD|38|2|cuius cornua de angulis procedebant operuitque illud aeneis lamminis
EXOD|38|3|et in usus eius paravit ex aere vasa diversa lebetas forcipes fuscinulas uncinos et ignium receptacula
EXOD|38|4|craticulamque eius in modum retis fecit aeneam et subter eam in altaris medio arulam
EXOD|38|5|fusis quattuor anulis per totidem retiaculi summitates ad inmittendos vectes ad portandum
EXOD|38|6|quos et ipsos fecit de lignis setthim et operuit lamminis aeneis
EXOD|38|7|induxitque in circulos qui in altaris lateribus eminebant ipsum autem altare non erat solidum sed cavum ex tabulis et intus vacuum
EXOD|38|8|fecit et labrum aeneum cum base sua de speculis mulierum quae excubabant in ostio tabernaculi
EXOD|38|9|et atrium in cuius australi plaga erant tentoria de bysso retorta cubitorum centum
EXOD|38|10|columnae aeneae viginti cum basibus suis capita columnarum et tota operis celatura argentea
EXOD|38|11|aeque ad septentrionalis plagam tentoria columnae basesque et capita columnarum eiusdem et mensurae et operis ac metalli erant
EXOD|38|12|in ea vero plaga quae occidentem respicit fuere tentoria cubitorum quinquaginta columnae decem cum basibus suis aeneae et capita columnarum celata argentea
EXOD|38|13|porro contra orientem quinquaginta cubitorum paravit tentoria
EXOD|38|14|e quibus quindecim cubitos columnarum trium cum basibus suis unum tenebat latus
EXOD|38|15|et in parte altera quia utraque introitum tabernaculi facit quindecim aeque cubitorum erant tentoria columnae tres et bases totidem
EXOD|38|16|cuncta atrii tentoria byssus torta texuerat
EXOD|38|17|bases columnarum fuere aeneae capita autem earum cum celaturis suis argentea sed et ipsas columnas atrii vestivit argento
EXOD|38|18|et in introitu eius opere plumario fecit tentorium ex hyacintho purpura vermiculo ac bysso retorta quod habebat viginti cubitos in longitudine altitudo vero quinque cubitorum erat iuxta mensuram quam cuncta atrii habebant tentoria
EXOD|38|19|columnae autem ingressus fuere quattuor cum basibus aeneis capitaque earum et celaturae argenteae
EXOD|38|20|paxillos quoque tabernaculi et atrii per gyrum fecit aeneos
EXOD|38|21|haec sunt instrumenta tabernaculi testimonii quae numerata sunt iuxta praeceptum Mosi in caerimonias Levitarum per manum Ithamar filii Aaron sacerdotis
EXOD|38|22|quas Beselehel filius Uri filii Hur de tribu Iuda Domino per Mosen iubente conpleverat
EXOD|38|23|iuncto sibi socio Hooliab filio Achisamech de tribu Dan qui et ipse artifex lignorum egregius fuit et polymitarius atque plumarius ex hyacintho purpura vermiculo et bysso
EXOD|38|24|omne aurum quod expensum est in opere sanctuarii et quod oblatum in donariis viginti novem talentorum fuit et septingentorum triginta siclorum ad mensuram sanctuarii
EXOD|38|25|oblatum est autem ab his qui transierant ad numerum a viginti annis et supra de sescentis tribus milibus et quingentis quinquaginta armatorum
EXOD|38|26|fuerunt praeterea centum talenta argenti e quibus conflatae sunt bases sanctuarii et introitus ubi velum pendet
EXOD|38|27|centum bases factae sunt de talentis centum singulis talentis per bases singulas supputatis
EXOD|38|28|de mille autem septingentis et septuaginta quinque fecit capita columnarum quas et ipsas vestivit argento
EXOD|38|29|aeris quoque oblata sunt talenta septuaginta duo milia et quadringenti supra sicli
EXOD|38|30|ex quibus fusae sunt bases in introitu tabernaculi testimonii et altare aeneum cum craticula sua omniaque vasa quae ad usum eius pertinent
EXOD|38|31|et bases atrii tam in circuitu quam in ingressu eius et paxilli tabernaculi atque atrii per gyrum
EXOD|39|1|de hyacintho vero et purpura vermiculo ac bysso fecit vestes quibus indueretur Aaron quando ministrabat in sanctis sicut praecepit Dominus Mosi
EXOD|39|2|fecit igitur superumerale de auro hyacintho et purpura coccoque bis tincto et bysso retorta
EXOD|39|3|opere polymitario inciditque bratteas aureas et extenuavit in fila ut possint torqueri cum priorum colorum subtemine
EXOD|39|4|duasque oras sibi invicem copulatas in utroque latere summitatum
EXOD|39|5|et balteum ex hisdem coloribus sicut praeceperat Dominus Mosi
EXOD|39|6|paravit et duos lapides onychinos adstrictos et inclusos auro et sculptos arte gemmaria nominibus filiorum Israhel
EXOD|39|7|posuitque eos in lateribus superumeralis in monumentum filiorum Israhel sicut praeceperat Dominus Mosi
EXOD|39|8|fecit et rationale opere polymito iuxta opus superumeralis ex auro hyacintho purpura coccoque bis tincto et bysso retorta
EXOD|39|9|quadrangulum duplex mensurae palmi
EXOD|39|10|et posuit in eo gemmarum ordines quattuor in primo versu erat sardius topazius zmaragdus
EXOD|39|11|in secundo carbunculus sapphyrus iaspis
EXOD|39|12|in tertio ligyrius achates amethistus
EXOD|39|13|in quarto chrysolitus onychinus berillus circumdati et inclusi auro per ordines suos
EXOD|39|14|ipsique lapides duodecim sculpti erant nominibus duodecim tribuum Israhel singuli per nomina singulorum
EXOD|39|15|fecerunt in rationali et catenulas sibi invicem coherentes de auro purissimo
EXOD|39|16|et duos uncinos totidemque anulos aureos porro anulos posuerunt in utroque latere rationalis
EXOD|39|17|e quibus penderent duae catenae aureae quas inseruerunt uncinis qui in superumeralis angulis eminebant
EXOD|39|18|haec et ante et retro ita conveniebant sibi ut superumerale et rationale mutuo necterentur
EXOD|39|19|stricta ad balteum et anulis fortius copulata quos iungebat vitta hyacinthina ne laxe fluerent et a se invicem moverentur sicut praecepit Dominus Mosi
EXOD|39|20|fecerunt quoque tunicam superumeralis totam hyacinthinam
EXOD|39|21|et capitium in superiori parte contra medium oramque per gyrum capitii textilem
EXOD|39|22|deorsum autem ad pedes mala punica ex hyacintho purpura vermiculo ac bysso retorta
EXOD|39|23|et tintinabula de auro mundissimo quae posuerunt inter mala granata in extrema parte tunicae per gyrum
EXOD|39|24|tintinabulum aureum et malum punicum quibus ornatus incedebat pontifex quando ministerio fungebatur sicut praecepit Dominus Mosi
EXOD|39|25|fecerunt et tunicas byssinas opere textili Aaron et filiis eius
EXOD|39|26|et mitras cum coronulis suis ex bysso
EXOD|39|27|feminalia quoque linea byssina
EXOD|39|28|cingulum vero de bysso retorta hyacintho purpura ac vermiculo distinctum arte plumaria sicut praecepit Dominus Mosi
EXOD|39|29|fecerunt et lamminam sacrae venerationis de auro purissimo scripseruntque in ea opere gemmario Sanctum Domini
EXOD|39|30|et strinxerunt eam cum mitra vitta hyacinthina sicut praecepit Dominus Mosi
EXOD|39|31|perfectum est igitur omne opus tabernaculi et tecti testimonii feceruntque filii Israhel cuncta quae praeceperat Dominus Mosi
EXOD|39|32|et obtulerunt tabernaculum et tectum et universam supellectilem anulos tabulas vectes columnas ac bases
EXOD|39|33|opertorium de pellibus arietum rubricatis et aliud operimentum de ianthinis pellibus
EXOD|39|34|velum arcam vectes propitiatorium
EXOD|39|35|mensam cum vasis et propositionis panibus
EXOD|39|36|candelabrum lucernas et utensilia eorum cum oleo
EXOD|39|37|altare aureum et unguentum thymiama ex aromatibus
EXOD|39|38|et tentorium in introitu tabernaculi
EXOD|39|39|altare aeneum retiaculum vectes et vasa eius omnia labrum cum basi sua tentoria atrii et columnas cum basibus suis
EXOD|39|40|tentorium in introitu atrii funiculosque illius et paxillos nihil ex vasis defuit quae in ministerium tabernaculi et in tectum foederis iussa sunt fieri
EXOD|39|41|vestes quoque quibus sacerdotes utuntur in sanctuario Aaron scilicet et filii eius
EXOD|39|42|obtulerunt filii Israhel sicut praeceperat Dominus
EXOD|39|43|quae postquam Moses cuncta vidit expleta benedixit eis
EXOD|40|1|locutusque est Dominus ad Mosen dicens
EXOD|40|2|mense primo die prima mensis eriges tabernaculum testimonii
EXOD|40|3|et pones in eo arcam dimittesque ante illam velum
EXOD|40|4|et inlata mensa pones super eam quae rite praecepta sunt candelabrum stabit cum lucernis suis
EXOD|40|5|et altare aureum in quo adoletur incensum coram arca testimonii tentorium in introitu tabernaculi pones
EXOD|40|6|et ante illud altare holocausti
EXOD|40|7|labrum inter altare et tabernaculum quod implebis aqua
EXOD|40|8|circumdabisque atrium tentoriis et ingressum eius
EXOD|40|9|et adsumpto unctionis oleo ungues tabernaculum cum vasis suis ut sanctificentur
EXOD|40|10|altare holocausti et omnia vasa eius
EXOD|40|11|labrum cum basi sua omnia unctionis oleo consecrabis ut sint sancta sanctorum
EXOD|40|12|adplicabisque Aaron et filios eius ad fores tabernaculi testimonii et lotos aqua
EXOD|40|13|indues sanctis vestibus ut ministrent mihi et unctio eorum in sacerdotium proficiat sempiternum
EXOD|40|14|fecitque Moses omnia quae praeceperat Dominus
EXOD|40|15|igitur mense primo anni secundi in prima die mensis conlocatum est tabernaculum
EXOD|40|16|erexitque illud Moses et posuit tabulas ac bases et vectes statuitque columnas
EXOD|40|17|et expandit tectum super tabernaculum inposito desuper operimento sicut Dominus imperarat
EXOD|40|18|posuit et testimonium in arca subditis infra vectibus et oraculum desuper
EXOD|40|19|cumque intulisset arcam in tabernaculum adpendit ante eam velum ut expleret Domini iussionem
EXOD|40|20|posuit et mensam in tabernaculo testimonii ad plagam septentrionalem extra velum
EXOD|40|21|ordinatis coram propositionis panibus sicut praeceperat Dominus Mosi
EXOD|40|22|posuit et candelabrum in tabernaculum testimonii e regione mensae in parte australi
EXOD|40|23|locatis per ordinem lucernis iuxta praeceptum Domini
EXOD|40|24|posuit et altare aureum sub tecto testimonii contra velum
EXOD|40|25|et adolevit super eo incensum aromatum sicut iusserat Dominus
EXOD|40|26|posuit et tentorium in introitu tabernaculi
EXOD|40|27|et altare holocausti in vestibulo testimonii offerens in eo holocaustum et sacrificia ut Dominus imperarat
EXOD|40|28|labrum quoque statuit inter tabernaculum testimonii et altare implens illud aqua
EXOD|40|29|laveruntque Moses et Aaron ac filii eius manus suas et pedes
EXOD|40|30|cum ingrederentur tectum foederis et accederent ad altare sicut praeceperat Dominus
EXOD|40|31|erexit et atrium per gyrum tabernaculi et altaris ducto in introitu eius tentorio postquam cuncta perfecta sunt
EXOD|40|32|operuit nubes tabernaculum testimonii et gloria Domini implevit illud
EXOD|40|33|nec poterat Moses ingredi tectum foederis nube operiente omnia et maiestate Domini coruscante quia cuncta nubes operuerat
EXOD|40|34|si quando nubes tabernaculum deserebat proficiscebantur filii Israhel per turmas suas
EXOD|40|35|si pendebat desuper manebant in eodem loco
EXOD|40|36|nubes quippe Domini incubabat per diem tabernaculo et ignis in nocte videntibus populis Israhel per cunctas mansiones suas
