DEUT|1|1|以下是 摩西 在 約旦河 東的曠野， 疏弗 對面的 亞拉巴 ，就是在 巴蘭 、 陀弗 、 拉班 、 哈洗錄 、 底撒哈 之間，向 以色列 眾人所說的話。
DEUT|1|2|從 何烈山 經過 西珥山 到 加低斯‧巴尼亞 要十一天的路程。
DEUT|1|3|第四十年十一月初一， 摩西 照耶和華所吩咐他一切有關 以色列 人的話，都告訴他們。
DEUT|1|4|那時，他已經擊敗了住 希實本 的 亞摩利 王 西宏 和住 亞斯她錄 、 以得來 的 巴珊 王 噩 。
DEUT|1|5|摩西 在 約旦河 東的 摩押 地講解這律法，說：
DEUT|1|6|「耶和華－我們的上帝在 何烈山 吩咐我們說：你們住在這山上已經夠久了。
DEUT|1|7|要起行，轉到 亞摩利 人的山區和附近的地區，就是 亞拉巴 、山區、 謝非拉 、 尼革夫 、沿海一帶， 迦南 人的地和 黎巴嫩 ，直到 大河 ，就是 幼發拉底河 。
DEUT|1|8|看，我將這地擺在你們面前。你們要進去得這地，就是耶和華向你們列祖 亞伯拉罕 、 以撒 、 雅各 起誓要賜給他們和他們後裔為業之地。」
DEUT|1|9|「那時，我對你們說：『我獨自一人無法承擔你們的事。
DEUT|1|10|耶和華－你們的上帝使你們增多。看哪，你們今日好像天上的星那樣多。
DEUT|1|11|惟願耶和華－你們列祖的上帝使你們更增加千倍，照他所應許你們的賜福給你們。
DEUT|1|12|但你們的擔子，你們的重任，以及你們的爭訟，我獨自一人怎能承擔呢？
DEUT|1|13|你們要按著各支派選出有智慧、明辨是非、為人所知的人來，我就立他們為你們的領袖。』
DEUT|1|14|你們回答我說：『你說要做的事很好！』
DEUT|1|15|我就將你們各支派的領袖，就是有智慧、為人所知的人，立他們為領袖，作你們各支派的千夫長、百夫長、五十夫長、十夫長等官長，來管理你們。
DEUT|1|16|「當時，我吩咐你們的審判官說：『你們聽訟，無論是弟兄之間的訴訟，或與寄居者之間的訴訟，都要秉公判斷。
DEUT|1|17|審判的時候不可看人的情面；無論大小，你們都要聽訟。不可因人而懼怕，因為審判是上帝的事。你們當中若有難斷的案件，可以呈到我這裏，讓我來聽訟。』
DEUT|1|18|那時，我已經把你們所當做的事都吩咐你們了。」
DEUT|1|19|「我們照著耶和華－我們上帝所吩咐的，從 何烈山 起行，經過你們所看見那一切大而可怕的曠野，往 亞摩利 人的山區去，到了 加低斯‧巴尼亞 。
DEUT|1|20|我對你們說：『你們已經到了耶和華－我們上帝所賜給我們的 亞摩利 人之山區。
DEUT|1|21|看，耶和華－你的上帝已將那地擺在你面前，你要照耶和華－你列祖的上帝所說的，上去得那地為業。不要懼怕，也不要驚惶。』
DEUT|1|22|你們都來到我這裏，說：『讓我們先派人去，為我們窺探那地，把我們上去該走的路線和該進的城鎮回報我們。』
DEUT|1|23|這話我看為美，就從你們中間選取十二個人，每支派一人。
DEUT|1|24|於是他們起身上山區去，到 以實各谷 ，窺探那地。
DEUT|1|25|他們的手帶著那地的一些果子，下到我們這裏，回報我們說：『耶和華－我們的上帝所賜給我們的是美地。』
DEUT|1|26|「你們卻不肯上去，竟違背了耶和華─你們上帝的指示，
DEUT|1|27|在帳棚內發怨言說：『耶和華因為恨我們，所以將我們從 埃及 地領出來，要把我們交在 亞摩利 人的手中，除滅我們。
DEUT|1|28|我們上哪裏去呢？我們的弟兄使我們膽戰心驚 ，說那裏的百姓比我們又大又高 ，那裏的城鎮又大，城牆又堅固，如天一樣高，並且我們在那裏看見 亞衲 族人。』
DEUT|1|29|我就對你們說：『不要驚惶，也不要怕他們。
DEUT|1|30|在你們前面行的耶和華－你們的上帝必為你們爭戰，正如他在 埃及 ，在你們眼前為你們所做的一樣；
DEUT|1|31|並且你們在曠野所行的一切路上，也看見了耶和華─你們的上帝背著你們，如同人背自己的兒子一樣，直到你們來到這地方。』
DEUT|1|32|你們在這事上卻不信耶和華─你們的上帝。
DEUT|1|33|他一路行在你們前面，為你們尋找安營的地方；他夜間在火中，日間在雲中，指示你們當走的路。」
DEUT|1|34|「耶和華聽見你們的怨言，就發怒，起誓說：
DEUT|1|35|『這邪惡世代的人，一個也不得看見我起誓要賜給你們列祖的美地；
DEUT|1|36|惟有 耶孚尼 的兒子 迦勒 必得看見，並且我要將他所踏過的地賜給他和他的子孫，因為他專心跟從我。』
DEUT|1|37|耶和華也因你們的緣故向我發怒，說：『你也不得進入那地。
DEUT|1|38|那侍候你， 嫩 的兒子 約書亞 必得進入那地。你要勉勵他，因為他要使 以色列 承受那地為業。
DEUT|1|39|你們的孩子，你們說要成為擄物的，就是今日尚不知善惡的兒女，必進入那地。我要將那地賜給他們，他們必得為業。
DEUT|1|40|至於你們，要轉回，從 紅海 的路往曠野去。』
DEUT|1|41|「你們回答我說：『我們得罪了耶和華！現在我們願遵照耶和華─我們上帝一切所吩咐的上去爭戰。』於是你們各人帶著兵器，以為很容易就能上到山區去。
DEUT|1|42|耶和華對我說：『你對他們說：不要上去，也不要爭戰，因我不在你們中間，恐怕你們在仇敵面前被擊敗。』
DEUT|1|43|我就告訴了你們，你們卻不聽從，竟違背耶和華的指示，擅自上到山區去。
DEUT|1|44|住在那山區的 亞摩利 人像蜂群一樣出來迎擊你們，追趕你們，在 西珥 擊敗你們，直到 何珥瑪 。
DEUT|1|45|你們就回來，在耶和華面前哭泣；耶和華卻不聽你們的聲音，也不向你們側耳。
DEUT|1|46|你們照著所停留的日子，在 加低斯 停留了許多日子。」
DEUT|2|1|「我們轉回，從 紅海 的路往曠野去，正如耶和華所吩咐我的。我們在 西珥山 繞行了許多日子。
DEUT|2|2|耶和華對我說：
DEUT|2|3|『你們繞行這山已經夠久了，要轉向北方。
DEUT|2|4|你要吩咐百姓說：你們弟兄 以掃 的子孫住在 西珥 ，你們要經過他們的邊界。他們必懼怕你們，但你們要分外謹慎。
DEUT|2|5|不可向他們挑戰；他們的地，連腳掌可踏之處，我都不給你們，因我已將 西珥山 賜給 以掃 為業。
DEUT|2|6|你們要用錢向他們買糧吃，也要用錢向他們買水喝。
DEUT|2|7|因為耶和華─你的上帝在你手裏所做的一切事上已賜福給你。你走這大曠野，他都知道。這四十年，耶和華─你的上帝與你同在，因此你一無所缺。』
DEUT|2|8|「於是，我們經過我們弟兄 以掃 子孫所住的 西珥 ，從 亞拉巴 的路，經過 以拉他 、 以旬‧迦別 ，轉向 摩押 曠野的路去。
DEUT|2|9|耶和華對我說：『不可侵犯 摩押 ，也不可向他們挑戰。他們的地，我不賜給你為業，因我已將 亞珥 賜給 羅得 的子孫為業。』
DEUT|2|10|先前， 以米 人住在那裏，百姓又大又多，像 亞衲 人一樣高大。
DEUT|2|11|他們跟 亞衲 人一樣，也算是 利乏音 人，但 摩押 人卻稱他們為 以米 人。
DEUT|2|12|從前， 何利 人也住在 西珥 ，但 以掃 的子孫把他們除滅，佔領了他們的地，接續他們在那裏居住，如同 以色列 在耶和華賜給他們為業之地所做的一樣。
DEUT|2|13|『現在，起來，過 撒烈溪 ！』於是我們過了 撒烈溪 。
DEUT|2|14|從離開 加低斯‧巴尼亞 到渡過 撒烈溪 ，這段時期共三十八年，直到這一代的戰士都從營中滅盡，正如耶和華向他們所起的誓。
DEUT|2|15|耶和華的手也攻擊他們，將他們從營中除滅，直到滅盡。
DEUT|2|16|「百姓中所有的戰士滅盡死亡以後，
DEUT|2|17|耶和華吩咐我說：
DEUT|2|18|『你今日要經過 摩押 的邊界 亞珥 ，
DEUT|2|19|走到 亞捫 人之地。不可侵犯他們，也不可向他們挑戰。 亞捫 人的地，我不賜給你們為業，因我已將那地賜給 羅得 的子孫為業。』
DEUT|2|20|那地也算是 利乏音 人之地，因為先前 利乏音 人住在那裏， 亞捫 人稱他們為 散送冥 人。
DEUT|2|21|那裏的百姓又大又多，像 亞衲 人一樣高大，但耶和華從 亞捫 人面前除滅他們， 亞捫 人就佔領他們的地，接續他們在那裏居住。
DEUT|2|22|這正如耶和華從前為住在 西珥 的 以掃 子孫，將 何利 人從他們面前除滅，使他們得了 何利 人的地，接續他們在那裏居住，直到今日一樣。
DEUT|2|23|亞衛 人先前住在鄉村直到 迦薩 ；從 迦斐託 出來的 迦斐託 人將 亞衛 人除滅，接續他們在那裏居住。
DEUT|2|24|你們起來往前去，過 亞嫩谷 。看哪，我已將 亞摩利 人 希實本 王 西宏 和他的地交在你手中，你要開始去得他的地為業，向他挑戰。
DEUT|2|25|從今日起，我要讓天下萬民因你驚慌懼怕，聽見你的名聲，就因你發顫傷慟。」
DEUT|2|26|「我從 基底莫 的曠野派遣使者到 希實本 王 西宏 那裏，用和平的話說：
DEUT|2|27|『求你讓我穿越你的地，我走路的時候，只走大路，不偏左右。
DEUT|2|28|你可以賣糧給我吃，賣水給我喝；只要讓我步行過去，
DEUT|2|29|就如住在 西珥 的 以掃 子孫和住在 亞珥 的 摩押 人待我一樣，等我過了 約旦河 ，進入耶和華－我們上帝所賜給我們的地。』
DEUT|2|30|但 希實本 王 西宏 不肯讓我們從他那裏經過，因為耶和華－你的上帝使他性情頑梗，內心剛硬，為要把他交在你手中，像今日一樣。
DEUT|2|31|耶和華對我說：『看，我已開始把 西宏 和他的地交給你了，你要開始得他的地為業。』
DEUT|2|32|「 西宏 和他的眾百姓出來迎擊我們，在 雅雜 與我們交戰。
DEUT|2|33|耶和華－我們的上帝把他交給我們，我們就殺了他和他的眾兒子，以及他所有的百姓。
DEUT|2|34|那時，我們奪了他一切的城鎮，毀滅各城的男人、女人、孩子，沒有留下一個倖存者。
DEUT|2|35|只有牲畜和所奪各城的財物，我們都取為自己的掠物。
DEUT|2|36|從 亞嫩谷 旁的 亞羅珥 和谷中的城，直到 基列 ，沒有一座城是高得我們不能攻取的；耶和華－我們的上帝把它們全都交給我們了。
DEUT|2|37|只有 亞捫 人之地， 雅博河 沿岸，以及山區的城鎮，你沒有挨近，這全是耶和華－我們上帝所吩咐的。」
DEUT|3|1|「我們又轉回，朝 巴珊 的路上去。 巴珊 王 噩 和他的眾百姓出來迎擊我們，在 以得來 與我們交戰。
DEUT|3|2|耶和華對我說：『不要怕他！因我已把他和他的眾百姓，以及他的地，都交在你手中；你要待他像從前待住在 希實本 的 亞摩利 王 西宏 一樣。』
DEUT|3|3|於是耶和華－我們的上帝也把 巴珊 王 噩 和他的眾百姓都交在我們手中；我們殺了他，沒有給他留下一個倖存者。
DEUT|3|4|那時，我們奪了他一切的城鎮，共六十座，沒有一座城不被我們所奪，這是 亞珥歌伯 的全境， 巴珊 王 噩 的國度。
DEUT|3|5|這些堅固的城都有高的城牆，有門有閂，此外，還有許多無城牆的鄉村。
DEUT|3|6|我們把這些都毀滅了，像從前待 希實本 王 西宏 一樣，毀滅各城的男人、女人、孩子；
DEUT|3|7|只有一切牲畜和城中的財物，我們取為自己的掠物。
DEUT|3|8|那時，我們從兩個 亞摩利 王的手裏把 約旦河 東邊的地奪過來，從 亞嫩谷 直到 黑門山 ，
DEUT|3|9|這 黑門山 ， 西頓 人稱為 西連 ， 亞摩利 人稱為 示尼珥 。
DEUT|3|10|我們奪了平原的各城、 基列 全地、 巴珊 全地，直到 撒迦 和 以得來 ，都是 巴珊 王 噩 國內的城鎮。
DEUT|3|11|利乏音 人所剩下的只有 巴珊 王 噩 。看哪，他的床是鐵床，按照人肘的度量，長九肘，寬四肘，現今不是在 亞捫 人的 拉巴 嗎？」
DEUT|3|12|「那時，我們得了這地。從 亞嫩谷 旁的 亞羅珥 起，連同 基列 山區的一半和境內的城鎮，我都給了 呂便 人和 迦得 人。
DEUT|3|13|基列 其餘的地和 巴珊 全地，就是 噩 的國度，我給了 瑪拿西 半支派。 亞珥歌伯 全境就是 巴珊 全地，也稱為 利乏音 人之地。
DEUT|3|14|瑪拿西 的子孫 睚珥 佔領了 亞珥歌伯 全境，直到 基述 人和 瑪迦 人的邊界，就按自己的名字稱這些地，就是 巴珊 ，為 哈倭特‧睚珥 ，直到今日。
DEUT|3|15|我又將 基列 給了 瑪吉 。
DEUT|3|16|我給了 呂便 人和 迦得 人從 基列 到 亞嫩谷 ，以谷的中央為界，直到 亞捫 人邊界的 雅博河 ；
DEUT|3|17|還有 亞拉巴 和靠近 約旦河 之地，從 基尼烈 直到 亞拉巴海 ，就是 鹽海 ，以及 毗斯迦山 斜坡的山腳東邊之地。
DEUT|3|18|「那時，我吩咐你們說：『耶和華－你們的上帝已將這地賜給你們為業；你們所有的勇士都要帶著兵器，在你們的弟兄 以色列 人前面過去。
DEUT|3|19|但你們的妻子、孩子、牲畜，可以住在我所賜給你們的各城裏，我知道你們有許多牲畜。
DEUT|3|20|等到耶和華讓你們的弟兄像你們一樣，得享太平，他們在 約旦河 另一邊，也得了耶和華－你們的上帝所賜給他們的地，你們各人才可以回到我所賜給你們為業之地。』
DEUT|3|21|那時，我吩咐 約書亞 說：『你親眼看見了耶和華－你們的上帝向這兩個王一切所做的事，耶和華也必向你所要去的各國照樣做。
DEUT|3|22|不要怕他們，因為那為你們爭戰的是耶和華－你們的上帝。』」
DEUT|3|23|「那時，我懇求耶和華說：
DEUT|3|24|『主耶和華啊，你已開始將你的偉大和你大能的手顯給你僕人看。在天上，在地下，有甚麼神明能像你行事，像你有大能的作為呢？
DEUT|3|25|求你讓我過去，看 約旦河 另一邊的美地，就是那佳美的山區和 黎巴嫩 。』
DEUT|3|26|但耶和華因你們的緣故向我發怒，不應允我。耶和華對我說：『你夠了吧！不要再向我提這事。
DEUT|3|27|你上 毗斯迦山 頂去，向東、西、南、北舉目，用你的眼睛觀看，因為你必不能過這 約旦河 。
DEUT|3|28|你卻要吩咐 約書亞 ，勉勵他，使他壯膽，因為他必在這百姓前面過去，使他們承受你所要觀看之地。』
DEUT|3|29|於是我們停留在 伯‧毗珥 對面的谷中。」
DEUT|4|1|「現在， 以色列 啊，聽我所教導你們的律例典章，要遵行，好使你們存活，得以進入耶和華－你們列祖之上帝所賜給你們的地，承受為業。
DEUT|4|2|我吩咐你們的話，你們不可加添，也不可刪減，好叫你們遵守耶和華－你們上帝的命令，就是我所吩咐你們的。
DEUT|4|3|你們已親眼看見耶和華因 巴力‧毗珥 所做的。凡隨從 巴力‧毗珥 的人，耶和華－你的上帝都從你中間除滅了。
DEUT|4|4|只有你們這緊緊跟隨耶和華－你們上帝的人，今日全都存活。
DEUT|4|5|看，我照著耶和華－我的上帝所吩咐我的，將律例和典章教導你們，使你們在所要進去得為業的地上遵行。
DEUT|4|6|你們要謹守遵行；這就是你們在萬民眼前的智慧和聰明。他們聽見這一切律例，必說：『這大國的人真是有智慧，有聰明！』
DEUT|4|7|哪一大國有神明與他們相近，像耶和華－我們的上帝在我們求告他的時候與我們相近呢？
DEUT|4|8|哪一大國有這樣公義的律例典章，像我今日在你們面前所頒佈的這一切律法呢？
DEUT|4|9|「但你要謹慎，殷勤保守你的心靈，免得忘記你親眼所看見的事，又免得在你一生的年日這些事離開你的心，總要把它們傳給你的子子孫孫。
DEUT|4|10|你在 何烈山 站在耶和華－你上帝面前的那日，耶和華對我說：『你為我召集百姓，我要叫他們聽見我的話，使他們活在世上的日子，可以學習敬畏我，又可以教導他們的兒女。』
DEUT|4|11|那時，你們近前來，站在山下；山上有火燃燒，直沖天頂，並有黑暗、密雲、幽暗。
DEUT|4|12|耶和華從火焰中對你們說話，你們聽見說話的聲音，只有聲音，卻沒有看見形像。
DEUT|4|13|他將所吩咐你們當守的約指示你們，就是十條誡命 ，並將誡命寫在兩塊石版上。
DEUT|4|14|那時，耶和華吩咐我將律例典章教導你們，使你們在所要過去得為業的地上遵行。」
DEUT|4|15|「所以，你們為自己的緣故要分外謹慎；因為耶和華在 何烈山 ，從火中對你們說話的那日，你們沒有看見任何形像。
DEUT|4|16|惟恐你們的行為敗壞，為自己雕刻任何形狀的偶像，無論是男像或女像，
DEUT|4|17|或地上任何走獸的像，或任何飛在空中有翅膀的鳥的像，
DEUT|4|18|或地上任何爬行動物的像，或地底下任何水中魚的像。
DEUT|4|19|又恐怕你向天舉目，看見耶和華－你的上帝為天下萬民所擺列的日月星辰，就是天上的萬象，就被誘惑去敬拜它們，事奉它們。
DEUT|4|20|耶和華將你們從 埃及 帶領出來，脫離鐵爐，是要你們成為他產業的子民，像今日一樣。
DEUT|4|21|「耶和華又因你們的緣故向我發怒，起誓不容我過 約旦河 ，不讓我進入耶和華－你上帝所賜你為業的那美地。
DEUT|4|22|我只好死在這地，不能過 約旦河 ；但你們必過去得那美地。
DEUT|4|23|你們要謹慎，免得忘記耶和華－你們的上帝與你們所立的約，為自己雕刻任何形狀的偶像，就是耶和華－你上帝所禁止的，
DEUT|4|24|因為耶和華－你的上帝是吞滅的火，是忌邪 的上帝。
DEUT|4|25|「你們在那地住久了，生子生孫，若行為敗壞，為自己雕刻任何形狀的偶像，行耶和華－你上帝眼中看為惡的事，惹他發怒，
DEUT|4|26|我今日呼天喚地向你們作見證，你們在過 約旦河 得為業的地上必迅速滅亡！你們在那地的日子必不長久，必全然滅絕。
DEUT|4|27|耶和華必將你們分散在萬民中；在耶和華領你們到的列國中，你們剩下的人丁稀少。
DEUT|4|28|在那裏，你們必事奉人手所造的神明，它們是木頭，是石頭，不能看，不能聽，不能吃，不能聞。
DEUT|4|29|你們在那裏必尋求耶和華－你的上帝。你若盡心盡性尋求他，就必尋見。
DEUT|4|30|日後你在患難中，當這一切的事臨到你，你必歸回耶和華－你的上帝，聽從他的話。
DEUT|4|31|耶和華－你的上帝是有憐憫的上帝，他不撇下你，不滅絕你，也不忘記他起誓與你列祖所立的約。
DEUT|4|32|「你去問，在你先前的時代，自從上帝造人在地上以來，從天這邊到天那邊，曾有過或聽過這樣的大事嗎？
DEUT|4|33|有哪些百姓聽見上帝在火中說話的聲音，像你聽見了還能存活呢？
DEUT|4|34|上帝何曾為自己嘗試從別的國中領出一國的子民來，用考驗、神蹟、奇事、戰爭、大能的手、伸出來的膀臂和大可畏的事，像耶和華－你們的上帝在 埃及 ，在你們眼前為你們所做的一切事呢？
DEUT|4|35|這是要顯給你看，使你知道，惟有耶和華他是上帝，除他以外，再沒有別的了。
DEUT|4|36|他從天上使你聽見他的聲音，為要教導你，又在地上使你看見他的烈火，並且聽見他從火中所說的話。
DEUT|4|37|因為他愛你的列祖，揀選他們的後裔 ，親自用大能領你出了 埃及 ，
DEUT|4|38|要將比你強大的列國從你面前趕出，領你進去，把他們的地賜你為業，像今日一樣。
DEUT|4|39|所以，今日你要知道，也要記在心裏，天上地下惟有耶和華他是上帝，再沒有別的了。
DEUT|4|40|我今日吩咐你的律例誡命，你要遵守，使你和你的後裔可以得福，並使你的日子一直在耶和華－你上帝賜你的地上得以長久。」
DEUT|4|41|「那時， 摩西 在 約旦河 東邊，向日出的方向，指定三座城，
DEUT|4|42|使那素無仇恨、無意中殺了鄰舍的兇手，可以逃到這三座城中的一座，就得存活：
DEUT|4|43|屬 呂便 人的是曠野平坦之地的 比悉 ，屬 迦得 人的是 基列 的 拉末 ，屬 瑪拿西 人的是 巴珊 的 哥蘭 。」
DEUT|4|44|這是 摩西 在 以色列 人面前頒佈的律法。
DEUT|4|45|這些法度、律例、典章是 摩西 在 以色列 人出 埃及 後對他們說的，
DEUT|4|46|在 約旦河 東 伯毗珥 對面的谷中，在住 希實本 的 亞摩利 王 西宏 之地；這 西宏 是 摩西 和 以色列 人出 埃及 後所擊殺的。
DEUT|4|47|他們得了他的地，又得了 巴珊 王 噩 的地，就是兩個 亞摩利 王，在 約旦河 東，向日出方向的地：
DEUT|4|48|從 亞嫩谷 旁的 亞羅珥 ，直到 西雲山 ，就是 黑門山 ，
DEUT|4|49|還有 約旦河 東的整個 亞拉巴 ，向日出方向，直到 亞拉巴海 ，靠近 毗斯迦山 斜坡的山腳。
DEUT|5|1|摩西 召集 以色列 眾人，對他們說：「 以色列 啊，要聽我今日在你們耳中所吩咐的律例典章，要學習，謹守遵行。
DEUT|5|2|耶和華－我們的上帝在 何烈山 與我們立約。
DEUT|5|3|這約耶和華不是與我們列祖立的，而是與我們，就是今日在這裏還活著的人立的。
DEUT|5|4|耶和華在山上，從火中，面對面與你們說話。
DEUT|5|5|那時我站在耶和華和你們之間，要將耶和華的話傳給你們，因為你們懼怕那火，沒有上山。他說：
DEUT|5|6|「『我是耶和華－你的上帝，曾將你從 埃及 地為奴之家領出來。
DEUT|5|7|「『除了我以外，你不可有別的神。
DEUT|5|8|「『不可為自己雕刻偶像，也不可做甚麼形像，彷彿上天、下地和地底下水中的百物。
DEUT|5|9|不可跪拜那些像，也不可事奉它們，因為我耶和華－你的上帝是忌邪 的上帝。恨我的，我必懲罰他們的罪，自父及子，直到三、四代；
DEUT|5|10|愛我、守我誡命的，我必向他們施慈愛，直到千代。
DEUT|5|11|「『不可妄稱耶和華－你上帝的名，因為妄稱耶和華名的，耶和華必不以他為無罪。
DEUT|5|12|「『當守安息日為聖日，正如耶和華－你上帝所吩咐的。
DEUT|5|13|六日要勞碌做你一切的工，
DEUT|5|14|但第七日是向耶和華－你的上帝當守的安息日。這一日，你和你的兒女、僕婢、牛、驢、牲畜，以及你城裏寄居的客旅，都不可做任何的工，使你的僕婢可以和你一樣休息。
DEUT|5|15|你要記念你在 埃及 地作過奴僕，耶和華－你的上帝用大能的手和伸出來的膀臂領你從那裏出來。因此，耶和華－你的上帝吩咐你守安息日。
DEUT|5|16|「『當孝敬父母，正如耶和華－你上帝所吩咐的，使你得福，並使你的日子在耶和華－你上帝所賜給你的地上得以長久。
DEUT|5|17|「『不可殺人。
DEUT|5|18|「『不可姦淫。
DEUT|5|19|「『不可偷盜。
DEUT|5|20|「『不可做假見證陷害你的鄰舍。
DEUT|5|21|「『不可貪戀你鄰舍的妻子；也不可貪圖你鄰舍的房屋、田地、僕婢、牛驢，以及他一切所有的。』
DEUT|5|22|「這些話是耶和華在山上，從火焰、密雲、幽暗中，大聲吩咐你們全會眾的，再沒有加添別的話了。他把這些話寫在兩塊石版上，交給我。
DEUT|5|23|山被火焰燒著，你們聽見從黑暗中發出的聲音，那時，你們各支派的領袖和長老都挨近我。
DEUT|5|24|你們說：『看哪，耶和華－我們的上帝將他的榮耀和他的偉大顯給我們看，我們也聽見他從火中發出的聲音。今日我們看到上帝與人說話，人還活著。
DEUT|5|25|現在這大火將要吞滅我們，我們何必死呢？若再聽見耶和華我們上帝的聲音，我們就必死。
DEUT|5|26|凡血肉之軀，有誰像我們一樣，聽見了永生上帝從火中講話的聲音還能活著呢？
DEUT|5|27|求你近前去，聽耶和華－我們上帝所要說的一切話，將耶和華－我們上帝對你說的話都傳給我們，我們就聽從遵行。』
DEUT|5|28|「你們對我說的話，耶和華都聽見了。耶和華對我說：『這百姓對你說的話，我聽見了；他們所說的都對。
DEUT|5|29|惟願他們存這樣的心敬畏我，常遵守我一切的誡命，使他們和他們的子孫永遠得福。
DEUT|5|30|你去對他們說：你們回帳棚去吧！
DEUT|5|31|至於你，可以站在我這裏，我要將一切誡命、律例、典章傳給你。你要教導他們，使他們在我賜他們為業的地上遵行。』
DEUT|5|32|所以，你們要照耶和華－你們上帝所吩咐的謹守遵行，不可偏離左右。
DEUT|5|33|你們要走耶和華－你們的上帝所吩咐的一切道路，使你們可以存活得福，並使你們的日子在所要承受的地上得以長久。」
DEUT|6|1|「這是耶和華－你們的上帝所吩咐要教導你們的誡命、律例、典章，叫你們在所要過去得為業的地上遵行，
DEUT|6|2|好叫你和你的子孫在一生的日子都敬畏耶和華－你的上帝，謹守他的一切律例、誡命，就是我所吩咐你的，使你的日子得以長久。
DEUT|6|3|以色列 啊，你要聽，要謹守遵行，使你可以在那流奶與蜜之地得福，人數極其增多，正如耶和華－你列祖的上帝所應許你的。
DEUT|6|4|「 以色列 啊，你要聽！耶和華－我們的上帝是獨一的主 。
DEUT|6|5|你要盡心、盡性、盡力愛耶和華－你的上帝。
DEUT|6|6|我今日吩咐你的這些話都要記在心上，
DEUT|6|7|也要殷勤教導你的兒女。無論你坐在家裏，走在路上，躺下，起來，都要吟誦。
DEUT|6|8|要繫在手上作記號，戴在額上 作經匣 ；
DEUT|6|9|又要寫在你房屋的門框上和你的城門上。
DEUT|6|10|「耶和華－你的上帝必領你進他向你列祖 亞伯拉罕 、 以撒 、 雅各 起誓要給你的地。那裏有又大又美的城鎮，不是你建造的；
DEUT|6|11|有裝滿各樣美物的房屋，不是你裝滿的；有挖成的水井，不是你挖的；有葡萄園、橄欖園，不是你栽植的；你吃了而且飽足。
DEUT|6|12|你要謹慎，免得你忘記領你從 埃及 地為奴之家出來的耶和華。
DEUT|6|13|你要敬畏耶和華－你的上帝，事奉他，奉他的名起誓。
DEUT|6|14|不可隨從別神，就是你們四圍民族的眾神明，
DEUT|6|15|因為在你中間的耶和華－你的上帝是忌邪 的上帝，恐怕耶和華－你上帝的怒氣向你發作，把你從地上除滅。
DEUT|6|16|「你們不可試探耶和華－你們的上帝，像你們在 瑪撒 那樣試探他。
DEUT|6|17|要謹慎遵守耶和華－你們上帝的誡命，和他所吩咐的法度、律例。
DEUT|6|18|耶和華眼中看為正直和美善的事，你都要遵行，使你得福，可以進去得耶和華向你列祖起誓應許的美地，
DEUT|6|19|可以從你面前趕出你所有的仇敵，正如耶和華所說的。
DEUT|6|20|「日後，你的兒子問你說：『耶和華－我們上帝吩咐你們的法度、律例、典章是甚麼意思呢？』
DEUT|6|21|你要告訴你的兒子說：『我們在 埃及 作過法老的奴僕，耶和華用大能的手將我們從 埃及 領出來。
DEUT|6|22|在我們眼前，他施行重大可怕的神蹟奇事對付 埃及 、法老和他的全家。
DEUT|6|23|他將我們從那裏領出來，為要領我們進入他向我們列祖起誓應許之地，把這地賜給我們。
DEUT|6|24|耶和華又吩咐我們遵行這一切的律例，敬畏耶和華－我們的上帝，使我們一生得福，得以存活，像今日一樣。
DEUT|6|25|我們若照耶和華－我們上帝所吩咐的，在他面前謹守遵行這一切誡命，這就是我們的義了。』」
DEUT|7|1|「耶和華－你的上帝領你進入你要得為業之地，從你面前趕出許多國家，就是比你更強大的七個國家： 赫 人、 革迦撒 人、 亞摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人。
DEUT|7|2|當耶和華－你的上帝把他們交給你，你擊殺他們的時候，你要完全消滅他們，不可與他們立約，也不可憐惜他們。
DEUT|7|3|不可與他們結親；不可將你的女兒嫁給他的兒子，也不可叫你的兒子娶他的女兒。
DEUT|7|4|因為他必使你的兒女離棄我，去事奉別神，以致耶和華的怒氣向你們發作，迅速將你除滅。
DEUT|7|5|你們卻要這樣處置他們：拆毀他們的祭壇，打碎他們的柱像，砍斷他們的 亞舍拉 ，用火焚燒他們雕刻的偶像。
DEUT|7|6|「因為你是屬於耶和華－你上帝神聖的子民；耶和華－你的上帝從地面上的萬民中揀選你，作自己寶貴的子民。
DEUT|7|7|耶和華專愛你們，揀選你們，並非因你們人數比任何民族多，其實你們的人數在各民族中是最少的。
DEUT|7|8|因為耶和華愛你們，又因要遵守他向你們列祖所起的誓，耶和華就用大能的手領你們出來，救贖你脫離為奴之家，脫離 埃及 王法老的手。
DEUT|7|9|所以，你知道耶和華－你的上帝，他是上帝，是信實的上帝。他向愛他、守他誡命的人守約施慈愛，直到千代；
DEUT|7|10|向恨他的人，他必當面報應，消滅他們。凡恨他的，他必當面報應，絕不遲延。
DEUT|7|11|所以，你要謹守我今日所吩咐你的誡命、律例、典章，遵行它們。」
DEUT|7|12|「你們若聽從這些典章，謹守遵行，耶和華－你的上帝必照他向你列祖所起的誓，對你守約，施慈愛。
DEUT|7|13|他必愛你，賜福給你，使你人數增多，也必在他向你列祖起誓要給你的地上賜福給你身所生的，你地所產的，你的五穀、新酒和新的油，以及你的牛犢、羔羊。
DEUT|7|14|你必蒙福勝過萬民；你沒有不育的男人和不孕的女人，牲畜也沒有不生育的。
DEUT|7|15|耶和華必使一切的疾病遠離你；你所知道 埃及 各樣的惡疾，他不加在你身上，反要加在所有恨你的人身上。
DEUT|7|16|你要吞滅耶和華－你的上帝交給你的各民族，你的眼目不可顧惜他們。你也不可事奉他們的神明，因為這必成為你的圈套。
DEUT|7|17|「你若心裏說，這些國的人數比我多，我怎能趕出他們呢？
DEUT|7|18|你不必怕他們，要牢牢記住耶和華－你上帝向法老和 埃及 全地所行的事，
DEUT|7|19|你親眼見過的大考驗、神蹟、奇事、大能的手和伸出來的膀臂，都是耶和華－你上帝領你出來所施行的。耶和華－你的上帝也必照樣處置你所懼怕的各民族，
DEUT|7|20|並且耶和華－你的上帝必派瘟疫 攻擊他們，直到那剩下而躲起來的人都從你面前滅亡。
DEUT|7|21|不要因他們驚恐，因為耶和華－你的上帝在你中間是大而可畏的上帝。
DEUT|7|22|耶和華－你的上帝必將這些國從你面前漸漸趕出；你不可迅速把他們消滅，免得野地的走獸多起來危害你。
DEUT|7|23|耶和華－你的上帝必將他們交給你，大大擾亂他們，直到他們被除滅。
DEUT|7|24|他又要將他們的君王交在你手中，你必從天下除去他們的名；必無一人能在你面前站立得住，直到你把他們除滅了。
DEUT|7|25|你們要用火焚燒他們神明的雕刻偶像；不可貪愛偶像上的金銀，也不可私自收起來，免得你因此陷入圈套，因為這是耶和華－你上帝所憎惡的。
DEUT|7|26|你不可把可憎之物帶進你的家，否則，你就像它一樣成為當毀滅的。你要徹底憎恨它，極其厭惡它，因為這是當毀滅的。」
DEUT|8|1|「我今日所吩咐你的一切誡命，你們要謹守遵行，好使你們存活，人數增多，可以進去得耶和華向你們列祖起誓應許的那地。
DEUT|8|2|你要記得，這四十年耶和華─你的上帝在曠野一路引導你，是要磨煉你，考驗你，為要知道你的心如何，是否願意遵守他的誡命。
DEUT|8|3|他磨煉你，任你飢餓，將你和你列祖所不認識的嗎哪賜給你吃，使你知道，人活著，不是單靠食物，乃是靠耶和華口裏所出的一切話。
DEUT|8|4|這四十年，你身上的衣服沒有穿破，你的腳也沒有腫。
DEUT|8|5|你心裏要知道，耶和華─你的上帝管教你，像人管教兒女一樣。
DEUT|8|6|你要謹守耶和華─你上帝的誡命，遵行他的道，敬畏他。
DEUT|8|7|「耶和華─你的上帝必領你進入美地，那地有河流，有泉源和深淵的水從谷中和山上流出。
DEUT|8|8|那地有小麥、大麥、葡萄樹、無花果樹、石榴樹，那地也有橄欖油和蜂蜜。
DEUT|8|9|那地沒有缺乏，你在那裏有食物吃，一無所缺；那地的石頭是鐵，山中可以挖銅。
DEUT|8|10|你吃得飽足，要稱頌耶和華─你的上帝，因為他將那美地賜給你。」
DEUT|8|11|「你要謹慎，免得忘記耶和華─你的上帝，不守他的誡命、典章、律例，就是我今日吩咐你的。
DEUT|8|12|免得你吃得飽足，建造上好的房屋，住在其中，
DEUT|8|13|你的牛羊增多，你的金銀增多，你擁有的一切全都增多，
DEUT|8|14|於是你的心高傲，忘記耶和華─你的上帝。他曾將你從 埃及 地為奴之家領出來，
DEUT|8|15|曾引領你經過那大而可怕的曠野，有火蛇、蠍子、乾旱無水之地。他也曾為你使水從堅硬的磐石中流出來，
DEUT|8|16|又在曠野將你列祖所不認識的嗎哪賜給你吃，為要磨煉你，考驗你，終久使你享福。
DEUT|8|17|你心裏說：『這財富是我的力量、我手的能力得來的。』
DEUT|8|18|你要記得耶和華─你的上帝，因為得財富的能力是他給你的，為要堅守他向你列祖起誓所立的約，像今日一樣。
DEUT|8|19|你若忘記耶和華─你的上帝，隨從別神，事奉它們，敬拜它們，我今日警告你們，你們必定滅亡。
DEUT|8|20|耶和華在你們面前怎樣使列國滅亡，你們也必照樣滅亡，因為你們不聽從耶和華─你們上帝的話。」
DEUT|9|1|「 以色列 啊，你要聽！你今日要過 約旦河 ，進去佔領比你更強大的列國，那裏的城鎮又大，城牆又堅固，如天一樣高。
DEUT|9|2|那裏的百姓是 亞衲 族人，又高又壯，是你所知道的；你也聽說過：『誰能在 亞衲 族人面前站立得住呢？』
DEUT|9|3|你今日應當知道，耶和華─你的上帝在你前面渡過去，如同吞噬的火，要除滅他們，並要在你面前將他們制伏，使你可以趕出他們，速速消滅他們，正如耶和華向你所說的。
DEUT|9|4|「耶和華─你的上帝將他們從你面前趕出以後，你心裏不可說：『耶和華領我得這地是因我的義。』其實，耶和華將這些國家從你面前趕出去是因他們的惡。
DEUT|9|5|你能進去得他們的地，並不是因你的義，也不是因你心裏正直，而是因這些國家的惡，耶和華─你的上帝才把他們從你面前趕出去，為了應驗耶和華向你列祖 亞伯拉罕 、 以撒 、 雅各 起誓應許的話。
DEUT|9|6|「你當知道，耶和華─你的上帝將這美地賜你為業，並不是因你的義；你本是硬著頸項的百姓。
DEUT|9|7|你要記得，不要忘記，你在曠野怎樣惹耶和華－你的上帝發怒。自從你出了 埃及 地的那日，直到你們來到這地方，你們常常悖逆耶和華。
DEUT|9|8|你們在 何烈山 惹耶和華發怒，耶和華對你們動怒，甚至要除滅你們。
DEUT|9|9|我上了山，要領受兩塊石版，就是耶和華與你們立約的版。那時我在山上住了四十晝夜，沒有吃飯，也沒有喝水。
DEUT|9|10|耶和華把那兩塊石版交給我，是上帝用指頭寫成的；版上是耶和華在大會的那一天，在山上從火中對你們所說的一切話。
DEUT|9|11|過了四十晝夜，耶和華把那兩塊石版，就是約版，交給我。
DEUT|9|12|耶和華對我說：『起來，趕快從這裏下去！因為你從 埃及 領出來的百姓已經敗壞了；他們這麼快偏離了我所吩咐的道，為自己鑄造偶像。』
DEUT|9|13|「耶和華對我說：『我看這百姓，看哪，他們是硬著頸項的百姓。
DEUT|9|14|你且由著我，我要除滅他們，從天下塗去他們的名，我要使你成為比他們更大更強的國。』
DEUT|9|15|於是我轉身下山，山上有火燃燒，兩塊約版在我雙手中。
DEUT|9|16|我觀看，看哪，你們得罪了耶和華－你們的上帝，為自己鑄成了一頭牛犢，迅速偏離了耶和華所吩咐你們的道，
DEUT|9|17|我拿著那兩塊石版，從我雙手中扔出去，在你們眼前把它們摔碎了。
DEUT|9|18|因為你們所犯的一切罪，做了耶和華眼中看為惡的事，惹他發怒，我就像從前一樣俯伏在耶和華面前四十晝夜，沒有吃飯，沒有喝水。
DEUT|9|19|我很害怕，因為耶和華向你們大發烈怒，要除滅你們。但那一次耶和華又應允了我。
DEUT|9|20|耶和華也向 亞倫 非常生氣，甚至要除滅他；那時我也為 亞倫 祈禱。
DEUT|9|21|我把那使你們犯罪所鑄的牛犢拿來，用火焚燒，搗碎後再磨成粉末，好像灰塵。我把這灰塵撒在從山上流下來的溪水中。
DEUT|9|22|「你們在 他備拉 、 瑪撒 、 基博羅‧哈他瓦 又惹耶和華發怒。
DEUT|9|23|耶和華叫你們離開 加低斯‧巴尼亞 ，說：『你們上去得我所賜給你們的地。』那時，你們違背了耶和華－你們上帝的指示，不信服他，不聽從他的話。
DEUT|9|24|自從我認識你們的日子以來，你們常常悖逆耶和華。
DEUT|9|25|「我因耶和華說要除滅你們，就在耶和華面前俯伏四十晝夜，像我以前俯伏一樣。
DEUT|9|26|我向耶和華祈禱，說：『主耶和華啊，求你不要滅絕你的百姓，你的產業。他們是你用大能救贖，用你強有力的手從 埃及 領出來的。
DEUT|9|27|求你記念你的僕人 亞伯拉罕 、 以撒 、 雅各 ，不看這百姓的頑梗、邪惡、罪愆，
DEUT|9|28|免得你領我們出來的那地之人說：耶和華因為不能將這百姓領進他所應許之地，又因恨他們，所以領他們出去，要在曠野殺他們。
DEUT|9|29|其實他們是你的百姓，你的產業，是你用大能和伸出的膀臂領出來的。』」
DEUT|10|1|「那時，耶和華對我說：『你要鑿出兩塊石版，和先前的一樣，上山到我這裏來。你也要造一個木櫃。
DEUT|10|2|我要把你先前摔碎的版上所寫的字，寫在這版上；你要把這版放在櫃裏。』
DEUT|10|3|於是我用金合歡木造了一個櫃子，又鑿出兩塊石版，和先前的一樣。我手裏拿著這兩塊版上山。
DEUT|10|4|耶和華將那大會之日、在山上從火中所吩咐你們的十條誡命，照先前所寫的寫在這版上。耶和華把它們交給我。
DEUT|10|5|我轉身下山，將這版放在我所造的櫃裏，現今這版還在那裏，正如耶和華所吩咐我的。
DEUT|10|6|（ 以色列 人從 比羅比尼‧亞干 起行，來到 摩西拉 ， 亞倫 死在那裏，就葬在那裏。他的兒子 以利亞撒 接續他擔任祭司的職分。
DEUT|10|7|他們從那裏起行，來到 谷歌大 ，又從 谷歌大 來到 約巴他 ，有溪水之地。
DEUT|10|8|那時，耶和華將 利未 支派分別出來，抬耶和華的約櫃，又侍立在耶和華面前事奉他，奉他的名祝福，直到今日。
DEUT|10|9|因此， 利未 沒有像他的弟兄有產業，耶和華是他的產業，正如耶和華－你上帝所應許他的。）
DEUT|10|10|「我又像先前一樣在山上停留了四十晝夜。這一次耶和華也應允我，不將你滅絕。
DEUT|10|11|耶和華對我說：『起來，走在百姓前面，領他們進去得我向他們列祖起誓要給他們的地。』」
DEUT|10|12|「 以色列 啊，現在耶和華－你的上帝向你要的是甚麼呢？只要你敬畏耶和華－你的上帝，遵行他一切的道，愛他，盡心盡性事奉耶和華－你的上帝，
DEUT|10|13|遵守耶和華的誡命律例，就是我今日所吩咐你的，為要使你得福。
DEUT|10|14|看哪，天和天上的天，地和地上所有的，都屬耶和華－你的上帝。
DEUT|10|15|然而，耶和華專愛你的列祖，愛他們，從萬民中揀選你們，就是他們的後裔，像今日一樣。
DEUT|10|16|所以你們的心要受割禮，不可再硬著頸項。
DEUT|10|17|因為耶和華－你們的上帝是萬神之神，萬主之主，是偉大、強有力、可畏的上帝，不看人的情面，也不受賄賂。
DEUT|10|18|他為孤兒寡婦伸冤，愛護寄居的，賜給他衣食。
DEUT|10|19|所以你們要愛護寄居的，因為你們在 埃及 地也作過寄居的。
DEUT|10|20|你要敬畏耶和華－你的上帝，事奉他，緊緊跟隨他，奉他的名起誓。
DEUT|10|21|他是你當讚美的，是你的上帝，為你做了大而可畏的事，這些是你親眼見過的。
DEUT|10|22|你的列祖七十人下 埃及 ，現在耶和華－你的上帝卻使你如同天上的星那樣多。」
DEUT|11|1|「你要愛耶和華－你的上帝，天天遵守他的吩咐、律例、典章、誡命。
DEUT|11|2|今日你們應當知道，而不是你們的兒女，因為他們不知道，也沒有見過耶和華─你們上帝的管教、他的偉大、他大能的手和伸出來的膀臂，
DEUT|11|3|以及他在 埃及 向 埃及 王法老和其全地所行的神蹟奇事；
DEUT|11|4|他怎樣對待 埃及 的軍隊、馬和戰車，他們追趕你們的時候，耶和華怎樣用 紅海 的水淹沒他們，消滅了他們，直到今日；
DEUT|11|5|他在曠野怎樣待你們，直到你們來到這地方，
DEUT|11|6|以及他怎樣待 呂便 子孫， 以利押 的兒子 大坍 、 亞比蘭 ，地怎樣在 以色列 人中開了裂口，吞了他們和他們的家眷，帳棚，以及跟他們在一起所有活著的。
DEUT|11|7|惟有你們親眼見過耶和華所做的一切大事。」
DEUT|11|8|「所以，你們要遵守我今日所吩咐的一切誡命，使你們剛強，可以進去得你們所要得的那地，就是你們將過河到那裏要得的，
DEUT|11|9|也使你們的日子，在耶和華向你們列祖起誓要給他們和他們後裔的地上得以長久，那是流奶與蜜之地。
DEUT|11|10|你要進去得為業的那地，不像你出來的 埃及 地。在 埃及 ，你撒種後，要用腳澆灌，像澆灌菜園一樣。
DEUT|11|11|你們要過去得為業的那地乃是有山有谷、天上的雨水滋潤之地，
DEUT|11|12|是耶和華－你上帝所眷顧的地；從歲首到年終，耶和華－你上帝的眼目時常看顧那地。
DEUT|11|13|「你們若留心聽從我今日所吩咐你們的誡命，愛耶和華－你們的上帝，盡心盡性事奉他，
DEUT|11|14|我 必按時降下雨水在你們的地上，就是秋雨和春雨，使你們可以收藏五穀、新酒和新的油，
DEUT|11|15|也必使田野為你的牲畜長出草來；這樣，你必吃得飽足。
DEUT|11|16|你們要謹慎，免得心受誘惑，轉去事奉別神，敬拜它們，
DEUT|11|17|以致耶和華的怒氣向你們發作，使天封閉不下雨，使地不出產，使你們在耶和華所賜給你們的美地上速速滅亡。
DEUT|11|18|「你們要將我這些話存在心裏，留在意念中，繫在手上作記號，戴在額上 作經匣。
DEUT|11|19|你們也要將這些話教導你們的兒女，無論坐在家裏，行在路上，躺下，起來，都要講論，
DEUT|11|20|又要寫在房屋的門框上和你的城門上。
DEUT|11|21|這樣，你們和你們子孫的日子必在耶和華向你們列祖起誓要給他們的地上得以增多，如天地之長久。
DEUT|11|22|你們若留心謹守遵行我所吩咐這一切的誡命，愛耶和華－你們的上帝，遵行他一切的道，緊緊跟隨他，
DEUT|11|23|他必從你們面前趕出這一切國家，你們也要佔領比你們更大更強的國家。
DEUT|11|24|凡你們腳掌所踏之地都必歸於你們；從曠野到 黎巴嫩 ，從 幼發拉底 大河，直到西邊的海，都要成為你們的疆土。
DEUT|11|25|必無一人能在你們面前站立得住；耶和華－你們的上帝必照他所說的，使懼怕驚恐臨到你們所踏的全地。
DEUT|11|26|「看，我今日將祝福與詛咒都陳明在你們面前。
DEUT|11|27|你們若聽從耶和華─你們上帝的誡命，就是我今日所吩咐你們的，就必蒙福。
DEUT|11|28|你們若不聽從耶和華─你們上帝的誡命，偏離我今日所吩咐你們的道，去隨從你們所不認識的別神，就必受詛咒。
DEUT|11|29|當耶和華－你的上帝領你進入要得為業的那地，你就要在 基利心山 上宣佈祝福，在 以巴路山 上宣佈詛咒。
DEUT|11|30|這二座山豈不是在 約旦河 的那邊，日落的方向，在住 亞拉巴 的 迦南 人之地， 吉甲 的前面，靠近 摩利 橡樹嗎？
DEUT|11|31|你們過 約旦河 ，進去得耶和華－你們的上帝所賜你們為業之地；當你們佔領它，在那地居住的時候，
DEUT|11|32|你們要謹守遵行我今日在你們面前頒佈的一切律例典章。」
DEUT|12|1|「你們活在世上的日子，在耶和華─你列祖的上帝所賜你為業的地上，你們要謹守遵行這些律例典章：
DEUT|12|2|你們佔領的國家所事奉他們眾神明的地方，無論是在高山，在小山，在一切的青翠樹下，你們要徹底毀壞；
DEUT|12|3|要拆毀他們的祭壇，打碎他們的柱像，用火焚燒他們的 亞舍拉 ，砍斷他們神明的雕刻偶像，並要從那地方除去他們的名。
DEUT|12|4|你們不可那樣敬拜耶和華－你們的上帝。
DEUT|12|5|但耶和華－你們的上帝在你們各支派中選擇何處作為立他名的居所，你們就要到那裏求問，
DEUT|12|6|將你們的燔祭、祭物、十一奉獻、手中的舉祭、還願祭、甘心祭，以及牛群羊群中頭生的，都帶到那裏。
DEUT|12|7|在那裏，你們和你們的全家都可以在耶和華─你們上帝的面前吃，並且因你們手所做的一切蒙耶和華－你的上帝賜福而歡樂。
DEUT|12|8|你們不可做像我們今日在這裏所做的，各人行自己眼中看為正的一切事；
DEUT|12|9|因為你們現在還沒有進入耶和華－你上帝所賜你的安息，所給你的產業。
DEUT|12|10|你們過了 約旦河 ，住在耶和華─你們上帝給你們承受為業的地；他又使你們得享太平，不受四圍一切仇敵擾亂，使你們安然居住。
DEUT|12|11|那時你們要將我所吩咐你們的燔祭、祭物、十一奉獻、手中的舉祭，和向耶和華許願的一切上好的祭，都帶到耶和華─你們上帝所選擇立他名的居所。
DEUT|12|12|你們和兒女、僕婢，以及住在你們城裏，沒有與你們一起分得產業的 利未 人，都要在耶和華－你們的上帝面前歡樂。
DEUT|12|13|你要謹慎，不可在自己所看中的各處獻燔祭。
DEUT|12|14|惟獨耶和華從你的一個支派中所選擇的地方，你要在那裏獻燔祭，在那裏遵行我一切所吩咐你的。
DEUT|12|15|「然而，你在各城裏都可以照著耶和華－你上帝所賜給你的福分，隨心所欲宰牲吃肉；無論潔淨的人不潔淨的人都可以吃，就如吃羚羊和鹿的肉一樣。
DEUT|12|16|只是血，你不可吃，要把它倒在地上，如同倒水一樣。
DEUT|12|17|你的五穀、新酒和新油的十分之一，或是牛群羊群中頭生的，或是你的許願祭、甘心祭和手中的舉祭，都不可在你的城裏吃，
DEUT|12|18|必須在耶和華－你的上帝面前吃，在耶和華－你上帝所選擇的地方，你和兒女、僕婢，以及住在你城裏的 利未 人都可以吃，並要因你手所做的一切，在耶和華－你上帝面前歡樂。
DEUT|12|19|你要謹慎，在你所住的地上，你永不可離棄 利未 人。
DEUT|12|20|「耶和華－你的上帝照他的應許擴張你疆土的時候，你心裏想要吃肉，說：『我要吃肉』，就可以隨心所欲吃肉。
DEUT|12|21|耶和華－你上帝選擇立他名的地方若離你太遠，你可以照我所吩咐的，將耶和華賜給你的牛羊取些宰了，隨心所欲在你的城裏吃。
DEUT|12|22|其實，就如吃羚羊和鹿的肉一樣，你要這樣吃它，無論潔淨的人不潔淨的人都可以一起吃。
DEUT|12|23|但是你要堅定，不可吃血，因為血是生命；不可將生命與肉一起吃。
DEUT|12|24|你不可吃血，要把它倒在地上，如同倒水一樣。
DEUT|12|25|不可吃血，好讓你和你的子孫可以得福，因為你行了耶和華眼中看為正的事。
DEUT|12|26|只是你分別為聖的物和你所還的願，都要帶到耶和華所選擇的地方去。
DEUT|12|27|你的燔祭，連肉帶血，都要獻在耶和華－你上帝的壇上。祭物的血要倒在耶和華－你上帝的壇上；肉你可以吃。
DEUT|12|28|你要謹守聽從我所吩咐的一切話，好讓你和你的子孫可以永遠得福，因為你行耶和華－你上帝眼中看為善、看為正的事。」
DEUT|12|29|「耶和華－你上帝把你要進去趕出的列國從你面前剪除，並且你得了他們的地為業居住，
DEUT|12|30|那時你要謹慎，在他們從你面前被除滅之後，你不可受引誘隨從他們，也不可求問他們的神明，說：『這些國家怎樣事奉他們的神明，我也要照樣做。』
DEUT|12|31|你不可向耶和華－你的上帝這樣做，因為他們向他們的神明做了耶和華所憎恨、所厭惡的一切事，甚至將自己的兒女用火焚燒，獻給他們的神明。
DEUT|12|32|凡我所吩咐你們的事，你們都要謹守遵行，不可加添，也不可刪減。」
DEUT|13|1|「你中間若有先知或是做夢的人起來，向你顯神蹟奇事，
DEUT|13|2|他對你說的神蹟奇事應驗了，說：『我們去隨從別神，事奉它們吧。』那是你不認識的。
DEUT|13|3|你不可聽那先知或是那做夢之人的話，因為這是耶和華－你們的上帝考驗你們，要知道你們是否盡心盡性愛耶和華－你們的上帝。
DEUT|13|4|你們要順從耶和華－你們的上帝，敬畏他，謹守他的誡命，聽從他的話，事奉他，緊緊跟隨他。
DEUT|13|5|那先知或那做夢的人要被處死，因為他出言悖逆那領你們出 埃及 地、救贖你脫離為奴之家的耶和華－你們的上帝，要引誘你離開耶和華－你上帝吩咐你要行的道。這樣，你就把惡從你中間除掉。
DEUT|13|6|「你的同胞兄弟，或是你的兒女，或是你懷中的妻，或是如同自己性命的朋友，若暗中引誘你，說：『我們去事奉別神吧。』那是你和你列祖所不認識的，
DEUT|13|7|你四圍列國的神明，無論是離你近或離你遠，從地這邊到地那邊，
DEUT|13|8|你都不可附和他，也不要聽從他。你的眼不可顧惜他，不可憐憫他，也不可袒護他。
DEUT|13|9|你務必殺他；你先下手，然後眾百姓才下手，把他處死。
DEUT|13|10|要用石頭打死他，因為他想引誘你離開那領你出 埃及 地為奴之家的耶和華－你的上帝。
DEUT|13|11|全 以色列 都要聽見而害怕，不敢在你中間再行這樣的惡事了。
DEUT|13|12|「若你聽見人說，在耶和華－你上帝所賜給你居住的城鎮中的一座，
DEUT|13|13|有些無賴之徒從你中間出來，引誘本城的居民，說：『我們去事奉別神吧。』那是你們不認識的，
DEUT|13|14|你就要調查，探聽，細心詢問。看哪，是真的，確實有這可憎的事在你中間發生，
DEUT|13|15|你務必用刀殺那城裏的居民，把城裏所有的，連牲畜都用刀滅盡。
DEUT|13|16|你要把從城裏所奪取的一切財物堆在廣場中，用火將那城和其中奪取的一切財物全燒給耶和華－你的上帝。那城要永遠成為廢墟，不得重建。
DEUT|13|17|那當毀滅的物一點都不可黏你的手，好讓耶和華轉回，不向你發烈怒，卻恩待你，憐憫你，照他向你列祖所起的誓使你人數增多；
DEUT|13|18|因為你聽從耶和華－你上帝的話，遵守我今日所吩咐你的一切誡命，行耶和華－你上帝眼中看為正的事。」
DEUT|14|1|「你們是耶和華─你們上帝的兒女。不可為了死人割劃自己，也不可使額上 光禿；
DEUT|14|2|因為你是屬於耶和華－你上帝神聖的子民，耶和華從地面上的萬民中揀選了你，作自己寶貴的子民。」
DEUT|14|3|「凡可憎的物， 你都不可吃。
DEUT|14|4|可吃的牲畜是：牛、綿羊、山羊、
DEUT|14|5|鹿、羚、麃子、野山羊、瞪羚、羚羊、山綿羊。
DEUT|14|6|凡蹄分兩瓣，分趾蹄而又反芻食物的牲畜，你們都可以吃。
DEUT|14|7|但那反芻或分蹄之中不可吃的是：駱駝、兔子、石獾，雖然反芻卻不分蹄，對你們是不潔淨的；
DEUT|14|8|豬，雖然分蹄卻不反芻，對你們也是不潔淨的。牠們的肉，你們一點都不可吃；牠們的屍體，你們也不可摸。
DEUT|14|9|「水中可吃的是這些：凡有鰭有鱗的都可以吃；
DEUT|14|10|凡無鰭無鱗的都不可吃，對你們是不潔淨的。
DEUT|14|11|「凡潔淨的鳥，你們都可以吃。
DEUT|14|12|不可吃的是：鵰、狗頭鵰、紅頭鵰、
DEUT|14|13|鸇、小鷹、鷂鷹的類群，
DEUT|14|14|各種烏鴉的類群、
DEUT|14|15|鴕鳥、夜鷹、魚鷹、鷹的類群、
DEUT|14|16|鴞鳥、貓頭鷹、角鴟、
DEUT|14|17|鵜鶘、禿鵰、鸕鶿、
DEUT|14|18|鸛、鷺鷥的類群、戴鵀與蝙蝠。
DEUT|14|19|凡有翅膀卻爬行的群聚動物對你們是不潔淨的，都不可吃。
DEUT|14|20|凡潔淨的鳥，你們都可以吃。
DEUT|14|21|「凡自然死去的動物，你們都不可吃，可以給城裏寄居的人吃，或賣給外人，因為你是屬於耶和華－你上帝神聖的子民。 「不可用母山羊的奶來煮牠的小山羊。」
DEUT|14|22|「每年，你務必從你播種的一切收成，田地所出產的，取十分之一獻上。
DEUT|14|23|要在耶和華－你上帝面前，就是他選擇那裏作為他名居所的地方，吃你所獻十分之一的五穀、新酒和新的油，以及牛群羊群中頭生的，好讓你天天學習敬畏耶和華－你的上帝。
DEUT|14|24|當耶和華－你的上帝賜福給你的時候，耶和華－你上帝選擇立他名的地方若離你太遠，路途太長，使你不能把這東西帶到那裏去，
DEUT|14|25|你可以把它換成銀子，把銀子包起來，拿在手中，往耶和華－你上帝所選擇的地方去。
DEUT|14|26|在那裏，你可以隨心所欲用銀子或買牛羊，或買清酒烈酒，或買任何你心所想的。你和你的全家要在耶和華－你上帝面前吃喝歡樂。
DEUT|14|27|「住在你城裏的 利未 人，你不可離棄他，因為他在你那裏沒有分得產業。
DEUT|14|28|每三年的最後一年，你要把那一年收成的十分之一取出來，積存在你的城中；
DEUT|14|29|那沒有與你一起分得產業的 利未 人，和城裏的寄居者，以及孤兒寡婦，都可以前來，吃得飽足，好讓耶和華－你的上帝在你手裏所做的一切事上賜福給你。」
DEUT|15|1|「每七年的最後一年，你要施行豁免。
DEUT|15|2|豁免的方式是這樣：凡債主要把手裏所借給鄰舍的全豁免，不可向鄰舍和弟兄追討，因為耶和華的豁免已經宣告了。
DEUT|15|3|你可以向外邦人追討；但你弟兄欠你的，無論是甚麼，你都要放手豁免。
DEUT|15|4|其實，在你中間不會有貧窮人；因為在耶和華－你上帝所賜你為業的地上，耶和華必大大賜福給你。
DEUT|15|5|只要你留心聽從耶和華－你上帝的話，謹守遵行我今日所吩咐你這一切的命令，
DEUT|15|6|因為耶和華－你的上帝會照他所應許你的賜福給你，你必借給許多國家，卻不需要去借貸；你要管轄許多國家，它們卻不能管轄你。
DEUT|15|7|「在耶和華－你上帝所賜給你的地上，任何一座城裏，你弟兄中若有一個貧窮人，你不可硬著心，袖手不幫助你貧窮的弟兄。
DEUT|15|8|你總要伸手幫助他，照他所缺乏的借給他，補他的不足。
DEUT|15|9|你要謹慎，不可心起惡念，說：『第七年的豁免年快到了』，你就冷眼看你貧窮的弟兄，甚麼都不給他。他若為你的緣故求告耶和華，你就有罪了。
DEUT|15|10|你要慷慨解囊，給他的時候不要心疼，因為耶和華－你的上帝必為這事，在你一切的工作上和你手所做的一切賜福給你。
DEUT|15|11|因為地上的貧窮人永遠不會斷絕，所以我吩咐你說：『總要伸手幫助你地上困苦貧窮的弟兄。』」
DEUT|15|12|「你弟兄中，若有一個 希伯來 男人或 希伯來 女人賣給你，已服事你六年，到了第七年就要讓他自由離開你。
DEUT|15|13|你讓他自由離開的時候，不可讓他空手而去，
DEUT|15|14|要從你的羊群、禾場、壓酒池中取一些，慷慨地送給他；耶和華－你的上帝怎樣賜福給你，你也要照樣給他。
DEUT|15|15|要記得你在 埃及 地作過奴僕，耶和華－你的上帝救贖了你。為此，我今日將這事吩咐你。
DEUT|15|16|他若對你說：『我不願意離開你』，因為他愛你和你的家，並且他在你那裏很好，
DEUT|15|17|你要拿錐子在門上穿透他的耳朵，他就永遠成為你的奴僕了。你待婢女也要這樣。
DEUT|15|18|你讓他從你那裏自由離開的時候，不要看作困難，因為他已服事你六年，相當於雇工雙倍的工錢。這樣，耶和華－你的上帝必在你所做的一切事上賜福給你。」
DEUT|15|19|「你牛群羊群中頭生的，凡是公的，都要分別為聖，歸給耶和華－你的上帝。頭生的牛，不可用牠來耕作；頭生的羊，不可剪牠的毛。
DEUT|15|20|這頭生的，你和你全家每年要到耶和華所選擇的地方，在耶和華－你上帝面前吃。
DEUT|15|21|這頭生的若有殘疾，瘸腿的或瞎眼的，若有任何嚴重缺陷，都不可獻給耶和華－你的上帝。
DEUT|15|22|你們可以在城裏吃，潔淨的人和不潔淨的人都可以吃，就如吃羚羊和鹿一樣。
DEUT|15|23|只是牠的血，你不可吃，要倒在地上，如同倒水一樣。」
DEUT|16|1|「你要守亞筆月，向耶和華－你的上帝守逾越節，因為在亞筆月，耶和華－你的上帝在夜間領你出 埃及 。
DEUT|16|2|你當在那裏，耶和華選擇作為他名居所的地方，從羊群牛群中，將逾越節的祭牲獻給耶和華－你的上帝。
DEUT|16|3|這祭牲不可和有酵的東西一起吃。因為你曾匆忙離開 埃及 地，你要吃無酵餅，就是困苦餅七日，好讓你一生的年日記得你從 埃及 地出來的那一日。
DEUT|16|4|在你全境內，七日不可見到酵母。第一日晚上所獻的肉，一點也不可留到早晨。
DEUT|16|5|你不可在耶和華－你上帝所賜的各城中，任何一座城裏，獻逾越節的祭，
DEUT|16|6|只可在那裏，耶和華－你上帝選擇作為他名居所的地方，在晚上日落的時候，就是你出 埃及 的時候，獻逾越節的祭。
DEUT|16|7|你要在耶和華－你上帝所選擇的地方把肉烤來吃，次日早晨就回到你的帳棚去。
DEUT|16|8|你要吃無酵餅六日，第七日要向耶和華－你的上帝守嚴肅會，不可做工。」
DEUT|16|9|「你要計算七個七日：從你用鐮刀開始收割莊稼時算起，一共七個七日。
DEUT|16|10|你要向耶和華－你的上帝守七七節，按照耶和華－你上帝所賜你的福，獻上你手裏的甘心祭。
DEUT|16|11|你和你的兒女、僕婢，以及住在你城裏的 利未 人、在你中間寄居的和孤兒寡婦，都要在那裏，耶和華－你上帝選擇作為他名居所的地方，在耶和華－你上帝面前歡樂。
DEUT|16|12|你要記得你在 埃及 作過奴僕，也要謹守遵行這些律例。」
DEUT|16|13|「你收藏了禾場和壓酒池的出產以後，就要守住棚節七日。
DEUT|16|14|在節期中，你和你的兒女、僕婢，以及住在你城裏的 利未 人、寄居的和孤兒寡婦，都要歡樂。
DEUT|16|15|在耶和華所選擇的地方，你要向耶和華－你的上帝守節七日，因為耶和華－你的上帝要在你一切的收成上和你手裏所做的一切賜福給你，你就非常歡樂。
DEUT|16|16|「你所有的男丁要在除酵節、七七節、住棚節，一年三次，在耶和華－你上帝所選擇的地方朝見他，不可空手朝見耶和華。
DEUT|16|17|各人要按自己手中的能力，照耶和華－你上帝所賜你的福，奉獻禮物。」
DEUT|16|18|「你要在耶和華－你上帝所賜的各城中，為各支派設立審判官和官長。他們要按公義的判斷審判百姓，
DEUT|16|19|不可屈枉正直，不可看人的情面，也不可接受賄賂，因為賄賂能使智慧人的眼睛變瞎，又能曲解義人的證詞。
DEUT|16|20|公正！你要追求公正，好使你存活，承受耶和華－你上帝所賜你的地。」
DEUT|16|21|「你為耶和華－你的上帝築壇，不可在壇旁栽種任何樹木作 亞舍拉 ，
DEUT|16|22|也不可為自己設立柱像，這是耶和華－你的上帝所憎恨的。」
DEUT|17|1|「凡有殘疾，有任何惡疾的牛羊，你都不可獻給耶和華－你的上帝，因為這是耶和華－你上帝所憎惡的。
DEUT|17|2|「在你中間，在耶和華－你上帝所賜你的各城中，任何一座城裏，若有男人或女人做了耶和華－你上帝眼中看為惡的事，違背了他的約，
DEUT|17|3|去事奉別神，敬拜它們，或拜太陽，或拜月亮，或拜天上的萬象，是我 不曾吩咐的。
DEUT|17|4|有人告訴你，你也聽見了，就要細心探聽。看哪，是真的，確實有這可憎的事在 以色列 中發生，
DEUT|17|5|你就要將行這惡事的男人或女人拉到城門外，用石頭把這男人或女人處死。
DEUT|17|6|要憑兩個證人或三個證人的口，才可以把他處死，不可只憑一個證人的口處死他。
DEUT|17|7|證人要先動手，然後眾百姓也動手把他處死。這樣，你就把惡從你中間除掉。
DEUT|17|8|「你城中若有難以判斷的案件，涉及流血，訴訟，或毆打等爭訟的事，你就要起來，上到那裏，耶和華－你上帝所選擇的地方，
DEUT|17|9|去見 利未 家的祭司和當時的審判官，求問他們，他們必將判決指示你。
DEUT|17|10|他們在耶和華所選擇的地方指示你的判決，你要執行，謹守遵行他們一切所教導你的。
DEUT|17|11|要按照所教導你的律法、所告訴你的典章去執行；他們指示你的判決，你不可偏離左右。
DEUT|17|12|若有人擅自行事，不聽從那侍立在耶和華－你上帝那裏事奉的祭司，或不聽從審判官，那人就要處死。這樣，你就把惡從 以色列 中除掉。
DEUT|17|13|眾百姓聽見了都要害怕，不再擅自行事了。」
DEUT|17|14|「你到了耶和華－你上帝所賜你的地，得了那地居住在其中的時候，若說：『我要立王治理我，像我四圍所有的國家一樣』，
DEUT|17|15|你一定要立耶和華－你上帝所揀選的人為你的王。要從你弟兄中立一人為你的王，不可立你弟兄之外的外邦人治理你。
DEUT|17|16|只是王不可為自己加添馬匹，也不可為加添馬匹使百姓回 埃及 去，因耶和華曾對你們說：『不可再回那條路去。』
DEUT|17|17|王不可為自己多立妃嬪，免得他的心偏離；也不可為自己多積金銀。
DEUT|17|18|他登了國度的王位之後，要在 利未 家的祭司面前，將這律法書為自己抄寫一份在書卷上。
DEUT|17|19|這書要存在他那裏，他一生的年日要誦讀，好使他學習敬畏耶和華－他的上帝，謹守遵行這律法書上的一切話和這些律例，
DEUT|17|20|免得他的心向弟兄高傲，偏離了這誡命，或向右或向左。這樣，他和他的子孫就可以長久作王治理 以色列 。」
DEUT|18|1|「 利未 家的祭司和 利未 全支派在 以色列 中沒有分得產業；他們可以吃耶和華的火祭，那是他的產業。
DEUT|18|2|他在弟兄中沒有產業；耶和華是他的產業，正如耶和華所應許他的。
DEUT|18|3|祭司從百姓當得的權益是這樣：凡獻牛或羊為祭物的，要把前腿、兩腮和胃給祭司。
DEUT|18|4|初收的五穀、新酒和新的油，以及初剪的羊毛，也要給他。
DEUT|18|5|因為耶和華－你的上帝從你眾支派中揀選他，使他和他子孫永遠奉耶和華的名侍立，事奉。
DEUT|18|6|「 利未 人若離開他在 以色列 中所居住的任何一座城，一心願意到耶和華所選擇的地方，
DEUT|18|7|就要在那裏奉耶和華－他上帝的名事奉，正如他的眾弟兄 利未 人在耶和華面前侍立一樣。
DEUT|18|8|除了賣祖產所得的以外，他們 要吃同等分量的祭物。」
DEUT|18|9|「你到了耶和華－你上帝所賜你之地，不可學那些國家行可憎惡的事。
DEUT|18|10|你中間不可有人使兒女經火，也不可有占卜的、觀星象的、行法術的 、行邪術的、
DEUT|18|11|施符咒的、招魂的、行巫術的和求問死人的。
DEUT|18|12|凡做這些事的都是耶和華所憎惡的；因這可憎惡的事，耶和華－你的上帝把他們從你面前趕出去。
DEUT|18|13|你要向耶和華－你的上帝作完全人。
DEUT|18|14|你所要趕出的那些國家都聽從觀星象的和占卜的，但是耶和華－你的上帝從來不准你這樣做。」
DEUT|18|15|「耶和華－你的上帝要從你弟兄中給你興起一位先知像我，你們要聽他。
DEUT|18|16|這正如你在 何烈山 大會的那日向耶和華－你的上帝所求的一切，說：『求你不要再叫我聽見耶和華－我上帝的聲音，也不要再叫我看見這大火，免得我死亡。』
DEUT|18|17|耶和華對我說：『他們說得對。
DEUT|18|18|我必在他們弟兄中給他們興起一位先知像你。我要將當說的話放在他口裏；他要將我一切所吩咐的都告訴他們。
DEUT|18|19|誰不聽從他奉我名所說的話，我必親自向他追究。
DEUT|18|20|若有先知擅自奉我的名說了我未曾吩咐他說的話，或是奉別神的名說話，那先知就必處死。』
DEUT|18|21|你心裏若說：『我們怎能知道那話是耶和華未曾吩咐的呢？』
DEUT|18|22|先知奉耶和華的名說話，所說的若沒有實現，或不應驗，這話就是耶和華未曾吩咐的，而是那先知擅自說的，你不必怕他。」
DEUT|19|1|「耶和華－你的上帝將列國剪除，他們的地耶和華－你上帝已賜給你，你又趕出他們，並且住在他們的城鎮和房屋，
DEUT|19|2|那時，你要在耶和華－你上帝所賜你為業的地上，為自己指定三座城。
DEUT|19|3|你要預備道路，將耶和華－你上帝使你承受為業的地分為三區，使任何一個殺人的可以逃到那裏去。
DEUT|19|4|「殺人的逃到那裏得以存活的案例是這樣：凡素無仇恨，無意中殺了鄰舍的，
DEUT|19|5|就如人與鄰舍同入林中伐木，手拿斧子一砍，本想砍下樹木，斧頭卻脫了把，飛落在鄰舍身上，以致那人死去，這人就可以逃到那些城中的一座，得以存活，
DEUT|19|6|免得報血仇的心中發火，去追趕那殺了人的，因為路途遙遠就能追上他，把他殺死。其實他是不該死的，因為他與被殺者素無仇恨。
DEUT|19|7|所以我吩咐你說，要為自己指定三座城。
DEUT|19|8|耶和華－你的上帝若照他向你列祖所起的誓擴張你的疆土，將所應許賜你列祖的全地給你，
DEUT|19|9|你若謹守遵行我今日所吩咐的這一切誡命，愛耶和華－你的上帝，天天遵行他的道，就要在這三座城之外，再添三座城，
DEUT|19|10|免得無辜人的血流在耶和華－你上帝所賜你為業的地中間，血就歸到你身上了。
DEUT|19|11|「若有人恨他的鄰舍，埋伏等著，起來擊殺他，把他殺死，然後逃到這些城中的一座，
DEUT|19|12|他本城的長老就要派人去，從那裏把他帶出來，交在報血仇者的手中，把他處死。
DEUT|19|13|你的眼不可顧惜他，要從 以色列 中除掉流無辜血的罪，使你得福。」
DEUT|19|14|「在耶和華－你上帝所賜你承受為業，所分得的地上，不可挪移你鄰舍的地界，因為這是前人所定的。」
DEUT|19|15|「人無論犯甚麼罪，作甚麼惡，不可單憑一個人的見證，總要憑兩個證人的口或三個證人的口才可定案。
DEUT|19|16|若有人懷惡意，起來作證，控告他人犯法，
DEUT|19|17|這兩個爭訟的人就要站在耶和華面前，和當時的祭司與審判官面前，
DEUT|19|18|審判官要細心調查。看哪，證人作的是偽證，要用偽證陷害弟兄，
DEUT|19|19|你們就要對付他如同他想要對付的弟兄一樣。這樣，你就把惡從你中間除掉。
DEUT|19|20|其他的人聽見就害怕，不敢在你中間再行這樣的惡事了。
DEUT|19|21|你的眼不可顧惜，要以命償命，以眼還眼，以牙還牙，以手還手，以腳還腳。」
DEUT|20|1|「你出去與仇敵作戰，若看見馬匹、戰車，以及比你更多的士兵，不要怕他們，因為領你出 埃及 地的耶和華－你的上帝與你同在。
DEUT|20|2|你們將要上陣的時候，祭司要來，向士兵宣告，
DEUT|20|3|對他們說：『 以色列 啊，要聽！你們今日將要與仇敵作戰，不要心驚膽戰，不要懼怕戰兢，也不要因他們驚慌，
DEUT|20|4|因為與你們同去的是耶和華－你們的上帝，他要為你們與仇敵作戰，拯救你們。』
DEUT|20|5|官長也要向士兵宣告說：『誰建了新的房屋尚未奉獻，他可以回家去，免得他陣亡，別人去奉獻。
DEUT|20|6|誰栽植了葡萄園尚未享用所結的果子，他可以回家去，免得他陣亡，別人去享用。
DEUT|20|7|誰與女子訂了婚尚未迎娶，他可以回家去，免得他陣亡，別人去娶。』
DEUT|20|8|官長要繼續對士兵說：『誰懼怕，心驚膽戰，可以回家去，免得他弟兄的心像他的心一樣消沉。』
DEUT|20|9|官長向士兵宣告完畢，軍官就率領士兵去了。
DEUT|20|10|「你來到一座城，要攻城之前，先向它宣告和平。
DEUT|20|11|那城若願意以和平回應，給你開城，城裏所有的人就要為你做苦工，服事你。
DEUT|20|12|若那城拒絕和平，卻要與你打仗，你就要圍困那城。
DEUT|20|13|耶和華－你的上帝把那城交在你手裏時，你就要用刀殺盡城裏的男丁。
DEUT|20|14|至於婦女、孩童、牲畜和城裏所有的，你都可以取為自己的掠物。從仇敵所掠奪的，就是耶和華－你上帝所賜給你的，你都可以享用。
DEUT|20|15|離你很遠的各城，就是不屬於這些國家的城鎮，你都要這樣對待他們。
DEUT|20|16|但是這些民族的城鎮，就是耶和華－你上帝所賜給你的產業，其中凡有氣息的，一個都不可存留。
DEUT|20|17|你要照耶和華－你上帝所吩咐的，將這些 赫 人、 亞摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人全都滅絕，
DEUT|20|18|免得他們教導你們去行一切可憎惡的事，就是他們向自己神明所行的，使你們得罪耶和華－你們的上帝。
DEUT|20|19|「你若圍困一座城，需要攻打許多日子才能奪取，就不可用斧頭砍壞樹木。你可以吃樹上的果子，卻不可把樹砍下來。田間的樹木豈是人，讓你去圍攻的嗎？
DEUT|20|20|只有那些你知道不能生產食物的樹才可以毀壞；你可以把它們砍下來造攻城的工具，攻打那與你打仗的城，直到把城攻下。」
DEUT|21|1|「在耶和華－你上帝所賜你為業的地上，若發現有人被殺，暴屍野地，不知道是誰殺的，
DEUT|21|2|長老和審判官 就要出去，從屍體那裏量起，量到四圍的城鎮，
DEUT|21|3|看哪一座城最靠近這屍體，那城的幾位長老就要取一頭未曾耕地、未曾負軛的母牛犢；
DEUT|21|4|那城的長老要把這母牛犢牽到流著溪水、未曾耕耘、未曾撒種的山谷去，在谷中打斷牠的頸項。
DEUT|21|5|利未 人祭司要近前來，因為耶和華－你的上帝揀選他們來事奉他，奉耶和華的名祝福，並且有任何的爭訟和毆打，都由他們的口判決。
DEUT|21|6|離屍體最近的那座城的每位長老要在山谷中，在頸項被打斷的母牛犢上面洗手，
DEUT|21|7|聲明說：『我們的手未曾流這人的血；我們的眼也未曾看見這事。
DEUT|21|8|耶和華啊，求你赦免你所救贖的百姓 以色列 ，不要讓無辜的血歸在你的百姓 以色列 中間。』這樣，他們流血的罪就必得赦免。
DEUT|21|9|你行了耶和華眼中看為正的事，就可以從你中間除掉無辜的血。」
DEUT|21|10|「你出去與仇敵作戰的時候，耶和華－你的上帝將他交在你手中，你就擄了他為俘虜。
DEUT|21|11|若你在被擄的人中看見美麗的女子，喜歡她，要娶她為妻，
DEUT|21|12|就可以帶她到你家去。她要剪頭髮，修指甲，
DEUT|21|13|脫去被擄時所穿的衣服，住在你家裏為自己父母哀哭一個月。然後，你就可以與她同房；你作她的丈夫，她作你的妻子。
DEUT|21|14|以後你若不喜歡她，就要讓她自由離開，絕不可為錢把她賣了，也不可把她當奴隸看待，因為你已經佔有過她。」
DEUT|21|15|「人若有兩個妻子，一個是他寵愛的，另一個是失寵的 ，她們都給他生了兒子，但長子是他失寵妻子生的；
DEUT|21|16|到了分產業給兒子的時候，不可將自己寵愛的妻子所生的兒子立為長子，在他失寵妻子所生的長子之上。
DEUT|21|17|他必須認失寵妻子所生的兒子為長子，在所有的產業中給他雙分，因為這兒子是他壯年時生的，長子的名分應當是他的。」
DEUT|21|18|「人若有頑梗忤逆的兒子，不聽從父母的話，他們雖然懲戒他，他還是不聽從他們，
DEUT|21|19|父母就要抓住他，帶他出去到當地的城門，本城的長老那裏，
DEUT|21|20|對本城的長老說：『我們這個兒子頑梗忤逆，不聽從我們的話，是貪食好酒的人。』
DEUT|21|21|然後，城裏的眾人就要用石頭將他打死。這樣，你就把惡從你中間除掉，全 以色列 聽見了都要害怕。」
DEUT|21|22|「人若犯了死罪被處死，你把他掛在木頭上，
DEUT|21|23|不可讓屍體留在木頭上過夜，一定要當日把他埋葬，因為被掛的人是上帝所詛咒的。你不可玷污耶和華－你上帝所賜你為業的地。」
DEUT|22|1|「你若看見弟兄的牛或羊迷了路，不可避開牠們，總要把牠們牽回來交給你的弟兄。
DEUT|22|2|你弟兄若離你遠，或是你不認識他，你就要牽到你家，留在你那裏，等你的弟兄來尋找就還給他。
DEUT|22|3|你弟兄所失落的，無論是驢，衣服，或任何東西，你若發現，都要這樣做，不能避開。
DEUT|22|4|你若看見你弟兄的牛或驢在路上跌倒了，不可避開牠們，總要幫助他把牛或驢拉起來。
DEUT|22|5|「婦女不可穿戴男子所穿戴的，男人也不可穿婦女的衣服，因為這樣做是耶和華－你上帝所憎惡的。
DEUT|22|6|「你若路上看見鳥窩，無論在樹上或地上，裏頭有小鳥或有蛋，母鳥伏在小鳥或蛋上，你不可連母鳥帶小鳥一起拿去。
DEUT|22|7|總要放母鳥走，只可以取小鳥。這樣你就可以享福，日子得以長久。
DEUT|22|8|「你若建造新房屋，要在屋頂安欄杆，免得有人從屋頂掉下來，血就歸於你家。
DEUT|22|9|「不可在你的葡萄園裏栽種別的種子，免得你栽種所結的和葡萄園的果子都成了聖物。
DEUT|22|10|不可並用牛和驢來耕地。
DEUT|22|11|不可穿羊毛和細麻混合做成的衣服。
DEUT|22|12|「你要在所披外衣的四個邊上縫繸子。」
DEUT|22|13|「人若娶妻，與她同房後恨惡她，
DEUT|22|14|捏造她行可恥的事，把醜名加在她身上，說：『我娶了這女人，親近她，卻發現她沒有貞潔的憑據』。
DEUT|22|15|女方的父母就要把這女子貞潔的憑據拿出去，到城門的本城長老那裏。
DEUT|22|16|女方的父親要對長老說：『我把女兒嫁給這人，他卻恨惡她，
DEUT|22|17|看哪，他捏造可恥的事，說：我發現你女兒沒有貞潔的憑據。但是，這就是我女兒貞潔的憑據。』父母要把那布鋪在本城長老的面前。
DEUT|22|18|那城的長老要拿住那人，懲罰他，
DEUT|22|19|罰他一百銀子，給女方的父親，因為他把醜名加在 以色列 一個少女身上。這女子仍是他的妻子，那人終身不可休她。
DEUT|22|20|但若這事是真的，找不到女子貞潔的憑據，
DEUT|22|21|他們就要把這女子帶到她父家的門口，城裏的人要用石頭打死她，因為她在父家犯了淫亂，在 以色列 中做了可恥的事。這樣，你就把惡從你中間除掉。
DEUT|22|22|「若發現有人與有夫之婦同寢，就要將姦夫淫婦一起處死。這樣，你就把惡從 以色列 中除掉。
DEUT|22|23|「若一女子是處女，已經許配了人，有男子在城裏遇見她，與她同寢，
DEUT|22|24|你們就要把這二人帶到那城的城門口，用石頭打死他們。處死女子是因為她雖然在城裏， 卻沒有喊叫；處死男子是因為他玷污了鄰舍的妻子。這樣，你就把惡從你中間除掉。
DEUT|22|25|「若有男子在野地遇見已經許配人的女子，抓住她與她同寢，只要處死那與女子同寢的男子。
DEUT|22|26|不可對女子處刑，這女子沒有該死的罪。這案件就好比人起來攻擊鄰舍，把他殺了一樣。
DEUT|22|27|因為男子是在野地遇見她，這已經許配了人的女子雖然喊叫，卻沒有人救她。
DEUT|22|28|「若有男子遇見沒有許配人的少女，抓住她與她同寢，被人發現，
DEUT|22|29|這男子就要拿五十銀子給女子的父親，並要娶她為妻，終身不可休她，因為他玷污了這女子。
DEUT|22|30|「人不可娶繼母為妻，不可掀開父親衣服的下邊 。」
DEUT|23|1|「凡外腎損傷的，或被閹割的，不可入耶和華的會。
DEUT|23|2|「私生子不可入耶和華的會；甚至到第十代，也不可入耶和華的會。
DEUT|23|3|「 亞捫 人或 摩押 人不可入耶和華的會；甚至到第十代，也永不可入耶和華的會。
DEUT|23|4|因為你們出 埃及 的時候，他們沒有拿食物和水在路上迎接你們，並且雇了 美索不達米亞 的 毗奪 人， 比珥 的兒子 巴蘭 來詛咒你。
DEUT|23|5|然而耶和華－你的上帝不願聽 巴蘭 ，耶和華－你的上帝為你使詛咒變為祝福，因為耶和華－你的上帝愛你。
DEUT|23|6|你一生一世永不可為他們求平安和福氣。
DEUT|23|7|「不可憎惡 以東 人，因為他是你的弟兄。不可憎惡 埃及 人，因為你曾在他的地上作過寄居的。
DEUT|23|8|他們所生的第三代子孫可以入耶和華的會。」
DEUT|23|9|「你出兵攻打敵人，要遠離一切惡事。
DEUT|23|10|「你中間若有人因夜間夢遺而不潔淨，就要出到營外，不可入營。
DEUT|23|11|到了傍晚，他要用水洗澡，等到日落才可以入營。
DEUT|23|12|「你要在營外劃定一個地方，你可以出去在那裏方便。
DEUT|23|13|在你器械中當有一把鍬；你出營外便溺以後，要用它挖洞，轉身掩蓋排泄物。
DEUT|23|14|因為耶和華－你的上帝在你營中走動，要拯救你，將仇敵交給你，所以你的營應當聖潔，免得他見你那裏有污穢之物就轉身離開你。」
DEUT|23|15|「你不可把從主人身邊逃到你那裏的奴僕，交回給他的主人，
DEUT|23|16|要讓他在你那裏與你同住，由他在你的城鎮中選擇一個自己喜歡的地方居住，不可欺負他。
DEUT|23|17|「 以色列 的女子中不可作神廟娼妓； 以色列 的男子中也不可作神廟娼妓。
DEUT|23|18|妓女和男娼 的賞金，都不可帶進耶和華－你上帝的殿中還願，因為兩者都是耶和華－你上帝所憎惡的。
DEUT|23|19|「你借給你弟兄的，無論是錢財是糧食，或任何可生利息的財物，都不可取利。
DEUT|23|20|借給外邦人可以取利，但借給你的弟兄就不可取利；好讓耶和華－你的上帝在你去得為業的地上和你手裏所做的一切，賜福給你。
DEUT|23|21|「你向耶和華－你的上帝許願，不可遲延還願，因為耶和華－你的上帝必定向你追討，你就有罪了。
DEUT|23|22|你若不許願，倒沒有罪。
DEUT|23|23|你嘴唇所說的，你親口承諾的，要照你甘心向耶和華－你上帝許的願謹守遵行。
DEUT|23|24|「你進入鄰舍的葡萄園，可以隨意吃葡萄，直到飽足，卻不可裝在器皿中。
DEUT|23|25|你進入鄰舍的莊稼中，可以用手摘麥穗，卻不可用鐮刀割取莊稼。」
DEUT|24|1|「人若娶妻，作了她的丈夫，發現她有不合宜的事不喜歡她，而寫休書交在她手中，打發她離開夫家，
DEUT|24|2|婦人若離開夫家以後，去嫁別人，
DEUT|24|3|後夫若恨惡她，寫休書交在她手中，打發她離開夫家，又或者娶她為妻的後夫死了，
DEUT|24|4|那休她的前夫就不可在婦人玷污之後再娶她為妻，因為這是耶和華所憎惡的。不可使耶和華－你上帝所賜為業之地蒙受玷污。
DEUT|24|5|「人若娶了新娘，不可從軍出征，也不可派他辦理任何事情。他可以在家清閒一年，使他所娶的妻快活。
DEUT|24|6|「不可拿人的石磨或上面的磨石作抵押，因為這是拿人的命作抵押。
DEUT|24|7|「若發現有人綁架 以色列 人中的一個弟兄，把他當奴隸對待，或把他賣了，那綁架人的就必處死。這樣，你就把惡從你中間除掉。
DEUT|24|8|「關於痲瘋 的災病，你們要謹慎，照 利未 家的祭司一切所指教你們的留心遵行。我怎樣吩咐他們，你們要照樣遵行。
DEUT|24|9|要記得，在你們出 埃及 後的路途中，耶和華－你的上帝向 米利暗 所做的事。
DEUT|24|10|「你借給鄰舍，無論是甚麼，不可進他家拿抵押品。
DEUT|24|11|要站在外面，等那借貸的人把抵押品拿出來交給你。
DEUT|24|12|他若是困苦的人，你不可用他的抵押品蓋著睡覺。
DEUT|24|13|日落的時候，總要把抵押品還給他，讓他用那件外衣蓋著睡覺，他就為你祝福。這在耶和華－你的上帝面前就是你的義行了。
DEUT|24|14|「困苦貧窮的雇工，無論是你的弟兄，或是住在你境內，在你城裏寄居的，你都不可欺負他 。
DEUT|24|15|要當日給他工錢，不可等到日落，因為他困苦，需要靠工錢過活，免得他因你的緣故求告耶和華，罪就歸於你了。
DEUT|24|16|「不可因兒子處死父親，也不可因父親處死兒子；各人要因自己的罪被處死。
DEUT|24|17|「不可對寄居的和孤兒屈枉正直，也不可拿寡婦的衣服作抵押。
DEUT|24|18|要記得你曾在 埃及 作過奴僕，耶和華－你的上帝從那裏救贖了你，所以我吩咐你遵行這事。
DEUT|24|19|「你在田間收割莊稼，若忘了一捆在田間，就不要再回去拿，要留給寄居的、孤兒和寡婦；好讓耶和華－你的上帝在你手裏所做的一切，賜福給你。
DEUT|24|20|你打了橄欖樹，枝上剩下的不可再打，要留給寄居的、孤兒和寡婦。
DEUT|24|21|你摘葡萄園的葡萄，掉落的不可拾取，要留給寄居的、孤兒和寡婦。
DEUT|24|22|你要記得你曾在 埃及 地作過奴僕，所以我吩咐你遵行這事。
DEUT|25|1|「人與人若有爭訟，要求審判，當宣判義人為義，惡人有罪的時候，
DEUT|25|2|惡人若該受責打，審判官就要叫他當著面，伏在地上，按他的罪照數責打。
DEUT|25|3|只能打四十下，不可加多；多過這數目就是在你眼中作賤你的弟兄了。
DEUT|25|4|「牛在踹穀的時候，不可籠住牠的嘴。」
DEUT|25|5|「兄弟住在一起，若其中一個死了，沒有兒子，死者的妻子就不可出去嫁給陌生人。她丈夫的兄弟應當盡兄弟的本分，娶她為妻，與她同房。
DEUT|25|6|婦人生的長子要歸在已故兄弟的名下，免得他的名在 以色列 中塗去了。
DEUT|25|7|那人若不情願娶他兄弟的妻子，他兄弟的妻子就要上到城門長老那裏，說：『我丈夫的兄弟拒絕在 以色列 中為他的兄弟留名，不願意為我盡兄弟的本分。』
DEUT|25|8|本城的長老就要召那人來，跟他談話。若他堅持說：『我不情願娶她。』
DEUT|25|9|他兄弟的妻子就要在長老眼前來到那人跟前，脫下他腳上的鞋，吐唾沫在他臉上，回應說：『凡不為兄弟建立家室的都要這樣待他。』
DEUT|25|10|在 以色列 中，他要以『脫鞋之家』聞名。」
DEUT|25|11|「若有人和弟兄爭鬥，其中一人的妻子近前去，為了救丈夫脫離那打丈夫之人的手，伸手抓住那人的下體，
DEUT|25|12|你就要砍斷婦人的手，你的眼不可顧惜。
DEUT|25|13|「你袋中不可有一大一小兩樣的法碼。
DEUT|25|14|你家裏不可有一大一小兩樣的伊法 。
DEUT|25|15|當用準確公正的法碼和伊法，好使你的日子在耶和華－你上帝所賜你的地上得以長久。
DEUT|25|16|因為行這一切不義之事的人都是耶和華－你上帝所憎惡的。」
DEUT|25|17|「你要記得你們出 埃及 的時候， 亞瑪力 在路上怎樣對待你，
DEUT|25|18|在路上迎擊你，趁你疲乏困倦時擊殺所有在你後面軟弱的人；並不敬畏上帝。
DEUT|25|19|所以，當耶和華－你的上帝使你不被四圍一切仇敵擾亂，在耶和華－你上帝賜你為業的地上得享平靜的時候，你要把 亞瑪力 的名從天下塗去；你不可忘記這事。」
DEUT|26|1|「你進去得了耶和華－你上帝所賜你為業的地，並且居住在那裏的時候，
DEUT|26|2|就要從耶和華－你上帝所賜你的地上，將收成的各種初熟土產取一些來，盛在筐子裏，帶到那裏，耶和華－你上帝選擇作為他名居所的地方，
DEUT|26|3|到當時的祭司那裏，對他說：『我今日向耶和華－你的上帝宣認，我已來到耶和華向我們列祖起誓要賜給我們的地。』
DEUT|26|4|祭司就從你手裏把筐子接過來，供在耶和華－你上帝的祭壇前。
DEUT|26|5|你要在耶和華－你上帝面前告白說：『我的祖先原是一個流亡的 亞蘭 人，帶著稀少的人丁下到 埃及 寄居。在那裏，他卻成了又大又強、人數眾多的國。
DEUT|26|6|埃及 人惡待我們，迫害我們，將苦工加在我們身上。
DEUT|26|7|於是我們哀求耶和華我們列祖的上帝。耶和華聽見我們的聲音，看見我們所受的困苦、勞役和欺壓，
DEUT|26|8|耶和華就用大能的手和伸出來的膀臂，以及大而可畏的事和神蹟奇事，領我們出了 埃及 ，
DEUT|26|9|將我們領進這地方，把這流奶與蜜之地賜給我們。
DEUT|26|10|耶和華啊，看哪，現在我把你所賜我地上初熟的土產供上。』隨後你要把筐子供在耶和華－你上帝面前，向耶和華－你的上帝下拜。
DEUT|26|11|你和 利未 人，以及在你中間寄居的，要因耶和華－你上帝所賜你和你家的一切福分歡樂。
DEUT|26|12|「每逢第三年，就是捐十分之一的那年，你從你一切土產中取了十分之一，要分給 利未 人、寄居的、孤兒和寡婦，使他們在你的城鎮中可以吃得飽足。
DEUT|26|13|你又要在耶和華－你上帝面前說：『我已將聖物從家裏拿出來，給了 利未 人、寄居的、孤兒和寡婦，是遵照你吩咐我的一切命令。你的命令，我沒有違背，也沒有忘記。
DEUT|26|14|我守喪的時候，沒有吃這聖物，不潔淨的時候，也沒有拿出來，又沒有把它獻給死人。我聽從了耶和華－我上帝的話，都照你一切所吩咐的做了。
DEUT|26|15|求你從天上，從你的聖所垂看，賜福給你的百姓 以色列 和你向我們列祖起誓所賜給我們的這片土地，就是流奶與蜜之地。』」
DEUT|26|16|「耶和華－你的上帝今日吩咐你遵行這些律例典章，所以你要盡心盡性謹守遵行。
DEUT|26|17|你今日宣認耶和華為你的上帝，承諾遵行他的道，謹守他的律例、誡命、典章，聽從他的話。
DEUT|26|18|耶和華今日照他所應許你的，也認你為他寶貴的子民，叫你謹守他的一切誡命，
DEUT|26|19|要使你得稱讚、美名、尊榮，超乎他所造的萬國之上，並且照他所應許的，使你歸耶和華－你的上帝為神聖的子民。」
DEUT|27|1|摩西 和 以色列 的眾長老吩咐百姓說：「你們要遵守我今日所吩咐的一切誡命。
DEUT|27|2|你們過了 約旦河 ，到耶和華－你上帝所賜給你的地，當日要豎立幾塊大石頭，塗上石灰。
DEUT|27|3|當你過了河，進入耶和華－你上帝所賜給你流奶與蜜之地，正如耶和華－你列祖的上帝所應許你的，你要把這律法的一切話寫在石頭上。
DEUT|27|4|你們過了 約旦河 ，就要在 基利心山 上照我今日所吩咐的，把這些石頭豎立起來，塗上石灰。
DEUT|27|5|你在那裏要為耶和華－你的上帝築一座石壇，卻不可動用鐵器在石頭上。
DEUT|27|6|要用沒有鑿過的石頭築耶和華－你上帝的壇，在壇上將燔祭獻給耶和華－你的上帝，
DEUT|27|7|又要獻平安祭，在那裏吃，在耶和華－你的上帝面前歡樂。
DEUT|27|8|你要將這律法的一切話清楚地寫在石頭上。」
DEUT|27|9|摩西 和 利未 家的祭司吩咐 以色列 眾人說：「 以色列 啊，你要靜默傾聽！你今日已成為耶和華－你上帝的子民了。
DEUT|27|10|你要聽從耶和華－你上帝的話，遵行他的誡命律例，就是我今日所吩咐你的。」
DEUT|27|11|當日， 摩西 吩咐百姓說：
DEUT|27|12|「你們過了 約旦河 ， 西緬 、 利未 、 猶大 、 以薩迦 、 約瑟 和 便雅憫 等支派的人要站在 基利心山 上為百姓祝福。
DEUT|27|13|呂便 、 迦得 、 亞設 、 西布倫 、 但 和 拿弗他利 等支派的人要站在 以巴路山 上宣佈詛咒。
DEUT|27|14|利未 人要大聲對 以色列 眾人說：
DEUT|27|15|「『凡製造耶和華所憎惡的偶像，無論是雕刻的，是鑄造的，就是工匠用手造的，或暗中設置的，這人必受詛咒！』眾百姓要回應說：『阿們！』
DEUT|27|16|「『輕慢父母的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|17|「『挪移鄰舍地界的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|18|「『引領瞎子走錯路的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|19|「『對寄居的、孤兒和寡婦屈枉正直的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|20|「『與繼母同寢的，必受詛咒！因為他掀開父親衣服的下邊。』眾百姓要說：『阿們！』
DEUT|27|21|「『與獸交合的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|22|「『與同父異母，或同母異父的姊妹同寢的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|23|「『與岳母同寢的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|24|「『暗中擊殺鄰舍的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|25|「『受賄賂擊殺人而流無辜之血的，必受詛咒！』眾百姓要說：『阿們！』
DEUT|27|26|「『不堅守遵行這律法之話的，必受詛咒！』眾百姓要說：『阿們！』」
DEUT|28|1|「你若留心聽從耶和華－你上帝的話，謹守遵行他的一切誡命，就是我今日所吩咐你的，他必使你超乎地上的萬國之上。
DEUT|28|2|你若聽從耶和華－你上帝的話，這一切的福氣必臨到你身上，追隨你：
DEUT|28|3|你在城裏必蒙福，在田間也必蒙福。
DEUT|28|4|你身所生的，你地所產的，你牲畜所生的，牛犢、羔羊，都必蒙福。
DEUT|28|5|你的筐子和你的揉麵盆都必蒙福。
DEUT|28|6|你出也蒙福，入也蒙福。
DEUT|28|7|「耶和華必使那起來攻擊你的仇敵在你面前潰敗。他們從一條路來攻擊你，必在你面前從七條路逃跑。
DEUT|28|8|在你倉房裏，以及你手所做的一切，耶和華必發令賜福給你。耶和華－你上帝也必在所賜你的地上賜福給你。
DEUT|28|9|你若謹守耶和華－你上帝的誡命，遵行他的道，他必照他向你所起的誓立你為自己神聖的子民。
DEUT|28|10|地上的萬民見你歸在耶和華的名下，就必懼怕你。
DEUT|28|11|在耶和華向你列祖起誓應許賜你的土地上，他必使你身所生的，牲畜所生的，地所產的，都豐富有餘。
DEUT|28|12|耶和華必為你敞開天上的寶庫，按時降雨在你的地上。他必賜福你手裏所做的一切。你必借給許多國家，卻不必去借貸。
DEUT|28|13|你若聽從耶和華－你上帝的誡命，就是我今日所吩咐你的，謹守遵行，耶和華就必使你作首不作尾，居上不居下，
DEUT|28|14|只要你不偏左右，不背離我今日所吩咐你的一切話，也不隨從別神，事奉它們。」
DEUT|28|15|「你若不聽從耶和華－你上帝的話，不謹守遵行他的一切誡命律例，就是我今日所吩咐你的，這一切的詛咒必臨到你身上，追隨你：
DEUT|28|16|你在城裏必受詛咒，在田間也必受詛咒。
DEUT|28|17|你的筐子和你的揉麵盆都必受詛咒。
DEUT|28|18|你身所生的，你地所產的，以及牛犢、羔羊，都必受詛咒。
DEUT|28|19|你出也受詛咒，入也受詛咒。
DEUT|28|20|耶和華因你作惡離棄他，必在你手裏所做的一切，使詛咒、困擾、責罰臨到你，直到你被除滅，直到你迅速滅亡。
DEUT|28|21|耶和華必使瘟疫緊貼著你，直到他把你從所進去得為業的地上滅絕。
DEUT|28|22|耶和華要用癆病、熱病、發炎、高燒、刀劍 、焚風 和霉爛攻擊你；這些要追趕你，直到你滅亡。
DEUT|28|23|你頭上的天要變成銅，下面的地要化為鐵。
DEUT|28|24|耶和華要使那降在你地上的雨變為灰塵，塵土從天落在你身上，直到你被除滅。
DEUT|28|25|「耶和華必使你在仇敵面前潰敗。你從一條路去攻擊他們，必從七條路逃跑。地上萬國必因你而驚駭。
DEUT|28|26|你的屍首必給空中的飛鳥和地上的走獸作食物，卻無人鬨趕。
DEUT|28|27|耶和華必用 埃及 人的瘡、潰瘍、癬和疥攻擊你，使你不得醫治。
DEUT|28|28|耶和華必用癲狂、眼瞎、心驚攻擊你。
DEUT|28|29|你必在午間摸索，好像盲人在黑暗中摸索。你的道路必不亨通，天天受人欺壓、搶奪，無人搭救。
DEUT|28|30|你聘了妻子，別人必與她同寢；你建了房屋，卻不得住在其內；你栽植了葡萄園，卻不得享用所結的果子。
DEUT|28|31|你的牛在你眼前宰了，你吃不到牠的肉；你的驢在你眼前被人搶奪，卻討不回來；你的羊被敵人拿走，無人幫助你。
DEUT|28|32|你的兒女被交給別國的民；你的眼目終日切望，甚至失明，你的手卻無能為力。
DEUT|28|33|你地所產的和你勞力所得的，必被你所不認識的百姓吃盡。你天天只被欺負，受壓制，
DEUT|28|34|甚至你因眼中所見的景象而瘋狂。
DEUT|28|35|耶和華必攻擊你，使你膝上腿上，從腳掌到頭頂，都長滿了毒瘡，無法醫治。
DEUT|28|36|「耶和華必將你和你所立統治你的王，領到你和你列祖不認識的國去；在那裏你必事奉別神，就是木頭和石頭。
DEUT|28|37|你在耶和華趕你到的萬民中，要令人驚駭，成為笑柄，被人譏誚。
DEUT|28|38|你撒在田裏的種子雖多，收的卻少，因為蝗蟲把它吃光了。
DEUT|28|39|你栽植修整葡萄園，卻沒有酒喝，也不得儲存，因為蟲子把它吃了。
DEUT|28|40|你全境有橄欖樹，卻得不到油抹身，因為你的橄欖都掉光了。
DEUT|28|41|你生兒育女，卻不屬於你，因為他們必被擄去。
DEUT|28|42|你所有的樹木和你地裏的出產必被蝗蟲吃盡了。
DEUT|28|43|在你中間寄居的必上升高過你，高而又高；你必下降，低而又低。
DEUT|28|44|他必借給你，你卻不能借給他；他必作首，你必作尾。
DEUT|28|45|這一切的詛咒必臨到你，追趕你，趕上你，直到把你除滅，因為你不聽從耶和華－你上帝的話，不遵守他吩咐的誡命律例。
DEUT|28|46|這些詛咒必在你和你後裔身上成為神蹟奇事，直到永遠！
DEUT|28|47|因為你富裕的時候，不以歡喜快樂的心事奉耶和華－你的上帝，
DEUT|28|48|所以你必在飢餓、乾渴、赤身、缺乏中事奉仇敵，那是耶和華派來攻擊你的。他必把鐵軛加在你的頸項上，直到把你除滅。
DEUT|28|49|耶和華要從遠方、地極之處帶一國來，如鷹飛來攻擊你；這國的語言，你聽不懂。
DEUT|28|50|這國的人面貌兇惡，不給長者面子，也不恩待年輕人。
DEUT|28|51|他們必吃你牲畜所生的和你土地所產的，直到你被除滅。你的五穀、新酒和新的油，以及牛犢、羔羊，他都不給你留下，直到使你滅亡。
DEUT|28|52|他們必在你的各城圍困你，直到你在全地所倚靠、高大堅固的城牆都倒塌。他們必在耶和華－你上帝所賜給你全地的各城圍困你。
DEUT|28|53|你在仇敵圍困的窘迫中，必吃你本身所生的，就是耶和華－你上帝所賜給你的兒女之肉。
DEUT|28|54|你中間，連那溫和文雅的人都必冷眼惡待自己的兄弟和懷中的妻子，以及他所剩下其餘的兒女，
DEUT|28|55|不把所吃兒女的肉分一點給他們任何一個人，因為在被仇敵圍困、陷入窘迫的各城中，他已經一無所剩了。
DEUT|28|56|你中間柔順嬌嫩的婦人，甚至因柔順嬌嫩腳不肯踏地的婦人，也必冷眼惡待她懷中的丈夫和自己的兒女。
DEUT|28|57|在被仇敵圍困、陷入窘迫的城鎮中，她因缺乏一切，就要暗中把從她兩腿中間出來的胞衣和所生下的兒女吃了。
DEUT|28|58|「這書上所寫律法的一切話，是叫你敬畏耶和華－你上帝尊榮可畏的名，你若不謹守遵行，
DEUT|28|59|耶和華就必將奇異的災害，就是嚴重持久的災害和長期難治的疾病，加在你和你後裔的身上。
DEUT|28|60|他必使你所畏懼、 埃及 一切的疾病臨到你，緊貼著你，
DEUT|28|61|沒有寫在這律法書上的各樣疾病、災害，耶和華也必降在你身上，直到你被除滅。
DEUT|28|62|你們雖然曾像天上的星那樣多，卻因不聽從耶和華－你上帝的話，所剩的人丁就稀少了。
DEUT|28|63|耶和華先前怎樣喜愛善待你們，使你們增多，耶和華也要照樣喜愛消滅你們，使你們滅絕。你們必從所要進去得為業的地上被拔除。
DEUT|28|64|耶和華必把你們分散在萬民中，從地的這邊到地的另一邊，在那裏你必事奉你和你列祖不認識的神明，就是木頭和石頭。
DEUT|28|65|在那些國中，你必得不到安寧，腳掌也沒有安歇之處；耶和華卻要使你在那裏心中發顫，眼目失明，精神沮喪。
DEUT|28|66|你的一生懸空不安；你晝夜恐懼，生命沒有保障。
DEUT|28|67|你因心中的恐懼，眼睛所見的景象，早晨必說：『但願現在是晚上！』晚上必說：『但願現在是早晨！』
DEUT|28|68|耶和華要用船把你送回 埃及 去，走那我曾告訴你不再看見的路；在那裏你們必賣身給你的仇敵作奴婢，卻沒有人要買。」
DEUT|29|1|耶和華在 何烈山 與 以色列 人立約以外，這是耶和華在 摩押 地吩咐 摩西 與 以色列 人立約的話。
DEUT|29|2|摩西 召全 以色列 來，對他們說：「耶和華在 埃及 地，在你們眼前向法老和他眾臣僕，以及他的全地所做的一切事，你們都看見了，
DEUT|29|3|就是你親眼看見的大考驗，那些神蹟和大奇事。
DEUT|29|4|但耶和華到今日還沒有使你們心能明白，眼能看見，耳能聽見。
DEUT|29|5|我領你們在曠野四十年，你們身上的衣服沒有穿破，腳上的鞋也沒有穿壞；
DEUT|29|6|你們沒有吃餅，也沒有喝清酒烈酒，好讓你們知道『我─耶和華是你們的上帝』。
DEUT|29|7|你們來到這地方， 希實本 王 西宏 和 巴珊 王 噩 出來迎擊我們，與我們交戰，我們擊敗了他們，
DEUT|29|8|取了他們的地，給 呂便 支派、 迦得 支派和 瑪拿西 半支派為業。
DEUT|29|9|所以你們要謹守這約的話，遵行它們，好使你們在一切所做的事上亨通。
DEUT|29|10|「今日你們全都要站在耶和華－你們的上帝面前，就是各領袖、族長 、長老、官長、 以色列 所有的男子、
DEUT|29|11|你們的妻子兒女、你營中寄居的，從為你砍柴到為你挑水的人，
DEUT|29|12|為要使你進入耶和華－你上帝的約，就是耶和華－你上帝今日向你起誓所立的；
DEUT|29|13|這樣，他今日要立你作他的子民，他作你的上帝，是照他向你所應許的，又照他向你列祖 亞伯拉罕 、 以撒 、 雅各 所起的誓。
DEUT|29|14|我不單單與你們立這約，起這誓，
DEUT|29|15|就是今日與我們一同站在耶和華－我們上帝面前的，而且也包括今日不在我們這裏的人。
DEUT|29|16|「你們知道，我們曾住過 埃及 地，也經過列國，從他們中間穿越。
DEUT|29|17|你們也見過他們的可憎之物，他們木、石、金、銀的偶像。
DEUT|29|18|惟恐你們中間有人，或男或女，或宗族或支派，今日心裏偏離耶和華－我們的上帝，去事奉那些國的神明，又怕你們中間有根長出苦菜和茵蔯來。
DEUT|29|19|這樣的人聽見這詛咒的話，心裏還慶幸，說：『我雖然隨著頑固的心行事，卻還是平安無事。』以致有水的和無水的都消滅了。
DEUT|29|20|耶和華必不願饒恕他；耶和華的怒氣與妒忌必向他如煙冒出，將這書上所寫的一切詛咒都加在他身上，耶和華也要從天下塗去他的名。
DEUT|29|21|耶和華又必照著寫在律法書上，約中的一切詛咒，將他從 以色列 眾支派中分別出來，使他遭受禍害。
DEUT|29|22|你們的後代，就是接續你們興起的子孫，和遠方來的外邦人，看見這地的災禍，以及耶和華所降於這地的疾病，
DEUT|29|23|遍地都被硫磺和鹽所侵蝕，不能耕種，沒有出產，連草都長不出來，好像耶和華在怒氣和憤怒中所傾覆的 所多瑪 、 蛾摩拉 、 押瑪 、 洗扁 一樣，
DEUT|29|24|萬國必說：『耶和華為甚麼向此地這樣做呢？為甚麼要大發烈怒呢？』
DEUT|29|25|人必說：『這是因為這地的人離棄了耶和華─他們列祖的上帝領他們出 埃及 地的時候與他們所立的約，
DEUT|29|26|去事奉別神，敬拜他們所不認識的神明，這是耶和華未曾允許的。
DEUT|29|27|所以耶和華的怒氣向這地發作，將這書上所寫的一切詛咒都降在這地上。
DEUT|29|28|耶和華在怒氣、憤怒、大惱恨中將他們從本地拔出來，扔到別的地上，像今日一樣。』
DEUT|29|29|「隱祕的事是屬耶和華─我們上帝的，但明顯的事是永遠屬我們和我們子孫的，為要叫我們遵行這律法上的一切話。」
DEUT|30|1|「當這一切的事，就是我擺在你面前的祝福和詛咒臨到你的時候，你在耶和華－你上帝趕逐你去的萬國中，心裏回想這些事，
DEUT|30|2|你和你的子孫若盡心盡性歸向耶和華－你的上帝，照我今日一切所吩咐你的，聽從他的話，
DEUT|30|3|耶和華－你的上帝就必憐憫你，使你這被擄的子民歸回。耶和華－你的上帝必轉回，從分散你到的萬民中把你召集回來。
DEUT|30|4|你就是被趕逐到天涯，耶和華－你的上帝也必從那裏召集你，從那裏領你回來。
DEUT|30|5|耶和華－你的上帝必領你進入你列祖所得的地，你必得著這地為業。他必善待你，使你增多，勝過你的列祖。
DEUT|30|6|耶和華－你的上帝要使你的心和你後裔的心受割禮，好叫你盡心盡性愛耶和華－你的上帝，使你可以存活。
DEUT|30|7|耶和華－你的上帝必將這一切詛咒加在你仇敵和恨惡你、迫害你的人身上。
DEUT|30|8|你必回轉，聽從耶和華的話，遵行他的一切誡命，就是我今日所吩咐你的。
DEUT|30|9|耶和華－你的上帝必使你手裏所做的一切，以及你身所生的，牲畜所生的，土地所產的都豐富有餘，而且順利；耶和華必再喜愛善待你，正如他喜愛你的列祖一樣，
DEUT|30|10|只要你聽從耶和華－你上帝的話，謹守這律法書上所寫的誡命律例，盡心盡性歸向耶和華－你的上帝。」
DEUT|30|11|「我今日所吩咐你的誡命，對你並不困難，也不太遠；
DEUT|30|12|不是在天上，使你說：『誰為我們上天去取來給我們，使我們聽了可以遵行呢？』
DEUT|30|13|也不是在海的那邊，使你說：『誰為我們渡海到另一邊，去取來給我們，使我們聽了可以遵行呢？』
DEUT|30|14|因這話離你很近，就在你口中，在你心裏，使你可以遵行。
DEUT|30|15|「看，我今日將生死禍福擺在你面前。
DEUT|30|16|我今日所吩咐你的 ，就是要愛耶和華－你的上帝，遵行他的道，謹守他的誡命、律例、典章，使你可以存活，增多，而且耶和華－你的上帝必在你所要進去得為業的地上賜福給你。
DEUT|30|17|倘若你的心偏離，不肯聽從，卻被引誘去敬拜別神，事奉它們，
DEUT|30|18|我今日向你們申明，你們必定滅亡；在你過 約旦河 進去得為業的地上，你的日子必不長久。
DEUT|30|19|我今日呼天喚地向你作見證：我已經將生與死，祝福與詛咒，擺在你面前。所以你要揀選生命，好使你和你的後裔都得存活。
DEUT|30|20|要愛耶和華－你的上帝，聽從他的話，緊緊跟隨他，因為他是你的生命，必使你的日子得以長久，可以在耶和華向你列祖 亞伯拉罕 、 以撒 、 雅各 起誓要給他們的地上居住。」
DEUT|31|1|摩西 去把這些話吩咐 以色列 眾人 ，
DEUT|31|2|對他們說：「我已經一百二十歲了，現在不能照常出入。耶和華曾對我說：『你不得過這 約旦河 。』
DEUT|31|3|耶和華－你的上帝必在你面前過河，把這些國從你面前除滅，你就必得他們的地。 約書亞 要在你面前過河，是照耶和華所吩咐的。
DEUT|31|4|耶和華必對待他們，如同從前待他所除滅的 亞摩利 人的王 西宏 與 噩 ，以及他們的國一樣。
DEUT|31|5|耶和華必將他們交在你們面前，你們要照我所吩咐的一切命令待他們。
DEUT|31|6|你們當剛強壯膽，不要害怕，也不要畏懼他們，因為耶和華－你的上帝必與你同去；他必不撇下你，也不丟棄你。」
DEUT|31|7|摩西 召了 約書亞 來，在 以色列 眾人眼前對他說：「你當剛強壯膽！因為你要和這百姓一同進入 耶和華向他們列祖起誓要給他們的地，你也要使他們承受那地為業。
DEUT|31|8|耶和華必在你前面行，他必親自與你同在，必不撇下你，也不丟棄你。你不要懼怕，也不要驚惶。」
DEUT|31|9|摩西 寫下這律法，交給抬耶和華約櫃的 利未 人祭司和 以色列 的眾長老。
DEUT|31|10|摩西 吩咐他們說：「每逢七年的最後一年，就是定期的豁免年，在住棚節的時候，
DEUT|31|11|當 以色列 眾人來到耶和華－你上帝所選擇的地方朝見他的時候，你要在 以色列 眾人面前念這律法給他們聽。
DEUT|31|12|要召集百姓，男人、女人、孩子，和在你城裏寄居的，叫他們都得以聽見，好學習敬畏耶和華－你們的上帝，謹守遵行這律法的一切話。
DEUT|31|13|他們的兒女，就是那未曾認識的，也可以聽，學習敬畏耶和華－你們的上帝；你們一生的日子，在你們過 約旦河 得為業的地上，都要這樣做。」
DEUT|31|14|耶和華對 摩西 說：「看哪，你的死期已近了。要召 約書亞 來，和你一起站在會幕裏，我好吩咐他。」於是 摩西 和 約書亞 去站在會幕裏。
DEUT|31|15|耶和華在會幕裏，在雲柱中顯現，雲柱停在會幕門口的上面。
DEUT|31|16|耶和華對 摩西 說：「看哪，你必和你的祖先同睡。這百姓要起來，在他們所要去的地上，在那地的人中，隨從外邦的神明行淫，離棄我，違背我與他們所立的約。
DEUT|31|17|那時，我的怒氣必向他們發作，我必離棄他們，轉臉不顧他們，以致他們被吞滅，並有許多的禍患災難臨到他們。在那日，人必說：『這些禍患臨到我，豈不是因為我的上帝不在我中間嗎？』
DEUT|31|18|在那日，因人偏向別神所行的一切惡事，我必定轉臉不顧。
DEUT|31|19|現在你們要寫下這首歌，教導 以色列 人，放在他們口中，使這首歌成為我指責 以色列 人的見證。
DEUT|31|20|因為我將他們領進我向他們列祖起誓應許那流奶與蜜之地，他們在那裏吃得飽足，長得肥胖，就偏向別神，事奉它們，藐視我，背棄我的約。
DEUT|31|21|當許多禍患災難臨到他們的時候，這首歌必在他們面前作見證，因為他們後裔的口必吟誦不忘。我未領他們到我所起誓應許之地以先，他們所懷的意念我都知道了。」
DEUT|31|22|當日 摩西 就寫了一首歌，教導 以色列 人。
DEUT|31|23|耶和華吩咐 嫩 的兒子 約書亞 說：「你當剛強壯膽，因為你必領 以色列 人進入我所起誓應許他們的地，我必與你同在。」
DEUT|31|24|當 摩西 把這律法的話寫完在書上，到完成的時候，
DEUT|31|25|摩西 吩咐抬耶和華約櫃的 利未 人說：
DEUT|31|26|「把這律法書拿來，放在耶和華－你們上帝的約櫃旁，可以在那裏作指責你們的見證。
DEUT|31|27|因為我知道你們是悖逆的，是硬著頸項的。看哪，我今日還活著與你們同在，你們尚且悖逆耶和華，何況我死後呢？
DEUT|31|28|你們要召集你們支派的眾長老和官長到我這裏來，我好把這些話說給他們聽，並且呼喚天地見證他們的不是。
DEUT|31|29|我知道我死後你們必全然敗壞，偏離我所吩咐你們的道。日後必有禍患臨到你們，因為你們做了耶和華眼中看為惡的事，以你們手中所做的惹他發怒。」
DEUT|31|30|摩西 把這首歌的話，從頭到尾吟誦給 以色列 全會眾聽。
DEUT|32|1|「諸天哪，要側耳聽我說話； 願地聆聽我口中的言語。
DEUT|32|2|我的教導要淋漓如雨， 我的言語要滴落如露， 如細雨降在嫩草上， 如甘霖降在蔬菜中。
DEUT|32|3|因為我要宣揚耶和華的名， 你們要把偉大歸給我們的上帝。
DEUT|32|4|「他是磐石，他的作為完全， 他一切所行的都公平； 他是信實無偽的上帝， 又公義，又正直。
DEUT|32|5|這乖僻彎曲的世代 向他行了敗壞的事； 因著他們的弊病， 不再是他的兒女。
DEUT|32|6|愚昧無知的百姓啊， 你們這樣報答耶和華嗎？ 他豈不是你的父，創造了你嗎？ 他造了你，堅立你。
DEUT|32|7|你當回想上古之日， 思念歷代之年； 問你的父親，他必告訴你； 問你的長者，他必向你述說。
DEUT|32|8|至高者將地業賜給列國， 將世人分開， 他按照神明 的數目， 為萬民劃定疆界。
DEUT|32|9|因為耶和華的份是他的百姓， 他的產業就是 雅各 。
DEUT|32|10|「耶和華在曠野之地， 在空曠，野獸吼叫之荒地遇見他， 就環繞他，看顧他， 保護他，如同保護眼中的瞳人。
DEUT|32|11|鷹怎樣攪動巢窩， 在雛鷹上面飛翔， 展開雙翅接住雛鷹， 背在兩翼之上，
DEUT|32|12|耶和華也照樣獨自引導他， 並無外邦神明與他同在。
DEUT|32|13|耶和華使他馳騁在地的高處， 他吃田間的出產； 耶和華使他從巖石中吃蜜， 從堅石中吸油，
DEUT|32|14|也吃牛的乳酪、羊的奶、 羔羊的脂肪， 巴珊 所出的公綿羊和山羊， 和上好的麥子。 你要喝葡萄汁釀的美酒。
DEUT|32|15|「 耶書崙 漸漸肥胖，能踼跳。 你長得肥胖，粗壯，豐潤。 他離棄造他的上帝， 輕看救他的磐石。
DEUT|32|16|他們用外邦神明惹上帝妒忌， 以可憎之物惹他發怒。
DEUT|32|17|他們祭祀鬼魔，而非上帝， 是他們不認識的神明， 是近來新興的， 是你們列祖所不畏懼的。
DEUT|32|18|你輕忽生你的磐石， 忘記生產你的上帝。
DEUT|32|19|「耶和華看見了， 因他兒女惹動他就拋棄他們，
DEUT|32|20|說：『我要轉臉離開他們， 看他們的結局如何。 他們是極乖謬的世代， 是不忠實的兒女。
DEUT|32|21|他們以那不是上帝的激起我妒忌， 以虛無的神明 惹我發怒。 我也要以不成國的激起你們嫉妒， 我要以愚頑的國惹起你們發怒。
DEUT|32|22|因為我的怒火焚燒， 直燒到極深的陰間， 吞噬地和地的出產， 連山的根基也燒著了。
DEUT|32|23|「『我要把禍患堆在他們身上， 我用盡我的箭射向他們：
DEUT|32|24|餓死人的饑荒、 灼人的熱症、 痛苦的災害。 我要叫野獸用牙齒咬他們， 叫土中爬行的用毒液害他們。
DEUT|32|25|外有刀劍使人喪亡， 內有驚恐， 少男少女是如此， 吃奶的、白髮的也是如此。
DEUT|32|26|我曾說，我要粉碎他們， 使他們的名 從人間消失。
DEUT|32|27|惟恐仇敵挑釁， 他們的敵人誤解， 說，我們的手得勝了， 這一切並非耶和華做的。』
DEUT|32|28|「因為他們是缺乏智謀的國家， 他們裏面毫無聰明。
DEUT|32|29|惟願他們有智慧，能明白這事， 他們就會想到自己的結局。
DEUT|32|30|若非他們的磐石賣了他們， 若非耶和華交出他們， 一人豈能追趕千人， 二人焉能使萬人逃跑呢？
DEUT|32|31|甚至我們的仇敵都承認， 他們的磐石不如我們的磐石。
DEUT|32|32|他們的葡萄樹是 所多瑪 的葡萄樹， 是 蛾摩拉 田園所長的； 他們的葡萄是毒葡萄， 整串都是苦的。
DEUT|32|33|他們的酒是大蛇的毒液， 是毒蛇劇烈的毒汁。
DEUT|32|34|「這豈不都存放在我這裏， 封存在我庫房中嗎？
DEUT|32|35|伸冤報應在我 ， 到了時候他們會失腳。 因為他們遭難的日子近了， 他們的厄運快要臨到。
DEUT|32|36|耶和華見他的百姓毫無能力， 無論是為奴的、自由的，都沒有存留， 就必為他們伸冤， 為自己的僕人發憐憫。
DEUT|32|37|他必說：『他們的神明， 他們所投靠的磐石，在哪裏呢？
DEUT|32|38|吃了他們祭牲脂肪的， 喝了他們澆酒祭之酒的， 叫那些神明站出來幫助你們， 作為你們的保障吧！
DEUT|32|39|「『如今，看！我，惟有我是上帝 ； 我以外並無別神。 我使人死，我使人活； 我擊傷人，也醫治人， 沒有人能從我手中救出來。
DEUT|32|40|我向天舉手， 我憑我的永生起誓說：
DEUT|32|41|我若磨我閃亮的刀， 我的手掌握審判權， 就必報復我的敵人， 報應那些恨我的人。
DEUT|32|42|我要使我的箭飲血而醉， 就是被殺被擄之人的血； 我的刀也要吃肉， 就是仇敵披髮頭顱 的肉。』
DEUT|32|43|「列國啊，當與耶和華的子民一同歡呼 ； 因為他要為他僕人 所流的血伸冤， 報應他的敵人 ， 救贖他的土地和他的子民 。」
DEUT|32|44|摩西 和 嫩 的兒子 約書亞 前來把這首歌的一切話吟誦給百姓聽。
DEUT|32|45|摩西 向 以色列 眾人吟誦完了這一切話，
DEUT|32|46|對他們說：「我今日以這一切話警戒你們，你們都要記在心中，要吩咐你們的子孫謹守遵行這律法上一切的話。
DEUT|32|47|因為這不是與你們無關的空話，而是你們的生命；因遵行這話，你們的日子必在你們過 約旦河 得為業的地上得以長久。」
DEUT|32|48|就在那日，耶和華吩咐 摩西 說：
DEUT|32|49|「你上 摩押 地的 亞巴琳山脈 ，到面對 耶利哥 的 尼波山 去，看我所要賜給 以色列 人為業的 迦南 地。
DEUT|32|50|你必死在你所登的山上，歸到你祖先 那裏，像你哥哥 亞倫 死在 何珥山 上，歸到他祖先 那裏一樣。
DEUT|32|51|因為你們在 以色列 人中得罪了我，在 尋 的曠野， 加低斯 的 米利巴 水那裏，在 以色列 人中沒有尊我為聖。
DEUT|32|52|我所賜給 以色列 人的地，你只可從對面觀看，卻不得進到那裏去。」
DEUT|33|1|這是神人 摩西 未死以前為 以色列 人的祝福。
DEUT|33|2|他說： 「耶和華從 西奈 來， 從 西珥 向他們顯現， 從 巴蘭山 發出光輝； 從萬萬聖者中來臨 ， 從他右手向他們發出烈火的律法 。
DEUT|33|3|他實在疼愛萬民。 他的眾聖徒都在你手中， 他們坐在你的腳下， 領受你的言語。」
DEUT|33|4|摩西 將律法傳給我們， 作為 雅各 會眾的產業。
DEUT|33|5|「耶和華 在 耶書崙 作王； 百姓的眾領袖和 以色列 各支派一同歡聚。
DEUT|33|6|願 呂便 存活，不致死亡， 雖然他的人丁稀少。
DEUT|33|7|關於 猶大 ，他這麼說： 『耶和華啊，求你垂聽 猶大 的聲音， 引導他歸回他的百姓中。 他曾用手為自己爭戰， 你必幫助他攻擊敵人。』
DEUT|33|8|關於 利未 ，他說： 『願你的土明和烏陵都在你的虔誠人那裏 。 你在 瑪撒 曾考驗他， 在 米利巴 水與他爭論。
DEUT|33|9|關於自己的父母，他說：我未曾關注。 他的弟兄，他不承認， 他的兒女，他也不認識， 因為 利未 人遵行你的話， 謹守你的約。
DEUT|33|10|他們將你的典章教導 雅各 ， 將你的律法教導 以色列 。 他們奉上香讓你聞， 把全牲的燔祭獻在你壇上。
DEUT|33|11|求耶和華賜福給他的財物 ， 悅納他手裏的工作。 求你刺透起來攻擊他的人的腰， 使那些恨惡他的人不再起來。』
DEUT|33|12|關於 便雅憫 ，他說： 『耶和華所親愛的必同耶和華安然居住， 耶和華終日庇護他， 他也住在耶和華兩肩之中 。』
DEUT|33|13|關於 約瑟 ，他說： 『願他的地蒙耶和華賜福， 得天上的甘露， 地下的泉源；
DEUT|33|14|得太陽下的美果， 月光中的佳穀；
DEUT|33|15|得古老山嶽的至寶， 永恆山嶺的寶物；
DEUT|33|16|得地的寶物和其中所充滿的， 得住在荊棘中者的喜悅。 願這些福都臨到 約瑟 的頭上， 臨到那與兄弟有分別之人的頭頂上。
DEUT|33|17|他是牛群中頭生的， 大有威嚴； 他的雙角是野牛的角， 用以牴觸萬民，直到地極。 這對角是 以法蓮 的萬萬， 這對角是 瑪拿西 的千千。』
DEUT|33|18|關於 西布倫 ，他說： 『 西布倫 哪，你出外可以歡喜。 以薩迦 啊，你在帳棚裏可以快樂。
DEUT|33|19|他們要召集萬民到山上， 在那裏獻公義的祭。 因為他們要吸取海裏的財富， 沙中隱藏的珍寶。』
DEUT|33|20|關於 迦得 ，他說： 『那使 迦得 擴張的，當受稱頌！ 迦得 臥如母獅， 撕裂膀臂和頭皮。
DEUT|33|21|他為自己看中了最好的， 因為那是為掌權者所存留的一份。 他與百姓的領袖同來 ， 執行耶和華的公義 和耶和華為 以色列 所立的典章。』
DEUT|33|22|關於 但 ，他說： 『 但 是小獅子， 從 巴珊 跳出來。』
DEUT|33|23|關於 拿弗他利 ，他說： 『 拿弗他利 啊，你享足恩寵， 滿得耶和華的福， 可以得西方和南方為業。』
DEUT|33|24|關於 亞設 ，他說： 『願 亞設 在眾子中蒙福 ， 願他得他弟兄的喜悅， 可以把腳蘸在油中。
DEUT|33|25|你的門閂是鐵的，是銅的。 只要你有多少日子，你就有多少力量 。』
DEUT|33|26|「 耶書崙 哪，沒有誰能比上帝！ 他騰雲，大顯威榮， 從天空來幫助你。
DEUT|33|27|亙古的上帝是避難所， 下面有永久的膀臂。 他從你面前趕走仇敵， 說：『毀滅吧！』
DEUT|33|28|因此， 以色列 獨自安然居住， 雅各 的泉源在五穀新酒之地， 他的天也滴下露水。
DEUT|33|29|以色列 啊，你有福了！ 蒙耶和華拯救的百姓啊，誰能像你？ 他是幫助你的盾牌， 是你威榮的刀劍。 你的仇敵要屈身就你； 你卻要踐踏他們的背脊 。」
DEUT|34|1|摩西 從 摩押 平原登上 尼波山 ，到了 耶利哥 對面的 毗斯迦山 頂。耶和華把全地指給他看：從 基列 到 但 ，
DEUT|34|2|拿弗他利 全地， 以法蓮 、 瑪拿西 的地， 猶大 全地直到西邊的海，
DEUT|34|3|尼革夫 ，從棕樹城 耶利哥 的平原到 瑣珥 。
DEUT|34|4|耶和華對他說：「這就是我向 亞伯拉罕 、 以撒 、 雅各 起誓應許之地，說：『我必將這地賜給你的後裔。』現在我使你親眼看見了，你卻不得過到那裏去。」
DEUT|34|5|於是耶和華的僕人 摩西 死在 摩押 地那裏，正如耶和華所說的。
DEUT|34|6|耶和華將他葬在 摩押 地， 伯‧毗珥 對面的谷中，只是到今日，沒有人知道他的墳墓。
DEUT|34|7|摩西 死的時候一百二十歲，眼目沒有昏花，力量沒有衰退。
DEUT|34|8|以色列 人在 摩押 平原為 摩西 哀哭了三十天，為 摩西 哀哭居喪的日期才結束。
DEUT|34|9|嫩 的兒子 約書亞 ，因為 摩西 曾為他按手，他就被智慧的靈充滿。 以色列 人聽從他，照著耶和華所吩咐 摩西 的去做。
DEUT|34|10|以後， 以色列 中再沒有興起一位先知像 摩西 的，他是耶和華面對面所認識的。
DEUT|34|11|耶和華差派他在 埃及 地，向法老和他的一切臣僕，以及他的全地，行了各樣神蹟奇事，
DEUT|34|12|又在 以色列 眾人眼前顯出大能的手，行了一切大而可畏的事。
