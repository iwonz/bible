COL|1|1|Павло, із волі Божої апостол Христа Ісуса, і брат Тимофій
COL|1|2|до святих і вірних братів у Христі, що в Колосах: благодать вам і мир від Бога, Отця нашого!
COL|1|3|Ми дякуємо Богові, Отцеві Господа нашого Ісуса Христа, завжди за вас молячись,
COL|1|4|прочувши про вашу віру в Христа Ісуса та про любов, яку маєте до всіх святих
COL|1|5|через надію, приготовану в небі для вас, що про неї давніше ви чули в слові істини Євангелії,
COL|1|6|що до вас прибула, і на цілому світі плодоносна й росте, як і в вас, з того дня, коли ви почули й пізнали благодать Божу в правді.
COL|1|7|Отак ви і навчилися від Епафра, улюбленого співробітника нашого, що за вас він вірний служитель Христа,
COL|1|8|що й виявив нам про вашу духовну любов.
COL|1|9|Через це то й ми з того дня, як почули, не перестаємо молитись за вас та просити, щоб для пізнання волі Його були ви наповнені всякою мудрістю й розумом духовним,
COL|1|10|щоб ви поводилися належно щодо Господа в усякому догодженні, в усякому доброму ділі приносячи плід і зростаючи в пізнанні Бога,
COL|1|11|зміцняючись усякою силою за могучістю слави Його для всякої витривалости й довготерпіння з радістю,
COL|1|12|дякуючи Отцеві, що вчинив нас достойними участи в спадщині святих у світлі,
COL|1|13|що визволив нас із влади темряви й переставив нас до Царства Свого улюбленого Сина,
COL|1|14|в Якім маємо відкуплення і прощення гріхів.
COL|1|15|Він є образ невидимого Бога, роджений перш усякого творива.
COL|1|16|Бо то Ним створено все на небі й на землі, видиме й невидиме, чи то престоли, чи то господства, чи то влади, чи то начальства, усе через Нього й для Нього створено!
COL|1|17|А Він є перший від усього, і все Ним стоїть.
COL|1|18|І Він Голова тіла, Церкви. Він початок, первороджений з мертвих, щоб у всьому Він мав першенство.
COL|1|19|Бо вгодно було, щоб у Нім перебувала вся повнота,
COL|1|20|і щоб Ним поєднати з Собою все, примиривши кров'ю хреста Його, через Нього, чи то земне, чи то небесне.
COL|1|21|І вас, що були колись відчужені й вороги думкою в злих учинках,
COL|1|22|тепер же примирив смертю в людськім тілі Його, щоб учинити вас святими, і непорочними, і неповинними перед Собою,
COL|1|23|якщо тільки пробуваєте в вірі тверді та сталі, і не відпадаєте від надії Євангелії, що ви чули її, яка проповідана всьому створінню під небом, якій я, Павло, став служителем.
COL|1|24|Тепер я радію в стражданнях своїх за вас, і доповнюю недостачу скорботи Христової в тілі своїм за тіло Його, що воно Церква;
COL|1|25|якій я став служителем за Божим зарядженням, що для вас мені дане, щоб виконати Слово Боже,
COL|1|26|Таємницю, заховану від віків і поколінь, а тепер виявлену Його святим,
COL|1|27|що їм Бог захотів показати, яке багатство слави цієї таємниці між поганами, а вона Христос у вас, надія слави!
COL|1|28|Його ми проповідуємо, нагадуючи кожній людині й навчаючи кожну людину всякої мудрости, щоб учинити кожну людину досконалою в Христі.
COL|1|29|У тому й працюю я, борючися силою Його, яка сильно діє в мені.
COL|2|1|Я хочу, щоб ви знали, яку велику боротьбу я маю за вас і за тих, хто в Лаодикії, і за всіх, хто не бачив мого тілесного обличчя.
COL|2|2|Хай потішаться їхні серця, у любові поєднані, для всякого багатства повного розуміння, для пізнання таємниці Бога, Христа,
COL|2|3|в Якому всі скарби премудрости й пізнання заховані.
COL|2|4|А це говорю, щоб ніхто вас не звів фальшивими доводами при суперечці.
COL|2|5|Бо хоч тілом я й неприсутній, та духом я з вами, і з радістю бачу ваш порядок та твердість вашої віри в Христа.
COL|2|6|Отже, як ви прийняли були Христа Ісуса Господа, так і в Ньому ходіть,
COL|2|7|бувши вкорінені й збудовані на Ньому, та зміцнені в вірі, як вас навчено, збагачуючись у ній з подякою.
COL|2|8|Стережіться, щоб ніхто вас не звів філософією та марною оманою за переданням людським, за стихіями світу, а не за Христом,
COL|2|9|бо в Ньому тілесно живе вся повнота Божества.
COL|2|10|І ви маєте в Нім повноту, а Він Голова всякої влади й начальства.
COL|2|11|Ви в Ньому були й обрізані нерукотворним обрізанням, скинувши людське тіло гріховне в Христовім обрізанні.
COL|2|12|Ви були з Ним поховані у хрищенні, у Ньому ви й разом воскресли через віру в силу Бога, що Він з мертвих Його воскресив.
COL|2|13|І вас, що мертві були в гріхах та в необрізанні вашого тіла, Він оживив разом із Ним, простивши усі гріхи,
COL|2|14|знищивши рукописання на нас, що наказами було проти нас, Він із середини взяв його та й прибив його на хресті,
COL|2|15|роззброївши влади й начальства, сміливо їх вивів на посміховисько, перемігши їх на хресті!
COL|2|16|Тож, хай ніхто вас не судить за їжу, чи за питво, чи за чергове свято, чи за новомісяччя, чи за суботи,
COL|2|17|бо це тінь майбутнього, а тіло Христове.
COL|2|18|Нехай вас не зводить ніхто удаваною покорою та службою Анголам, вдаючися до того, чого не бачив, нерозважно надимаючись своїм тілесним розумом,
COL|2|19|а не тримачись Голови, від Якої все тіло, суглобами й зв'язями з'єднане й зміцнене, росте зростом Божим.
COL|2|20|Отож, як ви вмерли з Христом для стихій світу, то чого ви, немов ті, хто в світі живе, пристаєте на постанови:
COL|2|21|не дотикайся, ані їж, ані рухай,
COL|2|22|бо то все знищиться, як уживати його, за приказами та наукою людською.
COL|2|23|Воно ж має вид мудрости в самовільній службі й покорі та в знесилюванні тіла, та не має якогось значення, хіба щодо насичення тіла.
COL|3|1|Отож, коли ви воскресли з Христом, то шукайте того, що вгорі, де сидить Христос по Божій правиці.
COL|3|2|Думайте про те, що вгорі, а не про те, що на землі.
COL|3|3|Бож ви вмерли, а життя ваше сховане в Бозі з Христом.
COL|3|4|Коли з'явиться Христос, наше життя, тоді з'явитеся з Ним у славі і ви.
COL|3|5|Отож, умертвіть ваші земні члени: розпусту, нечисть, пристрасть, лиху пожадливість та зажерливість, що вона ідолослуження,
COL|3|6|бо гнів Божий приходить за них на неслухняних.
COL|3|7|І ви поміж ними ходили колись, як жили поміж ними.
COL|3|8|Тепер же відкиньте і ви все оте: гнів, лютість, злобу, богозневагу, безсоромні слова з ваших уст.
COL|3|9|Не кажіть неправди один на одного, якщо скинули з себе людину стародавню з її вчинками,
COL|3|10|та зодягнулися в нову, що відновлюється для пізнання за образом Створителя її,
COL|3|11|де нема ані геллена, ані юдея, обрізання та необрізання, варвара, скита, раба, вільного, але все та в усьому Христос!
COL|3|12|Отож, зодягніться, як Божі вибранці, святі та улюблені, у щире милосердя, добротливість, покору, лагідність, довготерпіння.
COL|3|13|Терпіть один одного, і прощайте собі, коли б мав хто на кого оскарження. Як і Христос вам простив, робіть так і ви!
COL|3|14|А над усім тим зодягніться в любов, що вона союз досконалости!
COL|3|15|І нехай мир Божий панує у ваших серцях, до якого й були ви покликані в одному тілі. І вдячними будьте!
COL|3|16|Слово Христове нехай пробуває в вас рясно, у всякій премудрості. Навчайте та напоумляйте самих себе! Вдячно співайте у ваших серцях Господеві псалми, гімни, духовні пісні!
COL|3|17|І все, що тільки робите словом чи ділом, усе робіть у Ім'я Господа Ісуса, дякуючи через Нього Богові й Отцеві.
COL|3|18|Дружини, слухайтеся чоловіків своїх, як лицює то в Господі!
COL|3|19|Чоловіки, любіть дружин своїх, і не будьте суворі до них!
COL|3|20|Діти, будьте слухняні в усьому батькам, бо це Господеві приємне!
COL|3|21|Батьки, не дратуйте дітей своїх, щоб на дусі не впали вони!
COL|3|22|Раби, слухайтеся в усьому тілесних панів, і не працюйте тільки про людське око, немов підлещуючись, але в простоті серця, боячися Бога!
COL|3|23|І все, що тільки чините, робіть від душі, немов Господеві, а не людям!
COL|3|24|Знайте, що від Господа приймете в нагороду спадщину, бо служите ви Господеві Христові.
COL|3|25|А хто кривдить, той одержить за свою кривду. Бо не дивиться Бог на особу!
COL|4|1|Пани, виявляйте до рабів справедливість та рівність, і знайте, що й для вас є на небі Господь!
COL|4|2|Будьте тривалі в молитві, і пильнуйте з подякою в ній!
COL|4|3|Моліться разом і за нас, щоб Бог нам відчинив двері слова, звіщати таємницю Христову, що за неї я й зв'язаний,
COL|4|4|щоб з'явив я її, як звіщати належить мені.
COL|4|5|Поводьтеся мудро з чужими, використовуючи час.
COL|4|6|Слово ваше нехай буде завжди ласкаве, приправлене сіллю, щоб ви знали, як ви маєте кожному відповідати.
COL|4|7|Що зо мною, то все вам розповість Тихик, улюблений брат і вірний служитель і співробітник у Господі.
COL|4|8|Я саме на те його вислав до вас, щоб довідались ви про нас, і щоб ваші серця він потішив,
COL|4|9|із Онисимом, вірним та улюбленим братом, який з-поміж вас. Вони все вам розповідять, що діється тут.
COL|4|10|Поздоровлює вас Аристарх, ув'язнений разом зо мною, і Марко, небіж Варнавин, що про нього ви дістали накази; як прийде до вас, то прийміть його,
COL|4|11|теж Ісус, на прізвище Юст, вони із обрізаних. Для Божого Царства єдині вони співробітники, що були мені втіхою.
COL|4|12|Поздоровлює вас Епафрас, що з ваших, раб Христа Ісуса. Він завжди обстоює вас у молитвах, щоб ви досконалі були та наповнені всякою Божою волею.
COL|4|13|І я свідчу за нього, що він має велику горливість про вас та про тих, що знаходяться в Лаодикії та в Гієраполі.
COL|4|14|Вітає вас Лука, улюблений лікар, та Димас.
COL|4|15|Привітайте братів, що в Лаодикії, і Німфана, і Церкву домашню його.
COL|4|16|І як буде прочитаний лист цей у вас, то зробіть, щоб прочитаний був він також у Церкві Лаодикійській, а того, що написаний з Лаодикії, прочитайте і ви.
COL|4|17|Та скажіть Архіпові: Доглядай того служіння, що прийняв його в Господі, щоб ти його виконав!
COL|4|18|Привітання моєю рукою Павловою. Пам'ятайте про пута мої! Благодать Божа нехай буде з вами! Амінь.
