HEB|1|1|multifariam et multis modis olim Deus loquens patribus in prophetis
HEB|1|2|novissime diebus istis locutus est nobis in Filio quem constituit heredem universorum per quem fecit et saecula
HEB|1|3|qui cum sit splendor gloriae et figura substantiae eius portansque omnia verbo virtutis suae purgationem peccatorum faciens sedit ad dexteram Maiestatis in excelsis
HEB|1|4|tanto melior angelis effectus quanto differentius prae illis nomen hereditavit
HEB|1|5|cui enim dixit aliquando angelorum Filius meus es tu ego hodie genui te et rursum ego ero illi in Patrem et ipse erit mihi in Filium
HEB|1|6|et cum iterum introducit primogenitum in orbem terrae dicit et adorent eum omnes angeli Dei
HEB|1|7|et ad angelos quidem dicit qui facit angelos suos spiritus et ministros suos flammam ignis
HEB|1|8|ad Filium autem thronus tuus Deus in saeculum saeculi et virga aequitatis virga regni tui
HEB|1|9|dilexisti iustitiam et odisti iniquitatem propterea unxit te Deus Deus tuus oleo exultationis prae participibus tuis
HEB|1|10|et tu in principio Domine terram fundasti et opera manuum tuarum sunt caeli
HEB|1|11|ipsi peribunt tu autem permanebis et omnes ut vestimentum veterescent
HEB|1|12|et velut amictum involves eos et mutabuntur tu autem idem es et anni tui non deficient
HEB|1|13|ad quem autem angelorum dixit aliquando sede a dextris meis quoadusque ponam inimicos tuos scabillum pedum tuorum
HEB|1|14|nonne omnes sunt administratorii spiritus in ministerium missi propter eos qui hereditatem capient salutis
HEB|2|1|propterea abundantius oportet observare nos ea quae audivimus ne forte pereffluamus
HEB|2|2|si enim qui per angelos dictus est sermo factus est firmus et omnis praevaricatio et inoboedientia accepit iustam mercedis retributionem
HEB|2|3|quomodo nos effugiemus si tantam neglexerimus salutem quae cum initium accepisset enarrari per Dominum ab eis qui audierunt in nos confirmata est
HEB|2|4|contestante Deo signis et portentis et variis virtutibus et Spiritus Sancti distributionibus secundum suam voluntatem
HEB|2|5|non enim angelis subiecit orbem terrae futurum de quo loquimur
HEB|2|6|testatus est autem in quodam loco quis dicens quid est homo quod memor es eius aut filius hominis quoniam visitas eum
HEB|2|7|minuisti eum paulo minus ab angelis gloria et honore coronasti eum et constituisti eum super opera manuum tuarum
HEB|2|8|omnia subiecisti sub pedibus eius in eo enim quod ei omnia subiecit nihil dimisit non subiectum ei nunc autem necdum videmus omnia subiecta ei
HEB|2|9|eum autem qui modico quam angeli minoratus est videmus Iesum propter passionem mortis gloria et honore coronatum ut gratia Dei pro omnibus gustaret mortem
HEB|2|10|decebat enim eum propter quem omnia et per quem omnia qui multos filios in gloriam adduxerat auctorem salutis eorum per passiones consummare
HEB|2|11|qui enim sanctificat et qui sanctificantur ex uno omnes propter quam causam non confunditur fratres eos vocare dicens
HEB|2|12|nuntiabo nomen tuum fratribus meis in medio ecclesiae laudabo te
HEB|2|13|et iterum ego ero fidens in eum et iterum ecce ego et pueri mei quos mihi dedit Deus
HEB|2|14|quia ergo pueri communicaverunt sanguini et carni et ipse similiter participavit hisdem ut per mortem destrueret eum qui habebat mortis imperium id est diabolum
HEB|2|15|et liberaret eos qui timore mortis per totam vitam obnoxii erant servituti
HEB|2|16|nusquam enim angelos adprehendit sed semen Abrahae adprehendit
HEB|2|17|unde debuit per omnia fratribus similare ut misericors fieret et fidelis pontifex ad Deum ut repropitiaret delicta populi
HEB|2|18|in eo enim in quo passus est ipse temptatus potens est eis qui temptantur auxiliari
HEB|3|1|unde fratres sancti vocationis caelestis participes considerate apostolum et pontificem confessionis nostrae Iesum
HEB|3|2|qui fidelis est ei qui fecit illum sicut et Moses in omni domo illius
HEB|3|3|amplioris enim gloriae iste prae Mose dignus habitus est quanto ampliorem honorem habet domus qui fabricavit illam
HEB|3|4|omnis namque domus fabricatur ab aliquo qui autem omnia creavit Deus
HEB|3|5|et Moses quidem fidelis erat in tota domo eius tamquam famulus in testimonium eorum quae dicenda erant
HEB|3|6|Christus vero tamquam filius in domo sua quae domus sumus nos si fiduciam et gloriam spei usque ad finem firmam retineamus
HEB|3|7|quapropter sicut dicit Spiritus Sanctus hodie si vocem eius audieritis
HEB|3|8|nolite obdurare corda vestra sicut in exacerbatione secundum diem temptationis in deserto
HEB|3|9|ubi temptaverunt me patres vestri probaverunt et viderunt opera mea
HEB|3|10|quadraginta annos propter quod infensus fui generationi huic et dixi semper errant corde ipsi autem non cognoverunt vias meas
HEB|3|11|sicut iuravi in ira mea si introibunt in requiem meam
HEB|3|12|videte fratres ne forte sit in aliquo vestrum cor malum incredulitatis discedendi a Deo vivo
HEB|3|13|sed adhortamini vosmet ipsos per singulos dies donec hodie cognominatur ut non obduretur quis ex vobis fallacia peccati
HEB|3|14|participes enim Christi effecti sumus si tamen initium substantiae usque ad finem firmum retineamus
HEB|3|15|dum dicitur hodie si vocem eius audieritis nolite obdurare corda vestra quemadmodum in illa exacerbatione
HEB|3|16|quidam enim audientes exacerbaverunt sed non universi qui profecti sunt ab Aegypto per Mosen
HEB|3|17|quibus autem infensus est quadraginta annos nonne illis qui peccaverunt quorum cadavera prostrata sunt in deserto
HEB|3|18|quibus autem iuravit non introire in requiem ipsius nisi illis qui increduli fuerunt
HEB|3|19|et videmus quia non potuerunt introire propter incredulitatem
HEB|4|1|timeamus ergo ne forte relicta pollicitatione introeundi in requiem eius existimetur aliqui ex vobis deesse
HEB|4|2|etenim et nobis nuntiatum est quemadmodum et illis sed non profuit illis sermo auditus non admixtis fidei ex his quae audierunt
HEB|4|3|ingrediemur enim in requiem qui credidimus quemadmodum dixit sicut iuravi in ira mea si introibunt in requiem meam et quidem operibus ab institutione mundi factis
HEB|4|4|dixit enim quodam loco de die septima sic et requievit Deus die septima ab omnibus operibus suis
HEB|4|5|et in isto rursum si introibunt in requiem meam
HEB|4|6|quoniam ergo superest quosdam introire in illam et hii quibus prioribus adnuntiatum est non introierunt propter incredulitatem
HEB|4|7|iterum terminat diem quendam hodie in David dicendo post tantum temporis sicut supra dictum est hodie si vocem eius audieritis nolite obdurare corda vestra
HEB|4|8|nam si eis Iesus requiem praestitisset numquam de alio loqueretur posthac die
HEB|4|9|itaque relinquitur sabbatismus populo Dei
HEB|4|10|qui enim ingressus est in requiem eius etiam ipse requievit ab operibus suis sicut a suis Deus
HEB|4|11|festinemus ergo ingredi in illam requiem ut ne in id ipsum quis incidat incredulitatis exemplum
HEB|4|12|vivus est enim Dei sermo et efficax et penetrabilior omni gladio ancipiti et pertingens usque ad divisionem animae ac spiritus conpagum quoque et medullarum et discretor cogitationum et intentionum cordis
HEB|4|13|et non est ulla creatura invisibilis in conspectu eius omnia autem nuda et aperta sunt oculis eius ad quem nobis sermo
HEB|4|14|habentes ergo pontificem magnum qui penetraverit caelos Iesum Filium Dei teneamus confessionem
HEB|4|15|non enim habemus pontificem qui non possit conpati infirmitatibus nostris temptatum autem per omnia pro similitudine absque peccato
HEB|4|16|adeamus ergo cum fiducia ad thronum gratiae ut misericordiam consequamur et gratiam inveniamus in auxilio oportuno
HEB|5|1|omnis namque pontifex ex hominibus adsumptus pro hominibus constituitur in his quae sunt ad Deum ut offerat dona et sacrificia pro peccatis
HEB|5|2|qui condolere possit his qui ignorant et errant quoniam et ipse circumdatus est infirmitate
HEB|5|3|et propter eam debet quemadmodum et pro populo ita etiam pro semet ipso offerre pro peccatis
HEB|5|4|nec quisquam sumit sibi honorem sed qui vocatur a Deo tamquam Aaron
HEB|5|5|sic et Christus non semet ipsum clarificavit ut pontifex fieret sed qui locutus est ad eum Filius meus es tu ego hodie genui te
HEB|5|6|quemadmodum et in alio dicit tu es sacerdos in aeternum secundum ordinem Melchisedech
HEB|5|7|qui in diebus carnis suae preces supplicationesque ad eum qui possit salvum illum a morte facere cum clamore valido et lacrimis offerens et exauditus pro sua reverentia
HEB|5|8|et quidem cum esset Filius didicit ex his quae passus est oboedientiam
HEB|5|9|et consummatus factus est omnibus obtemperantibus sibi causa salutis aeternae
HEB|5|10|appellatus a Deo pontifex iuxta ordinem Melchisedech
HEB|5|11|de quo grandis nobis sermo et ininterpretabilis ad dicendum quoniam inbecilles facti estis ad audiendum
HEB|5|12|etenim cum deberetis magistri esse propter tempus rursum indigetis ut vos doceamini quae sint elementa exordii sermonum Dei et facti estis quibus lacte opus sit non solido cibo
HEB|5|13|omnis enim qui lactis est particeps expers est sermonis iustitiae parvulus enim est
HEB|5|14|perfectorum autem est solidus cibus eorum qui pro consuetudine exercitatos habent sensus ad discretionem boni ac mali
HEB|6|1|quapropter intermittentes inchoationis Christi sermonem ad perfectionem feramur non rursum iacientes fundamentum paenitentiae ab operibus mortuis et fidei ad Deum
HEB|6|2|baptismatum doctrinae inpositionis quoque manuum ac resurrectionis mortuorum et iudicii aeterni
HEB|6|3|et hoc faciemus siquidem permiserit Deus
HEB|6|4|inpossibile est enim eos qui semel sunt inluminati gustaverunt etiam donum caeleste et participes sunt facti Spiritus Sancti
HEB|6|5|gustaverunt nihilominus bonum Dei verbum virtutesque saeculi venturi
HEB|6|6|et prolapsi sunt renovari rursus ad paenitentiam rursum crucifigentes sibimet ipsis Filium Dei et ostentui habentes
HEB|6|7|terra enim saepe venientem super se bibens imbrem et generans herbam oportunam illis a quibus colitur accipit benedictionem a Deo
HEB|6|8|proferens autem spinas ac tribulos reproba est et maledicto proxima cuius consummatio in conbustionem
HEB|6|9|confidimus autem de vobis dilectissimi meliora et viciniora saluti tametsi ita loquimur
HEB|6|10|non enim iniustus Deus ut obliviscatur operis vestri et dilectionis quam ostendistis in nomine ipsius qui ministrastis sanctis et ministratis
HEB|6|11|cupimus autem unumquemque vestrum eandem ostentare sollicitudinem ad expletionem spei usque in finem
HEB|6|12|ut non segnes efficiamini verum imitatores eorum qui fide et patientia hereditabunt promissiones
HEB|6|13|Abrahae namque promittens Deus quoniam neminem habuit per quem iuraret maiorem iuravit per semet ipsum
HEB|6|14|dicens nisi benedicens benedicam te et multiplicans multiplicabo te
HEB|6|15|et sic longanimiter ferens adeptus est repromissionem
HEB|6|16|homines enim per maiorem sui iurant et omnis controversiae eorum finis ad confirmationem est iuramentum
HEB|6|17|in quo abundantius volens Deus ostendere pollicitationis heredibus inmobilitatem consilii sui interposuit iusiurandum
HEB|6|18|ut per duas res inmobiles quibus inpossibile est mentiri Deum fortissimum solacium habeamus qui confugimus ad tenendam propositam spem
HEB|6|19|quam sicut anchoram habemus animae tutam ac firmam et incedentem usque in interiora velaminis
HEB|6|20|ubi praecursor pro nobis introiit Iesus secundum ordinem Melchisedech pontifex factus in aeternum
HEB|7|1|hic enim Melchisedech rex Salem sacerdos Dei summi qui obviavit Abrahae regresso a caede regum et benedixit ei
HEB|7|2|cui decimas omnium divisit Abraham primum quidem qui interpretatur rex iustitiae deinde autem et rex Salem quod est rex pacis
HEB|7|3|sine patre sine matre sine genealogia neque initium dierum neque finem vitae habens adsimilatus autem Filio Dei manet sacerdos in perpetuum
HEB|7|4|intuemini autem quantus sit hic cui et decimam dedit de praecipuis Abraham patriarcha
HEB|7|5|et quidem de filiis Levi sacerdotium accipientes mandatum habent decimas sumere a populo secundum legem id est a fratribus suis quamquam et ipsi exierunt de lumbis Abrahae
HEB|7|6|cuius autem generatio non adnumeratur in eis decimas sumpsit Abraham et hunc qui habebat repromissiones benedixit
HEB|7|7|sine ulla autem contradictione quod minus est a meliore benedicitur
HEB|7|8|et hic quidem decimas morientes homines accipiunt ibi autem contestatus quia vivit
HEB|7|9|et ut ita dictum sit per Abraham et Levi qui decimas accipit decimatus est
HEB|7|10|adhuc enim in lumbis patris erat quando obviavit ei Melchisedech
HEB|7|11|si ergo consummatio per sacerdotium leviticum erat populus enim sub ipso legem accepit quid adhuc necessarium secundum ordinem Melchisedech alium surgere sacerdotem et non secundum ordinem Aaron dici
HEB|7|12|translato enim sacerdotio necesse est ut et legis translatio fiat
HEB|7|13|in quo enim haec dicuntur de alia tribu est de qua nullus altario praesto fuit
HEB|7|14|manifestum enim quod ex Iuda ortus sit Dominus noster in qua tribu nihil de sacerdotibus Moses locutus est
HEB|7|15|et amplius adhuc manifestum est si secundum similitudinem Melchisedech exsurgit alius sacerdos
HEB|7|16|qui non secundum legem mandati carnalis factus est sed secundum virtutem vitae insolubilis
HEB|7|17|contestatur enim quoniam tu es sacerdos in aeternum secundum ordinem Melchisedech
HEB|7|18|reprobatio quidem fit praecedentis mandati propter infirmitatem eius et inutilitatem
HEB|7|19|nihil enim ad perfectum adduxit lex introductio vero melioris spei per quam proximamus ad Deum
HEB|7|20|et quantum est non sine iureiurando alii quidem sine iureiurando sacerdotes facti sunt
HEB|7|21|hic autem cum iureiurando per eum qui dixit ad illum iuravit Dominus et non paenitebit tu es sacerdos in aeternum
HEB|7|22|in tantum melioris testamenti sponsor factus est Iesus
HEB|7|23|et alii quidem plures facti sunt sacerdotes idcirco quod morte prohiberentur permanere
HEB|7|24|hic autem eo quod maneat in aeternum sempiternum habet sacerdotium
HEB|7|25|unde et salvare in perpetuo potest accedentes per semet ipsum ad Deum semper vivens ad interpellandum pro eis
HEB|7|26|talis enim decebat ut nobis esset pontifex sanctus innocens inpollutus segregatus a peccatoribus et excelsior caelis factus
HEB|7|27|qui non habet cotidie necessitatem quemadmodum sacerdotes prius pro suis delictis hostias offerre deinde pro populi hoc enim fecit semel se offerendo
HEB|7|28|lex enim homines constituit sacerdotes infirmitatem habentes sermo autem iurisiurandi qui post legem est Filium in aeternum perfectum
HEB|8|1|capitulum autem super ea quae dicuntur talem habemus pontificem qui consedit in dextera sedis Magnitudinis in caelis
HEB|8|2|sanctorum minister et tabernaculi veri quod fixit Dominus et non homo
HEB|8|3|omnis enim pontifex ad offerenda munera et hostias constituitur unde necesse est et hunc habere aliquid quod offerat
HEB|8|4|si ergo esset super terram nec esset sacerdos cum essent qui offerrent secundum legem munera
HEB|8|5|qui exemplari et umbrae deserviunt caelestium sicut responsum est Mosi cum consummaret tabernaculum vide inquit omnia facito secundum exemplar quod tibi ostensum est in monte
HEB|8|6|nunc autem melius sortitus est ministerium quanto et melioris testamenti mediator est quod in melioribus repromissionibus sanctum est
HEB|8|7|nam si illud prius culpa vacasset non utique secundi locus inquireretur
HEB|8|8|vituperans enim eos dicit ecce dies veniunt dicit Dominus et consummabo super domum Israhel et super domum Iuda testamentum novum
HEB|8|9|non secundum testamentum quod feci patribus eorum in die qua adprehendi manum illorum ut educerem illos de terra Aegypti quoniam ipsi non permanserunt in testamento meo et ego neglexi eos dicit Dominus
HEB|8|10|quia hoc testamentum quod disponam domui Israhel post dies illos dicit Dominus dando leges meas in mentem eorum et in corde eorum superscribam eas et ero eis in Deum et ipsi erunt mihi in populum
HEB|8|11|et non docebit unusquisque proximum suum et unusquisque fratrem suum dicens cognosce Dominum quoniam omnes scient me a minore usque ad maiorem eorum
HEB|8|12|quia propitius ero iniquitatibus eorum et peccatorum illorum iam non memorabor
HEB|8|13|dicendo autem novum veteravit prius quod autem antiquatur et senescit prope interitum est
HEB|9|1|habuit quidem et prius iustificationes culturae et sanctum saeculare
HEB|9|2|tabernaculum enim factum est primum in quo inerant candelabra et mensa et propositio panum quae dicitur sancta
HEB|9|3|post velamentum autem secundum tabernaculum quod dicitur sancta sanctorum
HEB|9|4|aureum habens turibulum et arcam testamenti circumtectam ex omni parte auro in qua urna aurea habens manna et virga Aaron quae fronduerat et tabulae testamenti
HEB|9|5|superque eam cherubin gloriae obumbrantia propitiatorium de quibus non est modo dicendum per singula
HEB|9|6|his vero ita conpositis in priori quidem tabernaculo semper introibant sacerdotes sacrificiorum officia consummantes
HEB|9|7|in secundo autem semel in anno solus pontifex non sine sanguine quem offert pro sua et populi ignorantia
HEB|9|8|hoc significante Spiritu Sancto nondum propalatam esse sanctorum viam adhuc priore tabernaculo habente statum
HEB|9|9|quae parabola est temporis instantis iuxta quam munera et hostiae offeruntur quae non possunt iuxta conscientiam perfectum facere servientem
HEB|9|10|solummodo in cibis et in potibus et variis baptismis et iustitiis carnis usque ad tempus correctionis inpositis
HEB|9|11|Christus autem adsistens pontifex futurorum bonorum per amplius et perfectius tabernaculum non manufactum id est non huius creationis
HEB|9|12|neque per sanguinem hircorum et vitulorum sed per proprium sanguinem introivit semel in sancta aeterna redemptione inventa
HEB|9|13|si enim sanguis hircorum et taurorum et cinis vitulae aspersus inquinatos sanctificat ad emundationem carnis
HEB|9|14|quanto magis sanguis Christi qui per Spiritum Sanctum semet ipsum obtulit inmaculatum Deo emundabit conscientiam vestram ab operibus mortuis ad serviendum Deo viventi
HEB|9|15|et ideo novi testamenti mediator est ut morte intercedente in redemptionem earum praevaricationum quae erant sub priore testamento repromissionem accipiant qui vocati sunt aeternae hereditatis
HEB|9|16|ubi enim testamentum mors necesse est intercedat testatoris
HEB|9|17|testamentum enim in mortuis confirmatum est alioquin nondum valet dum vivit qui testatus est
HEB|9|18|unde ne primum quidem sine sanguine dedicatum est
HEB|9|19|lecto enim omni mandato legis a Mose universo populo accipiens sanguinem vitulorum et hircorum cum aqua et lana coccinea et hysopo ipsum quoque librum et omnem populum aspersit
HEB|9|20|dicens hic sanguis testamenti quod mandavit ad vos Deus
HEB|9|21|etiam tabernaculum et omnia vasa ministerii sanguine similiter aspersit
HEB|9|22|et omnia paene in sanguine mundantur secundum legem et sine sanguinis fusione non fit remissio
HEB|9|23|necesse est ergo exemplaria quidem caelestium his mundari ipsa autem caelestia melioribus hostiis quam istis
HEB|9|24|non enim in manufactis sanctis Iesus introiit exemplaria verorum sed in ipsum caelum ut appareat nunc vultui Dei pro nobis
HEB|9|25|neque ut saepe offerat semet ipsum quemadmodum pontifex intrat in sancta per singulos annos in sanguine alieno
HEB|9|26|alioquin oportebat eum frequenter pati ab origine mundi nunc autem semel in consummatione saeculorum ad destitutionem peccati per hostiam suam apparuit
HEB|9|27|et quemadmodum statutum est hominibus semel mori post hoc autem iudicium
HEB|9|28|sic et Christus semel oblatus ad multorum exhaurienda peccata secundo sine peccato apparebit expectantibus se in salutem
HEB|10|1|umbram enim habens lex bonorum futurorum non ipsam imaginem rerum per singulos annos hisdem ipsis hostiis quas offerunt indesinenter numquam potest accedentes perfectos facere
HEB|10|2|alioquin non cessassent offerri ideo quod nullam haberent ultra conscientiam peccati cultores semel mundati
HEB|10|3|sed in ipsis commemoratio peccatorum per singulos annos fit
HEB|10|4|inpossibile enim est sanguine taurorum et hircorum auferri peccata
HEB|10|5|ideo ingrediens mundum dicit hostiam et oblationem noluisti corpus autem aptasti mihi
HEB|10|6|holocaustomata et pro peccato non tibi placuit
HEB|10|7|tunc dixi ecce venio in capitulo libri scriptum est de me ut faciam Deus voluntatem tuam
HEB|10|8|superius dicens quia hostias et oblationes et holocaustomata et pro peccato noluisti nec placita sunt tibi quae secundum legem offeruntur
HEB|10|9|tunc dixit ecce venio ut faciam Deus voluntatem tuam aufert primum ut sequens statuat
HEB|10|10|in qua voluntate sanctificati sumus per oblationem corporis Christi Iesu in semel
HEB|10|11|et omnis quidem sacerdos praesto est cotidie ministrans et easdem saepe offerens hostias quae numquam possunt auferre peccata
HEB|10|12|hic autem unam pro peccatis offerens hostiam in sempiternum sedit in dextera Dei
HEB|10|13|de cetero expectans donec ponantur inimici eius scabillum pedum eius
HEB|10|14|una enim oblatione consummavit in sempiternum sanctificatos
HEB|10|15|contestatur autem nos et Spiritus Sanctus postquam enim dixit
HEB|10|16|hoc autem testamentum quod testabor ad illos post dies illos dicit Dominus dando leges meas in cordibus eorum et in mente eorum superscribam eas
HEB|10|17|et peccatorum et iniquitatium eorum iam non recordabor amplius
HEB|10|18|ubi autem horum remissio iam non oblatio pro peccato
HEB|10|19|habentes itaque fratres fiduciam in introitu sanctorum in sanguine Christi
HEB|10|20|quam initiavit nobis viam novam et viventem per velamen id est carnem suam
HEB|10|21|et sacerdotem magnum super domum Dei
HEB|10|22|accedamus cum vero corde in plenitudine fidei aspersi corda a conscientia mala et abluti corpus aqua munda
HEB|10|23|teneamus spei nostrae confessionem indeclinabilem fidelis enim est qui repromisit
HEB|10|24|et consideremus invicem in provocationem caritatis et bonorum operum
HEB|10|25|non deserentes collectionem nostram sicut est consuetudinis quibusdam sed consolantes et tanto magis quanto videritis adpropinquantem diem
HEB|10|26|voluntarie enim peccantibus nobis post acceptam notitiam veritatis iam non relinquitur pro peccatis hostia
HEB|10|27|terribilis autem quaedam expectatio iudicii et ignis aemulatio quae consumptura est adversarios
HEB|10|28|irritam quis faciens legem Mosi sine ulla miseratione duobus vel tribus testibus moritur
HEB|10|29|quanto magis putatis deteriora mereri supplicia qui Filium Dei conculcaverit et sanguinem testamenti pollutum duxerit in quo sanctificatus est et Spiritui gratiae contumeliam fecerit
HEB|10|30|scimus enim qui dixit mihi vindictam ego reddam et iterum quia iudicabit Dominus populum suum
HEB|10|31|horrendum est incidere in manus Dei viventis
HEB|10|32|rememoramini autem pristinos dies in quibus inluminati magnum certamen sustinuistis passionum
HEB|10|33|et in altero quidem obprobriis et tribulationibus spectaculum facti in altero autem socii taliter conversantium effecti
HEB|10|34|nam et vinctis conpassi estis et rapinam bonorum vestrorum cum gaudio suscepistis cognoscentes vos habere meliorem et manentem substantiam
HEB|10|35|nolite itaque amittere confidentiam vestram quae magnam habet remunerationem
HEB|10|36|patientia enim vobis necessaria est ut voluntatem Dei facientes reportetis promissionem
HEB|10|37|adhuc enim modicum quantulum qui venturus est veniet et non tardabit
HEB|10|38|iustus autem meus ex fide vivit quod si subtraxerit se non placebit animae meae
HEB|10|39|nos autem non sumus subtractionis in perditionem sed fidei in adquisitionem animae
HEB|11|1|est autem fides sperandorum substantia rerum argumentum non parentum
HEB|11|2|in hac enim testimonium consecuti sunt senes
HEB|11|3|fide intellegimus aptata esse saecula verbo Dei ut ex invisibilibus visibilia fierent
HEB|11|4|fide plurimam hostiam Abel quam Cain obtulit Deo per quam testimonium consecutus est esse iustus testimonium perhibente muneribus eius Deo et per illam defunctus adhuc loquitur
HEB|11|5|fide Enoch translatus est ne videret mortem et non inveniebatur quia transtulit illum Deus ante translationem enim testimonium habebat placuisse Deo
HEB|11|6|sine fide autem inpossibile placere credere enim oportet accedentem ad Deum quia est et inquirentibus se remunerator fit
HEB|11|7|fide Noe responso accepto de his quae adhuc non videbantur metuens aptavit arcam in salutem domus suae per quam damnavit mundum et iustitiae quae per fidem est heres est institutus
HEB|11|8|fide qui vocatur Abraham oboedivit in locum exire quem accepturus erat in hereditatem et exiit nesciens quo iret
HEB|11|9|fide moratus est in terra repromissionis tamquam in aliena in casulis habitando cum Isaac et Iacob coheredibus repromissionis eiusdem
HEB|11|10|expectabat enim fundamenta habentem civitatem cuius artifex et conditor Deus
HEB|11|11|fide et ipsa Sarra sterilis virtutem in conceptionem seminis accepit etiam praeter tempus aetatis quoniam fidelem credidit esse qui promiserat
HEB|11|12|propter quod et ab uno orti sunt et haec emortuo tamquam sidera caeli in multitudinem et sicut harena quae est ad oram maris innumerabilis
HEB|11|13|iuxta fidem defuncti sunt omnes isti non acceptis repromissionibus sed a longe eas aspicientes et salutantes et confitentes quia peregrini et hospites sunt supra terram
HEB|11|14|qui enim haec dicunt significant se patriam inquirere
HEB|11|15|et si quidem illius meminissent de qua exierunt habebant utique tempus revertendi
HEB|11|16|nunc autem meliorem appetunt id est caelestem ideo non confunditur Deus vocari Deus eorum paravit enim illis civitatem
HEB|11|17|fide obtulit Abraham Isaac cum temptaretur et unigenitum offerebat qui susceperat repromissiones
HEB|11|18|ad quem dictum est quia in Isaac vocabitur tibi semen
HEB|11|19|arbitrans quia et a mortuis suscitare potens est Deus unde eum et in parabola accepit
HEB|11|20|fide et de futuris benedixit Isaac Iacob et Esau
HEB|11|21|fide Iacob moriens singulis filiorum Ioseph benedixit et adoravit fastigium virgae eius
HEB|11|22|fide Ioseph moriens de profectione filiorum Israhel memoratus est et de ossibus suis mandavit
HEB|11|23|fide Moses natus occultatus est mensibus tribus a parentibus suis eo quod vidissent elegantem infantem et non timuerunt regis edictum
HEB|11|24|fide Moses grandis factus negavit se esse filium filiae Pharaonis
HEB|11|25|magis eligens adfligi cum populo Dei quam temporalis peccati habere iucunditatem
HEB|11|26|maiores divitias aestimans thesauro Aegyptiorum inproperium Christi aspiciebat enim in remunerationem
HEB|11|27|fide reliquit Aegyptum non veritus animositatem regis invisibilem enim tamquam videns sustinuit
HEB|11|28|fide celebravit pascha et sanguinis effusionem ne qui vastabat primitiva tangeret eos
HEB|11|29|fide transierunt mare Rubrum tamquam per aridam terram quod experti Aegyptii devorati sunt
HEB|11|30|fide muri Hiericho ruerunt circuiti dierum septem
HEB|11|31|fide Raab meretrix non periit cum incredulis excipiens exploratores cum pace
HEB|11|32|et quid adhuc dicam deficiet enim me tempus enarrantem de Gedeon Barac Samson Iepthae David et Samuhel et prophetis
HEB|11|33|qui per fidem devicerunt regna operati sunt iustitiam adepti sunt repromissiones obturaverunt ora leonum
HEB|11|34|extinxerunt impetum ignis effugerunt aciem gladii convaluerunt de infirmitate fortes facti sunt in bello castra verterunt exterorum
HEB|11|35|acceperunt mulieres de resurrectione mortuos suos alii autem distenti sunt non suscipientes redemptionem ut meliorem invenirent resurrectionem
HEB|11|36|alii vero ludibria et verbera experti insuper et vincula et carceres
HEB|11|37|lapidati sunt secti sunt temptati sunt in occisione gladii mortui sunt circumierunt in melotis in pellibus caprinis egentes angustiati adflicti
HEB|11|38|quibus dignus non erat mundus in solitudinibus errantes et montibus et speluncis et in cavernis terrae
HEB|11|39|et hii omnes testimonio fidei probati non acceperunt repromissionem
HEB|11|40|Deo pro nobis melius aliquid providente ut ne sine nobis consummarentur
HEB|12|1|ideoque et nos tantam habentes inpositam nubem testium deponentes omne pondus et circumstans nos peccatum per patientiam curramus propositum nobis certamen
HEB|12|2|aspicientes in auctorem fidei et consummatorem Iesum qui pro proposito sibi gaudio sustinuit crucem confusione contempta atque in dextera sedis Dei sedit
HEB|12|3|recogitate enim eum qui talem sustinuit a peccatoribus adversum semet ipsos contradictionem ut ne fatigemini animis vestris deficientes
HEB|12|4|nondum usque ad sanguinem restitistis adversus peccatum repugnantes
HEB|12|5|et obliti estis consolationis quae vobis tamquam filiis loquitur dicens fili mi noli neglegere disciplinam Domini neque fatigeris dum ab eo argueris
HEB|12|6|quem enim diligit Dominus castigat flagellat autem omnem filium quem recipit
HEB|12|7|in disciplina perseverate tamquam filiis vobis offert Deus quis enim filius quem non corripit pater
HEB|12|8|quod si extra disciplinam estis cuius participes facti sunt omnes ergo adulteri et non filii estis
HEB|12|9|deinde patres quidem carnis nostrae habuimus eruditores et reverebamur non multo magis obtemperabimus Patri spirituum et vivemus
HEB|12|10|et illi quidem in tempore paucorum dierum secundum voluntatem suam erudiebant nos hic autem ad id quod utile est in recipiendo sanctificationem eius
HEB|12|11|omnis autem disciplina in praesenti quidem videtur non esse gaudii sed maeroris postea autem fructum pacatissimum exercitatis per eam reddit iustitiae
HEB|12|12|propter quod remissas manus et soluta genua erigite
HEB|12|13|et gressus rectos facite pedibus vestris ut non claudicans erret magis autem sanetur
HEB|12|14|pacem sequimini cum omnibus et sanctimoniam sine qua nemo videbit Dominum
HEB|12|15|contemplantes ne quis desit gratiae Dei ne qua radix amaritudinis sursum germinans inpediat et per illam inquinentur multi
HEB|12|16|ne quis fornicator aut profanus ut Esau qui propter unam escam vendidit primitiva sua
HEB|12|17|scitote enim quoniam et postea cupiens hereditare benedictionem reprobatus est non enim invenit paenitentiae locum quamquam cum lacrimis inquisisset eam
HEB|12|18|non enim accessistis ad tractabilem et accensibilem ignem et turbinem et caliginem et procellam
HEB|12|19|et tubae sonum et vocem verborum quam qui audierunt excusaverunt se ne eis fieret verbum
HEB|12|20|non enim portabant quod dicebatur et si bestia tetigerit montem lapidabitur
HEB|12|21|et ita terribile erat quod videbatur Moses dixit exterritus sum et tremebundus
HEB|12|22|sed accessistis ad Sion montem et civitatem Dei viventis Hierusalem caelestem et multorum milium angelorum frequentiae
HEB|12|23|et ecclesiam primitivorum qui conscripti sunt in caelis et iudicem omnium Deum et spiritus iustorum perfectorum
HEB|12|24|et testamenti novi mediatorem Iesum et sanguinis sparsionem melius loquentem quam Abel
HEB|12|25|videte ne recusetis loquentem si enim illi non effugerunt recusantes eum qui super terram loquebatur multo magis nos qui de caelis loquentem nobis avertimur
HEB|12|26|cuius vox movit terram tunc modo autem repromittit dicens adhuc semel ego movebo non solum terram sed et caelum
HEB|12|27|quod autem adhuc semel dicit declarat mobilium translationem tamquam factorum ut maneant ea quae sunt inmobilia
HEB|12|28|itaque regnum inmobile suscipientes habemus gratiam per quam serviamus placentes Deo cum metu et reverentia
HEB|12|29|etenim Deus noster ignis consumens est
HEB|13|1|caritas fraternitatis maneat
HEB|13|2|hospitalitatem nolite oblivisci per hanc enim latuerunt quidam angelis hospitio receptis
HEB|13|3|mementote vinctorum tamquam simul vincti et laborantium tamquam et ipsi in corpore morantes
HEB|13|4|honorabile conubium in omnibus et torus inmaculatus fornicatores enim et adulteros iudicabit Deus
HEB|13|5|sint mores sine avaritia contenti praesentibus ipse enim dixit non te deseram neque derelinquam
HEB|13|6|ita ut confidenter dicamus Dominus mihi adiutor non timebo quid faciat mihi homo
HEB|13|7|mementote praepositorum vestrorum qui vobis locuti sunt verbum Dei quorum intuentes exitum conversationis imitamini fidem
HEB|13|8|Iesus Christus heri et hodie ipse et in saecula
HEB|13|9|doctrinis variis et peregrinis nolite abduci optimum enim est gratia stabiliri cor non escis quae non profuerunt ambulantibus in eis
HEB|13|10|habemus altare de quo edere non habent potestatem qui tabernaculo deserviunt
HEB|13|11|quorum enim animalium infertur sanguis pro peccato in sancta per pontificem horum corpora cremantur extra castra
HEB|13|12|propter quod et Iesus ut sanctificaret per suum sanguinem populum extra portam passus est
HEB|13|13|exeamus igitur ad eum extra castra inproperium eius portantes
HEB|13|14|non enim habemus hic manentem civitatem sed futuram inquirimus
HEB|13|15|per ipsum ergo offeramus hostiam laudis semper Deo id est fructum labiorum confitentium nomini eius
HEB|13|16|beneficientiae autem et communionis nolite oblivisci talibus enim hostiis promeretur Deus
HEB|13|17|oboedite praepositis vestris et subiacete eis ipsi enim pervigilant quasi rationem pro animabus vestris reddituri ut cum gaudio hoc faciant et non gementes hoc enim non expedit vobis
HEB|13|18|orate pro nobis confidimus enim quia bonam conscientiam habemus in omnibus bene volentes conversari
HEB|13|19|amplius autem deprecor vos hoc facere ut quo celerius restituar vobis
HEB|13|20|Deus autem pacis qui eduxit de mortuis pastorem magnum ovium in sanguine testamenti aeterni Dominum nostrum Iesum
HEB|13|21|aptet vos in omni bono ut faciatis voluntatem eius faciens in vobis quod placeat coram se per Iesum Christum cui gloria in saecula saeculorum amen
HEB|13|22|rogo autem vos fratres sufferatis verbum solacii etenim perpaucis scripsi vobis
HEB|13|23|cognoscite fratrem nostrum Timotheum dimissum cum quo si celerius venerit videbo vos
HEB|13|24|salutate omnes praepositos vestros et omnes sanctos salutant vos de Italia
HEB|13|25|gratia cum omnibus vobis amen
