JER|1|1|這些是 便雅憫 地 亞拿突城 的祭司， 希勒家 的兒子 耶利米 的話。
JER|1|2|亞們 的兒子 猶大 王 約西亞 在位第十三年，耶和華的話臨到 耶利米 。
JER|1|3|從 約西亞 的兒子 猶大 王 約雅敬 在位的時候，直到 約西亞 的兒子 猶大 王 西底家 在位的末年，就是第十一年五月間 耶路撒冷 被擄時，耶和華的話也常臨到 耶利米 。
JER|1|4|耶利米 說，耶和華的話臨到我，說：
JER|1|5|「我尚未將你造在母腹中，就已認識你； 你未出母胎，我已將你分別為聖， 派你作列國的先知。」
JER|1|6|我就說：「唉，主耶和華！看哪，我不知道怎麼說，因為我年輕。」
JER|1|7|耶和華對我說： 「不要說：『我年輕』， 因為我差遣你到誰那裏去，你都要去； 我吩咐你說甚麼話，你都要說。
JER|1|8|你不要怕他們， 因為我與你同在，要拯救你。 這是耶和華說的。」
JER|1|9|於是耶和華伸手按住我的口， 對我說： 「看哪，我已將我的話放在你口中。
JER|1|10|我今日立你在列邦列國之上， 為要拔出，拆毀，毀壞，傾覆， 又要建立，栽植。」
JER|1|11|耶和華的話臨到我，說：「 耶利米 ，你看見甚麼？」我說：「我看見一根杏樹枝。」
JER|1|12|耶和華對我說：「你看得不錯；因為我要看守 我的話，使它實現。」
JER|1|13|耶和華的話第二次臨到我，說：「你看見甚麼？」我說：「我看見一個水燒開的鍋，從北而傾。」
JER|1|14|耶和華對我說：「必有災禍從北方發出，臨到這地所有的居民。
JER|1|15|看哪，我要召北方列國的萬族。這是耶和華說的。他們要來，各安寶座在 耶路撒冷 的城門口，周圍攻擊城牆，又要攻擊 猶大 的一切城鎮。
JER|1|16|這百姓離棄我，向別神燒香，跪拜自己手所造的，我要針對這一切惡行，向他們宣讀我的判決。
JER|1|17|所以你當束腰，起來，將我所吩咐你的一切話都告訴他們；不要因他們驚惶，免得我使你在他們面前驚惶。
JER|1|18|看哪，我今日使你成為堅城、鐵柱、銅牆，對抗全地和 猶大 的君王、官長、祭司，並這地的百姓。
JER|1|19|他們要攻擊你，卻不能勝過你，因為我與你同在，要拯救你。這是耶和華說的。」
JER|2|1|耶和華的話臨到我，說：
JER|2|2|「你去向 耶路撒冷 居民的耳朵呼喊說，耶和華如此說： 『你年輕時的恩愛， 新婚時的愛情， 你怎樣在曠野， 在未耕種之地跟隨我， 我都記得。
JER|2|3|那時 以色列 歸耶和華為聖， 作為他初熟的土產； 凡吞吃它的必算為有罪， 災禍必臨到他們。 這是耶和華說的。』」
JER|2|4|雅各 家， 以色列 家的各族啊，當聽耶和華的話，
JER|2|5|耶和華如此說： 「你們的祖先看我有甚麼錯處， 竟遠離我，隨從那虛無的神明 ， 自己成為虛無呢？
JER|2|6|他們並不問： 『那領我們從 埃及 地上來， 引導我們走過曠野、沙漠有坑洞之地， 走過乾旱死蔭、無人經過、 無人居住之地的耶和華在哪裏呢？』
JER|2|7|我領你們進入肥沃之地， 使你們得吃其中的果子和美物； 你們進入時，卻使我的地玷污， 使我的產業成為可憎惡的。
JER|2|8|祭司從來不問：『耶和華在哪裏呢？』 傳講律法的不認識我， 官長違背我， 先知藉 巴力 說預言， 隨從無益的東西。」
JER|2|9|「我因此必與你們爭辯， 也與你們的子孫爭辯。 這是耶和華說的。
JER|2|10|你們且渡到 基提 海島察看， 派人往 基達 去留心查考， 看可曾有過這樣的事。
JER|2|11|豈有一國換了它的神明嗎？ 其實那不是神明！ 但我的百姓將他們的榮耀換了那無益的東西。
JER|2|12|諸天哪，要因此震驚， 顫慄，極其淒涼！ 這是耶和華說的。
JER|2|13|因為我的百姓做了兩件惡事： 離棄我這活水的泉源； 又為自己鑿出水池， 卻是破裂不能儲水的池子。」
JER|2|14|「 以色列 是僕人嗎？ 是家中生的奴僕嗎？ 為何成為掠物呢？
JER|2|15|少壯獅子向它咆哮，大聲吼叫， 使它的地荒蕪； 城鎮燒燬，無人居住。
JER|2|16|挪弗 人和 答比匿 人打破你的頭顱。
JER|2|17|這不是你自己招惹的嗎？ 不是因耶和華－你上帝引導你行路時， 你離棄了他嗎？
JER|2|18|現今你為何在 埃及 路上喝 西曷河 的水呢？ 為何在 亞述 路上喝 大河 的水呢？
JER|2|19|你自己的惡必懲治你， 你背道的事必責罰你。 由此可知可見，你離棄耶和華－你的上帝， 不存敬畏我的心， 實為惡事，為苦事； 這是萬軍之主耶和華說的。」
JER|2|20|「你 在古時折斷你的軛，解開你的繩索， 說：『我必不事奉耶和華 。』 你在各高岡上、各青翠的樹下屈身行淫。
JER|2|21|然而，我栽種你為上等的葡萄樹， 全用純正的種子； 你怎麼向我變為外邦葡萄樹的壞枝子呢？
JER|2|22|你雖用鹼、多用皂莢清洗， 你罪孽的痕跡仍顯在我面前。 這是主耶和華說的。
JER|2|23|你怎能說： 『我沒有玷污，沒有隨從 巴力 』？ 看看你在谷中所做的，思想你自己的所作所為； 你是快行的獨峰駝，狂奔亂闖。
JER|2|24|你是野驢，習慣曠野， 慾心發動時就呼吸急促， 發情時誰能使牠轉回呢？ 凡尋找牠的必不費力， 在牠的季節必能尋見牠。
JER|2|25|你不要弄到赤足而行， 喉嚨乾渴。 你卻說：『沒有用的， 我喜愛陌生人， 我必隨從他們。』」
JER|2|26|「賊被捉拿，怎樣羞愧， 以色列 家和他們的君王、官長、 祭司、先知也都照樣羞愧。
JER|2|27|他們向木頭說：『你是我的父』； 向石頭說：『你是生我的。』 他們以背向我， 不肯以面向我； 及至遭遇患難時卻說： 『起來拯救我們吧！』
JER|2|28|你為自己做的神明在哪裏呢？ 你遭遇患難的時候， 讓它們起來拯救你吧！ 猶大 啊，你神明的數目與你城的數目相等。
JER|2|29|「你們為何與我爭辯呢？ 你們都違背了我。 這是耶和華說的。
JER|2|30|我責打你們的兒女是徒然的， 他們不受管教。 你們自己的刀吞滅你們的先知， 好像殘害人的獅子。
JER|2|31|這世代的人哪， 你們要留意耶和華的話。 我向 以色列 豈是曠野， 或幽暗之地呢？ 我的百姓為何說： 『我們脫離約束，不再歸向你了』？
JER|2|32|少女豈能忘記她的妝飾呢？ 新娘豈能忘記她的美衣呢？ 我的百姓卻在無數的日子裏忘記了我！
JER|2|33|「你竟然如此精於求愛之道， 可把你的門徑教邪惡的女人！
JER|2|34|你衣服的邊上有無辜貧窮人的血， 其實你並未發現他們挖洞進屋偷竊 。 雖有這一切的事 ，
JER|2|35|你還說：『我無辜； 耶和華的怒氣必定轉離我了。』 看哪，我必審問你； 因你自己說：『我沒有犯罪。』
JER|2|36|你為何東奔西跑改變你的道路呢？ 你必因 埃及 蒙羞， 像從前因 亞述 蒙羞一樣。
JER|2|37|你也必兩手抱頭離開這裏； 因為耶和華已經棄絕你所倚靠的， 你不能因他們而得順利。」
JER|3|1|耶和華說 ：「人若休妻， 妻離他而去，做了別人的妻子， 前夫豈能再回到她那裏呢？ 那地豈不是大大污穢了嗎？ 但你和許多情郎行淫， 還是可以回到我這裏。 這是耶和華說的。
JER|3|2|你舉目向光禿的高地觀看， 何處沒有你的淫行呢？ 你坐在道路旁等候， 好像 阿拉伯 人在曠野埋伏， 你的淫行和邪惡使全地污穢了。
JER|3|3|因此甘霖停止， 春雨不降。 你還是一副娼妓之臉， 不顧羞恥。
JER|3|4|你不是才向我呼叫說： 『我父啊，你是我年輕時的密友，
JER|3|5|人豈永遠懷恨，長久存怒嗎？』 看哪，你雖這樣說，還是竭盡所能去行惡。」
JER|3|6|約西亞 王在位的時候，耶和華對我說：「你看見背道的 以色列 所做的嗎？她上到各高山，在各青翠的樹下行淫。
JER|3|7|我說：『她行這些事以後會回轉歸向我』，她卻不回轉。她奸詐的妹妹 猶大 也看見了。
JER|3|8|我看見背道的 以色列 行淫，我為這緣故給她休書休了她，她奸詐的妹妹 猶大 還不懼怕，也去行淫。
JER|3|9|因 以色列 輕忽了她的淫亂，與石頭和木頭行姦淫 ，她和這地就都污穢了 。
JER|3|10|雖有這一切的事，她奸詐的妹妹 猶大 還不一心歸向我，不過是假意歸我。這是耶和華說的。」
JER|3|11|耶和華對我說：「背道的 以色列 比奸詐的 猶大 還顯為義。
JER|3|12|你去向北方宣告這些話，說： 『背道的 以色列 啊，回來吧！ 這是耶和華說的。 我必不怒目看你們， 因為我是慈愛的， 這是耶和華說的。 我必不永遠懷怒；
JER|3|13|只要你承認你的罪孽， 就是違背耶和華－你的上帝， 在各青翠的樹下追逐外族的神明 ， 沒有聽從我的話。 這是耶和華說的。
JER|3|14|背道的兒女啊，回來吧！ 這是耶和華說的。 因為我作你們的丈夫， 要將你們從一城取一人， 從一族取兩人，帶到 錫安 。
JER|3|15|「『我必將合我心意的牧者賞賜給你們，他們要以知識和智慧牧養你們。
JER|3|16|你們在國中生養眾多的時候，那些日子，人必不再提說耶和華的約櫃，不追想，不記念，不覺缺少，也不再製造。這是耶和華說的。
JER|3|17|那時，人必稱 耶路撒冷 為耶和華的寶座；萬國聚集在那裏，為耶和華的名來到 耶路撒冷 ，他們必不再隨從自己頑梗的惡心行事。
JER|3|18|當那些日子， 猶大 家要和 以色列 家同行，從北方之地一同來到我所賜給你們祖先為業之地。』」
JER|3|19|我說，我多麼樂意把你列在兒女之中， 賜給你美地， 就是萬國中最美的產業。 我說，你會以「我父啊」稱呼我， 不再轉離而跟從我。
JER|3|20|以色列 家啊，你們向我行詭詐， 真像妻子行詭詐離開丈夫。 這是耶和華說的。
JER|3|21|有聲音從光禿的高地傳來， 就是 以色列 人哭泣懇求的聲音， 因為他們走彎曲之道， 忘記耶和華－他們的上帝。
JER|3|22|「你們這背道的兒女啊，回來吧！ 我要醫治你們背道的病。」 「看哪，我們來到你這裏， 因你是耶和華－我們的上帝。
JER|3|23|從小山來的真是枉然， 大山的喧嚷也是枉然 。 以色列 得救，誠然在乎耶和華－我們的上帝。
JER|3|24|「從我們幼年以來，那可恥之物 吞吃了我們祖先勞碌得來的，就是他們的羊群、牛群和他們的兒女。
JER|3|25|我們在羞恥中躺臥吧！願慚愧將我們遮蓋！因為從我們幼年以來，我們和我們的祖先都得罪了耶和華－我們的上帝，沒有聽從耶和華－我們上帝的話。」
JER|4|1|耶和華說：「 以色列 啊， 你若回轉，回轉歸向我， 若從我眼前除掉你可憎的偶像， 不再猶疑不定，
JER|4|2|憑誠實、公平、公義 指著永生的耶和華起誓； 列國就必因他蒙福， 也必因他誇耀。」
JER|4|3|耶和華對 猶大 人和 耶路撒冷 人如此說： 「你們要為自己開墾荒地， 不要撒種在荊棘裏。
JER|4|4|猶大 人和 耶路撒冷 的居民哪， 你們當自行割禮，歸耶和華， 將你們心裏的污穢 除掉； 免得我的憤怒因你們的惡行發作， 如火燃起， 甚至無人能熄滅！」
JER|4|5|你們要在 猶大 傳揚， 在 耶路撒冷 宣告，說： 「當在國中吹角，高聲呼叫說： 『你們當聚集！ 我們好進入堅固城！』
JER|4|6|應當向 錫安 豎立大旗。 逃吧，不要遲延， 因我必使災禍與大毀滅從北方來到。
JER|4|7|有獅子從密林中上來， 是毀壞列國的。 牠已動身出離本處， 要使你的地荒涼， 使你的城鎮變為廢墟，無人居住。
JER|4|8|因此，你們當腰束麻布，哭泣哀號， 因為耶和華的烈怒並未轉離我們。」
JER|4|9|耶和華說：「到那時，君王和領袖的心要失喪，祭司都要驚奇，先知都要詫異。」
JER|4|10|我說：「哀哉！主耶和華啊，你真是大大欺哄這百姓和 耶路撒冷 ，說：『你們必得平安。』其實刀劍已經抵住喉嚨了！」
JER|4|11|那時，必有話對這百姓和 耶路撒冷 說：「來自曠野光禿高地的熱風吹向我的百姓 ，不是為簸揚，也不是為揚淨。
JER|4|12|又有一陣比這更大的風向我颳來；現在，我要向他們宣讀我的判決。」
JER|4|13|看哪，他必如雲湧上； 他的戰車如旋風， 他的馬比鷹更快。 我們有禍了！ 我們敗落了！
JER|4|14|耶路撒冷 啊，你當洗去心中的惡， 使你可以得救。 惡念在你裏面要存到幾時呢？
JER|4|15|有聲音從 但 傳出， 有災禍從 以法蓮山 傳來。
JER|4|16|你們當傳給列國， 看哪，要向 耶路撒冷 報告： 「有圍攻的人從遠方來到， 向 猶大 的城鎮大聲喊叫。
JER|4|17|他們包圍 耶路撒冷 ， 好像看守田園的， 因為它背叛了我。 這是耶和華說的。
JER|4|18|你的作風和行為招惹這事； 這是你罪惡的結果， 實在是苦， 刺透了你的心！」
JER|4|19|我的肺腑啊，我的肺腑啊，我心疼痛！ 我的心在我裏面煩躁不安。 我不能靜默不言， 因我已聽見角聲和打仗的喊聲。
JER|4|20|毀壞的信息不斷傳來， 因為全地荒廢。 我的帳棚忽然毀壞， 我的幔子頃刻破裂。
JER|4|21|我看見大旗，聽見角聲， 要到幾時呢？
JER|4|22|「我的百姓愚頑，不認識我； 他們是愚昧無知的兒女， 有智慧行惡，沒有知識行善。」
JER|4|23|我觀看地， 看哪，地是空虛混沌； 我觀看天，天也無光。
JER|4|24|我觀看大山，看哪，盡都震動， 小山也都搖來搖去。
JER|4|25|我觀看，看哪，無人； 空中的飛鳥也都躲避。
JER|4|26|我觀看，看哪，肥田變為荒地； 所有城鎮在耶和華面前， 因他的烈怒都被拆毀。
JER|4|27|耶和華如此說：「全地必然荒涼， 我卻不毀滅淨盡。
JER|4|28|因此，地要悲哀， 天上也必黑暗； 因為我言已出，我意已定， 必不改變，也不由此轉回。」
JER|4|29|各城的人因騎兵和弓箭手的響聲就都逃跑， 進入密林，爬上磐石； 城鎮都被拋棄， 無人住在其中。
JER|4|30|你這被毀滅的啊， 你要做甚麼呢？ 你穿上朱紅衣服， 佩戴黃金飾物， 用眼影修飾眼睛， 徒然美化你自己。 戀慕你的卻藐視你， 尋索你的性命。
JER|4|31|我聽見彷彿婦人臨產的聲音， 好像生頭胎疼痛的聲音， 原來是 錫安 的聲音； 她喘著氣，伸開手： 「我有禍了！ 在殺人者跟前，我的心靈發昏。」
JER|5|1|你們要走遍 耶路撒冷 的街市， 在廣場尋找， 看是否有人行公平、求誠實； 若有，我就赦免這城。
JER|5|2|雖然他們說「我對永生的耶和華發誓」， 所起的誓實在是假的。
JER|5|3|耶和華啊，你的眼目不是在尋找誠實嗎？ 你擊打他們，他們卻不傷慟； 你摧毀他們，他們仍不領受管教。 他們使臉剛硬過於磐石， 不肯回頭。
JER|5|4|我說：「這些人實在是貧寒的， 他們是愚昧的， 因為不知道耶和華的作為， 也不知道他們上帝的法則。
JER|5|5|我要去見尊貴的人，向他們說話， 他們應該知道耶和華的作為， 知道他們上帝的法則。」 然而，這些人卻齊心將軛折斷， 掙開繩索。
JER|5|6|因此，林中的獅子必害死他們， 野地的狼必滅絕他們， 豹子在城外窺伺。 凡出城的必被撕碎， 因為他們的罪過極多， 背道的事也增加。
JER|5|7|我怎能赦免你呢？ 你的兒女離棄我， 又指著那不是上帝的起誓。 我使他們飽足， 他們就行姦淫， 居住 在娼妓家裏。
JER|5|8|他們如餵飽的馬，精力旺盛， 各向鄰舍的妻子吹哨。
JER|5|9|我豈不因這些事施行懲罰嗎？ 像這樣的國家，我豈能不報復呢？ 這是耶和華說的。
JER|5|10|你們要上去毀壞它的葡萄園， 但不可毀壞淨盡， 只可除掉其枝子， 因為不屬耶和華。
JER|5|11|以色列 家和 猶大 家向我大行詭詐。 這是耶和華說的。
JER|5|12|關乎耶和華他們說了虛謊的話： 「他不會的， 災禍必不臨到我們， 我們也不會遇見刀劍和饑荒。
JER|5|13|先知不過是一陣風， 道也不在他們裏面； 這災禍必臨到他們身上。」
JER|5|14|所以耶和華－萬軍之上帝如此說： 「因為他們說這話， 看哪，我必使我的話在你口中為火， 使這百姓為柴， 火便將他們燒滅。
JER|5|15|以色列 家啊， 看哪，我必使一國從遠方來攻擊你， 是強盛的國， 是古老的國； 他們的言語你不知道， 所說的話你不明白。 這是耶和華說的。
JER|5|16|他們的箭袋有如敞開的墳墓， 他們全都是勇士。
JER|5|17|他們必吃盡你的莊稼和糧食， 是你兒女該吃的 ； 必吃盡你的牛羊， 吃盡你的葡萄和無花果； 又必用刀劍毀壞你所倚靠的堅固城。
JER|5|18|「就是在那些日子，我也不會將你們毀滅淨盡。這是耶和華說的。
JER|5|19|百姓若說：『耶和華－我們的上帝為甚麼向我們行這一切事呢？』你就對他們說：『你們怎樣離棄我，在你們的地上事奉外邦神明，也必照樣在不屬你們的地上事奉外族人。』」
JER|5|20|當在 雅各 家傳揚， 在 猶大 宣告，說：
JER|5|21|「愚昧無知的百姓啊， 你們有眼不看， 有耳不聽， 現在當聽這話。
JER|5|22|你們難道不懼怕我嗎？ 在我面前還不戰兢嗎？ 這是耶和華說的。 我以沙為海的界限， 作永遠的條例，使它不得越過。 波浪洶湧，卻不能勝過； 怒濤澎湃，仍無法越過。
JER|5|23|但這百姓有背叛忤逆的心， 他們轉離而去。
JER|5|24|他們心裏並不說： 『我們應當敬畏耶和華－我們的上帝； 他按時賜雨，就是秋雨和春雨， 又為我們定收割的季節。』
JER|5|25|你們的罪孽使這些轉離你們， 你們的罪惡使你們不能得福。
JER|5|26|在我百姓當中有惡人， 他們埋伏，好像捕鳥的人在窺探 ； 他們設羅網陷害人。
JER|5|27|籠子怎樣裝滿雀鳥， 他們的屋裏也照樣充滿詭詐； 他們因此得以強大富足。
JER|5|28|他們肥胖光潤，作惡過甚， 不為人伸冤， 不為孤兒伸冤，使他們勝訴， 也不為貧窮人辯護。
JER|5|29|我豈不因這些事施行懲罰嗎？ 像這樣的國家，我豈能不報復呢？ 這是耶和華說的。
JER|5|30|「國中有令人驚駭、 恐怖的事發生，
JER|5|31|先知說假預言， 祭司把權柄抓在自己手上， 我的百姓也喜愛這樣， 到了結局你們要怎麼辦呢？」
JER|6|1|便雅憫 人哪，當逃離 耶路撒冷 ， 在 提哥亞 吹號角， 在 伯‧哈基琳 升信號， 因為有災禍與大毀滅從北方逼近。
JER|6|2|那秀美嬌嫩的 錫安 ， 我必剪除。
JER|6|3|牧人必引領羊群到它那裏， 在它周圍支搭帳棚， 各在自己的地方放牧。
JER|6|4|「你們要準備攻擊它。 起來吧，我們要趁正午上去。」 「哀哉！日已漸斜， 黃昏的影子拖長了。」
JER|6|5|「起來吧，我們要在夜間上去， 毀壞它的宮殿。」
JER|6|6|萬軍之耶和華如此說： 「你們要砍伐樹木， 建土堆攻打 耶路撒冷 ， 就是那該受罰的城 ， 其中盡是欺壓。
JER|6|7|井怎樣湧出水來， 這城也照樣湧出惡來； 其中常聽聞殘暴毀滅的事， 病痛損傷也常在我面前。
JER|6|8|耶路撒冷 啊，當受管教， 免得我心與你生疏， 免得我使你荒涼， 成為無人居住之地。」
JER|6|9|萬軍之耶和華如此說： 「他們洗劫 以色列 剩下的民， 如摘淨葡萄一樣； 現你的手如採收葡萄的人，在樹枝上採了又採 。」
JER|6|10|現在我可以向誰說話，警告誰，使他們聽呢？ 看哪，他們的耳朵未受割禮，不能聽見。 看哪，他們以耶和華的話為羞辱， 不以為喜悅。
JER|6|11|因此我被耶和華的憤怒充滿，難以忍受。 「你要把它倒在街上孩童 和成群的年輕人身上， 他們連夫帶妻， 年長者與高齡的人都必被擒拿。
JER|6|12|他們的房屋、田地， 和妻子都要一起轉歸別人， 我要伸手攻擊這地的居民。」 這是耶和華說的。
JER|6|13|「因為他們從最小的到最大的都貪圖不義之財， 從先知到祭司全都行事虛假。
JER|6|14|他們輕忽地醫治我百姓的損傷， 說：『平安了！平安了！』 其實沒有平安。
JER|6|15|他們行可憎之事，應當羞愧； 然而他們卻一點也不覺得羞愧， 也不知羞恥。 因此，他們必與仆倒的人一同仆倒， 我懲罰他們的時候， 他們必跌倒。」 這是耶和華說的。
JER|6|16|耶和華如此說： 「你們當站在路邊察看， 尋訪古老的路， 哪裏是完善的道路，就行走在其上； 這樣，你們自己必找到安息。 他們卻說：『我們不走。』
JER|6|17|我為你們設立守望的人， 要留心聽角聲。 他們卻說：『我們不聽。』
JER|6|18|因此，列國啊，當聽！ 會眾啊，要知道他們必遭遇的事。
JER|6|19|地啊，當聽！ 看哪，我必使災禍臨到這百姓， 是他們計謀所結的果子； 因為他們不肯留心聽我的話， 至於我的律法，他們也厭棄。
JER|6|20|從 示巴 來的乳香， 從遠方出的香菖蒲， 奉來給我有何用呢？ 你們的燔祭不蒙悅納； 你們的祭物，我也不喜悅。」
JER|6|21|所以耶和華如此說： 「看哪，我要將絆腳石放在這百姓面前； 父親和兒子要一同跌在其上， 鄰舍與朋友也都滅亡。」
JER|6|22|耶和華如此說： 「看哪，有一民族從北方而來； 有一大國被激起，從地極來到。
JER|6|23|他們拿弓和槍， 性情殘忍，不施憐憫； 他們的聲音如海浪澎湃。 錫安 哪， 他們都騎馬， 如上戰場的人擺陣攻擊你。」
JER|6|24|我們聽見這樣的風聲，手就發軟； 痛苦將我們抓住， 疼痛彷彿臨產的婦人。
JER|6|25|你們不要出到田野去， 也不要行走在路上， 因四圍有仇敵的刀劍和驚嚇。
JER|6|26|我的百姓 啊，應當腰束麻布，滾在灰中。 要悲傷，如喪獨子般痛痛哭號， 因為滅命的忽然臨到我們。
JER|6|27|我使你作我百姓的測試者 和考驗者 ， 使你知道並考驗他們的行為。
JER|6|28|他們極其悖逆， 到處毀謗人， 他們是銅是鐵， 全都敗壞了。
JER|6|29|風箱吹火，鉛被燒燬， 煉而又煉，終是徒然， 因為惡劣的還未除掉。
JER|6|30|人必稱他們為被拋棄的銀子， 因為耶和華已經拋棄了他們。
JER|7|1|耶和華的話臨到 耶利米 ，說：
JER|7|2|「你當站在耶和華殿的門口，在那裏宣講這話說：所有從這些門進來敬拜耶和華的 猶大 人哪，當聽耶和華的話。
JER|7|3|萬軍之耶和華－ 以色列 的上帝如此說：你們要改正你們的所作所為，我就使你們仍然居住這地 。
JER|7|4|不要倚靠虛謊的話，說：『這是耶和華的殿，是耶和華的殿，是耶和華的殿！』
JER|7|5|「你們若實在改正你們的所作所為，彼此誠然施行公平，
JER|7|6|不欺壓寄居的和孤兒寡婦，不在這地方流無辜人的血，也不隨從別神陷害自己，
JER|7|7|我就使你們仍然居住這地 ，就是我從古時所賜給你們祖先的地，從永遠到永遠。
JER|7|8|「看哪，你們倚靠虛謊無益的話語。
JER|7|9|你們豈可偷盜，殺害，姦淫，起假誓，向 巴力 燒香，隨從素不認識的別神，
JER|7|10|又來到這稱為我名下的殿，在我面前敬拜，說『我們平安無事』，為了要行這一切可憎的事呢？
JER|7|11|這稱為我名下的殿在你們眼中豈可看為賊窩呢？看哪，我真的都看見了。這是耶和華說的。
JER|7|12|你們到我的地方 示羅 去，就是我先前在那裏立為我名的居所，察看我因這百姓 以色列 的罪惡向那地方所行的事。
JER|7|13|現在，因你們行了這一切的事，我一再警戒你們，你們卻不聽從；我呼喚你們，你們也不回應。這是耶和華說的。
JER|7|14|所以我要向這稱為我名下、你們所倚靠的殿，與我所賜給你們和你們祖先的地這樣行，正如我從前向 示羅 所行的。
JER|7|15|我必將你們從我眼前趕出，正如趕出你們的眾弟兄，就是所有 以法蓮 的後裔。」
JER|7|16|「所以，你不要為這百姓祈禱；不要為他們呼求禱告，也不要為他們向我祈求，因我不聽你。
JER|7|17|他們在 猶大 城鎮和 耶路撒冷 街上所做的，你難道沒有看見嗎？
JER|7|18|孩子撿柴，父親燒火，婦女揉麵做餅，獻給天后，又向別神獻澆酒祭，惹我發怒。
JER|7|19|他們豈是惹我發怒呢？不是自己惹禍，以致臉上慚愧嗎？這是耶和華說的。
JER|7|20|所以主耶和華如此說：看哪，我必將我的怒氣和憤怒傾倒在這地方的人和牲畜身上、田野的樹木和地裏的出產上，它必燃燒，不會熄滅。」
JER|7|21|萬軍之耶和華－ 以色列 的上帝如此說：「你們要將燔祭加在你們的祭物上，又要吃肉；
JER|7|22|因為我將你們祖先從 埃及 地領出來的那日，燔祭和祭物的事我並沒有提說，也沒有吩咐他們。
JER|7|23|我只吩咐他們這一件事說：『你們當聽從我的話，我就作你們的上帝，你們也作我的子民。你們行走我所吩咐的一切道路，就可以得福。』
JER|7|24|他們卻不聽從，也不側耳而聽，竟隨從自己的計謀和頑梗的惡心去行，不進反退。
JER|7|25|自從你們祖先出 埃及 地的那日，直到今日，我每日一再差遣我的僕人眾先知到你們那裏去。
JER|7|26|你們卻不聽我，不側耳而聽，竟硬著頸項行惡，比你們的祖先更甚。
JER|7|27|「你要將這一切的話告訴他們，他們卻不聽你；呼喚他們，他們卻不回應。
JER|7|28|你要對他們說：『這就是不聽從耶和華－他們上帝的話、不領受訓誨的國民；誠信已從他們口中消失殆盡了。
JER|7|29|耶路撒冷 啊，要剪頭髮，扔掉它， 在光禿的高地唱哀歌， 因為耶和華棄絕、離棄了惹他發怒的世代。』」
JER|7|30|「 猶大 人行我眼中看為惡的事，將可憎之偶像立在稱為我名下的殿裏，玷污這殿。這是耶和華說的。
JER|7|31|他們在 欣嫩子谷 建造 陀斐特 的丘壇，要在火中焚燒自己的兒女。這並不是我所吩咐的，我心裏也從來沒有想過。
JER|7|32|因此，看哪，日子將到，這地方不再稱為 陀斐特 和 欣嫩子谷 ，反倒稱為 殺戮谷 。他們要在 陀斐特 埋葬屍首，甚至無處可葬。這是耶和華說的。
JER|7|33|並且這百姓的屍首要給空中的飛鳥和地上的走獸作食物，無人嚇走牠們。
JER|7|34|那時，我必止息 猶大 城鎮和 耶路撒冷 街上歡喜和快樂的聲音、新郎和新娘的聲音，因為這地必然荒蕪。」
JER|8|1|耶和華說：「那時，人必將 猶大 諸王和領袖的骸骨、祭司和先知的骸骨，以及 耶路撒冷 居民的骸骨，都從墳墓中取出來，
JER|8|2|散佈在太陽、月亮和天上眾星之下，就是他們從前所喜愛、所事奉、所隨從、所求問、所敬拜的。這些骸骨不被收殮，不被埋葬，必在地面上成為糞土。
JER|8|3|這邪惡家族所倖存的餘民，就是在我趕他們到的各處所剩下的 ，全都寧可選死不選活。這是萬軍之耶和華說的。」
JER|8|4|「你要對他們說，耶和華如此說： 人跌倒，不再起來嗎？ 人轉去，不再轉回來嗎？
JER|8|5|這 耶路撒冷 的百姓為何永久背道呢？ 他們抓住詭詐，不肯回頭。
JER|8|6|我留心聽，聽見他們說不誠實的話。 無人懊悔自己的惡行，說： 『我做的是甚麼呢？』 他們全都轉奔己路， 如馬直闖戰場。
JER|8|7|空中的鸛鳥知道自己的季節， 斑鳩、燕子與白鶴也守候當來的時令； 我的百姓卻不知道耶和華的法則。
JER|8|8|「你們怎麼說：『我們有智慧， 耶和華的律法在我們這裏』？ 看哪，其實文士的假筆舞弄虛假。
JER|8|9|智慧人慚愧，驚惶，被擒拿； 看哪，他們背棄耶和華的話， 還會有甚麼智慧呢？
JER|8|10|因此，我必將他們的妻子給別人， 將他們的田地給別人為業； 因為他們從最小的到最大的都貪圖不義之財， 從先知到祭司全都行事虛假。
JER|8|11|他們輕忽地醫治我百姓的損傷，說： 『平安了！平安了！』 其實沒有平安。
JER|8|12|他們行可憎之事，應當羞愧； 然而他們卻一點也不覺得羞愧， 又不知羞恥。 因此，他們必與仆倒的人一樣仆倒； 我懲罰他們的時候， 他們必跌倒。 這是耶和華說的。
JER|8|13|我必使他們全然滅絕； 葡萄樹上必沒有葡萄 ， 無花果樹上沒有果子， 葉子也必枯乾。 我所賜給他們的， 必離他們而去。 這是耶和華說的。」
JER|8|14|我們為何靜坐不動呢？ 我們當聚集，進入堅固城， 在那裏靜默不言； 因為耶和華－我們的上帝使我們靜默不言， 又將苦水給我們喝， 都因我們得罪了耶和華。
JER|8|15|我們指望平安， 卻得不著福氣； 指望痊癒的時刻， 看哪，受了驚惶。
JER|8|16|「從 但 那裏傳來敵人的馬噴氣的聲音， 壯馬發出嘶聲， 全地就都震動； 因為他們來吞滅這地和其上所有的， 吞滅這城與其中的居民。
JER|8|17|看哪，我必派蛇進到你們中間， 就是法術無法驅除的毒蛇， 牠們必咬你們。 這是耶和華說的。」
JER|8|18|憂愁時我尋找安慰 ， 我心在我裏面發昏。
JER|8|19|聽啊，是我百姓呼救的聲音從遠地傳來： 「耶和華不是在 錫安 嗎？ 錫安 的王不是在其中嗎？」 「他們為甚麼以自己雕刻的偶像 和外邦虛無的神明 惹我發怒呢？」
JER|8|20|「秋收已過，夏季已完， 我們還未得救！」
JER|8|21|因我百姓的損傷， 我也受了損傷。 我哀慟，驚惶將我抓住。
JER|8|22|在 基列 豈沒有乳香呢？ 在那裏豈沒有醫生呢？ 我百姓 為何得不著醫治呢？
JER|9|1|但願我的頭為水， 我的眼為淚水的泉源， 我好為我百姓 中被殺的人晝夜哭泣。
JER|9|2|惟願在曠野有旅客的客棧， 我好離開我的百姓而去； 因他們全都行姦淫， 是行詭詐的一黨。
JER|9|3|他們彎起舌頭像弓， 為要說謊話； 他們在國中增長勢力， 不是為誠信。 他們惡上加惡， 並不認識我。 這是耶和華說的。
JER|9|4|你們各人當謹防鄰舍， 不可信賴弟兄； 因為弟兄盡行欺騙， 鄰舍也都往來毀謗人。
JER|9|5|他們互相欺騙， 不說真話， 訓練自己的舌頭說謊， 竭盡所能地作惡。
JER|9|6|你居住在詭詐的人中； 他們因行詭詐 ，不願意認識我。 這是耶和華說的。
JER|9|7|所以萬軍之耶和華如此說： 「看哪，我要熬煉他們，考驗他們； 不然，為了我的百姓 ，我該如何行呢？
JER|9|8|他們的舌頭是毒箭，說話詭詐， 跟鄰舍口說平安， 心卻謀害他。
JER|9|9|我豈不因這些事向他們施行懲罰嗎？ 像這樣的國家，我豈能不報復呢？ 這是耶和華說的。」
JER|9|10|我要為山嶺哭泣悲哀， 為曠野的草場揚聲哀號； 因為都已枯焦，甚至無人經過。 牲畜的鳴叫聽不見， 空中的飛鳥和地上的走獸也都逃離。
JER|9|11|我必使 耶路撒冷 成為廢墟，為野狗的住處， 也必使 猶大 的城鎮荒廢，無人居住。
JER|9|12|誰是智慧人，可以明白這事？耶和華的口可向誰述說，使他傳講呢？這地為何毀滅，枯焦如曠野，無人經過呢？
JER|9|13|耶和華說：「因為這百姓離棄我在他們面前所設立的律法，不聽從我的話，不肯遵行，
JER|9|14|反隨從自己頑梗的心行事，照他們祖先所教訓的隨從諸 巴力 。」
JER|9|15|所以萬軍之耶和華－ 以色列 的上帝如此說：「看哪，我必將茵蔯給這百姓吃，又用苦水給他們喝。
JER|9|16|我要把他們分散在他們和他們祖宗所不認識的列國；我也要使刀劍追殺他們，直到將他們滅盡。」
JER|9|17|萬軍之耶和華如此說： 「你們要考慮， 將唱哀歌的婦女召來， 差人召善哭的婦女前來，
JER|9|18|叫她們速速為我們舉哀， 使我們淚眼汪汪， 使我們的眼皮湧出淚水。
JER|9|19|因為有哀聲從 錫安 傳來： 『我們竟然敗落！ 我們何等慚愧！ 我們撇下土地， 人拆毀了我們的房屋。』」
JER|9|20|婦女們哪，當聽耶和華的話， 領受他口中的言語； 當教導你們的女兒舉哀， 各人教導女伴唱哀歌。
JER|9|21|因為死亡從窗戶進來， 進入我們的宮殿， 從外邊剪除孩童， 從街上剪除少年。
JER|9|22|你當說，耶和華如此說： 人的屍首必倒在田野像糞土， 又像收割的人身後遺落的禾稼， 無人拾取。
JER|9|23|耶和華如此說：「智慧人不要因他的智慧誇口，勇士不要因他的力氣誇口，財主也不要因他的財富誇口；
JER|9|24|誇口的卻要誇自己有聰明，認識我是耶和華，知道我喜悅在世上施行慈愛、公平和公義。這是耶和華說的。
JER|9|25|「看哪，日子將到，這是耶和華說的，我要懲罰只在肉身受割禮的人，
JER|9|26|就是 埃及 、 猶大 、 以東 、 亞捫 人、 摩押 人，和住曠野所有剃鬢髮的人；因為列國都未受割禮， 以色列 全家心中也未受割禮。」
JER|10|1|以色列 家啊，要聽耶和華對你們所說的話，
JER|10|2|耶和華如此說： 「不要效法列國的行為， 任憑列國因天象驚惶， 你們不要驚惶。
JER|10|3|萬民的習俗是虛空的； 偶像 不過是從樹林中砍來的木頭， 是匠人用斧頭做成的手工。
JER|10|4|人用金銀妝飾它， 用釘子和錘子釘穩， 使它不動搖。
JER|10|5|偶像好像瓜田裏的稻草人， 不能說話，不能行走， 必須有人抬著。 不要怕它們， 因它們不能降禍， 也無力降福。」
JER|10|6|耶和華啊，沒有誰能與你相比！ 你本為大，你的名也大有能力。
JER|10|7|萬國的王啊，誰不敬畏你？ 敬畏你本是合宜的； 列國所有的智慧人中， 在他們一切的國度裏， 都沒有能與你相比的。
JER|10|8|他們如同畜牲，盡都愚昧。 偶像的訓誨算甚麼呢？ 偶像不過是木頭，
JER|10|9|錘煉的銀片是從 他施 來的， 金子則從 烏法 而來， 都是匠人和銀匠的手工； 又有藍色和紫色的衣服， 全都是巧匠的作品。
JER|10|10|惟耶和華是真上帝， 是活的上帝，是永遠的王。 他一發怒，大地震動； 他一惱恨，列國擔當不起。
JER|10|11|你們要對他們這樣說：「那些不是創造天地的神明，必從地上、從天下被除滅！」
JER|10|12|耶和華以能力創造大地， 以智慧建立世界， 以聰明鋪張穹蒼。
JER|10|13|他一出聲，天上就有眾水澎湃； 他使雲霧從地極上騰， 造電隨雨而閃， 從倉庫中吹出風來。
JER|10|14|人人都如同畜牲，毫無知識； 銀匠都因偶像羞愧， 他所鑄的偶像本是虛假， 它們裏面並無氣息。
JER|10|15|偶像都是虛無的， 是迷惑人的作品， 到受罰的時刻必被除滅。
JER|10|16|雅各 所得的福分不是這樣， 因主 是那創造萬有的， 以色列 是他產業的支派， 萬軍之耶和華是他的名。
JER|10|17|受圍困的居民哪，當收拾你的行囊， 離開這地。
JER|10|18|因為耶和華如此說： 「看哪，這一次，我必將此地的居民拋出去， 又必加害他們， 使他們覺悟 。」
JER|10|19|禍哉！我受損傷， 我的傷痕極其重大。 我卻說：「這真的是我必須忍受的痛苦。」
JER|10|20|我的帳棚毀壞， 我的繩索折斷， 我的兒女都離我而去，不在了。 再無人來支搭我的帳棚，掛起我的幔子。
JER|10|21|因為牧人如同畜牲， 沒有尋求耶和華， 所以不得順利； 他們的羊群也都分散了。
JER|10|22|有風聲！看哪，來了！ 有大擾亂從北方而來， 要使 猶大 的城鎮變為廢墟， 成為野狗的住處。
JER|10|23|耶和華啊，我知道人的道路不由自己， 行路的人也不能定自己的腳步。
JER|10|24|耶和華啊，求你按公平管教我， 不要在你的怒中懲治我， 免得你使我歸於無有。
JER|10|25|求你將憤怒傾倒在不認識你的列國中， 傾倒在不求告你名的各族上； 因為他們吞了 雅各 ，不但吞吃，而且滅絕， 使他的住處變為荒涼。
JER|11|1|耶和華的話臨到 耶利米 ，說：
JER|11|2|「當聽這約的話，告訴 猶大 人和 耶路撒冷 的居民，
JER|11|3|對他們說，耶和華－ 以色列 的上帝如此說：『不聽從這約之話的人必受詛咒。
JER|11|4|這約是我將你們祖先從 埃及 地領出來，脫離鐵爐的那日所吩咐他們的，說：你們要聽從我的話，照我所吩咐的一切去做。這樣，你們作我的子民，我也作你們的上帝，
JER|11|5|我好堅定我向你們列祖所起的誓，賞賜他們流奶與蜜之地，正如今日一樣。』」我就回應說：「耶和華啊，阿們！」
JER|11|6|耶和華對我說：「你要在 猶大 城鎮和 耶路撒冷 街市宣告這一切話，說：『當聽從遵行這約的話，
JER|11|7|因為我將你們祖先從 埃及 地領出來的那日，直到今日，都一再切切告誡他們說：當聽從我的話。
JER|11|8|他們卻不聽從，也不側耳而聽，竟隨從自己頑梗的惡心去行。我就使這約中一切詛咒的話臨到他們身上；這約是我吩咐他們遵行的，他們卻不遵行。』」
JER|11|9|耶和華對我說：「在 猶大 人和 耶路撒冷 居民中有同謀背叛的事。
JER|11|10|他們轉去效法他們祖先的惡行，不肯聽我的話，竟隨從別神，事奉它們。 以色列 家和 猶大 家違背了我與他們列祖所立的約。
JER|11|11|所以耶和華如此說：看哪，我必使災禍臨到他們，是他們不能逃脫的。他們向我哀求，我卻不聽。
JER|11|12|那時， 猶大 城鎮的人和 耶路撒冷 的居民要哀求他們燒香所供奉的神明；只是遭難的時候，這些神明一點也不能拯救他們。
JER|11|13|猶大 啊，你神明的數目與你城鎮的數目相等；你所築可恥的壇，就是向 巴力 燒香的壇 ，也與 耶路撒冷 街道的數目相等。
JER|11|14|「所以你不要為這百姓祈禱，也不要為他們呼求禱告，因為他們遭難向我哀求的時候，我必不應允。
JER|11|15|我所親愛的既多設惡謀，還能在我殿中做甚麼呢？你因作惡就喜樂，聖肉要離開你。
JER|11|16|從前耶和華給你起名叫青橄欖樹，又華美又結好果子；如今他用一聲巨響點火在其上，枝子就折斷了。
JER|11|17|「原來栽培你的萬軍之耶和華已經說要降禍給你，是因 以色列 家和 猶大 家行惡。他們向 巴力 燒香，惹我發怒，是自作自受。」
JER|11|18|耶和華指示我，我才知道； 你將他們所做的給我指明。
JER|11|19|我像柔順的羔羊被牽去宰殺， 並不知道他們設計謀害我： 「我們把樹連果子都滅了吧！ 把他從活人之地剪除， 使他的名不再被記得。」
JER|11|20|按公義判斷、察驗人肺腑心腸的萬軍之耶和華啊， 求你使我得見你在他們身上報仇， 因我已將我的案件向你稟明了。
JER|11|21|所以，耶和華論到尋索你命的 亞拿突 人如此說：「他們說：你不要奉耶和華的名說預言，免得你死在我們手中。
JER|11|22|所以萬軍之耶和華如此說：看哪，我必懲罰他們；他們的壯丁必被刀劍殺死，他們的兒女必因饑荒而死，
JER|11|23|他們當中必無任何倖存者；因為在他們受罰之年，我必使災禍臨到 亞拿突 人。」
JER|12|1|耶和華啊，我與你爭辯的時候， 你總是顯為義； 但有一件，我還要與你理論： 惡人的道路為何亨通呢？ 大行詭詐的為何得安逸呢？
JER|12|2|你栽培了他們， 他們也扎了根， 長大，而且結果。 他們的口與你相近， 心卻與你遠離。
JER|12|3|耶和華啊，你認識我，看見我， 你察驗我向你的心如何。 求你將他們拉出來， 如將宰的羊， 為殺戮的日子分別出來。
JER|12|4|這地悲哀， 一切田野的青草枯乾要到幾時呢？ 因其上居民的惡行， 牲畜和飛鳥都滅絕了。 因為他們說：「他看不見 我們的結局 。」
JER|12|5|「你與步行的人同跑， 尚且覺得累， 怎能與馬賽跑呢？ 你在安全之地尚且會跌倒 ， 在 約旦河 邊的叢林要怎麼辦呢？
JER|12|6|因為連你兄弟和你父家都以詭詐待你， 甚至在你後邊大聲喊叫。 雖然他們向你說好話， 你也不要相信他們。」
JER|12|7|我離棄了我的殿宇， 撇棄了我的產業， 將我心裏所親愛的交在她 仇敵手中。
JER|12|8|我的產業向我如林中的獅子， 出聲攻擊我， 因此我恨惡她。
JER|12|9|我的產業向我如斑點的鷙鳥， 有鷙鳥在四圍攻擊她。 你們去聚集田野的百獸， 叫牠們來吞吃吧！
JER|12|10|許多牧人毀壞我的葡萄園， 踐踏我的地產， 使我美好的地產變為荒涼的曠野。
JER|12|11|他們使地荒涼； 地既荒涼，就向我哀哭。 全地荒涼，卻無人在意。
JER|12|12|滅命的來到曠野中一切光禿的高地； 耶和華的刀從地這邊直到地那邊，盡行殺滅， 凡血肉之軀都不得平安。
JER|12|13|他們種的是麥子， 收的卻是荊棘； 辛辛苦苦卻無收穫。 因耶和華的烈怒， 你們必為自己的收成感到羞愧。
JER|12|14|耶和華如此說：「看哪，我要將所有的惡鄰拔出本地，他們曾佔據了我賜給 以色列 百姓所承受的產業；我也要將 猶大 家從他們中間拔出來。
JER|12|15|我拔出他們以後，必回轉過來憐憫他們，使他們歸回，各歸本業，各歸故土。
JER|12|16|他們若殷勤學習我百姓的道，指著我的名起誓：『我指著永生的耶和華起誓』，正如他們從前教我百姓指著 巴力 起誓，他們必在我百姓中得以建立。
JER|12|17|他們若是不聽，我必拔出那國，不但拔出，還要毀滅。這是耶和華說的。」
JER|13|1|耶和華對我如此說：「你去買一條麻布帶子，束在你腰上，不可把它泡在水裏。」
JER|13|2|我就照耶和華的話，買了一條帶子，束在我的腰上。
JER|13|3|耶和華的話第二次臨到我，說：
JER|13|4|「要拿你所買、在你腰上的帶子，起來往 幼發拉底河 去，把腰帶藏在那裏的磐石穴中。」
JER|13|5|我就去，照著耶和華命令我的，把腰帶藏在 幼發拉底河 邊。
JER|13|6|過了多日，耶和華對我說：「你起來往 幼發拉底河 去，把我命令你藏在那裏的腰帶取出來。」
JER|13|7|我就往 幼發拉底河 去，把那腰帶從我所藏的地方挖出來。看哪，腰帶已經破爛，毫無用處了。
JER|13|8|耶和華的話臨到我，說：
JER|13|9|「耶和華如此說：我要照樣敗壞 猶大 的驕傲和 耶路撒冷 的狂傲。
JER|13|10|這惡民不肯聽我的話，按自己頑梗的心而行，隨從別神，事奉敬拜它們；這惡民必像這腰帶，毫無用處。
JER|13|11|腰帶怎樣緊貼人的腰，照樣，我也曾使 以色列 全家和 猶大 全家緊貼著我，歸我為子民，使我得名聲，得頌讚，得榮耀；他們卻不肯聽從。這是耶和華說的。」
JER|13|12|「所以你要對他們說：『耶和華－ 以色列 的上帝如此說：各罈都要裝滿酒。』他們必對你說：『我們豈不知道各罈都要裝滿酒嗎？』
JER|13|13|你就對他們說：『耶和華如此說：看哪，我必使這地所有的居民，就是坐 大衛 寶座的君王、祭司和先知，並 耶路撒冷 所有的居民，都酩酊大醉。
JER|13|14|我要使他們彼此衝突，連父與子也互相衝突；我必不可憐，不顧惜，不憐憫，以致將他們滅絕。這是耶和華說的。』」
JER|13|15|你們當聽，當側耳而聽； 不可驕傲，因為耶和華已經吩咐了。
JER|13|16|當耶和華－你們的上帝 尚未使黑暗來臨， 在昏暗的山上 你們的腳未絆跌以前， 要將榮耀歸給他。 你們盼望光明， 他卻使光明變為死蔭， 成為幽暗。
JER|13|17|你們若不聽這話， 我的心必因你們的驕傲暗自哭泣； 我的眼必痛哭流淚， 因為耶和華的羊群被擄去了。
JER|13|18|你要對君王和太后說： 「你們當自卑，坐下； 因你們的王冠， 就是你們華美的冠冕已經掉落了 。」
JER|13|19|尼革夫 的城鎮都被關閉， 無人打開； 猶大 全被擄掠， 擄掠淨盡。
JER|13|20|你們要舉目觀看從北方來的人。 先前賜給你的羊群， 就是你所引以為榮的羊， 現今在哪裏呢？
JER|13|21|耶和華立你自己所教導的盟友， 立他們為頭來轄制你， 你還有甚麼話可說呢？ 痛苦豈不將你抓住像臨產的婦人嗎？
JER|13|22|你若心裏說：「這一切的事為何臨到我呢？」 是因你罪孽甚多。 你的下襬揭起， 你的腳跟受傷。
JER|13|23|古實 人豈能改變皮膚呢？ 豹豈能改變斑點呢？ 若能，你們這善於行惡的便能行善了。
JER|13|24|我必吹散他們， 如碎秸隨曠野的風飄動。
JER|13|25|這是你所當得的， 是我量給你的報應 ； 因為你忘記了我， 倚靠虛假 。 這是耶和華說的。
JER|13|26|我要揭起你的下襬， 蒙在你臉上， 顯露你的羞恥。
JER|13|27|你在田野的山上行姦淫， 發嘶聲，謀淫亂， 這些可憎之事我都看見了。 耶路撒冷 啊，你有禍了！ 你不肯潔淨 還要等到幾時呢？
JER|14|1|耶和華的話臨到 耶利米 ，論到旱災的事：
JER|14|2|「 猶大 悲哀，城門衰敗； 眾人坐在地上哀慟， 耶路撒冷 的哀聲上達。
JER|14|3|他們的貴族打發童僕去打水； 他們來到水池， 找不到水，就拿著空器皿， 蒙羞慚愧，抱頭而回。
JER|14|4|因為無雨降在地上，土地就乾裂， 農夫為此蒙羞抱頭。
JER|14|5|田野的母鹿因為無草 也撇棄才生的小鹿。
JER|14|6|野驢站在光禿的高地喘氣，好像野狗； 牠們的眼目因無草而失明。」
JER|14|7|耶和華啊，雖然我們的罪孽控告我們， 求你為你名的緣故行動吧！ 我們本是多次背道，得罪了你。
JER|14|8|以色列 所盼望，在患難時作他救主的啊， 你在這地為何像寄居的， 又如旅行的只住一夜呢？
JER|14|9|你為何像受驚嚇的人， 像不能救人的勇士呢？ 耶和華啊，你在我們中間， 我們是稱為你名下的人， 求你不要離開我們。
JER|14|10|耶和華論到這百姓如此說： 「這百姓喜愛遊蕩， 不約束自己的腳步， 所以耶和華不悅納他們。 現今他要記起他們的罪孽， 懲罰他們的罪惡。」
JER|14|11|耶和華又對我說：「不要為這百姓求福。
JER|14|12|他們禁食的時候，我不聽他們的呼求；他們獻燔祭和素祭，我也不悅納。我卻要用刀劍、饑荒、瘟疫滅絕他們。」
JER|14|13|我就說：「唉！主耶和華，看哪，那些先知常對他們說：『你們必不見刀劍，也不遭饑荒；耶和華要在這地方賞賜你們真正的平安。』」
JER|14|14|耶和華對我說：「那些先知託我的名說假預言，我並未差遣他們，沒有吩咐他們，也沒有對他們說話；他們向你們預言的是虛假的異象、占卜、虛無，以及心中的詭詐。
JER|14|15|所以耶和華如此說：『論到託我名說預言的那些先知，我並未差遣他們；他們說這地不會有刀劍、饑荒，其實那些先知自己必被刀劍、饑荒滅絕。
JER|14|16|聽他們說預言的百姓必因饑荒、刀劍被扔在 耶路撒冷 的街道上，無人埋葬。他們連妻子帶兒女，都是如此。我必將他們的惡倒在他們身上。』」
JER|14|17|你要向他們說這些話： 願我眼淚汪汪， 晝夜不息， 因為少女─我百姓 受了重大的打擊， 傷口極其嚴重。
JER|14|18|我若出到田間， 看哪，有被刀殺的； 我若進入城內， 看哪，有因饑荒患病的； 先知和祭司也在各地往來經商， 不知如何是好。
JER|14|19|你全然棄絕 猶大 嗎？ 你的心厭惡 錫安 嗎？ 你為何擊打我們，使我們無法得醫治呢？ 我們指望平安，卻得不著福氣； 指望痊癒，看哪，受了驚惶。
JER|14|20|耶和華啊，我們承認自己的罪惡 和我們祖先的罪孽， 因我們得罪了你。
JER|14|21|求你為你名的緣故， 不厭惡，不輕視你榮耀的寶座。 求你記念， 不要違背你與我們所立的約。
JER|14|22|外邦虛無的神明 中有能降雨的嗎？ 天能自降甘霖嗎？ 耶和華－我們的上帝啊，不是你嗎？ 我們要等候你， 因為這一切都是你所造的。
JER|15|1|耶和華對我說：「雖有 摩西 和 撒母耳 站在我面前，我的心也不顧惜這百姓。你把他們從我眼前趕出，叫他們出去吧！
JER|15|2|他們若問你說：『我們往哪裏去呢？』你就告訴他們，耶和華如此說： 『定為死亡的，必致死亡； 定為刀殺的，必被刀殺； 定為饑荒的，必遭饑荒； 定為擄掠的，必被擄掠。』」
JER|15|3|「我命定四樣災害臨到他們，就是刀劍殺戮、群狗拖拉、空中的飛鳥和地上的走獸吞吃毀滅。這是耶和華說的。
JER|15|4|我必使地上萬國因他們而驚駭，都因 希西家 的兒子 猶大 王 瑪拿西 在 耶路撒冷 所做的事。」
JER|15|5|耶路撒冷 啊，有誰同情你呢？ 有誰為你悲傷呢？ 有誰轉身問你安呢？
JER|15|6|你棄絕了我， 轉身退後； 因此我伸手攻擊你，毀滅你， 我已憐憫到厭煩了。 這是耶和華說的。
JER|15|7|我在境內各關口 用簸箕篩我的百姓， 使他們喪掉兒女， 又毀滅他們， 他們仍不轉離所行的道。
JER|15|8|他們的寡婦在我面前比海沙更多； 我使滅命者在正午來到， 攻擊年輕人的母親， 使痛苦驚嚇忽然臨到她身上。
JER|15|9|生過七個孩子的婦人衰弱； 尚在白晝，太陽忽然落下， 她就抱愧蒙羞。 我必當著敵人的面， 將他們當中的倖存者交給刀劍。 這是耶和華說的。
JER|15|10|我的母親哪，我有禍了！因你生我作全地爭相指控的人。我素來沒有借貸給人，人也沒有借貸給我，人人卻都咒罵我。
JER|15|11|耶和華說：「我必定釋放 你，使你得福氣。災禍苦難來臨時，我必使仇敵央求你。
JER|15|12|人豈能將銅與鐵，就是北方的鐵折斷呢？
JER|15|13|「我必因你在四境之內所犯的一切罪，將你的貨物財寶當掠物，白白地交出來 。
JER|15|14|我要使你的仇敵過去，到你所不認識的地方 ，因為你們要被我怒中所起的火焚燒。」
JER|15|15|耶和華啊，你是知道的； 求你記念我，眷顧我， 向迫害我的人為我報仇； 不要把我取去，因你不輕易發怒， 要知道我為你的緣故受了凌辱。
JER|15|16|耶和華－萬軍之上帝啊， 我得著你的話就把它們吃了， 你的話是我心中的歡喜快樂； 因我是稱為你名下的人。
JER|15|17|我並未坐在享樂人的會中歡樂； 因你的手，我就獨自靜坐， 你使我滿心憤慨。
JER|15|18|我的痛苦為何長久不止呢？ 我的傷痕為何無法可醫，不能痊癒呢？ 難道你以詭詐待我，像流乾的河道嗎？
JER|15|19|所以耶和華如此說：「你若回轉， 我就使你歸回， 站在我面前。 你若能將寶物和無用之物分別出來， 你就可以當作我的口。 他們必歸向你， 你卻不可歸向他們。
JER|15|20|我必使你向這百姓成為堅固的銅牆。 他們必攻擊你，卻不能勝過你； 因我與你同在，要拯救你，搭救你。 這是耶和華說的。
JER|15|21|我必搭救你脫離惡人的手， 救贖你脫離殘暴之人的手。」
JER|16|1|耶和華的話又臨到我，說：
JER|16|2|「你不可在這地方娶妻，為自己生兒育女。
JER|16|3|因為論到在這地方所生的兒女，又論到在這國中生他們的父母，耶和華如此說：
JER|16|4|他們必死於致命的疾病，無人哀哭，不得埋葬，在地上如糞土，因刀劍和饑荒而滅絕；他們的屍首必給空中的飛鳥和地上的走獸作食物。
JER|16|5|「耶和華如此說：不要進入喪家，不要去哀哭，也不要為他們悲傷，因我已使我的平安、慈愛、憐憫離開這百姓。這是耶和華說的。
JER|16|6|他們連大帶小，都必在這地死亡，不得埋葬。人必不為他們哀哭，不為他們割劃自己，也不剃光頭。
JER|16|7|有喪事，人不為他們擘餅 ，也不因死人安慰他們；他們喪父喪母，人也不給他們一杯酒安慰他們。
JER|16|8|你不可進入宴樂的家，與人同坐又吃又喝，
JER|16|9|因為萬軍之耶和華－ 以色列 的上帝如此說：看哪，你們還活著的日子，我必在你們眼前止息這地方歡喜和快樂的聲音、新郎和新娘的聲音。
JER|16|10|「你將這一切的話指示這百姓，他們若問你說：『耶和華為甚麼說，要降這大災禍攻擊我們呢？我們有甚麼罪孽呢？我們向耶和華－我們的上帝犯了甚麼罪呢？』
JER|16|11|你就對他們說：『因為你們祖先離棄了我，隨從別神，事奉敬拜它們，卻離棄我，不遵守我的律法。這是耶和華說的。
JER|16|12|你們行惡比你們祖先更甚，看哪，各人隨從自己頑梗的惡心行事，不聽從我。
JER|16|13|所以我必將你們從這地趕出，直趕到你們和你們祖先素不認識之地。你們在那裏晝夜必事奉別神，因為我必不再向你們施恩。』」
JER|16|14|「看哪，日子將到，人必不再指著那領 以色列 人從 埃及 地上來的永生耶和華起誓。這是耶和華說的。
JER|16|15|人卻要指著那領 以色列 人離開北方之地，離開他們被趕到的各國之永生的耶和華起誓；並且我要領他們歸回我從前賜給他們祖先之地。」
JER|16|16|「看哪，我要差派許多打魚的捕獲他們；以後，我也要派許多打獵的，從各山上、各岡上、各石穴中獵取他們。這是耶和華說的。
JER|16|17|因我的眼目察看他們一切的行為；他們不能在我面前遮掩，他們的罪孽也不能在我眼前隱藏。
JER|16|18|我要先加倍報應他們的罪孽和罪惡，因為他們以可憎之偶像的屍首使我的地玷污，使我的產業充斥可厭之物。」
JER|16|19|耶和華啊，你是我的力量， 是我的保障， 在患難之日是我的避難所。 列國的人必從地極來到你這裏，說： 「我們祖先所承受的， 不過是虛假，是虛空無益之物。
JER|16|20|人豈可為自己製造神明呢？ 其實它們不是神明。」
JER|16|21|「所以，看哪，我要使他們知道，就是這一次使他們知道我的手和我的能力。他們就知道我的名是耶和華了。」
JER|17|1|猶大 的罪是用鐵筆、用金剛石記錄的，銘刻在他們的心版和祭壇角上。
JER|17|2|他們的兒女思念他們在高岡上、青翠樹旁的祭壇和 亞舍拉 。
JER|17|3|我田野的山哪，因你在全境內的丘壇所犯的罪，我必使你的財富和一切的財寶成為掠物。
JER|17|4|因自己所做的 ，你必失去我所賜給你的產業。我也必使你在你所不認識的地服侍你的仇敵；因你們激起了我的怒火，直燒到永遠。
JER|17|5|耶和華如此說： 「倚靠人，以血肉為膀臂， 心中離棄耶和華的， 那人該受詛咒！
JER|17|6|他必像沙漠裏的矮樹， 不見福樂來到； 他要住在曠野乾旱之處， 無人居住的鹽地。
JER|17|7|倚靠耶和華、以耶和華為他所仰賴的， 那人有福了！
JER|17|8|他必像樹栽於水旁， 在河邊扎根， 炎熱來到，毫不察覺 ， 葉子仍必青翠； 在乾旱之年，一無掛慮， 並且結果不止。
JER|17|9|「人心比萬物都詭詐， 壞到極處， 誰能識透呢？
JER|17|10|我－耶和華是鑒察人心，考驗人肺腑的， 要按各人所行的和他做事的結果報應他。」
JER|17|11|那不按正道得財富的， 好像鷓鴣孵不是自己生的； 到了中年，財富必離開他， 終久他必成為愚頑人。
JER|17|12|我們的聖所是榮耀的寶座， 從太初就在高處。
JER|17|13|耶和華－ 以色列 的盼望啊， 凡離棄你的必蒙羞。 離我而去的， 他們必被寫在地裏， 因為他們離棄耶和華，這活水的泉源。
JER|17|14|耶和華啊，求你醫治我，我就痊癒， 拯救我，我便得救； 因你是我所讚美的。
JER|17|15|看哪，他們對我說： 「耶和華的話在哪裏呢？ 讓它應驗吧！」
JER|17|16|至於我，我並沒有逃避作牧人跟隨你 ， 也沒有想望那災殃的日子； 這是你所知道的。 我嘴唇所出的都在你面前。
JER|17|17|不要使我因你驚恐； 災禍來臨時，你是我的避難所。
JER|17|18|願那些迫害我的蒙羞， 卻不要使我蒙羞； 使他們驚惶， 卻不要使我驚惶； 願災禍的日子臨到他們， 以加倍的毀壞毀壞他們。
JER|17|19|耶和華對我如此說：「你去站在 猶大 君王出入的 平民門 ，和 耶路撒冷 的各城門口，
JER|17|20|對他們說：『你們這 猶大 君王、 猶大 眾人和 耶路撒冷 所有的居民，凡從這些城門進入的，都當聽耶和華的話。
JER|17|21|耶和華如此說：你們要謹慎，不可在安息日挑甚麼擔子進入 耶路撒冷 的城門，
JER|17|22|也不可在安息日從家中挑擔子出去。無論何工都不可做，只要以安息日為聖日，正如我所吩咐你們祖先的。』
JER|17|23|他們卻不聽從，也不側耳而聽，竟硬著頸項不聽，不肯領受訓誨。
JER|17|24|「你們若留意聽從我，在安息日不挑甚麼擔子進入這城的各門，只以安息日為聖日，在那日不做任何工作，這是耶和華說的，
JER|17|25|就必有坐 大衛 寶座的君王和領袖，與 猶大 人，並 耶路撒冷 的居民，或坐車，或騎馬，進入這城的各門，而且這城必存到永遠。
JER|17|26|也必有人從 猶大 城鎮和 耶路撒冷 四圍的各處，從 便雅憫 地、 謝非拉 、山區，並 尼革夫 而來，都帶燔祭和祭物，素祭和乳香，並感謝祭，到耶和華的殿去。
JER|17|27|你們若不聽從我，不以安息日為聖日，仍在安息日挑擔子進入 耶路撒冷 的各城門，我必在城門中點火；這火必燒燬 耶路撒冷 的宮殿，不會熄滅。」
JER|18|1|耶和華的話臨到 耶利米 ，說：
JER|18|2|「你起來，下到陶匠的家裏去，在那裏我要使你聽見我的話。」
JER|18|3|我就下到陶匠的家裏去，看哪，他在轉盤上做器皿。
JER|18|4|陶匠用泥做的器皿在他手中做壞了，他就用它另做別的器皿，照他看為好的去做。
JER|18|5|耶和華的話臨到我，說：
JER|18|6|「 以色列 家啊，我待你們豈不能像這陶匠弄泥嗎？ 以色列 家，看哪，泥在陶匠的手中怎樣，你們在我的手中也怎樣。這是耶和華說的。
JER|18|7|我何時論到一邦或一國說，要拔出、拆毀、毀壞；
JER|18|8|我所說的那一邦若回轉離開他們的惡，我就改變心意，不將我想要施行的災禍降與他們。
JER|18|9|我何時論到一邦或一國說，要建立、栽植；
JER|18|10|他們若行我眼中看為惡的事，不聽從我的話，我就改變心意，不將我所說的福氣賜給他們。
JER|18|11|現在你要對 猶大 人和 耶路撒冷 的居民說：『耶和華如此說：看哪，我捏塑災禍降給你們，定意懲罰你們。你們各人當回轉離開所行的惡道，改正你們的所作所為。』
JER|18|12|「他們卻說：『沒有用的，我們要照自己的計謀去行，各人要隨自己頑梗的惡心行事。』」
JER|18|13|「所以，耶和華如此說： 你們且往各國訪問， 有誰聽見這樣的事？ 少女 以色列 行了一件極恐怖的事。
JER|18|14|黎巴嫩 的雪豈能從田野 的磐石上融化呢？ 從遠處 流下的涼水豈能乾涸呢？
JER|18|15|我的百姓竟忘記我， 向那虛無的神明 燒香， 它們使百姓在所行的路上、在古道上絆跌， 去行未修築的斜路，
JER|18|16|他們的地就變為荒涼， 長久被人嘲笑； 凡經過這地的必驚駭搖頭。
JER|18|17|在仇敵面前，我必如東風颳散他們， 遭難的日子，我要以背向他們， 不以臉看他們。」
JER|18|18|他們說：「來吧！讓我們設計謀害 耶利米 ；因為我們有祭司講律法，有智慧人設謀略，有先知說預言，都未曾斷絕。來吧！讓我們用舌頭攻擊他，不要理他一切的話。」
JER|18|19|耶和華啊，求你留心聽我， 且聽那些指控我的人的話。
JER|18|20|人豈可以惡報善呢？ 他們竟挖坑要害我的性命！ 求你記念我站在你面前為他們說好話， 要使你的憤怒轉離他們。
JER|18|21|因此，願他們的兒女忍受饑荒， 願他們死於刀劍之手； 願他們的妻無子，且作寡婦， 願他們的男人被死亡所滅， 他們的壯丁在陣上被刀擊殺。
JER|18|22|你使敵軍忽然臨到他們的時候， 願人聽見哀聲從他們的屋內發出； 因他們挖坑要捉拿我， 暗設羅網要絆我的腳。
JER|18|23|耶和華啊，他們要殺我的那一切計謀， 你都知道。 求你不要赦免他們的罪孽， 也不要從你面前塗去他們的罪惡。 願他們在你面前跌倒， 願你在發怒的時候對付他們。
JER|19|1|耶和華如此說：「你去買陶匠的瓷瓶 ，你和 百姓中的長老、位尊的祭司
JER|19|2|出去到 欣嫩子谷 、 哈珥西 的門口，在那裏宣告我所吩咐你的話，
JER|19|3|說：『 猶大 君王和 耶路撒冷 的居民哪，當聽耶和華的話。萬軍之耶和華－ 以色列 的上帝如此說：看哪，我必使災禍臨到這地方，凡聽見的人都必耳鳴；
JER|19|4|因為他們和他們祖先，並 猶大 君王都離棄我，使這地方與我疏遠 ，在這裏向素不認識的別神燒香，又使這地方遍滿無辜人的血。
JER|19|5|他們建造 巴力 的丘壇，要在火中焚燒自己的兒女，作為燔祭獻給 巴力 。這不是我命令的，不是我吩咐的，我心裏也從來沒有想過。
JER|19|6|因此，看哪，日子將到，這地方不再稱為 陀斐特 和 欣嫩子谷 ，反倒稱為 殺戮谷 。這是耶和華說的。
JER|19|7|我要在這地方使 猶大 和 耶路撒冷 的計謀落空，也必使他們在仇敵面前倒在刀下，倒在尋索其命的人手下。我要把他們的屍首給空中的飛鳥和地上的走獸作食物。
JER|19|8|我必使這城令人驚駭嘲笑；凡路過的，必因這城所遭的災難驚駭嘲笑。
JER|19|9|仇敵和尋索其命的人追逼他們，使他們落在圍困窘迫之中，我必使他們各人吃自己兒女的肉和朋友的肉。』
JER|19|10|「你要在跟你同去的人眼前打碎那瓶，
JER|19|11|對他們說：『萬軍之耶和華如此說：我要打碎這百姓和這城，正如人打碎陶匠的器皿，不能再使其完整。他們要在 陀斐特 埋葬，甚至無處可葬。
JER|19|12|我必向這地方和其中的居民如此行，使這城與 陀斐特 一樣。這是耶和華說的。
JER|19|13|耶路撒冷 的房屋和 猶大 君王的宮殿，就是他們在其上向天上的萬象燒香、向別神獻澆酒祭的宮殿房屋，都必被玷污，和 陀斐特 一樣。』」
JER|19|14|耶利米 從耶和華差他去說預言的 陀斐特 回來，站在耶和華殿的院中對眾百姓說：
JER|19|15|「萬軍之耶和華－ 以色列 的上帝如此說：『看哪，我必使我所說的一切災禍臨到這城和屬它的城鎮，因為他們硬著頸項不聽我的話。』」
JER|20|1|音麥 的兒子 巴施戶珥 祭司作耶和華殿的總管，聽見 耶利米 預言這些事，
JER|20|2|就打 耶利米 先知，用耶和華殿裏 上便雅憫門 內的枷鎖，把他鎖在那裏。
JER|20|3|次日， 巴施戶珥 開枷釋放 耶利米 。於是 耶利米 對他說：「耶和華不叫你的名為 巴施戶珥 ，而叫你 瑪歌珥‧米撒畢 ，
JER|20|4|因耶和華如此說：『看哪，我要使你和你的眾朋友驚嚇；你們要親眼看見他們倒在仇敵的刀下。我必將 猶大 人全都交在 巴比倫 王的手中，他要把他們擄到 巴比倫 去，用刀殺他們。
JER|20|5|我要將這城中一切的貨財和勞碌得來的，並一切的珍寶，以及 猶大 君王所有的寶物，都交在仇敵手中。仇敵要搶奪他們，抓住他們，把他們帶到 巴比倫 去。
JER|20|6|你， 巴施戶珥 ，和所有住在你家中的人都必被擄；你和你的朋友，就是你向他們說假預言的，都要到 巴比倫 去，死在那裏，葬在那裏。』」
JER|20|7|耶和華啊，你欺哄了我， 我也被你欺哄了。 你比我強，並且得勝。 我終日成為笑柄， 人人都戲弄我。
JER|20|8|我每逢講話的時候，就哀嘆， 我喊叫：「有暴力和毀滅！」 因為耶和華的話終日成了我的凌辱和譏刺。
JER|20|9|我若說：「我不再提耶和華， 也不再奉他的名講論」， 我心裏便覺得 似乎有燒著的火悶在我骨中， 我忍受不住，不能自禁。
JER|20|10|我聽見許多的毀謗， 四圍都是驚嚇； 連我知己朋友都看著我跌倒： 「告他吧，我們要告他！ 或者他被引誘， 我們就能勝他， 在他身上報仇。」
JER|20|11|然而，耶和華與我同在， 好像可怕的勇士。 因此，迫害我的都絆跌， 不能得勝； 他們大大蒙羞， 由於行事沒有智慧， 必永遠受那不能忘懷的羞辱。
JER|20|12|考驗義人、察看人肺腑心腸的萬軍之耶和華啊， 求你使我得見你在他們身上報仇， 因我已將我的案件向你稟明了。
JER|20|13|你們要向耶和華唱歌！ 要讚美耶和華！ 因他救了窮人的性命 脫離惡人的手。
JER|20|14|願我出生的那日受詛咒！ 願我母親生我的那天不蒙福！
JER|20|15|報信給我父親說 「你得了兒子」， 使我父親甚歡喜的， 願那人受詛咒。
JER|20|16|願那人像耶和華所傾覆而不憐惜的城鎮； 願他早晨聽見哀聲， 中午聽見吶喊；
JER|20|17|因他沒有在我未出胎就把我殺了， 以致我母親成為我的墳墓， 她卻一直懷著胎 。
JER|20|18|我為何出胎見勞碌愁苦， 在羞愧中度盡我的年日呢？
JER|21|1|耶和華的話臨到 耶利米 。那時， 西底家 王差派 瑪基雅 的兒子 巴施戶珥 和 瑪西雅 的兒子 西番雅 祭司到他那裏去，說：
JER|21|2|「請你為我們求問耶和華，因為 巴比倫 王 尼布甲尼撒 前來攻擊我們；或者耶和華照他一切奇妙的作為待我們，使 巴比倫 王離開我們而去。」
JER|21|3|耶利米 對他們說：「你們當對 西底家 這樣說：
JER|21|4|『耶和華－ 以色列 的上帝如此說：看哪，我要使你們手中的兵器，就是你們與城外圍困你們的 巴比倫 王和 迦勒底 人打仗所用的兵器轉回來，把它們聚集在這城中。
JER|21|5|我要在怒氣、憤怒和大惱怒中，用伸出來的手和大能的膀臂，親自攻擊你們；
JER|21|6|又要擊打這城的居民，他們連人帶牲畜都必遭遇大瘟疫而死亡。
JER|21|7|以後，我要將 猶大 王 西底家 和他的臣僕百姓，就是在城內，從瘟疫、刀劍、饑荒中倖存的人，都交在 巴比倫 王 尼布甲尼撒 手中，交在仇敵和尋索其命的人手中。 巴比倫 王必用刀擊殺他們，不顧惜，不同情，不憐憫。這是耶和華說的。』
JER|21|8|「你要對這百姓說：『耶和華如此說：看哪，我將生命的路和死亡的路擺在你們面前。
JER|21|9|住在這城裏的必遭刀劍、饑荒、瘟疫而死；但出去投降圍困你們之 迦勒底 人的必得存活，保全自己的性命。
JER|21|10|我向這城板臉，降禍不降福；這城必交在 巴比倫 王的手中，他必用火焚燒。這是耶和華說的。』」
JER|21|11|「至於 猶大 王的家，你們當聽耶和華的話。
JER|21|12|大衛 家啊，耶和華如此說： 『每早晨你們要施行公平， 拯救被搶奪的脫離欺壓者的手， 免得我的憤怒因你們的惡行發作， 如火燃起，無人能熄滅。』
JER|21|13|住在山谷和平原磐石上的居民啊， 看哪，我與你們為敵， 因為你們說：『誰能下來攻擊我們？ 誰能進入我們的住處呢？』 這是耶和華說的。
JER|21|14|我必按你們行事的結果懲罰你們， 也必使火在 耶路撒冷 的林中燃起， 將四圍所有的盡行燒滅。 這是耶和華說的。」
JER|22|1|耶和華如此說：「你要下到 猶大 王的宮中，在那裏說這話，
JER|22|2|你要說：『坐 大衛 寶座的 猶大 王啊，你和你的臣僕，並進入這些城門的百姓，都當聽耶和華的話。
JER|22|3|耶和華如此說：你們要施行公平和公義，拯救被搶奪的脫離欺壓者的手，不可虧負寄居的和孤兒寡婦，不可用殘暴對待他們，也不可在這地方流無辜人的血。
JER|22|4|你們若切實遵行這話，就必有坐 大衛 寶座的君王和他的臣僕百姓，或坐車或騎馬，從這王宮的各門進入。
JER|22|5|你們若不聽這些話，我指著自己起誓，這王宮必變為廢墟。這是耶和華說的。』
JER|22|6|耶和華論到 猶大 王的家如此說： 「我看你如 基列 ， 如 黎巴嫩 的山頂； 然而，我必使你變為曠野， 成為無人居住的城鎮。
JER|22|7|我要預備施行毀滅的人， 各人佩帶兵器攻擊你； 他們要砍伐你佳美的香柏樹， 扔在火中。
JER|22|8|「許多國的百姓經過這城，就彼此談論說：『耶和華為何向這大城這樣做呢？』
JER|22|9|必有人回答說：『是因他們離棄了耶和華－他們上帝的約，事奉敬拜別神。』」
JER|22|10|不要為已死的人哀哭， 也不要為他悲傷， 卻要為離家外出的人大大哀哭； 因為他不再回來見自己的出生地。
JER|22|11|因為論到離開這地方的 約西亞 之子 猶大 王 沙龍 ，就是接續他父親 約西亞 作王的，耶和華這樣說：「他必不再回到這裏來，
JER|22|12|卻要死在被擄去的地方，必不得再見這地。」
JER|22|13|禍哉！那以不公義蓋房，以不公平造樓， 白白使鄰舍做工，卻不給工錢的人，
JER|22|14|他說：「我要為自己蓋寬敞的房，蓋高大的樓。」 他為它開窗戶， 以香柏木為牆板， 漆上丹紅色。
JER|22|15|難道你作王就是要蓋香柏木樓房爭勝的嗎？ 你的父親豈不是也吃也喝， 也施行公平和公義嗎？ 那時他得了福樂。
JER|22|16|他為困苦和貧窮的人伸冤， 那時就得了福樂。 認識我不就在此嗎？ 這是耶和華說的。
JER|22|17|你的眼和你的心卻專顧不義之財， 流無辜人的血， 行欺壓和殘暴。
JER|22|18|所以，耶和華論到 約西亞 的兒子 猶大 王 約雅敬 如此說： 人必不為他舉哀： 「哀哉，我的哥哥！ 哀哉，我的姊姊！」 也不為他舉哀： 「哀哉，我的主！ 哀哉，我主的榮華！」
JER|22|19|他被埋葬好像埋驢子一樣， 被拖出去，扔在 耶路撒冷 城門外。
JER|22|20|你要上 黎巴嫩 哀號， 在 巴珊 揚聲， 從 亞巴琳 哀號， 因為你所親愛的都毀滅了。
JER|22|21|你興盛的時候，我對你說話； 你卻說：「我不聽。」 你從年輕時就是這樣， 不肯聽我的話。
JER|22|22|你的牧人要被風吞吃， 你所親愛的必被擄去； 那時你必因你一切的惡行抱愧蒙羞。
JER|22|23|你這住 黎巴嫩 、在香柏樹上搭窩的， 有痛苦臨到你， 如疼痛臨到臨產的婦人， 那時你何等可憐 ！
JER|22|24|耶和華說：「 約雅敬 的兒子 猶大 王 哥尼雅 ，雖是我右手上帶印的戒指，我憑我的永生起誓，我必將你從其上摘下來。
JER|22|25|我要將你交在尋索你命的人和你所懼怕的人手中，就是 巴比倫 王 尼布甲尼撒 和 迦勒底 人手中。
JER|22|26|我也要將你和生你的母親趕到別國，不是你們出生的地方；你們必死在那裏，
JER|22|27|心中雖然很想歸回那地，卻不得歸回。」
JER|22|28|哥尼雅 這人是被輕看、遭毀壞的罐子， 是無人喜愛的器皿嗎？ 他和他的後裔為何被趕到素不認識之地呢？
JER|22|29|地啊，地啊，地啊，當聽耶和華的話！
JER|22|30|耶和華如此說： 「要把這人登記為無子， 是平生不得亨通的人； 因為他後裔中再無一人得亨通， 能坐在 大衛 的寶座上治理 猶大 。」
JER|23|1|耶和華說：「禍哉！那些殘害、趕散我草場之羊的牧人！」
JER|23|2|耶和華－ 以色列 的上帝論到那些牧養他百姓的牧人如此說：「你們趕散我的羊群，並未看顧他們；看哪，我必懲罰你們的惡行。這是耶和華說的。
JER|23|3|我要從我趕他們到的各國召集我羊群中剩餘的，領他們歸回本處；他們必生養眾多。
JER|23|4|我必設立牧人照管他們，牧養他們。他們不再懼怕，不再驚惶，沒有一個失喪的。這是耶和華說的。
JER|23|5|「看哪，日子將到，我要為 大衛 興起公義的苗裔； 他必掌王權，行事有智慧，在地上施行公平和公義。這是耶和華說的。
JER|23|6|在他的日子， 猶大 必得救， 以色列 也安然居住。他的名必稱為『耶和華－我們的義』。
JER|23|7|「看哪，日子將到，人必不再指著那領 以色列 人從 埃及 地上來的永生耶和華起誓。這是耶和華說的。
JER|23|8|人卻要指著那領 以色列 家的後裔離開北方之地、離開我趕他們到的各國的永生耶和華起誓。他們必住在本地。」
JER|23|9|論到那些先知， 我心在我裏面憂傷， 我的骨頭全都發顫； 因耶和華和他的聖言， 我像醉酒的人， 像被酒所勝的人。
JER|23|10|全地滿了犯姦淫的人！ 因妄自賭咒，地就悲哀， 曠野的草場都枯乾了。 他們所行的道是惡的； 他們的權力用得不對。
JER|23|11|連先知帶祭司都是褻瀆的， 就是在我殿中，我也看見他們的惡行。 這是耶和華說的。
JER|23|12|因此，他們的道路必像黑暗中的滑地， 他們必被追趕，仆倒在其上； 因為在他們受罰之年， 我必使災禍臨到他們。 這是耶和華說的。
JER|23|13|我在 撒瑪利亞 的先知中曾見狂妄的事； 他們藉 巴力 說預言， 使我的百姓 以色列 走迷了路。
JER|23|14|我在 耶路撒冷 的先知中曾見恐怖的事； 他們犯姦淫，行虛謊， 又堅固惡人的手， 無人回轉離開自己的惡行。 他們在我面前都像 所多瑪 ， 耶路撒冷 的居民都像 蛾摩拉 。
JER|23|15|因此，萬軍之耶和華論到先知如此說： 「看哪，我必使他們吃茵蔯， 喝苦水； 因為褻瀆的事出於 耶路撒冷 的先知，遍及各地。」
JER|23|16|萬軍之耶和華如此說：「你們不要聽這些先知向你們所說的預言。他們使你們成為虛無，所說的異象是出於自己的心，不是出於耶和華的口。
JER|23|17|他們常對藐視我的人說：『耶和華說：你們必享平安。』 又對一切按自己頑梗之心而行的人說：『災禍必不臨到你們。』」
JER|23|18|有誰站在耶和華的會中 察看並聽見他的話呢？ 有誰留心聽他的話呢？
JER|23|19|看哪！耶和華的暴風 在震怒中發出， 是旋轉的暴風， 必轉到惡人頭上。
JER|23|20|耶和華的怒氣必不轉消， 直到他心中所定的成就了，實現了。 末後的日子，你們要全然明白。
JER|23|21|我並未差遣那些先知， 他們竟自奔跑； 我沒有對他們說話， 他們竟自預言。
JER|23|22|他們若站在我的會中， 必使我的百姓聽我的話， 又使他們回轉離開惡道， 離開他們所行的惡。
JER|23|23|我是靠近你們的上帝，不是遙遠的上帝，不是嗎？ 這是耶和華說的。
JER|23|24|人豈能在隱密處藏身，使我看不見他呢？這是耶和華說的。我豈不遍滿天和地嗎？這是耶和華說的。
JER|23|25|我已聽見那些先知所說的，他們託我的名說假預言：「我做了夢！我做了夢！」
JER|23|26|所言虛假、心存詭詐的先知，他們這樣存心要到幾時呢？
JER|23|27|他們彼此述說所做的夢，想要使我的百姓忘記我的名，正如他們祖先因 巴力 忘記我的名一樣。
JER|23|28|得夢的先知可以述說那夢；領受我話的人可以誠實講我的話。糠秕怎能與麥子比較呢？這是耶和華說的。
JER|23|29|我的話豈不像火，又像能打碎磐石的大錘嗎？這是耶和華說的。
JER|23|30|看哪，那些先知各從鄰舍偷竊我的話，因此我必與他們為敵。這是耶和華說的。
JER|23|31|那些先知用自己的舌頭說是耶和華說的；看哪，我必與他們為敵。這是耶和華說的。
JER|23|32|那些以假夢為預言，又述說這夢，以謊言和魯莽使我百姓走迷了路的，看哪，我必與他們為敵。這是耶和華說的。我並未差遣他們，也沒有吩咐他們。他們對這百姓毫無益處。這是耶和華說的。
JER|23|33|無論是這百姓、是先知、是祭司，問你說：「耶和華有甚麼默示呢？」你就對他們說：「甚麼默示啊？ 我已撇棄你們了。這是耶和華說的。」
JER|23|34|凡說「耶和華的默示」的，無論是先知、是祭司、是百姓，我必懲罰那人和他的家。
JER|23|35|你們各人要對鄰舍、對弟兄如此說：「耶和華回答了甚麼？耶和華說了甚麼呢？」
JER|23|36|你們不可再提「耶和華的默示」，因為各人所說的話必成為自己的重擔 ；你們錯用了永生上帝、萬軍之耶和華－我們上帝的話。
JER|23|37|你們要對先知如此說：「耶和華回答了你甚麼？耶和華說了甚麼呢？」
JER|23|38|你們若說「耶和華的默示」，耶和華就必如此說：「我曾差人到你們那裏去，告訴你們不可說『耶和華的默示』這幾個字，你們卻說『耶和華的默示』；
JER|23|39|所以，看哪，我必忘記你們 ，將你們和我所賜給你們並你們祖先的城都撇棄了；
JER|23|40|又必使永遠的凌辱和長久的羞恥臨到你們，是不能忘記的。」
JER|24|1|巴比倫 王 尼布甲尼撒 將 約雅敬 的兒子 猶大 王 耶哥尼雅 和 猶大 的領袖，並工匠、鐵匠從 耶路撒冷 擄去，帶到 巴比倫 。這事以後，耶和華指給我看，看哪，有兩筐無花果放在耶和華殿前。
JER|24|2|一筐是極好的無花果，像是初熟的；一筐是極壞的無花果，壞得不能吃。
JER|24|3|耶和華對我說：「 耶利米 ，你看見甚麼？」我說：「我看見無花果，好的極好，壞的極壞，壞得不能吃。」
JER|24|4|於是耶和華的話臨到我，說：
JER|24|5|「耶和華－ 以色列 的上帝如此說：『被擄去的 猶大 人，就是我所打發離開這地到 迦勒底 人之地去的，我必看顧他們如這好的無花果，使他們得福樂。
JER|24|6|我要眷顧他們，使他們得福樂，領他們歸回這地。我也要建立他們，必不拆毀；栽植他們，必不拔出。
JER|24|7|我要賜給他們認識我的心，認識我是耶和華。他們要作我的子民，我要作他們的上帝，他們要一心歸向我。』」
JER|24|8|耶和華如此說：「我必將 猶大 王 西底家 和他的眾領袖，以及留在這地 耶路撒冷 剩餘的人，並住在 埃及 地的 猶大 人都交出來，好像那極壞、壞得不能吃的無花果。
JER|24|9|我必使他們在地上萬國中成為恐懼，成為災禍，在我趕逐他們到的各處成為凌辱、笑柄、譏笑、詛咒的對象。
JER|24|10|我必使刀劍、饑荒、瘟疫臨到他們，直到他們從我所賜給他們和他們祖先之地滅絕。」
JER|25|1|約西亞 的兒子 猶大 王 約雅敬 第四年，就是 巴比倫 王 尼布甲尼撒 的元年，耶和華論 猶大 眾百姓的話臨到 耶利米 。
JER|25|2|耶利米 先知就將這些話對 猶大 眾百姓和 耶路撒冷 所有的居民說：
JER|25|3|「從 亞們 的兒子 猶大 王 約西亞 十三年直到今日，在這二十三年中，常有耶和華的話臨到我；我也一再對你們傳講，只是你們不聽從。
JER|25|4|耶和華也曾一再差遣他的僕人眾先知到你們這裏來，只是你們不聽從，也不側耳而聽，
JER|25|5|說：『你們各人當回轉離開惡道和惡行，就可居住耶和華從古時所賜給你們和你們祖先之地，直到永遠。
JER|25|6|不可隨從別神，事奉敬拜它們，以你們手所做的惹我發怒；這樣，我就不會降災禍給你們。
JER|25|7|然而你們不聽從我，竟以手所做的惹我發怒，害了自己。這是耶和華說的。』」
JER|25|8|所以萬軍之耶和華如此說：「因為你們不聽我的話，
JER|25|9|看哪，我必召北方的眾族和我僕人 巴比倫 王 尼布甲尼撒 前來攻擊這地和這地的居民，並四圍所有的國民。我要將他們盡行滅絕，以致他們令人驚駭、嗤笑，並且永久荒涼 。這是耶和華說的。
JER|25|10|我又要止息他們歡喜和快樂的聲音、新郎和新娘的聲音、推磨的聲音和燈的亮光。
JER|25|11|這全地必然荒涼，令人驚駭。這些國家要服事 巴比倫 王七十年。
JER|25|12|七十年滿了以後，我必懲罰 巴比倫 王和那國，並 迦勒底 人之地，因他們的罪孽使那地永遠荒涼。這是耶和華說的。
JER|25|13|我也必使我向那地所說的話，就是所有記在這書上， 耶利米 向這些國家說的預言，都臨到那地。
JER|25|14|因為必有許多國家和大君王使 迦勒底 人作奴僕；我也必照他們的行為，按他們手所做的報應他們。」
JER|25|15|耶和華－ 以色列 的上帝對我如此說：「你從我手中拿這杯憤怒的酒，給我所差遣你去的各國的百姓喝。
JER|25|16|他們喝了就要東倒西歪，並要發狂，因我使刀劍臨到他們中間。」
JER|25|17|我就從耶和華的手中拿了這杯，給耶和華所差遣我去的各國的百姓喝，
JER|25|18|其中有 耶路撒冷 和 猶大 的城鎮，並 耶路撒冷 的君王與領袖；因此這城鎮荒涼，令人驚駭、嗤笑、詛咒，正如今日一樣。
JER|25|19|又有 埃及 王法老和他的臣僕、官長，以及他的眾百姓，
JER|25|20|並混居的各族和 烏斯 地的諸王，與 非利士 人之地的諸王，包括 亞實基倫 、 迦薩 、 以革倫 ，以及 亞實突 剩下的人，
JER|25|21|還有 以東 、 摩押 、 亞捫 人，
JER|25|22|推羅 的諸王、 西頓 的諸王、海的那邊沿海地區的諸王，
JER|25|23|底但 、 提瑪 、 布斯 ，和所有剃鬢髮的人，
JER|25|24|阿拉伯 的諸王、住曠野混居各族的諸王、
JER|25|25|心利 的諸王、 以攔 的諸王、 瑪代 的諸王、
JER|25|26|北方遠近的諸王，以及天下、地面上的萬國也一個一個都喝了，以後 示沙克 王也要喝。
JER|25|27|「你要對他們說：『萬軍之耶和華－ 以色列 的上帝如此說：你們要喝，且要喝醉，要嘔吐，且要跌倒，不再起來，都因我使刀劍臨到你們中間。』
JER|25|28|「他們若不肯從你手中拿這杯來喝，你就要對他們說：『萬軍之耶和華如此說：你們一定要喝！
JER|25|29|看哪，我既從稱為我名下的城起首施行災禍，你們能免去懲罰嗎？你們必不能免，因為我要命刀劍臨到地上所有的居民。這是萬軍之耶和華說的。』
JER|25|30|「所以你要向他們預言這一切的話，對他們說： 『耶和華從高天吼叫， 從聖所發出聲音， 向自己的羊群大聲吼叫； 他要向地上所有的居民吶喊， 像踹葡萄的人一樣。
JER|25|31|必有響聲達到地極， 因為耶和華與列國爭辯。 凡有血肉之軀的，他必審問； 至於惡人，他必交給刀劍。 這是耶和華說的。』
JER|25|32|「萬軍之耶和華如此說： 看哪，必有災禍發出，從這國到那國， 並有大暴風從地極颳起。
JER|25|33|「到那日，從地這邊到地那邊，都有耶和華所殺戮的人。必無人哀哭，不得收殮，不得埋葬，必在地面上成為糞土。
JER|25|34|「牧人哪，你們當哀號，呼喊； 羊群的領導者啊，你們要在灰中翻滾； 因為你們被宰殺、被分散 的日子已經來到。 你們要仆倒，好像珍貴的器皿打碎一樣。
JER|25|35|牧人無路可逃， 羊群的領導者也無法逃脫。
JER|25|36|聽啊，有牧人呼喊， 有羊群領導者哀號的聲音， 因為耶和華摧毀他們的草場。
JER|25|37|因耶和華猛烈的怒氣， 平安的羊圈都被肅清。
JER|25|38|他像獅子離開洞穴， 他們的地因兇猛的怒氣 和他強烈的怒氣，都變為荒涼。」
JER|26|1|約西亞 的兒子 猶大 王 約雅敬 登基時，有這話從耶和華臨到 耶利米 ，說：
JER|26|2|「耶和華如此說：你要站在耶和華殿的院內，對 猶大 所有城鎮的人，就是到耶和華的殿來禮拜的，傳講我所吩咐你的一切話，一字也不可刪減。
JER|26|3|或者他們肯聽從，各人回轉離開惡道，我就改變心意，不將我因他們所行的惡、想要施行的災禍降與他們。
JER|26|4|你要對他們說，耶和華如此說：『你們若不聽從我，不遵行我在你們面前所設立的律法，
JER|26|5|不聽從我一再差遣我僕人眾先知到你們那裏去所說的話，你們果然沒有聽從，
JER|26|6|我就必使這殿如 示羅 ，使這城成為地上萬國所詛咒的。』」
JER|26|7|耶利米 在耶和華殿中所說的這些話，祭司、先知與眾百姓都聽見了。
JER|26|8|耶利米 說完了耶和華吩咐他對眾百姓說的一切話，祭司、先知與眾百姓都來抓住他，說：「你該死！
JER|26|9|你為何假借耶和華的名預言，說這殿必如 示羅 ，這城必荒廢無人居住呢？」於是眾百姓都聚集在耶和華的殿中圍住 耶利米 。
JER|26|10|猶大 的官長們聽見這些事，就從王宮上到耶和華的殿，坐在耶和華殿 新門 的入口。
JER|26|11|祭司、先知對官長和眾百姓說：「這人該死，因為他說預言攻擊這城，正如你們親耳聽見的。」
JER|26|12|耶利米 就對官長和眾百姓說：「耶和華差遣我預言攻擊這殿和這城，傳講你們所聽見的這一切話。
JER|26|13|現在，要改正你們的所作所為，聽從耶和華－你們上帝的話，他就必改變心意，不把所說的災禍降與你們。
JER|26|14|至於我，看哪，我在你們手中，你們眼裏看甚麼是好的，是正確的，就那樣待我吧！
JER|26|15|但你們要確實知道，你們若把我處死，就使流無辜人血的罪歸給你們和這城，以及城裏的居民了；因為耶和華確實差遣我到你們這裏來，將這一切話傳到你們耳中。」
JER|26|16|官長和眾百姓對祭司和先知說：「這人是不該死的，因為他奉耶和華－我們上帝的名向我們說話。」
JER|26|17|國中的長老就有幾個人起來，對聚集的眾百姓說：
JER|26|18|「當 猶大 王 希西家 的日子，有 摩利沙 人 彌迦 對 猶大 眾百姓預言說： 『萬軍之耶和華如此說： 錫安 要被耕種像一塊田地， 耶路撒冷 要變為廢墟， 這殿的山必像叢林的高處。』
JER|26|19|「 猶大 王 希西家 和 猶大 人豈是把他處死呢？ 希西家 豈不是敬畏耶和華，懇求耶和華施恩嗎？耶和華就改變心意，不把所說的災禍降與他們。若處死這人，我們就做了大惡，害死自己了。」
JER|26|20|有一個人，就是 示瑪雅 的兒子 基列‧耶琳 人 烏利亞 ，也奉耶和華的名說預言；他說預言攻擊這城和這地，和 耶利米 所說的完全一樣。
JER|26|21|約雅敬 王和他所有的勇士、官長聽見了 烏利亞 的話，王想要把他處死。 烏利亞 聽見就懼怕，逃往 埃及 去了。
JER|26|22|約雅敬 王差 亞革波 的兒子 以利拿單 ，帶領幾個人前往 埃及 。
JER|26|23|他們將 烏利亞 從 埃及 帶出來，解送到 約雅敬 王那裏；王用刀殺了他，把他的屍首拋在平民的墳地中。
JER|26|24|然而， 沙番 的兒子 亞希甘 保護 耶利米 ，不將他交在百姓手中，以免他們把他處死。
JER|27|1|約西亞 的兒子 猶大 王 約雅敬 登基時，有這話從耶和華臨到 耶利米 ，說：
JER|27|2|「耶和華對我如此說：你要為自己做皮帶和木軛，套在你的頸項上，
JER|27|3|然後託那些來到 耶路撒冷 ，到 猶大 王 西底家 那裏的使節，把皮帶和木軛送到 以東 王、 摩押 王、 亞捫 王、 推羅 王、 西頓 王那裏，
JER|27|4|且囑咐他們轉達他們的主人。萬軍之耶和華－ 以色列 的上帝如此說，你們要對你們的主人這樣說：
JER|27|5|我用大能和伸出來的膀臂創造大地和地上的人民、牲畜。我看給誰合適，就把地給誰。
JER|27|6|現在我將全地都交在我僕人 巴比倫 王 尼布甲尼撒 手中，也把野地的走獸給他使用。
JER|27|7|列國都要服事他和他的子孫，直到他本國遭報的日期來到；那時，許多國家和大君王要使他作奴隸。
JER|27|8|「無論哪一邦、哪一國，不肯服事 巴比倫 王 尼布甲尼撒 ，不把頸項放在他的軛下，我必用刀劍、饑荒、瘟疫懲罰那邦，直到我藉 巴比倫 王的手毀滅他們。這是耶和華說的。
JER|27|9|至於你們，不可聽從你們的先知和占卜的、做夢的 、觀星象的，以及行邪術的；他們對你們說：『你們必不致服事 巴比倫 王。』
JER|27|10|他們向你們傳的是假預言，要叫你們遠離本地，以致我將你們趕出去，使你們滅亡。
JER|27|11|但哪一邦肯把頸項放在 巴比倫 王的軛下服事他，我必使那邦仍在本地存留，在那裏耕種居住。這是耶和華說的。」
JER|27|12|我就照這一切話對猶大王 西底家 說：「你們要把頸項放在 巴比倫 王的軛下，服事他和他的百姓，就得存活。
JER|27|13|你和你的百姓何必因刀劍、饑荒、瘟疫而死亡，像耶和華所論不肯服事 巴比倫 王的國家呢？
JER|27|14|不可聽那些先知對你們所說的話，他們說：『你們必不致服事 巴比倫 王』，其實他們向你們傳的是假預言。
JER|27|15|耶和華說：『我並未差遣他們，他們卻託我的名傳假預言，使我將你們和向你們說預言的那些先知趕出去，一同滅亡。』」
JER|27|16|我又對祭司和這眾百姓說：「耶和華如此說：你們不可聽那先知對你們所說的預言，他們說：『看哪，耶和華殿中的器皿快要從 巴比倫 帶回來』；其實他們向你們傳的是假預言。
JER|27|17|不可聽從他們，只管服事 巴比倫 王，就得存活。何必使這城變為廢墟呢？
JER|27|18|他們若真是先知，有耶和華的話臨到他們，讓他們祈求萬軍之耶和華，使耶和華殿中和 猶大 王宮內，並 耶路撒冷 剩下的器皿，不致被帶到 巴比倫 去。
JER|27|19|萬軍之耶和華這樣論柱子、銅海、盆座，並留在這城裏剩下的器皿，
JER|27|20|就是 巴比倫 王 尼布甲尼撒 擄掠 約雅敬 的兒子 猶大 王 耶哥尼雅 ，並 猶大 、 耶路撒冷 所有貴族時，沒有從 耶路撒冷 掠去 巴比倫 的器皿。
JER|27|21|論到那在耶和華殿中和 猶大 王宮內，並 耶路撒冷 剩下的器皿，萬軍之耶和華－ 以色列 的上帝如此說：
JER|27|22|它們必被帶到 巴比倫 ，存放在那裏，直到我眷顧 以色列 人，將這些器皿帶回歸還此地的日子。這是耶和華說的。」
JER|28|1|當年，就是 猶大 王 西底家 登基第四年五月， 押朔 的兒子 基遍 人 哈拿尼雅 先知，在耶和華的殿中當著祭司和眾百姓的面對我說：
JER|28|2|「萬軍之耶和華－ 以色列 的上帝如此說：我已經折斷 巴比倫 王的軛。
JER|28|3|二年之內，我要將 巴比倫 王 尼布甲尼撒 從這地擄掠到 巴比倫 的器皿，就是耶和華殿中的一切器皿，都帶回此地。
JER|28|4|我又要將 約雅敬 的兒子 猶大 王 耶哥尼雅 和被擄到 巴比倫 所有的 猶大 人帶回此地，因為我要折斷 巴比倫 王的軛。這是耶和華說的。」
JER|28|5|耶利米 先知當著祭司和站在耶和華殿裏眾百姓的面，對 哈拿尼雅 先知說：
JER|28|6|「阿們！願耶和華如此行，願耶和華實現你所預言的話，將耶和華殿中的器皿和所有被擄去的人從 巴比倫 帶回此地。
JER|28|7|然而我在你和眾百姓耳中所要說的話，你應當聽。
JER|28|8|從古以來，在你我以前的眾先知，向多國和大邦說預言，論到戰爭、災禍 、瘟疫的事。
JER|28|9|至於那預言平安的先知，到先知的話應驗的時候，人就知道他真是耶和華所差來的。」
JER|28|10|哈拿尼雅 先知就取下 耶利米 先知頸項上的軛，把它折斷。
JER|28|11|哈拿尼雅 又當著眾百姓的面說：「耶和華如此說：二年之內我必照樣從列國的頸項上折斷 巴比倫 王 尼布甲尼撒 的軛。」 耶利米 先知就離開了。
JER|28|12|哈拿尼雅 先知折斷 耶利米 先知頸項上的軛以後，耶和華的話臨到 耶利米 ，說：
JER|28|13|「你去告訴 哈拿尼雅 說，耶和華如此說：你折斷木軛，卻換來鐵軛！
JER|28|14|萬軍之耶和華－ 以色列 的上帝如此說：我已將鐵軛加在這些國的頸項上，使他們服事 巴比倫 王 尼布甲尼撒 。他們總要服事他，我也把野地的走獸給了他。」
JER|28|15|於是 耶利米 先知對 哈拿尼雅 先知說：「 哈拿尼雅 啊，你應當聽！耶和華並沒有差遣你，你竟使這百姓倚靠謊言。
JER|28|16|所以耶和華如此說：看哪，我要把你從地面上除掉，你今年必死，因為你向耶和華說了叛逆的話。」
JER|28|17|這樣， 哈拿尼雅 先知當年七月間就死了。
JER|29|1|耶利米 先知從 耶路撒冷 送信給被擄倖存的長老，以及祭司、先知，和 尼布甲尼撒 從 耶路撒冷 擄到 巴比倫 去的眾百姓。
JER|29|2|這是在 耶哥尼雅 王和太后、官員，並 猶大 和 耶路撒冷 的領袖，以及工匠、鐵匠都離開 耶路撒冷 之後。
JER|29|3|他藉 沙番 的兒子 以利亞薩 和 希勒家 的兒子 基瑪利 的手送去；他們二人是 猶大 王 西底家 差往 巴比倫 去見 巴比倫 王 尼布甲尼撒 的。
JER|29|4|信上說：「萬軍之耶和華－ 以色列 的上帝對所有被擄的，就是我使他們從 耶路撒冷 被擄到 巴比倫 去的人如此說：
JER|29|5|你們要建造房屋，住在其中；要開墾田園，吃園中所出產的；
JER|29|6|要娶妻生兒養女，為你們的兒子娶妻，使你們的女兒嫁人，生兒養女。你們要在那裏生養眾多，不可減少。
JER|29|7|我使你們被擄到的那城，你們要為那城求平安，為那城向耶和華祈求，因為那城得平安，你們也隨著得平安。
JER|29|8|萬軍之耶和華－ 以色列 的上帝如此說：不要被你們中間的先知和占卜的所誘惑，也不要聽信你們 所做的夢，
JER|29|9|因為他們託我的名對你們說假預言，我並未差遣他們。這是耶和華說的。
JER|29|10|「耶和華如此說：為 巴比倫 所定的七十年滿了以後，我要眷顧你們，向你們實現我的恩言，使你們歸回此地。
JER|29|11|我知道我向你們所懷的意念是賜平安的意念，不是降災禍的意念，要叫你們末後有指望。這是耶和華說的。
JER|29|12|你們呼求我，向我禱告，我就應允你們。
JER|29|13|你們尋求我，若專心尋求我，就必尋見。
JER|29|14|我必被你們尋見，也必使你們被擄的人歸回。這是耶和華說的。我必將你們從各國和我趕你們到的各處召集過來，又將你們帶回我使你們被擄離開的地方。這是耶和華說的。
JER|29|15|「你們說：『耶和華已在 巴比倫 為我們興起先知。』
JER|29|16|所以耶和華如此論坐 大衛 寶座的君王和住在這城裏所有的百姓，就是未曾與你們一同被擄的弟兄，
JER|29|17|萬軍之耶和華如此說：『看哪，我必使刀劍、饑荒、瘟疫臨到他們，使他們像極壞的無花果，壞得不能吃。
JER|29|18|我必用刀劍、饑荒、瘟疫追趕他們，使地上萬國因他們而驚駭；在我趕他們到的各國，令人詛咒、驚駭、嗤笑、羞辱。
JER|29|19|這是因為他們不聽從我先前一再差遣我僕人眾先知說的話。這是耶和華說的。你們 也一樣不聽。這是耶和華說的。』
JER|29|20|所以你們所有被擄去的，就是我從 耶路撒冷 放逐到 巴比倫 去的，當聽耶和華的話。
JER|29|21|萬軍之耶和華－ 以色列 的上帝論 哥賴雅 的兒子 亞哈 和 瑪西雅 的兒子 西底家 如此說：『他們託我的名向你們說假預言，看哪，我必把他們交在 巴比倫 王 尼布甲尼撒 的手中，他要在你們眼前殺害他們。
JER|29|22|在 巴比倫 所有被擄的 猶大 人必藉這二人賭咒說：願耶和華使你像 巴比倫 王在火中焚燒的 西底家 和 亞哈 一樣。
JER|29|23|這二人在 以色列 中做了醜事，與鄰舍的妻行淫，又假託我的名說我未曾吩咐他們的話。我知道這一切，也作見證。這是耶和華說的。』」
JER|29|24|「你要對 尼希蘭 人 示瑪雅 說：
JER|29|25|萬軍之耶和華－ 以色列 的上帝如此說：你曾用自己的名送信給 耶路撒冷 的眾百姓和 瑪西雅 的兒子 西番雅 祭司，並眾祭司，說：
JER|29|26|『耶和華已經立你 西番雅 為祭司，代替 耶何耶大 祭司，使耶和華的殿中有總管，好把所有狂妄自稱先知的人用枷枷住，用鎖鎖住。
JER|29|27|現在 亞拿突 人 耶利米 向你們自稱先知，你為甚麼不責備他呢？
JER|29|28|他送信給我們在 巴比倫 的人說：被擄的事必長久，你們要建造房屋，住在其中；要開墾田園，吃園中所出產的。』」
JER|29|29|西番雅 祭司就把這信念給 耶利米 先知聽。
JER|29|30|於是耶和華的話臨到 耶利米 ，說：
JER|29|31|「你當送信給所有被擄的人，說：『耶和華論到 尼希蘭 人 示瑪雅 說：因為 示瑪雅 向你們說預言，使你們倚靠謊言，而我並沒有差遣他，
JER|29|32|所以耶和華如此說：看哪，我必懲罰 尼希蘭 人 示瑪雅 和他的後裔，他必無一人存留住在這民中，也看不見我所要賞賜給我百姓的福樂，因為他向耶和華說了叛逆的話。這是耶和華說的。』」
JER|30|1|耶和華的話臨到 耶利米 ，說：
JER|30|2|「耶和華－ 以色列 的上帝如此說：你要將我對你說過的一切話都寫在書上。
JER|30|3|看哪，日子將到，我要使我的百姓 以色列 和 猶大 被擄的人歸回。這是耶和華說的。耶和華說：我要使他們回到我所賜給他們祖先之地，他們就得這地為業。」
JER|30|4|以下是耶和華論到 以色列 和 猶大 所說的話：
JER|30|5|耶和華如此說： 「我們聽見顫抖的聲音， 令人懼怕，沒有平安。
JER|30|6|你們且訪查看看， 男人會生孩子嗎？ 我怎麼看見人人都用手撐腰， 像臨產的婦人， 臉都發白了呢？
JER|30|7|哀哉！ 那日為大， 無日可比； 這是 雅各 遭難的時刻， 但他必從患難中得拯救。」
JER|30|8|萬軍之耶和華說：「到那日，我必折斷你頸項上仇敵的軛，拉斷你的皮帶。陌生人必不再使他作奴隸。
JER|30|9|他們卻要事奉耶和華－他們的上帝，事奉我為他們所興起的 大衛 王。」
JER|30|10|我的僕人 雅各 啊，不要懼怕； 以色列 啊，不要驚惶； 因我從遠方拯救你， 從被擄之地拯救你的後裔； 雅各 必回來得享平靜安逸， 無人能使他害怕。 這是耶和華說的。
JER|30|11|因我與你同在，要拯救你， 也要將那些國滅絕淨盡， 就是我趕你去的那些國； 卻不將你滅絕淨盡， 倒要從寬懲治你， 但絕不能不罰你。 這是耶和華說的。
JER|30|12|耶和華如此說： 「你的損傷無法醫治， 你的傷痕極其重大。
JER|30|13|無人為你的傷痛辯護， 也沒有可醫治你的良藥。
JER|30|14|你所親愛的都忘記你， 不來探望你。 我因你罪孽甚大，罪惡眾多， 曾藉仇敵加的傷害傷害你， 藉殘忍者懲治你。
JER|30|15|你為何因所受的損傷哀號呢？ 你的痛苦無法醫治。 我因你罪孽甚大，罪惡眾多， 曾將這些加在你身上。
JER|30|16|因此，凡吞吃你的必被吞吃， 你的敵人個個都被擄去； 擄掠你的必成為擄物， 我使搶奪你的成為掠物。
JER|30|17|我必使你痊癒， 醫好你的傷痕， 都因人稱你為被趕散的， 這是 錫安 ，是無人來探望的！ 這是耶和華說的。」
JER|30|18|耶和華如此說： 「看哪，我必使 雅各 被擄去的帳棚歸回， 也必顧惜他的住處。 城必建造在原有的廢墟上， 宮殿也必照樣有人居住。
JER|30|19|必有感謝和歡樂的聲音從其中發出， 我使他們增多，不致減少； 使他們尊榮，不致卑微。
JER|30|20|他們的兒女必如往昔； 他們的會眾堅立在我面前； 凡欺壓他們的，我必懲罰。
JER|30|21|他們的君王是他們自己的人， 掌權的必出自他們。 我要使他接近我， 他也要親近我； 不然，誰敢放膽親近我呢？ 這是耶和華說的。
JER|30|22|你們要作我的子民， 我要作你們的上帝。」
JER|30|23|看哪，耶和華的憤怒 如暴風已經發出； 是掃滅的暴風， 必轉到惡人的頭上。
JER|30|24|耶和華的烈怒必不轉消， 直到他心中所定的成就了，實現了； 末後的日子你們就會明白。
JER|31|1|耶和華說：「那時，我必作 以色列 各家的上帝，他們必作我的子民。」
JER|31|2|耶和華如此說： 「從刀劍生還的百姓 在曠野蒙恩； 以色列 尋找安歇之處。」
JER|31|3|耶和華從遠方向我顯現： 「我以永遠的愛愛你， 因此，我以慈愛吸引你。」
JER|31|4|少女 以色列 啊， 我要再建立你，你就得以建立； 你必再拿起手鼓， 隨著歡樂的舞者而出。
JER|31|5|你必在 撒瑪利亞 的山上栽葡萄園， 栽種的人栽種，而且享用。
JER|31|6|日子將到，守望的人必在 以法蓮 山上呼叫： 「起來吧！我們要上 錫安 ， 到耶和華－我們的上帝那裏去。」
JER|31|7|耶和華如此說： 「你們當為 雅各 歡樂歌唱， 為萬國中為首的歡呼。 當傳揚，頌讚說： 『耶和華啊， 求你拯救你的百姓 ， 拯救 以色列 的餘民。』
JER|31|8|看哪，我必將他們從北方之地領來， 從地極召集而來； 同他們來的有盲人、瘸子、孕婦、產婦； 他們必成群結隊回到這裏。
JER|31|9|他們要哭泣而來。 我要照他們懇求的引導他們， 使他們在河水旁行走正直的路， 他們在其上必不致絆跌； 因為我是 以色列 的父， 以法蓮 是我的長子。
JER|31|10|列國啊，要聽耶和華的話， 要在遠方的海島傳揚，說： 「趕散 以色列 的必召集他， 看守他，如牧人看守羊群。」
JER|31|11|因為耶和華救贖了 雅各 ， 救贖他脫離比他更強之人的手。
JER|31|12|他們來到 錫安 的高處歌唱， 因耶和華的宏恩而喜樂洋溢， 就是五穀、新酒和新的油， 並羔羊和牛犢。 他們必像有水澆灌的園子， 一點也不再有愁煩。
JER|31|13|那時，少女必歡樂跳舞； 年輕的、年老的，都一同歡樂； 因為我要使他們的悲哀變為歡喜， 並要安慰他們，使他們的愁煩轉為喜樂。
JER|31|14|我必以肥油使祭司的心滿足， 我的百姓也要因我的恩惠知足。 這是耶和華說的。
JER|31|15|耶和華如此說： 「在 拉瑪 聽見號咷痛哭的聲音， 是 拉結 哭她兒女，不肯因她兒女受安慰， 因為他們都不在了。」
JER|31|16|耶和華如此說： 「不要出聲哀哭， 你的眼目也不要流淚； 因你的辛勞必有報償， 他們必從仇敵之地歸回。 這是耶和華說的。
JER|31|17|你末後必有指望， 你的兒女必回到自己的疆土。 這是耶和華說的。
JER|31|18|我聽見 以法蓮 為自己悲嘆說： 『你管教我，我便受管教， 我如未馴服的牛犢。 求你使我回轉，我便回轉， 因為你是耶和華－我的上帝。
JER|31|19|我背離以後就懊悔， 受教以後就捶胸 ； 我因擔當年輕時的凌辱就抱愧蒙羞。』
JER|31|20|以法蓮 是我的愛子嗎？ 是我喜歡的孩子嗎？ 我每逢責備他，仍深顧念他。 因此，我的心腸牽掛著他， 我必要憐憫他。 這是耶和華說的。
JER|31|21|少女 以色列 啊， 當為自己設立路標， 為自己豎起指路牌。 要留心向著大道， 就是你曾走過的路； 你當回轉，回到你自己的城鎮。
JER|31|22|背道的女子啊， 你翻來覆去要到幾時呢？ 耶和華在地上造了一件新事， 就是女子護衛男子。」
JER|31|23|萬軍之耶和華－ 以色列 的上帝如此說：「我使被擄之人歸回的時候，他們在 猶大 地和其中的城鎮必再這樣說： 公義的居所啊，聖山哪， 願耶和華賜福給你。
JER|31|24|猶大 和 猶大 城鎮的人，耕地的和帶著群畜遊牧的人，都要一同住在其中。
JER|31|25|疲乏的人，我使他振作；愁煩的人，我使他滿足。」
JER|31|26|於是我醒了，我看到我睡得香甜。
JER|31|27|「看哪，日子將到，我要使人的後代和牲畜的種，在 以色列 家和 猶大 家繁衍。這是耶和華說的。
JER|31|28|我先前怎樣看守他們，為要拔出、拆毀、毀壞、傾覆、苦害，也必照樣看守他們，為要建立、栽植。這是耶和華說的。
JER|31|29|當那些日子，人不再說： 『父親吃了酸葡萄， 兒子牙齒就酸倒。』
JER|31|30|但各人要因自己的罪死亡；凡吃酸葡萄的，自己的牙必酸倒。
JER|31|31|「看哪，日子將到，我要與 以色列 家和 猶大 家另立新的約。這是耶和華說的。
JER|31|32|這約不像我拉著他們祖宗的手，領他們出 埃及 地的時候與他們所立的約。我雖作他們的丈夫，他們卻背了我的約。這是耶和華說的。
JER|31|33|那些日子以後，我與 以色列 家所立的約是這樣：我要將我的律法放在他們裏面，寫在他們心上。我要作他們的上帝，他們要作我的子民。這是耶和華說的。
JER|31|34|他們各人不再教導自己的鄰舍和弟兄說：『你該認識耶和華』，因為他們從最小的到最大的都必認識我。我要赦免他們的罪孽，不再記得他們的罪惡。這是耶和華說的。」
JER|31|35|耶和華使太陽白晝發光， 按定例使月亮和星辰照耀黑夜， 又攪動大海，使海中波浪澎湃， 萬軍之耶和華是他的名， 他如此說：
JER|31|36|「這些定例若能在我面前廢掉， 以色列 的後裔才會在我面前斷絕， 永遠不再成國。 這是耶和華說的。」
JER|31|37|耶和華如此說： 「若有人能測量上面的天， 探索下面地的根基， 我才會因 以色列 後裔所做的一切棄絕他們。 這是耶和華說的。」
JER|31|38|看哪，日子將到，這城必為耶和華而造，從 哈楠業樓 直到 角門 。這是耶和華說的。
JER|31|39|丈量的繩子要往外拉出，直到 迦立山 ，又轉到 歌亞 ；
JER|31|40|拋屍的全谷和倒灰之處，並一切田地，直到 汲淪溪 ，又到東邊 馬門 的角落，都要歸耶和華為聖；不再拔出，不再傾覆，直到永遠。
JER|32|1|猶大 王 西底家 第十年，就是 尼布甲尼撒 十八年，耶和華的話臨到 耶利米 。
JER|32|2|那時 巴比倫 王的軍隊圍困 耶路撒冷 ， 耶利米 先知被囚在 猶大 王宮中護衛兵的院內；
JER|32|3|因為 猶大 王 西底家 囚禁他，說：「你為甚麼預言耶和華如此說：『看哪，我要把這城交在 巴比倫 王的手中，他必攻下這城。
JER|32|4|猶大 王 西底家 必不能逃脫 迦勒底 人的手，定要交在 巴比倫 王手中，他要親眼看到 巴比倫 王，親口跟他說話。
JER|32|5|巴比倫 王要將 西底家 帶到 巴比倫 ； 西底家 必住在那裏，直到我懲罰 他的時候。你們雖與 迦勒底 人爭戰，卻不順利。這是耶和華說的。』」
JER|32|6|耶利米 說：「耶和華的話臨到我，說：
JER|32|7|『看哪，你叔父 沙龍 的兒子 哈拿篾 必到你這裏來，說：請你買我在 亞拿突 的那塊地，因為你有代贖的責任。』
JER|32|8|我叔父的兒子 哈拿篾 果然照耶和華的話來到護衛兵的院內，對我說：『請你買我在 便雅憫 境內、 亞拿突 的那塊地；因為它應該由你來承受，而且你也有代贖的責任。請你買下它吧！』我就知道這確是耶和華的話。
JER|32|9|「我便向我叔父的兒子 哈拿篾 買了 亞拿突 的那塊地，秤了十七舍客勒銀子給他。
JER|32|10|我在契上簽字，將契封緘，又請證人來，用天平把銀子秤給他。
JER|32|11|我又將按照法定條例所立的買契，就是封緘的那一張和敞開的那一張，
JER|32|12|在我叔父的兒子 哈拿篾 和簽字作證的人，並坐在護衛兵院內所有 猶大 人眼前，交給 瑪西雅 的孫子 尼利亞 的兒子 巴錄 。
JER|32|13|我在眾人眼前囑咐 巴錄 說：
JER|32|14|『萬軍之耶和華－ 以色列 的上帝如此說：你拿著這文件，就是封緘的和敞開的買契，把它們放在瓦器裏，以便長久保存。
JER|32|15|因為萬軍之耶和華－ 以色列 的上帝如此說：將來在這地必有人再購置房屋、田地和葡萄園。』」
JER|32|16|「我將買契交給 尼利亞 的兒子 巴錄 以後，就向耶和華禱告說：
JER|32|17|『唉！主耶和華，看哪，你曾用大能和伸出來的膀臂創造天和地，在你沒有難成的事。
JER|32|18|你施慈愛給千萬人，又將祖先的罪孽報應在他後世子孫身上。至大全能的上帝啊，萬軍之耶和華是你的名，
JER|32|19|你謀事有大略，行事有大能，注目觀看世人一切的舉動，為要照各人所做的和他做事的結果報應他。
JER|32|20|你在 埃及 地顯神蹟奇事，直到今日在 以色列 和世人中間也是如此，建立了自己的名聲，正如今日一樣。
JER|32|21|你用神蹟奇事、大能的手、伸出來的膀臂和大可畏的事，領你的百姓 以色列 出了 埃及 ，
JER|32|22|把這地賞賜給他們，就是你向他們列祖起誓應許要賜給他們的流奶與蜜之地。
JER|32|23|他們進入並取得這地，卻不聽從你的話，也不遵行你的律法。你吩咐他們所當行的，他們都不去行，因此你使這一切的災禍臨到他們。
JER|32|24|看哪，敵人已經來到，用土堆攻取這城；這城也因刀劍、饑荒、瘟疫被交在攻城的 迦勒底 人手中。你所說的話都應驗了，看哪，你也看見了。
JER|32|25|主耶和華啊，你卻對我說，要用銀子為自己買那塊地，又請人作證；其實這城已交在 迦勒底 人的手中了。』」
JER|32|26|耶和華的話臨到 耶利米 ，說：
JER|32|27|「看哪，我是耶和華，是凡有血肉之軀者的上帝，在我豈有難成的事嗎？
JER|32|28|耶和華如此說：看哪，我必將這城交給 迦勒底 人的手和 巴比倫 王 尼布甲尼撒 的手，他必攻取這城。
JER|32|29|攻城的 迦勒底 人必來放火焚燒這城和城裏的房屋；人曾在這房頂上向 巴力 燒香，向別神獻澆酒祭，惹我發怒。
JER|32|30|以色列 人和 猶大 人從年輕時，就專做我眼中看為惡的事。 以色列 人盡以手所做的惹我發怒。這是耶和華說的。
JER|32|31|這城自從建造的那日直到今日，常惹我的怒氣和憤怒，以致我將這城從我面前除掉；
JER|32|32|這是因 以色列 人和 猶大 人一切的邪惡，就是他們和他們的君王、官長、祭司、先知，並 猶大 人，以及 耶路撒冷 居民所做的，惹我發怒。
JER|32|33|他們以背向我，不以面向我；我雖然一再教導他們，他們卻不聽從，不領受訓誨，
JER|32|34|竟把可憎之偶像設立在稱為我名下的殿中，玷污了這殿。
JER|32|35|他們在 欣嫩子谷 建造 巴力 的丘壇，把自己的兒女經火獻給 摩洛 ；他們行這可憎的事，使 猶大 陷在罪裏，這並不是我吩咐的，我心裏也從來沒有想過。」
JER|32|36|現在論到這城，就是你們所說，已經因刀劍、饑荒、瘟疫被交在 巴比倫 王手中的，耶和華－ 以色列 的上帝如此說：
JER|32|37|「看哪，我曾在怒氣、憤怒和大惱怒中，將 以色列 人趕到各國；我必從那裏將他們召集出來，領他們回到此地，使他們安然居住。
JER|32|38|他們要作我的子民，我要作他們的上帝。
JER|32|39|我要使他們彼此同心同道，好叫他們永遠敬畏我，使他們和他們後世的子孫得享福樂。
JER|32|40|我要跟他們立永遠的約，要施恩給他們，絕不轉離；又要把敬畏我的心放在他們心裏，不離棄我。
JER|32|41|我必歡喜施恩給他們，盡心盡意、真誠地將他們栽於此地。
JER|32|42|「因為耶和華如此說：我怎樣使這一切大災禍臨到這百姓，也要照樣使我所應許他們的一切福樂都臨到他們。
JER|32|43|你們所說荒涼、無人、無牲畜，已交給 迦勒底 人手的這地，必有人購置田地。
JER|32|44|在 便雅憫 地、 耶路撒冷 四圍的各處、 猶大 的城鎮、山區的城鎮、 謝非拉 的城鎮，並 尼革夫 的城鎮，人必用銀子買田地，在契上簽字，將契封緘，找人作證，因為我必使被擄的人歸回。這是耶和華說的。」
JER|33|1|耶利米 還囚在護衛兵的院內，耶和華的話第二次臨到他，說：
JER|33|2|「成事的耶和華，塑造它為要建立它的耶和華，名為耶和華的那位如此說：
JER|33|3|『你求告我，我就應允你，並將你所不知道、又大又隱密的事指示你。
JER|33|4|論到這城中的房屋和 猶大 君王的宮殿，就是拆毀來擋圍城工事和刀劍的，耶和華－ 以色列 的上帝如此說：
JER|33|5|他們與 迦勒底 人爭戰，用我在怒氣和憤怒中所殺之人的屍首塞滿這房屋；我因他們一切的惡，轉臉不顧這城。
JER|33|6|看哪，我要使這城得以痊癒安舒，我要醫治他們，將豐盛的平安與信實顯明給他們。
JER|33|7|我也要使 猶大 被擄的和 以色列 被擄的人歸回，並要建立他們，如起初一樣。
JER|33|8|我要洗淨他們干犯我的一切罪，赦免他們干犯我、違背我的一切罪。
JER|33|9|這城在地上萬國面前要因我的緣故，以喜樂得名，得頌讚，得榮耀，因為他們聽見我所賞賜的一切福樂。他們因我向這城所施的一切福樂平安，就懼怕戰兢。」
JER|33|10|耶和華如此說：「你們論這地方，說是荒廢、無人、無牲畜之地，但在這荒涼、無人、無居民、無牲畜的 猶大 城鎮和 耶路撒冷 街上，必再聽見
JER|33|11|歡喜和快樂的聲音、新郎和新娘的聲音，並聽見有人說： 你們要稱謝萬軍之耶和華， 因耶和華本為善， 他的慈愛永遠長存！ 他們奉感謝祭到耶和華的殿中；因為我必使這地被擄的人歸回，如起初一樣。這是耶和華說的。」
JER|33|12|萬軍之耶和華如此說：「在這荒廢、無人、無牲畜之地，並其中所有的城鎮，必再有牧人的草場，可讓羊群躺臥在那裏。
JER|33|13|在山區的城鎮、 謝非拉 的城鎮、 尼革夫 的城鎮、 便雅憫 地、 耶路撒冷 四圍的各處和 猶大 的城鎮，必再有羊群從數點的人手下經過。這是耶和華說的。
JER|33|14|「看哪，日子將到，我應許 以色列 家和 猶大 家的恩言必然實現。這是耶和華說的。
JER|33|15|在那些日子、那時候，我必使 大衛 公義的苗裔長起來；他必在地上施行公平和公義。
JER|33|16|在那些日子， 猶大 必得救， 耶路撒冷 必安然居住，他的名必稱為『耶和華－我們的義』。
JER|33|17|「因為耶和華如此說： 大衛 家必永遠不斷有人坐在 以色列 家的寶座上；
JER|33|18|利未 家的祭司也不斷有人在我面前獻燔祭、燒素祭，時常辦理獻祭的事。」
JER|33|19|耶和華的話臨到 耶利米 ，說：
JER|33|20|「耶和華如此說：你們若能廢棄我所立白日黑夜的約，使白日黑夜不按時輪轉，
JER|33|21|就能廢棄我與我僕人 大衛 所立的約，使他沒有後裔在他的寶座上作王，並能廢棄我與事奉我的 利未 家的祭司所立的約。
JER|33|22|正如天上的萬象不能數算，海邊的塵沙不能斗量，我必照樣使我僕人 大衛 的後裔和事奉我的 利未 人多起來。」
JER|33|23|耶和華的話臨到 耶利米 ，說：
JER|33|24|「你沒有留意這百姓所說的話嗎？他們說：『耶和華所揀選的二族，他已經棄絕了。』他們這樣藐視我的百姓，不把他們當作國來看待。
JER|33|25|耶和華如此說：除非我沒有立白日黑夜之約，也未曾安排天和地的定例，
JER|33|26|否則我不會棄絕 雅各 的後裔和我僕人 大衛 的後裔，使 大衛 的後裔不再治理 亞伯拉罕 、 以撒 、 雅各 的後裔。我必使他們被擄的人歸回，也必憐憫他們。」
JER|34|1|巴比倫 王 尼布甲尼撒 率領他的全軍和地上他管轄的各國各邦，攻打 耶路撒冷 和 耶路撒冷 所有的城鎮。那時，耶和華的話臨到 耶利米 ，說：
JER|34|2|「耶和華－ 以色列 的上帝說，你去告訴 猶大 王 西底家 ，耶和華如此說：看哪，我要把這城交在 巴比倫 王的手中，他必用火焚燒。
JER|34|3|你必不能逃脫他的手，定被拿住，交在他手中。你要親眼看到 巴比倫 王，他要親口跟你說話，你也必到 巴比倫 去。
JER|34|4|猶大 王 西底家 啊，你一定要聽耶和華的話。耶和華論到你如此說：你必不死於刀下；
JER|34|5|必平安而終，人要為你焚燒，好像為你祖先，就是在你以前早先的王焚燒一樣。人要為你舉哀說：『哀哉！我主啊。』這話是我說的。這是耶和華說的。」
JER|34|6|於是， 耶利米 先知在 耶路撒冷 把這一切話告訴 猶大 王 西底家 。
JER|34|7|那時， 巴比倫 王的軍隊正攻打 耶路撒冷 ，又攻打 猶大 僅存的城鎮，就是 拉吉 和 亞西加 ；原來 猶大 的堅固城只剩下這兩座。
JER|34|8|西底家 王與 耶路撒冷 的眾百姓立約，要他們宣告自由，叫各人釋放自己的僕人和婢女，使 希伯來 的男人和女人得自由，誰也不可使他的 猶大 弟兄作奴僕。這事以後，耶和華的話臨到 耶利米 。
JER|34|9|
JER|34|10|所有前來立約的領袖和眾百姓都順從，各人釋放自己的僕人和婢女，使他們得自由，不再叫他們作奴僕。大家都順從，將僕婢釋放了。
JER|34|11|但後來他們又反悔，叫被釋放得自由的僕人婢女回來，強迫他們仍為僕婢。
JER|34|12|因此耶和華的話臨到 耶利米 ，說：
JER|34|13|「耶和華－ 以色列 的上帝如此說：我將你們祖先從 埃及 地為奴之家領出時，與他們立約說：
JER|34|14|『你的一個 希伯來 弟兄若賣給你，服事你六年，到第七年你們各人就要釋放他自由出去。』只是你們祖先不聽我，不側耳而聽。
JER|34|15|如今你們回轉，行我眼中看為正的事，各人向鄰舍宣告自由，並且在我面前、在稱為我名下的殿中立約。
JER|34|16|你們卻反悔，褻瀆我的名，各人叫所釋放得自由的僕人婢女回來，強迫他們仍為僕婢。
JER|34|17|所以耶和華如此說：你們不聽從我，各人不向弟兄鄰舍宣告自由。看哪！我要向你們宣告自由，把你們自由地交給刀劍、饑荒、瘟疫，並且使地上萬國因你們而驚駭。這是耶和華說的。
JER|34|18|那些違背我約的人，就是不遵守在我面前立約之話的，我要使他們成了那劈成兩半的牛犢，使人從切塊中經過：
JER|34|19|猶大 的領袖、 耶路撒冷 的領袖、官員、祭司，和從牛犢切塊中經過的這地的眾百姓，
JER|34|20|我必將他們交在仇敵和尋索其命的人手中；他們的屍首必給空中的飛鳥和地上的走獸作食物。
JER|34|21|我必將 猶大 王 西底家 和他的眾領袖交在仇敵和尋索其命的人手中，與那暫時離你們而去的 巴比倫 王軍隊的手中。
JER|34|22|看哪，我要吩咐他們回到這城，攻打這城，將城攻取，用火焚燒；我也要使 猶大 的城鎮變為廢墟，無人居住。這是耶和華說的。」
JER|35|1|當 約西亞 的兒子 約雅敬 作 猶大 王的時候，耶和華的話臨到 耶利米 ，說：
JER|35|2|「你去見 利甲 族的人，吩咐他們，領他們進入耶和華殿的一個房間，給他們酒喝。」
JER|35|3|我就帶 哈巴洗尼雅 的孫子 雅利米雅 的兒子 雅撒尼亞 ，和他的兄弟，並他所有的兒子，以及 利甲 全族的人，
JER|35|4|領他們到耶和華的殿，進入 伊基大利 的兒子神人 哈難 兒子們的房間；那房間靠近官長的房間，在 沙龍 之子門口的守衛 瑪西雅 的房間上面。
JER|35|5|於是我在 利甲 族的人面前擺設盛滿了酒的碗和杯，對他們說：「請喝酒。」
JER|35|6|他們卻說：「我們不喝酒，因為我們祖先 利甲 的兒子 約拿達 曾吩咐我們說：『你們與你們的子孫永不可喝酒，
JER|35|7|不可蓋房子，不可撒種，也不可栽葡萄園，連擁有都不可；但一生的年日要住帳棚，使你們的日子在寄居的地面上得以長久。』
JER|35|8|凡我們祖先 利甲 的兒子 約拿達 所吩咐我們的話，我們都聽從了。我們和我們的妻子兒女一生的年日都不喝酒，
JER|35|9|不蓋房子居住，我們也沒有葡萄園、田地和種子；
JER|35|10|但住在帳棚裏，聽從並遵行我們祖先 約拿達 所吩咐我們的一切話。
JER|35|11|巴比倫 王 尼布甲尼撒 上來攻打這地的時候，我們說：『來吧，我們到 耶路撒冷 去，躲避 迦勒底 的軍隊和 亞蘭 的軍隊。』這樣，我們才住在 耶路撒冷 。」
JER|35|12|耶和華的話臨到 耶利米 ，說：
JER|35|13|「萬軍之耶和華－ 以色列 的上帝如此說：你去對 猶大 人和 耶路撒冷 的居民說，你們不肯領受訓誨，聽從我的話嗎？這是耶和華說的。
JER|35|14|利甲 的兒子 約拿達 所吩咐他子孫不可喝酒的話，他們已經遵守了；他們因為聽從祖先的吩咐，直到今日都不喝酒。至於我，我一再警戒你們，你們卻不肯聽從我。
JER|35|15|我一再差遣我的僕人眾先知到你們那裏去，說：『你們各人當回頭離開惡道，改正行為，不再隨從事奉別神，如此，就必住在我所賜給你們和你們祖先的地上。』只是你們不側耳而聽，也不聽我。
JER|35|16|利甲 的兒子 約拿達 的子孫能遵守祖先所吩咐他們的命令，這百姓卻不肯聽從我！
JER|35|17|因此，耶和華－萬軍之上帝、 以色列 的上帝如此說：看哪，我要使我所說的一切災禍臨到 猶大 人和 耶路撒冷 所有的居民。因為我向他們說話，他們不聽從；我呼喚他們，他們也沒有回應。」
JER|35|18|耶利米 對 利甲 族的人說：「萬軍之耶和華－ 以色列 的上帝如此說：因你們聽從你們祖先 約拿達 的吩咐，謹守他的一切命令，照他所吩咐的去做，
JER|35|19|所以萬軍之耶和華－ 以色列 的上帝如此說： 利甲 的兒子 約拿達 必永遠不斷有人侍立在我面前。」
JER|36|1|約西亞 的兒子 猶大 王 約雅敬 第四年，有這話從耶和華臨到 耶利米 ，說：
JER|36|2|「你要取一書卷，把我對你所說攻擊 以色列 和 猶大 ，並各國的一切話，從我對你說話的那日，就是從 約西亞 的日子起直到今日，都寫在其上；
JER|36|3|或者 猶大 家聽見我想要降給他們的一切災禍，各人就回轉離開惡道，我就赦免他們的罪孽和罪惡。」
JER|36|4|耶利米 召了 尼利亞 的兒子 巴錄 來； 巴錄 就從 耶利米 口中，把耶和華對 耶利米 所說的一切話寫在書卷上。
JER|36|5|耶利米 吩咐 巴錄 說：「我被禁止，不能進耶和華的殿。
JER|36|6|所以你要趁禁食的日子進入耶和華的殿中，把耶和華的話，就是你從我口中寫在書卷上的話，念給百姓和所有從各城鎮前來的 猶大 人親耳聽；
JER|36|7|或者他們的懇求達到耶和華面前，各人回轉離開惡道，因為耶和華向這百姓所說要發的怒氣和憤怒實在很大。」
JER|36|8|尼利亞 的兒子 巴錄 就照 耶利米 先知所吩咐的一切去做，在耶和華殿中宣讀書卷上耶和華的話。
JER|36|9|約西亞 的兒子 猶大 王 約雅敬 第五年九月， 耶路撒冷 的眾百姓和那從 猶大 城鎮前來 耶路撒冷 的眾百姓，在耶和華面前宣告禁食，
JER|36|10|巴錄 就在耶和華殿的上院，靠近耶和華殿的 新門 口， 沙番 的兒子 基瑪利雅 文士的房間裏，宣讀書卷上 耶利米 的話給眾百姓親耳聽。
JER|36|11|沙番 的孫子 基瑪利雅 的兒子 米該亞 聽見書卷上耶和華的一切話，
JER|36|12|就下到王宮，進入書記的房間。看哪，所有的官長都坐在那裏，包括 以利沙瑪 文士、 示瑪雅 的兒子 第萊雅 、 亞革波 的兒子 以利拿單 、 沙番 的兒子 基瑪利雅 、 哈拿尼雅 的兒子 西底家 和其餘的官長。
JER|36|13|米該亞 向他們述說他所聽見的一切話，就是當 巴錄 向眾百姓宣讀那書卷時親耳聽見的。
JER|36|14|官長們就派 猶底 ，就是 古示 的曾孫， 示利米雅 的孫子， 尼探雅 的兒子到 巴錄 那裏，對他說：「你把你所念給百姓聽的書卷拿在手裏，到我們這裏來。」 尼利亞 的兒子 巴錄 就手拿書卷到他們那裏來。
JER|36|15|他們對他說：「請坐下，念給我們親耳聽。」 巴錄 就念給他們親耳聽。
JER|36|16|他們聽見這一切話就害怕，面面相覷，對 巴錄 說：「我們必須將這一切話稟告王。」
JER|36|17|他們問 巴錄 說：「請你告訴我們，你怎樣從他口中寫下這一切話呢？」
JER|36|18|巴錄 回答說：「他向我口述這一切話，我就用筆墨把它寫在書卷上。」
JER|36|19|眾官長對 巴錄 說：「你和 耶利米 要去躲起來，不可叫人知道你們躲在哪裏。」
JER|36|20|眾官長把書卷留在 以利沙瑪 文士的房間裏，然後進院見王，把這一切話說給王聽。
JER|36|21|王就派 猶底 去拿這書卷來；他就從 以利沙瑪 文士的房間內取來，念給王和侍立在王左右的眾官長親耳聽。
JER|36|22|那時正是九月，王坐在過冬的房屋裏，王前面有燃燒的火盆 。
JER|36|23|猶底 念了三、四段 ，王就用文士的刀把書卷割破，丟在火盆裏，直到全卷在火中燒盡了。
JER|36|24|王和聽見這一切話的臣僕都不懼怕，也不撕裂衣服。
JER|36|25|以利拿單 和 第萊雅 ，並 基瑪利雅 懇求王不要燒這書卷，王卻不聽。
JER|36|26|王吩咐王 的兒子 耶拉篾 、 亞斯列 的兒子 西萊雅 和 亞伯疊 的兒子 示利米雅 ，去捉拿 巴錄 文士和 耶利米 先知；耶和華卻將他們隱藏起來。
JER|36|27|王燒了有 巴錄 從 耶利米 口中所寫之話的書卷以後，耶和華的話臨到 耶利米 ，說：
JER|36|28|「你再取一書卷，將 猶大 王 約雅敬 所燒前一卷書上原有的一切話寫在上面。
JER|36|29|論到 猶大 王 約雅敬 你要說，耶和華如此說：你燒了這書卷，說：『你為甚麼在上面寫著， 巴比倫 王必要來毀滅這地，使這地絕了人民和牲畜呢？』
JER|36|30|所以耶和華論到 猶大 王 約雅敬 說：他後裔中必沒有人坐在 大衛 的寶座上；他的屍首必被拋棄，白天受炎熱，黑夜受寒霜。
JER|36|31|我必因他和他後裔，並他臣僕的罪孽懲罰他們。我要使我所說的一切災禍臨到他們和 耶路撒冷 的居民，並 猶大 人；只是他們不肯聽從。」
JER|36|32|於是， 耶利米 又取一書卷交給 尼利亞 的兒子 巴錄 文士，他就從 耶利米 的口中寫了 猶大 王 約雅敬 在火中所燒書卷上的一切話，另外又添了許多相仿的話。
JER|37|1|約西亞 的兒子 西底家 接續 約雅敬 的兒子 哥尼雅 作王，因為 巴比倫 王 尼布甲尼撒 立他在 猶大 地作王。
JER|37|2|但 西底家 、他的臣僕和這地的百姓都不聽從耶和華藉 耶利米 先知所說的話。
JER|37|3|西底家 王派 示利米雅 的兒子 猶甲 和 瑪西雅 的兒子 西番雅 祭司，去見 耶利米 先知，說：「求你為我們祈求耶和華－我們的上帝。」
JER|37|4|那時 耶利米 仍在百姓中進出，因為他們還沒有把他囚在監裏。
JER|37|5|法老的軍隊已經從 埃及 出來，那圍困 耶路撒冷 的 迦勒底 人聽見這風聲，就拔營離開 耶路撒冷 去了。
JER|37|6|耶和華的話臨到 耶利米 先知，說：
JER|37|7|「耶和華－ 以色列 的上帝如此說：你們要對派你們來求問我的 猶大 王如此說：『看哪，那出來幫助你們的法老軍隊必回 埃及 本國去。
JER|37|8|迦勒底 人必再來攻打這城，並要攻下，用火焚燒。
JER|37|9|耶和華如此說：你們不要自欺說「 迦勒底 人必定離開我們」，因為他們必不離開。
JER|37|10|你們即使擊敗與你們爭戰的 迦勒底 全軍，他們當中剩下受傷的人也必各自從帳棚裏起來，用火焚燒這城。』」
JER|37|11|迦勒底 的軍隊因躲避法老的軍隊，拔營離開 耶路撒冷 的時候，
JER|37|12|耶利米 離開 耶路撒冷 ，往 便雅憫 地去，要在那裏從百姓當中取得自己的地產。
JER|37|13|他到了 便雅憫門 ，那裏的守門官名叫 伊利雅 ，是 哈拿尼亞 的孫子， 示利米雅 的兒子，他逮捕 耶利米 先知，說：「你是去投降 迦勒底 人的！」
JER|37|14|耶利米 說：「你這是謊話，我並不是去投降 迦勒底 人。」 伊利雅 不聽 耶利米 的話，就逮捕他，把他帶到官長那裏。
JER|37|15|官長們惱怒 耶利米 ，打了他，把他囚在 約拿單 文士的房屋中，因為他們把這屋子當作監牢。
JER|37|16|耶利米 來到地牢，進入牢房，在那裏拘留多日。
JER|37|17|西底家 王差人提他出來，在自己的宮內私下問他說：「有甚麼話從耶和華臨到沒有？」 耶利米 說：「有！」又說：「你必被交在 巴比倫 王手中。」
JER|37|18|耶利米 又對 西底家 王說：「我在甚麼事上得罪你，或你的臣僕，或這百姓，你們竟將我囚在監裏呢？
JER|37|19|對你們預言『 巴比倫 王必不來攻擊你們和這地』的先知在哪裏呢？
JER|37|20|主－我的王啊，現在求你垂聽，允准我在你面前的懇求：不要把我送回 約拿單 文士的房屋中，免得我死在那裏。」
JER|37|21|於是 西底家 王下令，他們就把 耶利米 交在護衛兵的院中，每天從餅店街取一個餅給他，直到城中所有的餅都用盡了。這樣， 耶利米 仍拘留在護衛兵的院中。
JER|38|1|瑪坦 的兒子 示法提雅 、 巴施戶珥 的兒子 基大利 、 示利米雅 的兒子 猶甲 、 瑪基雅 的兒子 巴示戶珥 聽見 耶利米 對眾百姓所說的話，說：
JER|38|2|「耶和華如此說：留在這城裏的必遭刀劍、饑荒、瘟疫而死，但歸向 迦勒底 人的必得存活；至少能保全自己的性命，得以存活。
JER|38|3|耶和華如此說：這城必要交在 巴比倫 王軍隊的手中，他必攻下這城。」
JER|38|4|於是官長們對王說：「求你把這人處死，因他向城裏剩下的士兵和眾人說這樣的話，使他們的手發軟。這人不是為這百姓求平安，而是叫他們受災禍。」
JER|38|5|西底家 王說：「看哪，他在你們手中，王不能反對你們所做的事。」
JER|38|6|他們就拿住 耶利米 ，把他丟在王 的兒子 瑪基雅 的井裏；那口井在護衛兵的院中。他們用繩子把 耶利米 縋下去，井裏沒有水，只有淤泥， 耶利米 就陷在淤泥中。
JER|38|7|在王宮裏的太監 古實 人 以伯‧米勒 ，聽見他們把 耶利米 丟進井裏，那時王坐在 便雅憫門 前。
JER|38|8|以伯‧米勒 從王宮裏出來，對王說：
JER|38|9|「主－我的王啊，這些人向 耶利米 先知一味地行惡，把他丟在井裏；他在那裏必因飢餓而死，因為城裏不再有糧食了。」
JER|38|10|王就吩咐 古實 人 以伯‧米勒 說：「你從這裏帶領三十人，趁 耶利米 先知還沒死，把他從井裏拉上來。」
JER|38|11|於是 以伯‧米勒 帶領這些人同去，進入王宮，到庫房以下 ，從那裏取了些碎布和破衣服，用繩子縋下去，到井裏 耶利米 那裏。
JER|38|12|古實 人 以伯‧米勒 對 耶利米 說：「你用這些碎布和破衣服放在繩子上，墊你的腋下。」 耶利米 就照樣做。
JER|38|13|這樣，他們用繩子將 耶利米 從井裏拉上來。 耶利米 仍在護衛兵的院中。
JER|38|14|西底家 王差人將 耶利米 先知帶進耶和華殿的第三個門，到王那裏去。王對 耶利米 說：「我要問你一件事，你一點都不可向我隱瞞。」
JER|38|15|耶利米 對 西底家 說：「我若告訴你，你豈不是一定要把我處死嗎？我若勸你，你必不聽我。」
JER|38|16|西底家 王就私下對 耶利米 說：「我指著那造我們生命之永生的耶和華起誓：我必不把你處死，也不將你交在尋索你命的人手中。」
JER|38|17|耶利米 對 西底家 說：「耶和華－萬軍之上帝、 以色列 的上帝如此說：你若歸順 巴比倫 王的官長，你的命就必存活，這城也不致被火焚燒，你和你的全家都必存活。
JER|38|18|你若不歸順 巴比倫 王的官長，這城必交在 迦勒底 人手中。他們必用火焚燒，你也不得脫離他們的手。」
JER|38|19|西底家 王對 耶利米 說：「我怕那些投降 迦勒底 人的 猶大 人，恐怕 迦勒底 人把我交在他們手中，他們就戲弄我。」
JER|38|20|耶利米 說：「 迦勒底 人必不把你交出。求你聽從我對你所說耶和華的話，這樣對你有好處，你的命也必存活。
JER|38|21|你若不肯歸順，耶和華指示我的話是這樣：
JER|38|22|看哪， 猶大 王宮裏所留下來的婦女必被帶到 巴比倫 王的官長那裏。這些婦女要說： 你知己的朋友引誘你， 他們勝過你； 你的腳陷入淤泥， 他們卻離棄你。
JER|38|23|「人必將你的后妃和你的兒女帶到 迦勒底 人那裏；你也不得脫離他們的手，必被 巴比倫 王的手捉住，這城也必被火焚燒 。」
JER|38|24|西底家 對 耶利米 說：「不要讓人知道這些對話，你就不至於死。
JER|38|25|官長們若聽見我跟你說話，到你那裏對你說：『告訴我們，你對王說了甚麼話，王又向你說了甚麼；不可向我們隱瞞，否則我們就要殺你。』
JER|38|26|你就對他們說：『我在王面前懇求不要把我送回 約拿單 的房屋，免得我死在那裏。』」
JER|38|27|隨後官長們到 耶利米 那裏，問他，他就照王所吩咐的一切話回答他們。他們就不再問他，因為事情沒有洩漏。
JER|38|28|於是 耶利米 仍在護衛兵的院中，直到 耶路撒冷 被攻下的日子。當 耶路撒冷 被攻下時，他仍在那裏。
JER|39|1|猶大 王 西底家 第九年十月， 巴比倫 王 尼布甲尼撒 率領全軍前來圍困 耶路撒冷 。
JER|39|2|西底家 十一年四月初九日，城被攻破。
JER|39|3|耶路撒冷 被攻下的時候， 巴比倫 王的眾官長， 尼甲‧沙利薛 、 三甲‧尼波 、 撒西金 將軍 、 尼甲‧沙利薛 將軍 ，並 巴比倫 王其餘的官長都來坐在 中門 。
JER|39|4|猶大 王 西底家 和所有士兵看見他們，就在夜間從靠近王的花園、兩城牆中間的門逃跑出城，往 亞拉巴 逃去。
JER|39|5|迦勒底 的軍隊追趕他們，在 耶利哥 的平原追上 西底家 ，將他逮住，帶到 哈馬 地的 利比拉 、 巴比倫 王 尼布甲尼撒 那裏； 尼布甲尼撒 就判他的罪。
JER|39|6|在 利比拉 ， 巴比倫 王在 西底家 眼前殺了他的兒女； 巴比倫 王又殺了 猶大 所有的貴族，
JER|39|7|並且挖了 西底家 的眼睛，用銅鏈鎖住他，要帶到 巴比倫 去。
JER|39|8|迦勒底 人用火焚燒王宮和百姓的房屋，又拆毀 耶路撒冷 的城牆。
JER|39|9|那時， 尼布撒拉旦 護衛長把城裏所剩下的百姓和投降他的降民，以及其餘的百姓都擄到 巴比倫 去了。
JER|39|10|尼布撒拉旦 護衛長卻把百姓中一無所有的窮人留在 猶大 地，當時就賞給他們葡萄園和田地 。
JER|39|11|巴比倫 王 尼布甲尼撒 為了 耶利米 ，囑咐 尼布撒拉旦 護衛長：
JER|39|12|「你領他去，好好地看待他，切不可害他；他對你怎麼說，你就向他怎樣做。」
JER|39|13|尼布撒拉旦 護衛長和 尼布沙斯班 將軍 、 尼甲‧沙利薛 將軍 ，並 巴比倫 王眾官長，
JER|39|14|派人把 耶利米 從護衛兵的院中提出來，交給 沙番 的孫子， 亞希甘 的兒子 基大利 ，讓他自由進出屋子；於是 耶利米 住在百姓中間。
JER|39|15|耶利米 還囚在護衛兵院中的時候，耶和華的話臨到他，說：
JER|39|16|「你去告訴 古實 人 以伯‧米勒 說，萬軍之耶和華－ 以色列 的上帝如此說：看哪，我說降禍不降福的話必臨到這城，到那時必在你面前實現。
JER|39|17|到那日我必拯救你，你必不致交在你所怕的人手中。這是耶和華說的。
JER|39|18|我定要搭救你，你必不致倒在刀下，卻要保全自己的性命，因你倚靠我。這是耶和華說的。」
JER|40|1|耶利米 被鏈子鎖在 耶路撒冷 和 猶大 被擄到 巴比倫 的人中， 尼布撒拉旦 護衛長把他從 拉瑪 提出來，釋放他以後，耶和華的話臨到 耶利米 。
JER|40|2|護衛長提 耶利米 來，對他說：「耶和華－你的上帝曾說要降這災禍給此地。
JER|40|3|耶和華照他所說的做了，已使這災禍臨到；因你們得罪耶和華，不聽從他的話，所以這事臨到你們。
JER|40|4|看哪，現在我解開你手上的鏈子，你若看與我同往 巴比倫 去好，就可以去，我必厚待你；你若看與我同往 巴比倫 去不好，就不必去。看哪，全地在你面前，你以為哪裏美好，哪裏合宜，只管去吧
JER|40|5|─ 耶利米 尚未回去 ─你可以回到 巴比倫 王所立管理 猶大 城鎮的 沙番 的孫子， 亞希甘 的兒子 基大利 那裏去，在他那裏住在百姓當中。不然，你看哪裏合宜就可以去。」於是護衛長送他糧食和禮物，釋放了他。
JER|40|6|耶利米 就來到 米斯巴 ， 亞希甘 的兒子 基大利 那裏去，與他同住，住在留於境內的百姓當中。
JER|40|7|在鄉間所有的軍官和屬他們的人，聽見 巴比倫 王立了 亞希甘 的兒子 基大利 作當地的省長，並將沒有擄到 巴比倫 的男人、婦女、孩童和當地極窮的人全交給他，
JER|40|8|於是 尼探雅 的兒子 以實瑪利 ， 加利亞 的兩個兒子 約哈難 和 約拿單 ， 單戶篾 的兒子 西萊雅 ，並 尼陀法 人 以斐 的眾子， 瑪迦 人的兒子 耶撒尼亞 ，和屬他們的人，都來到 米斯巴 的 基大利 那裏。
JER|40|9|沙番 的孫子， 亞希甘 的兒子 基大利 向他們和屬他們的人起誓說：「不要怕服事 迦勒底 人，只管住在這地，服事 巴比倫 王，就可以得福。
JER|40|10|至於我，我要住在 米斯巴 ，侍候那些到我們這裏來的 迦勒底 人；只是你們當積蓄酒、油和夏天的果子，收藏在器皿裏，並住在你們所佔的城鎮中。」
JER|40|11|在 摩押 地和 亞捫 人當中，在 以東 地和各國，所有的 猶大 人聽見 巴比倫 王留下一些 猶大 人，並立 沙番 的孫子、 亞希甘 的兒子 基大利 管理他們，
JER|40|12|所有的 猶大 人就從被趕到的各處回來，到 猶大 地 米斯巴 的 基大利 那裏。他們積蓄了許多的酒，並夏天的果子。
JER|40|13|加利亞 的兒子 約哈難 和在鄉間的軍官來到 米斯巴 的 基大利 那裏，
JER|40|14|對他說：「 亞捫 人的王 巴利斯 派 尼探雅 的兒子 以實瑪利 來謀害你的命，你知道嗎？」 亞希甘 的兒子 基大利 卻不相信他們的話。
JER|40|15|加利亞 的兒子 約哈難 在 米斯巴 私下對 基大利 說：「求你容我去殺 尼探雅 的兒子 以實瑪利 ，必無人知道。何必讓他害你的命，使聚集到你這裏來的 猶大 人都分散，以致 猶大 剩餘的人都滅亡呢？」
JER|40|16|亞希甘 的兒子 基大利 對 加利亞 的兒子 約哈難 說：「你不可做這事，你所論 以實瑪利 的話是假的。」
JER|41|1|七月中，王的大臣，就是王室後裔 以利沙瑪 的孫子、 尼探雅 的兒子 以實瑪利 帶著十個人，來到 米斯巴 ， 亞希甘 的兒子 基大利 那裏；他們在 米斯巴 一同吃飯。
JER|41|2|尼探雅 的兒子 以實瑪利 和同他來的那十個人起來，用刀擊殺 沙番 的孫子， 亞希甘 的兒子 基大利 ，就是 巴比倫 王所立為當地省長的，把他殺死。
JER|41|3|以實瑪利 把所有在 米斯巴 與 基大利 一起的 猶大 人，以及他們在那裏所遇見的 迦勒底 人和士兵都殺了。
JER|41|4|他殺了 基大利 的第二天，還沒有人知道的時候，
JER|41|5|有八十人從 示劍 、 示羅 和 撒瑪利亞 前來，鬍鬚剃去，衣服撕裂，身體劃破，手拿素祭和乳香，要奉到耶和華的殿。
JER|41|6|尼探雅 的兒子 以實瑪利 從 米斯巴 出來迎接他們，隨走隨哭，遇見了他們，就對他們說：「你們可以到 亞希甘 的兒子 基大利 那裏。」
JER|41|7|他們到了城中， 尼探雅 的兒子 以實瑪利 和與他一起的人就把他們殺了，丟在坑裏。
JER|41|8|只是他們中間有十個人對 以實瑪利 說：「不要殺我們，因為我們有許多大麥、小麥、油和蜜藏在田間。」於是他住手，沒有在弟兄中間殺他們。
JER|41|9|以實瑪利 把那些因 基大利 事件所殺之人的屍首都丟在坑裏；這坑是從前 亞撒 王因怕 以色列 王 巴沙 所挖的。 尼探雅 的兒子 以實瑪利 把那些被殺的人填滿了坑。
JER|41|10|以實瑪利 把 米斯巴 剩下的人，就是眾公主和仍住在 米斯巴 所有的百姓都擄去，他們原是 尼布撒拉旦 護衛長交給 亞希甘 的兒子 基大利 的。 尼探雅 的兒子 以實瑪利 擄了他們，要到 亞捫 人那裏去。
JER|41|11|加利亞 的兒子 約哈難 和與他一起的軍官，聽見 尼探雅 的兒子 以實瑪利 所做的一切惡事，
JER|41|12|就帶領眾人前往，要和 尼探雅 的兒子 以實瑪利 爭戰，他們在 基遍 的大水池 旁遇見他。
JER|41|13|在 以實瑪利 那裏的眾人看見 加利亞 的兒子 約哈難 和與他一起的軍官，就都歡喜。
JER|41|14|這樣， 以實瑪利 從 米斯巴 所擄去的眾人都轉而歸向 加利亞 的兒子 約哈難 。
JER|41|15|尼探雅 的兒子 以實瑪利 和八個人脫離 約哈難 的手，逃到 亞捫 人那裏去。
JER|41|16|尼探雅 的兒子 以實瑪利 殺了 亞希甘 的兒子 基大利 ，從 米斯巴 把所有倖存的百姓、士兵、婦女、孩童、太監擄到 基遍 之後， 加利亞 的兒子 約哈難 和與他一起的軍官把他們都搶回來，
JER|41|17|帶到靠近 伯利恆 的 基羅特金罕 住下，要到 埃及 去，
JER|41|18|躲避 迦勒底 人。他們懼怕 迦勒底 人，因為 尼探雅 的兒子 以實瑪利 殺了 巴比倫 王所立管理那地的 亞希甘 的兒子 基大利 。
JER|42|1|眾軍官和 加利亞 的兒子 約哈難 ，並 何沙雅 的兒子 耶撒尼亞 以及眾百姓，從最小的到最大的都進前來，
JER|42|2|對 耶利米 先知說：「請你准我們在你面前祈求，為我們這倖存的人向耶和華－你的上帝禱告。我們本來眾多，現在剩下的極少，這是你親眼看見的。
JER|42|3|願耶和華－你的上帝指示我們當走的路，當做的事。」
JER|42|4|耶利米 先知對他們說：「我已經聽見了，看哪，我必照你們的話向耶和華－你們的上帝禱告。耶和華無論回答甚麼，我都必告訴你們，絕不隱瞞。」
JER|42|5|於是他們對 耶利米 說：「我們若不照耶和華－你上帝差遣你說的一切話去做，願耶和華在我們中間作真實可靠的見證。
JER|42|6|我們請你到耶和華－我們的上帝面前，他說的無論是好是歹，我們都必聽從；因為我們聽從耶和華－我們上帝的話，就可以得福。」
JER|42|7|過了十天，耶和華的話臨到 耶利米 。
JER|42|8|他就將 加利亞 的兒子 約哈難 和與他一起所有的軍官和百姓，從最小的到最大的都召來，
JER|42|9|對他們說：「你們請我到耶和華－ 以色列 的上帝面前為你們祈求，他如此說：
JER|42|10|『你們若仍留在這地，我就建立你們，必不拆毀；栽植你們，必不拔出；因我為所降與你們的災禍感到遺憾。
JER|42|11|不要怕你們所懼怕的 巴比倫 王。不要怕他！因為我與你們同在，要拯救你們脫離他的手。這是耶和華說的。
JER|42|12|我要向你們施憐憫，他 就憐憫你們，使你們歸回本地。』
JER|42|13|倘若你們說：『我們不留在這地』，不聽從耶和華－你們上帝的話，
JER|42|14|說：『我們不留在這地，卻要進入 埃及 地，在那裏我們看不見戰爭，聽不見角聲，也不致缺食挨餓；我們要住在那裏。』
JER|42|15|倖存的 猶大 人哪，你們現在要聽耶和華的話；萬軍之耶和華－ 以色列 的上帝如此說：『你們若定意進入 埃及 ，在那裏寄居，
JER|42|16|你們所懼怕的刀劍在 埃及 地必追上你們，你們所懼怕的饑荒在 埃及 要緊緊跟隨你們，你們必死在那裏。
JER|42|17|凡定意進入 埃及 在那裏寄居的，必遭刀劍、饑荒、瘟疫而死，無一人存留，得以逃脫我所降與他們的災禍。』
JER|42|18|「萬軍之耶和華－ 以色列 的上帝如此說：『我怎樣將我的怒氣和憤怒傾倒在 耶路撒冷 的居民身上，你們進入 埃及 的時候，我也必照樣將我的憤怒傾倒在你們身上，以致你們受辱罵、驚駭、詛咒、羞辱，並且不得再看見這地方。』
JER|42|19|倖存的 猶大 人哪，耶和華論到你們說：『不要進入 埃及 。』你們要確實知道，我今日已警戒你們了。
JER|42|20|你們行詭詐害自己；因為你們請我到耶和華－你們上帝那裏，說：『請你為我們向耶和華－我們的上帝禱告，你把耶和華－我們上帝所說的一切告訴我們，我們就必遵行。』
JER|42|21|我今日把這話告訴你們，你們卻不聽耶和華－你們上帝為這一切事差我到你們那裏所說的話。
JER|42|22|現在你們要確實知道，你們在所要去的寄居之地必遭刀劍、饑荒、瘟疫而死。」
JER|43|1|耶利米 向眾百姓說完了耶和華－他們上帝一切的話，就是耶和華－他們上帝差他去說的這一切話，
JER|43|2|何沙雅 的兒子 亞撒利雅 和 加利亞 的兒子 約哈難 ，以及所有狂傲的人，就對 耶利米 說：「你說謊！耶和華－我們的上帝並沒有差遣你說：『你們不可進入 埃及 ，在那裏寄居。』
JER|43|3|這是 尼利亞 的兒子 巴錄 挑唆你害我們，要把我們交在 迦勒底 人手中，使我們被殺或被擄到 巴比倫 去。」
JER|43|4|加利亞 的兒子 約哈難 和所有的軍官、百姓，都不肯聽從耶和華的話留在 猶大 地。
JER|43|5|加利亞 的兒子 約哈難 和所有的軍官卻將倖存的 猶大 人，就是從被趕到的各國回來，在 猶大 地寄居的男人、婦女、孩童和眾公主，並 尼布撒拉旦 護衛長留在 沙番 的孫子， 亞希甘 的兒子 基大利 那裏的眾人，與 耶利米 先知，以及 尼利亞 的兒子 巴錄 ，
JER|43|6|
JER|43|7|都帶入 埃及 地，到了 答比匿 ；這是因他們不肯聽從耶和華的話。
JER|43|8|在 答比匿 ，耶和華的話臨到 耶利米 ，說：
JER|43|9|「你要在 猶大 人眼前用手拿幾塊大石頭，藏在 答比匿 法老的宮門砌磚的石墩上，
JER|43|10|對他們說：『萬軍之耶和華－ 以色列 的上帝如此說：看哪，我必召我的僕人 巴比倫 王 尼布甲尼撒 前來，安置他的寶座在所藏的這些石頭上；他要在其上支搭華麗的帳幕。
JER|43|11|他要來攻擊 埃及 地： 定為死亡的，必致死亡； 定為擄掠的，必遭擄掠； 定為刀殺的，必被刀殺。
JER|43|12|我要用火點燃 埃及 眾神明的廟宇， 巴比倫 王要焚燒廟宇，擄去神像；他要圍住 埃及 地，好像牧人披上外衣，從那裏安然而去。
JER|43|13|他必打碎 埃及 地 伯‧示麥 的柱像，用火焚燒 埃及 眾神明的廟宇。』」
JER|44|1|有話臨到 耶利米 ，論到住 埃及 地所有的 猶大 人，就是住在 密奪 、 答比匿 、 挪弗 、 巴特羅 境內的 猶大 人，說：
JER|44|2|「萬軍之耶和華－ 以色列 的上帝如此說：我所降與 耶路撒冷 和 猶大 各城的一切災禍，你們都看見了。看哪，那些城鎮今日荒涼，無人居住；
JER|44|3|這是因居民所行的惡，去燒香事奉別神，就是他們和你們，以及你們列祖所不認識的神明，惹我發怒。
JER|44|4|我一再差遣我的僕人眾先知去，說：你們切不可行我所厭惡這可憎之事。
JER|44|5|他們卻不聽從，不側耳而聽，也不轉離惡事，仍向別神燒香。
JER|44|6|因此，我的怒氣和憤怒都傾倒出來，在 猶大 城鎮和 耶路撒冷 街市上燃起，以致它們都荒廢淒涼，正如今日一樣。
JER|44|7|現在耶和華－萬軍之上帝、 以色列 的上帝如此說：你們為何做這大惡自害己命，使你們的男人、婦女、孩童和吃奶的都從 猶大 剪除，不留一人呢？
JER|44|8|你們以手所做的，在寄居的 埃及 地向別神燒香，惹我發怒，使你們被剪除，在天下萬國中受詛咒羞辱。
JER|44|9|你們祖先的惡行， 猶大 諸王和后妃的惡行，你們自己和你們妻子的惡行，就是在 猶大 地和 耶路撒冷 街市上所做的，你們都忘了嗎？
JER|44|10|到如今你們還不懊悔，不懼怕，不肯遵行我在你們和你們祖先面前所設立的法度律例。
JER|44|11|「所以萬軍之耶和華－ 以色列 的上帝如此說：看哪，我必向你們變臉降災，剪除 猶大 眾人。
JER|44|12|我必使那定意進入 埃及 地、在那裏寄居的，就是倖存的 猶大 人，盡都滅絕。他們必在 埃及 地仆倒，因刀劍饑荒滅絕，從最小的到最大的都必遭刀劍饑荒而死，甚至受辱罵、驚駭、詛咒、羞辱。
JER|44|13|我怎樣用刀劍、饑荒、瘟疫懲罰 耶路撒冷 ，也必照樣懲罰那些住在 埃及 地的 猶大 人。
JER|44|14|那進入 埃及 地、在那裏寄居的，就是倖存的 猶大 人，都不得逃脫，也不得歸回 猶大 地。他們心中很想歸回，居住在那裏；但除了少數逃脫的以外，都不得歸回。」
JER|44|15|那些知道自己妻子向別神燒香的男人，與站在那裏的一大群婦女，就是住 埃及 地 巴特羅 所有的百姓，回答 耶利米 說：
JER|44|16|「論到你奉耶和華的名向我們所說的話，我們必不聽從。
JER|44|17|我們定要照我們口中所說的一切話去做，向天后燒香，獻澆酒祭，按著我們與我們祖先、君王、官長在 猶大 城鎮和 耶路撒冷 街市上素常所做的一樣；因為那時我們得以吃飽、享福樂，並未遇見災禍。
JER|44|18|自從我們停止向天后燒香，獻澆酒祭，我們倒缺乏這一切，又因刀劍饑荒滅絕。」
JER|44|19|婦女們說 ：「我們向天后燒香，獻澆酒祭，做天后像的餅供奉它，向它獻澆酒祭，難道我們的丈夫沒有參與嗎？」
JER|44|20|耶利米 對這樣回答他的男人和婦女說：
JER|44|21|「你們與你們祖先、君王、官長，以及這地的百姓，在 猶大 城鎮和 耶路撒冷 街市上所燒的香，耶和華豈不記得，放在他心上嗎？
JER|44|22|耶和華因你們所行的惡、所做可憎的事，不能再容忍，所以使你們的地荒涼，受驚駭詛咒，無人居住，正如今日一樣。
JER|44|23|你們燒香，得罪耶和華，不聽耶和華的話，不遵行他的律法、條例、法度，所以你們遭遇這災禍，正如今日一樣。」
JER|44|24|耶利米 又對眾百姓和婦女說：「所有在 埃及 地的 猶大 人哪，當聽耶和華的話。
JER|44|25|萬軍之耶和華－ 以色列 的上帝如此說：你們和你們的妻子口中說過、手裏做到，說：『我們定要向天后還願，向它燒香，獻澆酒祭。』現在你們儘管堅定所許的願，去還願吧！
JER|44|26|所有住 埃及 地的 猶大 人哪，當聽耶和華的話。耶和華說：看哪，我指著我至大的名起誓，在 埃及 全地，我的名必不再被 猶大 任何人的口呼喊：『我指著主－永生的耶和華起誓。』
JER|44|27|看哪，我看守他們，為要降禍不降福；在 埃及 地的 猶大 人必因刀劍、饑荒而滅亡，直到滅絕。
JER|44|28|從 埃及 地能脫離刀劍、歸回 猶大 地的人數很少。那進入 埃及 地、在那裏寄居的，就是倖存的 猶大 人，必知道是誰的話站得住，是我的話呢，還是他們的話。
JER|44|29|我在這地方懲罰你們，必有預兆，使你們知道我降禍給你們的話必站得住。這是耶和華說的。
JER|44|30|耶和華如此說：看哪，我必將 埃及 王 合弗拉 法老交在他仇敵和尋索其命的人手中，像我將 猶大 王 西底家 交在他仇敵和尋索其命的 巴比倫 王 尼布甲尼撒 手中一樣。」
JER|45|1|約西亞 的兒子 猶大 王 約雅敬 第四年， 尼利亞 的兒子 巴錄 把 耶利米 先知口中所說的話寫在書上； 耶利米 對 巴錄 說：
JER|45|2|「 巴錄 啊，耶和華－ 以色列 的上帝說：
JER|45|3|你曾說：『哀哉！耶和華使我愁上加愁，我因呻吟而困乏，不得安歇。』
JER|45|4|你要這樣告訴他，耶和華如此說：看哪，我所建立的，我必拆毀；我所栽植的，我必拔出；在全地我都如此行。
JER|45|5|你為自己圖謀大事嗎？不要圖謀！看哪，我必使災禍臨到凡有血肉之軀的。但你無論往哪裏去，我要保全你的性命。這是耶和華說的。」
JER|46|1|耶和華論列國的話臨到 耶利米 先知。
JER|46|2|論到 埃及 ，關於 埃及 王 尼哥 法老的軍隊，這軍隊安營在 幼發拉底河 邊的 迦基米施 ，是 巴比倫 王 尼布甲尼撒 在 約西亞 的兒子 猶大 王 約雅敬 第四年所打敗的。
JER|46|3|你們要預備大小盾牌， 往前上陣，
JER|46|4|套上車， 騎上馬！ 頂盔站立， 磨槍披甲！
JER|46|5|我為何看見他們驚惶， 轉身退後呢？ 他們的勇士打敗仗， 急忙逃跑，並不回頭； 四圍都有驚嚇！ 這是耶和華說的。
JER|46|6|不要容快跑的逃避， 也不要容勇士逃脫 ； 在北方 幼發拉底河 邊， 他們絆跌仆倒。
JER|46|7|這是誰，像 尼羅河 漲溢， 如江河的水翻騰呢？
JER|46|8|埃及 像 尼羅河 漲溢， 如江河的水翻騰。 它說：「我要漲溢遮蓋全地； 我要毀滅城鎮和其中的居民。
JER|46|9|馬匹啊，上去吧！ 戰車啊，要疾行！ 手拿盾牌的 古實 和 弗 的勇士， 擅長拉弓的 路德 人，前進吧！」
JER|46|10|那日是萬軍之主耶和華報仇的日子， 要向敵人報仇。 刀劍必吞吃飽足， 飲血滿足； 因為在北方 幼發拉底河 邊， 有祭物獻給萬軍之主耶和華。
JER|46|11|少女 埃及 啊， 要上 基列 去取乳香； 你雖服用許多藥， 還是徒然，不得治好。
JER|46|12|列國聽見你的羞辱， 遍地滿了你的哀聲； 勇士與勇士彼此相撞， 二人一起跌倒。
JER|46|13|以下是耶和華對 耶利米 先知說的話，論到 巴比倫 王 尼布甲尼撒 要來攻擊 埃及 地。
JER|46|14|你們要在 埃及 傳揚，在 密奪 報告， 在 挪弗 、 答比匿 宣告說： 「要擺好陣勢，預備作戰， 因為刀劍在你四圍施行吞滅。」
JER|46|15|你的壯士為何被掃除呢？ 他們站立不住， 因為耶和華驅逐他們；
JER|46|16|他使多人絆跌，彼此撞倒。 他們說：「起來，讓我們回到自己的同胞、 回到自己的出生地去， 好躲避欺壓的刀劍。」
JER|46|17|他們在那裏稱 埃及 王法老 為 「錯失良機的誇大者」。
JER|46|18|名為萬軍之耶和華的君王說： 我指著我的永生起誓： 「 尼布甲尼撒 來的時候， 必像眾山之中的 他泊 ， 像海邊的 迦密 。」
JER|46|19|住在 埃及 的啊， 要預備被擄時需用的物品； 因為 挪弗 必成為廢墟， 被燒燬，無人居住。
JER|46|20|埃及 是肥美的母牛犢； 但來自北方的牛虻來到了！來到了！
JER|46|21|它的傭兵好像圈裏的肥牛犢， 他們轉身退後， 一齊逃跑，站立不住； 因為他們遭難的日子、 受罰的時刻已經來臨。
JER|46|22|它的聲音好像蛇在滑行。 敵人要成隊而來，如砍伐樹木的人， 手拿斧頭攻擊它。
JER|46|23|雖然它的樹林不易穿過， 敵人卻要砍伐， 因敵人比蝗蟲還多，不可勝數。 這是耶和華說的。
JER|46|24|埃及 必然蒙羞， 被交在北方人的手中。
JER|46|25|萬軍之耶和華－ 以色列 的上帝說：「看哪，我要懲罰 挪 的 亞捫 和法老、 埃及 和它的神明，以及君王，也要懲罰法老和倚靠他的人。
JER|46|26|我要將他們交給尋索其命之人的手和 巴比倫 王 尼布甲尼撒 與他臣僕的手。但 埃及 日後必再有人居住，與從前一樣。這是耶和華說的。」
JER|46|27|我的僕人 雅各 啊，不要懼怕！ 以色列 啊，不要驚惶！ 因我要從遠方拯救你， 從被擄之地拯救你的後裔。 雅各 必回來，得享平靜安逸， 無人令他害怕。
JER|46|28|我的僕人 雅各 啊，不要懼怕！ 因我與你同在。 我要將那些國滅絕淨盡， 就是我趕你去的那些國； 卻不將你滅絕淨盡， 倒要從寬懲治你， 但絕不能不罰你。 這是耶和華說的。
JER|47|1|在法老攻擊 迦薩 之前，耶和華論 非利士 人的話臨到 耶利米 先知。
JER|47|2|耶和華如此說： 看哪，有水從北方漲起，成為漲溢的河， 要淹沒全地和其中所充滿的， 淹沒城和城裏的居民。 人必呼喊， 境內的居民都必哀號。
JER|47|3|一聽見敵人壯馬蹄踏的響聲、 戰車隆隆、車輪轟轟， 為父的手就發軟， 不能回頭看顧兒女。
JER|47|4|因為日子將到， 耶和華必毀滅所有 非利士 人， 剪除 推羅 、 西頓 僅存的幫助者； 他要毀滅 非利士 人、 迦斐託 海島剩餘的人。
JER|47|5|迦薩 成了光禿， 亞實基倫 歸於無有。 平原 中所剩的啊， 你割劃自己，要到幾時呢？
JER|47|6|耶和華的刀劍哪，你要到幾時才止息呢？ 要入鞘，安靜不動。
JER|47|7|耶和華吩咐它攻擊 亞實基倫 和海邊之地， 既已派定它，你 怎能靜止不動呢？
JER|48|1|論 摩押 。 萬軍之耶和華－ 以色列 的上帝如此說： 禍哉， 尼波 ！它要變為廢墟。 基列亭 蒙羞被攻取， 米斯迦 蒙羞被毀壞，
JER|48|2|摩押 不再被稱讚。 有人在 希實本 設計謀害它： 「來吧！我們將它剪除，使它不再成國。」 瑪得緬 哪，你也必靜默無聲； 刀劍必追趕你。
JER|48|3|從 何羅念 有哀號聲： 「荒涼！大毀滅！」
JER|48|4|「 摩押 毀滅了！」 它的孩童哀號，使人聽見。
JER|48|5|人上 魯希坡 隨走隨哭， 因為在 何羅念 的下坡聽見毀滅的哀聲。
JER|48|6|你們要奔逃，自救己命， 使你們的性命如曠野裏的矮樹 。
JER|48|7|你因倚靠自己所做的 和自己的財寶，必被攻取。 基抹 和屬它的祭司、官長也要一同被擄去。
JER|48|8|那行毀滅的要來到各城， 並無一城倖免。 山谷必敗落， 平原必毀壞， 正如耶和華所說的。
JER|48|9|你們要將翅膀給 摩押 ， 使它可以飛去 。 它的城鎮必荒涼， 無人居住。
JER|48|10|懶惰不肯為耶和華做事的，必受詛咒；禁止刀劍不見血的，必受詛咒。
JER|48|11|摩押 自幼年以來常享安逸， 如沉澱未被攪動的酒 ， 沒有從這器皿倒在那器皿， 也未曾被擄掠過。 因此，它的原味尚存， 香氣未變。
JER|48|12|看哪，日子將到，我必差倒酒的到它那裏去，將它倒出來；他們要倒空器皿，打碎罈子。這是耶和華說的。
JER|48|13|摩押 必因 基抹 羞愧，像 以色列 家因倚靠 伯特利 羞愧一樣。
JER|48|14|你們怎麼說： 「我們是勇士，是會打仗的壯士」呢？
JER|48|15|摩押 變為廢墟， 敵人上去佔它的城鎮。 它精良的壯丁都下去遭殺戮； 這是名為萬軍之耶和華的君王說的。
JER|48|16|摩押 的災殃臨近， 災難速速來到。
JER|48|17|凡在它四圍的和認識它名的， 都要為它悲傷，說： 那結實的杖和美好的棍， 竟然折斷了！
JER|48|18|底本 的居民哪， 要從你榮耀的座位上下來， 坐著忍受乾渴； 因毀滅 摩押 的人上來攻擊你， 毀壞了你的堡壘。
JER|48|19|住 亞羅珥 的啊， 要站在道路的邊上觀望， 問逃跑的男人和逃脫的女人說： 「發生了甚麼事呢」？
JER|48|20|摩押 因毀壞蒙羞； 你們要哀號呼喊， 要在 亞嫩 報告： 「 摩押 已成廢墟！」
JER|48|21|審判臨到平原之地的 何倫 、 雅雜 、 米法押 、
JER|48|22|底本 、 尼波 、 伯‧低比拉太音 、
JER|48|23|基列亭 、 伯‧迦末 、 伯‧米恩 、
JER|48|24|加略 、 波斯拉 和 摩押 地遠近所有的城鎮。
JER|48|25|摩押 的角砍斷了，膀臂折斷了。這是耶和華說的。
JER|48|26|你們要使 摩押 沉醉，因它向耶和華誇大。它要在自己所吐之物中打滾，又要被人嗤笑。
JER|48|27|以色列 不是你的笑柄嗎？它難道是在賊中被逮到，使你每逢提到它就搖頭的嗎？
JER|48|28|摩押 的居民哪， 要離開城鎮，住在山崖裏， 像鴿子在峽谷口上搭窩。
JER|48|29|我們聽聞 摩押 人的驕傲， 極其驕傲； 他們自高、自傲、 自我狂妄、居心自大。
JER|48|30|我知道他們的憤怒是虛空的， 他們誇大的話一無所成。 這是耶和華說的。
JER|48|31|因此，我要為 摩押 哀號， 為 摩押 全地呼喊； 人必為 吉珥‧哈列設 人嘆息。
JER|48|32|西比瑪 的葡萄樹啊，我為你哀哭， 甚於 雅謝 人的哀哭。 你的枝子蔓延過海， 直伸到 雅謝海 。 那行毀滅的已經臨到你夏天的果子和葡萄。
JER|48|33|肥田和 摩押 地的歡喜快樂都被奪去， 我使酒池不再流出酒來， 無人踹酒歡呼； 呼喊的聲音不再是歡呼。
JER|48|34|有哀聲從 希實本 達到 以利亞利 ，他們發的哀聲達到 雅雜 ；從 瑣珥 達到 何羅念 ，達到 伊基拉‧施利施亞 ，因為 寧林 的水必然乾涸。
JER|48|35|我必在 摩押 地使那在丘壇獻祭的，和那向他的神明燒香的都滅絕了。這是耶和華說的。
JER|48|36|因此，我的心為 摩押 哀鳴如簫，我的心為 吉珥‧哈列設 人哀哭； 摩押 人所得的財物都毀滅了。
JER|48|37|各人頭上光禿，鬍鬚剪短，手有劃傷，腰束麻布。
JER|48|38|在 摩押 的各房頂上和街市上到處有人哀哭，因我打碎 摩押 ，好像打碎無人喜愛的器皿。這是耶和華說的。
JER|48|39|打得粉碎了！他們要哀號了！ 摩押 要羞愧轉背了！這樣， 摩押 必受四圍的人嗤笑驚駭。
JER|48|40|耶和華如此說： 看哪，仇敵必如鷹展翅快飛， 攻擊 摩押 。
JER|48|41|加略 被攻取，堡壘也被佔據。 到那日， 摩押 的勇士心中疼痛如臨產的婦人。
JER|48|42|摩押 必被毀滅，不再成國， 因它向耶和華誇大。
JER|48|43|摩押 的居民哪， 驚嚇、陷阱、羅網都臨近你。 這是耶和華說的。
JER|48|44|躲過驚嚇的必墜入陷阱， 逃離陷阱的又被羅網纏住， 因我必使懲罰之年臨到 摩押 。 這是耶和華說的。
JER|48|45|逃難的人站在 希實本 的蔭下，筋疲力盡， 因為有火從 希實本 發出， 有火焰出自 西宏 ， 燒盡 摩押 的鬢角和鬧鬨人的頭頂。
JER|48|46|摩押 啊，你有禍了！ 屬 基抹 的百姓滅亡了！ 因你的兒子都被擄去， 你的女兒也被擄去。
JER|48|47|到末後，我卻要使 摩押 被擄的人歸回。 摩押 受審判的話到此為止。 這是耶和華說的。
JER|49|1|論 亞捫 人。 耶和華如此說： 以色列 沒有兒子嗎？ 沒有後嗣嗎？ 米勒公 為何承受 迦得 為業呢？ 屬它的百姓為何住其中的城鎮呢？
JER|49|2|看哪，日子將到，我必使人聽見打仗的喊聲， 攻擊 亞捫 人所住的 拉巴 的喊聲。 拉巴 要成為廢墟， 屬它的鄉鎮 要被火焚燒。 這是耶和華說的。 先前承受 以色列 為業的， 此時 以色列 倒要承受他們為業。 這是耶和華說的。
JER|49|3|希實本 哪，要哀號， 因為 愛 地已成荒地。 拉巴 的鄉鎮哪，要呼喊， 以麻布束腰； 要哭號，在籬笆中往來奔跑； 因 米勒公 和它的祭司、 官長要一同被擄去。
JER|49|4|背道的民 哪， 你為何因有山谷， 因有水流的山谷誇耀呢？ 為何倚靠自己的財寶，說： 「誰能來到我們這裏呢？」
JER|49|5|萬軍之主耶和華說： 看哪，我要使驚嚇從四圍的鄰邦臨到你們； 你們必被趕出， 各人一直往前， 無人收容難民。
JER|49|6|但後來，我卻要使被擄的 亞捫 人歸回。這是耶和華說的。
JER|49|7|論 以東 。 萬軍之耶和華如此說： 提幔 不再有智慧了嗎？ 聰明人的謀略都用盡了嗎？ 他們的智慧盡歸無有了嗎？
JER|49|8|底但 的居民哪，要轉身逃跑， 住在深密處； 因為我懲罰 以掃 的時候， 必使災殃臨到他。
JER|49|9|摘葡萄的若來到你那裏， 豈不留下幾串嗎？ 賊若夜間來到， 豈不是只毀壞他們要毀壞的嗎？
JER|49|10|我卻使 以掃 赤裸， 暴露他的藏身處； 他不能隱藏自己。 他的後裔、弟兄、鄰舍全都滅絕， 他也歸於無有。
JER|49|11|你撇下孤兒，我必保全他們的性命； 你的寡婦可以倚靠我。
JER|49|12|耶和華如此說：「看哪，既然原不該喝那杯的一定要喝，你能免去懲罰嗎？必不能免，一定要喝！
JER|49|13|我指著自己起誓， 波斯拉 必令人驚駭、受羞辱、被詛咒，並且全然荒廢。它所有的城鎮都要永遠成為廢墟。這是耶和華說的。」
JER|49|14|我從耶和華那裏聽見消息， 有使者被差往列國去，說： 「你們要聚集前來攻擊 以東 ， 要起來爭戰。」
JER|49|15|看哪，我使你在列國中為最小， 在世人中被藐視。
JER|49|16|住在山穴中盤據山頂的啊， 你被自己的聲勢與心中的狂傲所蒙蔽； 你雖如大鷹高高搭窩， 我卻要從那裏拉你下來。 這是耶和華說的。
JER|49|17|以東 必令人驚駭；凡經過的人都驚駭，又因它一切的災禍嗤笑。
JER|49|18|耶和華說：它要像 所多瑪 、 蛾摩拉 和鄰近的城鎮一樣傾覆，必無人住在那裏，也無人在其中寄居。
JER|49|19|看哪，就像獅子從 約旦河 邊的叢林上來，攻擊堅固的居所，我要在轉眼之間使 以東 人逃跑，離開這地。我揀選誰，就派誰治理這地。誰能像我呢？誰能召我出庭呢？ 有哪一個牧人能在我面前站得住呢？
JER|49|20|你們要聽耶和華攻擊 以東 所定的計劃和他攻擊 提幔 居民所定的旨意。他們羊群當中微弱的定要被拖走，他們的草場定要變為荒涼。
JER|49|21|因他們仆倒的聲音，地就震動，哀號的聲音傳到 紅海 那裏。
JER|49|22|看哪，仇敵必如大鷹飛起，展開翅膀攻擊 波斯拉 。到那日， 以東 的勇士心中疼痛如臨產的婦人。
JER|49|23|論 大馬士革 。 哈馬 和 亞珥拔 蒙羞， 因為他們聽見兇惡的消息就融化； 焦慮像海浪洶湧，不得平靜。
JER|49|24|大馬士革 發軟，轉身逃跑； 戰兢將它捉住， 痛苦憂愁將它抓住， 如臨產的婦人一樣。
JER|49|25|我所喜樂受稱讚的城， 怎能被撇棄 呢？
JER|49|26|它的壯丁必仆倒在街上， 當那日，戰士全都靜默無聲。 這是萬軍之耶和華說的。
JER|49|27|我必用火點燃 大馬士革 的城牆， 燒滅 便‧哈達 的宮殿。
JER|49|28|論 巴比倫 王 尼布甲尼撒 所攻打的 基達 和 夏瑣 諸國。 耶和華如此說： 迦勒底 人哪，起來上 基達 去， 毀滅東方人。
JER|49|29|人要奪去他們的帳棚和羊群， 人要帶走他們的幔子、一切器皿，和駱駝，佔為己有。 人向他們喊著說： 四圍都有驚嚇。
JER|49|30|夏瑣 的居民哪，要逃奔遠方， 住在深遠之處； 因為 巴比倫 王 尼布甲尼撒 設計謀害你們， 起意攻擊你們。 這是耶和華說的。
JER|49|31|迦勒底 人哪，起來！ 上到安逸無慮的國民那裏去， 他們是無門無閂、單獨居住的。 這是耶和華說的。
JER|49|32|他們的駱駝必成為掠物， 他們眾多的牲畜必成為擄物。 我要將剃鬢髮的人分散四方 ， 使災殃從四圍臨到他們。 這是耶和華說的。
JER|49|33|夏瑣 必成為野狗的住處， 永遠荒廢； 無人住在那裏， 也無人在其中寄居。
JER|49|34|猶大 王 西底家 登基的時候，耶和華論 以攔 的話臨到 耶利米 先知，說：
JER|49|35|「萬軍之耶和華如此說：看哪，我必折斷 以攔 人的弓，那是他們戰鬥的主力。
JER|49|36|我要使風從天的四方颳來，臨到 以攔 ，將他們分散四方。 以攔 被趕散的人沒有一國不到的。
JER|49|37|我必使 以攔 人在仇敵和尋索其命的人面前驚惶；我也必使災禍，就是我的烈怒臨到他們，又必使刀劍追殺他們，直到將他們滅盡。這是耶和華說的。
JER|49|38|我要在 以攔 設立我的寶座，在那裏除滅君王和官長。這是耶和華說的。
JER|49|39|「到末後，我卻要使被擄的 以攔 人歸回。這是耶和華說的。」
JER|50|1|以下是耶和華藉 耶利米 先知論 巴比倫 和 迦勒底 人之地所說的話。
JER|50|2|你們要在萬國中傳揚，宣告， 豎立大旗； 要宣告，不可隱瞞，說： 「 巴比倫 被攻取， 彼勒 蒙羞， 米羅達 驚惶。 巴比倫 的神像都蒙羞， 它的偶像都驚惶。」
JER|50|3|因有一國從北方上來攻擊它，使它的地荒涼，無人居住，連人帶牲畜都逃走了。
JER|50|4|在那日、在那時， 以色列 人要和 猶大 人同來，隨走隨哭，尋求耶和華－他們的上帝。這是耶和華說的。
JER|50|5|他們要問到 錫安 之路，又面向那裏，說：「來吧，他們要 在永不被遺忘的約中與耶和華聯合。」
JER|50|6|我的百姓成了失喪的羊，牧人使他們走迷了路，轉入叢山之間。他們從大山走到小山，竟忘了自己安歇之處。
JER|50|7|凡遇見他們的，就把他們吞滅。敵人說：「我們不算有罪；因他們得罪了那可作真正 居所的耶和華，就是他們祖先所仰望的耶和華。」
JER|50|8|「你們要逃離 巴比倫 ，要離開 迦勒底 人之地，像走在羊群前面的公山羊。
JER|50|9|看哪，因我必激起大國聯盟，帶領他們從北方來攻擊 巴比倫 ，他們要擺陣攻擊它，它必在那裏被攻取。他們的箭好像善射 勇士的箭，絕不徒然返回。
JER|50|10|迦勒底 要成為掠物，凡擄掠它的都必心滿意足。這是耶和華說的。」
JER|50|11|搶奪我產業的啊， 你們因歡喜快樂， 像踹穀 嬉戲的母牛犢， 又像發嘶聲的壯馬。
JER|50|12|你們的母親極其抱愧， 生你們的必然蒙羞。 看哪，她要列在諸國之末， 成為曠野、旱地、沙漠；
JER|50|13|因耶和華的憤怒， 巴比倫 必無人居住， 全然荒涼， 凡經過的都要受驚駭， 又因它所遭的災殃嗤笑。
JER|50|14|所有拉弓的啊，要在 巴比倫 的四圍擺陣， 射箭攻擊它， 不用愛惜箭枝， 因為它得罪了耶和華。
JER|50|15|要在它四圍吶喊： 「它已經投降， 堡壘坍塌了， 城牆拆毀了！」 這是耶和華所報的仇。 你們要向它報仇； 它怎樣待人，你們也要怎樣待它。
JER|50|16|你們要將 巴比倫 撒種的 和收割時拿鐮刀的全都剪除。 他們各人因躲避欺壓的刀劍， 必歸回本族，逃到本土。
JER|50|17|以色列 是打散的羊，被獅子趕散。首先是 亞述 王將他吞滅，末後是 巴比倫 王 尼布甲尼撒 折斷他的骨頭。
JER|50|18|所以萬軍之耶和華－ 以色列 的上帝如此說：「看哪，我必懲罰 巴比倫 王和他的地，像我從前懲罰 亞述 王一樣。
JER|50|19|我必領 以色列 回他自己的草場，他要在 迦密 和 巴珊 吃草，又在 以法蓮 山上和 基列 境內得以飽足。
JER|50|20|在那日、在那時，你尋找 以色列 的罪孽，一無所有；尋找 猶大 的罪惡，也無所得；因為我所留下的人，我必赦免。這是耶和華說的。」
JER|50|21|你要上去攻擊 米拉大翁 之地， 又攻擊 比割 的居民。 將他們追殺滅盡， 照我所吩咐你的一切去做。 這是耶和華說的。
JER|50|22|境內有打仗和大毀滅的響聲。
JER|50|23|全地的大錘竟然砍斷破壞！ 巴比倫 在列國中竟然荒涼！
JER|50|24|巴比倫 哪，我為你設下羅網， 你被纏住，竟不自覺。 你被尋著，也被捉住， 因為你對抗耶和華。
JER|50|25|耶和華已經打開軍械庫， 拿出他惱恨的兵器； 這是萬軍之主耶和華 在 迦勒底 人之地要做的事。
JER|50|26|你們要從極遠的邊界前來攻擊它 ， 要開它的倉廩， 將它堆起如高堆， 毀滅淨盡，絲毫不留。
JER|50|27|要殺它一切的牛犢， 使牠們下去遭殺戮。 他們有禍了， 因為他們的日子，就是他們受罰的時刻已經來到。
JER|50|28|從 巴比倫 之地逃出來的難民，在 錫安 揚聲宣告耶和華－我們的上帝要報仇，為他的聖殿報仇。
JER|50|29|你們要招集一切弓箭手來攻擊 巴比倫 ，在 巴比倫 四圍安營，不容一人逃脫。要照著它所做的報應它；它怎樣待人，你們也要怎樣待它，因為它向耶和華－ 以色列 的聖者狂傲。
JER|50|30|所以它的壯丁必仆倒在街上。當那日，它的士兵全都靜默無聲。這是耶和華說的。
JER|50|31|「看哪，你這狂傲的啊，我與你為敵， 因為你的日子， 我懲罰你的時刻已經來到。 這是萬軍之主耶和華說的。
JER|50|32|狂傲的必絆跌仆倒，無人扶起。 我必用火點燃他的城鎮， 將他四圍所有的盡行燒滅。」
JER|50|33|萬軍之耶和華如此說：「 以色列 人和 猶大 人一同受欺壓；凡擄掠他們的都緊緊抓住他們，不肯釋放。
JER|50|34|他們的救贖主大有能力，萬軍之耶和華是他的名。他必定為他們伸冤，使全地得享平靜；他卻要攪擾 巴比倫 的居民。」
JER|50|35|有刀劍臨到 迦勒底 人和 巴比倫 的居民， 臨到它的領袖與智慧人。 這是耶和華說的。
JER|50|36|有刀劍臨到矜誇的人， 他們就變為愚昧； 有刀劍臨到它的勇士， 他們就驚惶。
JER|50|37|有刀劍臨到它的馬匹、戰車， 和其中混居的各族， 他們變成與婦女一樣； 有刀劍臨到它的寶物， 寶物就被搶奪。
JER|50|38|有乾旱 臨到它的眾水， 它們就必乾涸； 因為這是雕刻偶像之地， 人因偶像顛狂 。
JER|50|39|所以野獸和土狼必住在那裏，鴕鳥也住在其中，永遠無人居住，世世代代無人定居。
JER|50|40|巴比倫 要像上帝所傾覆的 所多瑪 、 蛾摩拉 和鄰近的城鎮一樣，必無人住在那裏，也無人在其中寄居。這是耶和華說的。
JER|50|41|看哪，有一民族從北方而來， 有一大國和許多君王被激起，從地極來到。
JER|50|42|他們拿弓和槍， 性情殘忍，毫不留情； 他們的聲音像海浪澎湃。 巴比倫 啊， 他們騎著馬， 如上戰場的人擺列隊伍， 要攻擊你。
JER|50|43|巴比倫 王聽見他們的風聲， 手就發軟， 痛苦將他抓住， 彷彿臨產的婦人疼痛一般。
JER|50|44|「看哪，就像獅子從 約旦河 邊的叢林上來，攻擊堅固的居所，我要在轉眼之間使 迦勒底 人逃跑，離開這地。我揀選誰，就派誰治理這地。誰能像我呢？誰能召我出庭呢？有哪一個牧人能在我面前站得住呢？
JER|50|45|你們要聽耶和華攻擊 巴比倫 所定的計劃和他攻擊 迦勒底 人之地所定的旨意。他們羊群當中微弱的定要被拖走，他們的草場定要變為荒涼。
JER|50|46|因 巴比倫 被攻下的聲音，地就震動，人在列國都聽見呼喊的聲音。」
JER|51|1|耶和華如此說： 看哪，我必颳起毀滅的風， 攻擊 巴比倫 和住在 立加米 的人。
JER|51|2|我要差陌生人 來到 巴比倫 ， 他們要簸揚它，使它的地空無一物。 在它遭禍的日子， 他們要四圍攻擊它。
JER|51|3|不要叫拉弓的拉弓， 不要叫他佩戴盔甲 ； 不要憐惜 巴比倫 的壯丁， 要滅盡它的全軍。
JER|51|4|他們必在 迦勒底 人之地被殺仆倒， 在 巴比倫 的街市上被刺透。
JER|51|5|以色列 和 猶大 境內雖然充滿違背 以色列 聖者的罪， 卻沒有被他的上帝－萬軍之耶和華所遺棄。
JER|51|6|你們要奔逃，離開 巴比倫 ， 各救自己的性命！ 不要陷在它的罪孽中一同滅亡， 因為這是耶和華報仇的時刻， 他必向 巴比倫 施行報應。
JER|51|7|巴比倫 素來是耶和華手中的金杯， 使全地沉醉， 列國喝了它的酒就顛狂。
JER|51|8|巴比倫 忽然傾覆毀壞； 要為它哀號， 拿乳香來止它的疼痛， 或者可以治好。
JER|51|9|我們想醫治 巴比倫 ， 它卻未獲痊癒。 離開它吧！讓我們各人歸回本國， 因為它受的審判通於上天，達到穹蒼。
JER|51|10|耶和華已經彰顯出我們的義。 來吧！我們要在 錫安 傳揚耶和華－我們上帝的作為。
JER|51|11|你們要磨尖箭頭， 抓住盾牌。 論到 巴比倫 ，耶和華定意要毀滅它，所以激起 瑪代 君王的心；這是耶和華報仇，為他的聖殿報仇。
JER|51|12|你們要豎立大旗， 攻擊 巴比倫 的城牆； 要堅固瞭望臺， 派定守望的設下埋伏； 因為耶和華指著 巴比倫 居民所說的， 他不但這樣定意，也已成就。
JER|51|13|住在眾水之上多有財寶的啊， 你的結局已到！ 你貪婪之量已滿盈 ！
JER|51|14|萬軍之耶和華指著自己起誓說： 我必使人遍滿各處像蝗蟲一樣， 他們必吶喊攻擊你。
JER|51|15|耶和華以能力創造大地， 以智慧建立世界， 以聰明鋪張穹蒼。
JER|51|16|他一出聲，天上就有眾水澎湃； 他使雲霧從地極上騰， 造電隨雨而閃， 從倉庫中吹出風來。
JER|51|17|人人都如同畜牲，毫無知識； 銀匠都因偶像羞愧， 他所鑄的偶像本為虛假， 它們裏面並無氣息。
JER|51|18|它們都是虛無的， 是迷惑人的東西， 到它們受罰的時刻必被除滅。
JER|51|19|雅各 所得的福分不是這樣， 因主 是那創造萬有的， 以色列 是他產業的支派， 萬軍之耶和華是他的名。
JER|51|20|你是我爭戰的斧子和打仗的兵器。 我要用你打碎列邦， 毀滅列國；
JER|51|21|用你打碎馬和騎馬的， 打碎戰車和坐在其上的；
JER|51|22|用你打碎男人和女人， 打碎老人和少年， 打碎壯丁和少女；
JER|51|23|用你打碎牧人和他的羊群， 打碎農夫和他的一對耕牛， 打碎省長和官員。
JER|51|24|我必在你們眼前報復 巴比倫 人和 迦勒底 居民在 錫安 所做的一切惡事。這是耶和華說的。
JER|51|25|行毀滅的山，看哪，我與你為敵， 你毀滅全地， 我必伸手攻擊你， 將你從山巖滾下去， 使你成為燒燬了的山。 這是耶和華說的。
JER|51|26|人必不從你那裏取石頭為房角石， 也不取石頭來作根基， 因為你必永遠荒廢。 這是耶和華說的。
JER|51|27|你們要在境內豎立大旗， 在列邦中吹角， 使列邦預備攻擊 巴比倫 。 要招集 亞拉臘 、 米尼 、 亞實基拿 各國前來攻擊它， 派將軍攻擊它， 使馬匹上來如粗暴的蝗蟲；
JER|51|28|使列邦和 瑪代 君王，省長和官員， 他們所管的全地，都預備攻擊它。
JER|51|29|地必震動而移轉； 因耶和華向 巴比倫 旨意已確定， 要使 巴比倫 土地荒涼，無人居住。
JER|51|30|巴比倫 的勇士停止爭戰， 躲在堡壘之中。 他們的力氣耗盡， 他們變成與婦女一樣。 巴比倫 的住處焚燒， 門閂都折斷了。
JER|51|31|通報的彼此相遇， 送信的彼此相遇， 報告 巴比倫 王， 城的四方都被攻下了，
JER|51|32|渡口被佔據了， 蘆葦被火焚燒， 戰士都驚慌。
JER|51|33|萬軍之耶和華－ 以色列 的上帝如此說： 巴比倫 好像踹穀的禾場； 再過片時，它收割的時候就到了。
JER|51|34|巴比倫 王 尼布甲尼撒 吞滅我，壓碎我， 使我成為空器皿。 他如大魚將我吞下， 以我的美物充滿他的肚腹， 又把我趕出去。
JER|51|35|錫安 的居民要說： 願我和我骨肉之親所受的殘暴 歸給 巴比倫 。 耶路撒冷 人要說： 願我們所流的血 歸給 迦勒底 的居民。
JER|51|36|所以，耶和華如此說： 看哪，我必為你伸冤，為你報仇； 我必使 巴比倫 的海枯竭， 使它的泉源乾涸。
JER|51|37|巴比倫 必成為廢墟， 為野狗的住處， 令人驚駭、嗤笑， 並且無人居住。
JER|51|38|他們要像少壯獅子一同咆哮， 像小獅子吼叫。
JER|51|39|他們食慾一來的時候， 我必為他們擺設酒席， 使他們沉醉，好叫他們快樂； 他們睡了長覺，永不醒起。 這是耶和華說的。
JER|51|40|我必使他們像羔羊、 像公綿羊和公山羊被牽去宰殺。
JER|51|41|示沙克 竟然被攻取！ 全地所稱讚的被佔據！ 巴比倫 在列國中竟然變為荒涼！
JER|51|42|海水漲起，漫過 巴比倫 ； 澎湃的海浪遮蓋了它。
JER|51|43|它的城鎮變廢墟， 地變乾旱，成為沙漠， 成為無人居住、 無人經過之地。
JER|51|44|我要懲罰 巴比倫 的 彼勒 ， 使它吐出所吞之物。 列國必不再流歸到它那裏， 巴比倫 的城牆也必坍塌。
JER|51|45|我的子民哪，你們要離開 巴比倫 ！ 各人逃命，躲避耶和華的烈怒。
JER|51|46|不要因境內所聽見的風聲 心驚膽怯或懼怕； 因為這年有風聲傳來， 那年也有風聲傳來； 境內有殘暴的事， 官長攻擊官長。
JER|51|47|所以，看哪，日子將到， 我必懲罰 巴比倫 雕刻的偶像。 它的全地必然抱愧， 它被殺的人必仆倒在其上。
JER|51|48|那時，天地和其中所有的， 必因 巴比倫 歡呼， 因為行毀滅的要從北方來到它那裏。 這是耶和華說的。
JER|51|49|巴比倫 要因 以色列 被殺的人而仆倒， 正如全地被刺殺的人是因 巴比倫 仆倒一般。
JER|51|50|你們躲避刀劍的要快走， 不要站住！ 要在遠方懷念耶和華， 心中追想 耶路撒冷 。
JER|51|51|我們聽見辱罵就蒙羞，滿面慚愧， 因為外邦人進入耶和華殿的聖所。
JER|51|52|所以，看哪，日子將到， 我必懲罰 巴比倫 雕刻的偶像， 在全境內到處都有刺傷的人在呻吟。 這是耶和華說的。
JER|51|53|巴比倫 雖升到天上， 雖使它堅固的高處更堅固， 我也要差毀滅者到它那裏。 這是耶和華說的。
JER|51|54|有哀號的聲音從 巴比倫 出來， 有大毀滅從 迦勒底 人之地而來。
JER|51|55|耶和華使 巴比倫 變為廢墟， 使其中喧嘩的大聲滅絕。 仇敵彷彿眾水， 波浪澎湃，發出響聲；
JER|51|56|這是行毀滅的臨到 巴比倫 。 巴比倫 的勇士被捉住， 他們的弓折斷了； 因為耶和華是施行報應的上帝， 他必施行報應。
JER|51|57|我必使 巴比倫 的領袖、 智慧人、省長、官員和勇士都喝醉， 使他們永遠沉睡，不再醒起。 這是名為萬軍之耶和華的君王說的。
JER|51|58|萬軍之耶和華如此說： 巴比倫 寬闊的城牆要夷為平地， 它高大的城門必被火焚燒。 萬民所勞碌的必致虛空， 萬族所勞碌的被火焚燒， 他們都必困乏。
JER|51|59|猶大 王 西底家 在位第四年， 瑪西雅 的孫子， 尼利亞 的兒子 西萊雅 與王同去 巴比倫 ， 西萊雅 是王宮的大臣， 耶利米 先知有話吩咐他。
JER|51|60|耶利米 把一切要臨到 巴比倫 的災禍，就是論到 巴比倫 的這一切話，寫在一書卷上。
JER|51|61|耶利米 對 西萊雅 說：「你到了 巴比倫 ，務要宣讀這一切話，
JER|51|62|說：『耶和華啊，你曾論到這地方說：要剪除它，不再有人與牲畜居住此地，必永遠荒涼。』
JER|51|63|你讀完這書卷，就要把一塊石頭拴在其上，投入 幼發拉底河 中，
JER|51|64|說：『 巴比倫 因耶和華所要降與它的災禍，必如此沉下去，不再浮起來，百姓也必困乏。』」 耶利米 的話到此為止。
JER|52|1|西底家 登基的時候年二十一歲，在 耶路撒冷 作王十一年。他母親名叫 哈慕她 ，是 立拿 人 耶利米 的女兒。
JER|52|2|西底家 行耶和華眼中看為惡的事，像 約雅敬 所做的一切。
JER|52|3|因此，耶和華向 耶路撒冷 和 猶大 發怒，以致把他們從自己面前趕出去。 西底家 背叛 巴比倫 王，
JER|52|4|他作王第九年十月初十， 巴比倫 王 尼布甲尼撒 率領全軍前來攻擊 耶路撒冷 ，對著城安營，四圍築堡壘攻城，
JER|52|5|城被圍困，直到 西底家 王十一年。
JER|52|6|四月初九，城裏的饑荒非常嚴重，當地的百姓都沒有糧食。
JER|52|7|城被攻破，士兵全都在夜間從靠近王園兩城牆中間的門逃跑出城； 迦勒底 人正在四圍攻城，他們就往 亞拉巴 逃去。
JER|52|8|迦勒底 的軍隊追趕 西底家 王，在 耶利哥 的平原追上他。他的全軍都離開他潰散了。
JER|52|9|迦勒底 人就拿住王，帶他到 哈馬 地 利比拉 的 巴比倫 王那裏； 巴比倫 王就判他的罪。
JER|52|10|巴比倫 王在 西底家 眼前殺了他的兒女，又在 利比拉 殺了 猶大 全體的官長，
JER|52|11|並且挖了 西底家 的眼睛，用銅鏈鎖著他，帶到 巴比倫 去，將他囚在監裏，直到他死的日子。
JER|52|12|巴比倫 王 尼布甲尼撒 十九年五月初十，在 巴比倫 王面前侍立的 尼布撒拉旦 護衛長進入 耶路撒冷 ，
JER|52|13|他焚燒了耶和華的殿、王宮和 耶路撒冷 的房屋；用火焚燒所有大戶人家的房屋。
JER|52|14|跟隨護衛長的 迦勒底 全軍拆毀了 耶路撒冷 四圍的城牆。
JER|52|15|那時 尼布撒拉旦 護衛長將百姓中最窮的和城裏所剩下的百姓，並那些投降 巴比倫 王的人，以及剩下的工匠，都擄去了。
JER|52|16|但 尼布撒拉旦 護衛長留下一些當地最窮的人，叫他們修整葡萄園，耕種田地。
JER|52|17|耶和華殿的銅柱並殿內的盆座和銅海， 迦勒底 人都打碎了，把那些銅運到 巴比倫 去；
JER|52|18|他們又帶走鍋、鏟子、鉗子、盤子、勺子，和供奉用的一切銅器；
JER|52|19|杯、火盆、碗、鍋、燈臺、勺子、酒杯，無論金的銀的，護衛長都帶走了；
JER|52|20|還有 所羅門 為耶和華殿所造的兩根柱子、一面銅海，並座下的十二隻銅牛，這些器皿的銅多得無法可秤。
JER|52|21|至於柱子，這一根柱子高十八肘，厚四指，周圍十二肘，中間是空的；
JER|52|22|柱上有銅頂，每個銅頂高五肘；銅頂的周圍有網子和石榴，也都是銅的。另一根柱子與此相同，也有石榴。
JER|52|23|柱子四面有九十六個石榴，在網子周圍，總共有一百個石榴。
JER|52|24|護衛長拿住 西萊雅 大祭司、 西番亞 副祭司和門口的三個守衛，
JER|52|25|又從城中拿住一個管理士兵的官 ，並在城裏找到王面前的七個親信，和召募當地百姓之將軍的書記官，以及在城中找到的六十個當地百姓。
JER|52|26|尼布撒拉旦 護衛長把這些人帶到 利比拉 的 巴比倫 王那裏。
JER|52|27|巴比倫 王擊殺他們，在 哈馬 地的 利比拉 把他們處死。這樣， 猶大 人就被擄去離開本地。
JER|52|28|這是 尼布甲尼撒 所擄百姓的數目：他在位第七年擄去 猶大 人三千零二十三人；
JER|52|29|尼布甲尼撒 十八年從 耶路撒冷 擄去八百三十二人；
JER|52|30|尼布甲尼撒 二十三年， 尼布撒拉旦 護衛長擄去 猶大 人七百四十五人；共有四千六百人。
JER|52|31|巴比倫 王 以未‧米羅達 作王的元年，就是 猶大 王 約雅斤 被擄後三十七年十二月二十五日，他使 猶大 王 約雅斤 抬起頭來，提他出監，
JER|52|32|對他說好話，使他的位高過與他一同被擄、在 巴比倫 眾王的位；
JER|52|33|又給他脫了囚服，使他終身常在 巴比倫 王面前吃飯。
JER|52|34|巴比倫 王賜給他日常需用的食物，日日一份，終身都是這樣，直到他死的日子。
