JUDG|1|1|After the death of Joshua, the Israelites asked the LORD, "Who will be the first to go up and fight for us against the Canaanites?"
JUDG|1|2|The LORD answered, "Judah is to go; I have given the land into their hands."
JUDG|1|3|Then the men of Judah said to the Simeonites their brothers, "Come up with us into the territory allotted to us, to fight against the Canaanites. We in turn will go with you into yours." So the Simeonites went with them.
JUDG|1|4|When Judah attacked, the LORD gave the Canaanites and Perizzites into their hands and they struck down ten thousand men at Bezek.
JUDG|1|5|It was there that they found Adoni-Bezek and fought against him, putting to rout the Canaanites and Perizzites.
JUDG|1|6|Adoni-Bezek fled, but they chased him and caught him, and cut off his thumbs and big toes.
JUDG|1|7|Then Adoni-Bezek said, "Seventy kings with their thumbs and big toes cut off have picked up scraps under my table. Now God has paid me back for what I did to them." They brought him to Jerusalem, and he died there.
JUDG|1|8|The men of Judah attacked Jerusalem also and took it. They put the city to the sword and set it on fire.
JUDG|1|9|After that, the men of Judah went down to fight against the Canaanites living in the hill country, the Negev and the western foothills.
JUDG|1|10|They advanced against the Canaanites living in Hebron (formerly called Kiriath Arba) and defeated Sheshai, Ahiman and Talmai.
JUDG|1|11|From there they advanced against the people living in Debir (formerly called Kiriath Sepher).
JUDG|1|12|And Caleb said, "I will give my daughter Acsah in marriage to the man who attacks and captures Kiriath Sepher."
JUDG|1|13|Othniel son of Kenaz, Caleb's younger brother, took it; so Caleb gave his daughter Acsah to him in marriage.
JUDG|1|14|One day when she came to Othniel, she urged him to ask her father for a field. When she got off her donkey, Caleb asked her, "What can I do for you?"
JUDG|1|15|She replied, "Do me a special favor. Since you have given me land in the Negev, give me also springs of water." Then Caleb gave her the upper and lower springs.
JUDG|1|16|The descendants of Moses' father-in-law, the Kenite, went up from the City of Palms with the men of Judah to live among the people of the Desert of Judah in the Negev near Arad.
JUDG|1|17|Then the men of Judah went with the Simeonites their brothers and attacked the Canaanites living in Zephath, and they totally destroyed the city. Therefore it was called Hormah.
JUDG|1|18|The men of Judah also took Gaza, Ashkelon and Ekron-each city with its territory.
JUDG|1|19|The LORD was with the men of Judah. They took possession of the hill country, but they were unable to drive the people from the plains, because they had iron chariots.
JUDG|1|20|As Moses had promised, Hebron was given to Caleb, who drove from it the three sons of Anak.
JUDG|1|21|The Benjamites, however, failed to dislodge the Jebusites, who were living in Jerusalem; to this day the Jebusites live there with the Benjamites.
JUDG|1|22|Now the house of Joseph attacked Bethel, and the LORD was with them.
JUDG|1|23|When they sent men to spy out Bethel (formerly called Luz),
JUDG|1|24|the spies saw a man coming out of the city and they said to him, "Show us how to get into the city and we will see that you are treated well."
JUDG|1|25|So he showed them, and they put the city to the sword but spared the man and his whole family.
JUDG|1|26|He then went to the land of the Hittites, where he built a city and called it Luz, which is its name to this day.
JUDG|1|27|But Manasseh did not drive out the people of Beth Shan or Taanach or Dor or Ibleam or Megiddo and their surrounding settlements, for the Canaanites were determined to live in that land.
JUDG|1|28|When Israel became strong, they pressed the Canaanites into forced labor but never drove them out completely.
JUDG|1|29|Nor did Ephraim drive out the Canaanites living in Gezer, but the Canaanites continued to live there among them.
JUDG|1|30|Neither did Zebulun drive out the Canaanites living in Kitron or Nahalol, who remained among them; but they did subject them to forced labor.
JUDG|1|31|Nor did Asher drive out those living in Acco or Sidon or Ahlab or Aczib or Helbah or Aphek or Rehob,
JUDG|1|32|and because of this the people of Asher lived among the Canaanite inhabitants of the land.
JUDG|1|33|Neither did Naphtali drive out those living in Beth Shemesh or Beth Anath; but the Naphtalites too lived among the Canaanite inhabitants of the land, and those living in Beth Shemesh and Beth Anath became forced laborers for them.
JUDG|1|34|The Amorites confined the Danites to the hill country, not allowing them to come down into the plain.
JUDG|1|35|And the Amorites were determined also to hold out in Mount Heres, Aijalon and Shaalbim, but when the power of the house of Joseph increased, they too were pressed into forced labor.
JUDG|1|36|The boundary of the Amorites was from Scorpion Pass to Sela and beyond.
JUDG|2|1|The angel of the LORD went up from Gilgal to Bokim and said, "I brought you up out of Egypt and led you into the land that I swore to give to your forefathers. I said, 'I will never break my covenant with you,
JUDG|2|2|and you shall not make a covenant with the people of this land, but you shall break down their altars.' Yet you have disobeyed me. Why have you done this?
JUDG|2|3|Now therefore I tell you that I will not drive them out before you; they will be thorns in your sides and their gods will be a snare to you."
JUDG|2|4|When the angel of the LORD had spoken these things to all the Israelites, the people wept aloud,
JUDG|2|5|and they called that place Bokim. There they offered sacrifices to the LORD.
JUDG|2|6|After Joshua had dismissed the Israelites, they went to take possession of the land, each to his own inheritance.
JUDG|2|7|The people served the LORD throughout the lifetime of Joshua and of the elders who outlived him and who had seen all the great things the LORD had done for Israel.
JUDG|2|8|Joshua son of Nun, the servant of the LORD, died at the age of a hundred and ten.
JUDG|2|9|And they buried him in the land of his inheritance, at Timnath Heres in the hill country of Ephraim, north of Mount Gaash.
JUDG|2|10|After that whole generation had been gathered to their fathers, another generation grew up, who knew neither the LORD nor what he had done for Israel.
JUDG|2|11|Then the Israelites did evil in the eyes of the LORD and served the Baals.
JUDG|2|12|They forsook the LORD, the God of their fathers, who had brought them out of Egypt. They followed and worshiped various gods of the peoples around them. They provoked the LORD to anger
JUDG|2|13|because they forsook him and served Baal and the Ashtoreths.
JUDG|2|14|In his anger against Israel the LORD handed them over to raiders who plundered them. He sold them to their enemies all around, whom they were no longer able to resist.
JUDG|2|15|Whenever Israel went out to fight, the hand of the LORD was against them to defeat them, just as he had sworn to them. They were in great distress.
JUDG|2|16|Then the LORD raised up judges, who saved them out of the hands of these raiders.
JUDG|2|17|Yet they would not listen to their judges but prostituted themselves to other gods and worshiped them. Unlike their fathers, they quickly turned from the way in which their fathers had walked, the way of obedience to the LORD 's commands.
JUDG|2|18|Whenever the LORD raised up a judge for them, he was with the judge and saved them out of the hands of their enemies as long as the judge lived; for the LORD had compassion on them as they groaned under those who oppressed and afflicted them.
JUDG|2|19|But when the judge died, the people returned to ways even more corrupt than those of their fathers, following other gods and serving and worshiping them. They refused to give up their evil practices and stubborn ways.
JUDG|2|20|Therefore the LORD was very angry with Israel and said, "Because this nation has violated the covenant that I laid down for their forefathers and has not listened to me,
JUDG|2|21|I will no longer drive out before them any of the nations Joshua left when he died.
JUDG|2|22|I will use them to test Israel and see whether they will keep the way of the LORD and walk in it as their forefathers did."
JUDG|2|23|The LORD had allowed those nations to remain; he did not drive them out at once by giving them into the hands of Joshua.
JUDG|3|1|These are the nations the LORD left to test all those Israelites who had not experienced any of the wars in Canaan
JUDG|3|2|(he did this only to teach warfare to the descendants of the Israelites who had not had previous battle experience):
JUDG|3|3|the five rulers of the Philistines, all the Canaanites, the Sidonians, and the Hivites living in the Lebanon mountains from Mount Baal Hermon to Lebo Hamath.
JUDG|3|4|They were left to test the Israelites to see whether they would obey the LORD 's commands, which he had given their forefathers through Moses.
JUDG|3|5|The Israelites lived among the Canaanites, Hittites, Amorites, Perizzites, Hivites and Jebusites.
JUDG|3|6|They took their daughters in marriage and gave their own daughters to their sons, and served their gods.
JUDG|3|7|The Israelites did evil in the eyes of the LORD; they forgot the LORD their God and served the Baals and the Asherahs.
JUDG|3|8|The anger of the LORD burned against Israel so that he sold them into the hands of Cushan-Rishathaim king of Aram Naharaim, to whom the Israelites were subject for eight years.
JUDG|3|9|But when they cried out to the LORD, he raised up for them a deliverer, Othniel son of Kenaz, Caleb's younger brother, who saved them.
JUDG|3|10|The Spirit of the LORD came upon him, so that he became Israel's judge and went to war. The LORD gave Cushan-Rishathaim king of Aram into the hands of Othniel, who overpowered him.
JUDG|3|11|So the land had peace for forty years, until Othniel son of Kenaz died.
JUDG|3|12|Once again the Israelites did evil in the eyes of the LORD, and because they did this evil the LORD gave Eglon king of Moab power over Israel.
JUDG|3|13|Getting the Ammonites and Amalekites to join him, Eglon came and attacked Israel, and they took possession of the City of Palms.
JUDG|3|14|The Israelites were subject to Eglon king of Moab for eighteen years.
JUDG|3|15|Again the Israelites cried out to the LORD, and he gave them a deliverer-Ehud, a left-handed man, the son of Gera the Benjamite. The Israelites sent him with tribute to Eglon king of Moab.
JUDG|3|16|Now Ehud had made a double-edged sword about a foot and a half long, which he strapped to his right thigh under his clothing.
JUDG|3|17|He presented the tribute to Eglon king of Moab, who was a very fat man.
JUDG|3|18|After Ehud had presented the tribute, he sent on their way the men who had carried it.
JUDG|3|19|At the idols near Gilgal he himself turned back and said, "I have a secret message for you, O king." The king said, "Quiet!" And all his attendants left him.
JUDG|3|20|Ehud then approached him while he was sitting alone in the upper room of his summer palace and said, "I have a message from God for you." As the king rose from his seat,
JUDG|3|21|Ehud reached with his left hand, drew the sword from his right thigh and plunged it into the king's belly.
JUDG|3|22|Even the handle sank in after the blade, which came out his back. Ehud did not pull the sword out, and the fat closed in over it.
JUDG|3|23|Then Ehud went out to the porch; he shut the doors of the upper room behind him and locked them.
JUDG|3|24|After he had gone, the servants came and found the doors of the upper room locked. They said, "He must be relieving himself in the inner room of the house."
JUDG|3|25|They waited to the point of embarrassment, but when he did not open the doors of the room, they took a key and unlocked them. There they saw their Lord fallen to the floor, dead.
JUDG|3|26|While they waited, Ehud got away. He passed by the idols and escaped to Seirah.
JUDG|3|27|When he arrived there, he blew a trumpet in the hill country of Ephraim, and the Israelites went down with him from the hills, with him leading them.
JUDG|3|28|"Follow me," he ordered, "for the LORD has given Moab, your enemy, into your hands." So they followed him down and, taking possession of the fords of the Jordan that led to Moab, they allowed no one to cross over.
JUDG|3|29|At that time they struck down about ten thousand Moabites, all vigorous and strong; not a man escaped.
JUDG|3|30|That day Moab was made subject to Israel, and the land had peace for eighty years.
JUDG|3|31|After Ehud came Shamgar son of Anath, who struck down six hundred Philistines with an oxgoad. He too saved Israel.
JUDG|4|1|After Ehud died, the Israelites once again did evil in the eyes of the LORD.
JUDG|4|2|So the LORD sold them into the hands of Jabin, a king of Canaan, who reigned in Hazor. The commander of his army was Sisera, who lived in Harosheth Haggoyim.
JUDG|4|3|Because he had nine hundred iron chariots and had cruelly oppressed the Israelites for twenty years, they cried to the LORD for help.
JUDG|4|4|Deborah, a prophetess, the wife of Lappidoth, was leading Israel at that time.
JUDG|4|5|She held court under the Palm of Deborah between Ramah and Bethel in the hill country of Ephraim, and the Israelites came to her to have their disputes decided.
JUDG|4|6|She sent for Barak son of Abinoam from Kedesh in Naphtali and said to him, "The LORD, the God of Israel, commands you: 'Go, take with you ten thousand men of Naphtali and Zebulun and lead the way to Mount Tabor.
JUDG|4|7|I will lure Sisera, the commander of Jabin's army, with his chariots and his troops to the Kishon River and give him into your hands.'"
JUDG|4|8|Barak said to her, "If you go with me, I will go; but if you don't go with me, I won't go."
JUDG|4|9|"Very well," Deborah said, "I will go with you. But because of the way you are going about this, the honor will not be yours, for the LORD will hand Sisera over to a woman." So Deborah went with Barak to Kedesh,
JUDG|4|10|where he summoned Zebulun and Naphtali. Ten thousand men followed him, and Deborah also went with him.
JUDG|4|11|Now Heber the Kenite had left the other Kenites, the descendants of Hobab, Moses' brother-in-law, and pitched his tent by the great tree in Zaanannim near Kedesh.
JUDG|4|12|When they told Sisera that Barak son of Abinoam had gone up to Mount Tabor,
JUDG|4|13|Sisera gathered together his nine hundred iron chariots and all the men with him, from Harosheth Haggoyim to the Kishon River.
JUDG|4|14|Then Deborah said to Barak, "Go! This is the day the LORD has given Sisera into your hands. Has not the LORD gone ahead of you?" So Barak went down Mount Tabor, followed by ten thousand men.
JUDG|4|15|At Barak's advance, the LORD routed Sisera and all his chariots and army by the sword, and Sisera abandoned his chariot and fled on foot.
JUDG|4|16|But Barak pursued the chariots and army as far as Harosheth Haggoyim. All the troops of Sisera fell by the sword; not a man was left.
JUDG|4|17|Sisera, however, fled on foot to the tent of Jael, the wife of Heber the Kenite, because there were friendly relations between Jabin king of Hazor and the clan of Heber the Kenite.
JUDG|4|18|Jael went out to meet Sisera and said to him, "Come, my Lord, come right in. Don't be afraid." So he entered her tent, and she put a covering over him.
JUDG|4|19|"I'm thirsty," he said. "Please give me some water." She opened a skin of milk, gave him a drink, and covered him up.
JUDG|4|20|"Stand in the doorway of the tent," he told her. "If someone comes by and asks you, 'Is anyone here?' say 'No.'"
JUDG|4|21|But Jael, Heber's wife, picked up a tent peg and a hammer and went quietly to him while he lay fast asleep, exhausted. She drove the peg through his temple into the ground, and he died.
JUDG|4|22|Barak came by in pursuit of Sisera, and Jael went out to meet him. "Come," she said, "I will show you the man you're looking for." So he went in with her, and there lay Sisera with the tent peg through his temple-dead.
JUDG|4|23|On that day God subdued Jabin, the Canaanite king, before the Israelites.
JUDG|4|24|And the hand of the Israelites grew stronger and stronger against Jabin, the Canaanite king, until they destroyed him.
JUDG|5|1|On that day Deborah and Barak son of Abinoam sang this song:
JUDG|5|2|"When the princes in Israel take the lead, when the people willingly offer themselves- praise the LORD!
JUDG|5|3|"Hear this, you kings! Listen, you rulers! I will sing to the LORD, I will sing; I will make music to the LORD, the God of Israel.
JUDG|5|4|"O LORD, when you went out from Seir, when you marched from the land of Edom, the earth shook, the heavens poured, the clouds poured down water.
JUDG|5|5|The mountains quaked before the LORD, the One of Sinai, before the LORD, the God of Israel.
JUDG|5|6|"In the days of Shamgar son of Anath, in the days of Jael, the roads were abandoned; travelers took to winding paths.
JUDG|5|7|Village life in Israel ceased, ceased until I, Deborah, arose, arose a mother in Israel.
JUDG|5|8|When they chose new gods, war came to the city gates, and not a shield or spear was seen among forty thousand in Israel.
JUDG|5|9|My heart is with Israel's princes, with the willing volunteers among the people. Praise the LORD!
JUDG|5|10|"You who ride on white donkeys, sitting on your saddle blankets, and you who walk along the road, consider
JUDG|5|11|the voice of the singers at the watering places. They recite the righteous acts of the LORD, the righteous acts of his warriors in Israel. "Then the people of the LORD went down to the city gates.
JUDG|5|12|'Wake up, wake up, Deborah! Wake up, wake up, break out in song! Arise, O Barak! Take captive your captives, O son of Abinoam.'
JUDG|5|13|"Then the men who were left came down to the nobles; the people of the LORD came to me with the mighty.
JUDG|5|14|Some came from Ephraim, whose roots were in Amalek; Benjamin was with the people who followed you. From Makir captains came down, from Zebulun those who bear a commander's staff.
JUDG|5|15|The princes of Issachar were with Deborah; yes, Issachar was with Barak, rushing after him into the valley. In the districts of Reuben there was much searching of heart.
JUDG|5|16|Why did you stay among the campfires to hear the whistling for the flocks? In the districts of Reuben there was much searching of heart.
JUDG|5|17|Gilead stayed beyond the Jordan. And Dan, why did he linger by the ships? Asher remained on the coast and stayed in his coves.
JUDG|5|18|The people of Zebulun risked their very lives; so did Naphtali on the heights of the field.
JUDG|5|19|"Kings came, they fought; the kings of Canaan fought at Taanach by the waters of Megiddo, but they carried off no silver, no plunder.
JUDG|5|20|From the heavens the stars fought, from their courses they fought against Sisera.
JUDG|5|21|The river Kishon swept them away, the age-old river, the river Kishon. March on, my soul; be strong!
JUDG|5|22|Then thundered the horses' hoofs- galloping, galloping go his mighty steeds.
JUDG|5|23|'Curse Meroz,' said the angel of the LORD. 'Curse its people bitterly, because they did not come to help the LORD, to help the LORD against the mighty.'
JUDG|5|24|"Most blessed of women be Jael, the wife of Heber the Kenite, most blessed of tent-dwelling women.
JUDG|5|25|He asked for water, and she gave him milk; in a bowl fit for nobles she brought him curdled milk.
JUDG|5|26|Her hand reached for the tent peg, her right hand for the workman's hammer. She struck Sisera, she crushed his head, she shattered and pierced his temple.
JUDG|5|27|At her feet he sank, he fell; there he lay. At her feet he sank, he fell; where he sank, there he fell-dead.
JUDG|5|28|"Through the window peered Sisera's mother; behind the lattice she cried out, 'Why is his chariot so long in coming? Why is the clatter of his chariots delayed?'
JUDG|5|29|The wisest of her ladies answer her; indeed, she keeps saying to herself,
JUDG|5|30|'Are they not finding and dividing the spoils: a girl or two for each man, colorful garments as plunder for Sisera, colorful garments embroidered, highly embroidered garments for my neck- all this as plunder?'
JUDG|5|31|"So may all your enemies perish, O LORD! But may they who love you be like the sun when it rises in its strength." Then the land had peace forty years.
JUDG|6|1|Again the Israelites did evil in the eyes of the LORD, and for seven years he gave them into the hands of the Midianites.
JUDG|6|2|Because the power of Midian was so oppressive, the Israelites prepared shelters for themselves in mountain clefts, caves and strongholds.
JUDG|6|3|Whenever the Israelites planted their crops, the Midianites, Amalekites and other eastern peoples invaded the country.
JUDG|6|4|They camped on the land and ruined the crops all the way to Gaza and did not spare a living thing for Israel, neither sheep nor cattle nor donkeys.
JUDG|6|5|They came up with their livestock and their tents like swarms of locusts. It was impossible to count the men and their camels; they invaded the land to ravage it.
JUDG|6|6|Midian so impoverished the Israelites that they cried out to the LORD for help.
JUDG|6|7|When the Israelites cried to the LORD because of Midian,
JUDG|6|8|he sent them a prophet, who said, "This is what the LORD, the God of Israel, says: I brought you up out of Egypt, out of the land of slavery.
JUDG|6|9|I snatched you from the power of Egypt and from the hand of all your oppressors. I drove them from before you and gave you their land.
JUDG|6|10|I said to you, 'I am the LORD your God; do not worship the gods of the Amorites, in whose land you live.' But you have not listened to me."
JUDG|6|11|The angel of the LORD came and sat down under the oak in Ophrah that belonged to Joash the Abiezrite, where his son Gideon was threshing wheat in a winepress to keep it from the Midianites.
JUDG|6|12|When the angel of the LORD appeared to Gideon, he said, "The LORD is with you, mighty warrior."
JUDG|6|13|"But sir," Gideon replied, "if the LORD is with us, why has all this happened to us? Where are all his wonders that our fathers told us about when they said, 'Did not the LORD bring us up out of Egypt?' But now the LORD has abandoned us and put us into the hand of Midian."
JUDG|6|14|The LORD turned to him and said, "Go in the strength you have and save Israel out of Midian's hand. Am I not sending you?"
JUDG|6|15|"But Lord, "Gideon asked, "how can I save Israel? My clan is the weakest in Manasseh, and I am the least in my family."
JUDG|6|16|The LORD answered, "I will be with you, and you will strike down all the Midianites together."
JUDG|6|17|Gideon replied, "If now I have found favor in your eyes, give me a sign that it is really you talking to me.
JUDG|6|18|Please do not go away until I come back and bring my offering and set it before you." And the LORD said, "I will wait until you return."
JUDG|6|19|Gideon went in, prepared a young goat, and from an ephah of flour he made bread without yeast. Putting the meat in a basket and its broth in a pot, he brought them out and offered them to him under the oak.
JUDG|6|20|The angel of God said to him, "Take the meat and the unleavened bread, place them on this rock, and pour out the broth." And Gideon did so.
JUDG|6|21|With the tip of the staff that was in his hand, the angel of the LORD touched the meat and the unleavened bread. Fire flared from the rock, consuming the meat and the bread. And the angel of the LORD disappeared.
JUDG|6|22|When Gideon realized that it was the angel of the LORD, he exclaimed, "Ah, Sovereign LORD! I have seen the angel of the LORD face to face!"
JUDG|6|23|But the LORD said to him, "Peace! Do not be afraid. You are not going to die."
JUDG|6|24|So Gideon built an altar to the LORD there and called it The LORD is Peace. To this day it stands in Ophrah of the Abiezrites.
JUDG|6|25|That same night the LORD said to him, "Take the second bull from your father's herd, the one seven years old. Tear down your father's altar to Baal and cut down the Asherah pole beside it.
JUDG|6|26|Then build a proper kind of altar to the LORD your God on the top of this height. Using the wood of the Asherah pole that you cut down, offer the second bull as a burnt offering."
JUDG|6|27|So Gideon took ten of his servants and did as the LORD told him. But because he was afraid of his family and the men of the town, he did it at night rather than in the daytime.
JUDG|6|28|In the morning when the men of the town got up, there was Baal's altar, demolished, with the Asherah pole beside it cut down and the second bull sacrificed on the newly built altar!
JUDG|6|29|They asked each other, "Who did this?" When they carefully investigated, they were told, "Gideon son of Joash did it."
JUDG|6|30|The men of the town demanded of Joash, "Bring out your son. He must die, because he has broken down Baal's altar and cut down the Asherah pole beside it."
JUDG|6|31|But Joash replied to the hostile crowd around him, "Are you going to plead Baal's cause? Are you trying to save him? Whoever fights for him shall be put to death by morning! If Baal really is a god, he can defend himself when someone breaks down his altar."
JUDG|6|32|So that day they called Gideon "Jerub-Baal, "saying, "Let Baal contend with him," because he broke down Baal's altar.
JUDG|6|33|Now all the Midianites, Amalekites and other eastern peoples joined forces and crossed over the Jordan and camped in the Valley of Jezreel.
JUDG|6|34|Then the Spirit of the LORD came upon Gideon, and he blew a trumpet, summoning the Abiezrites to follow him.
JUDG|6|35|He sent messengers throughout Manasseh, calling them to arms, and also into Asher, Zebulun and Naphtali, so that they too went up to meet them.
JUDG|6|36|Gideon said to God, "If you will save Israel by my hand as you have promised-
JUDG|6|37|look, I will place a wool fleece on the threshing floor. If there is dew only on the fleece and all the ground is dry, then I will know that you will save Israel by my hand, as you said."
JUDG|6|38|And that is what happened. Gideon rose early the next day; he squeezed the fleece and wrung out the dew-a bowlful of water.
JUDG|6|39|Then Gideon said to God, "Do not be angry with me. Let me make just one more request. Allow me one more test with the fleece. This time make the fleece dry and the ground covered with dew."
JUDG|6|40|That night God did so. Only the fleece was dry; all the ground was covered with dew.
JUDG|7|1|Early in the morning, Jerub-Baal (that is, Gideon) and all his men camped at the spring of Harod. The camp of Midian was north of them in the valley near the hill of Moreh.
JUDG|7|2|The LORD said to Gideon, "You have too many men for me to deliver Midian into their hands. In order that Israel may not boast against me that her own strength has saved her,
JUDG|7|3|announce now to the people, 'Anyone who trembles with fear may turn back and leave Mount Gilead.'" So twenty-two thousand men left, while ten thousand remained.
JUDG|7|4|But the LORD said to Gideon, "There are still too many men. Take them down to the water, and I will sift them for you there. If I say, 'This one shall go with you,' he shall go; but if I say, 'This one shall not go with you,' he shall not go."
JUDG|7|5|So Gideon took the men down to the water. There the LORD told him, "Separate those who lap the water with their tongues like a dog from those who kneel down to drink."
JUDG|7|6|Three hundred men lapped with their hands to their mouths. All the rest got down on their knees to drink.
JUDG|7|7|The LORD said to Gideon, "With the three hundred men that lapped I will save you and give the Midianites into your hands. Let all the other men go, each to his own place."
JUDG|7|8|So Gideon sent the rest of the Israelites to their tents but kept the three hundred, who took over the provisions and trumpets of the others. Now the camp of Midian lay below him in the valley.
JUDG|7|9|During that night the LORD said to Gideon, "Get up, go down against the camp, because I am going to give it into your hands.
JUDG|7|10|If you are afraid to attack, go down to the camp with your servant Purah
JUDG|7|11|and listen to what they are saying. Afterward, you will be encouraged to attack the camp." So he and Purah his servant went down to the outposts of the camp.
JUDG|7|12|The Midianites, the Amalekites and all the other eastern peoples had settled in the valley, thick as locusts. Their camels could no more be counted than the sand on the seashore.
JUDG|7|13|Gideon arrived just as a man was telling a friend his dream. "I had a dream," he was saying. "A round loaf of barley bread came tumbling into the Midianite camp. It struck the tent with such force that the tent overturned and collapsed."
JUDG|7|14|His friend responded, "This can be nothing other than the sword of Gideon son of Joash, the Israelite. God has given the Midianites and the whole camp into his hands."
JUDG|7|15|When Gideon heard the dream and its interpretation, he worshiped God. He returned to the camp of Israel and called out, "Get up! The LORD has given the Midianite camp into your hands."
JUDG|7|16|Dividing the three hundred men into three companies, he placed trumpets and empty jars in the hands of all of them, with torches inside.
JUDG|7|17|"Watch me," he told them. "Follow my lead. When I get to the edge of the camp, do exactly as I do.
JUDG|7|18|When I and all who are with me blow our trumpets, then from all around the camp blow yours and shout, 'For the LORD and for Gideon.'"
JUDG|7|19|Gideon and the hundred men with him reached the edge of the camp at the beginning of the middle watch, just after they had changed the guard. They blew their trumpets and broke the jars that were in their hands.
JUDG|7|20|The three companies blew the trumpets and smashed the jars. Grasping the torches in their left hands and holding in their right hands the trumpets they were to blow, they shouted, "A sword for the LORD and for Gideon!"
JUDG|7|21|While each man held his position around the camp, all the Midianites ran, crying out as they fled.
JUDG|7|22|When the three hundred trumpets sounded, the LORD caused the men throughout the camp to turn on each other with their swords. The army fled to Beth Shittah toward Zererah as far as the border of Abel Meholah near Tabbath.
JUDG|7|23|Israelites from Naphtali, Asher and all Manasseh were called out, and they pursued the Midianites.
JUDG|7|24|Gideon sent messengers throughout the hill country of Ephraim, saying, "Come down against the Midianites and seize the waters of the Jordan ahead of them as far as Beth Barah." So all the men of Ephraim were called out and they took the waters of the Jordan as far as Beth Barah.
JUDG|7|25|They also captured two of the Midianite leaders, Oreb and Zeeb. They killed Oreb at the rock of Oreb, and Zeeb at the winepress of Zeeb. They pursued the Midianites and brought the heads of Oreb and Zeeb to Gideon, who was by the Jordan.
JUDG|8|1|Now the Ephraimites asked Gideon, "Why have you treated us like this? Why didn't you call us when you went to fight Midian?" And they criticized him sharply.
JUDG|8|2|But he answered them, "What have I accomplished compared to you? Aren't the gleanings of Ephraim's grapes better than the full grape harvest of Abiezer?
JUDG|8|3|God gave Oreb and Zeeb, the Midianite leaders, into your hands. What was I able to do compared to you?" At this, their resentment against him subsided.
JUDG|8|4|Gideon and his three hundred men, exhausted yet keeping up the pursuit, came to the Jordan and crossed it.
JUDG|8|5|He said to the men of Succoth, "Give my troops some bread; they are worn out, and I am still pursuing Zebah and Zalmunna, the kings of Midian."
JUDG|8|6|But the officials of Succoth said, "Do you already have the hands of Zebah and Zalmunna in your possession? Why should we give bread to your troops?"
JUDG|8|7|Then Gideon replied, "Just for that, when the LORD has given Zebah and Zalmunna into my hand, I will tear your flesh with desert thorns and briers."
JUDG|8|8|From there he went up to Peniel and made the same request of them, but they answered as the men of Succoth had.
JUDG|8|9|So he said to the men of Peniel, "When I return in triumph, I will tear down this tower."
JUDG|8|10|Now Zebah and Zalmunna were in Karkor with a force of about fifteen thousand men, all that were left of the armies of the eastern peoples; a hundred and twenty thousand swordsmen had fallen.
JUDG|8|11|Gideon went up by the route of the nomads east of Nobah and Jogbehah and fell upon the unsuspecting army.
JUDG|8|12|Zebah and Zalmunna, the two kings of Midian, fled, but he pursued them and captured them, routing their entire army.
JUDG|8|13|Gideon son of Joash then returned from the battle by the Pass of Heres.
JUDG|8|14|He caught a young man of Succoth and questioned him, and the young man wrote down for him the names of the seventy-seven officials of Succoth, the elders of the town.
JUDG|8|15|Then Gideon came and said to the men of Succoth, "Here are Zebah and Zalmunna, about whom you taunted me by saying, 'Do you already have the hands of Zebah and Zalmunna in your possession? Why should we give bread to your exhausted men?'"
JUDG|8|16|He took the elders of the town and taught the men of Succoth a lesson by punishing them with desert thorns and briers.
JUDG|8|17|He also pulled down the tower of Peniel and killed the men of the town.
JUDG|8|18|Then he asked Zebah and Zalmunna, "What kind of men did you kill at Tabor?Men like you," they answered, "each one with the bearing of a prince."
JUDG|8|19|Gideon replied, "Those were my brothers, the sons of my own mother. As surely as the LORD lives, if you had spared their lives, I would not kill you."
JUDG|8|20|Turning to Jether, his oldest son, he said, "Kill them!" But Jether did not draw his sword, because he was only a boy and was afraid.
JUDG|8|21|Zebah and Zalmunna said, "Come, do it yourself. 'As is the man, so is his strength.'" So Gideon stepped forward and killed them, and took the ornaments off their camels' necks.
JUDG|8|22|The Israelites said to Gideon, "Rule over us-you, your son and your grandson-because you have saved us out of the hand of Midian."
JUDG|8|23|But Gideon told them, "I will not rule over you, nor will my son rule over you. The LORD will rule over you."
JUDG|8|24|And he said, "I do have one request, that each of you give me an earring from your share of the plunder." (It was the custom of the Ishmaelites to wear gold earrings.)
JUDG|8|25|They answered, "We'll be glad to give them." So they spread out a garment, and each man threw a ring from his plunder onto it.
JUDG|8|26|The weight of the gold rings he asked for came to seventeen hundred shekels, not counting the ornaments, the pendants and the purple garments worn by the kings of Midian or the chains that were on their camels' necks.
JUDG|8|27|Gideon made the gold into an ephod, which he placed in Ophrah, his town. All Israel prostituted themselves by worshiping it there, and it became a snare to Gideon and his family.
JUDG|8|28|Thus Midian was subdued before the Israelites and did not raise its head again. During Gideon's lifetime, the land enjoyed peace forty years.
JUDG|8|29|Jerub-Baal son of Joash went back home to live.
JUDG|8|30|He had seventy sons of his own, for he had many wives.
JUDG|8|31|His concubine, who lived in Shechem, also bore him a son, whom he named Abimelech.
JUDG|8|32|Gideon son of Joash died at a good old age and was buried in the tomb of his father Joash in Ophrah of the Abiezrites.
JUDG|8|33|No sooner had Gideon died than the Israelites again prostituted themselves to the Baals. They set up Baal-Berith as their god and
JUDG|8|34|did not remember the LORD their God, who had rescued them from the hands of all their enemies on every side.
JUDG|8|35|They also failed to show kindness to the family of Jerub-Baal (that is, Gideon) for all the good things he had done for them.
JUDG|9|1|Abimelech son of Jerub-Baal went to his mother's brothers in Shechem and said to them and to all his mother's clan,
JUDG|9|2|"Ask all the citizens of Shechem, 'Which is better for you: to have all seventy of Jerub-Baal's sons rule over you, or just one man?' Remember, I am your flesh and blood."
JUDG|9|3|When the brothers repeated all this to the citizens of Shechem, they were inclined to follow Abimelech, for they said, "He is our brother."
JUDG|9|4|They gave him seventy shekels of silver from the temple of Baal-Berith, and Abimelech used it to hire reckless adventurers, who became his followers.
JUDG|9|5|He went to his father's home in Ophrah and on one stone murdered his seventy brothers, the sons of Jerub-Baal. But Jotham, the youngest son of Jerub-Baal, escaped by hiding.
JUDG|9|6|Then all the citizens of Shechem and Beth Millo gathered beside the great tree at the pillar in Shechem to crown Abimelech king.
JUDG|9|7|When Jotham was told about this, he climbed up on the top of Mount Gerizim and shouted to them, "Listen to me, citizens of Shechem, so that God may listen to you.
JUDG|9|8|One day the trees went out to anoint a king for themselves. They said to the olive tree, 'Be our king.'
JUDG|9|9|"But the olive tree answered, 'Should I give up my oil, by which both gods and men are honored, to hold sway over the trees?'
JUDG|9|10|"Next, the trees said to the fig tree, 'Come and be our king.'
JUDG|9|11|"But the fig tree replied, 'Should I give up my fruit, so good and sweet, to hold sway over the trees?'
JUDG|9|12|"Then the trees said to the vine, 'Come and be our king.'
JUDG|9|13|"But the vine answered, 'Should I give up my wine, which cheers both gods and men, to hold sway over the trees?'
JUDG|9|14|"Finally all the trees said to the thornbush, 'Come and be our king.'
JUDG|9|15|"The thornbush said to the trees, 'If you really want to anoint me king over you, come and take refuge in my shade; but if not, then let fire come out of the thornbush and consume the cedars of Lebanon!'
JUDG|9|16|"Now if you have acted honorably and in good faith when you made Abimelech king, and if you have been fair to Jerub-Baal and his family, and if you have treated him as he deserves-
JUDG|9|17|and to think that my father fought for you, risked his life to rescue you from the hand of Midian
JUDG|9|18|(but today you have revolted against my father's family, murdered his seventy sons on a single stone, and made Abimelech, the son of his slave girl, king over the citizens of Shechem because he is your brother)-
JUDG|9|19|if then you have acted honorably and in good faith toward Jerub-Baal and his family today, may Abimelech be your joy, and may you be his, too!
JUDG|9|20|But if you have not, let fire come out from Abimelech and consume you, citizens of Shechem and Beth Millo, and let fire come out from you, citizens of Shechem and Beth Millo, and consume Abimelech!"
JUDG|9|21|Then Jotham fled, escaping to Beer, and he lived there because he was afraid of his brother Abimelech.
JUDG|9|22|After Abimelech had governed Israel three years,
JUDG|9|23|God sent an evil spirit between Abimelech and the citizens of Shechem, who acted treacherously against Abimelech.
JUDG|9|24|God did this in order that the crime against Jerub-Baal's seventy sons, the shedding of their blood, might be avenged on their brother Abimelech and on the citizens of Shechem, who had helped him murder his brothers.
JUDG|9|25|In opposition to him these citizens of Shechem set men on the hilltops to ambush and rob everyone who passed by, and this was reported to Abimelech.
JUDG|9|26|Now Gaal son of Ebed moved with his brothers into Shechem, and its citizens put their confidence in him.
JUDG|9|27|After they had gone out into the fields and gathered the grapes and trodden them, they held a festival in the temple of their god. While they were eating and drinking, they cursed Abimelech.
JUDG|9|28|Then Gaal son of Ebed said, "Who is Abimelech, and who is Shechem, that we should be subject to him? Isn't he Jerub-Baal's son, and isn't Zebul his deputy? Serve the men of Hamor, Shechem's father! Why should we serve Abimelech?
JUDG|9|29|If only this people were under my command! Then I would get rid of him. I would say to Abimelech, 'Call out your whole army!'"
JUDG|9|30|When Zebul the governor of the city heard what Gaal son of Ebed said, he was very angry.
JUDG|9|31|Under cover he sent messengers to Abimelech, saying, "Gaal son of Ebed and his brothers have come to Shechem and are stirring up the city against you.
JUDG|9|32|Now then, during the night you and your men should come and lie in wait in the fields.
JUDG|9|33|In the morning at sunrise, advance against the city. When Gaal and his men come out against you, do whatever your hand finds to do."
JUDG|9|34|So Abimelech and all his troops set out by night and took up concealed positions near Shechem in four companies.
JUDG|9|35|Now Gaal son of Ebed had gone out and was standing at the entrance to the city gate just as Abimelech and his soldiers came out from their hiding place.
JUDG|9|36|When Gaal saw them, he said to Zebul, "Look, people are coming down from the tops of the mountains!" Zebul replied, "You mistake the shadows of the mountains for men."
JUDG|9|37|But Gaal spoke up again: "Look, people are coming down from the center of the land, and a company is coming from the direction of the soothsayers' tree."
JUDG|9|38|Then Zebul said to him, "Where is your big talk now, you who said, 'Who is Abimelech that we should be subject to him?' Aren't these the men you ridiculed? Go out and fight them!"
JUDG|9|39|So Gaal led out the citizens of Shechem and fought Abimelech.
JUDG|9|40|Abimelech chased him, and many fell wounded in the flight-all the way to the entrance to the gate.
JUDG|9|41|Abimelech stayed in Arumah, and Zebul drove Gaal and his brothers out of Shechem.
JUDG|9|42|The next day the people of Shechem went out to the fields, and this was reported to Abimelech.
JUDG|9|43|So he took his men, divided them into three companies and set an ambush in the fields. When he saw the people coming out of the city, he rose to attack them.
JUDG|9|44|Abimelech and the companies with him rushed forward to a position at the entrance to the city gate. Then two companies rushed upon those in the fields and struck them down.
JUDG|9|45|All that day Abimelech pressed his attack against the city until he had captured it and killed its people. Then he destroyed the city and scattered salt over it.
JUDG|9|46|On hearing this, the citizens in the tower of Shechem went into the stronghold of the temple of El-Berith.
JUDG|9|47|When Abimelech heard that they had assembled there,
JUDG|9|48|he and all his men went up Mount Zalmon. He took an ax and cut off some branches, which he lifted to his shoulders. He ordered the men with him, "Quick! Do what you have seen me do!"
JUDG|9|49|So all the men cut branches and followed Abimelech. They piled them against the stronghold and set it on fire over the people inside. So all the people in the tower of Shechem, about a thousand men and women, also died.
JUDG|9|50|Next Abimelech went to Thebez and besieged it and captured it.
JUDG|9|51|Inside the city, however, was a strong tower, to which all the men and women-all the people of the city-fled. They locked themselves in and climbed up on the tower roof.
JUDG|9|52|Abimelech went to the tower and stormed it. But as he approached the entrance to the tower to set it on fire,
JUDG|9|53|a woman dropped an upper millstone on his head and cracked his skull.
JUDG|9|54|Hurriedly he called to his armor-bearer, "Draw your sword and kill me, so that they can't say, 'A woman killed him.'" So his servant ran him through, and he died.
JUDG|9|55|When the Israelites saw that Abimelech was dead, they went home.
JUDG|9|56|Thus God repaid the wickedness that Abimelech had done to his father by murdering his seventy brothers.
JUDG|9|57|God also made the men of Shechem pay for all their wickedness. The curse of Jotham son of Jerub-Baal came on them.
JUDG|10|1|After the time of Abimelech a man of Issachar, Tola son of Puah, the son of Dodo, rose to save Israel. He lived in Shamir, in the hill country of Ephraim.
JUDG|10|2|He led Israel twenty-three years; then he died, and was buried in Shamir.
JUDG|10|3|He was followed by Jair of Gilead, who led Israel twenty-two years.
JUDG|10|4|He had thirty sons, who rode thirty donkeys. They controlled thirty towns in Gilead, which to this day are called Havvoth Jair.
JUDG|10|5|When Jair died, he was buried in Kamon.
JUDG|10|6|Again the Israelites did evil in the eyes of the LORD. They served the Baals and the Ashtoreths, and the gods of Aram, the gods of Sidon, the gods of Moab, the gods of the Ammonites and the gods of the Philistines. And because the Israelites forsook the LORD and no longer served him,
JUDG|10|7|he became angry with them. He sold them into the hands of the Philistines and the Ammonites,
JUDG|10|8|who that year shattered and crushed them. For eighteen years they oppressed all the Israelites on the east side of the Jordan in Gilead, the land of the Amorites.
JUDG|10|9|The Ammonites also crossed the Jordan to fight against Judah, Benjamin and the house of Ephraim; and Israel was in great distress.
JUDG|10|10|Then the Israelites cried out to the LORD, "We have sinned against you, forsaking our God and serving the Baals."
JUDG|10|11|The LORD replied, "When the Egyptians, the Amorites, the Ammonites, the Philistines,
JUDG|10|12|the Sidonians, the Amalekites and the Maonites oppressed you and you cried to me for help, did I not save you from their hands?
JUDG|10|13|But you have forsaken me and served other gods, so I will no longer save you.
JUDG|10|14|Go and cry out to the gods you have chosen. Let them save you when you are in trouble!"
JUDG|10|15|But the Israelites said to the LORD, "We have sinned. Do with us whatever you think best, but please rescue us now."
JUDG|10|16|Then they got rid of the foreign gods among them and served the LORD. And he could bear Israel's misery no longer.
JUDG|10|17|When the Ammonites were called to arms and camped in Gilead, the Israelites assembled and camped at Mizpah.
JUDG|10|18|The leaders of the people of Gilead said to each other, "Whoever will launch the attack against the Ammonites will be the head of all those living in Gilead."
JUDG|11|1|Jephthah the Gileadite was a mighty warrior. His father was Gilead; his mother was a prostitute.
JUDG|11|2|Gilead's wife also bore him sons, and when they were grown up, they drove Jephthah away. "You are not going to get any inheritance in our family," they said, "because you are the son of another woman."
JUDG|11|3|So Jephthah fled from his brothers and settled in the land of Tob, where a group of adventurers gathered around him and followed him.
JUDG|11|4|Some time later, when the Ammonites made war on Israel,
JUDG|11|5|the elders of Gilead went to get Jephthah from the land of Tob.
JUDG|11|6|"Come," they said, "be our commander, so we can fight the Ammonites."
JUDG|11|7|Jephthah said to them, "Didn't you hate me and drive me from my father's house? Why do you come to me now, when you're in trouble?"
JUDG|11|8|The elders of Gilead said to him, "Nevertheless, we are turning to you now; come with us to fight the Ammonites, and you will be our head over all who live in Gilead."
JUDG|11|9|Jephthah answered, "Suppose you take me back to fight the Ammonites and the LORD gives them to me-will I really be your head?"
JUDG|11|10|The elders of Gilead replied, "The LORD is our witness; we will certainly do as you say."
JUDG|11|11|So Jephthah went with the elders of Gilead, and the people made him head and commander over them. And he repeated all his words before the LORD in Mizpah.
JUDG|11|12|Then Jephthah sent messengers to the Ammonite king with the question: "What do you have against us that you have attacked our country?"
JUDG|11|13|The king of the Ammonites answered Jephthah's messengers, "When Israel came up out of Egypt, they took away my land from the Arnon to the Jabbok, all the way to the Jordan. Now give it back peaceably."
JUDG|11|14|Jephthah sent back messengers to the Ammonite king,
JUDG|11|15|saying: "This is what Jephthah says: Israel did not take the land of Moab or the land of the Ammonites.
JUDG|11|16|But when they came up out of Egypt, Israel went through the desert to the Red Sea and on to Kadesh.
JUDG|11|17|Then Israel sent messengers to the king of Edom, saying, 'Give us permission to go through your country,' but the king of Edom would not listen. They sent also to the king of Moab, and he refused. So Israel stayed at Kadesh.
JUDG|11|18|"Next they traveled through the desert, skirted the lands of Edom and Moab, passed along the eastern side of the country of Moab, and camped on the other side of the Arnon. They did not enter the territory of Moab, for the Arnon was its border.
JUDG|11|19|"Then Israel sent messengers to Sihon king of the Amorites, who ruled in Heshbon, and said to him, 'Let us pass through your country to our own place.'
JUDG|11|20|Sihon, however, did not trust Israel to pass through his territory. He mustered all his men and encamped at Jahaz and fought with Israel.
JUDG|11|21|"Then the LORD, the God of Israel, gave Sihon and all his men into Israel's hands, and they defeated them. Israel took over all the land of the Amorites who lived in that country,
JUDG|11|22|capturing all of it from the Arnon to the Jabbok and from the desert to the Jordan.
JUDG|11|23|"Now since the LORD, the God of Israel, has driven the Amorites out before his people Israel, what right have you to take it over?
JUDG|11|24|Will you not take what your god Chemosh gives you? Likewise, whatever the LORD our God has given us, we will possess.
JUDG|11|25|Are you better than Balak son of Zippor, king of Moab? Did he ever quarrel with Israel or fight with them?
JUDG|11|26|For three hundred years Israel occupied Heshbon, Aroer, the surrounding settlements and all the towns along the Arnon. Why didn't you retake them during that time?
JUDG|11|27|I have not wronged you, but you are doing me wrong by waging war against me. Let the LORD, the Judge, decide the dispute this day between the Israelites and the Ammonites."
JUDG|11|28|The king of Ammon, however, paid no attention to the message Jephthah sent him.
JUDG|11|29|Then the Spirit of the LORD came upon Jephthah. He crossed Gilead and Manasseh, passed through Mizpah of Gilead, and from there he advanced against the Ammonites.
JUDG|11|30|And Jephthah made a vow to the LORD: "If you give the Ammonites into my hands,
JUDG|11|31|whatever comes out of the door of my house to meet me when I return in triumph from the Ammonites will be the LORD 's, and I will sacrifice it as a burnt offering."
JUDG|11|32|Then Jephthah went over to fight the Ammonites, and the LORD gave them into his hands.
JUDG|11|33|He devastated twenty towns from Aroer to the vicinity of Minnith, as far as Abel Keramim. Thus Israel subdued Ammon.
JUDG|11|34|When Jephthah returned to his home in Mizpah, who should come out to meet him but his daughter, dancing to the sound of tambourines! She was an only child. Except for her he had neither son nor daughter.
JUDG|11|35|When he saw her, he tore his clothes and cried, "Oh! My daughter! You have made me miserable and wretched, because I have made a vow to the LORD that I cannot break."
JUDG|11|36|"My father," she replied, "you have given your word to the LORD. Do to me just as you promised, now that the LORD has avenged you of your enemies, the Ammonites.
JUDG|11|37|But grant me this one request," she said. "Give me two months to roam the hills and weep with my friends, because I will never marry."
JUDG|11|38|"You may go," he said. And he let her go for two months. She and the girls went into the hills and wept because she would never marry.
JUDG|11|39|After the two months, she returned to her father and he did to her as he had vowed. And she was a virgin. From this comes the Israelite custom
JUDG|11|40|that each year the young women of Israel go out for four days to commemorate the daughter of Jephthah the Gileadite.
JUDG|12|1|The men of Ephraim called out their forces, crossed over to Zaphon and said to Jephthah, "Why did you go to fight the Ammonites without calling us to go with you? We're going to burn down your house over your head."
JUDG|12|2|Jephthah answered, "I and my people were engaged in a great struggle with the Ammonites, and although I called, you didn't save me out of their hands.
JUDG|12|3|When I saw that you wouldn't help, I took my life in my hands and crossed over to fight the Ammonites, and the LORD gave me the victory over them. Now why have you come up today to fight me?"
JUDG|12|4|Jephthah then called together the men of Gilead and fought against Ephraim. The Gileadites struck them down because the Ephraimites had said, "You Gileadites are renegades from Ephraim and Manasseh."
JUDG|12|5|The Gileadites captured the fords of the Jordan leading to Ephraim, and whenever a survivor of Ephraim said, "Let me cross over," the men of Gilead asked him, "Are you an Ephraimite?" If he replied, "No,"
JUDG|12|6|they said, "All right, say 'Shibboleth.'" If he said, "Sibboleth," because he could not pronounce the word correctly, they seized him and killed him at the fords of the Jordan. Forty-two thousand Ephraimites were killed at that time.
JUDG|12|7|Jephthah led Israel six years. Then Jephthah the Gileadite died, and was buried in a town in Gilead.
JUDG|12|8|After him, Ibzan of Bethlehem led Israel.
JUDG|12|9|He had thirty sons and thirty daughters. He gave his daughters away in marriage to those outside his clan, and for his sons he brought in thirty young women as wives from outside his clan. Ibzan led Israel seven years.
JUDG|12|10|Then Ibzan died, and was buried in Bethlehem.
JUDG|12|11|After him, Elon the Zebulunite led Israel ten years.
JUDG|12|12|Then Elon died, and was buried in Aijalon in the land of Zebulun.
JUDG|12|13|After him, Abdon son of Hillel, from Pirathon, led Israel.
JUDG|12|14|He had forty sons and thirty grandsons, who rode on seventy donkeys. He led Israel eight years.
JUDG|12|15|Then Abdon son of Hillel died, and was buried at Pirathon in Ephraim, in the hill country of the Amalekites.
JUDG|13|1|Again the Israelites did evil in the eyes of the LORD, so the LORD delivered them into the hands of the Philistines for forty years.
JUDG|13|2|A certain man of Zorah, named Manoah, from the clan of the Danites, had a wife who was sterile and remained childless.
JUDG|13|3|The angel of the LORD appeared to her and said, "You are sterile and childless, but you are going to conceive and have a son.
JUDG|13|4|Now see to it that you drink no wine or other fermented drink and that you do not eat anything unclean,
JUDG|13|5|because you will conceive and give birth to a son. No razor may be used on his head, because the boy is to be a Nazirite, set apart to God from birth, and he will begin the deliverance of Israel from the hands of the Philistines."
JUDG|13|6|Then the woman went to her husband and told him, "A man of God came to me. He looked like an angel of God, very awesome. I didn't ask him where he came from, and he didn't tell me his name.
JUDG|13|7|But he said to me, 'You will conceive and give birth to a son. Now then, drink no wine or other fermented drink and do not eat anything unclean, because the boy will be a Nazirite of God from birth until the day of his death.'"
JUDG|13|8|Then Manoah prayed to the LORD: "O LORD, I beg you, let the man of God you sent to us come again to teach us how to bring up the boy who is to be born."
JUDG|13|9|God heard Manoah, and the angel of God came again to the woman while she was out in the field; but her husband Manoah was not with her.
JUDG|13|10|The woman hurried to tell her husband, "He's here! The man who appeared to me the other day!"
JUDG|13|11|Manoah got up and followed his wife. When he came to the man, he said, "Are you the one who talked to my wife?I am," he said.
JUDG|13|12|So Manoah asked him, "When your words are fulfilled, what is to be the rule for the boy's life and work?"
JUDG|13|13|The angel of the LORD answered, "Your wife must do all that I have told her.
JUDG|13|14|She must not eat anything that comes from the grapevine, nor drink any wine or other fermented drink nor eat anything unclean. She must do everything I have commanded her."
JUDG|13|15|Manoah said to the angel of the LORD, "We would like you to stay until we prepare a young goat for you."
JUDG|13|16|The angel of the LORD replied, "Even though you detain me, I will not eat any of your food. But if you prepare a burnt offering, offer it to the LORD." (Manoah did not realize that it was the angel of the LORD.)
JUDG|13|17|Then Manoah inquired of the angel of the LORD, "What is your name, so that we may honor you when your word comes true?"
JUDG|13|18|He replied, "Why do you ask my name? It is beyond understanding. "
JUDG|13|19|Then Manoah took a young goat, together with the grain offering, and sacrificed it on a rock to the LORD. And the LORD did an amazing thing while Manoah and his wife watched:
JUDG|13|20|As the flame blazed up from the altar toward heaven, the angel of the LORD ascended in the flame. Seeing this, Manoah and his wife fell with their faces to the ground.
JUDG|13|21|When the angel of the LORD did not show himself again to Manoah and his wife, Manoah realized that it was the angel of the LORD.
JUDG|13|22|"We are doomed to die!" he said to his wife. "We have seen God!"
JUDG|13|23|But his wife answered, "If the LORD had meant to kill us, he would not have accepted a burnt offering and grain offering from our hands, nor shown us all these things or now told us this."
JUDG|13|24|The woman gave birth to a boy and named him Samson. He grew and the LORD blessed him,
JUDG|13|25|and the Spirit of the LORD began to stir him while he was in Mahaneh Dan, between Zorah and Eshtaol.
JUDG|14|1|Samson went down to Timnah and saw there a young Philistine woman.
JUDG|14|2|When he returned, he said to his father and mother, "I have seen a Philistine woman in Timnah; now get her for me as my wife."
JUDG|14|3|His father and mother replied, "Isn't there an acceptable woman among your relatives or among all our people? Must you go to the uncircumcised Philistines to get a wife?" But Samson said to his father, "Get her for me. She's the right one for me."
JUDG|14|4|(His parents did not know that this was from the LORD, who was seeking an occasion to confront the Philistines; for at that time they were ruling over Israel.)
JUDG|14|5|Samson went down to Timnah together with his father and mother. As they approached the vineyards of Timnah, suddenly a young lion came roaring toward him.
JUDG|14|6|The Spirit of the LORD came upon him in power so that he tore the lion apart with his bare hands as he might have torn a young goat. But he told neither his father nor his mother what he had done.
JUDG|14|7|Then he went down and talked with the woman, and he liked her.
JUDG|14|8|Some time later, when he went back to marry her, he turned aside to look at the lion's carcass. In it was a swarm of bees and some honey,
JUDG|14|9|which he scooped out with his hands and ate as he went along. When he rejoined his parents, he gave them some, and they too ate it. But he did not tell them that he had taken the honey from the lion's carcass.
JUDG|14|10|Now his father went down to see the woman. And Samson made a feast there, as was customary for bridegrooms.
JUDG|14|11|When he appeared, he was given thirty companions.
JUDG|14|12|"Let me tell you a riddle," Samson said to them. "If you can give me the answer within the seven days of the feast, I will give you thirty linen garments and thirty sets of clothes.
JUDG|14|13|If you can't tell me the answer, you must give me thirty linen garments and thirty sets of clothes.Tell us your riddle," they said. "Let's hear it."
JUDG|14|14|He replied, "Out of the eater, something to eat; out of the strong, something sweet." For three days they could not give the answer.
JUDG|14|15|On the fourth day, they said to Samson's wife, "Coax your husband into explaining the riddle for us, or we will burn you and your father's household to death. Did you invite us here to rob us?"
JUDG|14|16|Then Samson's wife threw herself on him, sobbing, "You hate me! You don't really love me. You've given my people a riddle, but you haven't told me the answer.I haven't even explained it to my father or mother," he replied, "so why should I explain it to you?"
JUDG|14|17|She cried the whole seven days of the feast. So on the seventh day he finally told her, because she continued to press him. She in turn explained the riddle to her people.
JUDG|14|18|Before sunset on the seventh day the men of the town said to him, "What is sweeter than honey? What is stronger than a lion?" Samson said to them, "If you had not plowed with my heifer, you would not have solved my riddle."
JUDG|14|19|Then the Spirit of the LORD came upon him in power. He went down to Ashkelon, struck down thirty of their men, stripped them of their belongings and gave their clothes to those who had explained the riddle. Burning with anger, he went up to his father's house.
JUDG|14|20|And Samson's wife was given to the friend who had attended him at his wedding.
JUDG|15|1|Later on, at the time of wheat harvest, Samson took a young goat and went to visit his wife. He said, "I'm going to my wife's room." But her father would not let him go in.
JUDG|15|2|"I was so sure you thoroughly hated her," he said, "that I gave her to your friend. Isn't her younger sister more attractive? Take her instead."
JUDG|15|3|Samson said to them, "This time I have a right to get even with the Philistines; I will really harm them."
JUDG|15|4|So he went out and caught three hundred foxes and tied them tail to tail in pairs. He then fastened a torch to every pair of tails,
JUDG|15|5|lit the torches and let the foxes loose in the standing grain of the Philistines. He burned up the shocks and standing grain, together with the vineyards and olive groves.
JUDG|15|6|When the Philistines asked, "Who did this?" they were told, "Samson, the Timnite's son-in-law, because his wife was given to his friend." So the Philistines went up and burned her and her father to death.
JUDG|15|7|Samson said to them, "Since you've acted like this, I won't stop until I get my revenge on you."
JUDG|15|8|He attacked them viciously and slaughtered many of them. Then he went down and stayed in a cave in the rock of Etam.
JUDG|15|9|The Philistines went up and camped in Judah, spreading out near Lehi.
JUDG|15|10|The men of Judah asked, "Why have you come to fight us?We have come to take Samson prisoner," they answered, "to do to him as he did to us."
JUDG|15|11|Then three thousand men from Judah went down to the cave in the rock of Etam and said to Samson, "Don't you realize that the Philistines are rulers over us? What have you done to us?" He answered, "I merely did to them what they did to me."
JUDG|15|12|They said to him, "We've come to tie you up and hand you over to the Philistines." Samson said, "Swear to me that you won't kill me yourselves."
JUDG|15|13|"Agreed," they answered. "We will only tie you up and hand you over to them. We will not kill you." So they bound him with two new ropes and led him up from the rock.
JUDG|15|14|As he approached Lehi, the Philistines came toward him shouting. The Spirit of the LORD came upon him in power. The ropes on his arms became like charred flax, and the bindings dropped from his hands.
JUDG|15|15|Finding a fresh jawbone of a donkey, he grabbed it and struck down a thousand men.
JUDG|15|16|Then Samson said, "With a donkey's jawbone I have made donkeys of them. With a donkey's jawbone I have killed a thousand men."
JUDG|15|17|When he finished speaking, he threw away the jawbone; and the place was called Ramath Lehi.
JUDG|15|18|Because he was very thirsty, he cried out to the LORD, "You have given your servant this great victory. Must I now die of thirst and fall into the hands of the uncircumcised?"
JUDG|15|19|Then God opened up the hollow place in Lehi, and water came out of it. When Samson drank, his strength returned and he revived. So the spring was called En Hakkore, and it is still there in Lehi.
JUDG|15|20|Samson led Israel for twenty years in the days of the Philistines.
JUDG|16|1|One day Samson went to Gaza, where he saw a prostitute. He went in to spend the night with her.
JUDG|16|2|The people of Gaza were told, "Samson is here!" So they surrounded the place and lay in wait for him all night at the city gate. They made no move during the night, saying, "At dawn we'll kill him."
JUDG|16|3|But Samson lay there only until the middle of the night. Then he got up and took hold of the doors of the city gate, together with the two posts, and tore them loose, bar and all. He lifted them to his shoulders and carried them to the top of the hill that faces Hebron.
JUDG|16|4|Some time later, he fell in love with a woman in the Valley of Sorek whose name was Delilah.
JUDG|16|5|The rulers of the Philistines went to her and said, "See if you can lure him into showing you the secret of his great strength and how we can overpower him so we may tie him up and subdue him. Each one of us will give you eleven hundred shekels of silver."
JUDG|16|6|So Delilah said to Samson, "Tell me the secret of your great strength and how you can be tied up and subdued."
JUDG|16|7|Samson answered her, "If anyone ties me with seven fresh thongs that have not been dried, I'll become as weak as any other man."
JUDG|16|8|Then the rulers of the Philistines brought her seven fresh thongs that had not been dried, and she tied him with them.
JUDG|16|9|With men hidden in the room, she called to him, "Samson, the Philistines are upon you!" But he snapped the thongs as easily as a piece of string snaps when it comes close to a flame. So the secret of his strength was not discovered.
JUDG|16|10|Then Delilah said to Samson, "You have made a fool of me; you lied to me. Come now, tell me how you can be tied."
JUDG|16|11|He said, "If anyone ties me securely with new ropes that have never been used, I'll become as weak as any other man."
JUDG|16|12|So Delilah took new ropes and tied him with them. Then, with men hidden in the room, she called to him, "Samson, the Philistines are upon you!" But he snapped the ropes off his arms as if they were threads.
JUDG|16|13|Delilah then said to Samson, "Until now, you have been making a fool of me and lying to me. Tell me how you can be tied." He replied, "If you weave the seven braids of my head into the fabric on the loom and tighten it with the pin, I'll become as weak as any other man." So while he was sleeping, Delilah took the seven braids of his head, wove them into the fabric
JUDG|16|14|and tightened it with the pin. Again she called to him, "Samson, the Philistines are upon you!" He awoke from his sleep and pulled up the pin and the loom, with the fabric.
JUDG|16|15|Then she said to him, "How can you say, 'I love you,' when you won't confide in me? This is the third time you have made a fool of me and haven't told me the secret of your great strength."
JUDG|16|16|With such nagging she prodded him day after day until he was tired to death.
JUDG|16|17|So he told her everything. "No razor has ever been used on my head," he said, "because I have been a Nazirite set apart to God since birth. If my head were shaved, my strength would leave me, and I would become as weak as any other man."
JUDG|16|18|When Delilah saw that he had told her everything, she sent word to the rulers of the Philistines, "Come back once more; he has told me everything." So the rulers of the Philistines returned with the silver in their hands.
JUDG|16|19|Having put him to sleep on her lap, she called a man to shave off the seven braids of his hair, and so began to subdue him. And his strength left him.
JUDG|16|20|Then she called, "Samson, the Philistines are upon you!" He awoke from his sleep and thought, "I'll go out as before and shake myself free." But he did not know that the LORD had left him.
JUDG|16|21|Then the Philistines seized him, gouged out his eyes and took him down to Gaza. Binding him with bronze shackles, they set him to grinding in the prison.
JUDG|16|22|But the hair on his head began to grow again after it had been shaved.
JUDG|16|23|Now the rulers of the Philistines assembled to offer a great sacrifice to Dagon their god and to celebrate, saying, "Our god has delivered Samson, our enemy, into our hands."
JUDG|16|24|When the people saw him, they praised their god, saying, "Our god has delivered our enemy into our hands, the one who laid waste our land and multiplied our slain."
JUDG|16|25|While they were in high spirits, they shouted, "Bring out Samson to entertain us." So they called Samson out of the prison, and he performed for them. When they stood him among the pillars,
JUDG|16|26|Samson said to the servant who held his hand, "Put me where I can feel the pillars that support the temple, so that I may lean against them."
JUDG|16|27|Now the temple was crowded with men and women; all the rulers of the Philistines were there, and on the roof were about three thousand men and women watching Samson perform.
JUDG|16|28|Then Samson prayed to the LORD, "O Sovereign LORD, remember me. O God, please strengthen me just once more, and let me with one blow get revenge on the Philistines for my two eyes."
JUDG|16|29|Then Samson reached toward the two central pillars on which the temple stood. Bracing himself against them, his right hand on the one and his left hand on the other,
JUDG|16|30|Samson said, "Let me die with the Philistines!" Then he pushed with all his might, and down came the temple on the rulers and all the people in it. Thus he killed many more when he died than while he lived.
JUDG|16|31|Then his brothers and his father's whole family went down to get him. They brought him back and buried him between Zorah and Eshtaol in the tomb of Manoah his father. He had led Israel twenty years.
JUDG|17|1|Now a man named Micah from the hill country of Ephraim
JUDG|17|2|said to his mother, "The eleven hundred shekels of silver that were taken from you and about which I heard you utter a curse-I have that silver with me; I took it." Then his mother said, "The LORD bless you, my son!"
JUDG|17|3|When he returned the eleven hundred shekels of silver to his mother, she said, "I solemnly consecrate my silver to the LORD for my son to make a carved image and a cast idol. I will give it back to you."
JUDG|17|4|So he returned the silver to his mother, and she took two hundred shekels of silver and gave them to a silversmith, who made them into the image and the idol. And they were put in Micah's house.
JUDG|17|5|Now this man Micah had a shrine, and he made an ephod and some idols and installed one of his sons as his priest.
JUDG|17|6|In those days Israel had no king; everyone did as he saw fit.
JUDG|17|7|A young Levite from Bethlehem in Judah, who had been living within the clan of Judah,
JUDG|17|8|left that town in search of some other place to stay. On his way he came to Micah's house in the hill country of Ephraim.
JUDG|17|9|Micah asked him, "Where are you from?I'm a Levite from Bethlehem in Judah," he said, "and I'm looking for a place to stay."
JUDG|17|10|Then Micah said to him, "Live with me and be my father and priest, and I'll give you ten shekels of silver a year, your clothes and your food."
JUDG|17|11|So the Levite agreed to live with him, and the young man was to him like one of his sons.
JUDG|17|12|Then Micah installed the Levite, and the young man became his priest and lived in his house.
JUDG|17|13|And Micah said, "Now I know that the LORD will be good to me, since this Levite has become my priest."
JUDG|18|1|In those days Israel had no king. And in those days the tribe of the Danites was seeking a place of their own where they might settle, because they had not yet come into an inheritance among the tribes of Israel.
JUDG|18|2|So the Danites sent five warriors from Zorah and Eshtaol to spy out the land and explore it. These men represented all their clans. They told them, "Go, explore the land." The men entered the hill country of Ephraim and came to the house of Micah, where they spent the night.
JUDG|18|3|When they were near Micah's house, they recognized the voice of the young Levite; so they turned in there and asked him, "Who brought you here? What are you doing in this place? Why are you here?"
JUDG|18|4|He told them what Micah had done for him, and said, "He has hired me and I am his priest."
JUDG|18|5|Then they said to him, "Please inquire of God to learn whether our journey will be successful."
JUDG|18|6|The priest answered them, "Go in peace. Your journey has the LORD 's approval."
JUDG|18|7|So the five men left and came to Laish, where they saw that the people were living in safety, like the Sidonians, unsuspecting and secure. And since their land lacked nothing, they were prosperous. Also, they lived a long way from the Sidonians and had no relationship with anyone else.
JUDG|18|8|When they returned to Zorah and Eshtaol, their brothers asked them, "How did you find things?"
JUDG|18|9|They answered, "Come on, let's attack them! We have seen that the land is very good. Aren't you going to do something? Don't hesitate to go there and take it over.
JUDG|18|10|When you get there, you will find an unsuspecting people and a spacious land that God has put into your hands, a land that lacks nothing whatever."
JUDG|18|11|Then six hundred men from the clan of the Danites, armed for battle, set out from Zorah and Eshtaol.
JUDG|18|12|On their way they set up camp near Kiriath Jearim in Judah. This is why the place west of Kiriath Jearim is called Mahaneh Dan to this day.
JUDG|18|13|From there they went on to the hill country of Ephraim and came to Micah's house.
JUDG|18|14|Then the five men who had spied out the land of Laish said to their brothers, "Do you know that one of these houses has an ephod, other household gods, a carved image and a cast idol? Now you know what to do."
JUDG|18|15|So they turned in there and went to the house of the young Levite at Micah's place and greeted him.
JUDG|18|16|The six hundred Danites, armed for battle, stood at the entrance to the gate.
JUDG|18|17|The five men who had spied out the land went inside and took the carved image, the ephod, the other household gods and the cast idol while the priest and the six hundred armed men stood at the entrance to the gate.
JUDG|18|18|When these men went into Micah's house and took the carved image, the ephod, the other household gods and the cast idol, the priest said to them, "What are you doing?"
JUDG|18|19|They answered him, "Be quiet! Don't say a word. Come with us, and be our father and priest. Isn't it better that you serve a tribe and clan in Israel as priest rather than just one man's household?"
JUDG|18|20|Then the priest was glad. He took the ephod, the other household gods and the carved image and went along with the people.
JUDG|18|21|Putting their little children, their livestock and their possessions in front of them, they turned away and left.
JUDG|18|22|When they had gone some distance from Micah's house, the men who lived near Micah were called together and overtook the Danites.
JUDG|18|23|As they shouted after them, the Danites turned and said to Micah, "What's the matter with you that you called out your men to fight?"
JUDG|18|24|He replied, "You took the gods I made, and my priest, and went away. What else do I have? How can you ask, 'What's the matter with you?'"
JUDG|18|25|The Danites answered, "Don't argue with us, or some hot-tempered men will attack you, and you and your family will lose your lives."
JUDG|18|26|So the Danites went their way, and Micah, seeing that they were too strong for him, turned around and went back home.
JUDG|18|27|Then they took what Micah had made, and his priest, and went on to Laish, against a peaceful and unsuspecting people. They attacked them with the sword and burned down their city.
JUDG|18|28|There was no one to rescue them because they lived a long way from Sidon and had no relationship with anyone else. The city was in a valley near Beth Rehob. The Danites rebuilt the city and settled there.
JUDG|18|29|They named it Dan after their forefather Dan, who was born to Israel-though the city used to be called Laish.
JUDG|18|30|There the Danites set up for themselves the idols, and Jonathan son of Gershom, the son of Moses, and his sons were priests for the tribe of Dan until the time of the captivity of the land.
JUDG|18|31|They continued to use the idols Micah had made, all the time the house of God was in Shiloh.
JUDG|19|1|In those days Israel had no king. Now a Levite who lived in a remote area in the hill country of Ephraim took a concubine from Bethlehem in Judah.
JUDG|19|2|But she was unfaithful to him. She left him and went back to her father's house in Bethlehem, Judah. After she had been there four months,
JUDG|19|3|her husband went to her to persuade her to return. He had with him his servant and two donkeys. She took him into her father's house, and when her father saw him, he gladly welcomed him.
JUDG|19|4|His father-in-law, the girl's father, prevailed upon him to stay; so he remained with him three days, eating and drinking, and sleeping there.
JUDG|19|5|On the fourth day they got up early and he prepared to leave, but the girl's father said to his son-in-law, "Refresh yourself with something to eat; then you can go."
JUDG|19|6|So the two of them sat down to eat and drink together. Afterward the girl's father said, "Please stay tonight and enjoy yourself."
JUDG|19|7|And when the man got up to go, his father-in-law persuaded him, so he stayed there that night.
JUDG|19|8|On the morning of the fifth day, when he rose to go, the girl's father said, "Refresh yourself. Wait till afternoon!" So the two of them ate together.
JUDG|19|9|Then when the man, with his concubine and his servant, got up to leave, his father-in-law, the girl's father, said, "Now look, it's almost evening. Spend the night here; the day is nearly over. Stay and enjoy yourself. Early tomorrow morning you can get up and be on your way home."
JUDG|19|10|But, unwilling to stay another night, the man left and went toward Jebus (that is, Jerusalem), with his two saddled donkeys and his concubine.
JUDG|19|11|When they were near Jebus and the day was almost gone, the servant said to his master, "Come, let's stop at this city of the Jebusites and spend the night."
JUDG|19|12|His master replied, "No. We won't go into an alien city, whose people are not Israelites. We will go on to Gibeah."
JUDG|19|13|He added, "Come, let's try to reach Gibeah or Ramah and spend the night in one of those places."
JUDG|19|14|So they went on, and the sun set as they neared Gibeah in Benjamin.
JUDG|19|15|There they stopped to spend the night. They went and sat in the city square, but no one took them into his home for the night.
JUDG|19|16|That evening an old man from the hill country of Ephraim, who was living in Gibeah (the men of the place were Benjamites), came in from his work in the fields.
JUDG|19|17|When he looked and saw the traveler in the city square, the old man asked, "Where are you going? Where did you come from?"
JUDG|19|18|He answered, "We are on our way from Bethlehem in Judah to a remote area in the hill country of Ephraim where I live. I have been to Bethlehem in Judah and now I am going to the house of the LORD. No one has taken me into his house.
JUDG|19|19|We have both straw and fodder for our donkeys and bread and wine for ourselves your servants-me, your maidservant, and the young man with us. We don't need anything."
JUDG|19|20|"You are welcome at my house," the old man said. "Let me supply whatever you need. Only don't spend the night in the square."
JUDG|19|21|So he took him into his house and fed his donkeys. After they had washed their feet, they had something to eat and drink.
JUDG|19|22|While they were enjoying themselves, some of the wicked men of the city surrounded the house. Pounding on the door, they shouted to the old man who owned the house, "Bring out the man who came to your house so we can have sex with him."
JUDG|19|23|The owner of the house went outside and said to them, "No, my friends, don't be so vile. Since this man is my guest, don't do this disgraceful thing.
JUDG|19|24|Look, here is my virgin daughter, and his concubine. I will bring them out to you now, and you can use them and do to them whatever you wish. But to this man, don't do such a disgraceful thing."
JUDG|19|25|But the men would not listen to him. So the man took his concubine and sent her outside to them, and they raped her and abused her throughout the night, and at dawn they let her go.
JUDG|19|26|At daybreak the woman went back to the house where her master was staying, fell down at the door and lay there until daylight.
JUDG|19|27|When her master got up in the morning and opened the door of the house and stepped out to continue on his way, there lay his concubine, fallen in the doorway of the house, with her hands on the threshold.
JUDG|19|28|He said to her, "Get up; let's go." But there was no answer. Then the man put her on his donkey and set out for home.
JUDG|19|29|When he reached home, he took a knife and cut up his concubine, limb by limb, into twelve parts and sent them into all the areas of Israel.
JUDG|19|30|Everyone who saw it said, "Such a thing has never been seen or done, not since the day the Israelites came up out of Egypt. Think about it! Consider it! Tell us what to do!"
JUDG|20|1|Then all the Israelites from Dan to Beersheba and from the land of Gilead came out as one man and assembled before the LORD in Mizpah.
JUDG|20|2|The leaders of all the people of the tribes of Israel took their places in the assembly of the people of God, four hundred thousand soldiers armed with swords.
JUDG|20|3|(The Benjamites heard that the Israelites had gone up to Mizpah.) Then the Israelites said, "Tell us how this awful thing happened."
JUDG|20|4|So the Levite, the husband of the murdered woman, said, "I and my concubine came to Gibeah in Benjamin to spend the night.
JUDG|20|5|During the night the men of Gibeah came after me and surrounded the house, intending to kill me. They raped my concubine, and she died.
JUDG|20|6|I took my concubine, cut her into pieces and sent one piece to each region of Israel's inheritance, because they committed this lewd and disgraceful act in Israel.
JUDG|20|7|Now, all you Israelites, speak up and give your verdict."
JUDG|20|8|All the people rose as one man, saying, "None of us will go home. No, not one of us will return to his house.
JUDG|20|9|But now this is what we'll do to Gibeah: We'll go up against it as the lot directs.
JUDG|20|10|We'll take ten men out of every hundred from all the tribes of Israel, and a hundred from a thousand, and a thousand from ten thousand, to get provisions for the army. Then, when the army arrives at Gibeah in Benjamin, it can give them what they deserve for all this vileness done in Israel."
JUDG|20|11|So all the men of Israel got together and united as one man against the city.
JUDG|20|12|The tribes of Israel sent men throughout the tribe of Benjamin, saying, "What about this awful crime that was committed among you?
JUDG|20|13|Now surrender those wicked men of Gibeah so that we may put them to death and purge the evil from Israel." But the Benjamites would not listen to their fellow Israelites.
JUDG|20|14|From their towns they came together at Gibeah to fight against the Israelites.
JUDG|20|15|At once the Benjamites mobilized twenty-six thousand swordsmen from their towns, in addition to seven hundred chosen men from those living in Gibeah.
JUDG|20|16|Among all these soldiers there were seven hundred chosen men who were left-handed, each of whom could sling a stone at a hair and not miss.
JUDG|20|17|Israel, apart from Benjamin, mustered four hundred thousand swordsmen, all of them fighting men.
JUDG|20|18|The Israelites went up to Bethel and inquired of God. They said, "Who of us shall go first to fight against the Benjamites?" The LORD replied, "Judah shall go first."
JUDG|20|19|The next morning the Israelites got up and pitched camp near Gibeah.
JUDG|20|20|The men of Israel went out to fight the Benjamites and took up battle positions against them at Gibeah.
JUDG|20|21|The Benjamites came out of Gibeah and cut down twenty-two thousand Israelites on the battlefield that day.
JUDG|20|22|But the men of Israel encouraged one another and again took up their positions where they had stationed themselves the first day.
JUDG|20|23|The Israelites went up and wept before the LORD until evening, and they inquired of the LORD. They said, "Shall we go up again to battle against the Benjamites, our brothers?" The LORD answered, "Go up against them."
JUDG|20|24|Then the Israelites drew near to Benjamin the second day.
JUDG|20|25|This time, when the Benjamites came out from Gibeah to oppose them, they cut down another eighteen thousand Israelites, all of them armed with swords.
JUDG|20|26|Then the Israelites, all the people, went up to Bethel, and there they sat weeping before the LORD. They fasted that day until evening and presented burnt offerings and fellowship offerings to the LORD.
JUDG|20|27|And the Israelites inquired of the LORD. (In those days the ark of the covenant of God was there,
JUDG|20|28|with Phinehas son of Eleazar, the son of Aaron, ministering before it.) They asked, "Shall we go up again to battle with Benjamin our brother, or not?" The LORD responded, "Go, for tomorrow I will give them into your hands."
JUDG|20|29|Then Israel set an ambush around Gibeah.
JUDG|20|30|They went up against the Benjamites on the third day and took up positions against Gibeah as they had done before.
JUDG|20|31|The Benjamites came out to meet them and were drawn away from the city. They began to inflict casualties on the Israelites as before, so that about thirty men fell in the open field and on the roads-the one leading to Bethel and the other to Gibeah.
JUDG|20|32|While the Benjamites were saying, "We are defeating them as before," the Israelites were saying, "Let's retreat and draw them away from the city to the roads."
JUDG|20|33|All the men of Israel moved from their places and took up positions at Baal Tamar, and the Israelite ambush charged out of its place on the west of Gibeah.
JUDG|20|34|Then ten thousand of Israel's finest men made a frontal attack on Gibeah. The fighting was so heavy that the Benjamites did not realize how near disaster was.
JUDG|20|35|The LORD defeated Benjamin before Israel, and on that day the Israelites struck down 25,100 Benjamites, all armed with swords.
JUDG|20|36|Then the Benjamites saw that they were beaten. Now the men of Israel had given way before Benjamin, because they relied on the ambush they had set near Gibeah.
JUDG|20|37|The men who had been in ambush made a sudden dash into Gibeah, spread out and put the whole city to the sword.
JUDG|20|38|The men of Israel had arranged with the ambush that they should send up a great cloud of smoke from the city,
JUDG|20|39|and then the men of Israel would turn in the battle. The Benjamites had begun to inflict casualties on the men of Israel (about thirty), and they said, "We are defeating them as in the first battle."
JUDG|20|40|But when the column of smoke began to rise from the city, the Benjamites turned and saw the smoke of the whole city going up into the sky.
JUDG|20|41|Then the men of Israel turned on them, and the men of Benjamin were terrified, because they realized that disaster had come upon them.
JUDG|20|42|So they fled before the Israelites in the direction of the desert, but they could not escape the battle. And the men of Israel who came out of the towns cut them down there.
JUDG|20|43|They surrounded the Benjamites, chased them and easily overran them in the vicinity of Gibeah on the east.
JUDG|20|44|Eighteen thousand Benjamites fell, all of them valiant fighters.
JUDG|20|45|As they turned and fled toward the desert to the rock of Rimmon, the Israelites cut down five thousand men along the roads. They kept pressing after the Benjamites as far as Gidom and struck down two thousand more.
JUDG|20|46|On that day twenty-five thousand Benjamite swordsmen fell, all of them valiant fighters.
JUDG|20|47|But six hundred men turned and fled into the desert to the rock of Rimmon, where they stayed four months.
JUDG|20|48|The men of Israel went back to Benjamin and put all the towns to the sword, including the animals and everything else they found. All the towns they came across they set on fire.
JUDG|21|1|The men of Israel had taken an oath at Mizpah: "Not one of us will give his daughter in marriage to a Benjamite."
JUDG|21|2|The people went to Bethel, where they sat before God until evening, raising their voices and weeping bitterly.
JUDG|21|3|"O LORD, the God of Israel," they cried, "why has this happened to Israel? Why should one tribe be missing from Israel today?"
JUDG|21|4|Early the next day the people built an altar and presented burnt offerings and fellowship offerings.
JUDG|21|5|Then the Israelites asked, "Who from all the tribes of Israel has failed to assemble before the LORD?" For they had taken a solemn oath that anyone who failed to assemble before the LORD at Mizpah should certainly be put to death.
JUDG|21|6|Now the Israelites grieved for their brothers, the Benjamites. "Today one tribe is cut off from Israel," they said.
JUDG|21|7|"How can we provide wives for those who are left, since we have taken an oath by the LORD not to give them any of our daughters in marriage?"
JUDG|21|8|Then they asked, "Which one of the tribes of Israel failed to assemble before the LORD at Mizpah?" They discovered that no one from Jabesh Gilead had come to the camp for the assembly.
JUDG|21|9|For when they counted the people, they found that none of the people of Jabesh Gilead were there.
JUDG|21|10|So the assembly sent twelve thousand fighting men with instructions to go to Jabesh Gilead and put to the sword those living there, including the women and children.
JUDG|21|11|"This is what you are to do," they said. "Kill every male and every woman who is not a virgin."
JUDG|21|12|They found among the people living in Jabesh Gilead four hundred young women who had never slept with a man, and they took them to the camp at Shiloh in Canaan.
JUDG|21|13|Then the whole assembly sent an offer of peace to the Benjamites at the rock of Rimmon.
JUDG|21|14|So the Benjamites returned at that time and were given the women of Jabesh Gilead who had been spared. But there were not enough for all of them.
JUDG|21|15|The people grieved for Benjamin, because the LORD had made a gap in the tribes of Israel.
JUDG|21|16|And the elders of the assembly said, "With the women of Benjamin destroyed, how shall we provide wives for the men who are left?
JUDG|21|17|The Benjamite survivors must have heirs," they said, "so that a tribe of Israel will not be wiped out.
JUDG|21|18|We can't give them our daughters as wives, since we Israelites have taken this oath: 'Cursed be anyone who gives a wife to a Benjamite.'
JUDG|21|19|But look, there is the annual festival of the LORD in Shiloh, to the north of Bethel, and east of the road that goes from Bethel to Shechem, and to the south of Lebonah."
JUDG|21|20|So they instructed the Benjamites, saying, "Go and hide in the vineyards
JUDG|21|21|and watch. When the girls of Shiloh come out to join in the dancing, then rush from the vineyards and each of you seize a wife from the girls of Shiloh and go to the land of Benjamin.
JUDG|21|22|When their fathers or brothers complain to us, we will say to them, 'Do us a kindness by helping them, because we did not get wives for them during the war, and you are innocent, since you did not give your daughters to them.'"
JUDG|21|23|So that is what the Benjamites did. While the girls were dancing, each man caught one and carried her off to be his wife. Then they returned to their inheritance and rebuilt the towns and settled in them.
JUDG|21|24|At that time the Israelites left that place and went home to their tribes and clans, each to his own inheritance.
JUDG|21|25|In those days Israel had no king; everyone did as he saw fit.
