PS|1|1|Блажен муж, що за радою несправедливих не ходить, і не стоїть на дорозі грішних, і не сидить на сидінні злоріків,
PS|1|2|та в Законі Господнім його насолода, і про Закон Його вдень та вночі він роздумує!
PS|1|3|І він буде, як дерево, над водним потоком посаджене, що родить свій плід своєдчасно, і що листя не в'яне його, і все, що він чинить, щаститься йому!
PS|1|4|Не так ті безбожні, вони як полова, що вітер її розвіває!
PS|1|5|Ось тому то не встоять безбожні на суді, ані грішники у зборі праведних,
PS|1|6|дорогу бо праведних знає Господь, а дорога безбожних загине!
PS|2|1|Чого то племена бунтують, а народи задумують марне?
PS|2|2|Земні царі повстають, і князі нараджуються разом на Господа та на Його Помазанця:
PS|2|3|Позриваймо ми їхні кайдани, і поскидаймо із себе їхні пута!
PS|2|4|Але Той, Хто на небесах пробуває посміється, Владика їх висміє!
PS|2|5|Він тоді в Своїм гніві промовить до них, і настрашить їх Він у Своїм пересерді:
PS|2|6|Я ж помазав Свого Царя на Сіон, святу гору Свою.
PS|2|7|Я хочу звістити постанову: Промовив до Мене Господь: Ти Мій Син, Я сьогодні Тебе породив.
PS|2|8|Жадай Ти від Мене, і дам Я народи Тобі, як спадщину Твою, володіння ж Твоє аж по кінці землі!
PS|2|9|Ти їх повбиваєш залізним жезлом, потовчеш їх, як посуд ганчарський...
PS|2|10|А тепер помудрійте, царі, навчіться ви, судді землі:
PS|2|11|Служіть Господеві зо страхом, і радійте з тремтінням!
PS|2|12|Шануйте Сина, щоб Він не розгнівався, і щоб вам не загинути в дорозі, бо гнів Його незабаром запалиться. Блаженні усі, хто на Нього надіється!
PS|3|1|Псалом Давидів, як він утікав був від перед Авесаломом, своїм сином. (3-2) Господи, як багато моїх ворогів, як багато стають проти мене!
PS|3|2|(3-3) Багато-хто кажуть про душу мою: Йому в Бозі спасіння нема! Села.
PS|3|3|(3-4) Але, Господи, щит Ти для мене та слава моя, і мою голову Ти підіймаєш!
PS|3|4|(3-5) Своїм голосом кличу до Господа, і Він озветься зо святої Своєї гори. Села.
PS|3|5|(3-6) Я лягаю і сплю, і пробуджуюся, бо Господь підпирає мене,
PS|3|6|(3-7) і я не побоюсь десяти тисяч люду, які проти мене навколо отаборились!
PS|3|7|(3-8) Устань же, о Господи! Спаси мене, Боже мій, бо Ти разиш усіх ворогів моїх в щоку, зуби грішникам крушиш!
PS|3|8|(3-9) Спасіння від Господа, і над народом Твоїм Твоє благословення! Села.
PS|4|1|Для дириґетна хору. На струнніх знаряддях. Псалом Давидів. (4-2) Коли кличу, озвися до мене, Боже правди моєї, Ти простір для мене робив у тісноті... Помилуй мене, і почуй молитву мою!
PS|4|2|(4-3) Людські сини, доки слава моя буде ганьбитись? Доки будете марне любити, шукати неправди? Села.
PS|4|3|(4-4) і знайте, що святого для Себе Господь відділив, почує Господь, як я кликати буду до Нього!
PS|4|4|(4-5) Гнівайтеся, та не грішіть; на ложах своїх розмишляйте у ваших серцях, та й мовчіть! Села.
PS|4|5|(4-6) Жертви правди приносьте, і надійтесь на Господа.
PS|4|6|(4-7) Багато-хто кажуть: Хто нам покаже добро? Підійми ж на нас, Господи, світло Свого лиця!
PS|4|7|(4-8) Ти даєш більшу радість у серці моїм, ніж у них, як помножилося їхнє збіжжя та їхнє вино молоде.
PS|4|8|(4-9) У спокої я ляжу, і засну, бо Ти, Господи, єдиний даєш мені жити безпечно!
PS|5|1|Для дириґетна хору. До флейти. Псалом Давидів. (5-2) Почуй, Господи, мову мою, стогнання моє зрозумій.
PS|5|2|(5-3) Прислухайсь до голосу зойку мого, о мій Царю та Боже Ти мій, як до Тебе молитися буду!
PS|5|3|(5-4) Ти слухаєш, Господи, ранком мій голос, ранком молитися буду до Тебе та буду чекати,
PS|5|4|(5-5) бо Бог Ти не той, що несправедливости хоче, зло не буде в Тобі пробувати!
PS|5|5|(5-6) Перед очима Твоїми не втримаються гультяї, всіх злочинців ненавидиш Ти.
PS|5|6|(5-7) Погубиш Ти неправдомовців, кровожерну й підступну людину обридить Господь.
PS|5|7|(5-8) А я в ласці великій Твоїй до дому Твого ввійду, до Храму святого Твого вклонюся в страху Твоїм.
PS|5|8|(5-9) Провадь мене, Господи, в правді Своїй задля моїх ворогів, і вирівняй передо мною дорогу Свою,
PS|5|9|(5-10) бо в їхніх устах нема правди, нутро їхнє приносить нещастя, гріб відкритий їхнє горло, свій язик вони роблять гладеньким!
PS|5|10|(5-11) Признай їх за винних, о Боже, через свої заміри хай упадуть, за їхні великі злочинства відкинь їх від Себе, бо вони проти Тебе бунтують!
PS|5|11|(5-12) А всі, хто надію на Тебе складають, хай тішаться, будуть вічно співати вони, і Ти їх охорониш, і будуть радіти Тобою, хто любить ім'я Твоє!
PS|5|12|(5-13) Бо Ти, Господи, благословлятимеш праведного, милістю вкриєш його, як щитом!
PS|6|1|Для дириґетна хору. На струнніх знаряддях. На октаву. Псалом Давидів. (6-2) Не карай мене, Господи, в гніві Своїм, не завдавай мені кари в Своїм пересерді!
PS|6|2|(6-3) Помилуй мене, Господи, я ж бо слабий, уздоров мене, Господи, бо тремтять мої кості,
PS|6|3|(6-4) і душа моя сильно стривожена, а ти, Господи, доки?
PS|6|4|(6-5) Вернися, о Господи, визволи душу мою, ради ласки Своєї спаси Ти мене!
PS|6|5|(6-6) Бож у смерті нема пам'ятання про Тебе, у шеолі ж хто буде хвалити Тебе?
PS|6|6|(6-7) Змучився я від стогнання свого, щоночі постелю свою обмиваю слізьми, сльозами своїми окроплюю ложе своє!...
PS|6|7|(6-8) Моє око зів'яло з печалі, постаріло через усіх ворогів моїх...
PS|6|8|(6-9) Відступіться від мене, усі беззаконники, бо почув Господь голос мого плачу!
PS|6|9|(6-10) Благання моє Господь вислухає, молитву мою Господь прийме,
PS|6|10|(6-11) усі мої вороги посоромлені будуть, і будуть настрашені дуже: хай вернуться, і будуть вони посоромлені зараз!
PS|7|1|Жалібна пісня Давидова, яку він співав Господеві в справі веніямінівця Куща.
PS|7|2|(7-3) щоб ворог моєї душі не розшарпав, як лев, що кості ламає, й ніхто не рятує!
PS|7|3|(7-4) Господи, Боже мій, коли я таке учинив, коли є беззаконня в долонях моїх,
PS|7|4|(7-5) коли я доброчинцеві злом відплатив, і без причини ограбував свого противника,
PS|7|5|(7-6) ворог нехай переслідує душу мою, і нехай дожене, і нехай до землі він потопче життя моє, і хай мою славу оберне на порох! Села.
PS|7|6|(7-7) Устань же, о Господи, в гніві Своїм, понесися на лютість моїх ворогів, і до мене скеруй постанову Свою, яку Ти заповів!
PS|7|7|(7-8) і громада народів оточить Тебе, і над нею вернися на висоту!
PS|7|8|(7-9) Господь судить людей, суди ж мене, Господи, за моєю правотою й за моєю невинністю.
PS|7|9|(7-10) Нехай злоба безбожних скінчиться, а Ти зміцни праведного, бо вивідуєш Ти серця й нирки, о праведний Боже!
PS|7|10|(7-11) Щит мій у Бозі, Який чистих серцем спасає.
PS|7|11|(7-12) Бог Суддя справедливий, і щоденно на злого Бог гнівається,
PS|7|12|(7-13) коли хто не навернеться, буде гострити меча Свого Він, Свого лука натягне й наставить його,
PS|7|13|(7-14) і йому приготовив смертельні знаряддя, Він зробить огнистими стріли Свої.
PS|7|14|(7-15) Ото, беззаконня зачне нечестивий, і завагітніє безправ'ям, і породить неправду.
PS|7|15|(7-16) Він рова копав, і його викопав, і впав сам до ями, яку приготовив,
PS|7|16|(7-17) обернеться зло його на його голову, і на маківку зійде його беззаконня!
PS|7|17|(7-18) Я ж Господа буду хвалити за Його правдою, і буду виспівувати Ймення Всевишнього Господа!
PS|8|1|Для дириґетна хору. На інструменті ґатійськім. Псалом Давидів. (8-2) Господи, Владико наш, яке то величне на цілій землі Твоє Ймення, Слава Твоя понад небесами!
PS|8|2|(8-3) З уст дітей й немовлят учинив Ти хвалу ради Своїх ворогів, щоб знищити противника й месника.
PS|8|3|(8-4) Коли бачу Твої небеса діло пальців Твоїх, місяця й зорі, що Ти встановив,
PS|8|4|(8-5) то що є людина, що Ти пам'ятаєш про неї, і син людський, про якого Ти згадуєш?
PS|8|5|(8-6) А однак учинив Ти його мало меншим від Бога, і славою й величчю Ти коронуєш його!
PS|8|6|(8-7) Учинив Ти його володарем творива рук Своїх, все під ноги йому вмістив:
PS|8|7|(8-8) худобу дрібну та биків, їх усіх, а також степових звірів диких,
PS|8|8|(8-9) птаство небесне та риби морські, і все, що морськими дорогами ходить!
PS|8|9|(8-10) Господи, Боже наш, яке то величне на цілій землі Твоє Ймення!
PS|9|1|Для дириґетна хору. На спів: „На смерть сина". Псалом Давидів. (9-2) Хвалитиму Господа усім серцем своїм, розповім про всі чуда Твої!
PS|9|2|(9-3) Я буду радіти, і тішитись буду Тобою, і буду виспівувати Ймення Твоє, о Всевишній!
PS|9|3|(9-4) Як будуть назад відступати мої вороги, то спіткнуться і вигинуть перед обличчям Твоїм!
PS|9|4|(9-5) Бо суд мій і справу мою розсудив Ти, Ти на троні суддевім сидів, Судде праведний!
PS|9|5|(9-6) Докорив Ти народам, безбожного знищив, ім'я їхнє Ти витер на вічні віки!
PS|9|6|(9-7) О вороже мій, руйнування твої закінчились на вічність, ти й міста повалив був, і згинула з ними їхня пам'ять!
PS|9|7|(9-8) Та буде Господь пробувати навіки, Він для суду поставив престола Свого,
PS|9|8|(9-9) і вселенну Він буде судити по правді, справедливістю буде судити народи.
PS|9|9|(9-10) і твердинею буде Господь для пригніченого, в час недолі притулком.
PS|9|10|(9-11) і на Тебе надіятись будуть усі, що ім'я Твоє знають, бо не кинув Ти, Господи, тих, хто шукає Тебе!
PS|9|11|(9-12) Співайте Господеві, що сидить на Сіоні, між народами розповідайте про чини Його,
PS|9|12|(9-13) бо карає Він вчинки криваві, про них пам'ятає, і не забуває Він зойку убогих!
PS|9|13|(9-14) Помилуй мене, Господи, поглянь на страждання моє від моїх ненависників, Ти, що мене підіймаєш із брам смерти,
PS|9|14|(9-15) щоб я розповідав про всю славу Твою, у брамах Сіонської доні я буду радіти спасінням Твоїм!
PS|9|15|(9-16) Народи попадали в яму, яку самі викопали, до пастки, яку заховали, нога їхня схоплена.
PS|9|16|(9-17) Господь знаний, Він суд учинив, спіткнувсь нечестивий у вчинку своєї руки! Гра на струнах. Села.
PS|9|17|(9-18) Попрямують безбожні в шеол, всі народи, що Бога забули,
PS|9|18|(9-19) бож не навіки забудеться бідний, надія убогих не згине назавжди!
PS|9|19|(9-20) Устань же, о Господи, хай людина не перемагає, нехай перед лицем Твоїм засуджені будуть народи!
PS|9|20|(9-21) Накинь, Господи, пострах на них, нехай знають народи, що вони тільки люди! Села.
PS|10|1|Для чого стоїш Ти, о Господи, здалека, в час недолі ховаєшся?
PS|10|2|Безбожний в своїм гордуванні женеться за вбогим, хай схоплені будуть у підступах, які замишляли вони!
PS|10|3|Бо жаданням своєї душі нечестивий пишається, а ласун проклинає, зневажає він Господа.
PS|10|4|У гордощах каже безбожний, що Він не слідкує, бо Бога нема, оце всі його помисли!...
PS|10|5|Сильні дороги його повсякчасно, від нього суди Твої високо, тим то віддмухує він ворогів своїх...
PS|10|6|Сказав він у серці своєму: Я не захитаюсь, бо лиха навіки не буде мені...
PS|10|7|Уста його повні прокляття й обмани та зради, під його язиком злочинство й переступ.
PS|10|8|Причаївшись, сидить на подвір'ях, мордує невинного, його очі слідкують за вбогим...
PS|10|9|В укритті він чатує, як лев той у зарості, чатує схопити убогого, хапає убогого й тягне його в свою сітку...
PS|10|10|Припадає, знижається він, і попадають убогі в його міцні кігті...
PS|10|11|Безбожний говорить у серці своїм: Бог забув, заховав Він обличчя Своє, не побачить ніколи.
PS|10|12|Устань же, о Господи Боже, руку Свою підійми, не забудь про убогих!
PS|10|13|Чому нечестивий ображує Бога і говорить у серці своїм, що Ти не слідкуєш?
PS|10|14|Але Ти все бачиш, бо спостерігаєш злочинство та утиск, щоб віддати Своєю рукою! На Тебе слабий опирається, Ти сироті помічник.
PS|10|15|Зламай же рамено безбожному, і злого скарай за неправду його, аж більше не знайдеш його!
PS|10|16|Господь Цар на вічні віки, із землі Його згинуть погани!
PS|10|17|Бажання понижених чуєш Ти, Господи, серця їх зміцняєш, їх вислуховує ухо Твоє,
PS|10|18|щоб дати суд сироті та пригніченому, щоб більш не страшив чоловік із землі!
PS|11|1|Для дириґетна хору. Давидів. Я надіюсь на Господа, як же кажете ви до моєї душі: Відлітай ти на гору свою, немов птах?
PS|11|2|Бо ось, нечестиві натягують лука, міцно ставлять стрілу свою на тятиву, щоб у темряві до простосердих стріляти...
PS|11|3|Як основи зруйновано, що тоді праведний зробить?
PS|11|4|Господь у святім Своїм храмі, Господь престол Його на небесах, бачать очі Його, повіки Його випробовують людських синів!
PS|11|5|Господь випробовує праведного, а безбожного й того, хто любить насилля, ненавидить душа Його!
PS|11|6|Він спустить дощем на безбожних горюче вугілля, огонь, і сірку, і вітер гарячий, це частка їхньої чаші.
PS|11|7|Бо Господь справедливий, кохає Він правду, праведний бачить обличчя Його!
PS|12|1|Для дириґетна хору. На октаву. Псалом Давидів. (12-2) Спаси мене, Господи, бо нема вже побожного, з-поміж людських синів позникали вже вірні!
PS|12|2|(12-3) Марноту говорять один до одного, їхні уста облесні, і серцем подвійним говорять...
PS|12|3|(12-4) Нехай підітне Господь уста облесливі та язика чванькуватого
PS|12|4|(12-5) тим, хто говорить: Своїм язиком будем сильні, наші уста при нас, хто ж буде нам пан?
PS|12|5|(12-6) Через утиск убогих, ради стогону бідних тепер Я повстану, говорить Господь, поставлю в безпеці того, на кого розтягують сітку!
PS|12|6|(12-7) Господні слова слова чисті, як срібло, очищене в глинянім горні, сім раз перетоплене!
PS|12|7|(12-8) Ти, Господи, їх пильнуватимеш, і будеш навіки нас стерегти перед родом оцим!
PS|12|8|(12-9) Безбожні кружляють навколо, бо нікчемність між людських синів підіймається.
PS|13|1|Для дириґетна хору. Псалом Давидів. (13-2) Доки, Господи, будеш мене забувати назавжди, доки будеш ховати від мене обличчя Своє?
PS|13|2|(13-3) Як довго я буду складати в душі своїй болі, у серці своїм щодня смуток? Як довго мій ворог підноситись буде над мене?
PS|13|3|(13-4) Зглянься, озвися до мене, о Господи, Боже мій! Просвітли мої очі, щоб на смерть не заснув я!
PS|13|4|(13-5) Щоб мій неприятель не сказав: Я його переміг! Щоб мої вороги не раділи, як я захитаюсь!
PS|13|5|(13-6) Я надію на милість Твою покладаю, моє серце радіє спасінням Твоїм!
PS|13|6|(13-7) Я буду співати Господеві, бо Він добродійство для мене вчинив...
PS|14|1|Для дириґетна хору. Давидів. Безумний говорить у серці своїм: Нема Бога! Зіпсулись вони, і обридливий чинять учинок, нема доброчинця!...
PS|14|2|Господь дивиться з неба на людських синів, щоб побачити, чи є там розумний, що Бога шукає.
PS|14|3|Усе повідступало, разом стали бридкими вони, нема доброчинця, нема ні одного!...
PS|14|4|Чи ж не розуміють всі ті, хто чинить безправ'я, хто мій люд поїдає? Вони хліб Господній їдять, та не кличуть Його...
PS|14|5|Тоді настрашилися страхом вони, бо Бог в праведнім роді.
PS|14|6|Раду вбогого ганьбите ви, та Господь охорона йому.
PS|14|7|Аби то Він дав із Сіону спасіння ізраїлеві! Як долю Своєму народу поверне Господь, то радітиме Яків, втішатися буде ізраїль!
PS|15|1|Псалом Давидів. Господи, хто може перебувати в наметі Твоїм? Хто мешкати може на святій Твоїй горі?
PS|15|2|Той, хто в невинності ходить, і праведність чинить, і правду говорить у серці своїм,
PS|15|3|хто не обмовляє своїм язиком, і злого не чинить для друга свого, і свого ближнього не зневажає!
PS|15|4|Обридливий погорджений в очах його, і він богобійних шанує, присягає, для себе хоча б і на зло, і дотримує;
PS|15|5|не дає свого срібла на лихву, і не бере на невинного підкупу. Хто чинить таке, ніколи той не захитається!
PS|16|1|Золота пісня Давадова. Хорони мене, Боже, я бо до Тебе вдаюся!
PS|16|2|Я сказав Господеві: Ти Бог мій, добро моє тільки в Тобі!
PS|16|3|До святих, які на землі, що шляхетні вони, до них все жадання моє!
PS|16|4|Нехай множаться смутки для тих, хто набув собі інших богів, я не буду приносить їм ливної жертви із крови, і їхніх імен не носитиму в устах своїх!
PS|16|5|Господь то частина спадку мого та чаші моєї, Ти долю мою підпираєш!
PS|16|6|Частки припали для мене в хороших місцях, і гарна для мене спадщина моя!
PS|16|7|Благословляю я Господа, що радить мені, навіть ночами навчають мене мої нирки.
PS|16|8|Уявляю я Господа перед собою постійно, бо Він по правиці моїй, й я не буду захитаний!
PS|16|9|Через те моє серце радіє та дух веселиться, і тіло моє спочиває безпечно!
PS|16|10|Бо Ти не опустиш моєї душі до шеолу, не попустиш Своєму святому побачити тління!
PS|16|11|Дорогу життя Ти покажеш мені: радість велика з Тобою, завжди блаженство в правиці Твоїй!
PS|17|1|Молитва Давидова. Вислухай, Господи, правду мою, послухай благання моє! Почуй молитву мою із уст необлудних!
PS|17|2|Від Твого лиця нехай вирок мій вийде, а очі Твої нехай бачать мою правоту!
PS|17|3|Ти випробував моє серце, навістив уночі, перетопив Ти мене, й не знайшов чогось злого. і роздумував я, щоб лихе з моїх уст не виходило,
PS|17|4|а в людських ділах, за словом уст Твоїх, я стерігся доріг гнобителя.
PS|17|5|Зміцняй стопи мої на дорогах Твоїх, щоб кроки мої не хиталися!
PS|17|6|Я кличу до Тебе, бо відповіси мені, Боже, нахили Своє ухо до мене, вислухай мову мою,
PS|17|7|покажи дивну милість Свою, Спасителю тих, хто вдається до Тебе від заколотників проти правиці Твоєї.
PS|17|8|Хорони Ти мене, як зіницю Свою, дочку ока, у тіні Своїх крил заховай Ти мене
PS|17|9|від безбожних, що гублять мене, смертельні мої вороги оточили мене!
PS|17|10|Товщем замкнули вони своє серце, уста їхні говорять бундючно.
PS|17|11|Вороги оточили тепер наші кроки, наставили очі свої, щоб мене повалити на землю...
PS|17|12|із них кожен подібний до лева, що шарпати прагне, й як левчук, що сидить в укритті...
PS|17|13|Устань же, о Господи, його попередь, кинь його на коліна! Мечем Своїм душу мою збережи від безбожного,
PS|17|14|від людей рукою Своєю, Господи, від людей цього світу, що частка їхня в цьому житті, що Ти скарбом Своїм наповняєш їхнє черево! Ситі їхні сини, останок же свій для дітей вони лишать.
PS|17|15|А я в правді побачу обличчя Твоє, і, збудившись, насичусь Твоєю подобою!
PS|18|1|Для дириґента хору. Раба Господнього Давида, коли він промовив до Господа слова цієї пісні того дня, як Господь урятував його з руки всіх його ворогів та від руки Саула, (18-2) то він проказав: Полюблю Тебе, Господи, сило моя,
PS|18|2|(18-3) Господь моя скеля й твердиня моя, і Він мій Спаситель! Мій Бог моя скеля, сховаюсь я в ній, Він щит мій, і ріг Він спасіння мого, Він башта моя!
PS|18|3|(18-4) Я кличу: Преславний Господь, і я визволений від своїх ворогів!
PS|18|4|(18-5) Тенета смертельні мене оточили, і потоки велійяала лякають мене!
PS|18|5|(18-6) Тенета шеолу мене оточили, і пастки смертельні мене попередили.
PS|18|6|(18-7) В тісноті своїй кличу до Господа, і до Бога свого я взиваю, Він почує мій голос із храму Свого, і доходить мій зойк до лиця Його в уші Йому!
PS|18|7|(18-8) Захиталась земля й затремтіла, і затряслись і хитались підвалини гір, бо Він запалився від гніву:
PS|18|8|(18-9) із ніздер Його бухнув дим, з Його ж уст пожирущий огонь, і жар запалився від Нього!
PS|18|9|(18-10) Він небо простяг і спустився, а хмара густа під ногами Його.
PS|18|10|(18-11) Усівся Він на херувима й летів, і на вітрових крилах понісся...
PS|18|11|(18-12) Поклав темряву Він як заслону Свою, довкілля Його то темрява вод, а мешкання Його густі хмари!
PS|18|12|(18-13) Від блиску, що був перед Ним, град і жар огняний пройшли хмари Його...
PS|18|13|(18-14) і Господь загримів у небесах, і Всевишній Свій голос подав, град і жар огняний!
PS|18|14|(18-15) Він послав Свої стріли, та їх розпорошив, і стрілив Він блискавками, та їх побентежив.
PS|18|15|(18-16) Показалися річища водні, і відкрились основи вселенної, від сваріння Твого, о Господи, від подиху вітру із ніздер Твоїх...
PS|18|16|(18-17) Він простяг з висоти Свою руку, узяв Він мене, витяг мене з вод великих,
PS|18|17|(18-18) він мене врятував від мого потужного ворога, і від моїх ненависників, бо сильніші від мене вони!
PS|18|18|(18-19) Напали на мене вони в день нещастя мого, та Господь був моїм опертям,
PS|18|19|(18-20) і на місце розлоге Він вивів мене, Він мене врятував, бо вподобав мене!
PS|18|20|(18-21) Нехай Господь зробить мені за моєю справедливістю, хай заплатить мені згідно з чистістю рук моїх,
PS|18|21|(18-22) бо беріг я дороги Господні, і від Бога свого я не відступив,
PS|18|22|(18-23) бо всі Його присуди передо мною, і не відкидав я від себе Його постанов!
PS|18|23|(18-24) і був я із Ним непорочний, і стерігся своєї провини,
PS|18|24|(18-25) і Господь заплатив був мені за моєю справедливістю, згідно з чистістю рук моїх перед очима Його.
PS|18|25|(18-26) із справедливим поводишся Ти справедливо, із чесним по-чесному,
PS|18|26|(18-27) із чистим поводишся чисто, а з лукавим за лукавством його,
PS|18|27|(18-28) бо народ із біди Ти спасаєш, а очі зухвалі принижуєш,
PS|18|28|(18-29) бо Ти світиш мого світильника, Господь Бог мій, освітлює Він мою темряву!
PS|18|29|(18-30) Бо з Тобою поб'ю я ворожого відділа, і з Богом своїм проберусь через мур.
PS|18|30|(18-31) Бог непорочна дорога Його, слово Господнє очищене, щит Він для всіх, хто вдається до Нього!
PS|18|31|(18-32) Бо хто Бог, окрім Господа? і хто скеля, крім нашого Бога?
PS|18|32|(18-33) Цей Бог мене силою оперезав, і дорогу мою учинив непорочною,
PS|18|33|(18-34) Він зробив мої ноги, мов у лані, і ставить мене на висотах моїх,
PS|18|34|(18-35) мої руки навчає до бою, і на рамена мої лука мідяного напинає.
PS|18|35|(18-36) і дав Ти мені щит спасіння Свого, а правиця Твоя підпирає мене, і чинить великим мене Твоя поміч.
PS|18|36|(18-37) Ти чиниш широким мій крок підо мною, і стопи мої не спіткнуться.
PS|18|37|(18-38) Женуся я за ворогами своїми, і їх дожену, і не вернуся, аж поки не винищу їх,
PS|18|38|(18-39) я їх потрощу, й вони встати не зможуть, повпадають під ноги мої!
PS|18|39|(18-40) Ти ж для бою мене підперізуєш силою, валиш під мене моїх ворохобників.
PS|18|40|(18-41) Повернув Ти до мене плечима моїх ворогів, і понищу ненависників я своїх!
PS|18|41|(18-42) Кричали вони, та немає спасителя, взивали до Господа, і не відповів їм.
PS|18|42|(18-43) і я їх зітру, як той порох на вітрі, як болото на вулицях, їх потопчу!
PS|18|43|(18-44) Ти від бунту народу мене бережеш, Ти робиш мене головою племенам, мені будуть служити народи, яких я не знав!
PS|18|44|(18-45) На вістку про мене слухняні мені, до мене чужинці підлещуються,
PS|18|45|(18-46) в'януть чужинці і тремтять у твердинях своїх...
PS|18|46|(18-47) Живий Господь, і благословенна будь, скеле моя, і нехай Бог спасіння мойого звеличиться,
PS|18|47|(18-48) Бог, що помсти за мене дає, і що народи під мене підбив,
PS|18|48|(18-49) що рятує мене від моїх ворогів, Ти звеличив мене над повстанців на мене, спасаєш мене від насильника!
PS|18|49|(18-50) Тому то хвалю Тебе, Господи, серед народів, і Йменню Твоєму співаю!
PS|18|50|(18-51) Ти Своєму цареві спасіння побільшуєш, і милість вчиняєш Своєму помазанцеві Давиду й насінню його аж навіки.
PS|19|1|Для дириґетна хору. Псалом Давидів. (19-2) Небо звіщає про Божую славу, а про чин Його рук розказує небозвід.
PS|19|2|(19-3) Оповіщує день дневі слово, а ніч ночі показує думку,
PS|19|3|(19-4) без мови й без слів, не чутний їхній голос,
PS|19|4|(19-5) та по цілій землі пішов відголос їхній, і до краю вселенної їхні слова! Для сонця намета поставив у них,
PS|19|5|(19-6) а воно, немов той молодий, що виходить із-під балдахину свого, воно тішиться, мов той герой, щоб пробігти дорогу!
PS|19|6|(19-7) Вихід його з краю неба, а обіг його аж на кінці його, і від спеки його ніщо не заховається.
PS|19|7|(19-8) Господній Закон досконалий, він зміцнює душу. Свідчення Господа певне, воно недосвідченого умудряє.
PS|19|8|(19-9) Справедливі Господні накази, бо серце вони звеселяють. Заповідь Господа чиста, вона очі просвітлює.
PS|19|9|(19-10) Страх Господа чистий, він навіки стоїть. Присуди Господа правда, вони справедливі всі разом,
PS|19|10|(19-11) дорожчі вони понад золото і понад безліч щирого золота, і солодші за мед і за сік щільниковий,
PS|19|11|(19-12) і раб Твій у них бережкий, а в дотриманні їх нагорода велика.
PS|19|12|(19-13) А помилки хто зрозуміє? Від таємних очисть Ти мене,
PS|19|13|(19-14) і від свавільців Свого раба заховай, нехай не панують вони надо мною, тоді непорочним я буду, і від провини великої буду очищений.
PS|19|14|(19-15) Нехай будуть із волі Твоєї слова моїх уст, а думки мого серця перед лицем Твоїм, Господи, скеле моя й мій Спасителю!
PS|20|1|Для дириґетна хору. Псалом Давидів. (20-2) В день недолі озветься до тебе Господь, ім'я Бога Якового зробить сильним тебе!
PS|20|2|(20-3) Він пошле тобі поміч із святині, і з Сіону тебе підіпре!
PS|20|3|(20-4) Усі жертви твої пам'ятати Він буде, і буде вважати твоє цілопалення ситим. Села.
PS|20|4|(20-5) Він дасть тобі, як твоє серце бажає, і виповнить цілий твій задум!
PS|20|5|(20-6) Ми будем радіти спасінням Твоїм, і підіймемо прапор в ім'я Бога нашого, нехай Господь виконає всі прохання твої!
PS|20|6|(20-7) Тепер я пізнав, що спасає Господь помазанця Свого, дає йому відповідь з неба святого Свого могутніми чинами помічної правиці Своєї.
PS|20|7|(20-8) Одні колесницями хваляться, а інші кіньми, а ми будем хвалитись ім'ям Господа, нашого Бога:
PS|20|8|(20-9) вони похилились і впали, а ми стоїмо та ростемо на силах!
PS|20|9|(20-10) Господи, спаси! Хай озветься нам Цар у день нашого кликання!
PS|21|1|Для дириґетна хору. Псалом Давидів. (21-2) Господи, силою Твоєю веселиться цар, і спасінням Твоїм як він сильно радіє!
PS|21|2|(21-3) Ти йому дав бажання серця його, і прохання уст його не відмовив. Села.
PS|21|3|(21-4) Бо Ти його випередив благословеннями добра, на голову йому поклав корону зо щирого золота.
PS|21|4|(21-5) Життя він у Тебе просив, і дав Ти йому довголіття на вічні віки!
PS|21|5|(21-6) Слава велика його при Твоїй допомозі, хвалу та величність кладеш Ти на нього,
PS|21|6|(21-7) бо Ти вчиниш його благословенням вічним, звеселиш його радістю, як буде він разом з Тобою!
PS|21|7|(21-8) Цар має надію на Господа, у ласці Всевишнього не захитається він.
PS|21|8|(21-9) Знайде рука Твоя всіх ворогів Твоїх, знайде правиця Твоя Твоїх ненависників.
PS|21|9|(21-10) На час гніву Свого Ти їх учиниш огненною піччю, Господь гнівом Своїм їх понищить, і огонь пожере їх.
PS|21|10|(21-11) Ти вигубиш плід їхній із землі, а їхнє насіння з-поміж синів людських.
PS|21|11|(21-12) Бо нещастя на Тебе вони простягли, замишляли злу думку, якої здійснити не зможуть,
PS|21|12|(21-13) бо Ти їх обернеш плечима до нас, на тятивах Своїх міцно стріли поставиш на них.
PS|21|13|(21-14) Піднесися ж, о Господи, в силі Своїй, а ми будем співати й хвалити могутність Твою!
PS|22|1|Для дириґетна хору. На спів: „Ланя зорі досвітньої". Псалом Давидів. (22-2) Боже мій, Боже мій, нащо мене Ти покинув? Далекі слова мого зойку від спасіння мого!...
PS|22|2|(22-3) Мій Боже, взиваю я вдень, та Ти не озвешся, і кличу вночі, і спокою немає мені!
PS|22|3|(22-4) Та Ти Святий, пробуваєш на хвалах ізраїлевих!
PS|22|4|(22-5) На Тебе надіялись наші батьки, надіялися і Ти визволив їх.
PS|22|5|(22-6) До Тебе взивали вони і спасені були, на Тебе надіялися і не посоромились.
PS|22|6|(22-7) А я червяк, а не чоловік, посміховище людське й погорда в народі.
PS|22|7|(22-8) Всі, хто бачить мене, насміхаються з мене, розкривають роти, головою хитають!
PS|22|8|(22-9) Покладався на Господа він, хай же рятує його, нехай Той його визволить, він бо Його уподобав!
PS|22|9|(22-10) Бо з утроби Ти вивів мене, Ти безпечним мене учинив був на персах матері моєї!
PS|22|10|(22-11) На Тебе з утроби я зданий, від утроби матері моєї Ти мій Бог!
PS|22|11|(22-12) Не віддаляйся від мене, бо горе близьке, бо нема мені помічника!
PS|22|12|(22-13) Багато биків оточили мене, башанські бугаї обступили мене,
PS|22|13|(22-14) на мене розкрили вони свої пащі, як лев, що шматує й ричить!
PS|22|14|(22-15) Я розлитий, немов та вода, і всі кості мої поділились, стало серце моє, немов віск, розтопилось в моєму нутрі.
PS|22|15|(22-16) Висохла сила моя, як лушпиння, і прилип мій язик до мого піднебіння, і в порох смертельний поклав Ти мене.
PS|22|16|(22-17) Бо пси оточили мене... обліг мене натовп злочинців, прокололи вони мої руки та ноги мої...
PS|22|17|(22-18) Я висох, рахую всі кості свої, а вони придивляються й бачать нещастя в мені!
PS|22|18|(22-19) Вони ділять для себе одежу мою, а про шату мою жеребка вони кидають...
PS|22|19|(22-20) А Ти, Господи, не віддаляйся, Допомого моя, поспіши ж мені на оборону!
PS|22|20|(22-21) Від меча збережи мою душу, одиначку мою з руки пса!
PS|22|21|(22-22) Спаси мене від пащі лев'ячої, а вбогу мою від рогів буйволів.
PS|22|22|(22-23) Я звіщатиму Ймення Твоє своїм браттям, буду хвалити Тебе серед збору!
PS|22|23|(22-24) Хто боїться Господа, прославляйте Його, увесь Яковів роде шануйте Його, страхайтесь Його, все насіння ізраїлеве,
PS|22|24|(22-25) бо Він не погордував і не зневажив страждання убогого, і від нього обличчя Свого не сховав, а почув, як він кликав до Нього!
PS|22|25|(22-26) Від Тебе повстане хвала моя в зборі великім, принесу свої жертви в присутності тих, хто боїться Його,
PS|22|26|(22-27) будуть їсти покірні і ситими стануть, хвалитимуть Господа ті, хто шукає Його, буде жить серце ваше навіки!
PS|22|27|(22-28) Усі кінці землі спам'ятають, і до Господа вернуться, і вклоняться перед обличчям Його всі племена народів,
PS|22|28|(22-29) бо царство Господнє, і Він Пан над народами!
PS|22|29|(22-30) Будуть їсти й поклоняться всі багачі на землі, перед обличчям Його на коліна попадають всі, хто до пороху сходить і не може себе оживити!
PS|22|30|(22-31) Буде потомство служити Йому, й залічене буде навіки у Господа.
PS|22|31|(22-32) Прийдуть і будуть звіщать Його правду народові, який буде народжений, що Він це вчинив!
PS|23|1|Псалом Давидів. Господь то мій Пастир, тому в недостатку не буду,
PS|23|2|на пасовиськах зелених оселить мене, на тихую воду мене запровадить!
PS|23|3|Він душу мою відживляє, провадить мене ради Ймення Свого по стежках справедливости.
PS|23|4|Коли я піду хоча б навіть долиною смертної темряви, то не буду боятися злого, бо Ти при мені, Твоє жезло й Твій посох вони мене втішать!
PS|23|5|Ти передо мною трапезу зготовив при моїх ворогах, мою голову Ти намастив був оливою, моя чаша то надмір пиття!
PS|23|6|Тільки добро й милосердя мене супроводити будуть по всі дні мого життя, а я пробуватиму в домі Господньому довгі часи!
PS|24|1|Псалом Давидів. Господня земля, і все, що на ній, вселенна й мешканці її,
PS|24|2|бо заклав Він її на морях, і на річках її встановив.
PS|24|3|Хто зійде на гору Господню, і хто буде стояти на місці святому Його?
PS|24|4|У кого чисті руки та щиреє серце, і хто не нахиляв на марноту своєї душі, і хто не присягав на обману,
PS|24|5|нехай носить він благословення від Господа, а праведність від Бога спасіння свого!
PS|24|6|Таке покоління усіх, хто шукає Його, хто прагне обличчя Твого, Боже Яковів! Села.
PS|24|7|Піднесіте верхи свої, брами, і будьте відчинені, входи відвічні, і ввійде Цар слави!
PS|24|8|Хто ж то Цар слави? Господь сильний й могутній, Господь, що потужний в бою!
PS|24|9|Піднесіте верхи свої, брами, і піднесіте, входи відвічні, і ввійде Цар слави!
PS|24|10|Хто ж то Він, той Цар слави? Господь Саваот Він Цар слави! Села.
PS|25|1|Давидів. До Тебе підношу я, Господи, душу свою,
PS|25|2|Боже мій, я на Тебе надіюсь, нехай же я не засоромлюсь, нехай не радіють мої вороги ради мене!
PS|25|3|Не будуть також посоромлені всі, хто на Тебе надіється, та нехай посоромляться ті, хто на Тебе встає надаремно!
PS|25|4|Дороги Твої дай пізнати мені, Господи, стежками Своїми мене попровадь,
PS|25|5|провадь мене в правді Своїй і навчи Ти мене, бо Ти Бог спасіння мого, кожен день я на Тебе надіюсь!
PS|25|6|Пам'ятай милосердя Своє, о мій Господи, і ласки Свої, бо відвічні вони!
PS|25|7|Гріхи молодечого віку мого та провини мої не пригадуй, пам'ятай мене, Господи, в ласці Своїй через добрість Свою!
PS|25|8|Господь добрий та праведний, тому грішних навчає в дорозі,
PS|25|9|Він провадить покірних у правді, і лагідних навчає дороги Своєї!
PS|25|10|Всі Господні стежки милосердя та правда для тих, хто Його заповіта й свідоцтва додержує.
PS|25|11|Ради Ймення Свого, о Господи, прости мені прогріх, великий бо він!
PS|25|12|Хто той чоловік, що боїться він Господа? Він наставить його на дорогу, котру має вибрати:
PS|25|13|душа його житиме в щасті, і насіння його вспадку землю!
PS|25|14|Приязнь Господня до тих, хто боїться Його, і Свій заповіт Він звістить їм.
PS|25|15|Мої очі постійно до Господа, бо Він з пастки витягує ноги мої.
PS|25|16|Обернися до мене й помилуй мене, я ж бо самітний та бідний!
PS|25|17|Муки серця мого поширились, визволь мене з моїх утисків!
PS|25|18|Подивися на горе моє та на муку мою, і прости всі гріхи мої!
PS|25|19|Подивись на моїх ворогів, як їх стало багато, вони лютою ненавистю ненавидять мене!...
PS|25|20|Пильнуй же моєї душі та мене хорони, щоб не бути мені засоромленим, бо надіюсь на Тебе!
PS|25|21|Невинність та правда нехай оточають мене, бо надіюсь на Тебе!
PS|25|22|Визволи, Боже, ізраїля від усіх його утисків!
PS|26|1|Давидів. Суди мене, Господи, бо ходив я в своїй непорочності, і надіявсь на Господа, тому не спіткнуся!
PS|26|2|Перевір мене, Господи, і випробуй мене, перетопи мої нирки та серце моє,
PS|26|3|бо перед очима моїми Твоє милосердя, і в правді Твоїй я ходив.
PS|26|4|Не сидів я з людьми неправдивими, і не буду ходити з лукавими,
PS|26|5|я громаду злочинців зненавидів, і з грішниками я сидіти не буду.
PS|26|6|Умию в невинності руки свої, й обійду Твого, Господи, жертівника,
PS|26|7|щоб хвалу Тобі голосно виголосити, та звістити про всі чуда Твої.
PS|26|8|Господи, полюбив я оселю дому Твого, і місце перебування слави Твоєї.
PS|26|9|Не губи Ти моєї душі з нечестивими, та мого життя з кровожерами,
PS|26|10|що в руках їх злодійство, що їхня правиця наповнена підкупом.
PS|26|11|А я буду ходити в своїй непорочності, визволь мене та помилуй мене!
PS|26|12|Нога моя стала на рівному місці, на зборах я благословлятиму Господа!
PS|27|1|Давидів. Господь моє світло й спасіння моє, кого буду боятись? Господь то твердиня мого життя, кого буду лякатись?
PS|27|2|Коли будуть зближатись до мене злочинці, щоб жерти їм тіло моє, мої напасники та мої вороги, вони спотикнуться й попадають!...
PS|27|3|коли проти мене розложиться табір, то серце моє не злякається, коли проти мене повстане війна, я надіятись буду на те, на поміч Його!
PS|27|4|Одного прошу я від Господа, буду жадати того, щоб я міг пробувати в Господньому домі по всі дні свого життя, щоб я міг оглядати Господню приємність і в храмі Його пробувати!
PS|27|5|бо Він заховає мене дня нещастя в Своїй скинії, сховає мене потаємно в Своєму наметі, на скелю мене проведе!
PS|27|6|А тепер піднесеться моя голова понад ворогами моїми навколо мене, і я в Його скинії буду приносити жертви при відзвуках сурм, і я буду співати та грати Господеві!
PS|27|7|Почуй, Господи, голос мій, коли кличу, і помилуй мене, і озвися до мене!
PS|27|8|За Тебе промовило серце моє: Шукайте Мого лиця! тому, Господи, буду шукати обличчя Твого:
PS|27|9|не ховай же від мене обличчя Свого, у гніві Свого раба не відкинь! Ти був мені поміч, не кидай мене, і не лишай мене, Боже спасіння мого,
PS|27|10|бо мій батько та мати моя мене кинули, та Господь прийме мене!
PS|27|11|Дорогу Свою покажи мені, Господи, і провадь мене стежкою рівною, ради моїх ворогів!
PS|27|12|Не видай мене на сваволю моїх ворогів, бо повстали на мене ті свідки облудні та неправдомовці,
PS|27|13|немов би не вірував я, що в країні життя я побачу Господнє добро!
PS|27|14|Надійся на Господа, будь сильний, і хай буде міцне твоє серце, і надійся на Господа!
PS|28|1|Давидів. До Тебе я кличу, о Господи скеле моя, не будь же безмовним до мене, бо коли Ти замовкнеш до мене, я стану подібний до тих, що сходять до гробу...
PS|28|2|Почуй голос благання мого, як я кличу до Тебе, коли руки свої я підношу до храму святого Твого!
PS|28|3|Не хапай мене з грішними й тими, хто чинить безправство, хто плете своїм ближнім про мир, але зло в їхнім серці!
PS|28|4|Віддай їм за їхнім учинком, і за злом їхніх учинків, згідно з ділом їхніх рук Ти їм дай, верни їм заслужене ними,
PS|28|5|бо вони не вдивляються в чинність Господню й діла Його рук, нехай їх поруйнує, й нехай не будує Він їх!
PS|28|6|Благословенний Господь, бо Він почув голос благання мого!
PS|28|7|Господь моя сила та щит мій, на нього надіялось серце моє, й Він мені допоміг, і втішилося моє серце, і співом своїм я прославлю Його!
PS|28|8|Господь сила народу Свого, і захист спасіння Свого помазанця!
PS|28|9|Спаси Свій народ, і поблагослови спадщину Свою, і спаси їх, і піднось їх навіки!
PS|29|1|Псалом Давидів. Дайте Господу, Божі сини, дайте Господу славу та силу!
PS|29|2|Дайте Господу славу імення Його, у препишній святині впадіть перед Господом!
PS|29|3|Голос Господній над водами, Бог слави гримить, Господь над великими водами!
PS|29|4|Голос Господній із силою, голос Господній з величністю.
PS|29|5|Голос Господній ламає кедрини, голос Господній торощить кедрини ливанські.
PS|29|6|Він примусить скакати Ливан як теля, та Сиріон, мов молоду антилопу.
PS|29|7|Голос Господній викрешує полум'я огняне,
PS|29|8|голос Господній пустиню тремтіти примушує, Господь чинить пустелю Кадеша тремтячою.
PS|29|9|Голос Господній примушує лані тремтіти, й ліси обнажає, а в храмі Його все належне Йому виголошує: Слава!
PS|29|10|Господь пробував в час потопу, і буде Господь пробувати повік віку Царем!
PS|29|11|Господь подасть силу народу Своєму, Господь поблагословить миром народ Свій!
PS|30|1|Псалом Давидів. Пісня освячення дому. (30-2) Буду тебе величати, о Господи, бо Ти з глибини мене витяг, і не потішив моїх ворогів ради мене!
PS|30|2|(30-3) Господи, Боже мій, я кликав до Тебе, і мене вздоровив Ти.
PS|30|3|(30-4) Господи, вивів Ти душу мою із шеолу, Ти мене оживив, щоб в могилу не сходити мені!
PS|30|4|(30-5) Співайте Господеві, святії Його, й славте пам'ять святині Його!
PS|30|5|(30-6) Бо хвилю триває Він у гніві Своїм, все життя в Своїй ласці: буває увечорі плач, а радість на ранок!
PS|30|6|(30-7) А я говорив був у мирі своєму: Я не захитаюсь навіки!
PS|30|7|(30-8) Господи, в ласці Своїй Ти поставив мене на горі моїх сил. Як лице Своє Ти заховав, то збентежився я.
PS|30|8|(30-9) До Тебе я кличу, о Господи, і благаю я Господа:
PS|30|9|(30-10) Яка користь із крови моєї, коли я до гробу зійду? Чи хвалити Тебе буде порох? Чи він виявить правду Твою?
PS|30|10|(30-11) Почуй, Господи, і помилуй мене, Господи, будь мені помічником!
PS|30|11|(30-12) Ти перемінив мені плач мій на радість, жалобу мою розв'язав, і підперезав мене радістю,
PS|30|12|(30-13) щоб славу співала людина Тобі й не замовкла! Господи, Боже мій, повік славити буду Тебе!
PS|31|1|Для дириґетна хору. Псалом Давидів. (31-2) На Тебе надіюсь я, Господи, хай не буду повік засоромлений, визволь мене в Своїй правді!
PS|31|2|(31-3) Нахили Своє ухо до мене, скоро мене порятуй, стань для мене могутньою скелею, домом твердині, щоб спас Ти мене!
PS|31|3|(31-4) Бо ти скеля моя та твердиня моя, і ради Ймення Свого Ти будеш провадити мене й керувати мене!
PS|31|4|(31-5) Ти витягнеш з пастки мене, що на мене таємно поставили, бо Ти сила моя!
PS|31|5|(31-6) У руку Твою доручаю я духа свого, і Ти мене визволиш, Господи, Боже правди!
PS|31|6|(31-7) Я зненавидив всіх, хто шанує бовванів марних, я ж надіюсь на Господа.
PS|31|7|(31-8) Я буду радіти та тішитися в Твоїй милості, що побачив Ти горе моє, що приглянувся Ти до скорботи моєї душі,
PS|31|8|(31-9) і мене не віддав в руку ворога, на місці розлогім поставив Ти ноги мої!
PS|31|9|(31-10) Помилуй мене, Господи, бо тісно мені, від горя вже виснажилось моє око, душа моя й нутро моє,
PS|31|10|(31-11) бо скінчилось життя моє в смутку, а роки мої у квилінні, моя сила спіткнулася через мій гріх, і виснажились мої кості!
PS|31|11|(31-12) Я в усіх ворогів своїх став посміховищем, надто сусідам своїм, і страхіттям знайомим моїм, хто бачить надворі мене утікають від мене!
PS|31|12|(31-13) Я забутий у серці, немов той небіжчик, став я немов та розбита посудина...
PS|31|13|(31-14) Бо чую багато шептання, страхання навколо, як змовляються разом на мене, вони замишляють забрати мою душу,
PS|31|14|(31-15) а я покладаю надію на Тебе, о Господи, я кажу: Ти мій Бог!
PS|31|15|(31-16) В Твою руку кладу свою долю, Ти ж визволь мене від руки ворогів моїх і моїх переслідників!
PS|31|16|(31-17) Хай засяє обличчя Твоє на Твого раба, та спаси мене в ласці Своїй,
PS|31|17|(31-18) Господи, щоб не бути мені посоромленим, що кличу до Тебе! Нехай посоромлені будуть безбожні, хай замовкнуть та йдуть до шеолу,
PS|31|18|(31-19) нехай заніміють облудні уста, що гидоту говорять на праведного із пихою й погордою!
PS|31|19|(31-20) Яка величезна Твоя доброта, яку заховав Ти для тих, хто боїться Тебе, яку приготовив для тих, хто на Тебе надіється перед людськими синами!
PS|31|20|(31-21) Ти їх у заслоні обличчя Свого заховаєш від людських тенет, Ти їх від лихих язиків у наметі сховаєш!
PS|31|21|(31-22) Благословенний Господь, що вчинив мені милість чудовну Свою в оборонному місті!
PS|31|22|(31-23) А я говорив у своїм побентеженні: Я відрізаний з-перед очей Твоїх! Та дійсно Ти вислухав голос благання мого, коли я до Тебе взивав...
PS|31|23|(31-24) Любіть Господа, усі святії Його, стереже Господь вірних, а гордому з лишком відплачує.
PS|31|24|(31-25) Будьте сильні, і хай буде міцне ваше серце, усі, хто надію покладає на Господа!
PS|32|1|Давидів. Пісня навчальна. Блаженний, кому подарований злочин, кому гріх закрито,
PS|32|2|блаженна людина, що Господь їй гріха не залічить, що нема в її дусі лукавства!
PS|32|3|Коли я мовчав, спорохнявіли кості мої в цілоденному зойку моєму,
PS|32|4|бо рука Твоя вдень та вночі надо мною тяжить, і волога моя обернулась на літню посуху! Села.
PS|32|5|Я відкрив Тобі гріх свій, і не сховав був провини своєї. Я сказав був: Признаюся в проступках своїх перед Господом! і провину мого гріха Ти простив. Села.
PS|32|6|Тому кожен побожний відповідного часу молитися буде до Тебе, і навіть велика навала води не досягне до нього!
PS|32|7|Ти покрова моя, Ти від утиску будеш мене стерегти, Ти обгорнеш мене радістю спасіння! Села.
PS|32|8|Я зроблю тебе мудрим, і буду навчати тебе у дорозі, якою ти будеш ходити, Я дам тобі раду, Моє око вважає на тебе!
PS|32|9|Не будьте, як кінь, як той мул нерозумні, що їх треба приборкати оздобою їхньою вудилом і вуздечкою, як до тебе вони не зближаються.
PS|32|10|Багато хворіб на безбожного, хто ж надію свою покладає на Господа того милість оточує!
PS|32|11|Веселітесь у Господі, і тіштеся, праведні, і співайте із радістю, всі щиросерді!
PS|33|1|Співайте із радістю, праведні в Господі, бо щирим лицює хвала!
PS|33|2|Хваліть Господа гуслами, співайте Йому з десятиструнною арфою,
PS|33|3|заспівайте Йому нову пісню, гарно заграйте Йому з гуком сурем,
PS|33|4|бо щире Господнєє слово, і кожен чин Його вірний!
PS|33|5|Правду та суд Він кохає, і Господньої милости повна земля!
PS|33|6|Словом Господнім учинене небо, а подихом уст Його все його військо.
PS|33|7|Воду морську збирає Він, мов би до міху, безодні складає в коморах.
PS|33|8|Буде боятися Господа ціла земля, всі мешканці всесвіту будуть лякатись Його,
PS|33|9|бо сказав Він і сталось, наказав і з'явилось.
PS|33|10|Господь раду поганів понищить, понівечить мислі народів,
PS|33|11|а задум Господній навіки стоятиме, думки Його серця на вічні віки!
PS|33|12|Блаженний той люд, що Богом у нього Господь, блаженний народ, що Він вибрав його на спадок Собі!
PS|33|13|Господь споглядає з небес, і бачить усіх синів людських,
PS|33|14|приглядається з місця оселі Своєї до всіх, хто замешкує землю:
PS|33|15|Хто створив серце кожного з них, наглядає всі їхні діла!
PS|33|16|Немає царя, що його многість війська спасає, не врятується велетень великістю сили,
PS|33|17|для спасіння той кінь ненадійний, і великістю сили своєї він не збереже,
PS|33|18|ось око Господнє на тих, хто боїться Його, хто надію на милість Його покладає,
PS|33|19|щоб рятувати життя їхнє від смерти, і щоб за час голоду їх оживляти!
PS|33|20|Душа наша надію складає на Господа, Він наша поміч і щит наш,
PS|33|21|бо Ним радується наше серце, бо на Ймення святеє Його ми надію кладемо!
PS|33|22|Нехай Твоя милість, о Господи, буде на нас, коли покладаємо надію на Тебе!
PS|34|1|Давидів, коли він удавав був причинного перед Авімелехом, що вигнав його, і той пішов. (34-2) Я благословлятиму Господа кожного часу, хвала Йому завсіди в устах моїх!
PS|34|2|(34-3) Душа моя буде хвалитися Господом, хай це почують слухняні, і нехай звеселяться!
PS|34|3|(34-4) Зо мною звеличуйте Господа, і підносьте ім'я Його разом!
PS|34|4|(34-5) Шукав я був Господа, і Він озвався до мене, і від усіх небезпек мене визволив.
PS|34|5|(34-6) Приглядайтесь до Нього й засяєте, і не посоромляться ваші обличчя!
PS|34|6|(34-7) Цей убогий взивав, і Господь його вислухав, і від усіх його бід його визволив.
PS|34|7|(34-8) Ангол Господній табором стає кругом тих, хто боїться його, і визволює їх.
PS|34|8|(34-9) Скуштуйте й побачте, який добрий Господь, блаженна людина, що надію на Нього кладе!
PS|34|9|(34-10) Бійтеся Господа, всі святії Його, бо ті, що бояться Його, недостатку не мають!
PS|34|10|(34-11) Левчуки бідні й голодні, а ті, хто пошукує Господа, недостатку не чують в усьому добрі.
PS|34|11|(34-12) Ходіть, діти, послухайте мене, страху Господнього я вас навчу!
PS|34|12|(34-13) Хто та людина, що хоче життя, що любить дні довгі, щоб бачити добро?
PS|34|13|(34-14) Свого язика бережи від лихого, а уста свої від говорення підступу.
PS|34|14|(34-15) Відступися від злого і добре чини, миру шукай і женися за ним!
PS|34|15|(34-16) Очі Господні на праведних, уші ж Його на їхній зойк,
PS|34|16|(34-17) Господнє лице на злочинців, щоб винищити їхню пам'ять з землі.
PS|34|17|(34-18) Коли праведні кличуть, то їх чує Господь, і з усіх утисків їхніх визволює їх.
PS|34|18|(34-19) Господь зламаносердим близький, і впокорених духом спасає.
PS|34|19|(34-20) Багато лихого для праведного, та його визволяє Господь з них усіх:
PS|34|20|(34-21) Він пильнує всі кості його, із них жодна не зламається!
PS|34|21|(34-22) Зло безбожному смерть заподіє, і винними будуть усі, хто ненавидить праведного.
PS|34|22|(34-23) Господь визволить душу рабів Своїх, і винні не будуть усі, хто вдається до Нього!
PS|35|1|Давидів. Судися, о Господи, з тими, хто судиться зо мною воюй з тими, хто зо мною воює,
PS|35|2|візьми малого й великого щита, і встань мені на допомогу!
PS|35|3|Дістань списа, і дорогу замкни моїм напасникам, скажи до моєї душі: Я спасіння твоє!
PS|35|4|Нехай засоромляться й будуть поганьблені ті, хто чатує на душу мою; хай відступлять назад і нехай посоромляться ті, хто лихо мені замишляє.
PS|35|5|Бодай вони стали, немов та полова на вітрі, і Ангол Господній нехай їх жене;
PS|35|6|нехай буде дорога їхна темна й сковзька, і Ангол Господній нехай їх жене,
PS|35|7|бо вони безпричинно тенета свої розставляють на мене, яму копають безвинно на душу мою!
PS|35|8|Нехай нагла загибіль, якої не знає, на нього спаде, і сітка його, яку він наставив, хай зловить його у нагле нещастя, бодай він до нього упав!
PS|35|9|А душа моя в Господі буде радіти, звеселиться Його допомогою!
PS|35|10|Скажуть усі мої кості: Господи, хто подібний до Тебе? Ти рятуєш убогого від сильнішого над нього, покірного та бідаря від його дерія.
PS|35|11|Свідки встають неправдиві, чого я не знав питають мене,
PS|35|12|віддають мені злом за добро, осирочують душу мою!
PS|35|13|А я, як вони хворували були, зодягався в верету, душу свою мучив постом, молитва ж моя поверталась на лоно моє...
PS|35|14|Як приятель, буцім то брат він для мене, так я ходив, ніби був я в жалобі по матері, був я засмучений, схилений...
PS|35|15|А вони, як упав я, радіють та сходяться, напасники проти мене збираються, я ж не знаю про те; кричать, і не вмовкають,
PS|35|16|з дармоїдами та пересмішниками скрегочуть на мене своїми зубами...
PS|35|17|Господи, чи довго Ти будеш дивитись на це? Відверни мою душу від їхніх зубів, від отих левчуків одиначку мою!
PS|35|18|Я буду Тебе прославляти на зборах великих, буду Тебе вихваляти в численнім народі!
PS|35|19|Нехай з мене не тішаться ті, хто ворогує на мене безвинно, нехай ті не моргають очима, хто мене без причини ненавидить,
PS|35|20|бо говорять вони не про мир, але на спокійних у краї облудні слова вимишляють,
PS|35|21|свої уста на мене вони розкривають, говорять: Ага, ага! Наші очі це бачили!
PS|35|22|Ти бачив це, Господи, не помовчи ж, Господи, не віддаляйся від мене!
PS|35|23|Устань, і збудися на суд мій, Боже мій і Господи мій, на суперечку мою,
PS|35|24|розсуди Ти мене до Своїй справедливості, Господи, Боже мій, і нехай через мене не тішаться,
PS|35|25|нехай не говорять у серці своїм: Ага, його маємо ми, хай не кажуть вони: Ми його проковтнули...
PS|35|26|Нехай посоромляться та застидаються разом, хто з мого нещастя радіє, бодай вбрались у сором та в ганьбу, хто рота свого розкриває на мене!
PS|35|27|Хай співають та звеселяються ті, хто бажає мені правоти, і нехай кажуть завжди: Хай буде великий Господь, що миру бажає Своєму рабові!
PS|35|28|А язик мій звіщатиме правду Твою, славу Твою кожен день!
PS|36|1|Для диригенту хору. Раба Господнього Давида. (36-2) Грішне слово безбожного в серці моїм: Нема страху Божого перед очима його,
PS|36|2|(36-3) бо в очах своїх він до себе підлещується, щоб буцім то гріх свій знайти, щоб зненавидіти.
PS|36|3|(36-4) Слова його уст то марнота й обмана, перестав він бути мудрим, щоб чинити добро.
PS|36|4|(36-5) Беззаконство задумує він на постелі своїй, стає на дорозі недобрій, не цурається злого.
PS|36|5|(36-6) Господи, аж до небес милосердя Твоє, аж до хмар Твоя вірність,
PS|36|6|(36-7) Твоя справедливість немов гори Божі, Твої суди безодня велика, людину й худобу спасаєш Ти, Господи!
PS|36|7|(36-8) Яка дорога Твоя милість, о Боже, і ховаються людські сини в тіні Твоїх крил:
PS|36|8|(36-9) вони з ситости дому Твого напоюються, і Ти їх напуваєш з потока Своїх солодощів,
PS|36|9|(36-10) бо в Тебе джерело життя, в Твоїм світлі побачимо світло!
PS|36|10|(36-11) Продовж Свою милість на тих, хто знає Тебе, а правду Свою на людей щиросердих!
PS|36|11|(36-12) Нога пишних нехай не наступить на мене, і безбожна рука нехай не викидає мене!
PS|36|12|(36-13) Попадали там беззаконники, повалено їх і встати не зможуть.
PS|37|1|Давидів. Не розпалюйся гнівом своїм на злочинців, не май заздрости до беззаконних,
PS|37|2|бо вони, як трава, будуть скоро покошені, і мов та зелена билина пов'януть!
PS|37|3|Надійся на Господа й добре чини, землю замешкуй та правди дотримуй!
PS|37|4|Хай Господь буде розкіш твоя, і Він сповнить тобі твого серця бажання!
PS|37|5|На Господа здай дорогу свою, і на Нього надію клади, і Він зробить,
PS|37|6|і Він випровадить, немов світло, твою справедливість, а правду твою немов південь.
PS|37|7|Жди Господа мовчки й на Нього надійся, не розпалюйся гнівом на того, хто щасливою чинить дорогу свою, на людину, що виконує задуми злі.
PS|37|8|Повстримайсь від гніву й покинь пересердя, не розпалюйся лютістю, щоб чинити лиш зло,
PS|37|9|бо витяті будуть злочинці, а ті, хто вповає на Господа землю вспадкують!
PS|37|10|А ще трохи й не буде безбожного, і будеш дивитись на місце його і не буде його,
PS|37|11|а покірні вспадкують землю, і зарозкошують миром великим!
PS|37|12|Лихе замишляє безбожний на праведного, і скрегоче на нього своїми зубами,
PS|37|13|та Господь посміється із нього, бачить бо Він, що наближується його день!
PS|37|14|Безбожні меча добувають та лука свого натягають, щоб звалити нужденного й бідного, щоб порізати людей простої дороги,
PS|37|15|та ввійде їхній меч до їхнього власного серця, і поламані будуть їхні луки!
PS|37|16|Краще мале справедливого, ніж велике багатство безбожних, і то багатьох,
PS|37|17|бо зламані будуть рамена безбожних, а справедливих Господь підпирає!
PS|37|18|Знає Господь дні невинних, а їхня спадщина пробуде навіки,
PS|37|19|за лихоліття не будуть вони посоромлені, і за днів голоду ситими будуть.
PS|37|20|Бо загинуть безбожні, і Господні вороги, як овечий той лій, заникнуть, у димі заникнуть вони!
PS|37|21|Позичає безбожний і не віддає, а праведний милість висвідчує та роздає,
PS|37|22|бо благословенні від Нього вспадкують землю, а прокляті від Нього понищені будуть!
PS|37|23|Від Господа кроки людини побожної ставляться міцно, і Він любить дорогу її;
PS|37|24|коли ж упаде, то не буде покинена, бо руку її підпирає Господь.
PS|37|25|Я був молодий і постарівся, та не бачив я праведного, щоб опущений був, ні нащадків його, щоб хліба просили.
PS|37|26|Кожен день виявляє він милість та позичає, і над потомством його благословення.
PS|37|27|Ухиляйся від злого та добре чини, та й навіки живи!
PS|37|28|Бо любить Господь справедливість, і Він богобійних Своїх не покине, вони будуть навіки бережені, а насіння безбожних загине!
PS|37|29|Успадкують праведні землю, і повік будуть жити на ній.
PS|37|30|Уста праведного кажуть мудрість, язик же його промовляє про право,
PS|37|31|Закон Бога його в його серці, кроки його не спіткнуться.
PS|37|32|А безбожний чатує на праведного, і пильнує забити його,
PS|37|33|та Господь не зоставить його в руках того, і несправедливим не вчинить його, коли буде судити його.
PS|37|34|Надійся на Господа, та держися дороги Його, і піднесе Він тебе, щоб успадкувати землю, ти бачитимеш, як понижені будуть безбожні.
PS|37|35|Я бачив безбожного, що збуджував пострах, що розкоренився, немов саморосле зелене те дерево,
PS|37|36|та він проминув, й ось немає його, і шукав я його, й не знайшов!
PS|37|37|Бережи неповинного та дивися на праведного, бо людині спокою належить майбутність,
PS|37|38|переступники ж разом понищені будуть, майбутність безбожних загине!
PS|37|39|А спасіння праведних від Господа, Він їхня твердиня за час лихоліття,
PS|37|40|і Господь їм поможе та їх порятує, визволить їх від безбожних і їх збереже, бо вдавались до Нього вони!
PS|38|1|Псалом Давидів. На пам'ятку. (38-2) Господи, не карай мене в гніві Своїм, і не завдавай мені кари в Своїм пересерді,
PS|38|2|(38-3) бо прошили мене Твої стріли, і рука Твоя тяжко спустилась на мене...
PS|38|3|(38-4) Від гніву Твого нема цілого місця на тілі моїм, немає спокою в костях моїх через мій гріх,
PS|38|4|(38-5) бо провини мої переросли мою голову, як великий тягар, вони тяжчі над сили мої,
PS|38|5|(38-6) смердять та гниють мої рани з глупоти моєї...
PS|38|6|(38-7) Скорчений я, і над міру похилений, цілий день я тиняюсь сумний,
PS|38|7|(38-8) бо нутро моє повне запалення, і в тілі моїм нема цілого місця...
PS|38|8|(38-9) Обезсилений я й перемучений тяжко, ридаю від стогону серця свого...
PS|38|9|(38-10) Господи, всі бажання мої перед Тобою, зідхання ж моє не сховалось від Тебе.
PS|38|10|(38-11) Сильно тріпочеться серце моє, опустила мене моя сила, навіть ясність очей моїх і вона не зо мною...
PS|38|11|(38-12) Друзі мої й мої приятелі поставали здаля від моєї біди, а ближні мої поставали оподаль...
PS|38|12|(38-13) Тенета розставили ті, хто чатує на душу мою, а ті, хто бажає нещастя мені, говорять прокляття, і ввесь день вимишляють зрадливе!
PS|38|13|(38-14) А я, мов глухий, вже не чую, і мов той німий, який уст своїх не відкриває...
PS|38|14|(38-15) і я став, мов людина, що нічого не чує і в устах своїх оправдання не має,
PS|38|15|(38-16) бо на Тебе надіюся я, Господи, Ти відповіси, Господи, Боже мій!
PS|38|16|(38-17) Бо сказав я: Нехай не потішаться з мене, нехай не несуться вони понад мене, коли послизнеться нога моя!
PS|38|17|(38-18) Бо я до упадку готовий, і передо мною постійно недуга моя,
PS|38|18|(38-19) бо провину свою визнаю, журюся гріхом своїм я!
PS|38|19|(38-20) А мої вороги проживають, міцніють, і без причини помножилися мої недруги...
PS|38|20|(38-21) Ті ж, хто відплачує злом за добро, обчорнюють мене, бо женусь за добром...
PS|38|21|(38-22) Не покинь мене, Господи, Боже мій, не віддаляйся від мене,
PS|38|22|(38-23) поспіши мені на допомогу, Господи, Ти спасіння моє!
PS|39|1|Для дириґетна хору. Єдутуна. Псалом Давидів. (39-2) Я сказав: Пильнувати я буду дороги свої, щоб своїм язиком не грішити, накладу я вуздечку на уста свої, поки передо мною безбожний.
PS|39|2|(39-3) Занімів я в мовчанні, замовк про добро, а мій біль був подражнений.
PS|39|3|(39-4) Розпалилося серце моє у моєму нутрі, палає огонь від мого роздумування... Я став говорити своїм язиком:
PS|39|4|(39-5) Повідоми мене, Господи, про кінець мій та про днів моїх міру, яка то вона, нехай знаю, коли я помру!
PS|39|5|(39-6) Ось відміряв долонею Ти мої дні, а мій вік як ніщо проти Тебе, і тільки марнота сама кожна людина жива! Села.
PS|39|6|(39-7) У темноті лиш ходить людина, клопочеться тільки про марне: громадить вона, та не знає, хто звозити буде оте!
PS|39|7|(39-8) А тепер на що маю надіятись, Господи? Надія моя на Тебе вона!
PS|39|8|(39-9) Від усіх моїх прогріхів визволи мене, не чини мене посміхом для нерозумного!
PS|39|9|(39-10) Занімів я та уст своїх не відкриваю, бо Ти те вчинив,
PS|39|10|(39-11) забери Ти від мене Свій доторк, від порази Твоєї руки я кінчаюсь...
PS|39|11|(39-12) Ти караєш людину докорами за беззаконня, Ти знищив, як міль, привабність її, кожна людина направду марнота! Села.
PS|39|12|(39-13) Вислухай, Господи, молитву мою, і почуй благання моє, не будь мовчазний до моєї сльози, бо приходько я в Тебе, мандрівник, як батьки мої всі!
PS|39|13|(39-14) Відверни гнів від мене і я підкріплюся, перше ніж відійду, і не буде мене!
PS|40|1|Для дириґетна хору. Псалом Давидів. (40-2) Непохитно надіюсь на Господа, і Він прихилився до мене, і благання моє Він почув.
PS|40|2|(40-3) Витяг мене Він із згубної ями, із багна болотистого, і поставив на скелі ноги мої, і зміцнив мої стопи,
PS|40|3|(40-4) і дав пісню нову в мої уста, для нашого Бога хвалу, нехай бачать багато-хто й пострах хай мають, і хай вони мають надію, на Господа!
PS|40|4|(40-5) Блаженна людина, що Бога вчинила своєю твердинею, і не зверталась до пишних та тих, що вони до неправди схиляються!
PS|40|5|(40-6) Багато вчинив Ти, о Господи, Боже мій, Твої чуда й думки Твої тільки про нас, нема Тобі рівного! Я хотів би все це показати й про це розказати, та воно численніше, щоб можна його розповісти.
PS|40|6|(40-7) Жертви й приношення Ти не схотів, Ти розкрив мені уші, цілопалення й жертви покутної Ти не жадав.
PS|40|7|(40-8) Тоді я сказав: Ось я прийшов із звоєм книжки, про мене написаної.
PS|40|8|(40-9) Твою волю чинити, мій Боже, я хочу, і Закон Твій у мене в серці.
PS|40|9|(40-10) Я проповідував правду в великому зборі, ото, своїх уст не ув'язнюю я, Господи, знаєш Ти,
PS|40|10|(40-11) справедливість Твою не ховав я в середині серця свого, про вірність Твою та спасіння Твоє я звіщав, не таїв я про милість Твою та про правду Твою на великім зібранні.
PS|40|11|(40-12) Тому, Господи, не ув'язни милосердя Свого від мене, а милість та правда Твоя нехай завжди мене стережуть,
PS|40|12|(40-13) бо нещастя без ліку мене оточили, беззаконня мої досягли вже мене, так що й бачити не можу, вони численнішими стали за волосся на моїй голові, і серце моє опустило мене...
PS|40|13|(40-14) Зволь спасти мене, Господи, Господи, поспіши ж бо на поміч мені,
PS|40|14|(40-15) нехай посоромлені будуть, і хай зганьблені будуть усі, хто шукає моєї душі, щоб схопити її! Нехай подадуться назад, і нехай посоромлені будуть, хто бажає для мене лихого!
PS|40|15|(40-16) Бодай скам'яніли від сорому ті, хто говорить до мене: Ага! Ага!
PS|40|16|(40-17) Нехай тішаться та веселяться Тобою всі ті, хто шукає Тебе та хто любить спасіння Твоє, нехай завжди говорять: Хай буде великий Господь!
PS|40|17|(40-18) А я вбогий та бідний, за мене подбає Господь: моя поміч і мій оборонець то Ти, Боже мій, не спізняйся!
PS|41|1|Для дириґетна хору. Псалом Давидів. (41-2) Блаженний, хто дбає про вбогого, в день нещастя Господь порятує його!
PS|41|2|(41-3) Господь берегтиме його та його оживлятиме, буде блаженний такий на землі, і Він не видасть його на поталу його ворогам!
PS|41|3|(41-4) На ложі недуги подасть йому сили Господь, усе ложе йому перемінить в недузі його.
PS|41|4|(41-5) Я промовив був: Господи, май же Ти милість до мене, вилікуй душу мою, бо я перед Тобою згрішив!
PS|41|5|(41-6) Вороги мої кажуть на мене лихе: Коли вмре та загине імення його?
PS|41|6|(41-7) А коли хто приходить відвідати, мовить марне: його серце збирає для себе лихе, і як вийде надвір, то говорить про те...
PS|41|7|(41-8) Всі мої вороги між собою шепочуться разом на мене, на мене лихе замишляють:
PS|41|8|(41-9) Негідна річ тисне його, а що він поклався то більше не встане!...
PS|41|9|(41-10) Навіть приятель мій, на якого надіявся я, що мій хліб споживав, підняв проти мене п'яту!
PS|41|10|(41-11) Але, Господи, помилуй мене, і мене підійми, і я їм відплачу,
PS|41|11|(41-12) із того довідаюся, що Ти любиш мене, коли надо мною сурмити не буде мій ворог.
PS|41|12|(41-13) А я через невинність мою Ти підсилиш мене, і перед обличчям Своїм ти поставиш навіки мене!
PS|41|13|(41-14) Благословенний Господь, Бог ізраїлів, від віку й до віку! Амінь і амінь!
PS|42|1|Для дириґетна хору. Псалом навчальний, синів Кореєвих. (42-2) Як лине той олень до водних потоків, так лине до Тебе, о Боже, душа моя,
PS|42|2|(42-3) душа моя спрагнена Бога, Бога Живого! Коли я прийду й появлюсь перед Божим лицем?
PS|42|3|(42-4) Сльоза моя стала для мене поживою вдень та вночі, коли кажуть мені цілий день: Де твій Бог?
PS|42|4|(42-5) Як про це пригадаю, то душу свою виливаю, як я многолюдді ходив, і водив їх до Божого дому, із голосом співу й подяки святкового натовпу...
PS|42|5|(42-6) Чого, душе моя, ти сумуєш, і чого ти в мені непокоїшся? Май надію на Бога, бо я Йому буду ще дякувати за спасіння Його!
PS|42|6|(42-7) Мій Боже, душа моя тужить в мені, бо я пам'ятаю про Тебе з країни Йордану й Гермону, із гори із Міц'ар.
PS|42|7|(42-8) Прикликає безодня безодню на гуркіт Твоїх водоспадів, усі вали Твої й хвилі Твої перейшли надо мною.
PS|42|8|(42-9) Удень виявляє Господь Свою милість, уночі ж Його пісня зо мною, молитва до Бога мого життя!
PS|42|9|(42-10) Повім я до Бога: Ти Скеле моя, чому Ти про мене забув? Чого я блукаю сумний через утиск ворожий?
PS|42|10|(42-11) Ніби кості ламають мені, коли вороги мої лають мене, коли кажуть мені цілий день: Де твій Бог?
PS|42|11|(42-12) Чого, душе моя, ти сумуєш, і чого ти в мені непокоїшся? Май надію на Бога, бо я Йому буду ще дякувати за спасіння Його, мого Бога!
PS|43|1|Розсуди мене, Боже, й справуйся за справу мою із людьми небогобійними, визволь мене від людини обмани та кривди!
PS|43|2|Бож Бог Ти моєї твердині, чого ж Ти покинув мене? Чого я блукаю сумний через утиск ворожий?
PS|43|3|Пошли Своє світло та правду Свою, вони мене будуть провадити, вони запровадять мене до Твоєї святої гори та до місць пробування Твого.
PS|43|4|і нехай я дістанусь до Божого жертівника, до Бога розради й потіхи моєї, і буду на арфі хвалити Тебе, Боже, Боже Ти мій!
PS|43|5|Чого, душе моя, ти сумуєш, і чого ти в мені непокоїшся? Май надію на Бога, бо я Йому буду ще дякувати за спасіння Його, мого Бога!
PS|44|1|Для дириґетна хору. Синів Кореєвих. Псалом навчальний. (44-2) Боже, своїми ушима ми чули, наші батьки нам оповідали: велике Ти діло вчинив за їхніх днів, за днів стародавніх:
PS|44|2|(44-3) Ти вигнав поганів Своєю рукою, а їх осадив, понищив народи, а їх Ти поширив!
PS|44|3|(44-4) Не мечем бо своїм вони землю посіли, і їхнє рамено їм не помогло, а правиця Твоя та рамено Твоє, та Світло обличчя Твого, бо Ти їх уподобав!
PS|44|4|(44-5) Ти Сам Цар мій, о Боже, звели ж про спасіння для Якова:
PS|44|5|(44-6) Тобою поб'ємо своїх ворогів, ім'ям Твоїм будемо топтати повсталих на нас,
PS|44|6|(44-7) бо я буду надіятися не на лука свого, і мій меч не поможе мені,
PS|44|7|(44-8) але Ти нас спасеш від противників наших, і наших ненависників засоромиш!
PS|44|8|(44-9) Ми хвалимось Богом щодня, і повіки ім'я Твоє славимо, Села,
PS|44|9|(44-10) та однак Ти покинув і нас засоромив, і вже не виходиш із нашими військами:
PS|44|10|(44-11) Ти вчинив, що від ворога ми обернулись назад, а наші ненависники грабували собі наш маєток...
PS|44|11|(44-12) Ти віддав нас на поїд, немов тих овечок, і нас розпорошив посеред народів,
PS|44|12|(44-13) Ти за безцін продав Свій народ, і ціни йому не побільшив!
PS|44|13|(44-14) Ти нас нашим сусідам віддав на зневагу, на наругу та посміх для наших околиць,
PS|44|14|(44-15) Ти нас учинив за прислів'я поганам, і головою хитають народи на нас...
PS|44|15|(44-16) Передо мною щоденно безчестя моє, і сором вкриває обличчя моє,
PS|44|16|(44-17) через голос того, хто лає мене й проклинає, через ворога й месника...
PS|44|17|(44-18) Прийшло було все це на нас, та ми не забули про Тебе, й заповіту Твого не порушили,
PS|44|18|(44-19) не вступилось назад наше серце, і не відхилився наш крок від Твоєї дороги!
PS|44|19|(44-20) Хоч у місце шакалів Ти випхнув був нас, і прикрив був нас смертною тінню,
PS|44|20|(44-21) чи й тоді ми забули ім'я Бога нашого, і руки свої простягнули до Бога чужого?
PS|44|21|(44-22) Таж про те Бог довідається, бо Він знає таємності серця,
PS|44|22|(44-23) що нас побивають за Тебе щоденно, пораховано нас, як овечок жертовних...
PS|44|23|(44-24) Прокинься ж, для чого Ти, Господи, спиш? Пробудися, не кидай назавжди!
PS|44|24|(44-25) Для чого обличчя Своє Ти ховаєш, забуваєш про нашу недолю та нашу тісноту?
PS|44|25|(44-26) Бо душа наша знижилася аж до пороху, а живіт наш приліг до землі...
PS|44|26|(44-27) Устань же, о Помоче наша, і викупи нас через милість Свою!
PS|45|1|Для дириґетна хору. На „Лілеї". Синів Кореєвих. Псалом навчальний. Пісня любови. (45-2) Моє серце бринить добрим словом, проказую я: Для Царя мої твори, мій язик мов перо скорописця!
PS|45|2|(45-3) Ти кращий від людських синів, в Твоїх устах розлита краса та добро, тому благословив Бог навіки Тебе.
PS|45|3|(45-4) Прив'яжи до стегна Свого, Сильний, Свого меча, красу Свою та величність Свою,
PS|45|4|(45-5) і в величності Своїй сідай, та й верхи помчися за справи правди, і лагідности та справедливости, і навчить Тебе страшних чинів правиця Твоя!
PS|45|5|(45-6) Твої стріли нагострені, а від них під Тобою народи попадають, у серце Царських ворогів.
PS|45|6|(45-7) Престол Твій, о Боже, на вічні віки, берло правди берло Царства Твого.
PS|45|7|(45-8) Ти полюбив справедливість, а беззаконня зненавидів, тому намастив Тебе Бог, Твій Бог, оливою радости понад друзів Твоїх.
PS|45|8|(45-9) Миро, алое й кассія всі шати Твої, а з палат із слонової кости струни Тебе звеселили.
PS|45|9|(45-10) Серед скарбів Твоїх царські дочки, по правиці Твоїй стала цариця в офірському щирому золоті.
PS|45|10|(45-11) Слухай, дочко, й побач, і нахили своє ухо, і забудь свій народ і дім батька свого!
PS|45|11|(45-12) А Цар буде жадати твоєї краси, бо Він твій Господь, а ти до землі Йому кланяйся.
PS|45|12|(45-13) А Тирська дочка прийде з даром, будуть благати тебе найбагатші з народу.
PS|45|13|(45-14) Вся оздоба царської дочки усередині, шата ж її погаптована золотом.
PS|45|14|(45-15) У шати гаптовані вбрану провадять її до Царя, за нею дівчата, подруги її, до Тебе проваджені.
PS|45|15|(45-16) Провадять їх з радощами та потіхою, у палату царську вони війдуть.
PS|45|16|(45-17) Замість батьків Твоїх будуть сини Твої, їх по цілій землі Ти поставиш володарями.
PS|45|17|(45-18) Я буду ім'я Твоє згадувати по всіх поколіннях, тому то народи по вічні віки Тебе славити будуть!
PS|46|1|Для дириґетна хору. Синів Кореєвих. На спів „Аламот". Пісня. (46-2) Бог для нас охорона та сила, допомога в недолях, що часто трапляються,
PS|46|2|(46-3) тому не лякаємось ми, як трясеться земля, і коли гори зсуваються в серце морів!
PS|46|3|(46-4) Шумлять і киплять Його води, через велич Його тремтять гори. Села.
PS|46|4|(46-5) Річка, відноги її веселять місто Боже, найсвятіше із місць пробування Всевишнього.
PS|46|5|(46-6) Бог серед нього, нехай не хитається, Бог поможе йому, коли ранок настане.
PS|46|6|(46-7) Шуміли народи, хиталися царства, а Він голос подав Свій і земля розпливлася.
PS|46|7|(46-8) З нами Господь Саваот, наша твердиня Бог Яковів. Села.
PS|46|8|(46-9) ідіть, оглядайте Господні діла, які руйнування вчинив на землі!
PS|46|9|(46-10) Аж до краю землі припиняє Він війни, ламає Він лука й торощить списа, палить огнем колесниці!
PS|46|10|(46-11) Вгамуйтесь та знайте, що Бог Я, піднесусь між народами, піднесусь на землі!
PS|46|11|(46-12) З нами Господь Саваот, наша твердиня Бог Яковів! Села.
PS|47|1|Для дириґетна хору. Синів Кореєвих. Псалом. (47-2) Всі народи, плещіть у долоні, покликуйте Богові голосом радости,
PS|47|2|(47-3) грізний бо Всевишній Господь, Цар великий всієї землі!
PS|47|3|(47-4) Він народи під нас підбиває, а поган нам під ноги,
PS|47|4|(47-5) Він нашу спадщину для нас вибирає, величність для Якова, що його полюбив. Села.
PS|47|5|(47-6) Бог виступає при радісних окриках, Господь при голосі рога.
PS|47|6|(47-7) Співайте Богові нашому, співайте, співайте Цареві нашому, співайте,
PS|47|7|(47-8) бо Бог Цар усієї землі, співайте навчальний псалом!
PS|47|8|(47-9) Бог зацарював над народами, Бог сів на святому Своєму престолі!
PS|47|9|(47-10) Зібрались владики народів, народ Бога Авраамового, як Божі щити на землі, між ними Він сильно звеличений!
PS|48|1|Пісня. Псалом синів Кореєвих. (48-2) Великий Господь і прославлений вельми в місті нашого Бога, на святій Своїй горі!
PS|48|2|(48-3) Препишна країна, розрада всієї землі, то Сіонська гора, на північних околицях, місто Царя можновладного!
PS|48|3|(48-4) Бог у храмах Своїх, за твердиню Він знаний.
PS|48|4|(48-5) Бо царі ось зібрались, ішли вони разом,
PS|48|5|(48-6) але, як побачили, то здивувались, полякалися та й розпорошились...
PS|48|6|(48-7) Обгорнув їх там страх, немов біль породіллю;
PS|48|7|(48-8) Ти східнім вітром розбив кораблі ті Таршіські.
PS|48|8|(48-9) Як ми чули, так бачили в місті Господа Саваота, у місті нашого Бога, Бог міцно поставить навіки його! Села.
PS|48|9|(48-10) Розмишляли ми, Боже, про милість Твою серед храму Твого.
PS|48|10|(48-11) Як ім'я Твоє, Боже, так слава Твоя аж по кінці землі, справедливости повна правиця Твоя!
PS|48|11|(48-12) Нехай веселиться Сіонська гора, Юдині дочки хай тішаться через Твої правосуддя.
PS|48|12|(48-13) Оточіте Сіон й обступіте його, полічіть його башти,
PS|48|13|(48-14) зверніте увагу на вала його, високість палати його пообмірюйте, щоб розповісти поколінню наступному,
PS|48|14|(48-15) бо Цей Бог то наш Бог на вічні віки, Він буде провадити нас аж до смерти!
PS|49|1|Для дириґетна хору. Синів Кореєвих. Псалом. (49-2) Слухайте це, всі народи, візьміть до ушей, усі мешканці всесвіту,
PS|49|2|(49-3) і людські сини й сини мужів, разом багатий та вбогий,
PS|49|3|(49-4) мої уста казатимуть мудрість, думка ж серця мого розумність,
PS|49|4|(49-5) нахилю своє ухо до приказки, розв'яжу свою загадку лірою!
PS|49|5|(49-6) Чому маю боятись у день лихоліття, як стане круг мене неправда моїх ошуканців,
PS|49|6|(49-7) які на багатство своє покладають надію, і своїми достатками хваляться?
PS|49|7|(49-8) Але жодна людина не викупить брата, не дасть його викупу Богові,
PS|49|8|(49-9) бо викуп їхніх душ дорогий, і не перестане навіки,
PS|49|9|(49-10) щоб міг він ще жити навіки й не бачити гробу!
PS|49|10|(49-11) Та люди побачать, що мудрі вмирають так само, як гинуть невіглас та неук, і лишають для інших багатство своє...
PS|49|11|(49-12) Вони думають, ніби доми їхні навіки, місця їхнього замешкання з роду до роду, іменами своїми звуть землі,
PS|49|12|(49-13) та не зостається в пошані людина, подібна худобі, що гине!
PS|49|13|(49-14) Така їхня дорога глупота для них, та за ними йдуть ті, хто кохає їхню думку. Села.
PS|49|14|(49-15) Вони зійдуть в шеол, і смерть їх пасе, немов вівці, а праведники запанують над ними від рання; подоба їхня знищиться, шеол буде мешканням для них...
PS|49|15|(49-16) Та визволить Бог мою душу із влади шеолу, бо Він мене візьме! Села.
PS|49|16|(49-17) Не лякайся, коли багатіє людина, коли збільшується слава дому її,
PS|49|17|(49-18) бо, вмираючи, не забере вона всього, її слава не піде за нею!
PS|49|18|(49-19) Хоч вона свою душу за життя свого хвалить, і славлять тебе, як для себе ти чиниш добро,
PS|49|19|(49-20) вона прийде до роду батьків своїх, що світла вони не побачать навіки!
PS|49|20|(49-21) Людина в пошані, але нерозумна, подібна худобі, що гине!
PS|50|1|Псалом Асафів. Прорік Бог над Богами Господь, і землю покликав від схід сонця і аж до заходу його.
PS|50|2|із Сіону, корони краси, Бог явився в промінні!
PS|50|3|Приходить наш Бог, і не буде мовчати: палючий огонь перед Ним, а круг Нього все буриться сильно!
PS|50|4|Він покличе згори небеса, і землю народ Свій судити:
PS|50|5|Позбирайте для Мене побожних Моїх, що над жертвою склали заповіта зо Мною.
PS|50|6|і небеса звістять правду Його, що Бог Він суддя. Села.
PS|50|7|Слухай же ти, Мій народе, бо буду ось Я говорити, ізраїлеві, і буду свідчить на тебе: Бог, Бог твій Я!
PS|50|8|Я буду картати тебе не за жертви твої, бо все передо Мною твої цілопалення,
PS|50|9|не візьму Я бичка з твого дому, ні козлів із кошар твоїх,
PS|50|10|бо належить Мені вся лісна звірина та худоба із тисячі гір,
PS|50|11|Я знаю все птаство гірське, і звір польовий при Мені!
PS|50|12|Якби був Я голодний, тобі б не сказав, бо Моя вся вселенна й усе, що на ній!
PS|50|13|Чи Я м'ясо бичків споживаю, і чи п'ю кров козлів?
PS|50|14|Принось Богові в жертву подяку, і виконуй свої обітниці Всевишньому,
PS|50|15|і до Мене поклич в день недолі, Я тебе порятую, ти ж прославиш Мене!
PS|50|16|А до грішника Бог промовляє: Чого про устави Мої розповідаєш, і чого заповіта Мого на устах своїх носиш?
PS|50|17|Ти ж науку зненавидів, і поза себе слова Мої викинув.
PS|50|18|Як ти злодія бачив, то бігав із ним, і з перелюбниками накладав.
PS|50|19|Свої уста пускаєш на зло, і язик твій оману плете.
PS|50|20|Ти сидиш, проти брата свого наговорюєш, поголоски пускаєш про сина своєї матері...
PS|50|21|Оце ти робив, Я ж мовчав, і ти думав, що Я такий самий, як ти. Тому буду картати тебе, і виложу все перед очі твої!
PS|50|22|Зрозумійте ж це ви, що забуваєте Бога, щоб Я не схопив, бо не буде кому рятувати!
PS|50|23|Хто жертву подяки приносить, той шанує Мене; а хто на дорогу Свою уважає, Боже спасіння йому покажу!
PS|51|1|Для дириґетна хору. Псалом Давидів. (51-3) Помилуй мене, Боже, з великої милости Твоєї, і з великого милосердя Свого загладь беззаконня мої!
PS|51|2|(51-4) Обмий мене зовсім з мого беззаконня, й очисти мене від мого гріха,
PS|51|3|(51-5) бо свої беззаконня я знаю, а мій гріх передо мною постійно.
PS|51|4|(51-6) Тобі, одному Тобі я згрішив, і перед очима Твоїми лукаве вчинив, тому справедливий Ти будеш у мові Своїй, бездоганний у суді Своїм.
PS|51|5|(51-7) Отож я в беззаконні народжений, і в гріху зачала мене мати моя.
PS|51|6|(51-8) Ото, полюбив єси правду в глибинах, і в таємних речах виявляєш премудрість мені.
PS|51|7|(51-9) Очисти ісопом мене, і буду я чистий, обмий Ти мене і я стану біліший від снігу.
PS|51|8|(51-10) Дай почути мені втіху й радість, і радітимуть кості, що Ти покрушив.
PS|51|9|(51-11) Обличчя Своє заховай від гріхів моїх, і всі беззаконня мої позагладжуй.
PS|51|10|(51-12) Серце чисте створи мені, Боже, і тривалого духа в моєму нутрі віднови.
PS|51|11|(51-13) Не відкинь мене від Свого лиця, й не бери Свого Духа Святого від мене.
PS|51|12|(51-14) Верни мені радість спасіння Твого, і з лагідним духом підтримай мене.
PS|51|13|(51-15) Я буду навчати беззаконців доріг Твоїх, і навернуться грішні до Тебе.
PS|51|14|(51-16) Визволь мене від переступу кровного, Боже, Боже спасіння мого, мій язик нехай славить Твою справедливість!
PS|51|15|(51-17) Господи, відкрий мої уста, і язик мій звістить Тобі хвалу,
PS|51|16|(51-18) бо Ти жертви не прагнеш, а дам цілопалення, то не любе воно Тобі буде.
PS|51|17|(51-19) Жертва Богові зламаний дух; серцем зламаним та упокореним Ти не погордуєш, Боже!
PS|51|18|(51-20) Ущаслив Своїм благоволінням Сіон, збудуй мури для Єрусалиму,
PS|51|19|(51-21) тоді Ти полюбиш Собі жертви правди, цілопалення та приношення, тоді покладуть на Твій вівтар тельців!
PS|52|1|Для дириґетна хору. Псалом навчальний Давидів. (52-3) Чого хвалишся злом, о могутній? Цілий день Божа милість зо мною.
PS|52|2|(52-4) Замишляє лукавство язик твій, як та бритва нагострена ти, що чиниш обману!
PS|52|3|(52-5) Ти зло полюбив над добро, а неправду більш, як правду казати, Села,
PS|52|4|(52-6) ти любиш усякі шкідливі слова, ти язику обманний!
PS|52|5|(52-7) Отож, Бог зруйнує назавжди тебе, тебе викине й вирве з намету тебе, й тебе викоренить із країни життя. Села.
PS|52|6|(52-8) і побачать це праведні, й будуть боятись, і будуть сміятися з нього:
PS|52|7|(52-9) Ось муж, що Бога не чинить своєю твердинею, та на великість багатства свого покладає надію, втікає до злого свого...
PS|52|8|(52-10) А я як зелена оливка у Божому домі, надіюсь на Божую милість на вічні віки!
PS|52|9|(52-11) Буду славити вічно Тебе, що вчинив Ти оце, і про ймення Твоє буду звіщати побожним Твоїм, що добре воно!
PS|53|1|Для дириґетна хору. На „Махалат". Навчальний псалом. Давидів. (53-2) Безумний говорить у серці своїм: Нема Бога! Зіпсулись вони, і несправедливість обридливу чинять, нема доброчинця!...
PS|53|2|(53-3) Бог зорить із неба на людських синів, щоб побачити, чи є там розумний, що Бога шукає.
PS|53|3|(53-4) Усі повідступали, разом стали огидними, нема доброчинця, нема ні одного!...
PS|53|4|(53-5) Чи ж не розуміють оті, хто беззаконня вчиняє, що мій люд поїдають? Вони споживають хліб Божий, та не кличуть Його!
PS|53|5|(53-6) Тоді настрашилися страхом вони, хоч страху не було, бо розсипав Бог кості того, хто тебе оточив був, ти їх посоромив, бо ними погордував Бог!
PS|53|6|(53-7) Аби то Він дав із Сіону спасіння ізраїлеві! Як долю Свого народу поверне Господь, то радітиме Яків, утішатися буде ізраїль!
PS|54|1|Для дириґетна хору. На неґінах. Псалом навчальний Давидів, (54-2) як зіфіяни прийшли були та сказали Саулові: „Ось Давид поміж нами ховається!" (54-3) Спаси мене, Боже, іменням Своїм, і міццю Своєю мене оправдай!
PS|54|2|(54-4) Вислухай, Боже, молитву мою, нахили Своє ухо до слів моїх уст,
PS|54|3|(54-5) бо чужинці повстали на мене, розбишаки ж шукають моєї душі, вони Бога не ставили перед собою. Села.
PS|54|4|(54-6) Ось Бог помагає мені, Господь серед тих, хто підтримує душу мою.
PS|54|5|(54-7) Хай повернеться зло на моїх ворогів, Своєю правдою винищи їх.
PS|54|6|(54-8) В добровільному дарі я жертву Тобі принесу, ім'я Твоє, Господи, славити буду, що добре воно,
PS|54|7|(54-9) бо мене воно визволило від усяких нещасть, і я бачу занепад моїх ворогів!
PS|55|1|Для дириґетна хору. На неґінах. Псалом навчальний Давидів. (55-2) Вислухай, Боже, молитву мою й від благання мого не ховайся!
PS|55|2|(55-3) Прислухайсь до мене й подай мені відповідь, я блукаю у смутку своїм і стогну,
PS|55|3|(55-4) від крику ворожого, від утисків грішного, бо гріх накидають на мене вони, і в гніві мене переслідують...
PS|55|4|(55-5) Тремтить моє серце в мені, і страхи смертельні напали на мене,
PS|55|5|(55-6) страх та тремтіння на мене найшли, і тривога мене обгорнула...
PS|55|6|(55-7) казав я: Коли б я мав крила, немов та голубка, то я полетів би й спочив!
PS|55|7|(55-8) Отож, помандрую далеко, пробуватиму я на пустині. Села.
PS|55|8|(55-9) Поспішу собі, щоб утекти перед вітром бурхливим та бурею...
PS|55|9|(55-10) Вигуби, Господи, та погуби язика їхнього, бо в місті я бачив насильство та сварку,
PS|55|10|(55-11) вони ходять удень та вночі коло нього на мурах його, а гріх та неправда всередині в ньому,
PS|55|11|(55-12) нещастя всередині в ньому, а з вулиць його не виходять насилля й обмана,
PS|55|12|(55-13) бож не ворог злорічить на мене, це я переніс би, і не ненависник мій побільшивсь надо мною, я сховався б від нього,
PS|55|13|(55-14) але ти, чоловік мені рівня, мій приятель близький і знайомий мені,
PS|55|14|(55-15) з яким солодко щиру розмову провадимо, і ходимо до Божого дому серед бурхливого натовпу...
PS|55|15|(55-16) Нехай же впаде на них смерть, нехай зійдуть вони до шеолу живими, бо зло в їхнім мешканні, у їхній середині!
PS|55|16|(55-17) Я кличу до Бога, і Господь урятує мене:
PS|55|17|(55-18) увечорі, вранці й опівдні я скаржусь й зідхаю, і Він вислухає мого голосу!
PS|55|18|(55-19) У мирі Він викупить душу мою, щоб до мене вони не зближались, бо багато було їх на мене!
PS|55|19|(55-20) Бог вислухає, і їм Той відповість, Хто відвіку сидить на престолі, Села, бо немає у них перемін, і Бога вони не бояться,
PS|55|20|(55-21) ворог витягнув руки свої проти тих, що в спокої жили з ним, він зганьбив заповіта свого,
PS|55|21|(55-22) його уста гладенькі, як масло, та сварка у серці його, від оливи м'якіші слова його, та вони як мечі ті оголені!...
PS|55|22|(55-23) Свого тягара поклади ти на Господа, і тебе Він підтримає, Він ніколи не дасть захитатися праведному!
PS|55|23|(55-24) А Ти їх, Боже мій, поскидаєш до ями погибелі! Люди чинів кривавих й обмани, бодай своїх днів вони не дожили навіть до половини, а я покладаю надію на Тебе!
PS|56|1|Для дириґетна хору. На „Німа голубка в далечині". Золотий Давидів псалом, коли филистимляни захопили були його в Ґаті. (56-2) Помилуй мене, Боже, бо топче мене чоловік, цілий день він воює та тисне мене!
PS|56|2|(56-3) Чатують мої вороги цілий день, бо багато таких, що воюють завзято на мене!
PS|56|3|(56-4) Того дня, коли страх обгортає мене, я надію на Тебе кладу,
PS|56|4|(56-5) я в Бозі хвалитиму слово Його, на Бога надію кладу, й не боюся, що тіло учинить мені?
PS|56|5|(56-6) Цілий день біль приносять слова мої, усі їхні думки проти мене на зло:
PS|56|6|(56-7) слідкують, ховаються, пильнують вони мої стопи... Як чатують на душу мою,
PS|56|7|(56-8) так Ти через гріх віджени їх, пониж, Боже, людей в Своїм гніві!
PS|56|8|(56-9) Полічив Ти тиняння моє, помісти ж мої сльози перед Собою, чи ж вони не записані в книзі Твоїй?
PS|56|9|(56-10) Тоді то мої вороги повтікають назад, того дня, як я кликати буду. Те я знаю, що Бог при мені,
PS|56|10|(56-11) і в Бозі я справу свою докінчу, докінчу я в Господі справу!
PS|56|11|(56-12) На Бога надію кладу й не боюсь, що людина учинить мені?
PS|56|12|(56-13) На мені зостаються, о Боже, присяги Тобі, та для Тебе я виповню жертви хвали.
PS|56|13|(56-14) Як Ти спас мою душу від смерти, то хіба ж не спасеш моїх ніг від падіння, щоб у світлі життя я ходив перед Богом?
PS|57|1|Для дириґетна хору. На спів: „Не вигуби". Золотий псалом Давидів, коли він утікав від Саула в печеру. (57-2) Помилуй мене, Боже, помилуй мене, бо до Тебе вдається душа моя, і в тіні Твоїх крил я сховаюсь, аж поки нещастя мине!
PS|57|2|(57-3) Я кличу до Бога Всевишнього, до Бога, що чинить для мене добро.
PS|57|3|(57-4) Він пошле з небес і врятує мене, Він поганьбить того, хто чатує на мене. Села. Бог пошле Свою милість та правду Свою
PS|57|4|(57-5) на душу мою. Знаходжуся я серед левів, що людських синів пожирають, їхні зуби як спис той та стріли, а їхній язик гострий меч.
PS|57|5|(57-6) Піднесися ж, о Боже, над небо, а слава Твоя над всією землею!
PS|57|6|(57-7) Вороги приготовили пастку для стіп моїх, душу мою нахилили, вони викопали вовчу яму для мене, і попадали в неї самі! Села.
PS|57|7|(57-8) Моє серце зміцнилося, Боже, зміцнилося серце моє, я буду співати та славити Тебе!
PS|57|8|(57-9) Збудися ж ти, хвало моя, пробудися ж ти, арфо та цитро, я буду будити досвітню зорю!
PS|57|9|(57-10) Я буду Тебе вихваляти, о Господи, серед народів, я буду співати Тобі між племенами,
PS|57|10|(57-11) бо Твоє милосердя велике воно аж до неба, а правда Твоя аж до хмар!
PS|57|11|(57-12) Піднесися ж, о Боже, над небо, а слава Твоя над всією землею!
PS|58|1|Для дириґетна хору. На спів: „Не вигуби". Золотий псалом Давидів. (58-2) Чи ж то справді ви, можні, говорите правду, чи людських синів слушно судите?
PS|58|2|(58-3) Отже, у серці ви чините кривди, дорогу насильства рук ваших торуєте ви на землі.
PS|58|3|(58-4) Від лоня ще матернього вже віддалені несправедливі, з утроби ще матерньої заблудилися неправдомовці,
PS|58|4|(58-5) їхня отрута така, як отрута зміїна, як отрута глухої гадюки, що ухо своє затуляє,
PS|58|5|(58-6) що не слухає голосу заклиначів, чарівника, в чарах вправного!
PS|58|6|(58-7) Поруйнуй, Боже, зуби їхні в їхніх устах, левчукам розбий, Господи, щелепи,
PS|58|7|(58-8) нехай розпливуться, немов та вода, що собі розтікається, хай пов'януть вони, як трава по дорозі,
PS|58|8|(58-9) бодай стали, немов той слимак, що в своїй слизоті розпускається, щоб сонця не бачили, як мертвий отой плід у жінки!
PS|58|9|(58-10) Поки почують тернину запалену ваші горшки, нехай буря її рознесе, чи свіжу, чи спалену!
PS|58|10|(58-11) А праведний тішитись буде, бо помсту побачить, у крові безбожного стопи свої він обмиє!
PS|58|11|(58-12) і скаже людина: Поправді є плід справедливому, справді є Бог, суддя на землі!
PS|59|1|Для дириґетна хору. На спів: „Не вигуби". Золотий псалом Давидів, коли послав був Саул, і стерегли його дім. щоб убити його. (59-2) Визволь мене від моїх ворогів, о мій Боже, від напасників моїх охорони Ти мене!
PS|59|2|(59-3) Визволь мене від злочинців, і спаси мене від кровожерних,
PS|59|3|(59-4) бо ось причаїлись на душу мою, на мене збираються сильні, не моя в тім провина, о Господи, і не мій гріх!
PS|59|4|(59-5) Без моєї провини вони он збігаються та готуються, устань же назустріч мені та побач!
PS|59|5|(59-6) і Ти, Господи, Боже Саваоте, Боже ізраїлів, збудися, щоб покарати всіх поган, і не помилуй нікого із зрадників злих! Села.
PS|59|6|(59-7) Надвечір вони повертаються, скиглять, як пес, і перебігають по місту,
PS|59|7|(59-8) й ось слова вивергають устами своїми, мечі в їхніх губах, та хто це почує...
PS|59|8|(59-9) Але посмієшся з них, Господи, і всіх поган засоромиш!
PS|59|9|(59-10) Твердине моя, я Тебе пильнуватиму, бо Бог оборона моя!
PS|59|10|(59-11) Мій Бог, Його милість мене попередила, Бог учинить мені, що побачу падіння своїх ворогів!
PS|59|11|(59-12) Не вбивай їх, щоб народ мій цього не забув, міццю Своєю розвій їх і зниж їх, о щите наш, Господи!
PS|59|12|(59-13) Гріх їхніх уст слово губ їхніх, і нехай вони схоплені будуть своєю пихою, і за клятву й брехню, яку кажуть!
PS|59|13|(59-14) У гніві їх знищ, знищ і хай їх не буде, і хай знають вони, що царює Бог в Якові, аж до кінців землі! Села.
PS|59|14|(59-15) А надвечір вони повертаються, скиглять, як пес, і перебігають по місту.
PS|59|15|(59-16) Вони вештатись будуть, щоб їсти, коли ж не наїдяться, то скаржитись будуть.
PS|59|16|(59-17) А я буду співати про силу Твою, буду радісно вранці хвалити Твою милість, бо для мене Ти був в день недолі моєї твердинею й захистом!
PS|59|17|(59-18) Твердине моя, до Тебе співати я буду, бо Бог оборона моя, милостивий мій Боже!
PS|60|1|Для дириґетна хору. На спів: „Лілея свідчення". Золотий псалом Давидів для навчання, (60-2) коли він підпалив був Арам двух річок і Арам Цови, і вернувся Йоав і побив Едома в Соляній долині, дванадцять тисяч. (60-3) Боже, покинув Ти нас, розпорошив Ти нас, Ти нагнівався був, повернися ж до нас!
PS|60|2|(60-4) Ти землею затряс, і її розірвав, уздоров же уламки її, бо вона захиталась!
PS|60|3|(60-5) Ти вчинив, що народ Твій побачив тяжке, напоїв нас отрутним вином...
PS|60|4|(60-6) Ти дав прапора тим, хто боїться Тебе, щоб збирались вони перед правдою. Села.
PS|60|5|(60-7) Щоб любі Твої були визволені, Своєю правицею допоможи, й обізвися до нас!
PS|60|6|(60-8) У святині Своїй Бог промовив: Нехай розвеселюсь, розділю Я Сихем і долину Суккотську поміряю!
PS|60|7|(60-9) Належить Мені Ґілеад, Мені Манасія, а Єфрем охорона Моїй голові, Юда берло Моє.
PS|60|8|(60-10) Моав то мідниця Мого миття, на Едом узуттям Своїм кину, филистею, вигукуй для Мене із радістю!
PS|60|9|(60-11) Хто мене запровадить до міста твердинного, хто до Едому мене попровадить?
PS|60|10|(60-12) Хіба ж Ти покинув нас, Боже, і серед нашого війська не вийдеш вже, Боже?
PS|60|11|(60-13) Подай же нам поміч на ворога, людська бо поміч марнота!
PS|60|12|(60-14) Ми мужність виявимо в Бозі, і Він потопче противників наших!
PS|61|1|Для дириґетна хору. На струннім інструменті. Псалом Давидів. (61-2) Вислухай, Боже, благання моє, почуй же молитву мою,
PS|61|2|(61-3) я кличу до Тебе від краю землі, коли серце моє омліває! На скелю, що вища від мене, мене попровадь,
PS|61|3|(61-4) бо для мене Ти став пристановищем, баштою сильною супроти ворога!
PS|61|4|(61-5) Хай я оселюся навіки в наметі Твоїм, в укритті Твоїх крил заховаюся, Села,
PS|61|5|(61-6) бо Ти, Боже, почув обітниці мої, Ти дав спадщину тим, хто Ймення Твого боїться!
PS|61|6|(61-7) Цареві примнож дні до днів, продовж роки йому немов вічні віки,
PS|61|7|(61-8) нехай він перед Божим лицем пробуває навіки, хай милість та правда його стережуть!
PS|61|8|(61-9) Отак буду співати я завжди про Ймення Твоє, виконувати буду щоденно обіти свої!
PS|62|1|Для дириґетна хору. Для Єдутуна. Псалом Давидів. (62-2) Тільки від Бога чекай у мовчанні, о душе моя, від Нього спасіння моє!
PS|62|2|(62-3) Тільки Він моя скеля й спасіння моє, Він твердиня моя, тому не захитаюся дуже!
PS|62|3|(62-4) Доки будете ви нападати на людину? Усі хочете ви розтрощити її, немов мур той похилений, мов би паркан той валющий!
PS|62|4|(62-5) Вони тільки й думають, як би зіпхнути її з висоти, вони полюбили неправду: благословляють своїми устами, в своєму ж нутрі проклинають!... Села.
PS|62|5|(62-6) Тільки від Бога чекай у мовчанні, о душе моя, бо від Нього надія моя!
PS|62|6|(62-7) Тільки Він моя скеля й спасіння моє, Він твердиня моя, тому не захитаюсь!
PS|62|7|(62-8) У Бозі спасіння моє й моя слава, скеля сили моєї, моє пристановище в Бозі!
PS|62|8|(62-9) Мій народе, кожного часу надійтесь на Нього, серце своє перед Ним виливайте, Бог для нас пристановище! Села.
PS|62|9|(62-10) Справді, людські сини як та пара, сини й вищих мужів обмана: як узяти на вагу вони легші від пари всі разом!
PS|62|10|(62-11) Не надійтесь на утиск, і не пишайтесь грабунком; як багатство росте, не прикладайте свого серця до нього!
PS|62|11|(62-12) Один раз Бог сказав, а двічі я чув, що сила у Бога!
PS|62|12|(62-13) і в Тебе, о Господи, милість, бо відплачуєш кожному згідно з ділами його!
PS|63|1|Псалом Давидів, коли був він у пустині юдейській. (63-2) Боже Ти Бог мій, я шукаю від рання Тебе, душа моя прагне до Тебе, тужить тіло моє за Тобою в країні пустельній і вимученій без води...
PS|63|2|(63-3) Я так приглядався до Тебе в святині, щоб бачити силу Твою й Твою славу,
PS|63|3|(63-4) ліпша бо милість Твоя над життя, й мої уста Тебе прославляють!
PS|63|4|(63-5) Так я буду в житті своїм благословляти Тебе, ради Ймення Твого буду руки свої підіймати!
PS|63|5|(63-6) Насичується, ніби лоєм і товщем, душа моя, а уста мої хвалять губами співними.
PS|63|6|(63-7) Як згадаю Тебе на постелі своїй, розмишляю про Тебе в сторожах нічних:
PS|63|7|(63-8) що став Ти на поміч для мене, в тіні ж Твоїх крил я співатиму!
PS|63|8|(63-9) Пригорнулась до Тебе душа моя, правиця Твоя підпирає мене.
PS|63|9|(63-10) Вороги ж мою душу шукають для згуби, нехай западуться до споду землі,
PS|63|10|(63-11) нехай помордовані будуть мечем, бодай стали шакалам поживою!
PS|63|11|(63-12) А цар звеселиться у Бозі, буде хвалений кожен, хто йому присягає, будуть бо замкнені уста лжемовцям!
PS|64|1|Для дириґетна хору. Псалом Давидів. (64-2) Вислухай, Боже, мій голос, як скаржуся я, від страху ворожого душу мою хорони!
PS|64|2|(64-3) Заховай мене від потаємного збору злочинців, від крику свавільців,
PS|64|3|(64-4) які нагострили свого язика, як меча, натягнули стрілу свою словом гірким,
PS|64|4|(64-5) щоб таємно стріляти в невинного, вони нагло стрілятимуть в нього, і не будуть боятись!...
PS|64|5|(64-6) У злій справі зміцняють себе, змовляються пастки таємно розставити, кажуть: Хто буде їх бачити?
PS|64|6|(64-7) Вони кривди ховають... Загинемо, як задум їхній сповниться, бо нутро чоловіка та серце глибоке!
PS|64|7|(64-8) Але вчинить Бог, що стріла на них стрілить, і нагло поранені будуть,
PS|64|8|(64-9) і вчинить, що їхній язик допадеться до них, і будуть хитати головою усі, хто спогляне на них!...
PS|64|9|(64-10) і всі люди боятися будуть, і будуть розказувати про чин Бога, і діло Його зрозуміють!
PS|64|10|(64-11) і праведний Господом буде радіти, і буде вдаватись до Нього, і будуть похвалені всі простосерді!
PS|65|1|Для дириґетна хору. Псалом Давидів. Пісня. Уся земле, покликуйте Богові:
PS|65|2|Тобі, Боже, належиться слава в Сіоні, і Тобі має відданий бути обіт!
PS|65|3|Ти, що молитви вислухуєш, всяке тіло до Тебе приходить!
PS|65|4|Справи грішні зробились сильніші від нас, Ти наші гріхи пробачаєш!
PS|65|5|Блаженний, кого вибираєш Ти та наближаєш, в оселях Твоїх спочивати той буде! наситимось ми добром дому Твого, найсвятішим із храму Твого!
PS|65|6|Грізні речі Ти відповідаєш нам правдою, Боже, Спасителю наш, надіє всіх кінців землі та сущих далеко на морі,
PS|65|7|що гори ставиш Своєю силою, підперезаний міццю,
PS|65|8|що втихомирюєш гуркіт морів, їхніх хвиль та галас народів...
PS|65|9|і будуть боятись ознак Твоїх мешканці кінців землі. Ти розвеселяєш країну, де вихід поранку й де вечір.
PS|65|10|Ти відвідуєш землю та поїш її, Ти збагачуєш щедро її, повний води потік Божий, Ти збіжжя готуєш її, бо Ти так приготовив її!
PS|65|11|Ти ріллю її насичуєш вогкістю, вирівнюєш груддя її, розпускаєш дощами її, Ти благословляєш рослинність її!
PS|65|12|Ти добром Своїм рік вкороновуєш, і стежки Твої краплями товщу течуть!
PS|65|13|Пасовиська пустині спливаються краплями, і радістю підперезались узгір'я! (65-14) Луги зодягнулись отарами, а долини покрилися збіжжям, гукають вони та співають!
PS|66|1|Для дириґетна хору. Пісня. Псалом. Уся земле, покликуйте Богові,
PS|66|2|виспівуйте честь Його Йменню, честь для слави Його покладіть!
PS|66|3|Скажіть Богу: Які Твої вчинки грізні! Через силу велику Твою Твої вороги піддадуться Тобі,
PS|66|4|вся земля буде падати до ніг Твоїх, і співати Тобі буде, оспівувати Ймення Твоє! Села.
PS|66|5|ідіть і погляньте на Божі діла, Він грізний у ділах проти людських синів!
PS|66|6|Він на суходіл змінив море, й переходили річку ногою, там раділи ми в Ньому!
PS|66|7|Він царює навіки Своєю могутністю, очі Його між народами зорять, нехай не несуться відступники! Села.
PS|66|8|Благословляйте, народи, нашого Бога, і голос слави Його розголошуйте,
PS|66|9|що зберіг при житті нашу душу, і не дав нозі нашій спіткнутись,
PS|66|10|бо Ти, Боже, нас випробовував, Ти нас перетопив, як срібло перетоплюється...
PS|66|11|Ти нас до в'язниці впровадив, Ти пута поклав нам на стегна,
PS|66|12|Ти їздити дав був людині по головах наших, ми ввійшли до огню й до води, але на широкі місця Ти нас вивів!
PS|66|13|Увійду я до дому Твого з цілопаленнями, обіти свої Тобі виплачу ті,
PS|66|14|що їх вимовили мої губи й сказали були мої уста в тісноті моїй!
PS|66|15|Цілопалення ситих тельців піднесу Тобі з димом кадильним баранячим, приготую биків із козлами. Села.
PS|66|16|ідіть, і послухайте, всі богобійні, а я розкажу, що Він учинив для моєї душі:
PS|66|17|До Нього я кликав устами своїми, і хвали Йому під моїм язиком!
PS|66|18|Коли б беззаконня я бачив у серці своїм, то Господь не почув би мене,
PS|66|19|але Бог почув, і вислухав голос моєї молитви!
PS|66|20|Благословенний Бог, Який не відкинув моєї молитви й Свого милосердя від мене!
PS|67|1|Для дириґетна хору. На струнних знаряддях. Псалом. Пісня. (67-2) Нехай Бог помилує нас, і хай поблагословить, хай засяє над нами обличчям Своїм, Села,
PS|67|2|(67-3) щоб пізнати дорогу Твою на землі, посеред народів усіх спасіння Твоє!
PS|67|3|(67-4) Хай Тебе вихваляють народи, о Боже, хай славлять Тебе всі народи!
PS|67|4|(67-5) Нехай веселяться й співають племена, бо Ти правдою судиш народи й племена ведеш на землі! Села.
PS|67|5|(67-6) Хай Тебе вихваляють народи, о Боже, хай славлять Тебе всі народи!
PS|67|6|(67-7) Земля врожай свій дала, Бог поблагословив нас, наш Бог!
PS|67|7|(67-8) Нехай благословляє нас Бог, і всі кінці землі хай бояться Його!
PS|68|1|Для дириґетна хору. Псалом Давидів. Пісня. (68-2) Нехай воскресне Бог, і розпорошаться вороги Його, і нехай від лиця Його повтікають Його ненависники!
PS|68|2|(68-3) Як дим розвівається, так їх розвій, як топиться віск від огню, отак несправедливі загинуть перед Божим лицем!
PS|68|3|(68-4) А праведні будуть радіти, і будуть тішитися перед Богом, і веселитися в радості будуть!
PS|68|4|(68-5) Співайте Богові, виспівуйте Йменню Його, рівняйте дорогу Тому, Хто їде на хмарах, Господь Йому Ймення, та перед Ним веселіться!
PS|68|5|(68-6) Сиротам батько й вдовицям суддя, то Бог у святому мешканні Своїм!
PS|68|6|(68-7) Бог самітних уводить до дому, витягує в'язнів з кайданів, тільки відступники мешкати будуть у спаленій сонцем землі!
PS|68|7|(68-8) Боже, коли перед народом Своїм Ти виходив, коли йшов Ти пустинею, Села,
PS|68|8|(68-9) то тряслася земля, також капало небо було перед Богом, Сінай затремтів перед Богом, Богом ізраїля!
PS|68|9|(68-10) Дощ добродійний спускаєш Ти краплями, Боже, на спадок Свій перемучений міцно поставив його.
PS|68|10|(68-11) У ньому сиділо Твоє многолюддя, у Своїй доброті все готуєш Ти бідному, Боже!
PS|68|11|(68-12) Господь дає слово; провісниць велика многота:
PS|68|12|(68-13) Царі військ утікають, утікають, пані ж дому розділює здобич.
PS|68|13|(68-14) Коли ви спочиваєте між обійстями то крила голубки покриті сріблом, а пера її зеленкавістю золота.
PS|68|14|(68-15) Коли Всемогутній царів розпорошував в Краї, то сніг Ти спускав на Цалмоні.
PS|68|15|(68-16) Гора Божа Башанська гора, гора верхогір'я гора та Башанська.
PS|68|16|(68-17) Верхогір'я, чого заздрісно дивитеся на ту гору, що Бог зажадав на мешкання Своє, і Господь буде мешкати там завжди?
PS|68|17|(68-18) Колесниць Божих дві десятьтисячки, тисячі багатократні, Господь із Сінаю прибув до святині.
PS|68|18|(68-19) Ти піднявся був на висоту, полонених набрав, узяв дари ради людини, і відступники мешкати будуть у Господа Бога також.
PS|68|19|(68-20) Благословенний Господь, тягарі Він щоденно нам носить, Бог наше спасіння! Села.
PS|68|20|(68-21) Бог для нас Бог спасіння, і в Господа Владики виходи смерти!
PS|68|21|(68-22) Але розторощить Бог голову Своїх ворогів, маківку, вкриту волоссям, того, хто в гріхах своїх ходить!
PS|68|22|(68-23) Промовив Господь: Я спроваджу з Башану тебе, з глибин моря спроваджу,
PS|68|23|(68-24) щоб ти ногу свою мив у крові, щоб язик твоїх псів мав частину свою в ворогів!
PS|68|24|(68-25) Походи Твої, Боже, бачено, походи Бога мого у святині мого Царя:
PS|68|25|(68-26) Попереду йшли співаки, потому грачі, посеред дівчат, що бряжчали на бубнах:
PS|68|26|(68-27) Благословляйте на зборах Бога, Господа, ви, хто від джерел ізраїля!
PS|68|27|(68-28) Там Веніямин молодий, їхній володар, князі Юди, їхні полки, князі Завулона, князі Нефталима.
PS|68|28|(68-29) Твій Бог наказав тобі силу, будь силою, Боже, того, кого нам учинив!
PS|68|29|(68-30) із храму Твого на Єрусалимі царі привезуть Тобі дара.
PS|68|30|(68-31) Погрози звірині в очереті, череді волів разом з телятами людськими, понищ тих, хто кавалками срібла милується, розпорош ті народи, що воєн бажають!
PS|68|31|(68-32) Прийдуть з Єгипту посли, і руки свої Куш простягне до Бога.
PS|68|32|(68-33) Царства землі, співайте Богові, виспівуйте Господа, Села,
PS|68|33|(68-34) що їздить в відвічному небі небес. Ось Він загримить Своїм голосом, голосом сильним.
PS|68|34|(68-35) Визнайте Богові силу, величність Його над ізраїлем, а в хмарах потуга Його!
PS|68|35|(68-36) Бог грізний у святинях Своїх, Бог ізраїлів Він, що народові дає силу й міць, Бог благословенний!
PS|69|1|Для дириґетна хору. На спів: „Лелії". Давидів. (69-2) Спаси мене, Боже, бо води вже аж до душі підійшли!
PS|69|2|(69-3) Я загруз у глибокім багні, і нема на чім стати, ввійшов я до водних глибин, і мене залила течія!
PS|69|3|(69-4) Я змучився в крику своїм, висохло горло моє, очі мої затуманились від виглядання надії від Бога мого!...
PS|69|4|(69-5) Тих, хто мене без причини ненавидить, стало більш, як волосся на моїй голові, набралися сили мої вороги, що безвинно мене переслідують, чого не грабував, те вертаю!
PS|69|5|(69-6) Боже, Ти знаєш глупоту мою, а гріхи мої перед Тобою не сховані!
PS|69|6|(69-7) Нехай через мене не матимуть стиду оті, хто на Тебе надіється, Господи, Господи Саваоте; нехай через мене не матимуть сорому ті, хто шукає Тебе, Боже ізраїлів,
PS|69|7|(69-8) бо я ради Тебе зневагу ношу, ганьба покрила обличчя моє!...
PS|69|8|(69-9) Для братів своїх став я відчужений, і чужий для синів своєї матері,
PS|69|9|(69-10) бо ревність до дому Твойого з'їдає мене, і зневаги Твоїх зневажальників спадають на мене,
PS|69|10|(69-11) і постом я виплакав душу свою, а це сталось мені на зневагу...
PS|69|11|(69-12) За одежу надів я верету, і за приказку став я для них:
PS|69|12|(69-13) про мене балакають ті, хто в брамі сидить, і пісні тих, хто п'янке попиває...
PS|69|13|(69-14) А я молитва моя до Тебе, Господи, в часі Твоєї зичливости; в многоті милосердя Твойого подай мені відповідь про певність спасіння Твого,
PS|69|14|(69-15) визволь з болота мене, щоб я не втопився, щоб я урятований був від своїх ненависників та від глибокости вод!
PS|69|15|(69-16) Хай мене не заллє водяна течія, і хай глибінь мене не проковтне, і нехай своїх уст не замкне надо мною безодня!
PS|69|16|(69-17) Обізвися до мене, о Господи, в міру доброї ласки Своєї, в міру великости Свого милосердя звернися до мене,
PS|69|17|(69-18) і обличчя Свого не ховай від Свого раба, бо тісно мені, озвися ж небаром до мене,
PS|69|18|(69-19) наблизись до моєї душі, порятуй же її, ради моїх ворогів відкупи Ти мене!...
PS|69|19|(69-20) Ти знаєш наругу мою, і мій сором та ганьбу мою, перед Тобою всі мої вороги!
PS|69|20|(69-21) Моє серце зламала наруга, і невигойний мій сором: я чекав співчуття та немає його, і потішителів та не знайшов!
PS|69|21|(69-22) і жовчі поклали у мій хліб потішення, а в спразі моїй оцтом мене напували...
PS|69|22|(69-23) Бодай пасткою стала їм їхня трапеза, а їхні учти тенетами,
PS|69|23|(69-24) бодай їхні очі потемніли, щоб їм не бачити, а їхні клуби хай завжди хитаються!
PS|69|24|(69-25) Вилий на них Свою ревність, а полум'я гніву Твого нехай їх доганяє!
PS|69|25|(69-26) Нехай їхнє село опустошене буде, хай мешканця в їхніх наметах не буде!
PS|69|26|(69-27) Бо кого Ти був збив, вони ще переслідують, і побільшують муки раненим Тобою...
PS|69|27|(69-28) Додай же гріха на їхній гріх, щоб вони не ввійшли в справедливість Твою,
PS|69|28|(69-29) нехай скреслені будуть із книги життя, і хай не будуть записані з праведними!...
PS|69|29|(69-30) А я бідний та хворий, але, Боже, спасіння Твоє мене чинить могутнім,
PS|69|30|(69-31) і я піснею буду хвалити ім'я Боже, співом вдячним Його величатиму!
PS|69|31|(69-32) і буде для Господа краща вона від вола, від бика, що роги він має, що копита роздвоєні має.
PS|69|32|(69-33) Побачать слухняні, і будуть радіти, хто ж Бога шукає нехай оживе ваше серце,
PS|69|33|(69-34) бо до вбогих Господь прислухається, і в'язнями Своїми не гордує Він!
PS|69|34|(69-35) Нехай хвалять Його небеса та земля, море й усе, що в них рухається,
PS|69|35|(69-36) бо спасе Бог Сіона, і збудує для Юди міста, і замешкають там, і вспадкують його,
PS|69|36|(69-37) і нащадки рабів Його посядуть його, й ті, хто любить ім'я Його, житимуть в нім!
PS|70|1|Для дириґетна хору. Давидів. На пам'ятку. (70-2) Поквапся спасти мене, Боже, Господи, поспішися ж на поміч мені!
PS|70|2|(70-3) Нехай посоромлені будуть, і хай застидаються ті, хто шукає моєї душі, щоб схопити її! Нехай подадуться назад, і нехай посоромлені будуть усі, хто бажає для мене лихого!
PS|70|3|(70-4) Бодай повернулися з соромом ті, хто говорить на мене: Ага! Ага!
PS|70|4|(70-5) Нехай тішаться та веселяться Тобою усі, хто шукає Тебе, та хто любить спасіння Твоє, і хай завжди говорять: Хай буде великий Господь!
PS|70|5|(70-6) А я вбогий та бідний, поспіши ж Ти до Мене, о Боже: моя поміч і мій оборонець то Ти, Боже мій, не спізняйся!
PS|71|1|До Тебе вдаюся я, Господи, хай же не буду повік засоромлений!
PS|71|2|визволь мене через правду Свою, і звільни мене, нахили Своє ухо до мене, й спаси мене,
PS|71|3|стань для мене за скелю мешкальну, куди міг би я завжди ховатись! Ти наказав рятувати мене, бо Ти скеля моя та твердиня моя!
PS|71|4|Боже мій, визволь мене від руки беззаконного, від руки того, хто кривдить та гнобить мене,
PS|71|5|Ти бо, Владико, надія моя, Господи, Ти охорона моя від юнацького віку мого!
PS|71|6|На Тебе оперся я був від народження, від утроби моєї матері Ти охорона моя, в Тобі моя слава постійно!
PS|71|7|Я став багатьом, як дивовище, та Ти сильна моя охорона!
PS|71|8|Уста мої повні Твоєї хвали, увесь день Твоєї величности!
PS|71|9|Не кидай мене на час старости, коли зменшиться сила моя, не лиши Ти мене,
PS|71|10|бо мої вороги проти мене змовляються, а ті, що чатують на душу мою нараджаються разом,
PS|71|11|говорячи: Бог покинув його, доганяйте й хапайте його, бо нема, хто б його врятував!...
PS|71|12|Не віддалюйся, Боже, від мене, Боже мій поспішися ж на поміч мені!
PS|71|13|Нехай посоромляться, хай позникають усі, хто ненавидить душу мою, бодай зодяглися в наругу та в сором усі, хто прагне для мене лихого!
PS|71|14|А я буду постійно надіятись, і славу Твою над усе я помножу!
PS|71|15|Уста мої оповідатимуть правду Твою, про спасіння Твоє увесь день, бо числа їх не знаю,
PS|71|16|буду славити вчинки великі всевладного Господа, згадаю про правду Твою, єдино Твою!
PS|71|17|Боже, навчав Ти мене від юнацтва мого, і аж дотепер я звіщаю про чуда Твої.
PS|71|18|А Ти, Боже, не кидай мене аж до старости та сивини, поки я не звіщу про рамено Твоє поколінню, і кожному, хто тільки прийде про чини великі Твої!
PS|71|19|Бо Твоя справедливість, о Боже, сягає аж до високости, Боже, що речі великі вчинив, хто рівний Тобі?
PS|71|20|Ти мені показав був великі та люті нещастя, та знов Ти оживиш мене, і з безодень землі мене знову Ти витягнеш,
PS|71|21|Ти збільшиш величність мою, і знову потішиш мене!
PS|71|22|А я буду на арфі хвалити Тебе, Твою правду, мій Боже, із гуслами буду співати Тобі, Святий Ти ізраїлів!
PS|71|23|Нехай співом радіють уста мої, бо буду співати Тобі я та душа моя, яку Ти врятував!
PS|71|24|Шепоче про правду Твою мій язик цілий день, бо посоромлені, бо поганьблені всі, хто шукає лихого для мене!
PS|72|1|Соломонів. Боже, Свої суди цареві подай, а Свою справедливість для сина царевого,
PS|72|2|хай він правдою судить народа Твого, а вбогих Твоїх справедливістю!
PS|72|3|Нехай гори приносять народові мир, а пагірки правду.
PS|72|4|Він судитиме вбогих народу, помагатиме бідним, і тиснути буде гнобителя!
PS|72|5|Будуть боятися Тебе, поки сонця, і поки місяця, з роду до роду!
PS|72|6|Він зійде, як дощ на покіс, немов краплі, що зрошують землю!
PS|72|7|Праведний буде цвісти в його дні, а спокій великий аж поки світитиме місяць,
PS|72|8|і він запанує від моря до моря, і від Ріки аж до кінців землі!
PS|72|9|Мешканці пустинь на коліна попадають перед обличчям його, а його вороги будуть порох лизати...
PS|72|10|Царі Таршішу та островів дадуть дари, принесуть царі Шеви та Севи дарунки!
PS|72|11|і впадуть перед ним усі царі, і будуть служити йому всі народи,
PS|72|12|бо визволить він бідаря, що голосить, та вбогого, що немає собі допомоги!
PS|72|13|Він змилується над убогим та бідним, і спасе душу бідних,
PS|72|14|від кривди й насилля врятує їхню душу, їхня кров дорога буде в очах його!
PS|72|15|і буде він жити, і дасть йому з золота Шеви, і завжди молитися буде за нього, буде благословляти його кожен день!
PS|72|16|На землі буде збіжжя багато, на гірському верху зашумить, як Ливан, його плід, і народ зацвіте по містах, як трава на землі!
PS|72|17|Хай ім'я його буде навіки, хай росте, поки сонця, наймення його, нехай благословляються ним, будуть хвалити його всі народи!
PS|72|18|Благословен Господь Бог, Бог ізраїлів, єдиний, що чуда вчиняє,
PS|72|19|і благословенне навіки ім'я Його слави, і хай Його слава всю землю наповнить! Амінь і амінь!
PS|72|20|Скінчились молитви Давида, сина Єссея.
PS|73|1|Псалом Асафів. Поправді Бог добрий ізраїлеві, Бог для щиросердих!
PS|73|2|А я, мало не послизнулися ноги мої, мало не посковзнулися стопи мої,
PS|73|3|бо лихим я завидував, бачивши спокій безбожних,
PS|73|4|бо не мають страждання до смерти своєї, і здорове їхнє тіло,
PS|73|5|на людській роботі нема їх, і разом із іншими людьми не зазнають вони вдарів.
PS|73|6|Тому то пиха їхню шию оздоблює, зодягає їх шата насилля,
PS|73|7|вилазять їм очі від жиру, бажання їхнього серця збулися,
PS|73|8|сміються й злосливо говорять про утиск, говорять бундючно:
PS|73|9|свої уста до неба підносять, а їхній язик по землі походжає!...
PS|73|10|Тому то туди Його люди звертаються, і щедро беруть собі воду
PS|73|11|та й кажуть: Хіба Бог те знає, і чи має Всевишній відомість,
PS|73|12|як он ті безбожні й безпечні на світі збільшили багатство своє?
PS|73|13|Направду, надармо очистив я серце своє, і в невинності вимив руки свої,
PS|73|14|і ввесь день я побитий, і щоранку покараний...
PS|73|15|Коли б я сказав: Буду так говорить, як вони, то спроневірився б я поколінню синів Твоїх.
PS|73|16|і роздумував я, щоб пізнати оте, та трудне воно в очах моїх,
PS|73|17|аж прийшов я в Божу святиню, і кінець їхній побачив:
PS|73|18|направду, Ти їх на слизькому поставив, на спустошення кинув Ти їх!
PS|73|19|Як вони в одній хвилі спустошені, згинули, пощезали від страхів!
PS|73|20|Немов сном по обудженні, Господи, образом їхнім погордиш, мов сном по обудженні!
PS|73|21|Бо болить моє серце, і в нутрі моїм коле,
PS|73|22|а я немов бидло й не знаю, я перед Тобою худобою став!...
PS|73|23|Та я завжди з Тобою, Ти держиш мене за правицю,
PS|73|24|Ти Своєю порадою водиш мене, і потому до слави Ти візьмеш мене!
PS|73|25|Хто є мені на небесах, окрім Тебе? А я при Тобі на землі не бажаю нічого!
PS|73|26|Гине тіло моє й моє серце, та Бог скеля серця мого й моя доля навіки,
PS|73|27|бо погинуть ось ті, хто бокує від Тебе, понищиш Ти кожного, хто відступить від Тебе!
PS|73|28|А я, близькість Бога для мене добро, на Владику, на Господа свою певність складаю, щоб звіщати про всі Твої чини!
PS|74|1|Псалом навчальний, Асафів. Нащо, Боже, назавжди Ти нас опустив, чого розпалився Твій гнів на отару Твого пасовиська?
PS|74|2|Спогадай про громаду Свою, яку Ти віддавна набув, про племено спадку Свого, що його Ти був викупив, про ту гору Сіон, що на ній оселився,
PS|74|3|підійми ж Свої стопи до вічних руїн, бо ворог усе зруйнував у святині!...
PS|74|4|Ревіли Твої вороги у святині Твоїй, умістили знаки за ознаки свої,
PS|74|5|виглядало то так, якби хто догори підіймав був сокири в гущавині дерева...
PS|74|6|А тепер її різьби ураз розбивають вони молотком та сокирами,
PS|74|7|Святиню Твою на огонь віддали, оселю Твого Ймення аж дощенту збезчестили...
PS|74|8|Сказали вони в своїм серці: Зруйнуймо їх разом! і спалили в краю всі місця Божих зборів...
PS|74|9|Наших ознак ми не бачимо, нема вже пророка, і між нами немає такого, хто знає, аж доки це буде...
PS|74|10|Аж доки, о Боже, гнобитель знущатися буде, зневажатиме ворог навіки ім'я Твоє?
PS|74|11|Для чого притримуєш руку Свою та правицю Свою? З середини лоня Свого їх понищ!
PS|74|12|А Ти, Боже, віддавна мій Цар, Ти чиниш спасіння посеред землі!
PS|74|13|Розділив Ти був море Своєю потугою, побив голови зміям на водах,
PS|74|14|Ти левіятанові голову був поторощив, його Ти віддав був на їжу народові пустині,
PS|74|15|Ти був розділив джерело та потік, Ти висушив ріки великі!
PS|74|16|Твій день, а також Твоя ніч, приготовив Ти світло та сонце,
PS|74|17|всі границі землі Ти поставив, Ти літо та зиму створив!
PS|74|18|Пам'ятай же про це: ворог знущається з Господа, а народ нерозумний зневажує Ймення Твоє!
PS|74|19|Не віддай звірині душі Своєї горлиці, живої Твоїх бідарів не забудь же назавжди!
PS|74|20|Споглянь же на Свій заповіт, бо темноти землі повні мешкань насилля!
PS|74|21|Нехай не відходить пригноблений посоромленим, бідний та вбогий нехай прославляють імення Твоє!
PS|74|22|Встань же, о Боже, судися за справу Свою, пам'ятай про щоденну наругу Свою від безумного!
PS|74|23|Не забудь же про вереск Своїх ворогів, про галас бунтівників проти Тебе, що завжди зростає!
PS|75|1|Для дириґетна хору. „Не вигуби!" Псалом Асафів. Пісня. (75-2) Прославляємо, Боже, Тебе, прославляєм, бо близьке Твоє Ймення! Оповідають про чуда Твої.
PS|75|2|(75-3) Коли прийде година означена, то Я буду судити справедливо.
PS|75|3|(75-4) Розтопилась земля, і всі її мешканці, та стовпи її зміцнюю Я. Села.
PS|75|4|(75-5) Я сказав до лихих: Не шалійте, а безбожним: Не підіймайте ви рога!
PS|75|5|(75-6) Не підіймайте ви рога свого догори, не говоріть твердошийно,
PS|75|6|(75-7) бо не від сходу, і не від заходу, і не від пустині надійде повищення,
PS|75|7|(75-8) але судить Бог: того Він понижує, а того повищує,
PS|75|8|(75-9) бо чаша в Господній руці, а шумливе вино повне мішаного, і наливає Він з нього, усі ж беззаконні землі виссуть та вип'ють лиш дріжджі її!
PS|75|9|(75-10) А я буду звіщати навіки, співатиму Богові Якова,
PS|75|10|(75-11) відрубаю всі роги безбожних, роги праведного піднесуться!
PS|76|1|Для дириґетна хору. На неґінах. Псалом Асафів. Пісня. (76-2) Бог знаний у Юді, Його Ймення велике в ізраїлі!
PS|76|2|(76-3) У Салимі намет Його, а мешкання Його на Сіоні,
PS|76|3|(76-4) Він там поламав стріли луку, щита та меча, та війну! Села.
PS|76|4|(76-5) Ти осяйний, потужніший за гори відвічні.
PS|76|5|(76-6) Обдерто людей сильносердих, задрімали вони своїм сном, і не знайшли своїх рук усі мужі військові...
PS|76|6|(76-7) Від сваріння Твого, Боже Яковів, оглушується колесниця та кінь:
PS|76|7|(76-8) Ти Ти грізний, і хто перед обличчям Твоїм устоїть часу гніву Твого?...
PS|76|8|(76-9) Як звіщаєш Ти суд із небес, то боїться й стихає земля,
PS|76|9|(76-10) як встає Бог на суд, щоб спасти всіх покірних землі! Села.
PS|76|10|(76-11) Бо й гнів людський Тебе вихваляє, решту ж гніву Ти поясом в'яжеш.
PS|76|11|(76-12) Присягайте й виконуйте Господу, Богові вашому, усі, хто Його оточає, хай приносять дарунка Грізному:
PS|76|12|(76-13) Він духа вельмож впокоряє, страшний Він для земних царів!
PS|77|1|Для дириґетна хору. Псалом Асафів. (77-2) Мій голос до Бога, й я кликати буду, мій голос до Бога, й почує мене!
PS|77|2|(77-3) В день недолі моєї шукаю я Господа, до Нього рука моя витягнена вночі й не зомліє, не хоче душа моя бути потішена:
PS|77|3|(77-4) згадаю про Бога й зідхаю, розважаю й мій дух омліває! Села.
PS|77|4|(77-5) Ти держиш повіки очей моїх, я побитий і не говорю...
PS|77|5|(77-6) Пригадую я про дні давні, про роки відвічні,
PS|77|6|(77-7) свою пісню вночі я пригадую, говорю з своїм серцем, а мій дух розважає:
PS|77|7|(77-8) Чи навіки покине Господь, і вже більш не вподобає?
PS|77|8|(77-9) Чи навіки спинилася милість Його? Чи скінчилося слово Його в рід і рід?
PS|77|9|(77-10) Чи Бог милувати позабув? Чи гнівом замкнув Він Своє милосердя? Села.
PS|77|10|(77-11) і промовив був я: То страждання моє переміна правиці Всевишнього.
PS|77|11|(77-12) Пригадаю я вчинки Господні, як чудо Твоє я згадаю віддавна,
PS|77|12|(77-13) і буду я думати про кожен Твій чин, і про вчинки Твої оповім!
PS|77|13|(77-14) Боже, святая дорога Твоя, котрий бог великий, як Бог наш?
PS|77|14|(77-15) Ти Той Бог, що чуда вчиняє, Ти виявив силу Свою між народами,
PS|77|15|(77-16) Ти визволив люд Свій раменом, синів Якова й Йосипа! Села.
PS|77|16|(77-17) Тебе бачили води, о Боже, Тебе бачили води й тремтіли, затряслися й безодні.
PS|77|17|(77-18) Лилася струмком вода з хмар, тучі видали грім, також там і сям Твої стріли літали.
PS|77|18|(77-19) Гуркіт грому Твого на небесному колі, й блискавки освітили вселенну, тремтіла й тряслася земля!
PS|77|19|(77-20) Через море дорога Твоя, а стежка Твоя через води великі, і не видно було Твоїх стіп.
PS|77|20|(77-21) Ти провадив народ Свій, немов ту отару, рукою Мойсея та Аарона.
PS|78|1|Пісня навчальна Асафова. Послухай, мій люду, науки моєї, нахиліть своє ухо до слів моїх уст,
PS|78|2|нехай я відкрию уста свої приказкою, нехай стародавні прислів'я я висловлю!
PS|78|3|Що ми чули й пізнали, і що розповідали батьки наші нам,
PS|78|4|того не сховаємо від їхніх синів, будемо розповідати про славу Господню аж до покоління останнього, і про силу Його та про чуда Його, які Він учинив!
PS|78|5|Він поставив засвідчення в Якові, а Закона поклав ув ізраїлі, про які наказав був Він нашим батькам завідомити про них синів їхніх,
PS|78|6|щоб знало про це покоління майбутнє, сини, що народжені будуть, устануть і будуть розповідати своїм дітям.
PS|78|7|і положать на Бога надію свою, і не забудуть діл Божих, Його ж заповіді берегтимуть.
PS|78|8|і не стануть вони, немов їхні батьки, поколінням непокірливим та бунтівничим, поколінням, що серця свого не поставило міцно, і що дух його Богу невірний.
PS|78|9|Сини Єфрема, озброєні лучники, повернулися взад у день бою:
PS|78|10|вони не берегли заповіту Божого, а ходити в Законі Його відреклися,
PS|78|11|і забули вони Його чини та чуда Його, які їм показав.
PS|78|12|Він чудо вчинив був для їхніх батьків ув єгипетськім краї, на полі Цоанськім:
PS|78|13|Він море розсік, і їх перепровадив, а воду поставив, як вал;
PS|78|14|і провадив їх хмарою вдень, а сяйвом огню цілу ніч;
PS|78|15|на пустині Він скелі розсік, і щедро усіх напоїв, як з безодні.
PS|78|16|Він витягнув із скелі потоки, і води текли, немов ріки.
PS|78|17|Та грішили вони проти Нього ще далі, і в пустині гнівили Всевишнього,
PS|78|18|і Бога вони випробовували в своїм серці, для душ своїх їжі бажаючи.
PS|78|19|і вони говорили насупроти Бога й казали: Чи Бог зможе в пустині трапезу зготовити?
PS|78|20|Тож ударив у скелю і води линули, і полилися потоки! Чи Він зможе також дати хліба? Чи Він наготує м'ясива народові Своєму?
PS|78|21|Тому то почув це Господь та й розгнівався, і огонь запалав проти Якова, і проти ізраїля теж знявся гнів,
PS|78|22|бо не вірували вони в Бога, і на спасіння Його не надіялись.
PS|78|23|А Він хмарам згори наказав, і відчинив двері неба,
PS|78|24|і спустив, немов дощ, на них манну для їжі, і збіжжя небесне їм дав:
PS|78|25|Хліб ангольський їла людина, Він послав їм поживи до ситости!
PS|78|26|Крім цього, Він східнього вітра порушив на небі, і міццю Своєю привів полудневого вітра,
PS|78|27|і дощем на них м'ясо пустив, немов порох, а птаство крилате, як морський пісок,
PS|78|28|і спустив його серед табору його, коло наметів його.
PS|78|29|і їли вони та й наситились дуже, Він їм їхнє бажання приніс!
PS|78|30|Та ще не вдовольнили жадання свого, ще їхня їжа була в їхніх устах,
PS|78|31|а гнів Божий піднявся на них, та й побив їхніх ситих, і вибранців ізраїлевих повалив...
PS|78|32|Проте ще й далі грішили вони та не вірили в чуда Його,
PS|78|33|і Він докінчив у марноті їхні дні, а їхні літа у страху.
PS|78|34|Як Він їх побивав, то бажали Його, і верталися, й Бога шукали,
PS|78|35|і пригадували, що Бог їхня скеля, і Бог Всевишній то їхній Викупитель.
PS|78|36|і своїми устами влещували Його, а своїм язиком лжу сплітали Йому,
PS|78|37|бо їхнє серце не міцно стояло при Нім, і не були вони вірні в Його заповіті...
PS|78|38|Та він, Милосердний, гріх прощав і їх не губив, і часто відвертав Свій гнів, і не будив усю Свою лютість,
PS|78|39|і Він пам'ятав, що вони тільки тіло, вітер, який переходить і не повертається!
PS|78|40|Скільки вони прогнівляли Його на пустині, зневажали Його на степу!
PS|78|41|і все знову та знов випробовували вони Бога, і зневажали Святого ізраїлевого,
PS|78|42|вони не пам'ятали руки Його з дня, як Він вибавив їх із недолі,
PS|78|43|як в Єгипті чинив Він знамена Свої, а на полі Цоанському чуда Свої,
PS|78|44|і в кров обернув річки їхні та їхні потоки, щоб вони не пили...
PS|78|45|Він послав був на них рої мух, і їх жерли вони, і жаб і вони їх губили.
PS|78|46|А врожай їхній віддав був Він гусені, а їхню працю сарані.
PS|78|47|Виноград їхній Він градом побив, а приморозком їхні шовковиці.
PS|78|48|і Він градові віддав їхній скот, а блискавкам череди їхні.
PS|78|49|Він послав був на них Свій гнів запальний, і лютість, й обурення, й утиск, наслання злих анголів.
PS|78|50|Він дорогу зрівняв був для гніву Свого, їхні душі не стримав від смерти, життя ж їхнє віддав моровиці.
PS|78|51|і побив Він усіх перворідних в Єгипті, первістків сили в наметах Хамових.
PS|78|52|і повів Він, немов ту отару, народ Свій, і їх попровадив, як стадо, в пустині.
PS|78|53|і провадив безпечно Він їх, і вони не боялись, а море накрило було ворогів їхніх.
PS|78|54|і Він їх привів до границі святині Своєї, до тієї гори, що правиця Його набула.
PS|78|55|і народи Він повиганяв перед їхнім обличчям, і кинув для них жеребка про спадок, і в їхніх наметах племена ізраїлеві оселив.
PS|78|56|Та й далі вони випробовували та гнівили Всевишнього Бога, і Його постанов не додержували,
PS|78|57|і відступали та зраджували, немов їхні батьки відвернулись, як обманливий лук.
PS|78|58|і жертівниками своїми гнівили Його, і дрочили Його своїми фіґурами.
PS|78|59|Бог почув усе це і розгнівався, і сильно обридивсь ізраїлем,
PS|78|60|і покинув оселю в Шіло, скинію ту, що вмістив був посеред людей,
PS|78|61|і віддав до неволі Він силу Свою, а величність Свою в руку ворога...
PS|78|62|і віддав для меча Свій народ, і розгнівався був на спадщину Свою:
PS|78|63|його юнаків огонь пожирав, а дівчатам його не співали весільних пісень,
PS|78|64|його священики від меча полягли, і не плакали вдови його.
PS|78|65|Та небавом збудився Господь, немов зо сну, як той велет, що ніби вином був підкошений,
PS|78|66|і вдарив Своїх ворогів по озадку, вічну ганьбу їм дав!
PS|78|67|Та Він погордив намет Йосипів, і племена Єфремового не обрав,
PS|78|68|а вибрав Собі плем'я Юдине, гору Сіон, що її полюбив!
PS|78|69|і святиню Свою збудував Він, як місце високе, як землю, що навіки її вґрунтував.
PS|78|70|і вибрав Давида, Свого раба, і від кошар його взяв,
PS|78|71|від кітних овечок його Він привів, щоб Якова пас він, народа Свого, та ізраїля, спадок Свій,
PS|78|72|і він пас їх у щирості серця свого, і провадив їх мудрістю рук своїх!
PS|79|1|Псалом Асафів. Боже, погани ввійшли до спадку Твого, занечистили храм Твій святий, Єрусалим на руїни змінили!
PS|79|2|Рабів Твоїх трупи вони віддали на поживу для птаства небесного, тіло Твоїх богобійних звірині земній...
PS|79|3|Вони розливали їхню кров, немов воду, в околицях Єрусалиму, і не було погребальників!...
PS|79|4|Ми стали за ганьбу для наших сусідів, за наругу та посміх для наших околиць...
PS|79|5|Аж доки, о Господи, гніватись будеш назавжди, доки буде палати Твій гнів, як огонь?
PS|79|6|Вилий Свій гнів на людей, що Тебе не пізнали, і на царства, що Ймення Твого не кличуть,
PS|79|7|бо вони з'їли Якова, а мешкання його опустошили!
PS|79|8|Не пам'ятай гріхів предківських нам, нехай попередить нас скоро Твоє милосердя, бо ми зовсім ослабли!...
PS|79|9|Поможи нам, Боже нашого спасіння, ради слави Ймення Твого, і збережи нас, і прости наші гріхи ради Ймення Свого!
PS|79|10|Чого будуть казати погани: Де їхній Бог? Нехай в наших очах між народами стане відомою помста за пролиту кров Твоїх рабів,
PS|79|11|нехай перед лице Твоє дійде стогін в'язня! За великістю сили рамена Твого збережи на смерть прирокованих!
PS|79|12|А нашим сусідам верни семикратно на лоно їхнє їхню наругу, якою Тебе зневажали, о Господи!
PS|79|13|А ми, Твій народ і отара Твого пасовиська, будем дякувати Тобі вічно, будем оповідати про славу Твою з роду в рід!
PS|80|1|Для дириґетна хору. На „Лілеї". Свідоцтво. Псалом Асафів. (80-2) Пастирю ізраїлів, послухай же, Ти, що провадиш, немов ту отару, Йосипа, що на Херувимах сидиш, появися
PS|80|2|(80-3) перед обличчям Єфрема, і Веніямина, і Манасії! Пробуди Свою силу, і прийди, щоб спасти нас!
PS|80|3|(80-4) Боже, приверни нас, і хай засяє обличчя Твоє, й ми спасемось!
PS|80|4|(80-5) Господи, Боже Саваоте, доки будеш Ти гніватися на молитву народу Свого?
PS|80|5|(80-6) Ти вчинив був, що їли вони слізний хліб, і їх напоїв Ти сльозами великої міри...
PS|80|6|(80-7) Ти нас положив суперечкою нашим сусідам, і насміхаються з нас неприятелі наші...
PS|80|7|(80-8) Боже Саваоте, приверни нас, і хай засяє обличчя Твоє, й ми спасемось!
PS|80|8|(80-9) Виноградину Ти переніс із Єгипту, Ти вигнав народи й її посадив,
PS|80|9|(80-10) Ти випорожнив перед нею, і закоренила коріння своє, й переповнила край,
PS|80|10|(80-11) гори покрилися тінню її, а віття її Божі кедри,
PS|80|11|(80-12) аж до моря галузки її посилаєш, а парості її до ріки!
PS|80|12|(80-13) Але нащо вилім зробив Ти в горожі її, і всі нищать її, хто проходить дорогою?
PS|80|13|(80-14) Гризе її вепр лісовий, і звірина польова виїдає її!
PS|80|14|(80-15) Боже Саваоте, вернися ж, споглянь із небес і побач, і відвідай цього виноградника,
PS|80|15|(80-16) і охорони його, якого насадила правиця Твоя, і галузку, яку Ти для Себе зміцнив!
PS|80|16|(80-17) В огні виноградина спалена, відтята, гинуть від свару обличчя Твого,
PS|80|17|(80-18) нехай буде рука Твоя над мужем Твоєї правиці, на людському сині, якого зміцнив Ти Собі!
PS|80|18|(80-19) А ми не відступимо від Тебе, Ти нас оживиш, і ми будемо ім'я Твоє кликати!
PS|80|19|(80-20) Господи, Боже Саваоте, приверни нас, і хай засяє обличчя Твоє, й ми спасемось!
PS|81|1|Для дириґетна хору. На ґітійськім знарядді. Асафів. (81-2) Співайте Богові, нашій твердині, покликуйте Богові Якова,
PS|81|2|(81-3) заспівайте пісню, і заграйте на бубні, на цитрі приємній із гуслами,
PS|81|3|(81-4) засурміть у сурму в новомісяччя, на повні в день нашого свята,
PS|81|4|(81-5) бо це право ізраїлеві, Закон Бога Якова!
PS|81|5|(81-6) На свідчення в Йосипі Він учинив його, як пішов був на землю єгипетську. Почув був там мову, якої не знав:
PS|81|6|(81-7) Рамена його Я звільнив з тягару, від коша його руки звільнились.
PS|81|7|(81-8) Ти був кликав у недолі, й я видер тебе, Я відповідаю тобі в укритті громовім, Я випробував був тебе над водою Мериви. Села.
PS|81|8|(81-9) Слухай же ти, Мій народе, і хай Я засвідчу тобі, о ізраїлю, коли б ти послухав Мене:
PS|81|9|(81-10) нехай бога чужого у тебе не буде, і не кланяйся богу сторонньому!
PS|81|10|(81-11) Я Господь, Бог твій, що з краю єгипетського тебе вивів, відчини свої уста і Я їх наповню!
PS|81|11|(81-12) Але Мій народ не послухався був Мого голосу, не згодився зо Мною ізраїль,
PS|81|12|(81-13) і Я їх пустив ради впертости їхнього серця, нехай вони йдуть за своїми порадами!
PS|81|13|(81-14) Коли б Мій народ був послухав Мене, коли б був ізраїль ходив по дорогах Моїх,
PS|81|14|(81-15) ще мало і Я похилив би був їхніх ворогів, і руку Свою повернув би був Я на противників їхніх!
PS|81|15|(81-16) Ненависники Господа йому б покорились, і був би навіки їхній час,
PS|81|16|(81-17) і Я жиром пшениці його годував би, і медом із скелі тебе б насищав!
PS|82|1|Псалом Асафів. Бог на Божім зібранні стоїть, серед богів Він судить:
PS|82|2|Аж доки ви будете несправедливо судити, і доки будете ви підіймати обличчя безбожних? Села.
PS|82|3|Розсудіте нужденного та сироту, оправдайте убогого та бідаря,
PS|82|4|порятуйте нужденного та бідака, збережіть з руки несправедливих!
PS|82|5|Не пізнали та не зрозуміли, у темряві ходять вони... Всі основи землі захитались...
PS|82|6|Я сказав був: Ви боги, і сини ви Всевишнього всі,
PS|82|7|та однак повмираєте ви, як людина, і попадаєте, як кожен із вельмож.
PS|82|8|Устань же, о Боже, та землю суди, бо у владі Твоїй всі народи!
PS|83|1|Пісня. Псалом Асафів. (83-2) Боже, не будь мовчазним, не мовчи, і не будь Ти спокійним, о Боже,
PS|83|2|(83-3) бо ось зашуміли Твої вороги, а Твої ненависники голови попідіймали!
PS|83|3|(83-4) Вони проти народу Твого хитрий задум видумують, і нараджуються проти тих, кого Ти бережеш!
PS|83|4|(83-5) Вони кажуть: Ходіть но, та знищимо їх з-між народів, і згадуватись більш не буде імення ізраїля!
PS|83|5|(83-6) Бо вони однодушно нарадилися, проти Тебе умови складають,
PS|83|6|(83-7) намети Едома й ізмаїльтян, Моав та агаряни,
PS|83|7|(83-8) Ґевал і Аммон, і Амалик, Филистея з мешканцями Тиру.
PS|83|8|(83-9) і Ашшур поєднався був з ними, вони синам Лотовим стали раменом. Села.
PS|83|9|(83-10) Зроби їм, як Мідіянові, як Сісері, як Явінові в долині Кішон,
PS|83|10|(83-11) при Ен-Дорі вони були знищені, стали погноєм землі!
PS|83|11|(83-12) Поклади їх та їхніх вельмож, як Орева, й як Зеева, й як Зеваха, й як Цалмунну, усіх їхніх князів,
PS|83|12|(83-13) що казали були: Візьмімо на спадок для себе помешкання Боже!
PS|83|13|(83-14) Боже мій, бодай стали вони, немов порох у вихрі, як солома на вітрі!
PS|83|14|(83-15) Як огонь палить ліс, й як запалює полум'я гори,
PS|83|15|(83-16) так Ти їх пожени Своїм вихром, і настраш Своєю бурею!
PS|83|16|(83-17) Наповни обличчя їхнє соромом, і хай шукають вони Твоє Ймення, о Господи!
PS|83|17|(83-18) Нехай будуть вони засоромлені, й завжди хай будуть настрашені, і хай застидаються, й хай вони згинуть!
PS|83|18|(83-19) і нехай вони знають, що Ти, Твоє Ймення Господь, Сам Ти, Всевишній, на цілій землі!
PS|84|1|Для дириґетна хору. На ґітійськомім знарядді. Синів Кореєвих. Псалом. (84-2) Які любі оселі Твої, Господи Саваоте!
PS|84|2|(84-3) Затужена та омліває душа моя за подвір'ями Господа, моє серце та тіло моє линуть до Бога Живого!
PS|84|3|(84-4) і пташка знаходить домівку, і кубло собі ластівка, де кладе пташенята свої, при жертівниках Твоїх, Господи Саваоте, Царю мій і Боже мій!
PS|84|4|(84-5) Блаженні, хто мешкає в домі Твоїм, вони будуть повіки хвалити Тебе! Села.
PS|84|5|(84-6) Блаженна людина, що в Тобі має силу свою, блаженні, що в їхньому серці дороги до Тебе,
PS|84|6|(84-7) ті, що через долину Плачу переходять, чинять її джерелом, і дощ ранній дає благословення!
PS|84|7|(84-8) Вони ходять від сили до сили, і показуються перед Богом у Сіоні.
PS|84|8|(84-9) Господи, Боже Саваоте, послухай молитву мою, почуй, Боже Яковів! Села.
PS|84|9|(84-10) Щите наш, поглянь же, о Боже, і придивись до обличчя Свого помазанця!
PS|84|10|(84-11) Ліпший бо день на подвір'ях Твоїх, аніж тисяча в іншому місці, я б вибрав сидіти при порозі дому Бога мого, аніж жити в наметах безбожности!
PS|84|11|(84-12) Бо сонце та щит Господь, Бог! Господь дає милість та славу, добра не відмовляє усім, хто в невинності ходить.
PS|84|12|(84-13) Господи Саваоте, блаженна людина, що на Тебе надіється!
PS|85|1|Для дириґетна хору. Синів Кореєвих. Псалом. (85-2) Ти вподобав Собі Свою землю, о Господи, долю Якову Ти повернув,
PS|85|2|(85-3) Ти провину народу Свого простив, увесь гріх їхній покрив! Села.
PS|85|3|(85-4) Ти гнів Свій увесь занехав, Ти повстримав Свій гнів від палючої лютости!
PS|85|4|(85-5) Поверни нас до Себе, о Боже нашого спасіння, а Свій гнів проти нас поторощ!
PS|85|5|(85-6) Чи навіки Ти гніватись будеш на нас, і протягнеш Свій гнів з роду в рід?
PS|85|6|(85-7) Отож, Ти оживиш нас знову, і буде радіти народ Твій Тобою!
PS|85|7|(85-8) Покажи нам, о Господи, милість Свою, і подай нам спасіння Своє,
PS|85|8|(85-9) нехай я почую, що каже Бог, Господь, бо говорить Він Мир! народові Своєму й Своїм святим, і нехай до безумства вони не вертаються!
PS|85|9|(85-10) Справді, спасіння Його близьке тим, хто боїться Його, щоб слава Його була в нашій землі.
PS|85|10|(85-11) Милість та правда спіткаються, справедливість та мир поцілуються,
PS|85|11|(85-12) правда з землі виростає, а справедливість із небес визирає.
PS|85|12|(85-13) і Господь дасть добро, а земля наша дасть урожай свій.
PS|85|13|(85-14) Справедливість ходитиме перед обличчям Його, і кроки свої на дорогу поставить.
PS|86|1|Молитва Давидова. Нахили, Господи, ухо Своє і вислухай мене, бо я бідний та вбогий!
PS|86|2|Бережи мою душу, бо я богобійний, спаси Ти, мій Боже, Свого раба, що на Тебе надію кладе!
PS|86|3|Змилосердься до мене, о Господи, бо я кличу до Тебе ввесь день,
PS|86|4|потіш душу Свого раба, бо до Тебе підношу я, Господи, душу мою,
PS|86|5|бо Ти, Господи, добрий і вибачливий, і многомилостивий для всіх, хто кличе до Тебе!
PS|86|6|Почуй же, о Господи, молитву мою, і вислухай голос благання мого,
PS|86|7|в день недолі своєї я кличу до Тебе, бо Ти обізвешся до мене!
PS|86|8|Нема, Господи, поміж богами такого, як Ти, і чинів нема, як чини Твої!
PS|86|9|Всі народи, яких Ти створив, поприходять і попадають перед лицем Твоїм, Господи, та ім'я Твоє славити будуть,
PS|86|10|великий бо Ти, та чуда вчиняєш, Ти Бог єдиний!
PS|86|11|Дорогу Свою покажи мені, Господи, і я буду ходити у правді Твоїй, приєднай моє серце боятися Ймення Твого!
PS|86|12|Я буду всім серцем своїм вихваляти Тебе, Господи, Боже Ти мій, і славити буду повіки ім'я Твоє,
PS|86|13|велика бо милість Твоя надо мною, і вирвав Ти душу мою від шеолу глибокого!
PS|86|14|Боже, злочинці повстали на мене, а натовп гнобителів прагне моєї душі, і перед собою не ставлять Тебе...
PS|86|15|А Ти, Господи, Бог щедрий і милосердний, довготерпеливий і многомилостивий, і справедливий,
PS|86|16|зглянься на мене, й помилуй мене, подай же Своєму рабові Свою силу, і спаси сина Своєї невільниці!
PS|86|17|Учини мені знака на добре, і нехай це побачать мої ненависники, і хай засоромлені будуть, бо Ти, Господи, мені допоміг та мене звеселив!
PS|87|1|Синів Кореєвих. Псалом. Пісня. Основа його на горах святих,
PS|87|2|Господь любить брами Сіону понад усі селища Яковові.
PS|87|3|Славне розповідають про тебе, місто Боже! Села.
PS|87|4|Тим, хто знає мене, нагадаю про Рагав та про Вавилон; ось Филистея та Тир з Кушем кажуть: Отой народився був там.
PS|87|5|і про Сіон говоритимуть: Той і той народився був у ньому, й Сам Всевишній зміцняє його!
PS|87|6|Господь буде лічити у книзі народів: Оцей народився був там! Села.
PS|87|7|і співають у танку вони: У Тобі всі джерела мої!
PS|88|1|Пісня. Псалом. Синів Кореєвих. Для дириґетна хору. На „Махалат лефннот". Пісня навчальна Гемана езрахеяннина. (88-2) Господи, Боже спасіння мого, вдень я кличу й вночі я перед Тобою:
PS|88|2|(88-3) хай молитва моя дійде перед обличчя Твоє, нахили Своє ухо до зойку мого,
PS|88|3|(88-4) душа бо моя наситилась нещастями, а життя моє зблизилося до шеолу!
PS|88|4|(88-5) Я до тих прирахований став, що в могилу відходять, я став, немов муж той безсилий...
PS|88|5|(88-6) Я кинений серед померлих, немов оті трупи, що в гробі лежать, що про них Ти не згадуєш більш, і потяті вони від Твоєї руки...
PS|88|6|(88-7) Умістив Ти мене в глибочезну могилу, до пітьми в глибинах.
PS|88|7|(88-8) На мене лягла Твоя лють, і Ти всіма Своїми ламаннями мучив мене... Села.
PS|88|8|(88-9) Віддалив Ти від мене знайомих моїх, учинив Ти мене за огиду для них... Я замкнений і не виходжу,
PS|88|9|(88-10) стемніло з біди моє око... Я кожного дня Тебе кличу, о Господи, простягаю до Тебе руки свої!...
PS|88|10|(88-11) Чи Ти чудо вчиниш померлим? Чи трупи встануть і будуть хвалити Тебе? Села.
PS|88|11|(88-12) Хіба милість Твоя буде в гробі звіщатись, а вірність Твоя в аввадоні?
PS|88|12|(88-13) Чи познається в темряві чудо Твоє, а в краю забуття справедливість Твоя?
PS|88|13|(88-14) Та я кличу до Тебе, о Господи, і вранці молитва моя Тебе випереджує...
PS|88|14|(88-15) Для чого, о Господи, кидаєш душу мою, ховаєш від мене обличчя Своє?
PS|88|15|(88-16) Нужденний я та помираю відмалку, переношу страхіття Твої, я ослаблений став...
PS|88|16|(88-17) Перейшли надо мною Твої пересердя, страхіття Твої зруйнували мене,
PS|88|17|(88-18) вони оточають мене, як вода, увесь день, вони разом мене облягають...
PS|88|18|(88-19) друга й приятеля віддалив Ти від мене, знайомі мої як та темрява!...
PS|89|1|Навчальна пісня Етана езрахеяннина. (89-2) Про милості Господа буду співати повіки, я буду звіщати устами своїми про вірність Твою з роду в рід!
PS|89|2|(89-3) Бо я був сказав: Буде навіки збудована милість, а небо Ти вірність Свою встановляєш на нім.
PS|89|3|(89-4) Я склав заповіта з вибранцем Своїм, присягнув Я Давидові, Моєму рабові:
PS|89|4|(89-5) Встановлю Я навіки насіння твоє, а твій трон Я збудую на вічні віки! Села.
PS|89|5|(89-6) і небо хвалитиме, Господи, чудо Твоє, також вірність Твою на зібранні святих,
PS|89|6|(89-7) бо хто в небі подібний до Господа? Хто подібний до Господа серед Божих синів?
PS|89|7|(89-8) Бог дуже страшний у зібранні святих, і грізний Він на ціле довкілля Своє!
PS|89|8|(89-9) Господи, Боже Саваоте, хто сильний, як Ти, Господи? А вірність Твоя на довкіллі Твоїм!
PS|89|9|(89-10) Ти пануєш над силою моря, коли підіймаються хвилі, Ти їх втихомирюєш.
PS|89|10|(89-11) Ти стиснув Рагава, як трупа, і сильним раменом Своїм розпорошив Своїх ворогів.
PS|89|11|(89-12) Твої небеса, Твоя теж земля, вселенна і все, що на ній, Ти їх заложив!
PS|89|12|(89-13) Північ та південє Ти їх створив, Фавор та Хермон співають про Ймення Твоє.
PS|89|13|(89-14) Могутнє рамено Твоє, рука Твоя сильна, висока правиця Твоя!
PS|89|14|(89-15) Справедливість та право підстава престолу Твого, милість та правда обличчя Твоє випереджують!
PS|89|15|(89-16) Блаженний народ, що знає він поклик святковий, Господи, вони ходять у світлі обличчя Твого!
PS|89|16|(89-17) Радіють вони цілий день Твоїм іменням, і підвищуються Твоєю справедливістю,
PS|89|17|(89-18) бо окраса їхньої сили то Ти, а Твоєю зичливістю ріг наш підноситься,
PS|89|18|(89-19) бо щит наш Господній, а цар наш від Святого ізраїлевого!
PS|89|19|(89-20) Тоді богобійним Своїм промовляв Ти в об'явленні та говорив: Я поклав допомогу на сильного, Я вибранця підніс із народу:
PS|89|20|(89-21) знайшов Я Давида, Свого раба, Я його намастив Своєю святою оливою,
PS|89|21|(89-22) щоб із ним була сильна рука Моя, а рамено Моє вміцнило його!
PS|89|22|(89-23) Ворог на нього не нападе, а син беззаконня не буде його переслідувати,
PS|89|23|(89-24) його ворогів поб'ю перед обличчям його, і вдарю його ненависників!
PS|89|24|(89-25) із ним Моя вірність та милість Моя, а Йменням Моїм його ріг піднесеться,
PS|89|25|(89-26) і Я покладу його руку на море, і на ріки правицю його.
PS|89|26|(89-27) Він Мене буде звати: Отець Ти мій, Бог мій, і скеля спасіння мого!
PS|89|27|(89-28) Я вчиню його теж перворідним, найвищим над земних царів.
PS|89|28|(89-29) Свою милість для нього навіки сховаю, і Мій заповіт йому вірний,
PS|89|29|(89-30) і насіння його покладу Я навіки, а трона його як дні неба!
PS|89|30|(89-31) Коли ж його діти покинуть Закона Мого, і не будуть держатись наказів Моїх,
PS|89|31|(89-32) коли ізневажать Мої постанови, і не будуть держатись наказів Моїх,
PS|89|32|(89-33) тоді палицею навіщу їхню провину, та поразами їхнє беззаконня!
PS|89|33|(89-34) А ласки Своєї від нього Я не заберу, і не зраджу його в Своїй вірності,
PS|89|34|(89-35) не збезчещу Свого заповіту, а що було з уст Моїх вийшло, того не зміню!
PS|89|35|(89-36) Одне в Своїй святості Я присягнув, не повім Я неправди Давидові:
PS|89|36|(89-37) повік буде насіння його, а престол його передо Мною як сонце,
PS|89|37|(89-38) як місяць, він буде стояти повіки, і Свідок на хмарі правдивий... Села.
PS|89|38|(89-39) А Ти опустив та обридив, розгнівався Ти на Свого помазанця,
PS|89|39|(89-40) Ти неважливим зробив заповіта Свого раба, Ти скинув на землю корону його,
PS|89|40|(89-41) всю горожу його поламав, твердині його обернув на руїну!...
PS|89|41|(89-42) Всі грабують його, хто проходить дорогою, він став для сусідів своїх посміховищем...
PS|89|42|(89-43) Підніс Ти правицю його переслідувачів, усіх його ворогів Ти потішив,
PS|89|43|(89-44) і Ти відвернув вістря шаблі його... у війні ж не підтримав його...
PS|89|44|(89-45) Ти слави позбавив його, а трона його повалив був на землю,
PS|89|45|(89-46) скоротив Ти був дні його молодости, розтягнув над ним сором! Села.
PS|89|46|(89-47) Доки, Господи, будеш ховатись назавжди, доки буде палати Твій гнів, як огонь?
PS|89|47|(89-48) Пам'ятай же про мене, яка довгота життя людського? Для чого створив Ти всіх людських синів на ніщо?
PS|89|48|(89-49) Котрий чоловік буде жити, а смерти на бачитиме, збереже свою душу від сили шеолу? Села.
PS|89|49|(89-50) Де Твої перші милості, Господи, що їх присягав Ти Давидові у Своїй вірності?
PS|89|50|(89-51) Згадай, Господи, про ганьбу рабів Своїх, яку я ношу в своїм лоні від усіх великих народів,
PS|89|51|(89-52) якою Твої вороги зневажають, о Господи, і кроки Твого помазанця безславлять!
PS|89|52|(89-53) Благословенний навіки Господь! Амінь і амінь!
PS|90|1|Молитва Мойсея, чоловіка Божого. Господи, пристановищем нашим Ти був з роду в рід!
PS|90|2|Перше ніж гори народжені, і поки Ти витворив землю та світ, то від віку й до віку Ти Бог!
PS|90|3|Ти людину вертаєш до пороху, і кажеш: Вернітеся, людські сини!
PS|90|4|Бо в очах Твоїх тисяча літ, немов день той вчорашній, який проминув, й як сторожа нічна...
PS|90|5|Пустив Ти на них течію, вони стали, як сон, вони, як трава, що минає:
PS|90|6|уранці вона розцвітає й росте, а на вечір зів'яне та сохне!
PS|90|7|Бо від гніву Твого ми гинемо, і пересердям Твоїм перестрашені,
PS|90|8|Ти наші провини поклав перед Себе, гріхи ж нашої молодости на світло Свого лиця!
PS|90|9|Бо всі наші дні промайнули у гніві Твоїм, скінчили літа ми свої, як зідхання...
PS|90|10|Дні літ наших у них сімдесят літ, а при силах вісімдесят літ, і гордощі їхні страждання й марнота, бо все швидко минає, і ми відлітаємо...
PS|90|11|Хто відає силу гніву Твого? А Твоє пересердя як страх перед Тобою!
PS|90|12|Навчи нас лічити отак наші дні, щоб ми набули серце мудре!
PS|90|13|Привернися ж, о Господи, доки терпітимемо? і пожалій Своїх рабів!
PS|90|14|Насити нас уранці Своїм милосердям, і ми будемо співати й радіти по всі наші дні!
PS|90|15|Порадуй же нас за ті дні, коли Ти впокоряв нас, за ті роки, що в них ми зазнали лихого!
PS|90|16|Нехай виявиться Твоє діло рабам Твоїм, а величність Твоя їхнім синам,
PS|90|17|і хай буде над нами благовоління Господа, Бога нашого, і діло рук наших утверди нам, і діло рук наших утверди його!
PS|91|1|Хто живе під покровом Всевишнього, хто в тіні Всемогутнього мешкає,
PS|91|2|той скаже до Господа: Охороно моя та твердине моя, Боже мій, я надіюсь на Нього!
PS|91|3|Бо Він тебе вирве з тенет птахолова, з моровиці згубної,
PS|91|4|Він пером Своїм вкриє тебе, і під крильми Його заховаєшся ти! Щит та лук Його правда.
PS|91|5|Не будеш боятися страху нічного, ані стріли, що вдень пролітає,
PS|91|6|ані зарази, що в темряві ходить, ані моровиці, що нищить опівдні,
PS|91|7|впаде тисяча з боку від тебе, і десять тисяч праворуч від тебе, до тебе ж не дійде!...
PS|91|8|Тільки своїми очима подивишся, і заплату безбожним попобачиш,
PS|91|9|бо Господа, охорону мою, Всевишнього ти учинив за своє пристановище!
PS|91|10|Тебе зло не спіткає, і до намету твого вдар не наблизиться,
PS|91|11|бо Своїм Анголам Він накаже про тебе, щоб тебе пильнували на всіх дорогах твоїх,
PS|91|12|на руках вони будуть носити тебе, щоб не вдарив об камінь своєї ноги!
PS|91|13|На лева й вужа ти наступиш, левчука й крокодила ти будеш топтати!
PS|91|14|Що бажав він Мене, то його збережу, зроблю його сильним, бо знає ім'я Моє він;
PS|91|15|як він Мене кликатиме, то йому відповім, Я з ним буду в недолі, врятую його та прославлю його,
PS|91|16|і довгістю днів Я насичу його, і він бачити буде спасіння Моє!
PS|92|1|Псалом. Пісня на день суботній. (92-2) То добре, щоб дякувати Господеві й виспівувати Ймення Твоє, о Всевишній,
PS|92|2|(92-3) вранці розповідати про милість Твою, а ночами про правду Твою
PS|92|3|(92-4) на десятиструнній й на арфі, на лютні та гуслах,
PS|92|4|(92-5) бо потішив мене Ти, о Господи, вчинком Своїм, про діла Твоїх рук я співаю!
PS|92|5|(92-6) Які то величні діла Твої, Господи, дуже глибокі думки Твої,
PS|92|6|(92-7) нерозумна людина не знає, а недоумок не зрозуміє того!
PS|92|7|(92-8) Коли несправедливі ростуть, як трава, і цвітуть всі злочинці, то на те, щоб навіки були вони знищені,
PS|92|8|(92-9) а Ти, Господи, на висоті повік-віку!
PS|92|9|(92-10) Бо ось вороги Твої, Господи, бо ось вороги Твої згинуть, розпорошаться всі беззаконники!
PS|92|10|(92-11) і Ти рога мого підніс немов в однорожця, мене намастив Ти оливою свіжою.
PS|92|11|(92-12) і дивилося око моє на занепад моїх ворогів, тих злочинців, що на мене встають, почують про це мої уші!
PS|92|12|(92-13) Зацвіте справедливий, як пальма, і виженеться, немов кедр на Ливані,
PS|92|13|(92-14) посаджені в домі Господнім цвітуть на подвір'ях нашого Бога,
PS|92|14|(92-15) іще в сивині вони будуть цвісти, будуть ситі та свіжі,
PS|92|15|(92-16) щоб розповідати, що щирий Господь, моя скеля, і в Ньому неправди нема!
PS|93|1|Царює Господь, зодягнувся у велич, зодягнувся Господь, оперезався Він силою, і міцно поставлений всесвіт, щоб не захитався!
PS|93|2|Престол Твій поставлений міцно спрадавна, від вічности Ти!
PS|93|3|Ріки піднесли, о Господи, ріки піднесли свій гуркіт, ріки будуть підносити шум від удару їхніх хвиль,
PS|93|4|та над гуркіт великих тих вод, над морські потужнії хвилі, могутніший Господь у висоті!
PS|93|5|Свідоцтва Твої дуже певні, а дому Твоєму належиться святість, о Господи, на довгії дні!
PS|94|1|Бог помсти Господь, Бог помсти з'явився,
PS|94|2|піднесися, о Судде землі, бундючним заплату віддай!
PS|94|3|Аж доки безбожні, о Господи, аж доки безбожні втішатися будуть?
PS|94|4|Доки будуть верзти, говорити бундючно, доки будуть пишатись злочинці?
PS|94|5|Вони тиснуть народ Твій, о Господи, а спадок Твій вони мучать...
PS|94|6|Вдову та чужинця вбивають вони, і мордують сиріт
PS|94|7|та й говорять: Не бачить Господь, і не завважить Бог Яковів...
PS|94|8|Зрозумійте це ви, нерозумні в народі, а ви, убогі на розум, коли наберетеся глузду?
PS|94|9|Хіба Той, що ухо щепив, чи Він не почує? Хіба Той, що око створив, чи Він не побачить?
PS|94|10|Хіба Той, що карає народи, чи Він не скартає, Він, що навчає людину знання?
PS|94|11|Господь знає всі людські думки, що марнота вони!
PS|94|12|Блаженний той муж, що його Ти караєш, о Господи, і з Закону Свого навчаєш його,
PS|94|13|щоб його заспокоїти від лиходення, аж поки не викопана буде яма безбожному,
PS|94|14|бо Господь не опустить народу Свого, а спадку Свого не полишить,
PS|94|15|бо до праведности суд повернеться, а за ним всі невинного серця!
PS|94|16|Хто встане зо мною навпроти злостивих, хто встане зо мною навпроти злочинців?
PS|94|17|Коли б не Господь мені в поміч, то душа моя трохи була б не лягла в царство смерти!...
PS|94|18|Коли я кажу: Похитнулась нога моя, то, Господи, милість Твоя підпирає мене!
PS|94|19|Коли мої думки болючі в нутрі моїм множаться, то розради Твої веселять мою душу!
PS|94|20|Чи престол беззаконня з Тобою з'єднається, той, що гріх учиняє над право?
PS|94|21|Збираються проти душі справедливого, і чисту кров винуватять.
PS|94|22|і Господь став для мене твердинею, і мій Бог став за скелю притулку мого,
PS|94|23|і Він їхню силу на них повернув, і злом їхнім їх нищить, їх нищить Господь, Бог наш!
PS|95|1|Ходіть, заспіваймо Господеві, покликуймо радісно скелі спасіння нашого,
PS|95|2|хвалою обличчя Його випереджуймо, співаймо для Нього пісні,
PS|95|3|бо Господь Бог великий, і великий Він Цар над богами всіма,
PS|95|4|що в Нього в руці глибини землі, і Його верхогір'я гірські,
PS|95|5|що море Його, і вчинив Він його, і руки Його суходіл уформували!
PS|95|6|Прийдіть, поклонімося, і припадім, на коліна впадім перед Господом, що нас учинив!
PS|95|7|Він наш Бог, а ми люди Його пасовиська й отара руки Його. Сьогодні, коли Його голос почуєте,
PS|95|8|не робіте твердим серця вашого, мов при Мериві, немов на пустині в день спроби,
PS|95|9|коли ваші батьки Мене брали на спробу, Мене випробовували, також бачили діло Моє.
PS|95|10|Сорок літ був огидним Мені оцей рід, й Я сказав: Цей народ блудосерді вони, й не пізнали доріг Моїх,
PS|95|11|тому заприсягся Я в гніві Своїм, що до місця Мого відпочинку не ввійдуть вони!
PS|96|1|Співайте для Господа пісню нову, уся земле, співайте для Господа!
PS|96|2|Співайте для Господа, благословляйте ім'я Його, з дня на день сповіщайте спасіння Його!
PS|96|3|Розповідайте про славу Його між поганами, про чуда Його між усіми народами,
PS|96|4|бо великий Господь і прославлений вельми, Він грізний понад богів усіх!
PS|96|5|Бо всі боги народів божки, а Господь створив небеса,
PS|96|6|перед лицем Його слава та велич, сила й краса у святині Його!
PS|96|7|Дайте Господу, роди народів, дайте Господу славу та силу,
PS|96|8|дайте Господу славу ймення Його, жертви приносьте і входьте в подвір'я Його!
PS|96|9|Додолу впадіть ув оздобі святій перед Господом, тремтіть перед обличчям Його, уся земле,
PS|96|10|сповістіть між народами: Царює Господь! Він вселенну зміцнив, щоб не захиталась, Він буде судити людей справедливо!
PS|96|11|Хай небо радіє, і хай веселиться земля, нехай гримить море й усе, що у нім,
PS|96|12|нехай поле радіє та все, що на ньому! Нехай заспівають тоді всі дерева лісні,
PS|96|13|перед Господнім лицем, бо гряде Він, бо землю судити гряде, Він за справедливістю буде судити вселенну, і народи по правді Своїй!
PS|97|1|Царює Господь: хай радіє земля, нехай веселяться численні острови!
PS|97|2|Хмара та морок круг Нього, справедливість та право підстава престолу Його.
PS|97|3|Огонь іде перед лицем Його, і ворогів Його палить навколо.
PS|97|4|Освітили вселенну Його блискавиці, те бачить земля та тремтить!
PS|97|5|Гори, як віск, розтопилися перед обличчям Господнім, перед обличчям Господа всієї землі.
PS|97|6|Небо розповідає про правду Його, й бачать славу Його всі народи.
PS|97|7|Нехай посоромлені будуть усі, хто ідолам служить, хто божками вихвалюється! Додолу впадіть перед Ним, усі боги!
PS|97|8|Почув і звеселився Сіон, і потішились Юдині дочки через Твої присуди, Господи,
PS|97|9|бо над усією землею Найвищий Ти, Господи, над богами всіма Ти піднесений сильно!
PS|97|10|Хто Господа любить, ненавидьте зло! Хто рятує душі святих Своїх, Той визволить їх із руки несправедливих.
PS|97|11|Світло сіється для справедливого, а для простосердих розрада.
PS|97|12|Радійте, праведні, Господом, і славте Його святу пам'ять!
PS|98|1|Псалом. Співайте для Господа пісню нову, бо Він чуда вчинив! Йому помогла правиця Його та святе рамено Його.
PS|98|2|Спасіння Своє Господь виявив, перед очима народів відкрив Свою правду.
PS|98|3|Пам'ятає Він Якову милість Свою, й Свою вірність для дому ізраїля. Бачать всі кінці землі те спасіння, що чинить наш Бог.
PS|98|4|Уся земле, викликуйте Господу, покликуйте радісно, і співайте та грайте!
PS|98|5|Грайте Господеві на гуслах, на гуслах і піснопінням,
PS|98|6|на сурмах і голосом рогу викликуйте перед обличчям Царя Цього й Господа!
PS|98|7|Нехай шумить море й усе, що у ньому, вселенна й мешканці її,
PS|98|8|ріки хай плещуть в долоні, разом радіють хай гори
PS|98|9|перед обличчям Господнім, бо Він землю судити гряде: Він за справедливістю буде судити вселенну, і народи по правді!
PS|99|1|Царює Господь, і народи тремтять, сидить на Херувимах, і трясеться земля!
PS|99|2|Великий Господь на Сіоні, і піднесений Він над усіма народами!
PS|99|3|Хай ім'я Твоє славлять, велике й грізне воно!
PS|99|4|А сила Царя любить право, справедливість Ти міцно поставив, Ти Якову право та правду вчинив!
PS|99|5|Звеличуйте Господа, нашого Бога, і вклоняйтесь підніжкові ніг Його, Він бо Святий!
PS|99|6|Мойсей й Аарон серед священиків Його, а Самуїл серед тих, що кличуть імення Його. Вони кликали до Господа, і Він вислухав їх,
PS|99|7|у стовпі хмари до них говорив. Вони зберігали свідоцтва Його й постанови, що Він дав був для них.
PS|99|8|Господи, Боже наш, Ти вислуховував їх, Ти був для них Богом вибачливим, але мстився за їхні діла.
PS|99|9|Звеличуйте Господа, нашого Бога, і вклоняйтеся перед горою святою Його, бо Святий Господь, Бог наш!
PS|100|1|Вдячний псалом. Уся земле, покликуйте Господу!
PS|100|2|Служіть Господеві із радістю, перед обличчя Його підійдіте зо співом!
PS|100|3|Знайте, що Господь Бог Він, Він нас учинив, і Його ми, Його ми народ та отара Його пасовиська.
PS|100|4|Увійдіть в Його брами з подякуванням, на подвір'я Його з похвалою! Виславляйте Його, ім'я Його благословляйте,
PS|100|5|бо добрий Господь, Його милість навіки, а вірність Його з роду в рід!
PS|101|1|Псалом Давидів. Я виспівувати буду про милість та суд, я буду співати до Тебе, о Господи,
PS|101|2|придивлятимуся до дороги невинного. Коли прийдеш до мене? Я буду ходити в невинності серця свого серед дому мого,
PS|101|3|не поставлю я перед очима своїми речі нікчемної, діло відступства ненавиджу, не приляже до мене воно,
PS|101|4|перекірливе серце відходить від мене, лихого не знаю!
PS|101|5|Хто таємно обчорнює ближнього свого, я знищу того, високоокого й гордосердого, його не стерплю!
PS|101|6|Мої очі на вірних землі, щоб сиділи зо мною. Хто ходить дорогою невинного, той буде служити мені.
PS|101|7|Обманець не сяде в середині дому мого, і міцно не стане навпроти очей моїх неправдомовець!
PS|101|8|Всіх безбожних землі буду нищити кожного ранку, щоб з міста Господнього вигубити всіх злочинців!
PS|102|1|Молитва вбогого, коли він слабне та перед Господнім лицем виливає мову свою. (102-2) Господи, вислухай молитву мою, і благання моє нехай дійде до Тебе!
PS|102|2|(102-3) Не ховай від мене обличчя Свого, в день недолі моєї схили Своє ухо до мене, в день благання озвися небавом до мене!
PS|102|3|(102-4) Бо минають, як дим, мої дні, а кості мої немов висохли в огнищі...
PS|102|4|(102-5) Як трава та побите та висохло серце моє, так що я забував їсти хліб свій...
PS|102|5|(102-6) Від зойку стогнання мого прилипли до тіла мого мої кості...
PS|102|6|(102-7) Уподобився я пеликанові пустині, я став, як той пугач руїн!
PS|102|7|(102-8) Я безсонний, і став, немов пташка самотня на дасі...
PS|102|8|(102-9) Увесь день ображають мене вороги мої, ті, хто з мене кепкує, заприсяглись проти мене!
PS|102|9|(102-10) і попіл я їм, немов хліб, а напої свої із плачем перемішую,
PS|102|10|(102-11) через гнів Твій та лютість Твою, бо підняв був мене Ти та й кинув мене...
PS|102|11|(102-12) Мої дні як похилена тінь, а я сохну, немов та трава!
PS|102|12|(102-13) А Ти, Господи, будеш повік пробувати, а пам'ять Твоя з роду в рід.
PS|102|13|(102-14) Ти встанеш та змилуєшся над Сіоном, бо час учинити йому милосердя, бо прийшов речінець,
PS|102|14|(102-15) бо раби Твої покохали й каміння його, і порох його полюбили!
PS|102|15|(102-16) і будуть боятись народи Господнього Ймення, а всі земні царі слави Твоєї.
PS|102|16|(102-17) Бо Господь побудує Сіона, появиться в славі Своїй.
PS|102|17|(102-18) До молитви забутих звернеться Він, і молитви їхньої не осоромить.
PS|102|18|(102-19) Запишеться це поколінню майбутньому, і народ, який створений буде, хвалитиме Господа,
PS|102|19|(102-20) бо споглянув Він із високости святої Своєї, Господь зорив на землю з небес,
PS|102|20|(102-21) щоб почути зідхання ув'язненого, щоб на смерть прирокованих визволити,
PS|102|21|(102-22) щоб розповідати про Ймення Господнє в Сіоні, а в Єрусалимі про славу Його,
PS|102|22|(102-23) коли разом зберуться народи й держави служити Господеві.
PS|102|23|(102-24) Мою силу в дорозі Він виснажив, дні мої скоротив...
PS|102|24|(102-25) Я кажу: Боже мій, не бери Ти мене в половині днів моїх! Твої роки на вічні віки.
PS|102|25|(102-26) Колись землю Ти був заклав, а небо то чин Твоїх рук,
PS|102|26|(102-27) позникають вони, а Ти будеш стояти... і всі вони, як одежа, загинуть, Ти їх зміниш, немов те вбрання, і минуться вони...
PS|102|27|(102-28) Ти ж Той Самий, а роки Твої не закінчаться!
PS|102|28|(102-29) Сини Твоїх рабів будуть жити, а їхнє насіння стоятиме міцно перед обличчям Твоїм!
PS|103|1|Давидів. Благослови, душе моя, Господа, і все нутро моє святе Ймення Його!
PS|103|2|Благослови, душе моя, Господа, і не забувай за всі добродійства Його!
PS|103|3|Всі провини Твої Він прощає, всі недуги твої вздоровляє.
PS|103|4|Від могили життя твоє Він визволяє, Він милістю та милосердям тебе коронує.
PS|103|5|Він бажання твоє насичає добром, відновиться, мов той орел, твоя юність!
PS|103|6|Господь чинить правду та суд для всіх переслідуваних.
PS|103|7|Він дороги Свої об'явив був Мойсеєві, діла Свої дітям ізраїлевим.
PS|103|8|Щедрий і милосердний Господь, довготерпеливий і многомилостивий.
PS|103|9|Не завжди на нас ворогує, і не навіки заховує гнів.
PS|103|10|Не за нашими прогріхами Він поводиться з нами, і відплачує нам не за провинами нашими.
PS|103|11|Бо як високо небо стоїть над землею, велика така Його милість до тих, хто боїться Його,
PS|103|12|як далекий від заходу схід, так Він віддалив від нас наші провини!
PS|103|13|Як жалує батько дітей, так Господь пожалівся над тими, хто боїться Його,
PS|103|14|бо знає Він створення наше, пам'ятає, що ми порох:
PS|103|15|чоловік як трава дні його, немов цвіт польовий так цвіте він,
PS|103|16|та вітер перейде над ним і немає його, і вже місце його не пізнає його...
PS|103|17|А милість Господня від віку й до віку на тих, хто боїться Його, і правда Його над синами синів,
PS|103|18|що Його заповіта додержують, і що пам'ятають накази Його, щоб виконувати їх!
PS|103|19|Господь міцно поставив на Небі престола Свого, а Царство Його над усім володіє.
PS|103|20|Благословіть Господа, Його Анголи, велетні сильні, що виконуєте Його слово, щоб слухати голосу слів Його!
PS|103|21|Благословіть Господа, усі сили небесні Його, слуги Його, що чините волю Його!
PS|103|22|Благословіть Господа, всі діла Його, на всіх місцях царювання Його! Благослови, душе моя, Господа!
PS|104|1|Благослови, душе моя, Господа! Господи, Боже мій, Ти вельми великий, зодягнувся Ти в велич та в славу!
PS|104|2|Зодягає Він світло, як шати, небеса простягає, немов би завісу.
PS|104|3|Він ставить на водах палати Свої, хмари кладе за Свої колесниці, ходить на крилах вітрових!
PS|104|4|Він чинить вітри за Своїх посланців, палючий огонь за Своїх слуг.
PS|104|5|Землю Ти вґрунтував на основах її, щоб на вічні віки вона не захиталась,
PS|104|6|безоднею вкрив Ти її, немов шатою. Стала вода над горами,
PS|104|7|від погрози Твоєї вона втекла, від гуркоту грому Твого побігла вона,
PS|104|8|виходить на гори та сходить в долини, на місце, що Ти встановив був для неї.
PS|104|9|Ти границю поклав, щоб її вона не перейшла, щоб вона не вернулася землю покрити.
PS|104|10|Він джерела пускає в потоки, що пливуть між горами,
PS|104|11|напувають вони всю пільну звірину, ними дикі осли гасять спрагу свою.
PS|104|12|Птаство небесне над ними живе, видає воно голос з-посеред галузок.
PS|104|13|Він напоює гори з палаців Своїх, із плоду чинів Твоїх земля сититься.
PS|104|14|Траву для худоби вирощує, та зеленину для праці людині, щоб хліб добувати з землі,
PS|104|15|і вино, що серце людині воно звеселяє, щоб більш від оливи блищало обличчя, і хліб, що серце людині зміцняє.
PS|104|16|Насичуються Господні дерева, ті кедри ливанські, що Ти насадив,
PS|104|17|що там кубляться птахи, бузько, кипариси мешкання його.
PS|104|18|Гори високі для диких козиць, скелі сховище скельним звіринам.
PS|104|19|і місяця Він учинив для означення часу, сонце знає свій захід.
PS|104|20|Темноту Ти наводиш і ніч настає, в ній порушується вся звірина лісна,
PS|104|21|ричать левчуки за здобичею та шукають від Бога своєї поживи.
PS|104|22|Сонце ж засвітить вони повтікають, та й кладуться по норах своїх.
PS|104|23|Людина виходить на працю свою, й на роботу свою аж до вечора.
PS|104|24|Які то численні діла Твої, Господи, Ти мудро вчинив їх усіх, Твого творива повна земля!
PS|104|25|Ось море велике й розлогошироке, там повзюче, й числа їм немає, звірина мала та велика!
PS|104|26|Ходять там кораблі, там той левіятан, якого створив Ти, щоб бавитися йому в морі.
PS|104|27|Вони всі чекають Тебе, щоб Ти часу свого поживу їм дав.
PS|104|28|Даєш їм збирають вони, руку Свою розкриваєш добром насичаються.
PS|104|29|Ховаєш обличчя Своє то вони перелякані, забираєш їм духа вмирають вони, та й вертаються до свого пороху.
PS|104|30|Посилаєш Ти духа Свого вони творяться, і Ти відновляєш обличчя землі.
PS|104|31|Нехай буде слава Господня навіки, хай ділами Своїми радіє Господь!
PS|104|32|Він погляне на землю й вона затремтить, доторкнеться до гір і димують вони!
PS|104|33|Я буду співати Господеві в своєму житті, буду грати для Бога мого, аж поки живу!
PS|104|34|Буде приємна Йому моя мова, я Господом буду радіти!
PS|104|35|Нехай згинуть грішні з землі, а безбожні немає вже їх! Благослови, душе моя, Господа! Алілуя!
PS|105|1|Дякуйте Господу, кличте ім'я Його, серед народів звіщайте про чини Його!
PS|105|2|Співайте Йому, грайте Йому, говоріть про всі чуда Його!
PS|105|3|Хваліться святим Його Йменням, хай тішиться серце шукаючих Господа!
PS|105|4|Пошукуйте Господа й силу Його, лице Його завжди шукайте!
PS|105|5|Пам'ятайте про чуда Його, які Він учинив, про ознаки Його та про присуди уст Його,
PS|105|6|ви, насіння Авраама, раба Його, сини Яковові, вибранці Його!
PS|105|7|Він Господь, Бог наш, по цілій землі Його присуди!
PS|105|8|Він пам'ятає навіки Свого заповіта, те слово, яке наказав був на тисячу родів,
PS|105|9|що склав Він його з Авраамом, і присягу Свою для ісака.
PS|105|10|Він поставив її за Закона для Якова, ізраїлеві заповітом навіки,
PS|105|11|говорячи: Я дам тобі Край ханаанський, частину спадщини для вас!
PS|105|12|Тоді їх було невелике число, нечисленні були та приходьки на ній,
PS|105|13|і ходили вони від народу до народу, від царства до іншого люду.
PS|105|14|Не дозволив нікому Він кривдити їх, і за них Він царям докоряв:
PS|105|15|Не доторкуйтеся до Моїх помазанців, а пророкам Моїм не робіте лихого!
PS|105|16|і покликав Він голод на землю, всяке хлібне стебло поламав.
PS|105|17|Перед їхнім обличчям Він мужа послав, за раба Йосип проданий був.
PS|105|18|Кайданами мучили ноги його, залізо пройшло в його тіло,
PS|105|19|аж до часу виповнення слова Його, слово Господнє його було виявило.
PS|105|20|Цар послав і його розв'язав, володар народів і його був звільнив.
PS|105|21|Він настановив його паном над домом своїм, і володарем над усім маєтком своїм,
PS|105|22|щоб в'язнив він його можновладців по волі своїй, а старших його умудряв.
PS|105|23|і ізраїль прибув до Єгипту, і Яків замешкав у Хамовім краї.
PS|105|24|А народ Свій Він сильно розмножив, і зробив був ряснішим його від його ворогів.
PS|105|25|Він перемінив їхнє серце, щоб народа Його ненавиділи, щоб брались на хитрощі проти рабів Його.
PS|105|26|Він послав був Мойсея, Свого раба, Аарона, що вибрав його,
PS|105|27|вони положили були серед них Його речі знаменні, та чуда у Хамовім краї.
PS|105|28|Він темноту наслав і потемніло, і вони не противились слову Його.
PS|105|29|Він перемінив їхню воду на кров, і вморив їхню рибу.
PS|105|30|Їхній край зароївся був жабами, навіть в покоях царів їхніх.
PS|105|31|Він сказав й прибули рої мух, воші в цілому обширі їхньому.
PS|105|32|Він градом зробив їхній дощ, палючий огонь на їхню землю.
PS|105|33|і Він повибивав виноград їхній та фіґове дерево їхнє, і деревину на обширі їхньому повиломлював.
PS|105|34|Він сказав і найшла сарана та гусінь без ліку,
PS|105|35|усю ярину в їхнім краї пожерла, і плід землі їхньої з'їла.
PS|105|36|і Він повбивав усіх первістків в їхньому краї, початок усякої їхньої сили.
PS|105|37|і Він випровадив їх у сріблі та в золоті, і серед їхніх племен не було, хто б спіткнувся.
PS|105|38|Єгипет радів, коли вийшли вони, бо страх перед ними напав був на них.
PS|105|39|Він хмару простяг на заслону, а огонь на освітлення ночі.
PS|105|40|Зажадав був ізраїль і Він перепелиці наслав, і хлібом небесним Він їх годував.
PS|105|41|Відчинив був Він скелю й линула вода, потекли були ріки в пустинях,
PS|105|42|бо Він пам'ятав за святе Своє слово, за Авраама, Свого раба.
PS|105|43|і Він з радістю вивів народ Свій, зо співом вибранців Своїх,
PS|105|44|і їм землю народів роздав, і посіли вони працю людів,
PS|105|45|щоб виконували Його заповіді, та закони Його берегли! Алілуя!
PS|106|1|Алілуя! Дякуйте Господу, добрий бо Він, бо навіки Його милосердя!
PS|106|2|Хто розкаже про велич Господню, розповість усю славу Його?
PS|106|3|Блаженні, хто держиться права, хто чинить правду кожного часу!
PS|106|4|Згадай мене, Господи, в ласці Своїй до народу Свого, відвідай мене спасінням Своїм,
PS|106|5|щоб побачити добре вибранців Твоїх, щоб я тішився радощами Твого народу, і хвалився зо спадком Твоїм!
PS|106|6|Ми згрішили з батьками своїми, скривили, неправдиве чинили...
PS|106|7|Не зважали на чуда Твої батьки наші в Єгипті, многоти Твоїх ласк не пригадували й бунтувались над морем, над морем Червоним.
PS|106|8|Та Він ради Ймення Свого їх спас, щоб виявити Свою силу.
PS|106|9|Він кликнув на море Червоне і висохло, і Він їх повів через морські глибини, немов по пустині!...
PS|106|10|і Він спас їх з руки неприятеля, визволив їх з руки ворога,
PS|106|11|і закрила вода супротивників їхніх, жоден з них не зостався!
PS|106|12|Тоді то в слова Його ввірували, виспівували Йому славу.
PS|106|13|Та скоро забули вони Його чин, не чекали поради Його,
PS|106|14|і палали в пустині жаданням, і Бога в пустині ізнов випробовували,
PS|106|15|і Він їхнє жадання їм дав, але худість послав в їхню душу...
PS|106|16|Та Мойсею позаздрили в таборі, й Ааронові, святому Господньому.
PS|106|17|Розкрилась земля і Датана поглинула, Авіронові збори накрила,
PS|106|18|і огонь запалав на їхніх зборах, і полум'я те попалило безбожних...
PS|106|19|Зробили тельця на Хориві, і били поклони бовванові вилитому,
PS|106|20|і змінили вони свою славу на образ вола, що траву пожирає,
PS|106|21|забули про Бога, свого Спасителя, що велике в Єгипті вчинив,
PS|106|22|у землі Хамовій чуда, страшні речі над морем Червоним...
PS|106|23|і сказав Він понищити їх, коли б не Мойсей, вибранець Його, що став був у виломі перед обличчям Його відвернути Його гнів, щоб не шкодив!
PS|106|24|Погордили землею жаданою, не повірили слову Його,
PS|106|25|і ремствували по наметах своїх, неслухняні були до Господнього голосу.
PS|106|26|і Він підійняв Свою руку на них, щоб їх повалити в пустині,
PS|106|27|і щоб повалити їхнє потомство посеред народів, та щоб розпорошити їх по країнах!
PS|106|28|і служили Ваалові пеорському, й їли вони жертви мертвих,
PS|106|29|і ділами своїми розгнівали Бога, тому вдерлась зараза між них!
PS|106|30|і встав тоді Пінхас та й розсудив, і зараза затрималась,
PS|106|31|і йому пораховано в праведність це, з роду в рід аж навіки.
PS|106|32|і розгнівали Бога вони над водою Меріви, і через них стало зле для Мойсея,
PS|106|33|бо духа його засмутили, і він говорив нерозважно устами своїми...
PS|106|34|Вони не познищували тих народів, що Господь говорив їм про них,
PS|106|35|і помішались з поганами, та їхніх учинків навчились.
PS|106|36|і божищам їхнім служили, а ті пасткою стали для них...
PS|106|37|і приносили в жертву синів своїх, а дочок своїх демонам,
PS|106|38|і кров чисту лили, кров синів своїх і дочок своїх, що їх у жертву приносили божищам ханаанським. і через кривавий переступ земля посквернилась,
PS|106|39|і стали нечисті вони через учинки свої, і перелюб чинили ділами своїми...
PS|106|40|і проти народу Свого запалав гнів Господній, і спадок Його Йому став огидним,
PS|106|41|і віддав їх у руку народів, і їхні ненависники панували над ними,
PS|106|42|і їхні вороги їх гнобили, і вони впокорилися під їхню руку...
PS|106|43|Багато разів Він визволював їх, але вони вперті були своїм задумом, і пригноблено їх через їхню провину!
PS|106|44|Та побачив Він їхню тісноту, коли почув їхні благання,
PS|106|45|і Він пригадав їм Свого заповіта, і пожалував був за Своєю великою милістю,
PS|106|46|і збудив милосердя до них між усіма, що їх полонили!
PS|106|47|Спаси нас, о Господи, Боже наш, і нас позбирай з-між народів, щоб дякувати Йменню святому Твоєму, щоб Твоєю хвалитися славою!
PS|106|48|Благословенний Господь, Бог ізраїлів звіку й навіки! і ввесь народ нехай скаже: Амінь! Алілуя!
PS|107|1|Дякуйте Господу, добрий бо Він, бо навіки Його милосердя!
PS|107|2|хай так скажуть ті всі, що Господь урятував їх, що визволив їх з руки ворога,
PS|107|3|і з країв їх зібрав, від сходу й заходу, від півночі й моря!
PS|107|4|Блудили вони по пустині дорогою голою, осілого міста не знаходили,
PS|107|5|голодні та спрагнені, і в них їхня душа омлівала...
PS|107|6|і в недолі своїй вони Господа кликали, і Він визволяв їх від утисків їхніх!
PS|107|7|і Він їх попровадив дорогою простою, щоб до міста осілого йшли.
PS|107|8|Нехай же подяку складуть Господеві за милість Його, та за чуда Його синам людським,
PS|107|9|бо наситив Він спрагнену душу, а душу голодну наповнив добром!
PS|107|10|Ті, хто перебував був у темряві та в смертній тіні, то в'язні біди та заліза,
PS|107|11|бо вони спротивлялися Божим словам, і відкинули раду Всевишнього.
PS|107|12|Та Він упокорив їхнє серце терпінням, спіткнулись вони і ніхто не поміг,
PS|107|13|і в недолі своїй вони Господа кликали, і Він визволяв їх від утисків їхніх!
PS|107|14|і Він вивів їх з темряви й мороку, їхні ж кайдани сторощив.
PS|107|15|Нехай же подяку складуть Господеві за милість Його, та за чуда Його синам людським,
PS|107|16|бо Він поламав мідні двері, і засуви залізні зрубав!
PS|107|17|Нерозумні страждали за грішну дорогу свою й за свої беззаконня.
PS|107|18|Душа їхня від усякої їжі відверталася, і дійшли вони аж до брам смерти,
PS|107|19|і в недолі своїй вони Господа кликали, і Він визволяв їх від утисків їхніх,
PS|107|20|Він послав Своє слово та їх уздоровив, і їх урятував з їхньої хвороби!
PS|107|21|Нехай же подяку складуть Господеві за милість Його та за чуда Його синам людським,
PS|107|22|і хай жертви подяки приносять, і хай розповідають зо співом про чини Його!
PS|107|23|Ті, хто по морю пливе кораблями, хто чинить зайняття своє на великій воді,
PS|107|24|вони бачили чини Господні та чуда Його в глибині!
PS|107|25|Він скаже і буря зривається, і підносяться хвилі Його,
PS|107|26|до неба вони підіймаються, до безодні спадають, у небезпеці душа їхня хвилюється!
PS|107|27|Вони крутяться й ходять вперед та назад, як п'яний, і вся їхня мудрість бентежиться!
PS|107|28|Та в недолі своїй вони Господа кликали, і Він визволяв їх від утисків їхніх!
PS|107|29|Він змінює бурю на тишу, і стихають їхні хвилі,
PS|107|30|і раділи, що втихли вони, і Він їх привів до бажаної пристані.
PS|107|31|Нехай же подяку складуть Господеві за милість, та за чуда Його синам людським!
PS|107|32|Нехай величають Його на народньому зборі, і нехай вихваляють Його на засіданні старших!
PS|107|33|Він обертає річки в пустиню, а водні джерела на суходіл,
PS|107|34|плодючу землю на солончак через злобу мешканців її.
PS|107|35|Він пустиню обертає в водне болото, а землю суху в джерело,
PS|107|36|і голодних садовить Він там, а вони ставлять місто на мешкання,
PS|107|37|і поля засівають, і виноградники садять, і отримують плід урожаю!
PS|107|38|і благословляє Він їх, і сильно розмножуються, і одержують плід урожаю!
PS|107|39|Та змаліли вони й похилилися з утиску злого та з смутку.
PS|107|40|Виливає Він ганьбу на можних, і блудять вони без дороги в пустині,
PS|107|41|а вбогого Він підіймає з убозтва, і розмножує роди, немов ту отару.
PS|107|42|Це бачать правдиві й радіють, і закриває уста свої всяке безправ'я.
PS|107|43|Хто мудрий, той все це завважить, і познають вони милосердя Господнє!
PS|108|1|Пісня. Псалом Давидів. (108-2) Моє серце зміцнилося, Боже, я буду співати та славити разом з своєю хвалою!
PS|108|2|(108-3) Збудися ж ти, арфо та цитро, я буду будити досвітню зорю!
PS|108|3|(108-4) Я буду Тебе вихваляти, о Господи, серед народів, і буду співати Тобі між племенами,
PS|108|4|(108-5) бо більше від неба Твоє милосердя, а правда Твоя аж до хмар!
PS|108|5|(108-6) Піднесися ж, о Боже, над небо, а слава Твоя над усією землею!
PS|108|6|(108-7) Щоб любі Твої були визволені, Своєю правицею допоможи й обізвися до нас!
PS|108|7|(108-8) У святині Своїй Бог промовив: Нехай Я звеселюся, розділю Я Сихем, і долину Суккотську поміряю.
PS|108|8|(108-9) Належить Мені Ґілеад, і Мені Манасія, а Єфрем охорона Моєї голови, Юда берло Моє.
PS|108|9|(108-10) Моав то мідниця Мого миття, на Едом узуттям Своїм кину, над Филистеєю буду погукувати!
PS|108|10|(108-11) Хто мене запровадить до міста твердинного, хто до Едому мене приведе?
PS|108|11|(108-12) Хіба ж Ти покинув нас, Боже, і серед нашого війська не вийдеш вже, Боже?
PS|108|12|(108-13) Подай же нам поміч на ворога, людська бо поміч марнота!
PS|108|13|(108-14) Ми мужність покажемо в Бозі, і Він потопче противників наших!
PS|109|1|Для дириґетна хору. Псалом Давидів. Боже слави моєї, не будь мовчазливий,
PS|109|2|бо мої вороги порозкривали на мене уста нечестиві та пельки лукаві, язиком неправдивим говорять зо мною!
PS|109|3|і вони оточили мене словами ненависти, і без причини на мене воюють,
PS|109|4|обмовляють мене за любов мою, а я молюся за них,
PS|109|5|вони віддають мені злом за добро, і ненавистю за любов мою!
PS|109|6|Постав же над ним нечестивого, і по правиці його сатана нехай стане!
PS|109|7|Як буде судитись нехай вийде винним, молитва ж його бодай стала гріхом!
PS|109|8|Нехай дні його будуть короткі, хай інший маєток його забере!
PS|109|9|Бодай діти його стали сиротами, а жінка його удовою!
PS|109|10|і хай діти його все мандрують та жебрають, і нехай вони просять у тих, хто їх руйнував!
PS|109|11|Бодай їм тенета розставив лихвар на все, що його, і нехай розграбують чужі його працю!
PS|109|12|Щоб до нього ніхто милосердя не виявив, і бодай не було його сиротам милости!
PS|109|13|Щоб на знищення стали нащадки його, бодай було скреслене в другому роді ім'я їхнє!
PS|109|14|Беззаконня батьків його хай пам'ятається в Господа, і хай не стирається гріх його матері!
PS|109|15|Нехай будуть вони перед Господом завжди, а Він нехай вирве з землі їхню пам'ять,
PS|109|16|ворог бо не пам'ятав милосердя чинити, і напастував був людину убогу та бідну, та серцем засмучену, щоб убивати її!
PS|109|17|Полюбив він прокляття, бодай же на нього воно надійшло! і не хотів благословення, щоб воно віддалилось від нього!
PS|109|18|Зодягнув він прокляття, немов свою одіж, просякло воно, як вода, в його нутро, та в кості його, мов олива!
PS|109|19|Бодай воно стало йому за одежу, в яку зодягнеться, і за пояс, що завжди він ним підпережеться!
PS|109|20|Це заплата від Господа тим, хто мене обмовляє, на душу мою наговорює зло!
PS|109|21|А Ти Господи, Владико, зо мною зроби ради Ймення Свого, що добре Твоє милосердя, мене порятуй,
PS|109|22|бо я вбогий та бідний, і зранене серце моє в моїм нутрі!...
PS|109|23|Я ходжу, мов та тінь, коли хилиться день, немов сарана я відкинений!
PS|109|24|Коліна мої знесилилися з посту, і вихудло тіло моє з недостачі оливи,
PS|109|25|і я став для них за посміховище, коли бачать мене, головою своєю хитають...
PS|109|26|Поможи мені, Господи, Боже мій, за Своїм милосердям спаси Ти мене!
PS|109|27|і нехай вони знають, що Твоя це рука, що Ти, Господи, все це вчинив!
PS|109|28|Нехай проклинають вони, Ти ж поблагослови! Вони повстають, та нехай засоромлені будуть, а раб Твій радітиме!
PS|109|29|Хай зодягнуться ганьбою ті, хто мене обмовляє, і хай вони сором свій вдягнуть, як шату!
PS|109|30|Я устами своїми хвалитиму голосно Господа, і між багатьма Його славити буду,
PS|109|31|бо стоїть на правиці убогого Він для спасіння від тих, хто осуджує душу його!
PS|110|1|Псалом Давидів. Промовив Господь Господеві моєму: Сядь праворуч Мене, доки не покладу Я Твоїх ворогів за підніжка ногам Твоїм!
PS|110|2|Господь із Сіону пошле берло сили Своєї, пануй Ти поміж ворогами Своїми!
PS|110|3|Народ Твій готовий у день військового побору Твого, в оздобах святині із лоня зірниці прилине для Тебе, немов та роса, Твоя молодість.
PS|110|4|Поклявся Господь, і не буде жаліти: Ти священик навіки за чином Мелхиседековим.
PS|110|5|По правиці Твоїй розторощить Владика царів у день гніву Свого,
PS|110|6|Він буде судити між народами, землю виповнить трупами, розторощить Він голову в краї великім...
PS|110|7|Буде пити з струмка на дорозі, тому то підійме Він голову!
PS|111|1|Алілуя! Буду славити Господа з повного серця, в колі праведних та на згромадженні!
PS|111|2|Великі Господні діла, вони пожадані для всіх, хто їх любить!
PS|111|3|Його діло краса та величність, а правда Його пробуває навіки!
PS|111|4|Він пам'ятку чудам Своїм учинив, милостивий та щедрий Господь!
PS|111|5|Поживу дає Він для тих, хто боїться Його, заповіта Свого пам'ятає повік!
PS|111|6|Силу чинів Своїх об'явив Він народові Своєму, щоб спадщину народів їм дати.
PS|111|7|Діла рук Його правда та право, всі накази Його справедливі,
PS|111|8|вони кріпкі на вічні віки, вони зроблені вірністю і правотою!
PS|111|9|Послав Він Своєму народові визволення, заповіта Свого поставив навіки, святе та грізне Його Ймення!
PS|111|10|Початок премудрости страх перед Господом, добрий розум у тих, хто виконує це, Його слава навіки стоїть!
PS|112|1|Алілуя! Блажен муж, що боїться Господа, що заповіді Його любить!
PS|112|2|Буде сильним насіння його на землі, буде поблагословлений рід безневинних!
PS|112|3|Багатство й достаток у домі його, а правда його пробуває навіки!
PS|112|4|Світло сходить у темряві для справедливих, Він ласкавий, і милостивий, і праведний!
PS|112|5|Добрий муж милостивий та позичає, удержує справи свої справедливістю,
PS|112|6|і навіки він не захитається, у вічній пам'яті праведний буде!
PS|112|7|Не боїться він звістки лихої, його серце міцне, надію складає на Господа!
PS|112|8|Уміцнене серце його не боїться, бо він бачить нещастя поміж ворогами своїми!
PS|112|9|Він щедро убогим дає, його правда навіки стоїть, його ріг підіймається в славі!
PS|112|10|Це бачить безбожний та гнівається, скрегоче зубами своїми та тане... Бажання безбожних загине!
PS|113|1|Алілуя! Хваліте, Господні раби, хваліть ім'я Господа!
PS|113|2|Нехай буде благословенне Господнє ім'я відтепер і навіки!
PS|113|3|Від сходу сонця аж до заходу його прославляйте Господнє ім'я!
PS|113|4|Господь підіймається над усі народи, Його слава понад небеса!
PS|113|5|Хто подібний до Господа, нашого Бога, що мешкає на висоті,
PS|113|6|та знижується, щоб побачити те, що на небесах і на землі?
PS|113|7|Бідаря Він підводить із пороху, зо сміття підіймає нужденного,
PS|113|8|щоб його посадити з вельможними, з вельможними люду Його!
PS|113|9|Він неплідну в домі садовить за радісну матір дітей! Алілуя!
PS|114|1|Як виходив ізраїль з Єгипту, від народу чужого дім Яковів,
PS|114|2|Юда став за святиню Йому, а ізраїль Його пануванням!
PS|114|3|Побачило море все це і побігло, Йордан повернувся назад!
PS|114|4|Гори скакали, немов баранці, а пагірки немов ті ягнята!
PS|114|5|Що тобі, море, що ти втікаєш? Йордане, що ти повернувся назад?
PS|114|6|Чого скачете, гори, немов баранці, а пагірки мов ті ягнята?
PS|114|7|Тремти, земле, перед Господнім лицем, перед лицем Бога Якова,
PS|114|8|що скелю обертає в озеро водне, а кремінь на водне джерело!
PS|115|1|(114-9) Не нам, Господи, не нам, але Йменню Своєму дай славу за милість Твою, за правду Твою!
PS|115|2|(114-10) Пощо мають казати народи: Де ж то їхній Бог?
PS|115|3|(114-11) А Бог наш на небі, усе, що хотів, учинив.
PS|115|4|(114-12) Їхні божки срібло й золото, діло рук людських:
PS|115|5|(114-13) вони мають уста й не говорять, очі мають вони і не бачать,
PS|115|6|(114-14) мають уші й не чують, мають носа й без нюху,
PS|115|7|(114-15) мають руки та не дотикаються, мають ноги й не ходять, своїм горлом вони не говорять!
PS|115|8|(114-16) Нехай стануть такі, як вони, ті, хто їх виробляє, усі, хто надію на них покладає!
PS|115|9|(114-17) ізраїлю, надію складай лиш на Господа: Він їм поміч та щит їм!
PS|115|10|(114-18) Аароновий доме, надійтесь на Господа: Він їм поміч та щит їм!
PS|115|11|(114-19) Ті, що Господа боїтеся, надійтесь на Господа: Він їм поміч та щит їм!
PS|115|12|(114-20) Господь пам'ятає про нас, нехай поблагословить! Нехай поблагословить ізраїлів дім, нехай поблагословить Він дім Ааронів!
PS|115|13|(114-21) Нехай поблагословить Він тих, хто має до Господа страх, малих та великих!
PS|115|14|(114-22) Нехай вас розмножить Господь, вас і ваших дітей!
PS|115|15|(114-23) Благословенні ви в Господа, що вчинив небо й землю!
PS|115|16|(114-24) Небо, небо для Господа, а землю віддав синам людським!
PS|115|17|(114-25) Не мертві хвалитимуть Господа, ані ті всі, хто сходить у місце мовчання,
PS|115|18|(114-26) а ми благословлятимемо Господа відтепер й аж навіки! Алілуя!
PS|116|1|(115-1) Люблю я Господа, бо Він почув голос мій у благаннях моїх,
PS|116|2|(115-2) бо Він нахилив Своє ухо до мене, і я кликатиму в свої дні!
PS|116|3|(115-3) Болі смерти мене оточили і знайшли мене муки шеолу, нещастя та смуток знайшов я!
PS|116|4|(115-4) А я в ім'я Господа кличу: О Господи, визволи ж душу мою!
PS|116|5|(115-5) Господь милостивий та справедливий, і наш Бог милосердний!
PS|116|6|(115-6) Пильнує Господь недосвідчених, став я нужденний, та Він допоможе мені!
PS|116|7|(115-7) Вернися, о душе моя, до свого відпочинку, бо Господь робить добре тобі,
PS|116|8|(115-8) бо від смерти Ти визволив душу мою, від сльози моє око, ногу мою від спотикання.
PS|116|9|(115-9) Я ходитиму перед обличчям Господнім на землях живих!
PS|116|10|(116-1) Я вірив, коли говорив: Я сильно пригнічений!
PS|116|11|(116-2) Я сказав був у поспіху: Кожна людина говорить неправду!
PS|116|12|(116-3) Чим я відплачу Господеві за всі добродійства Його на мені?
PS|116|13|(116-4) Я чашу спасіння прийму, і прикличу Господнє ім'я!
PS|116|14|(116-5) Присяги свої Господеві я виконаю перед усім народом Його!
PS|116|15|(116-6) Дорога в очах Господа смерть богобійних Його!
PS|116|16|(116-7) О Господи, я бо Твій раб, я Твій раб, син Твоєї невільниці, Ти кайдани мої розв'язав!
PS|116|17|(116-8) Я жертву подяки Тобі принесу, і Господнім ім'ям буду кликати!
PS|116|18|(116-9) Присяги свої Господеві я виконаю перед усім народом Його,
PS|116|19|(116-10) на подвір'ях Господнього дому, посеред тебе, о Єрусалиме! Алілуя!
PS|117|1|Хваліть Господа, всі племена, прославляйте Його, всі народи,
PS|117|2|бо зміцнилось Його милосердя над нами, а правда Господня навіки! Алілуя!
PS|118|1|Дякуйте Господу, добрий бо Він, бо навіки Його милосердя!
PS|118|2|Нехай скаже ізраїль, бо навіки Його милосердя!
PS|118|3|Нехай скаже дім Ааронів, бо навіки Його милосердя!
PS|118|4|Нехай скажуть ті, хто боїться Господа, бо навіки Його милосердя!
PS|118|5|У тісноті я кликав до Господа, і простором озвався до мене Господь!
PS|118|6|Зо мною Господь не боюся нікого, що зробить людина мені?
PS|118|7|Господь серед тих, що мені помагають, і побачу загибіль своїх ненависників.
PS|118|8|Краще вдаватись до Господа, ніж надіятися на людину,
PS|118|9|краще вдаватись до Господа, ніж надіятися на вельможних!
PS|118|10|Всі народи мене оточили, я ж Господнім ім'ям їх понищив!
PS|118|11|Оточили мене й обступили мене, я ж Господнім ім'ям їх понищив!
PS|118|12|Оточили мене немов бджоли, та погасли вони, як терновий огонь, я бо Господнім ім'ям їх понищив!
PS|118|13|Дошкульно попхнув ти мене на падіння, та Господь спас мене!
PS|118|14|Господь моя сила та пісня, і став Він спасінням мені!
PS|118|15|Голос співу й спасіння в наметах між праведників: Господня правиця виконує чуда!
PS|118|16|Правиця Господня підноситься, правиця Господня виконує чуда!
PS|118|17|Не помру, але житиму, і буду звіщати про чини Господні!
PS|118|18|Покарати мене покарав був Господь, та смерти мені не завдав.
PS|118|19|Відчиніте мені брами правди, я ними ввійду, буду славити Господа!
PS|118|20|Це брама Господня, праведники в неї входять.
PS|118|21|Я буду хвалити Тебе, бо озвався до мене, і став Ти спасінням мені!
PS|118|22|Камінь, що його будівничі відкинули, той наріжним став каменем,
PS|118|23|від Господа сталося це, і дивне воно в очах наших!
PS|118|24|Це день, що його створив Господь, радіймо та тішмося в нім!
PS|118|25|Просимо, Господи, спаси! Просимо, Господи, пощасти!
PS|118|26|Благословен, хто гряде у Господнє ім'я! Благословляємо вас із Господнього дому!
PS|118|27|Господь Бог, і засяяв Він нам. Прив'яжіте святковую жертву шнурами аж до наріжників жертівника!
PS|118|28|Ти мій Бог, і я буду Тебе прославляти, мій Боже, я буду Тебе величати!
PS|118|29|Дякуйте Господу, добрий бо Він, бо навіки Його милосердя!
PS|119|1|Блаженні непорочні в дорозі, що ходять Законом Господнім!
PS|119|2|Блаженні, хто держить свідоцтва Його, хто шукає Його всім серцем,
PS|119|3|і хто кривди не робить, хто ходить путями Його!
PS|119|4|Ти видав накази Свої, щоб виконувати пильно.
PS|119|5|Коли б же дороги мої були певні, щоб держатись Твоїх постанов,
PS|119|6|не буду тоді засоромлений я, як буду дивитись на всі Твої заповіді!
PS|119|7|Щирим серцем я буду Тебе прославляти, як навчуся законів Твоїх справедливих.
PS|119|8|Я буду держатись Твоїх постанов, не кидай же зовсім мене!
PS|119|9|Чим додержить юнак у чистоті свою стежку? Як держатиметься Твоїх слів!
PS|119|10|Цілим серцем своїм я шукаю Тебе, не дай же мені заблудитися від Твоїх заповідей!
PS|119|11|Я в серці своїм заховав Твоє слово, щоб мені не грішити проти Тебе.
PS|119|12|Благословен єси, Господи, навчи мене постанов Своїх!
PS|119|13|Устами своїми я розповідаю про всі присуди уст Твоїх.
PS|119|14|З дороги свідоцтв Твоїх радію я, як маєтком великим.
PS|119|15|Про накази Твої розмовлятиму я, і на стежки Твої буду дивитись.
PS|119|16|Я буду радіти Твоїми постановами, слова Твого не забуду!
PS|119|17|Своєму рабові пощасти, щоб я жив, і я буду держатися слова Твого!
PS|119|18|Відкрий мої очі, і хай чуда Закону Твого я побачу!
PS|119|19|На землі я приходько, Своїх заповідей не ховай Ти від мене!
PS|119|20|Омліває душа моя з туги за Твоїми законами кожного часу...
PS|119|21|Насварив Ти проклятих отих гордунів, що вхиляються від Твоїх заповідей.
PS|119|22|Відверни Ти від мене зневагу та сором, бо держуся свідоцтв Твоїх я!
PS|119|23|Теж вельможі сидять та на мене змовляються, та Твій раб про постанови Твої розмовляє,
PS|119|24|і свідоцтва Твої то потіха моя, то для мене дорадники!
PS|119|25|Душа моя гнеться до пороху, за словом Своїм оживи Ти мене!
PS|119|26|Про дороги свої я казав, і почув Ти мене, навчи Ти мене постанов Своїх!
PS|119|27|Дай мені розуміти дорогу наказів Твоїх, і про чуда Твої я звіщатиму.
PS|119|28|Розпливає зо смутку душа моя, постав мене згідно зо словом Своїм!
PS|119|29|Дорогу неправди від мене відсунь, і дай мені з ласки Своєї Закона!
PS|119|30|Я вибрав путь правди, закони Твої біля себе поставив.
PS|119|31|До свідоцтв Твоїх я приєднався, Господи, не посором же мене!
PS|119|32|Буду бігти шляхом Твоїх заповідей, бо пошириш Ти серце моє.
PS|119|33|Путь Своїх постанов покажи мені, Господи, і я буду держатись її до кінця!
PS|119|34|Дай мені зрозуміти, і нехай я держуся Закону Твого, і всім серцем я буду триматись його!
PS|119|35|Провадь мене стежкою Твоїх заповідей, бо в ній я знайшов уподобу.
PS|119|36|Серце моє прихили до свідоцтв Твоїх, а не до користи.
PS|119|37|Відверни мої очі, щоб марноти не бачили, на дорозі Своїй оживи Ти мене!
PS|119|38|Для Свого раба сповни слово Своє, що на страх Твій воно.
PS|119|39|Відверни Ти від мене зневагу, якої боюся, бо добрі закони Твої.
PS|119|40|Ось я прагну наказів Твоїх, оживи мене правдою Своєю!
PS|119|41|і хай зійде на мене, о Господи, милість Твоя, спасіння Твоє, згідно з словом Твоїм,
PS|119|42|і нехай відповім я тому, хто словом ганьбить мене, бо надіюсь на слово Твоє!
PS|119|43|і не відіймай з моїх уст слова правди ніколи, бо я жду Твоїх присудів!
PS|119|44|А я буду держатися завжди Закону Твого, на вічні віки!
PS|119|45|і буду ходити в широкості, бо наказів Твоїх я шукаю.
PS|119|46|і буду я перед царями звіщати про свідоцтва Твої, й не зазнаю я сорому!
PS|119|47|і буду я розкошувати Твоїми заповідями, бо їх полюбив,
PS|119|48|і я руки свої простягну до Твоїх заповідей, бо їх полюбив, і буду роздумувати про Твої постанови!
PS|119|49|Пам'ятай про те слово Своєму рабові, що його наказав Ти чекати мені.
PS|119|50|Це розрада моя в моїм горі, як слово Твоє оживляє мене.
PS|119|51|Гордуни насміхалися з мене занадто, та я не відступив від Закону Твого!
PS|119|52|Твої присуди я пам'ятаю відвіку, о Господи, і радію!
PS|119|53|Буря мене обгорнула через нечестивих, що Закона Твого опускають!
PS|119|54|Співи для мене Твої постанови у домі моєї мандрівки.
PS|119|55|Я вночі пам'ятаю ім'я Твоє, Господи, і держуся Закону Твого!
PS|119|56|Оце сталось мені, бо наказів Твоїх я держуся.
PS|119|57|Я сказав: Моя доля, о Господи, щоб держатись мені Твоїх слів.
PS|119|58|Я благаю Тебе цілим серцем: Учини мені милість за словом Своїм!
PS|119|59|Я розважив дороги свої, й до свідоцтв Твоїх ноги свої звернув.
PS|119|60|Я спішу й не барюся виконувати Твої заповіді.
PS|119|61|Тенета безбожних мене оточили, та я не забув про Закона Твого.
PS|119|62|Опівночі встаю я, щоб скласти подяку Тобі за присуди правди Твоєї.
PS|119|63|Я приятель всім, хто боїться Тебе, й хто накази Твої береже!
PS|119|64|Милосердя Твого, о Господи, повна земля, навчи Ти мене Своїх постанов!
PS|119|65|Ти з рабом Своїм добре зробив, Господи, за словом Своїм.
PS|119|66|Навчи мене доброго розуму та познавання, бо в заповіді Твої вірую я!
PS|119|67|Доки я не страждав, блудив був, та тепер я держусь Твого слова.
PS|119|68|Ти добрий, і чиниш добро, навчи Ти мене Своїх постанов!
PS|119|69|Гордуни вимишляють на мене неправду, а я цілим серцем держуся наказів Твоїх.
PS|119|70|Зробилось нечуле, як лій, їхнє серце, а я розкошую з Закону Твого.
PS|119|71|Добре мені, що я змучений був, щоб навчитися Твоїх постанов!
PS|119|72|Ліпший для мене Закон Твоїх уст, аніж тисячі золота й срібла.
PS|119|73|Руки Твої створили мене й збудували мене, подай мені розуму, й хай я навчусь Твоїх заповідей!
PS|119|74|Хто боїться Тебе, ті побачать мене та й зрадіють, бо я Твого слова чекаю!
PS|119|75|Знаю я, Господи, що справедливі були Твої присуди, і справедливо мене понижав Ти.
PS|119|76|Нехай буде милість Твоя на розраду мені, за словом Твоїм до Свого раба.
PS|119|77|Нехай зійде на мене Твоє милосердя, й я житиму, бо Закон Твій розрада моя.
PS|119|78|Нехай гордуни посоромлені будуть, бо робили нечесно, а я буду роздумувати про накази Твої.
PS|119|79|До мене повернуться ті, хто боїться Тебе, і пізнають свідоцтва Твої.
PS|119|80|Нехай серце моє буде чисте в Твоїх постановах, щоб я не посоромився!
PS|119|81|Душа моя слабне від туги за спасінням Твоїм, чекаю я слова Твого!
PS|119|82|За словом Твоїм гаснуть очі мої та питають: Коли Ти потішиш мене?...
PS|119|83|Хоч я став, як той міх у диму, та Твоїх постанов не забув.
PS|119|84|Скільки днів для Твого раба? Коли присуда зробиш моїм переслідникам?
PS|119|85|Гордуни покопали були мені ями, що не за Законом Твоїм.
PS|119|86|Усі Твої заповіді справедливі; неправдиво мене переслідують, допоможи Ти мені!
PS|119|87|Малощо не погубили мене на землі, та я не покинув наказів Твоїх!
PS|119|88|Оживи Ти мене за Своїм милосердям, і я буду триматися свідчення уст Твоїх!
PS|119|89|Навіки, о Господи, слово Твоє в небесах пробуває.
PS|119|90|З роду в рід Твоя правда; Ти землю поставив і стала вона,
PS|119|91|усі за Твоїми судами сьогодні стоять, бо раби Твої всі.
PS|119|92|Коли б не Закон Твій, розрада моя, то я був би загинув в недолі своїй!
PS|119|93|Я повік не забуду наказів Твоїх, бо Ти ними мене оживляєш.
PS|119|94|Твій я, спаси Ти мене, бо наказів Твоїх я шукаю!
PS|119|95|Чекають безбожні забити мене, а я про свідоцтва Твої розважаю.
PS|119|96|Я бачив кінець усього досконалого, але Твоя заповідь вельми широка!
PS|119|97|Як я кохаю Закона Твого, цілий день він розмова моя!
PS|119|98|Твоя заповідь робить мудрішим мене від моїх ворогів, вона бо навіки моя!
PS|119|99|Я став розумніший за всіх своїх учителів, бо свідоцтва Твої то розмова моя!
PS|119|100|Став я мудріший за старших, бо держуся наказів Твоїх!
PS|119|101|Я від кожної злої дороги повстримую ноги свої, щоб держатися слова Твого.
PS|119|102|Я не ухиляюся від Твоїх присудів, Ти бо навчаєш мене.
PS|119|103|Яке то солодке слово Твоє для мого піднебіння, солодше від меду воно моїм устам!
PS|119|104|Від наказів Твоїх я мудріший стаю, тому то ненавиджу всяку дорогу неправди!
PS|119|105|Для моєї ноги Твоє слово світильник, то світло для стежки моєї.
PS|119|106|Я присяг і дотримаю, що буду держатися присудів правди Твоєї.
PS|119|107|Перемучений я аж занадто, за словом Своїм оживи мене, Господи!
PS|119|108|Хай же будуть приємні Тобі жертви уст моїх, Господи, і навчи Ти мене Своїх присудів!
PS|119|109|У небезпеці душа моя завжди, але я Закону Твого не забув.
PS|119|110|Безбожні поставили пастку на мене, та я не зблудив від наказів Твоїх.
PS|119|111|Я навіки свідоцтва Твої вспадкував, бо вони радість серця мого.
PS|119|112|Я серце своє нахилив, щоб чинити Твої постанови, повік, до кінця.
PS|119|113|Сумнівне ненавиджу я, а Закона Твого покохав.
PS|119|114|Ти моя охорона та щит мій, чекаю я слова Твого.
PS|119|115|Відступіться від мене, злочинці, і я буду держатися заповідей мого Бога!
PS|119|116|За словом Своїм підіпри Ти мене, і я житиму, і в надії моїй не завдай мені сорому!
PS|119|117|Підкріпи Ти мене і спасуся, і я буду дивитися завжди в Твої постанови!
PS|119|118|Ти погорджуєш усіма, хто від Твоїх постанов відступає, бо хитрощі їхні неправда.
PS|119|119|Всіх безбожних землі відкидаєш, як жужель, тому покохав я свідоцтва Твої.
PS|119|120|Зо страху Твого моє тіло тремтить, й я боюсь Твоїх присудів!
PS|119|121|Я право та правду чиню, щоб мене не віддав Ти моїм переслідникам.
PS|119|122|Поручи Ти на добре Свого раба, щоб мене гордуни не гнобили.
PS|119|123|Гаснуть очі мої за спасінням Твоїм та за словом правди Твоєї.
PS|119|124|Учини ж Ти Своєму рабові за Своїм милосердям, і навчи Ти мене Своїх постанов!
PS|119|125|Я раб Твій, і зроби мене мудрим, і свідоцтва Твої буду знати!
PS|119|126|Це для Господа час, щоб діяти: Закона Твого уневажнили.
PS|119|127|Тому я люблю Твої заповіді більш від золота й щирого золота.
PS|119|128|Тому всі накази Твої уважаю за слушні, а кожну дорогу неправди ненавиджу!
PS|119|129|Чудові свідоцтва Твої, тому то душа моя держиться їх.
PS|119|130|Вхід у слова Твої світло дає, недосвідчених мудрими робить.
PS|119|131|Я уста свої розкриваю й повітря ковтаю, бо чую жадобу до Твоїх заповідей.
PS|119|132|Обернися до мене та будь милостивий мені, Як чиниш Ти тим, хто кохає імення Твоє.
PS|119|133|Своїм словом зміцни мої кроки, і не дай панувати надо мною ніякому прогріхові.
PS|119|134|Від людського утиску визволь мене, і нехай я держуся наказів Твоїх!
PS|119|135|Хай засяє лице Твоє на Твого раба, і навчи Ти мене уставів Своїх!
PS|119|136|Пливуть водні потоки з очей моїх, бо Твого Закону не додержують...
PS|119|137|Ти праведний, Господи, і прямі Твої присуди,
PS|119|138|бо Ти наказав справедливі свідоцтва Свої й щиру правду!
PS|119|139|Нищить мене моя ревність, бо мої вороги позабували слова Твої.
PS|119|140|Вельми очищене слово Твоє, і Твій раб його любить.
PS|119|141|Я малий і погорджений, та не забуваю наказів Твоїх.
PS|119|142|Правда Твоя правда вічна, а Закон Твій то істина.
PS|119|143|Недоля та утиск мене обгорнули, але Твої заповіді моя розкіш!
PS|119|144|Правда свідоцтв Твоїх вічна, подай мені розуму, й буду я жити!
PS|119|145|Цілим серцем я кличу: почуй мене, Господи, і я буду держатись уставів Твоїх!
PS|119|146|Я кличу до Тебе, спаси Ти мене, і я буду держатись свідоцтв Твоїх!
PS|119|147|Світанок я випередив та й вже кличу, Твого слова чекаю.
PS|119|148|Мої очі сторожі нічні випереджують, щоб про слово Твоє розмовляти.
PS|119|149|Почуй же мій голос з Свого милосердя, о Господи, оживи Ти мене з Свого присуду!
PS|119|150|Наближаться ті, що за чином ганебним ганяють, від Закону Твого далекі,
PS|119|151|та близький Ти, о Господи, а всі Твої заповіді справедливість!
PS|119|152|Віддавна я знаю свідоцтва Твої, бо навіки Ти їх заклав!
PS|119|153|Подивись на недолю мою та мене порятуй, бо я не забуваю Закону Твого!
PS|119|154|Вступися за справу мою й мене визволи, за словом Своїм оживи Ти мене!
PS|119|155|Від безбожних спасіння далеке, бо вони не шукають Твоїх постанов.
PS|119|156|Велике Твоє милосердя, о Господи, оживи Ти мене з Свого присуду!
PS|119|157|Багато моїх переслідників та ворогів моїх, але від свідоцтв Твоїх не відхиляюсь!
PS|119|158|Бачив я зрадників й бридився ними, бо не держать вони Твого слова.
PS|119|159|Подивися: люблю я накази Твої, за милосердям Своїм оживи мене, Господи!
PS|119|160|Правда підвалина слова Твого, а присуди правди Твоєї навіки.
PS|119|161|Безневинно вельможі мене переслідують, та серце моє Твого слова боїться.
PS|119|162|Радію я словом Твоїм, ніби здобич велику знайшов.
PS|119|163|Я неправду ненавиджу й бриджуся нею, покохав я Закона Твого!
PS|119|164|Сім раз денно я славлю Тебе через присуди правди Твоєї.
PS|119|165|Мир великий для тих, хто кохає Закона Твого, і не мають вони спотикання.
PS|119|166|На спасіння Твоє я надіюся, Господи, і Твої заповіді виконую.
PS|119|167|Душа моя держить свідоцтва Твої, і я сильно люблю їх.
PS|119|168|Я держуся наказів Твоїх та свідоцтв Твоїх, бо перед Тобою мої всі дороги!
PS|119|169|Благання моє хай наблизиться перед лице Твоє, Господи, за словом Своїм подай мені розуму!
PS|119|170|Нехай прийде молитва моя перед лице Твоє, за словом Своїм мене визволь!
PS|119|171|Нехай уста мої вимовляють хвалу, бо уставів Своїх Ти навчаєш мене.
PS|119|172|Хай язик мій звіщатиме слово Твоє, бо всі Твої заповіді справедливість.
PS|119|173|Нехай буде рука Твоя в поміч мені, бо я вибрав накази Твої.
PS|119|174|Я прагну спасіння Твого, о Господи, а Закон Твій то розкіш моя!
PS|119|175|Хай душа моя буде жива, і хай славить Тебе, а Твій присуд нехай допоможе мені!
PS|119|176|Я блукаю, немов та овечка загублена, пошукай же Свого раба, бо я не забув Твоїх заповідей!...
PS|120|1|Пісня прочан. Я кликав до Господа в горі своїм, і Він мене вислухав,
PS|120|2|Господи, визволь же душу мою від губи неправдивої, від язика зрадливого!
PS|120|3|Що Тобі дасть, або що для Тебе додасть лукавий язик?
PS|120|4|Загострені стріли потужного із ялівцевим вугіллям!
PS|120|5|Горе мені, що замешкую в Мешеху, що живу із шатрами Кедару!
PS|120|6|Довго душа моя перебувала собі разом з тими, хто ненавидить мир:
PS|120|7|я за мир, та коли говорю, то вони за війну!
PS|121|1|Пісня прочан. Свої очі я зводжу на гори, звідки прийде мені допомога,
PS|121|2|мені допомога від Господа, що вчинив небо й землю!
PS|121|3|Він не дасть захитатись нозі твоїй, не здрімає твій Сторож:
PS|121|4|оце не дрімає й не спить Сторож ізраїлів!
PS|121|5|Господь то твій Сторож, Господь твоя тінь при правиці твоїй,
PS|121|6|удень сонце не вдарить тебе, ані місяць вночі!
PS|121|7|Господь стерегтиме тебе від усякого зла, стерегтиме Він душу твою,
PS|121|8|Господь стерегтиме твій вихід та вхід відтепер аж навіки!
PS|122|1|Пісня прочан. Давидова. Я радів, як казали мені: Ходімо до дому Господнього!
PS|122|2|Ноги наші стояли в воротях Твоїх, Єрусалиме.
PS|122|3|Єрусалиме, збудований ти як те місто, що злучене разом,
PS|122|4|куди сходять племена, племена Господні, щоб свідчити ізраїлеві, щоб іменню Господньому дякувати!
PS|122|5|Бо то там на престолах для суду сидять, на престолах дому Давидового.
PS|122|6|Миру бажайте для Єрусалиму: Нехай будуть безпечні, хто любить тебе!
PS|122|7|Нехай буде мир у твоїх передмур'ях, безпека в палатах твоїх!
PS|122|8|Ради братті моєї та друзів моїх я буду казати: Мир тобі!
PS|122|9|Ради дому Господа, нашого Бога, я буду шукати для тебе добра!
PS|123|1|Пісня прочан. Свої очі я зводжу до Тебе, що на небесах пробуваєш!
PS|123|2|Ото бо, як очі рабів до руки їх панів, як очі невільниці до руки її пані, отак наші очі до Господа, нашого Бога, аж поки не змилується Він над нами!
PS|123|3|Помилуй нас, Господи, помилуй нас, бо погорди ми досить наситились!
PS|123|4|Душа наша наситилась досить собі: від безпечних наруги, від пишних погорди!...
PS|124|1|Пісня прочан. Давидова. Коли б не Господь, що був з нами нехай но ізраїль повість!
PS|124|2|коли б не Господь, що був з нами, як повстала була на нас людина,
PS|124|3|то нас поковтали б живцем, коли розпалився на нас їхній гнів,
PS|124|4|то нас позаливала б вода, душу нашу потік перейшов би,
PS|124|5|душу нашу тоді перейшла б та бурхлива вода!
PS|124|6|Благословенний Господь, що не дав нас на здобич для їхніх зубів!
PS|124|7|Душа наша, як птах, урятувалась із сільця птахоловів, сільце розірвалось, а ми врятувались!
PS|124|8|Наша поміч ув імені Господа, що вчинив небо й землю!
PS|125|1|Пісня прочан. Ті, хто надію складає на Господа, вони як Сіонська гора, яка не захитається, яка буде стояти повік!
PS|125|2|Єрусалим, гори круг нього, а Господь круг народу Свого відтепер й аж навіки!
PS|125|3|Не спочине бо берло нечестя на долі тих праведних, щоб праведні не простягли своїх рук до неправди.
PS|125|4|Зроби ж, Господи, добре для добрих, та для простосердих!
PS|125|5|Тих же, що збочують на свої манівці, нехай їх провадить Господь разом із беззаконцями! Мир на ізраїля!
PS|126|1|Пісня прочан. Як вертався Господь із полоном Сіону, то були ми немов би у сні...
PS|126|2|Наші уста тоді були повні веселощів, а язик наш співання! Казали тоді між народами: Велике вчинив Господь з ними!
PS|126|3|Велике вчинив Господь з нами, були радісні ми!
PS|126|4|Вернися ж із нашим полоном, о Господи, немов ті джерела, на південь!
PS|126|5|Хто сіє з слізьми, зо співом той жне:
PS|126|6|все ходить та плаче, хто носить торбину насіння на посів, та вернеться з співом, хто носить снопи свої!
PS|127|1|Пісня прочан. Соломонова. Коли дому Господь не будує, даремно працюють його будівничі при ньому! Коли міста Господь не пильнує, даремно сторожа чуває!
PS|127|2|Даремно вам рано вставати, допізна сидіти, їсти хліб загорьований, Він і в спанні подасть другові Своєму!
PS|127|3|Діти спадщина Господнє, плід утроби нагорода!
PS|127|4|Як стріли в руках того велетня, так і сини молоді:
PS|127|5|блаженний той муж, що сагайдака свого ними наповнив, не будуть такі посоромлені, коли в брамі вони говоритимуть із ворогами!
PS|128|1|Пісня прочан. Блажен кожен, хто боїться Господа, хто ходить путями Його!
PS|128|2|Коли труд своїх рук будеш їсти, блажен ти, і добре тобі!
PS|128|3|Твоя жінка в кутах твого дому як та виноградина плідна, твої діти навколо твого стола немов саджанці ті оливкові!
PS|128|4|Оце так буде поблагословлений муж, що боїться він Господа!
PS|128|5|Нехай поблагословить тебе Господь із Сіону, і побачиш добро Єрусалиму по всі дні свого життя,
PS|128|6|і побачиш онуків своїх! Мир на ізраїля!
PS|129|1|Пісня прочан. Багато гнобили мене від юнацтва мого, нехай но ізраїль повість!
PS|129|2|Багато гнобили мене від юнацтва мого, та мене не подужали!
PS|129|3|Орали були на хребті моїм плугатарі, поклали вони довгі борозни,
PS|129|4|та Господь справедливий, Він шнури безбожних порвав!
PS|129|5|Нехай посоромлені будуть, і хай повідступають назад усі ті, хто Сіона ненавидить!
PS|129|6|Бодай стали вони, як трава на дахах, що всихає вона, поки виросте,
PS|129|7|що нею жмені своєї жнець не наповнить, ані оберемка свого в'язальник,
PS|129|8|і не скаже прохожий до них: Благословення Господнє на вас, благословляємо вас ім'ям Господа!
PS|130|1|Пісня прочан. З глибини я взиваю до Тебе, о Господи:
PS|130|2|Господи, почуй же мій голос! Нехай уші Твої будуть чулі на голос благання мого!
PS|130|3|Якщо, Господи, будеш зважати на беззаконня, хто встоїть, Владико?
PS|130|4|Бо в Тебе пробачення, щоб боятись Тебе...
PS|130|5|Я надіюсь на Господа, має надію душа моя, і на слово Його я вповаю.
PS|130|6|Виглядає душа моя Господа більш, ніж поранку сторожа, що до ранку вона стереже.
PS|130|7|Хай надію складає ізраїль на Господа, бо з Господом милість, і велике визволення з Ним,
PS|130|8|і ізраїля визволить Він від усіх його прогріхів!
PS|131|1|Пісня прочан. Давидова. Господи, серце моє не пишнилось, і очі мої не підносились, і я не ганявсь за речами, що більші й дивніші над мене!
PS|131|2|Таж я втихомирював і заспокоював душу свою, як дитя, від перс мами своєї відлучене, як дитина відлучена в мене душа моя!
PS|131|3|Хай надію складає ізраїль на Господа відтепер аж навіки!
PS|132|1|Пісня прочан. Згадай, Господи, про Давида, про всі його муки,
PS|132|2|що клявсь Господеві, присягався був Сильному Якова:
PS|132|3|Не ввійду я в намет свого дому, не зійду я на ложе постелі своєї,
PS|132|4|не дам сну своїм очам, дрімання повікам своїм,
PS|132|5|аж поки не знайду я для Господа місця, місця перебування для Сильного Якова!
PS|132|6|Ось ми чули про Нього в Ефрафі, на Яарських полях ми знайшли Його.
PS|132|7|Увійдім же в мешкання Його, поклонімось підніжкові ніг Його!
PS|132|8|Встань же Господи, йди до Свого відпочинку, Ти й ковчег сили Твоєї!
PS|132|9|Священики Твої хай зодягнуться в правду, і будуть співати Твої богобійні!
PS|132|10|Ради Давида, Свого раба, не відвертай лиця від Свого помазанця.
PS|132|11|Господь присягнув був Давидові правду, і не відступить від неї: Від плоду утроби твоєї Я посаджу на престолі твоїм!
PS|132|12|Якщо будуть синове твої пильнувати Мого заповіта й свідоцтва Мого, що його Я навчатиму їх, то й сини їхні на вічні віки будуть сидіти на троні твоїм!
PS|132|13|Бо вибрав Сіона Господь, уподобав його на оселю Собі:
PS|132|14|То місце Мого відпочинку на вічні віки, пробуватиму тут, бо його уподобав,
PS|132|15|поживу його щедро благословлю, і хлібом убогих його нагодую!
PS|132|16|Священиків його зодягну у спасіння, а його богобійні співатимуть радісно.
PS|132|17|Я там вирощу рога Давидового, для Свого помазанця вготую світильника,
PS|132|18|ворогів його соромом позодягаю, а на ньому корона його буде сяяти!
PS|133|1|Пісня прочан. Давидова. Оце яке добре та гарне яке, щоб жити братам однокупно!
PS|133|2|Воно як та добра олива на голову, що спливає на бороду, Ааронову бороду, що спливає на кінці одежі його!
PS|133|3|Воно як хермонська роса, що спадає на гори Сіону, бо там наказав Господь благословення, повіквічне життя!
PS|134|1|Пісня прочан. Поблагословіть оце Господа, всі раби Господні, що по ночах у домі Господньому ви стоїте!
PS|134|2|Ваші руки здійміть до святині, і Господа благословіть!
PS|134|3|Нехай поблагословить тебе із Сіону Господь, що вчинив небо й землю!
PS|135|1|Алілуя! Хваліте Господнє ім'я, хваліте, Господні раби,
PS|135|2|що стоїте в домі Господньому, на подвір'ях дому нашого Бога!
PS|135|3|Хваліть Господа, бо добрий Господь, співайте іменню Його, бо приємне воно,
PS|135|4|бо вибрав Господь собі Якова, ізраїля на власність Свою!
PS|135|5|Знаю бо я, що Господь і Владика наш більший від богів усіх!
PS|135|6|Все, що хоче Господь, те Він чинить на небі та на землі, на морях та по всяких глибинах!
PS|135|7|Підіймає Він хмари від краю землі, блискавиці вчинив для дощу, випроваджує вітер з запасів Своїх.
PS|135|8|Він позабивав перворідних Єгипту, від людини аж до скотини.
PS|135|9|Він послав між Єгипет ознаки та чуда, на фараона і на рабів всіх його.
PS|135|10|Він уразив багато народів, і потужних царів повбивав:
PS|135|11|Сигона, царя амореян, і Оґа, Башану царя, та всіх ханаанських царів.
PS|135|12|і Він дав їхню землю спадщиною, на спадок ізраїлеві, Своєму народові.
PS|135|13|Господи, Ймення Твоє віковічне, Господи, пам'ять Твоя з роду в рід!
PS|135|14|Бо буде судити Господь Свій народ, та змилосердиться Він над Своїми рабами.
PS|135|15|Божки людів то срібло та золото, діло рук людських:
PS|135|16|вони мають уста й не говорять, очі мають вони і не бачать,
PS|135|17|мають уші й не чують, в їхніх устах нема віддиху!
PS|135|18|Нехай стануть такі, як вони, ті, хто їх виробляє, усі, хто надію на них покладає!
PS|135|19|Доме ізраїлів, благословіть Господа! Аароновий доме, благословіть Господа!
PS|135|20|Доме Левіїв, благословіть Господа! Хто боїться Господа, благословіть Господа!
PS|135|21|Благословенний Господь від Сіону, що мешкає в Єрусалимі! Алілуя!
PS|136|1|Дякуйте Господу, добрий бо Він, бо навіки Його милосердя!
PS|136|2|Дякуйте Богу богів, бо навіки Його милосердя!
PS|136|3|Дякуйте Владиці владик, бо навіки Його милосердя!
PS|136|4|Тому, хто чуда великі Єдиний вчиняє, бо навіки Його милосердя!
PS|136|5|Хто розумом небо вчинив, бо навіки Його милосердя!
PS|136|6|Хто землю простяг над водою, бо навіки Його милосердя!
PS|136|7|Хто світила великі вчинив, бо навіки Його милосердя!
PS|136|8|сонце, щоб вдень панувало воно, бо навіки Його милосердя!
PS|136|9|місяця й зорі, щоб вони панували вночі, бо навіки Його милосердя!
PS|136|10|Хто Єгипет побив був у їхніх перворідних, бо навіки Його милосердя!
PS|136|11|і ізраїля вивів з-між них, бо навіки Його милосердя!
PS|136|12|рукою міцною й раменом простягненим, бо навіки Його милосердя!
PS|136|13|Хто море Червоне розтяв на частини, бо навіки Його милосердя!
PS|136|14|і серед нього ізраїля перепровадив, бо навіки Його милосердя!
PS|136|15|і фараона та війська його вкинув у море Червоне, бо навіки Його милосердя!
PS|136|16|Хто провадив народ Свій в пустині, бо навіки Його милосердя!
PS|136|17|Хто великих царів повбивав, бо навіки Його милосердя!
PS|136|18|і потужних царів перебив, бо навіки Його милосердя!
PS|136|19|Сигона, царя амореян, бо навіки Його милосердя!
PS|136|20|і Оґа, Башану царя, бо навіки Його милосердя!
PS|136|21|і Хто землю їхню дав на спадщину, бо навіки Його милосердя!
PS|136|22|на спадок ізраїлеві, Своєму рабові, бо навіки Його милосердя!
PS|136|23|Хто про нас пам'ятав у пониженні нашім, бо навіки Його милосердя!
PS|136|24|і від ворогів наших визволив нас, бо навіки Його милосердя!
PS|136|25|Хто кожному тілові хліба дає, бо навіки Його милосердя!
PS|136|26|Дякуйте Богу небесному, бо навіки Його милосердя!
PS|137|1|Над річками Вавилонськими, там ми сиділи та й плакали, коли згадували про Сіона!
PS|137|2|На вербах у ньому повісили ми свої арфи,
PS|137|3|співу бо пісні від нас там жадали були поневолювачі наші, а веселощів наші мучителі: Заспівайте но нам із Сіонських пісень!
PS|137|4|Як же зможемо ми заспівати Господнюю пісню в землі чужинця?
PS|137|5|Якщо я забуду за тебе, о Єрусалиме, хай забуде за мене правиця моя!
PS|137|6|Нехай мій язик до мого піднебіння прилипне, якщо я не буду тебе пам'ятати, якщо не поставлю я Єрусалима над радість найвищу свою!...
PS|137|7|Пам'ятай же, о Господи, едомським синам про день Єрусалиму, як кричали вони: Руйнуйте, руйнуйте аж до підвалин його!...
PS|137|8|Вавилонськая дочко, що маєш і ти ограбована бути, блажен, хто заплатить тобі за твій чин, що ти нам заподіяла!
PS|137|9|Блажен, хто ухопить та порозбиває об скелю і твої немовлята!...
PS|138|1|Давидів. Прославляю Тебе цілим серцем своїм, перед богами співаю Тобі!
PS|138|2|Вклоняюсь до храму святого Твого, і славлю імення Твоє за Твоє милосердя й за правду Твою, бо звеличив Ти був над усе Своє Ймення та слово Своє!
PS|138|3|Удень, як взиваю, почуєш мене, підбадьорюєш силою душу мою!
PS|138|4|Усі земні царі прославлять Тебе, Господи, будуть, бо почують вони слово уст Твоїх,
PS|138|5|і будуть співати про Господні дороги, бо слава Господня велика,
PS|138|6|бо високий Господь, але бачить низького, а гордого Він пізнає іздалека!
PS|138|7|Якщо серед тісноти піду, Ти оживиш мене, на лютість моїх ворогів пошлеш руку Свою, і правиця Твоя допоможе мені,
PS|138|8|для мене Господь оце виконає! Твоя милість, о Господи, вічна, чинів Своєї руки не полиш!
PS|139|1|Для дириґетна хору. Псалом Давидів. Господи, випробував Ти мене та й пізнав,
PS|139|2|Ти знаєш сидіння моє та вставання моє, думку мою розумієш здалека.
PS|139|3|Дорогу мою та лежання моє виміряєш, і Ти всі путі мої знаєш,
PS|139|4|бо ще слова нема на моїм язиці, а вже, Господи, знаєш те все!
PS|139|5|Оточив Ти мене ззаду й спереду, і руку Свою надо мною поклав.
PS|139|6|Дивне знання над моє розуміння, високе воно, я його не подолаю!
PS|139|7|Куди я від Духа Твого піду, і куди я втечу від Твого лиця?
PS|139|8|Якщо я на небо зійду, то Ти там, або постелюся в шеолі ось Ти!
PS|139|9|Понесуся на крилах зірниці, спочину я на кінці моря,
PS|139|10|то рука Твоя й там попровадить мене, і мене буде тримати правиця Твоя!
PS|139|11|Коли б я сказав: Тільки темрява вкриє мене, і ніч світло для мене,
PS|139|12|то мене не закриє від Тебе і темрява, і ніч буде світити, як день, і темнота як світло!
PS|139|13|Бо Ти вчинив нирки мої, Ти виткав мене в утробі матері моєї,
PS|139|14|Прославляю Тебе, що я дивно утворений! Дивні діла Твої, і душа моя відає вельми про це!
PS|139|15|і кості мої не сховались від Тебе, бо я вчинений був в укритті, я витканий був у глибинах землі!
PS|139|16|Мого зародка бачили очі Твої, і до книги Твоєї записані всі мої члени та дні, що в них були вчинені, коли жодного з них не було...
PS|139|17|Які дорогі мені стали думки Твої, Боже, як побільшилося їх число,
PS|139|18|перелічую їх, численніші вони від піску! Як пробуджуюся, то я ще з Тобою.
PS|139|19|Якби, Боже, вразив Ти безбожника, а ви, кровожерці, відступітесь від мене!
PS|139|20|Вони називають підступно Тебе, Твої вороги на марноту пускаються!
PS|139|21|Отож, ненавиджу Твоїх ненависників, Господи, і Твоїх заколотників бриджусь:
PS|139|22|повною ненавистю я ненавиджу їх, вони стали мені ворогами!...
PS|139|23|Випробуй, Боже, мене, і пізнай моє серце, досліди Ти мене, і пізнай мої задуми,
PS|139|24|і побач, чи не йду я дорогою злою, і на вічну дорогу мене попровадь!
PS|140|1|Для дириґетна хору. Псалом Давидів. (140-2) Визволь мене від людини лихої, о Господи, бережи мене від насильника,
PS|140|2|(140-3) що в серці своїм замишляють злі речі, що війни щодня викликають!
PS|140|3|(140-4) Вони гострять свого язика, як той вуж, отрута гадюча під їхніми устами! Села.
PS|140|4|(140-5) Пильнуй мене, Господи, від рук нечестивого, бережи мене від насильника, що задумали стопи мої захитати...
PS|140|5|(140-6) Чванливі сховали на мене тенета та шнури, розтягли свою сітку при стежці, сільця розмістили на мене! Села.
PS|140|6|(140-7) Я сказав Господеві: Ти Бог мій, почуй же, о Господи, голос благання мого!
PS|140|7|(140-8) Господи, Владико мій, сило мого спасіння, що в день бою покрив мою голову,
PS|140|8|(140-9) не виконай, Господи, бажань безбожного, не здійсни його задуму! Села.
PS|140|9|(140-10) Бодай голови не піднесли всі ті, хто мене оточив, бодай зло їхніх уст їх покрило!
PS|140|10|(140-11) Хай присок на них упаде, нехай кине Він їх до огню, до провалля, щоб не встали вони!...
PS|140|11|(140-12) Злоязична людина щоб міцною вона не була на землі, людина насильства бодай лихо спіймало її, щоб попхнути на погибіль!
PS|140|12|(140-13) Я знаю, що зробить Господь правосуддя убогому, присуд правдивий для бідних,
PS|140|13|(140-14) тільки праведні дякувати будуть іменню Твоєму, невинні сидітимуть перед обличчям Твоїм!
PS|141|1|Псалом Давидів. Господи, кличу до Тебе, поспішися до мене, почуй же мій голос, як кличу до Тебе!
PS|141|2|Нехай стане молитва моя як кадило перед лицем Твоїм, підношення рук моїх як жертва вечірня!
PS|141|3|Поклади, Господи, сторожу на уста мої, стережи двері губ моїх!
PS|141|4|Не дай нахилятися серцю моєму до речі лихої, щоб учинки робити безбожністю, із людьми, що чинять переступ, і щоб не ласувався я їхніми присмаками!
PS|141|5|Як праведний вразить мене, то це милість, а докорить мені, це олива на голову, її не відкине моя голова, бо ще і молитва моя проти їхнього зла.
PS|141|6|Їхні судді по скелі розкидані, та слова мої вчують, бо приємні вони...
PS|141|7|Як дрова рубають й розколюють їх на землі, так розкидані наші кістки над отвором шеолу.
PS|141|8|Бо до Тебе, о Господи, Владико, мої очі, на Тебе надіюсь не зруйновуй мого життя!
PS|141|9|Бережи Ти від пастки мене, що на мене поставили, та від тенет переступників!
PS|141|10|Хай безбожні попадають разом до сітки своєї, а я промину!
PS|142|1|Псалом навчальний, Давида, коли був у печері. Молитва. (142-2) Мій голос до Господа, я кличу, мій голос до Господа, я благаю!
PS|142|2|(142-3) Перед обличчям Його виливаю я мову свою, про недолю свою я розказую перед обличчям Його,
PS|142|3|(142-4) коли омліває мій дух у мені. А Ти знаєш дорогу мою: на дорозі, якою ходжу, пастку для мене сховали!
PS|142|4|(142-5) Праворуч поглянь і побач: немає нікого знайомого, загинув притулок від мене, ніхто не питає за душу мою...
PS|142|5|(142-6) Я кличу до Тебе, о Господи, я кажу: Ти моє пристановище, доля моя у країні живих!
PS|142|6|(142-7) Прислухайся ж Ти до благання мого, бо зробився я зовсім нужденний! Визволь мене від моїх переслідників, бо стали сильніші від мене вони!
PS|142|7|(142-8) Виведи душу мою із в'язниці, щоб славити Ймення Твоє! Праведні оточать мене, як учиниш добро надо мною!
PS|143|1|Псалом Давидів. Господи, вислухай молитву мою, почуй благання моє в Своїй вірності, у правді Своїй обізвися до мене!
PS|143|2|і на суд не вступай із рабом Своїм, бо жоден живий перед обличчям Твоїм справедливим не буде!
PS|143|3|Бо неприятель переслідує душу мою, топче живую мою до землі... Посадив мене в темряву, як мерців цього світу!
PS|143|4|Омліває мій дух у мені, кам'яніє в нутрі моїм серце моє...
PS|143|5|Я згадую дні стародавні, над усіми Твоїми чинами роздумую, говорю про діла Твоїх рук.
PS|143|6|Я руки свої простягаю до Тебе, душа моя прагне Тебе, як води пересохла земля! Села.
PS|143|7|Поспіши мене вислухати, Господи, дух мій кінчається! Не ховай Ти від мене обличчя Свого, і нехай я не буду подібний до тих, хто сходить до гробу!
PS|143|8|Об'яви мені вранці Своє милосердя, бо на Тебе надіюсь, повідом Ти мене про дорогу, якою я маю ходити, бо до Тебе підношу я душу свою!
PS|143|9|Урятуй мене, Господи, від моїх ворогів, бо до Тебе вдаюся!
PS|143|10|Навчи мене волю чинити Твою, бо Ти Бог мій, добрий Дух Твій нехай попровадить мене по рівній землі!
PS|143|11|Ради Ймення Свого, о Господи, оживи мене, Своєю правдою виведи душу мою від недолі!
PS|143|12|А в Своїм милосерді понищ моїх ворогів, і вигуби всіх, хто ненавидить душу мою, бо я раб Твій!
PS|144|1|Давидів. Благословенний Господь, моя скеля, що руки мої Він навчає до бою, пальці мої до війни!
PS|144|2|Він моє милосердя й твердиня моя, фортеця моя та моя охорона мені, Він мій щит, і я до Нього вдаюся, Він мій народ підбиває під мене!
PS|144|3|Господи, що то людина, що знаєш її, що то син людський, що зважаєш на нього?
PS|144|4|Людина стала до пари подібна, її дні як та тінь проминуща!
PS|144|5|Господи, нахили Своє небо, й зійди, доторкнися до гір, і вони задимують!
PS|144|6|Заблищи блискавицею, й їх розпорош, пошли Свої стріли, і їх побентеж!
PS|144|7|Пошли з висоти Свою руку, й мене порятуй, і визволь мене з вод великих, від руки чужинців,
PS|144|8|що їхні уста промовляють неправду, а їхня правиця правиця зрадлива!
PS|144|9|Боже, я пісню нову заспіваю Тобі, на арфі десятиструнній заграю Тобі,
PS|144|10|що Ти перемогу царям подаєш, що рятуєш Давида, Свого раба, від лихого меча!
PS|144|11|Порятуй же мене й збережи Ти мене від руки чужинців, що їхні уста промовляють марноту, а їхня правиця правиця зрадлива,
PS|144|12|щоб були сини наші, немов саджанці, виплекані в їхній молодості, наші дочки немов ті наріжні стовпи, витесані на окрасу палати!
PS|144|13|Повні наші комори, вони видають найрізніше, котяться тисячами наші вівці та кози, десятками тисяч по наших подвір'ях розплоджуються!
PS|144|14|Ситі наші бики, немає пригод і немає хвороби, і на вулицях наших нема нарікань!
PS|144|15|Блаженний народ, що йому так ведеться, блаженний народ, що Господь йому Бог!
PS|145|1|Хвала Давидова. Я буду Тебе величати, о Боже мій, Царю, і благословлятиму Ймення Твоє повік-віку!
PS|145|2|Я кожного дня Тебе благословлятиму, і хвалитиму Ймення Твоє повік-віку!
PS|145|3|Великий Господь і прославлений вельми, і недослідиме величчя Його!
PS|145|4|Рід родові буде хвалити діла Твої, і будуть могутність Твою виявляти!
PS|145|5|Про пишну славу величчя Твого, про справи чудовні Твої розповім!
PS|145|6|Будуть казати про силу грізних Твоїх чинів, а про велич Твою розповім я про неї.
PS|145|7|Пам'ять про добрість велику Твою сповіщатимуть, і будуть співати про правду Твою!
PS|145|8|Щедрий і милосердний Господь, довготерпеливий й многомилостивий,
PS|145|9|Господь добрий до всіх, а Його милосердя на всі Його творива!
PS|145|10|Тебе, Господи, славити будуть усі Твої творива, а святі Твої Тебе благословлятимуть,
PS|145|11|про славу Царства Твого звіщатимуть, про могутність Твою говоритимуть,
PS|145|12|щоб людським синам об'явити про могутність Його та про славу величчя Царства Його!
PS|145|13|Царство Твоє царство всіх віків, а влада Твоя по всі роди!
PS|145|14|Господь підпирає всіх падаючих, усіх зігнутих Він випростовує!
PS|145|15|Очі всіх уповають на Тебе, і Ти їм поживу даєш своєчасно,
PS|145|16|Ти руку Свою відкриваєш, і все, що живе, Ти зичливо годуєш!
PS|145|17|Господь справедливий на кожній дорозі Своїй, і милостивий у всіх Своїх учинках,
PS|145|18|Господь близький всім, хто взиває до Нього, хто правдою кличе Його!
PS|145|19|Волю тих, хто боїться Його, Він сповняє, і благання їх чує та їм помагає,
PS|145|20|Господь береже тих усіх, хто любить Його, а безбожних усіх Він понищить!
PS|145|21|Славу Господню уста мої будуть звіщати, і благословлятиме кожне тіло святе Його Ймення на віки віків!
PS|146|1|Алілуя! Хвали, душе моя, Господа,
PS|146|2|хвалитиму Господа, поки живу, співатиму Богу моєму, аж поки існую!
PS|146|3|Не надійтесь на князів, на людського сина, бо в ньому спасіння нема:
PS|146|4|вийде дух його і він до своєї землі повертається, того дня його задуми гинуть!
PS|146|5|Блаженний, кому його поміч Бог Яковів, що надія його на Господа, Бога його,
PS|146|6|що небо та землю вчинив, море й усе, що є в них, що правди пильнує навіки,
PS|146|7|правосуддя вчиняє покривдженим, що хліба голодним дає! Господь в'язнів розв'язує,
PS|146|8|Господь очі сліпим відкриває, Господь випростовує зігнутих, Господь милує праведних!
PS|146|9|Господь обороняє приходьків, сироту та вдовицю підтримує, а дорогу безбожних викривлює!
PS|146|10|Хай царює навіки Господь, Бог твій, Сіоне, із роду у рід! Алілуя!
PS|147|1|Хваліть Господа, добрий бо Він, виспівуйте нашому Богу, приємний бо Він, Йому подобає хвала!
PS|147|2|Господь Єрусалима будує, збирає вигнанців ізраїлевих.
PS|147|3|Він зламаносердих лікує, і їхні рани болючі обв'язує,
PS|147|4|вираховує Він число зорям, і кожній із них дає ймення.
PS|147|5|Великий Господь наш, та дужий на силі, Його мудрости міри нема!
PS|147|6|Господь підіймає слухняних, безбожних понижує аж до землі.
PS|147|7|Дайте відповідь Господу нашому вдячною піснею, заграйте для нашого Бога на гуслах:
PS|147|8|Він хмарами небо вкриває, приготовлює дощ для землі, оброщує гори травою,
PS|147|9|худобі дає її корм, воронятам чого вони кличуть!
PS|147|10|Не в силі коня уподоба Його, і не в членах людини Його закохання,
PS|147|11|Господь любить тих, хто боїться Його, хто надію складає на милість Його!
PS|147|12|Хвали Господа, Єрусалиме, прославляй Свого Бога, Сіоне,
PS|147|13|бо зміцняє Він засуви брам твоїх, синів твоїх благословляє в тобі,
PS|147|14|чинить мир у границі твоїй, годує тебе пшеницею щирою,
PS|147|15|посилає на землю наказа Свого, дуже швидко летить Його Слово!
PS|147|16|Дає сніг, немов вовну, розпорошує паморозь, буцім то порох,
PS|147|17|Він кидає лід Свій, немов ті кришки, і перед морозом Його хто устоїть?
PS|147|18|Та Він пошле Своє слово, та й розтопить його, Своїм вітром повіє, вода потече!
PS|147|19|Своє слово звіщає Він Якову, постанови Свої та Свої правосуддя ізраїлю:
PS|147|20|для жодного люду Він так не зробив, той не знають вони правосуддя Його! Алілуя!
PS|148|1|Алілуя! Хваліте Господа з небес, хваліте Його в висоті!
PS|148|2|Хваліте Його, всі Його Анголи, хваліте Його, усі війська Його:
PS|148|3|Хваліте Його, сонце й місяцю, хваліте Його, усі зорі ясні!
PS|148|4|Хваліте Його, небеса із небес, та води, що над небесами!
PS|148|5|Нехай Господа хвалять вони, бо Він наказав, і створились вони,
PS|148|6|Він їх поставив на вічні віки, дав наказа, і не переступлять його!
PS|148|7|Хваліть Господа також з землі: риби великі й безодні усі,
PS|148|8|огонь та град, сніг та туман, вітер бурхливий, що виконує слово Його,
PS|148|9|гори та пагірки всі, плідне дерево та всі кедрини,
PS|148|10|звірина й вся худоба, все плазуюче та птаство крилате,
PS|148|11|земні царі й всі народи, князі та всі судді землі,
PS|148|12|юнаки та дівиці, старі разом із дітьми,
PS|148|13|нехай усі хвалять Господнє ім'я, бо Його тільки Ймення звеличилось, величність Його на землі й небесах!
PS|148|14|Він рога народу Своєму підніс! Слава всім богобійним Його, дітям ізраїлевим, народові, що до Нього близький! Алілуя!
PS|149|1|Алілуя! Заспівайте для Господа пісню нову, Йому слава на зборах святих!
PS|149|2|Хай ізраїль радіє Творцем своїм, хай Царем своїм тішаться діти Сіону!
PS|149|3|Нехай славлять ім'я Його танцем, нехай вигравають для Нього на бубні та гуслах,
PS|149|4|бо знаходить Господь уподобу в народі Своїм, прикрашає покірних спасінням!
PS|149|5|Хай радіють у славі святі, хай співають на ложах своїх,
PS|149|6|прославлення Бога на їхніх устах, а меч обосічний ув їхніх руках,
PS|149|7|щоб чинити між племенами помсту, між народами кари,
PS|149|8|щоб їхніх царів пов'язати кайданами, а їхніх вельмож ланцюгами,
PS|149|9|щоб між ними чинити суд написаний! Він величність для всіх богобійних! Алілуя!
PS|150|1|Алілуя! Хваліть Бога в святині Його, хваліте Його на могутнім Його небозводі!
PS|150|2|Хваліте Його за чини могутні Його, хваліте Його за могутню величність Його!
PS|150|3|Хваліте Його звуком трубним, хваліте Його на арфі та гуслах!
PS|150|4|Хваліте Його на бубні та танцем, хваліте Його на струнах та флейті!
PS|150|5|Хваліте Його на цимбалах дзвінких, хваліте Його на цимбалах гучних!
PS|150|6|Все, що дихає, хай Господа хвалить! Алілуя!
