EXOD|1|1|以色列 的眾兒子各帶著家眷，和 雅各 一同來到 埃及 ，他們的名字如下：
EXOD|1|2|呂便 、 西緬 、 利未 、 猶大 、
EXOD|1|3|以薩迦 、 西布倫 、 便雅憫 、
EXOD|1|4|但 、 拿弗他利 、 迦得 、 亞設 。
EXOD|1|5|凡從 雅各 生的，共有七十人。那時， 約瑟 已經在 埃及 。
EXOD|1|6|約瑟 和他所有的兄弟，以及那一代的人都死了。
EXOD|1|7|然而， 以色列 人生養眾多，繁衍昌盛，極其強盛，遍滿了那地。
EXOD|1|8|有一位不認識 約瑟 的新王興起，統治 埃及 。
EXOD|1|9|他對自己的百姓說：「看哪， 以色列 人的百姓比我們還多，又比我們強盛。
EXOD|1|10|來吧，讓我們機巧地待他們，恐怕他們增多起來，將來若有戰爭，他們就聯合我們的仇敵來攻擊我們，然後離開這地去了。」
EXOD|1|11|於是 埃及 人派監工管轄他們，用勞役苦待他們。他們為法老建造儲貨城，就是 比東 和 蘭塞 。
EXOD|1|12|可是越苦待他們，他們就越發增多，更加繁衍， 埃及 人就因 以色列 人愁煩。
EXOD|1|13|埃及 人嚴厲地強迫 以色列 人做工，
EXOD|1|14|使他們因苦工而生活痛苦；無論是和泥，是做磚，是做田間各樣的工，一切的工 埃及 人都嚴厲地對待他們。
EXOD|1|15|埃及 王又對 希伯來 的接生婆，一個名叫 施弗拉 ，另一個名叫 普阿 的說：
EXOD|1|16|「你們為 希伯來 婦人接生，臨盆的時候要注意 ，若是男的，就把他殺了，若是女的，就讓她活。」
EXOD|1|17|但是接生婆敬畏上帝，不照 埃及 王的吩咐去做，卻讓男孩活著。
EXOD|1|18|埃及 王召了接生婆來，對她們說：「你們為甚麼做這事，讓男孩活著呢？」
EXOD|1|19|接生婆對法老說：「因為 希伯來 婦人與 埃及 婦人不同； 希伯來 婦人健壯，接生婆還沒有到，她們已經生產了。」
EXOD|1|20|上帝恩待接生婆； 以色列 人增多起來，極其強盛。
EXOD|1|21|接生婆因為敬畏上帝，上帝就叫她們成立家室。
EXOD|1|22|法老吩咐他的眾百姓說：「把所生的 每一個男孩都丟到 尼羅河 裏去，讓所有的女孩存活。」
EXOD|2|1|有一個 利未 家的人娶了一個 利未 女子為妻。
EXOD|2|2|那女人懷孕，生了一個兒子，見他俊美，就把他藏了三個月，
EXOD|2|3|後來不能再藏，就取了一個蒲草箱，抹上柏油和樹脂，將孩子放在裏面，把箱子擱在 尼羅河 邊的蘆葦中。
EXOD|2|4|孩子的姊姊遠遠站著，要知道他究竟會怎樣。
EXOD|2|5|法老的女兒來到 尼羅河 邊洗澡，她的女僕們在河邊行走。她看見在蘆葦中的箱子，就派一個使女把它拿來。
EXOD|2|6|她打開箱子，看見那孩子。看哪，男孩在哭，她就可憐他，說：「這是 希伯來 人的一個孩子。」
EXOD|2|7|孩子的姊姊對法老的女兒說：「我去叫一個 希伯來 婦人來作奶媽，替你乳養這孩子，好嗎？」
EXOD|2|8|法老的女兒對她說：「去吧！」那女孩就去叫了孩子的母親來。
EXOD|2|9|法老的女兒對她說：「你把這孩子抱去，替我乳養這孩子，我必給你工錢。」那婦人就把孩子接過來，乳養他。
EXOD|2|10|孩子長大了，婦人把他帶到法老的女兒那裏，就作了她的兒子。她給孩子起名叫 摩西 ，說：「因我把他從水裏拉出來。」
EXOD|2|11|過了一段日子， 摩西 長大了，他出去到他同胞那裏，看見他們的勞役。他看見一個 埃及 人打他的同胞，一個 希伯來 人。
EXOD|2|12|他左右觀看，見沒有人，就把 埃及 人打死了，藏在沙土裏。
EXOD|2|13|第二天他出去，看哪，有兩個 希伯來 人在打架，他就對那兇惡的人說：「你為甚麼打你同族的人呢？」
EXOD|2|14|那人說：「誰立你作我們的領袖和審判官呢？難道你要殺我，像殺那 埃及 人一樣嗎？」 摩西 就懼怕，說：「這事一定是讓人知道了。」
EXOD|2|15|法老聽見這事，就設法要殺 摩西 。於是 摩西 逃走，躲避法老，到了 米甸 地，坐在井旁。
EXOD|2|16|米甸 的祭司有七個女兒；她們來打水，打滿了槽，要給父親的羊群喝水。
EXOD|2|17|有一些牧羊人來，把她們趕走， 摩西 卻起來幫助她們，取水給她們的羊群喝。
EXOD|2|18|她們回到父親 流珥 那裏；他說：「今日你們為何這麼快就回來了呢？」
EXOD|2|19|她們說：「有一個 埃及 人來救我們脫離牧羊人的手，他甚至打水給我們的羊群喝。」
EXOD|2|20|他對女兒們說：「那人在哪裏？你們為甚麼撇下他呢？去請他來吃飯吧！」
EXOD|2|21|摩西 願意和那人同住， 那人就把女兒 西坡拉 給 摩西 為妻。
EXOD|2|22|西坡拉 生了一個兒子， 摩西 給他起名叫 革舜 ，因他說：「我在外地作了寄居者。」
EXOD|2|23|過了許多年， 埃及 王死了。 以色列 人因做苦工，就嘆息哀求；他們因苦工所發出的哀聲達於上帝。
EXOD|2|24|上帝聽見他們的哀聲，就記念他與 亞伯拉罕 、 以撒 、 雅各 所立的約。
EXOD|2|25|上帝看顧 以色列 人，上帝是知道的 。
EXOD|3|1|摩西 牧放他岳父 米甸 祭司 葉特羅 的羊群，他領羊群往曠野的那一邊去，到了上帝的山，就是 何烈山 。
EXOD|3|2|耶和華的使者在荊棘的火焰中向他顯現。 摩西 觀看，看哪，荊棘在火中焚燒，卻沒有燒燬。
EXOD|3|3|摩西 說：「我要轉過去看這大異象，這荊棘為何沒有燒燬呢？」
EXOD|3|4|耶和華見 摩西 轉過去看，上帝就從荊棘裏呼叫他說：「 摩西 ！ 摩西 ！」他說：「我在這裏。」
EXOD|3|5|上帝說：「不要靠近這裏。把你腳上的鞋脫下來，因為你所站的地方是聖地」。
EXOD|3|6|他又說：「我是你父親的上帝，是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。」 摩西 蒙上臉，因為怕看上帝。
EXOD|3|7|耶和華說：「我確實看見了我百姓在 埃及 所受的困苦，我也聽見了他們因受監工苦待所發的哀聲；我確實知道他們的痛苦。
EXOD|3|8|我下來是要救他們脫離 埃及 人的手，領他們從那地上來，到美好與寬闊之地，到流奶與蜜之地，就是 迦南 人、 赫 人、 亞摩利 人、 比利洗 人、 希未 人、 耶布斯 人之地。
EXOD|3|9|現在，看哪， 以色列 人的哀聲達到我這裏，我也看見 埃及 人怎樣欺壓他們。
EXOD|3|10|現在，你去，我要差派你到法老那裏，把我的百姓 以色列 人從 埃及 領出來。」
EXOD|3|11|摩西 對上帝說：「我是甚麼人，竟能去見法老，把 以色列 人從 埃及 領出來呢？」
EXOD|3|12|上帝說：「我必與你同在。這就是我差派你去，給你的憑據：你把百姓從 埃及 領出來之後，你們必在這山上事奉上帝。」
EXOD|3|13|摩西 對上帝說：「看哪，我到 以色列 人那裏，對他們說：『你們祖宗的上帝差派我到你們這裏來。』他們若對我說：『他叫甚麼名字？』我要對他們說甚麼呢？」
EXOD|3|14|上帝對 摩西 說：「我是自有永有的」；又說：「你要對 以色列 人這樣說：『那自有永有的差派我到你們這裏來。』」
EXOD|3|15|上帝又對 摩西 說：「你要對 以色列 人這樣說：『耶和華－你們祖宗的上帝，就是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝差派我到你們這裏來。』這是我的名，直到永遠；這也是我的稱號 ，直到萬代。
EXOD|3|16|你去召集 以色列 的長老，對他們說：『耶和華－你們祖宗的上帝，就是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝向我顯現，說：我實在眷顧了你們，眷顧你們在 埃及 的遭遇。
EXOD|3|17|我也曾說：要把你們從 埃及 的困苦中領出來，往 迦南 人、 赫 人、 亞摩利 人、 比利洗 人、 希未 人、 耶布斯 人的地去，就是到流奶與蜜之地。』
EXOD|3|18|他們必聽你的話。你和 以色列 的長老要到 埃及 王那裏，對他說：『耶和華－ 希伯來 人的上帝向我們顯現，現在求你讓我們往曠野去，走三天的路程，為要向耶和華我們的上帝獻祭。』
EXOD|3|19|我知道若不用大能的手， 埃及 王不會放你們走。
EXOD|3|20|因此，我必伸出我的手，在 埃及 施行我一切的神蹟，擊打這地，然後，他才放你們走。
EXOD|3|21|我必使 埃及 人看得起你們，你們離開的時候就不至於空手而去。
EXOD|3|22|每一個婦女必向她的鄰舍，以及寄居在她家裏的女人，索取金器、銀器和衣裳，給你們的兒女穿戴。這樣你們就掠奪了 埃及 人。」
EXOD|4|1|摩西 回答說：「看哪！他們不會信我，也不會聽我的話，因為他們必說：『耶和華並沒有向你顯現。』」
EXOD|4|2|耶和華對 摩西 說：「你手裏的是甚麼？」他說：「是杖。」
EXOD|4|3|耶和華說：「把它丟在地上！」他一丟在地上，杖就變成一條蛇； 摩西 逃走避開牠。
EXOD|4|4|耶和華對 摩西 說：「伸出手來，拿住牠的尾巴─ 摩西 就伸出手，抓住牠，牠就在 摩西 的手掌中變為杖─
EXOD|4|5|為了要使他們信耶和華他們祖宗的上帝，就是 亞伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝，曾向你顯現了。」
EXOD|4|6|耶和華又對他說：「把手放進懷裏。」他就把手放進懷裏。當他把手抽出來，看哪，手竟然長了痲瘋 ，像雪一樣白。
EXOD|4|7|耶和華說：「把手放回懷裏─他就把手放回懷裏。當他把手從懷裏再抽出來，看哪，手復原了，與全身的肉一樣─
EXOD|4|8|倘若他們不信你，也不聽第一個神蹟的聲音，他們會信第二個神蹟的聲音。
EXOD|4|9|倘若他們不信這兩個神蹟，不聽你的話，你就從 尼羅河 裏取些水，倒在乾的地上。你從 尼羅河 裏所取的水必在乾地上變成血。」
EXOD|4|10|摩西 對耶和華說：「主啊，求求你，我並不是一個能言善道的人，以前這樣，就是你對僕人說話以後也是這樣，因為我是拙口笨舌的。」
EXOD|4|11|耶和華對他說：「誰造人的口呢？誰使人口啞、耳聾、目明、眼瞎呢？豈不是我－耶和華嗎？
EXOD|4|12|現在，去吧，我必賜你口才，指教你應當說的。」
EXOD|4|13|摩西 說：「主啊，求求你，你要藉著誰的手，就差派誰去吧！」
EXOD|4|14|耶和華的怒氣向 摩西 發作，說：「你不是有一個哥哥 利未 人 亞倫 嗎？我知道他是個能言善道的人。看哪，他正出來迎接你。他一見到你，心裏就歡喜。
EXOD|4|15|你要跟他說話，把話放在他的口裏，我要賜你口才，也要賜他口才，又要教你們做當做的事。
EXOD|4|16|他要替你向百姓說話；他要當你的口，你要當他的上帝。
EXOD|4|17|你手裏要拿這杖，用它來行神蹟。」
EXOD|4|18|於是， 摩西 回到他岳父 葉特羅 那裏，對他說：「請你讓我回 埃及 我同胞那裏，看他們還在不在。」 葉特羅 對 摩西 說：「平平安安地去吧！」
EXOD|4|19|耶和華在 米甸 對 摩西 說：「你要回 埃及 去，因為那些尋索你命的人都死了。」
EXOD|4|20|摩西 就帶著妻子和兩個兒子，讓他們騎上驢，回 埃及 地去。 摩西 手裏拿著上帝的杖。
EXOD|4|21|耶和華對 摩西 說：「你回到 埃及 去的時候，要留意將我交在你手中的一切奇事行在法老面前。但我要任憑他的心剛硬，他必不放百姓走。
EXOD|4|22|你要對法老說：『耶和華如此說： 以色列 是我的兒子，我的長子。
EXOD|4|23|我對你說過：放我的兒子走，好事奉我。你還是不肯放他走。看哪，我要殺你頭生的兒子。』」
EXOD|4|24|在路上住宿的地方，耶和華遇見 摩西 ，想要殺他。
EXOD|4|25|西坡拉 就拿一塊火石，割下她兒子的包皮，碰觸 摩西 的腳，說：「你真是我血的新郎了。」
EXOD|4|26|這樣，耶和華才放了他。那時， 西坡拉 說：「你因割禮就是血的新郎 了」。
EXOD|4|27|耶和華對 亞倫 說：「你往曠野去迎接 摩西 。」他就去，在上帝的山遇見 摩西 ，就親他。
EXOD|4|28|摩西 將耶和華差派他所說的話和吩咐他所行的神蹟都告訴了 亞倫 。
EXOD|4|29|摩西 和 亞倫 就去召集 以色列 的眾長老。
EXOD|4|30|亞倫 將耶和華對 摩西 所說的一切話述說了一遍，又在百姓眼前行了那些神蹟，
EXOD|4|31|百姓就信了。他們聽見耶和華眷顧 以色列 人，鑒察他們的困苦，就低頭敬拜。
EXOD|5|1|後來， 摩西 和 亞倫 去對法老說：「耶和華－ 以色列 的上帝這樣說：『放我的百姓走，好讓他們在曠野向我守節。』」
EXOD|5|2|法老說：「耶和華是誰，要我聽他的話，讓 以色列 人去？我不認識耶和華，也不放 以色列 人走！」
EXOD|5|3|他們說：「 希伯來 人的上帝已向我們顯現了。求你讓我們往曠野去，走三天的路程，向耶和華我們的上帝獻祭，免得他用瘟疫、刀劍攻擊我們。」
EXOD|5|4|埃及 王對他們說：「 摩西 、 亞倫 ！你們為甚麼叫百姓不做工呢？去，服你們的勞役吧！」
EXOD|5|5|他又說：「看哪，這地的 以色列 人如今這麼多，你們竟然叫他們歇下勞役！」
EXOD|5|6|當天，法老吩咐監工和工頭說：
EXOD|5|7|「你們不可照以前一樣提供草給百姓做磚，要叫他們自己去撿草。
EXOD|5|8|他們平時做磚的數目，你們仍舊向他們要，一點不可減少，因為他們是懶惰的，所以才呼求說：『讓我們去向我們的上帝獻祭。』
EXOD|5|9|你們要把更重的工作加在這些人身上，使他們在其中勞碌，不去理會謊言。」
EXOD|5|10|監工和工頭出來對百姓說：「法老這樣說：『我不給你們草，
EXOD|5|11|你們自己在哪裏能找到草，就往哪裏去找吧！但你們的工作一點也不可減少。』」
EXOD|5|12|於是，百姓分散在 埃及 全地，撿碎秸當草用。
EXOD|5|13|監工催逼他們，說：「你們每天要做完一天的工，與先前有草一樣。」
EXOD|5|14|法老的監工擊打他們所派的 以色列 工頭，說：「為甚麼昨天和今天你們沒有按照以前做磚的數目，完成你們的工作呢？」
EXOD|5|15|以色列 人的工頭來哀求法老說：「為甚麼這樣待你的僕人呢？
EXOD|5|16|監工不把草給僕人，並且對我們說：『做磚吧！』看哪，你僕人挨了打，其實是你百姓的錯。」
EXOD|5|17|法老卻說：「懶惰，你們真是懶惰！所以你們說：『讓我們去向耶和華獻祭吧。』
EXOD|5|18|現在，去做工吧！草是不會給你們，磚卻要如數交納。」
EXOD|5|19|以色列 人的工頭聽見「你們每天做磚的工作一點也不可減少」，就知道惹上禍了。
EXOD|5|20|他們離開法老出來，正遇見 摩西 和 亞倫 站在那裏等候他們，
EXOD|5|21|就向他們說：「願耶和華鑒察你們，施行判斷，因為你們使我們在法老和他臣僕面前有了臭名，把刀遞在他們手中來殺我們。」
EXOD|5|22|摩西 回到耶和華那裏，說：「主啊，你為甚麼苦待這百姓呢？為甚麼差派我呢？
EXOD|5|23|自從我到法老那裏，奉你的名說話，他就苦待這百姓，你卻一點也沒有拯救你的百姓。」
EXOD|6|1|耶和華對 摩西 說：「現在你必看見我向法老所行的事，使他因我大能的手放 以色列 人走，因我大能的手把他們趕出他的地。」
EXOD|6|2|上帝吩咐 摩西 ，對他說：「我是耶和華。
EXOD|6|3|我從前向 亞伯拉罕 、 以撒 、 雅各 顯現為全能的上帝；至於我的名耶和華，我未曾讓他們知道。
EXOD|6|4|我要與他們堅立我的約，要把 迦南 地，他們寄居的地賜給他們。
EXOD|6|5|我聽見 以色列 人被 埃及 人奴役的哀聲，我就記念我的約。
EXOD|6|6|所以你要對 以色列 人說：『我是耶和華；我要除去 埃及 人加給你們的勞役，救你們脫離他們的奴役。我要用伸出來的膀臂，藉嚴厲的懲罰救贖你們。
EXOD|6|7|我要以你們為我的百姓，我也要作你們的上帝。我除去 埃及 人加給你們的勞役，你們就知道我是耶和華你們的上帝。
EXOD|6|8|我起誓應許給 亞伯拉罕 、 以撒 、 雅各 的地，我要領你們進去，將那地賜給你們為業。我是耶和華。』」
EXOD|6|9|摩西 把這話告訴 以色列 人，但是他們因心裏愁煩，又因苦工，就不肯聽 摩西 的話。
EXOD|6|10|耶和華吩咐 摩西 說：
EXOD|6|11|「你去對 埃及 王法老說，讓 以色列 人離開他的地。」
EXOD|6|12|摩西 在耶和華面前說：「看哪， 以色列 人尚且不聽我，法老怎麼會聽我這不會講話的人呢？」
EXOD|6|13|耶和華吩咐 摩西 和 亞倫 ，命令他們到 以色列 人和 埃及 王法老那裏，把 以色列 人從 埃及 地領出來。
EXOD|6|14|以色列 人族長的名字如下： 以色列 長子 呂便 的兒子是 哈諾 、 法路 、 希斯倫 、 迦米 ；這是 呂便 的家族。
EXOD|6|15|西緬 的兒子是 耶母利 、 雅憫 、 阿轄 、 雅斤 、 瑣轄 ，和 迦南 女子生的兒子 掃羅 ；這是 西緬 的家族。
EXOD|6|16|以下是 利未 的兒子按著家譜的名字： 革順 、 哥轄 、 米拉利 。 利未 一生的歲數是一百三十七歲。
EXOD|6|17|革順 的兒子按著家族是 立尼 、 示每 。
EXOD|6|18|哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 、 烏薛 。 哥轄 一生的歲數是一百三十三歲。
EXOD|6|19|米拉利 的兒子是 抹利 和 母示 ；這是 利未 按著家譜的家族。
EXOD|6|20|暗蘭 娶了他父親的妹妹 約基別 為妻，她為他生了 亞倫 和 摩西 。 暗蘭 一生的歲數是一百三十七歲。
EXOD|6|21|以斯哈 的兒子是 可拉 、 尼斐 、 細基利 。
EXOD|6|22|烏薛 的兒子是 米沙利 、 以利撒反 、 西提利 。
EXOD|6|23|亞倫 娶了 亞米拿達 的女兒， 拿順 的妹妹， 以利沙巴 為妻，她為他生了 拿答 、 亞比戶 、 以利亞撒 、 以他瑪 。
EXOD|6|24|可拉 的兒子是 亞惜 、 以利加拿 、 亞比亞撒 ；這是 可拉 的家族。
EXOD|6|25|亞倫 的兒子 以利亞撒 娶了 普鐵 的一個女兒為妻，她為他生了 非尼哈 。這是 利未 人按著家族的族長。
EXOD|6|26|這就是曾聽見耶和華說「把 以色列 人按著隊伍從 埃及 地領出來」的 亞倫 和 摩西 ，
EXOD|6|27|對 埃及 王法老說要將 以色列 人從 埃及 領出來的，也是這 摩西 和 亞倫 。
EXOD|6|28|當耶和華在 埃及 地對 摩西 說話的時候，
EXOD|6|29|耶和華對 摩西 說：「我是耶和華；我對你所說的一切話，你都要告訴 埃及 王法老。」
EXOD|6|30|摩西 在耶和華面前說：「看哪，我是不會講話的人，法老怎麼會聽我呢？」
EXOD|7|1|耶和華對 摩西 說：「我使你在法老面前像上帝一樣，你的哥哥 亞倫 是你的代言人 。
EXOD|7|2|凡我所吩咐你的，你都要說。你的哥哥 亞倫 要對法老說，讓 以色列 人離開他的地。
EXOD|7|3|我要使法老的心固執，我也要在 埃及 地多行神蹟奇事。
EXOD|7|4|法老必不聽從你們，因此我要伸手嚴厲地懲罰 埃及 ，把我的軍隊，就是我的百姓 以色列 人從 埃及 地領出來。
EXOD|7|5|我伸手攻擊 埃及 ，把 以色列 人從他們中間領出來的時候， 埃及 人就知道我是耶和華。」
EXOD|7|6|摩西 和 亞倫 就去做；他們照耶和華吩咐的去做了。
EXOD|7|7|摩西 和 亞倫 與法老說話的時候， 摩西 八十歲， 亞倫 八十三歲。
EXOD|7|8|耶和華對 摩西 和 亞倫 說：
EXOD|7|9|「法老若吩咐你們說：『你們行一件奇事吧！』你就對 亞倫 說：『把杖丟在法老面前！杖會變成蛇。』」
EXOD|7|10|摩西 和 亞倫 到法老那裏去，照耶和華所吩咐的去做。 亞倫 把杖丟在法老和他臣僕面前，杖就變成蛇。
EXOD|7|11|法老也召了智慧人和行邪術的人來，這些 埃及 術士也用邪術照樣做。
EXOD|7|12|他們各人丟下自己的杖，杖就變成蛇；但 亞倫 的杖吞了他們的杖。
EXOD|7|13|法老心裏剛硬，不聽 摩西 和 亞倫 ，正如耶和華所說的。
EXOD|7|14|耶和華對 摩西 說：「法老心硬，不肯放百姓走。
EXOD|7|15|明天早晨你要到法老那裏去，看哪，他出來往水邊去，你要到 尼羅河 邊去迎見他，手裏拿著那根變過蛇的杖。
EXOD|7|16|你要對他說：『耶和華－ 希伯來 人的上帝差派我到你這裏，說：放我的百姓走，到曠野事奉我。看哪，到如今你還是不聽。
EXOD|7|17|耶和華如此說：看哪，我要用我手裏的杖擊打 尼羅河 中的水，水就變成血；這樣，你就知道我是耶和華。
EXOD|7|18|河裏的魚必死，河也要發臭， 埃及 人就厭惡喝這河裏的水。』」
EXOD|7|19|耶和華對 摩西 說：「你要對 亞倫 說：『拿你的杖，伸出你的手在 埃及 所有的水上，在他們的江、河、池塘，所有水聚集的地方上，叫水變成血。在 埃及 全地，無論在木器中，石器中，都必有血。』」
EXOD|7|20|摩西 和 亞倫 就照耶和華所吩咐的去做。 亞倫 在法老和他臣僕眼前舉杖擊打 尼羅河 裏的水，河裏的水都變成血了。
EXOD|7|21|河裏的魚死了，河也臭了， 埃及 人就不能喝這河裏的水； 埃及 遍地都有了血。
EXOD|7|22|但是， 埃及 的術士也用邪術照樣做了；法老心裏剛硬，不聽 摩西 和 亞倫 ，正如耶和華所說的。
EXOD|7|23|法老轉身回宮去，並不把這事放在心上。
EXOD|7|24|所有的 埃及 人都沿著 尼羅河 邊挖掘，要找水喝，因為他們不能喝河裏的水。
EXOD|7|25|耶和華擊打 尼羅河 後，過了七天。
EXOD|8|1|耶和華對 摩西 說：「你要到法老那裏，對他說：『耶和華如此說：放我的百姓走，好事奉我。
EXOD|8|2|你若不肯放他們走，看哪，我必以青蛙之災擊打你的疆土。
EXOD|8|3|尼羅河 要滋生青蛙；這青蛙要上來進你的宮殿和你的臥房，上你的床榻，進你臣僕的房屋，上你百姓的身上，進你的爐灶和你的揉麵盆。
EXOD|8|4|這些青蛙要跳上你、你百姓和你眾臣僕的身上。』」
EXOD|8|5|耶和華對 摩西 說：「你要對 亞倫 說：『伸出你手裏的杖在江、河、池塘上，把青蛙帶上 埃及 地來。』」
EXOD|8|6|亞倫 伸手在 埃及 的眾水上，青蛙就上來，遮滿了 埃及 地。
EXOD|8|7|術士也用他們的邪術照樣去做，把青蛙帶上 埃及 地。
EXOD|8|8|法老召 摩西 和 亞倫 來，說：「請你們祈求耶和華使這些青蛙離開我和我的百姓，我就讓這百姓去向耶和華獻祭。」
EXOD|8|9|摩西 對法老說：「悉聽尊便，告訴我何時為你、你臣僕和你的百姓祈求，使青蛙被剪除，離開你和你的宮殿，只留在 尼羅河 裏。」
EXOD|8|10|他說：「明天。」 摩西 說：「就照你的話吧，為要叫你知道沒有像耶和華我們上帝的，
EXOD|8|11|青蛙必會離開你、你宮殿、你臣僕和你的百姓，只留在 尼羅河 裏。」
EXOD|8|12|於是 摩西 和 亞倫 離開法老出去。 摩西 為了青蛙的事呼求耶和華，因為他帶來青蛙攪擾法老。
EXOD|8|13|耶和華就照 摩西 的請求去做；在屋裏、院中、田間的青蛙都死了。
EXOD|8|14|眾人把青蛙聚攏成堆，地就發出臭氣。
EXOD|8|15|但法老見災禍舒緩了，就硬著心，不聽從他們，正如耶和華所說的。
EXOD|8|16|耶和華對 摩西 說：「你要對 亞倫 說：『伸出你的杖擊打地上的塵土，使塵土在 埃及 全地變成蚊子 。』」
EXOD|8|17|他們就照樣做了。 亞倫 伸出他手裏的杖，擊打地上的塵土，人和牲畜身上就有了蚊子； 埃及 全地的塵土都變成蚊子了。
EXOD|8|18|術士也用邪術要照樣產生蚊子，卻做不成。於是人和牲畜的身上都有了蚊子。
EXOD|8|19|術士對法老說：「這是上帝的手指。」法老心裏剛硬，不聽 摩西 和 亞倫 ，正如耶和華所說的。
EXOD|8|20|耶和華對 摩西 說：「你要清早起來，站在法老面前。看哪，法老來到水邊，你就對他說：『耶和華如此說：放我的百姓走，好事奉我。
EXOD|8|21|你若不放我的百姓走，看哪，我要派成群的蒼蠅到你、你臣僕和你百姓身上，進你的宮殿； 埃及 人的房屋和他們所住的地都要滿了成群的蒼蠅。
EXOD|8|22|那一日，我必把我百姓所住的 歌珊 地分別出來，使那裏沒有成群的蒼蠅，好叫你知道我─耶和華是在全地之中。
EXOD|8|23|我要施行救贖，區隔我的百姓和你的百姓。明天必有這神蹟。』」
EXOD|8|24|耶和華就這樣做了。大群的蒼蠅進入法老的宮殿和他臣僕的房屋；在 埃及 全地，地就因這成群的蒼蠅毀壞了。
EXOD|8|25|法老召了 摩西 和 亞倫 來，說：「去，在此地向你們的上帝獻祭。」
EXOD|8|26|摩西 說：「這樣做是不妥的，因為我們要獻給耶和華－我們上帝的祭物是 埃及 人所厭惡的；看哪，我們在 埃及 人眼前獻他們所厭惡的，他們豈不拿石頭打死我們嗎？
EXOD|8|27|我們要遵照耶和華－我們上帝所吩咐我們的，往曠野去，走三天路程，向他獻祭。」
EXOD|8|28|法老說：「我可以放你們走，在曠野向耶和華－你們的上帝獻祭，只是不可走得太遠。你們要為我祈禱。」
EXOD|8|29|摩西 說：「看哪，我要從你這裏出去祈求耶和華，使成群的蒼蠅明天離開法老、法老的臣僕和法老的百姓；法老卻不可再欺騙，不讓百姓去向耶和華獻祭。」
EXOD|8|30|於是 摩西 離開法老，去祈求耶和華。
EXOD|8|31|耶和華就照 摩西 的請求去做，使成群的蒼蠅離開法老、他的臣僕和他的百姓，一隻也沒有留下。
EXOD|8|32|但這一次法老又硬著心，不放百姓走。
EXOD|9|1|耶和華對 摩西 說：「你要到法老那裏，對他說：『耶和華－ 希伯來 人的上帝如此說：放我的百姓走，好事奉我。
EXOD|9|2|你若不肯放他們走，仍要強留他們，
EXOD|9|3|看哪，耶和華的手必以嚴重的瘟疫加在你田間的牲畜上，就是在馬、驢、駱駝、牛群和羊群的身上。
EXOD|9|4|耶和華卻要分別 以色列 的牲畜和 埃及 的牲畜，凡屬 以色列 人的，一隻都不死。』」
EXOD|9|5|耶和華就設定時間，說：「明天耶和華必在此地行這事。」
EXOD|9|6|第二天，耶和華行了這事。 埃及 的牲畜全都死了，只是 以色列 人的牲畜，一隻都沒有死。
EXOD|9|7|法老派人去，看哪， 以色列 人的牲畜連一隻都沒有死。可是法老硬著心，不放百姓走。
EXOD|9|8|耶和華對 摩西 和 亞倫 說：「你們從爐裏滿滿捧出爐灰， 摩西 要在法老眼前把它撒在空中。
EXOD|9|9|這灰要在 埃及 全地變成塵土，使 埃及 全地的人和牲畜身上起泡生瘡。」
EXOD|9|10|摩西 和 亞倫 取了爐灰，站在法老面前。 摩西 把它撒在空中，人和牲畜的身上就起泡生瘡了。
EXOD|9|11|因為這瘡，術士在 摩西 面前站立不住，術士和所有 埃及 人的身上都生了瘡。
EXOD|9|12|但耶和華任憑法老的心剛硬，不聽 摩西 和 亞倫 ，正如耶和華對 摩西 所說的。
EXOD|9|13|耶和華對 摩西 說：「你要清早起來，站在法老面前，對他說：『耶和華－ 希伯來 人的上帝如此說：放我的百姓走，好事奉我。
EXOD|9|14|因為這一次我要使一切的災禍臨到你自己，你臣僕和你百姓的身上，為要叫你知道在全地沒有像我的。
EXOD|9|15|現在，我若伸手用瘟疫攻擊你和你的百姓，你就會從地上除滅了。
EXOD|9|16|然而，我讓你存活，是為了要使你看見我的大能，並要使我的名傳遍全地。
EXOD|9|17|可是你仍然向我的百姓自高自大，不放他們走。
EXOD|9|18|看哪，明天大約這時候，我必使大量的冰雹降下，這是從 埃及 立國直到如今沒有出現過的。
EXOD|9|19|現在，你要派人把你的牲畜和你田間一切所有的帶去躲避；任何在田間，無論是人是牲畜沒有回到屋內的，冰雹必降在他們身上，他們就必死。』」
EXOD|9|20|法老的臣僕中，懼怕耶和華這話的，就讓他的奴僕和牲畜逃進屋裏。
EXOD|9|21|但那不把耶和華這話放在心上的，就把他的奴僕和牲畜留在田裏。
EXOD|9|22|耶和華對 摩西 說：「你向天伸出你的手，使冰雹降在 埃及 全地，降在 埃及 地的人和牲畜身上，以及田間各樣菜蔬上。」
EXOD|9|23|摩西 向天伸杖，耶和華就打雷下雹，有火降到地上；耶和華下雹在 埃及 地上。
EXOD|9|24|那時，有雹，也有火在雹中閃爍，極其嚴重；自從 埃及 立國以來，全地沒有像這樣的。
EXOD|9|25|在 埃及 全地，冰雹擊打田間所有的人和牲畜，擊打一切的菜蔬，也打壞了田間一切的樹木。
EXOD|9|26|惟獨 以色列 人所住的 歌珊 地沒有冰雹。
EXOD|9|27|法老差派人去召 摩西 和 亞倫 來，對他們說：「這一次我犯罪了。耶和華是公義的；我和我的百姓是邪惡的。
EXOD|9|28|請你們祈求耶和華，因上帝的雷轟和冰雹已經夠了。我要放你們走，你們不用再留下來了。」
EXOD|9|29|摩西 對他說：「我一出城就向耶和華舉起雙手；雷必止住，也不再有冰雹，叫你知道地是屬於耶和華的。
EXOD|9|30|至於你和你的臣僕，我知道你們仍然不敬畏耶和華上帝。」
EXOD|9|31|那時，亞麻和大麥被摧毀了，因為大麥已經吐穗，亞麻也開了花。
EXOD|9|32|只是小麥和粗麥沒有被摧毀，因為它們還沒有長成。
EXOD|9|33|摩西 離開法老出了城，向耶和華舉起雙手，雷和雹就止住，雨也不再下在地上了。
EXOD|9|34|法老見雨、雹、雷止住，又再犯罪；他和他的臣僕都硬著心。
EXOD|9|35|法老的心剛硬，不放 以色列 人走，正如耶和華藉著 摩西 所說的。
EXOD|10|1|耶和華對 摩西 說：「你要到法老那裏，因我使他硬著心，也使他臣僕硬著心，為要在他們中間 顯出我的這些神蹟來，
EXOD|10|2|並要叫你將我嚴厲對付 埃及 的事，和在他們中間所行的神蹟，傳於兒子和孫子的耳中，好叫你們知道我是耶和華。」
EXOD|10|3|摩西 和 亞倫 就到法老那裏，對他說：「耶和華－ 希伯來 人的上帝這樣說：『你在我面前不肯謙卑要到幾時呢？放我的百姓走，好事奉我。
EXOD|10|4|你若不肯放我的百姓走，看哪，明天我要使蝗蟲進入你的境內，
EXOD|10|5|遮滿地面 ，甚至地也看不見了。牠們要吃那冰雹後所剩，就是留給你們的；並且要吃那生長在田間的一切樹木。
EXOD|10|6|你的宮殿和你眾臣僕的房屋，以及一切 埃及 人的房屋，都要被蝗蟲佔滿；你祖宗和你祖宗的祖宗在世以來，直到今日都沒有見過。』」 摩西 就轉身離開法老出去。
EXOD|10|7|法老的臣僕對法老說：「這傢伙成為我們的羅網要到幾時呢？讓這些人去事奉耶和華－他們的上帝吧！ 埃及 快要滅亡了，你還不知道嗎？」
EXOD|10|8|於是 摩西 和 亞倫 被召回來見法老。法老對他們說：「去，事奉耶和華－你們的上帝吧！但要去的是哪些人呢？」
EXOD|10|9|摩西 說：「我們要帶著年老的和年少的同去，要帶著我們的兒子和女兒，以及我們的羊群牛群一起去，因為我們要向耶和華守節。」
EXOD|10|10|法老對他們說：「願耶和華與你們同在吧！我若讓你們帶著你們的孩子同去，看，災禍就在你們面前 ！
EXOD|10|11|不可都去！你們壯年人去事奉耶和華吧，因為這是你們所求的。」於是法老把他們從自己面前趕出去。
EXOD|10|12|耶和華對 摩西 說：「你向 埃及 地伸出你的手，使蝗蟲上到 埃及 地，吃地上冰雹後所剩一切的植物。」
EXOD|10|13|摩西 就向 埃及 地伸杖；整整一晝一夜，耶和華使東風颳在 埃及 地上，到了早晨，東風把蝗蟲颳了來。
EXOD|10|14|蝗蟲上到 埃及 全地，落在 埃及 全境，非常厲害；蝗蟲這麼多，是空前絕後的。
EXOD|10|15|蝗蟲遮滿地面，地上一片黑暗。牠們吃盡了地上一切的植物和冰雹過後所剩樹上的果子。 埃及 全地，無論是樹木，是田間的植物，連一點綠的也沒有留下。
EXOD|10|16|於是法老急忙召了 摩西 和 亞倫 來，說：「我得罪了耶和華－你們的上帝，又得罪了你們。
EXOD|10|17|現在求你，就這一次，饒恕我的罪，祈求耶和華－你們的上帝救我脫離這次的死亡。」
EXOD|10|18|摩西 就離開法老，去祈求耶和華。
EXOD|10|19|耶和華轉變風向，使強勁的西風吹來，把蝗蟲颳起，吹入 紅海 ；在 埃及 全境連一隻也沒有留下。
EXOD|10|20|但耶和華任憑法老的心剛硬，不放 以色列 人走。
EXOD|10|21|耶和華對 摩西 說：「你向天伸出你的手，使黑暗籠罩 埃及 地；這黑暗甚至可以摸得到。」
EXOD|10|22|摩西 向天伸出他的手，濃密的黑暗就籠罩了 埃及 全地三天之久。
EXOD|10|23|三天內，人人彼此看不見，誰也不敢起身離開原地；但所有 以色列 人住的地方卻有光。
EXOD|10|24|法老就召 摩西 來，說：「去，事奉耶和華吧！只是你們的羊群牛群要留下來。你們的孩子可以和你們同去。」
EXOD|10|25|摩西 說：「你必須把祭物和燔祭牲交在我們手中，讓我們可以向耶和華我們的上帝獻祭。
EXOD|10|26|我們的牲畜也要與我們同去，連一蹄也不留下，因為我們要從牲畜中挑選來事奉耶和華－我們的上帝。未到那裏之前，我們還不知道要用甚麼來事奉耶和華。」
EXOD|10|27|但耶和華任憑法老的心剛硬，法老不肯放他們走。
EXOD|10|28|法老對 摩西 說：「離開我去吧！你要小心，不要再見我的面，因為再見我面的那日，你就必死！」
EXOD|10|29|摩西 說：「就照你說的，我也不要再見你的面了！」
EXOD|11|1|耶和華對 摩西 說：「我要再降一個災禍給法老和 埃及 ，然後他必讓你們離開這裏。他放你們走的時候，一定會趕你們全都離開這裏。
EXOD|11|2|你要傳於百姓耳中，叫他們男的女的各向鄰舍索取金器銀器。」
EXOD|11|3|耶和華使 埃及 人看得起他的百姓 ，並且 摩西 在 埃及 地，在法老臣僕和百姓眼中看為偉大。
EXOD|11|4|摩西 說：「耶和華如此說：『約到半夜，我必出去走遍 埃及 。
EXOD|11|5|凡在 埃及 地，從坐寶座的法老到推磨 的婢女所生的長子，以及一切頭生的牲畜，都必死。
EXOD|11|6|埃及 全地必有大大的哀號，這將是空前絕後的。
EXOD|11|7|至於 以色列 人中，無論是人是牲畜，連狗也不敢向他們吠叫，使你們知道耶和華區別 埃及 和 以色列 。』
EXOD|11|8|你所有的這些臣僕都要下到我這裏，向我下拜說：『請你和跟從你的百姓都離開吧！』然後我才離開。」於是， 摩西 氣憤憤地離開法老出去了。
EXOD|11|9|耶和華對 摩西 說：「法老必不聽你們，為了要使我在 埃及 地多行奇事。」
EXOD|11|10|摩西 和 亞倫 在法老面前行了這一切奇事，但耶和華任憑法老的心剛硬，不讓 以色列 人離開他的地。
EXOD|12|1|耶和華在 埃及 地對 摩西 和 亞倫 說：
EXOD|12|2|「你們要以本月為正月，為一年之首。
EXOD|12|3|你們要吩咐 以色列 全會眾說：本月初十，各人要按著家庭 取羔羊，一家一隻羔羊。
EXOD|12|4|若一家的人太少，吃不了一隻羔羊，就要按照人數和隔壁的鄰舍共取一隻；你們要按每人的食量來估算羔羊。
EXOD|12|5|你們要從綿羊或山羊中取一隻無殘疾、一歲的公羔羊，
EXOD|12|6|要把牠留到本月十四日；那日黃昏的時候， 以色列 全會眾要把羔羊宰了。
EXOD|12|7|他們要取一些血，塗在他們吃羔羊的房屋兩邊的門框上和門楣上。
EXOD|12|8|當晚要吃羔羊的肉；要用火烤了，與無酵餅和苦菜一起吃。
EXOD|12|9|不可吃生的，或用水煮的，要把羔羊連頭帶腿和內臟用火烤了吃。
EXOD|12|10|一點也不可留到早晨；若有留到早晨的，要用火燒了。
EXOD|12|11|你們要這樣吃羔羊：腰間束帶，腳上穿鞋，手中拿杖，快快地吃。這是耶和華的逾越。
EXOD|12|12|因為那夜我要走遍 埃及 地，把 埃及 地一切頭生的，無論是人是牲畜，都擊殺了；我要對 埃及 所有的神明施行審判。我是耶和華。
EXOD|12|13|這血要在你們所住的房屋上作記號；我一見這血，就逾越你們。我擊打 埃及 地的時候，災殃必不臨到你們身上施行毀滅。」
EXOD|12|14|「你們要記念這日，世世代代守這日為耶和華的節日，作為你們永遠的定例。
EXOD|12|15|你們要吃無酵餅七日。第一日要把酵從你們各家中除去，因為從第一日到第七日，任何吃有酵之物的，必從 以色列 中剪除。
EXOD|12|16|第一日當有聖會，第七日也當有聖會。在這兩日，任何工作都不可做，只能預備各人的食物，這是惟一可做的工作。
EXOD|12|17|你們要守除酵節，因為我在這一日把你們的軍隊從 埃及 地領出來。所以，你們要世世代代守這日，立為永遠的定例。
EXOD|12|18|從正月十四日晚上，直到二十一日晚上，你們要吃無酵餅。
EXOD|12|19|在你們各家中，七日之內不可有酵，因為凡吃有酵之物的，無論是寄居的，是本地的，必從 以色列 的會中剪除。
EXOD|12|20|任何有酵的物，你們都不可吃；在你們一切的住處要吃無酵餅。」
EXOD|12|21|於是， 摩西 召了 以色列 的眾長老來，對他們說：「你們要為家人取羔羊，把逾越的羔羊宰了。
EXOD|12|22|要拿一把牛膝草，蘸盆裏的血，把盆裏的血塗在門楣上和兩邊的門框上。直到早晨你們誰也不可出自己家裏的門。
EXOD|12|23|因為耶和華要走遍 埃及 ，施行擊殺，他看見血在門楣上和兩邊的門框上，耶和華就必逾越那門，不讓滅命者進你們的家，施行擊殺。
EXOD|12|24|你們要守這命令，作為你們和你們子孫永遠的定例。
EXOD|12|25|日後，你們到了耶和華所應許賜給你們的那地，就要守這禮儀。
EXOD|12|26|你們的兒女對你們說：『這禮儀是甚麼意思呢？』
EXOD|12|27|你們就說：『這是獻給耶和華逾越節的祭物。當耶和華擊殺 埃及 人的時候，他逾越了 以色列 人在 埃及 的房屋，救了我們各家。』」於是百姓低頭敬拜。
EXOD|12|28|以色列 人就去做；他們照耶和華吩咐 摩西 和 亞倫 的去做了。
EXOD|12|29|到了半夜，耶和華把 埃及 地所有頭生的，就是從坐寶座的法老，到關在牢裏的人的長子，以及一切頭生的牲畜，盡都殺了。
EXOD|12|30|法老和他眾臣僕，以及所有的 埃及 人，都在夜間起來了。在 埃及 有大大的哀號，因為沒有一家不死人的。
EXOD|12|31|夜間，法老召了 摩西 和 亞倫 來，說：「起來！你們和 以色列 人，都離開我的百姓出去，照你們所說的，去事奉耶和華吧！
EXOD|12|32|照你們所說的，連羊群牛群也帶走，也為我祝福吧！」
EXOD|12|33|埃及 人催促百姓趕快離開那地，因為 埃及 人說：「我們都快死了。」
EXOD|12|34|百姓就拿著沒有發酵的生麵，把揉麵盆包在衣服中，扛在肩上。
EXOD|12|35|以色列 人照 摩西 的話去做，向 埃及 人索取金器、銀器和衣裳。
EXOD|12|36|耶和華使 埃及 人看得起他的百姓， 埃及 人就給了他們所要的。他們就掠奪了 埃及 人。
EXOD|12|37|以色列 人從 蘭塞 起程，往 疏割 去。除了小孩，步行的男人約有六十萬。
EXOD|12|38|又有許多不同族群的人，以及眾多的羊群牛群，和他們一同上去。
EXOD|12|39|他們用 埃及 帶出來的生麵烤成無酵餅。這生麵是沒有發酵的；因為他們被催促離開 埃及 ，不能耽延，就沒有為自己預備食物。
EXOD|12|40|以色列 人住在 埃及 共四百三十年。
EXOD|12|41|正滿四百三十年的那一天，耶和華的全軍從 埃及 地出來了。
EXOD|12|42|這是向耶和華守的夜，他領他們出 埃及 地；這是 以色列 眾人世世代代要向耶和華守的夜。
EXOD|12|43|耶和華對 摩西 和 亞倫 說：「逾越節的條例是這樣：外邦人不可吃這羔羊。
EXOD|12|44|但是你們用銀子買來，又受過割禮的奴僕可以吃。
EXOD|12|45|寄居的和雇工都不可吃。
EXOD|12|46|應當在一個屋子裏吃，不可把肉帶到屋外，骨頭一根也不可折斷。
EXOD|12|47|以色列 全會眾都要守這禮儀。
EXOD|12|48|若有外人寄居在你那裏，要向耶和華守逾越節，他所有的男子務要先受割禮，然後才可以當他是本地人，容許他守這禮儀。但未受割禮的都不可吃這羔羊。
EXOD|12|49|本地人和寄居在你們中間的外人當守同一個條例。」
EXOD|12|50|以色列 眾人就去做，他們照耶和華吩咐 摩西 和 亞倫 的去做了。
EXOD|12|51|正當那日，耶和華將 以色列 人按著他們的隊伍從 埃及 地領了出來。
EXOD|13|1|耶和華吩咐 摩西 說：
EXOD|13|2|「頭生的要分別為聖歸我； 以色列 中凡頭生的，無論是人是牲畜，都是我的。」
EXOD|13|3|摩西 對百姓說：「你們要記念從 埃及 為奴之家出來的這日，因為耶和華用大能的手將你們從這地領出來。有酵之物都不可吃。
EXOD|13|4|亞筆月的這一日你們走出來了。
EXOD|13|5|將來耶和華領你進 迦南 人、 赫 人、 亞摩利 人、 希未 人、 耶布斯 人之地，就是他向你祖宗起誓應許給你的那流奶與蜜之地，那時你要在這一個月守這禮儀。
EXOD|13|6|你要吃無酵餅七日，在第七日要向耶和華守節。
EXOD|13|7|這七日之內，要吃無酵餅；在你的全境內不可見有酵之物，也不可見酵母。
EXOD|13|8|當那日，你要告訴你的兒子說：『這樣做是因為耶和華在我出 埃及 的時候為我所做的事。』
EXOD|13|9|這要在你手上作記號，在你額上 作紀念，使耶和華的教導常在你口中，因為耶和華用大能的手將你從 埃及 領出來。
EXOD|13|10|所以你每年要按著日期守這條例。」
EXOD|13|11|「當耶和華照他向你和你祖宗所起的誓將你領進 迦南 人之地，把那地賜給你的時候，
EXOD|13|12|你要將一切頭生的獻給耶和華；你牲畜中頭生的，公的都歸耶和華。
EXOD|13|13|然而，凡頭生的驢，你要用羔羊贖回；若不贖牠，就要打斷牠的頸項。你兒子中的長子都要贖出來。
EXOD|13|14|日後，你的兒子問你說：『這是甚麼意思？』你就說：『耶和華用大能的手將我們從 埃及 為奴之家領出來。
EXOD|13|15|那時法老固執，不肯放我們走，耶和華就把 埃及 地所有頭生的，無論是人是牲畜，都殺了。因此，我把一切頭生的公的牲畜獻給耶和華為祭，卻將所有頭生的兒子贖出來。
EXOD|13|16|這要在你手上作記號，在你額上作經匣 ，因為耶和華用大能的手將我們從 埃及 領出來。』」
EXOD|13|17|法老放百姓走的時候， 非利士 人之地的路雖近，上帝卻不領他們從那裏走，因為上帝說：「恐怕百姓遇見戰爭就後悔，轉回 埃及 去。」
EXOD|13|18|上帝領百姓繞道而行，走曠野的路到 紅海 。 以色列 人出 埃及 地，都帶著兵器上去 。
EXOD|13|19|摩西 把 約瑟 的骸骨一起帶走；因為 約瑟 曾叫 以色列 人鄭重地起誓，對他們說：「上帝必定眷顧你們，你們要把我的骸骨從這裏一起帶上去。」
EXOD|13|20|他們從 疏割 起程，在曠野邊上的 以倘 安營。
EXOD|13|21|耶和華走在他們前面，日間用雲柱引領他們的路，夜間用火柱照亮他們，使他們日夜都可以行走。
EXOD|13|22|日間的雲柱，夜間的火柱，總不離開百姓的面前。
EXOD|14|1|耶和華吩咐 摩西 說：
EXOD|14|2|「你吩咐 以色列 人轉回，要在 比‧哈希錄 前面， 密奪 和海的中間， 巴力‧洗分 的前面安營。你們要在對面，靠近海邊安營。
EXOD|14|3|以色列 人這樣做，法老必說：『他們在此地迷了路，曠野把他們困住了。』
EXOD|14|4|我要任憑法老的心剛硬，他要追趕他們。我必在法老和他全軍身上得榮耀， 埃及 人就知道我是耶和華。」於是 以色列 人照樣做了。
EXOD|14|5|有人報告 埃及 王說：「百姓逃跑了！」法老和他的臣僕對百姓改變了心意，說：「我們放 以色列 人走，不再服事我們，我們怎麼會做這種事呢？」
EXOD|14|6|法老就預備戰車，帶領他的軍兵同去，
EXOD|14|7|他帶了六百輛特選的戰車和 埃及 所有的戰車，每輛都有軍官。
EXOD|14|8|耶和華任憑 埃及 王法老的心剛硬，他就追趕 以色列 人； 以色列 人卻抬起頭 來出去了。
EXOD|14|9|埃及 人追趕他們，法老一切的馬匹、戰車、戰車長，與軍兵就在海邊上，靠近 比‧哈希錄 ，在 巴力‧洗分 的前面，在他們安營的地方追上了。
EXOD|14|10|法老逼近的時候， 以色列 人舉目，看哪， 埃及 人追來了，就非常懼怕， 以色列 人向耶和華哀求。
EXOD|14|11|他們對 摩西 說：「難道 埃及 沒有墳地，你要把我們帶來死在曠野嗎？你為甚麼這樣待我們，將我們從 埃及 領出來呢？
EXOD|14|12|我們在 埃及 豈沒有對你說過，不要攪擾我們，讓我們服事 埃及 人嗎？因為服事 埃及 人總比死在曠野好。」
EXOD|14|13|摩西 對百姓說：「不要怕，要站穩，看耶和華今天向你們所要施行的拯救，因為你們今天所看見的 埃及 人必永遠不再看見了。
EXOD|14|14|耶和華必為你們爭戰，你們要安靜！」
EXOD|14|15|耶和華對 摩西 說：「你為甚麼向我哀求呢？你吩咐 以色列 人往前走。
EXOD|14|16|你舉手向海伸杖，把水分開。 以色列 人要下到海中，走在乾地上。
EXOD|14|17|看哪，我要任憑 埃及 人的心剛硬，他們就跟著下去。我要在法老和他的全軍、戰車、戰車長身上得榮耀。
EXOD|14|18|我在法老和他的戰車、戰車長身上得榮耀的時候， 埃及 人就知道我是耶和華。」
EXOD|14|19|在 以色列 營前行走的上帝的使者移動，走到他們後面；雲也從他們的前面移動，站在他們後面。
EXOD|14|20|它來到 埃及 營和 以色列 營的中間：一邊有雲和黑暗，另一邊它照亮夜晚，整夜彼此不得接近。
EXOD|14|21|摩西 向海伸手，耶和華就用強勁的東風，使海水在一夜間退去，海就成了乾地；水分開了。
EXOD|14|22|以色列 人下到海中，走在乾地上，水在他們左右成了牆壁。
EXOD|14|23|埃及 人追趕他們，法老一切的馬匹、戰車和戰車長都跟著下到海中。
EXOD|14|24|破曉時分，耶和華從雲柱、火柱中瞭望 埃及 的軍兵，使 埃及 的軍兵混亂。
EXOD|14|25|他使他們的車輪脫落 ，難以前行， 埃及 人說：「我們從 以色列 人面前逃跑吧！因耶和華為他們作戰，攻擊 埃及 了。」
EXOD|14|26|耶和華對 摩西 說：「你要向海伸手，使水回流到 埃及 人，他們的戰車和戰車長身上。」
EXOD|14|27|摩西 就向海伸手，到了天亮的時候，海恢復原狀。 埃及 人逃避水的時候，耶和華把他們推入海中。
EXOD|14|28|海水回流，淹沒了戰車和戰車長，以及那些跟著 以色列 人下到海中的法老全軍，連一個也沒有剩下。
EXOD|14|29|以色列 人卻在海中走乾地，水在他們的左右成了牆壁。
EXOD|14|30|那一日，耶和華拯救 以色列 脫離 埃及 人的手。 以色列 人看見 埃及 人死在海邊。
EXOD|14|31|以色列 人看見耶和華向 埃及 人所施展的大能，百姓就敬畏耶和華，並且信服耶和華和他的僕人 摩西 。
EXOD|15|1|那時， 摩西 和 以色列 人向耶和華唱這歌，說： 「我要向耶和華歌唱，因他大大得勝， 將馬和騎馬的投在海中。
EXOD|15|2|耶和華是我的力量，是我的詩歌， 他也成了我的拯救。 這是我的上帝，我要讚美他； 我父親的上帝，我要尊崇他。
EXOD|15|3|耶和華是戰士； 耶和華是他的名。
EXOD|15|4|「法老的戰車、軍兵，他已拋在海中； 法老精選的軍官都沉於 紅海 。
EXOD|15|5|深水淹沒他們； 他們好像石頭墜到深處。
EXOD|15|6|耶和華啊，你的右手施展能力，大顯榮耀； 耶和華啊，你的右手摔碎仇敵。
EXOD|15|7|你大發威嚴，摧毀了你的敵人； 你發出烈怒，吞滅他們如同碎秸。
EXOD|15|8|因你鼻中的氣，水就聚成堆， 大水豎立如壘， 海的中心深水凝結。
EXOD|15|9|仇敵說：『我要追趕，我要追上， 我要分擄物，在他們身上滿足我的心願， 我要拔刀，親手毀滅他們。』
EXOD|15|10|你用風一吹，海水就淹沒他們； 他們像鉛沉在大水之中。
EXOD|15|11|「耶和華啊，眾神明中，誰能像你？ 誰能像你，至聖至榮， 可頌可畏，施行奇事！
EXOD|15|12|你伸出右手， 地就吞滅他們。
EXOD|15|13|「你以慈愛引領你所救贖的百姓； 你以能力引導他們到你的聖所。
EXOD|15|14|萬民聽見就戰抖； 疼痛抓住 非利士 的居民。
EXOD|15|15|那時， 以東 的族長驚惶， 摩押 的英雄被戰兢抓住， 迦南 所有的居民都融化。
EXOD|15|16|驚駭恐懼臨到他們； 耶和華啊，因你膀臂的大能， 他們如石頭寂靜不動， 等候你百姓過去， 等候你所贖的百姓過去。
EXOD|15|17|你要將他們領進去，栽在你產業的山上， 耶和華啊，就是你為自己所造的住處， 主啊，就是你手所建立的聖所。
EXOD|15|18|耶和華必作王，直到永永遠遠！」
EXOD|15|19|法老的馬匹、戰車和戰車長下到海中，耶和華使海水回流到他們身上； 以色列 人卻走在海中的乾地上。
EXOD|15|20|那時， 米利暗 女先知， 亞倫 的姊姊，手裏拿著鈴鼓；眾婦女也跟她出去打鼓跳舞。
EXOD|15|21|米利暗 回應他們： 「你們要歌頌耶和華，因他大大得勝， 將馬和騎馬的投在海中。」
EXOD|15|22|摩西 領 以色列 人從 紅海 起程，到了 書珥 的曠野，在曠野走了三天，找不到水。
EXOD|15|23|到了 瑪拉 ，他們不能喝 瑪拉 的水，因為水是苦的；所以那地名叫 瑪拉 。
EXOD|15|24|百姓就向 摩西 發怨言，說：「我們喝甚麼呢？」
EXOD|15|25|摩西 呼求耶和華，耶和華指示他一棵樹 。他把樹丟在水裏，水就變甜了。 耶和華在那裏為他們定了律例、典章，在那裏考驗他們。
EXOD|15|26|他說：「你若留心聽從耶和華－你上帝的話，行我眼中看為正的事，側耳聽我的誡令，遵守我一切的律例，我就不將所加於 埃及 人的疾病加在你身上，因為我是醫治你的耶和華。」
EXOD|15|27|他們到了 以琳 ，在那裏有十二股水泉，七十棵棕樹；他們就在那裏的水邊安營。
EXOD|16|1|以色列 全會眾從 以琳 起程，在出 埃及 之後第二個月十五日到了 以琳 和 西奈 中間， 汛 的曠野。
EXOD|16|2|以色列 全會眾在曠野向 摩西 和 亞倫 發怨言。
EXOD|16|3|以色列 人對他們說：「我們寧願在 埃及 地死在耶和華手中！那時我們坐在肉鍋旁，吃餅得飽。你們卻將我們領出來，到這曠野，要叫這全會眾都餓死啊！」
EXOD|16|4|耶和華對 摩西 說：「看哪，我要從天降食物給你們。百姓可以出去，每天收集當天的分量。這樣，我就可以考驗他們是否遵行我的指示。
EXOD|16|5|到第六天，他們預備食物，所收集的分量要比每天所收的多一倍。」
EXOD|16|6|摩西 和 亞倫 對 以色列 眾人說：「到了晚上，你們就知道是耶和華將你們從 埃及 地領出來的。
EXOD|16|7|早晨，你們要看見耶和華的榮耀，因為耶和華聽見你們向他所發的怨言了。我們算甚麼，你們竟然向我們發怨言呢？」
EXOD|16|8|摩西 又說：「耶和華晚上必給你們肉吃，早晨必給你們食物得飽，因為耶和華已經聽見你們向他所發的怨言。我們算甚麼呢？你們的怨言不是向我們發的，而是向耶和華發的。」
EXOD|16|9|摩西 對 亞倫 說：「你對 以色列 全會眾說：『你們來到耶和華面前，因為他已經聽見你們的怨言了。』」
EXOD|16|10|亞倫 正對 以色列 全會眾說話的時候，他們轉向曠野，看哪，耶和華的榮光在雲中顯現。
EXOD|16|11|耶和華吩咐 摩西 說：
EXOD|16|12|「我已經聽見 以色列 人的怨言了。你要對他們說：『到黃昏的時候 ，你們要吃肉，早晨也必有食物得飽。你們就知道我是耶和華－你們的上帝。』」
EXOD|16|13|到了晚上，有鵪鶉上來，遮滿營地；早晨，營地周圍有一層露水。
EXOD|16|14|那一層露水蒸發之後，看哪，曠野的表面出現了小圓物，好像地上的薄霜一樣。
EXOD|16|15|以色列 人看見了，不知道是甚麼，就彼此說：「這是甚麼？ 」 摩西 對他們說：「這是耶和華給你們吃的食物。
EXOD|16|16|耶和華所吩咐的是這樣：『你們每個人要按自己的食量收集，各人要為帳棚裏的人收集，按照人口數每個人一俄梅珥。』」
EXOD|16|17|以色列 人就照樣去做；有的收多，有的收少。
EXOD|16|18|用俄梅珥量一量，多收的沒有餘，少收的也沒有缺；各人都按著自己的食量收集。
EXOD|16|19|摩西 對他們說：「任何人都不可以把所收的留到早晨。」
EXOD|16|20|然而他們不聽從 摩西 ，當中有人把食物留到早晨，食物就生蟲發臭了。 摩西 就向他們發怒。
EXOD|16|21|他們每日早晨按著各人的食量收集；太陽一發熱，食物就融化了。
EXOD|16|22|到第六天，他們收集了雙倍的食物，每個人二俄梅珥。會眾的官長來告訴 摩西 ，
EXOD|16|23|摩西 對他們說：「耶和華吩咐：『明天是安息日，是向耶和華守的聖安息日。你們要烤的就烤，要煮的就煮，所剩下的都留到早晨。』」
EXOD|16|24|他們就照 摩西 的吩咐把剩下的留到早晨，這些食物既不發臭，裏頭也沒有生蟲。
EXOD|16|25|摩西 說：「你們今天就吃這些吧！因為今天是向耶和華守的安息日，你們在野外必找不著食物了。
EXOD|16|26|六天可以收集，第七天是安息日，這一天甚麼也沒有了。」
EXOD|16|27|第七天，百姓中有人出去收，甚麼也找不著。
EXOD|16|28|耶和華對 摩西 說：「你們不肯遵守我的誡令和教導，要到幾時呢？
EXOD|16|29|你們看，耶和華既然將安息日賜給你們，所以第六天他就賜給你們兩天的食物，第七天各人都要留在自己的地方，不許任何人從這裏出去。」
EXOD|16|30|於是百姓在第七天安息了。
EXOD|16|31|以色列 家給這食物取名叫嗎哪，它的樣子像芫荽子，顏色是白的，吃起來像和蜜的薄餅。
EXOD|16|32|摩西 說：「耶和華所吩咐的是這樣：『要裝滿一俄梅珥的嗎哪留給你們的後代，使他們可以看見我領你們出 埃及 地的時候，在曠野所給你們吃的食物。』」
EXOD|16|33|摩西 對 亞倫 說：「你拿一個罐子，裝滿一俄梅珥的嗎哪，存在耶和華面前，留給你們的後代。」
EXOD|16|34|耶和華怎麼吩咐 摩西 ， 亞倫 就照樣做，把嗎哪存留作見證 。
EXOD|16|35|以色列 人吃嗎哪共四十年，直到進入有人居住的地方；他們吃嗎哪，直到 迦南 地的邊境。
EXOD|16|36|一俄梅珥是一伊法的十分之一。
EXOD|17|1|以色列 全會眾遵照耶和華的吩咐，從 汛 的曠野一段一段地往前行。他們在 利非訂 安營，但百姓沒有水喝。
EXOD|17|2|百姓就與 摩西 爭鬧，說：「給我們水喝吧！」 摩西 對他們說：「你們為甚麼與我爭鬧呢？你們為甚麼試探耶和華呢？」
EXOD|17|3|百姓在那裏口渴要喝水，就向 摩西 發怨言，說：「你為甚麼把我們從 埃及 領出來，使我們和我們的兒女，以及牲畜都渴死呢？」
EXOD|17|4|摩西 就呼求耶和華說：「我要怎樣對待這百姓呢？他們差一點就要拿石頭打死我了。」
EXOD|17|5|耶和華對 摩西 說：「你帶著 以色列 的幾個長老，走在百姓前面，手裏拿著你先前擊打 尼羅河 的杖，去吧！
EXOD|17|6|看哪，我要在 何烈 的磐石那裏，站在你面前。你要擊打磐石，水就會從磐石流出來，給百姓喝。」 摩西 就在 以色列 的長老眼前這樣做了。
EXOD|17|7|他給那地方起名叫 瑪撒 ，又叫 米利巴 ，因為 以色列 人在那裏爭鬧，並且試探耶和華，說：「耶和華是否在我們中間呢？」
EXOD|17|8|那時， 亞瑪力 來到 利非訂 ，和 以色列 爭戰。
EXOD|17|9|摩西 對 約書亞 說：「你為我們選出人來，出去和 亞瑪力 爭戰。明天我要站在山頂上，手裏拿著上帝的杖。」
EXOD|17|10|於是， 約書亞 照著 摩西 對他所說的話去做，和 亞瑪力 爭戰。 摩西 、 亞倫 和 戶珥 都上了山頂。
EXOD|17|11|摩西 何時舉手， 以色列 就得勝；何時垂手， 亞瑪力 就得勝。
EXOD|17|12|但 摩西 的雙手沉重，他們就搬一塊石頭來放在他下面，他就坐在上面。 亞倫 與 戶珥 扶著他的手，一個在這邊，一個在那邊，他的手就穩住，直到日落。
EXOD|17|13|約書亞 用刀打敗了 亞瑪力 和他的百姓。
EXOD|17|14|耶和華對 摩西 說：「你要把這事記錄在書上作紀念，又念給 約書亞 聽：我要把 亞瑪力 的名字從天下全然塗去。」
EXOD|17|15|摩西 築了一座壇，起名叫「耶和華尼西 」。
EXOD|17|16|他說：「我指著耶和華的寶座發誓 ，耶和華必世世代代和 亞瑪力 爭戰。」
EXOD|18|1|摩西 的岳父， 米甸 祭司 葉特羅 ，聽見上帝為 摩西 和為他百姓 以色列 所行的一切事，就是耶和華將 以色列 從 埃及 領了出來。
EXOD|18|2|摩西 的岳父 葉特羅 帶著 西坡拉 ，就是 摩西 先前送回家的妻子，
EXOD|18|3|又帶著她的兩個兒子：一個名叫 革舜 ，因為 摩西 說：「我在外地作了寄居者」；
EXOD|18|4|另一個名叫 以利以謝 ，因為他說：「我父親的上帝幫助我，救我脫離法老的刀。」
EXOD|18|5|摩西 的岳父 葉特羅 帶著 摩西 的妻子和兩個兒子來到上帝的山，就是 摩西 在曠野安營的地方。
EXOD|18|6|他對 摩西 說：「我是 你岳父 葉特羅 ，帶著你的妻子和兩個兒子來到你這裏。」
EXOD|18|7|摩西 迎接他的岳父，向他下拜，親他，彼此問安，然後進入帳棚。
EXOD|18|8|摩西 將耶和華為 以色列 的緣故向法老和 埃及 人所行的一切事，他們在路上遭遇的一切艱難，以及耶和華怎樣搭救他們，都述說給他的岳父聽。
EXOD|18|9|葉特羅 因耶和華待 以色列 的一切恩惠，就是拯救他們脫離 埃及 人的手，就非常喜樂。
EXOD|18|10|葉特羅 說：「耶和華是應當稱頌的，他救了你們脫離 埃及 人和法老的手，將這百姓從 埃及 人的手裏救出來 。
EXOD|18|11|現在，從 埃及 人狂傲地對待 以色列 人這件事上，我知道耶和華比萬神更大。」
EXOD|18|12|摩西 的岳父 葉特羅 把燔祭和祭物獻給上帝。 亞倫 和 以色列 的眾長老都來了，與 摩西 的岳父在上帝面前吃飯。
EXOD|18|13|第二天， 摩西 坐著審判百姓，百姓從早到晚站在 摩西 的旁邊。
EXOD|18|14|摩西 的岳父看見他為百姓所做的一切事，就說：「你為百姓所做的，這是甚麼事呢？你為甚麼獨自一人坐著，而眾百姓從早到晚都站在你旁邊呢？」
EXOD|18|15|摩西 對岳父說：「這是因為百姓到我這裏來求問上帝。
EXOD|18|16|他們有事的時候，就到我這裏來，我就在雙方之間作判決；我又叫他們知道上帝的律例和法度。」
EXOD|18|17|摩西 的岳父對他說：「你這樣做不好。
EXOD|18|18|你和這些與你在一起的百姓都必疲憊，因為這事太重，你獨自一人做不了。
EXOD|18|19|現在，聽我的話，我給你出個主意，願上帝與你同在。你要代替百姓到上帝面前，將事件帶到上帝那裏，
EXOD|18|20|又要用律例和法度警戒他們，指示他們當行的道，當做的事。
EXOD|18|21|你也要從百姓中選出有才能的人，敬畏上帝、誠實可靠、恨惡不義之財的人，派他們作千夫長、百夫長、五十夫長、十夫長來管理百姓。
EXOD|18|22|他們要隨時審判百姓；重大的事要送到你這裏，小事就由他們自行判決。這樣，你就可以輕省一些，他們可以與你分擔。
EXOD|18|23|你若這樣做，上帝也這樣吩咐你，你就能承受得住，眾百姓也可以和睦地回到自己的地方。」
EXOD|18|24|摩西 聽了他岳父的話，照著他所說的一切去做。
EXOD|18|25|摩西 從 以色列 人中選出有才能的人，立他們為百姓的領袖，作千夫長、百夫長、五十夫長、十夫長。
EXOD|18|26|他們隨時審判百姓：難斷的事就送到 摩西 那裏，各樣小事就由他們自行判決。
EXOD|18|27|於是， 摩西 給他的岳父送行，他就回到本地去了。
EXOD|19|1|以色列 人出 埃及 地以後，第三個月的初一，就在那一天他們來到了 西奈 的曠野。
EXOD|19|2|他們從 利非訂 起程，來到 西奈 的曠野，在那裏的山下安營。
EXOD|19|3|摩西 到上帝那裏，耶和華從山上呼喚他說：「你要這樣告訴 雅各 家，對 以色列 人說：
EXOD|19|4|『我向 埃及 人所行的事，你們都看見了， 我如鷹將你們背在翅膀上，帶你們來歸我。
EXOD|19|5|如今你們若真的聽從我的話，遵守我的約，就要在萬民中作屬我的子民 ，因為全地都是我的。
EXOD|19|6|你們要歸我作祭司的國度，為神聖的國民。』這些話你要告訴 以色列 人。」
EXOD|19|7|摩西 去召了百姓中的長老來，將耶和華吩咐他的話當面告訴他們。
EXOD|19|8|百姓都同聲回答：「凡耶和華所說的，我們一定遵行。」 摩西 就將百姓的話回覆耶和華。
EXOD|19|9|耶和華對 摩西 說：「看哪，我要在密雲中臨到你那裏，叫百姓在我與你說話的時候可以聽見，就可以永遠相信你了。」於是， 摩西 將百姓的話稟告耶和華。
EXOD|19|10|耶和華對 摩西 說：「你往百姓那裏去，使他們今天明天分別為聖，又叫他們洗衣服。
EXOD|19|11|第三天要預備好，因為第三天耶和華要在眾百姓眼前降臨在 西奈山 。
EXOD|19|12|你要在山的周圍給百姓劃定界限，說：『你們當謹慎，不可上山去，也不可摸山的邊界。凡摸這山的，必被處死。
EXOD|19|13|不可用手碰他，要用石頭打死，或射死；無論是人是牲畜，都不可活。』到角聲拉長的時候，他們才可到山腳來。」
EXOD|19|14|摩西 下山到百姓那裏去，使他們分別為聖，他們就洗衣服。
EXOD|19|15|他對百姓說：「第三天要預備好；不可親近女人。」
EXOD|19|16|到了第三天早晨，山上有雷轟、閃電和密雲，並且角聲非常響亮，營中的百姓盡都戰抖。
EXOD|19|17|摩西 率領百姓出營迎見上帝，都站在山下。
EXOD|19|18|西奈山 全山冒煙，因為耶和華在火中降臨山上。山的煙霧上騰，彷彿燒窯，整座山劇烈震動。
EXOD|19|19|角聲越來越響， 摩西 說話，上帝以聲音回答他。
EXOD|19|20|耶和華降臨在 西奈山 頂上，耶和華召 摩西 上山頂， 摩西 就上去了。
EXOD|19|21|耶和華對 摩西 說：「你下去警告百姓，免得他們闖過來看耶和華，就會有許多人死亡。
EXOD|19|22|那些親近耶和華的祭司也要把自己分別為聖，免得耶和華忽然出來擊殺他們。」
EXOD|19|23|摩西 對耶和華說：「百姓不能上 西奈山 ，因為你已經警告我們說：『要在山的周圍劃定界限，使山成聖。』」
EXOD|19|24|耶和華對他說：「下去吧，你要和 亞倫 一起上來；只是祭司和百姓不可闖上來到耶和華這裏，免得耶和華忽然出來擊殺他們。」
EXOD|19|25|於是， 摩西 下到百姓那裏告訴他們。
EXOD|20|1|上帝吩咐這一切的話，說：
EXOD|20|2|「我是耶和華－你的上帝，曾將你從 埃及 地為奴之家領出來。
EXOD|20|3|「除了我以外，你不可有別的神。
EXOD|20|4|「不可為自己雕刻偶像，也不可做甚麼形像，彷彿上天、下地和地底下水中的百物。
EXOD|20|5|不可跪拜那些像，也不可事奉它們，因為我耶和華─你的上帝是忌邪 的上帝。恨我的，我必懲罰他們的罪，自父及子，直到三、四代；
EXOD|20|6|愛我，守我誡命的，我必向他們施慈愛，直到千代。
EXOD|20|7|「不可妄稱耶和華－你上帝的名，因為妄稱耶和華名的，耶和華必不以他為無罪。
EXOD|20|8|「當記念安息日，守為聖日。
EXOD|20|9|六日要勞碌做你一切的工，
EXOD|20|10|但第七日是向耶和華─你的上帝當守的安息日。這一日你和你的兒女、奴僕、婢女、牲畜，以及你城裏寄居的客旅，都不可做任何的工。
EXOD|20|11|因為六日之內，耶和華造天、地、海和其中的萬物，第七日就安息了；所以耶和華賜福與安息日，定為聖日。
EXOD|20|12|「當孝敬父母，使你的日子在耶和華－你上帝所賜你的地上得以長久。
EXOD|20|13|「不可殺人。
EXOD|20|14|「不可姦淫。
EXOD|20|15|「不可偷盜。
EXOD|20|16|「不可做假見證陷害你的鄰舍。
EXOD|20|17|「不可貪戀你鄰舍的房屋；不可貪戀你鄰舍的妻子、奴僕、婢女、牛驢，以及他一切所有的。」
EXOD|20|18|眾百姓見雷轟、閃電、角聲、山上冒煙，百姓看見 就都戰抖，遠遠站著。
EXOD|20|19|他們對 摩西 說：「請你向我們說話，我們必聽；不要讓上帝向我們說話，免得我們死亡。」
EXOD|20|20|摩西 對百姓說：「不要害怕；因為上帝降臨是要考驗你們，要你們敬畏他，不致犯罪。」
EXOD|20|21|於是百姓遠遠站著，但 摩西 卻挨近上帝所在的幽暗中。
EXOD|20|22|耶和華對 摩西 說：「你要向 以色列 人這樣說：『你們親自看見我從天上向你們說話了。
EXOD|20|23|你們不可為我製造偶像，不可為自己造任何金銀的神像。
EXOD|20|24|你要為我築一座土壇，在上面獻牛羊為燔祭和平安祭。凡在我叫你記念我名的地方，我必到那裏賜福給你。
EXOD|20|25|你若為我築一座石壇，不可用鑿過的石頭，因為你在石頭上動了工具，就使壇污穢了。
EXOD|20|26|你不可用臺階上我的壇，免得露出你的下體來。』」
EXOD|21|1|「你在百姓面前所要立的典章是這樣：
EXOD|21|2|「你若買 希伯來 人作奴僕，他服事你六年，第七年他可以自由，白白地離去。
EXOD|21|3|他若單身來就可以單身去；他若是有妻子的，他的妻子可以同他離去。
EXOD|21|4|若他主人給他娶了妻，妻子為他生了兒子或女兒，妻子和兒女要歸主人，他要獨自離去。
EXOD|21|5|倘若奴僕聲明：『我愛我的主人和我的妻子兒女，不願意自由離去。』
EXOD|21|6|他的主人就要帶他到審判官 前，再帶他到門或門框那裏，用錐子穿他的耳朵，他就要永遠服事主人。
EXOD|21|7|「人若賣女兒作婢女，婢女不可像男的奴僕那樣離去。
EXOD|21|8|主人若選定她歸自己，後來看不順眼，就要允許她贖身；主人既然對她失信，就沒有權柄把她賣給外邦人。
EXOD|21|9|主人若選定她給自己的兒子，就當照女兒的規矩對待她。
EXOD|21|10|若另娶一個，她的飲食、衣服和房事不可減少。
EXOD|21|11|若不向她行這三樣，她就可以白白離去，不必付贖金。」
EXOD|21|12|「打人致死的，必被處死。
EXOD|21|13|他若不是出於預謀 ，而是上帝交在他手中，我就設立一個地方，讓他可以逃到那裏。
EXOD|21|14|人若蓄意用詭計殺了他的鄰舍，就是逃到我的壇那裏，也當把他捉去處死。
EXOD|21|15|「打父母的，必被處死。
EXOD|21|16|「誘拐人口的，無論是把人賣了，或是扣留在他手中，必被處死。
EXOD|21|17|「咒罵父母的，必被處死。
EXOD|21|18|「人若彼此爭吵，一個用石頭或拳頭打另一個，被打的人沒有死去，卻要躺臥在床，
EXOD|21|19|若他還能起來扶杖行走，那打他的可免處刑，卻要賠償他不能工作的損失，並要把他完全醫好。
EXOD|21|20|「人若用棍子打奴僕或婢女，當場死在他的手下，他必受報應。
EXOD|21|21|若能撐過一兩天，主人就不必受懲罰，因為那是他的財產。
EXOD|21|22|「人若彼此打鬥，傷害有孕的婦人，以致胎兒掉了出來，隨後卻無別的傷害，那傷害她的人，總要按婦人的丈夫所提出的，照審判官所裁定的賠償。
EXOD|21|23|若有別的傷害，就要以命抵命，
EXOD|21|24|以眼還眼，以牙還牙，以手還手，以腳還腳，
EXOD|21|25|以灼傷還灼傷，以損傷還損傷，以鞭打還鞭打。
EXOD|21|26|「人若打奴僕或婢女的眼睛，毀了一隻，就要因他的眼讓他自由離去。
EXOD|21|27|若打掉了奴僕或婢女的一顆牙，就要因他的牙讓他自由離去。」
EXOD|21|28|「牛若牴死男人或女人，總要用石頭打死那牛，卻不可吃牠的肉；牛的主人可免處刑。
EXOD|21|29|倘若那牛向來是牴人的，牛的主人雖然受過警告，仍不把牠拴好，以致把男人或女人牴死，牛要用石頭打死，主人也要被處死。
EXOD|21|30|若罰他付贖命的賠款，他就要照所罰的數目贖他的命。
EXOD|21|31|牛若牴了男孩或女孩，也要照這條例處理。
EXOD|21|32|牛若牴了奴僕或婢女，就要把三十舍客勒銀子給他的主人，牛要用石頭打死。
EXOD|21|33|「人若敞開井口，或挖井不蓋住它，有牛或驢掉進井裏，
EXOD|21|34|井的主人要拿錢賠償牲畜的主人，死牲畜要歸自己。
EXOD|21|35|「人的牛若牴死鄰舍的牛，他們就要賣了那活牛，平分價錢；也要平分死牛。
EXOD|21|36|若這牛向來是以好牴人出名的，主人竟不把牛拴好，他必要以牛賠牛，死牛卻歸自己。」
EXOD|22|1|「人若偷牛或羊，無論是宰了或賣了，他就要以五牛賠一牛， 四羊賠一羊。
EXOD|22|2|賊挖洞，若被發現而被打死，打的人沒有流血的罪。
EXOD|22|3|若太陽已經出來，打的人就有流血的罪。賊總要賠償，若他一無所有，就要被賣來還他所偷的東西。
EXOD|22|4|若發現他所偷的，無論是牛、驢，或羊，在他手中還活著，他就要加倍賠償。
EXOD|22|5|「人若在田間或葡萄園裏牧放牲畜，任憑牲畜上別人田裏去吃 ，他就要拿自己田間和葡萄園裏上好的賠償。
EXOD|22|6|「若火冒出，延燒到荊棘，以致將堆積的禾捆，直立的莊稼，或田地，都燒盡了，那點火的必要賠償。
EXOD|22|7|「人若將銀錢或物件託鄰舍保管，東西從這人的家中被偷去，若找到了賊，賊要加倍賠償；
EXOD|22|8|若找不到賊，這家的主人就要到審判官 那裏，聲明 自己沒有伸手拿鄰舍的物件。
EXOD|22|9|「關於任何侵害的案件，無論是為牛、驢、羊、衣服，或任何失物，有一人說：『這是我的』，雙方就要將案件帶到審判官面前，審判官定誰有罪，誰就要加倍賠償給他的鄰舍。
EXOD|22|10|「人將驢、牛、羊，或別的牲畜託鄰舍看管，若牲畜死亡，受了傷，或被搶走，無人看見，
EXOD|22|11|雙方要在耶和華前起誓，受託人要表明自己沒有伸手拿鄰舍的東西，原主要接受誓言，受託人不必賠償。
EXOD|22|12|牲畜若從受託人那裏被偷去，他就要賠償原主；
EXOD|22|13|若被野獸撕碎，受託人要帶回來作證據，被撕碎的就不必賠償。
EXOD|22|14|「人若向鄰舍借牲畜 ，所借的或傷或死，原主沒有在場，借的人總要賠償。
EXOD|22|15|若原主在場，借的人不必賠償；若是租用的，只要付租金 。」
EXOD|22|16|「人若引誘沒有訂婚的處女，與她同寢，他就必須交出聘禮，娶她為妻。
EXOD|22|17|若女子的父親堅決不將女子給他，他就要按著處女的聘禮交出錢來。
EXOD|22|18|「行邪術的女人，不可讓她存活。
EXOD|22|19|「凡與獸交合的，必被處死。
EXOD|22|20|「向別神獻祭，不單單獻給耶和華的，那人必要滅絕。
EXOD|22|21|「不可虧待寄居的，也不可欺壓他，因為你們在 埃及 地也作過寄居的。
EXOD|22|22|不可苛待寡婦和孤兒；
EXOD|22|23|若你確實苛待他，他向我苦苦哀求，我一定會聽他的呼求，
EXOD|22|24|並要發烈怒，用刀殺你們，使你們的妻子成為寡婦，兒女成為孤兒。
EXOD|22|25|「我的子民中有困苦人在你那裏，你若借錢給他，不可如放債的向他取利息。
EXOD|22|26|你果真拿了鄰舍的外衣作抵押，也要在日落前還給他；
EXOD|22|27|因為他只有這一件用來作被子，是他蔽體的衣服。他還可以拿甚麼睡覺呢？當他哀求我，我就應允，因為我是有恩惠的。
EXOD|22|28|「不可毀謗上帝；也不可詛咒你百姓的領袖。
EXOD|22|29|「不可遲延獻你的莊稼、酒和油 。 「要將你頭生的兒子歸給我。
EXOD|22|30|你的牛羊也要照樣做：七天當跟著牠母親，第八天你要把牠歸給我。
EXOD|22|31|「你們要分別為聖歸給我。因此，田間被野獸撕裂的肉，你們不可吃，要把它丟給狗。」
EXOD|23|1|「不可散佈謠言；不可與惡人連手作惡意的見證。
EXOD|23|2|不可附和群眾作惡；不可在訴訟中附和群眾歪曲公正，作歪曲的見證；
EXOD|23|3|也不可在訴訟中偏袒貧寒人。
EXOD|23|4|「若遇見你仇敵的牛或驢迷了路，務必牽回來交給他。
EXOD|23|5|若看見恨你的人的驢被壓在重馱之下，不可走開，務要和他一同卸下驢的重馱。
EXOD|23|6|「不可在貧窮人的訴訟中屈枉正直。
EXOD|23|7|當遠離誣告的事。不可殺害無辜和義人，因我必不以惡人為義。
EXOD|23|8|不可接受賄賂，因為賄賂能使明眼人變瞎，又能曲解義人的證詞。
EXOD|23|9|「不可欺壓寄居的，因為你們在 埃及 地作過寄居的，知道寄居者的心情。」
EXOD|23|10|「六年你要耕種田地，收集地的出產。
EXOD|23|11|只是第七年你要讓地歇息，不耕不種，使你百姓中的貧窮人有吃的；他們吃剩的，野獸可以吃。你的葡萄園和橄欖園也要照樣辦理。
EXOD|23|12|「六日你要做工，第七日要安息，使牛、驢可以歇息，也讓你使女的兒子和寄居的可以恢復精力。
EXOD|23|13|「凡我對你們說的話，你們都要謹守。別神的名，你不可提，也不可用口說給人聽。」
EXOD|23|14|「一年三次，你要向我守節。
EXOD|23|15|你要守除酵節，照我所吩咐你的，在亞筆月內所定的日期吃無酵餅七天，因為你是在這月離開了 埃及 。誰也不可空手來朝見我。
EXOD|23|16|你要守收割節，收田間所種、勞碌所得初熟之物。你年底收藏田間勞碌所得時，要守收藏節。
EXOD|23|17|所有的男丁都要一年三次朝見主耶和華。
EXOD|23|18|「不可將我祭牲的血和有酵之物一同獻上，也不可將我節期中祭牲的脂肪留到早晨。
EXOD|23|19|「要把地裏最好的初熟之物帶到耶和華－你上帝的殿中。 「不可用母山羊的奶來煮牠的小山羊。」
EXOD|23|20|「看哪，我要差遣使者在你前面，在路上保護你，領你到我所預備的地方。
EXOD|23|21|你們要在他面前謹慎，聽從他的話。不可抗拒 他，否則他必不赦免你們的過犯，因為我的名在他身上。
EXOD|23|22|「你若真的聽從他的話，照我一切所說的去做，我就以你的仇敵為仇敵，以你的敵人為敵人。
EXOD|23|23|「我的使者要走在你前面，領你到 亞摩利 人、 赫 人、 比利洗 人、 迦南 人、 希未 人、 耶布斯 人那裏，我必將他們除滅。
EXOD|23|24|你不可跪拜事奉他們的神明，也不可隨從他們的習俗，卻要徹底廢除，完全打碎他們的柱像。
EXOD|23|25|你們要事奉耶和華－你們的上帝，他必賜福給你的糧食和水，也必從你中間除去疾病。
EXOD|23|26|你境內必沒有流產的、不生育的。我要使你享滿你年日的數目。
EXOD|23|27|凡你所到的地方，我要使那裏的眾百姓在你面前驚慌失措，又要使你所有的仇敵轉身逃跑。
EXOD|23|28|我要派瘟疫 在你的前面，把 希未 人、 迦南 人、 赫 人從你面前趕出去。
EXOD|23|29|我不在一年之內把他們從你面前趕出去，恐怕地會荒廢，野地的走獸增多危害你。
EXOD|23|30|我要逐漸把他們從你面前趕出去，直到你的人數增多，承受那地為業。
EXOD|23|31|我要定你的疆界，從 紅海 直到 非利士海 ，從曠野直到 大河 。我要把那地的居民交在你手中，你要把他們從你面前趕出去。
EXOD|23|32|不可跟他們和他們的神明立約。
EXOD|23|33|他們不可住在你的地上，免得他們使你得罪我。你若事奉他們的神明，必成為你的圈套。」
EXOD|24|1|耶和華對 摩西 說：「你和 亞倫 、 拿答 、 亞比戶 ，以及 以色列 長老中的七十人，都要上到耶和華這裏來，遠遠地下拜。
EXOD|24|2|只有 摩西 可以接近耶和華，其他的人卻不可接近；百姓也不可和他一同上來。」
EXOD|24|3|摩西 下山，向百姓陳述耶和華一切的命令和典章。眾百姓齊聲說：「耶和華所吩咐的一切，我們都必遵行。」
EXOD|24|4|摩西 將耶和華一切的命令都寫下來。 他清早起來，在山腳築了一座壇，按著 以色列 十二支派立了十二根石柱。
EXOD|24|5|他差派 以色列 的年輕人去獻燔祭，又宰牛獻給耶和華為平安祭。
EXOD|24|6|摩西 將血的一半盛在盆中，另一半灑在壇上。
EXOD|24|7|然後，他拿起約書來，念給百姓聽。他們說：「耶和華所吩咐的一切，我們都必遵行，也必聽從。」
EXOD|24|8|摩西 把血灑在百姓身上，說：「看哪！這是立約的血，是耶和華按照這一切的命令和你們立約的憑據。」
EXOD|24|9|摩西 、 亞倫 、 拿答 、 亞比戶 ，以及 以色列 長老中的七十人都上去，
EXOD|24|10|看見了 以色列 的上帝。在他的腳下，彷彿有藍寶石鋪道，明淨如天。
EXOD|24|11|他不把手伸在 以色列 領袖的身上。他們瞻仰上帝，又吃又喝。
EXOD|24|12|耶和華對 摩西 說：「你上山到我這裏來，就在那裏，我要將石版，就是我所寫的律法和誡命賜給你，使你可以教導他們。」
EXOD|24|13|摩西 和他的助手 約書亞 站起來； 摩西 上了上帝的山。
EXOD|24|14|摩西 對長老們說：「你們在這裏等我們，直到我們再回到你們這裏。看哪， 亞倫 和 戶珥 與你們同在。誰有訴訟，可以去找他們。」
EXOD|24|15|摩西 上山，有雲彩把山遮蓋。
EXOD|24|16|耶和華的榮耀駐在 西奈山 ，雲彩遮蓋了山六天，第七天他從雲中呼叫 摩西 。
EXOD|24|17|耶和華的榮耀在山頂上，在 以色列 人眼前，形狀如吞噬的火。
EXOD|24|18|摩西 進入雲中，登上了山。 摩西 在山上四十晝夜。
EXOD|25|1|耶和華吩咐 摩西 說：
EXOD|25|2|「你要吩咐 以色列 人獻禮物給我。凡甘心樂意獻給我的禮物，你們都可以收下。
EXOD|25|3|要從他們收的禮物是：金、銀、銅，
EXOD|25|4|藍色、紫色、朱紅色紗 ，細麻，山羊毛，
EXOD|25|5|染紅的公羊皮、精美的皮料，金合歡木，
EXOD|25|6|點燈的油，做膏油的香料、做香的香料，
EXOD|25|7|紅瑪瑙與寶石，可以鑲嵌在以弗得和胸袋上。
EXOD|25|8|他們要為我造聖所，使我住在他們中間。
EXOD|25|9|你們要按照我指示你的，帳幕和其中一切器具的樣式，照樣去做。」
EXOD|25|10|「他們要用金合歡木做一個櫃子，長二肘半，寬一肘半，高一肘半。
EXOD|25|11|你要把它裏裏外外包上純金，四圍要鑲上金邊。
EXOD|25|12|要鑄造四個金環，安在櫃子的四腳上；這邊兩個環，那邊兩個環。
EXOD|25|13|要用金合歡木做兩根槓，包上金子。
EXOD|25|14|要把槓穿過櫃旁的環，以便抬櫃。
EXOD|25|15|這槓要留在櫃的環內，不可抽出來。
EXOD|25|16|要把我所要賜給你的法版 放在櫃裏。
EXOD|25|17|要用純金做一個櫃蓋 ，長二肘半，寬一肘半。
EXOD|25|18|要造兩個用金子錘出的基路伯，從櫃蓋的兩端錘出它們。
EXOD|25|19|這端錘出一個基路伯，那端錘出一個基路伯；從櫃蓋的兩端錘出兩個基路伯。
EXOD|25|20|二基路伯的翅膀要向上張開，用翅膀遮住櫃蓋，臉要彼此相對；基路伯的臉要朝向櫃蓋。
EXOD|25|21|要把櫃蓋安在櫃的上邊，又要把我所要賜給你的法版放在櫃裏。
EXOD|25|22|我要在那裏與你相會，並要從法版之櫃的櫃蓋上，兩個基路伯的中間，將我要吩咐 以色列 人的一切事告訴你。」
EXOD|25|23|「你要用金合歡木做一張供桌，長二肘，寬一肘，高一肘半，
EXOD|25|24|把它包上純金，四圍鑲上金邊。
EXOD|25|25|供桌的四圍各做一掌寬的邊緣，邊緣周圍要鑲上金邊。
EXOD|25|26|要為供桌做四個金環，把環安在四個桌腳的四角上。
EXOD|25|27|環要靠近邊緣，以便穿槓抬供桌。
EXOD|25|28|要用金合歡木做兩根槓，包上金子，用來抬供桌。
EXOD|25|29|要用純金做桌上的盤、碟，以及澆酒祭的壺和杯。
EXOD|25|30|要把供餅擺在桌上，常在我面前。」
EXOD|25|31|「要造一座用純金錘出的燈臺。燈臺的座、幹、杯、花萼和花瓣，都要和燈臺接連一塊。
EXOD|25|32|燈臺兩旁要伸出六根枝子：這邊三根，那邊三根。
EXOD|25|33|這邊枝子上有三個杯，形狀像杏花，有花萼有花瓣；那邊枝子上也有三個杯，形狀像杏花，有花萼有花瓣。從燈臺伸出來的六根枝子都是如此。
EXOD|25|34|燈臺本身要有四個杯，形狀像杏花，有花萼有花瓣。
EXOD|25|35|燈臺的第一對枝子下面有花萼，燈臺的第二對枝子下面有花萼，燈臺的第三對枝子下面也有花萼；燈臺伸出的六根枝子都是如此。
EXOD|25|36|花萼和枝子都要和燈臺接連一塊，全是從一塊純金錘出來的。
EXOD|25|37|要做燈臺的七盞燈，燈要點燃，照亮前面。
EXOD|25|38|要用純金做燈剪和燈盤。
EXOD|25|39|做燈臺和這一切的器具要用一他連得純金。
EXOD|25|40|要謹慎，照著在山上指示你的樣式去做。」
EXOD|26|1|「你要用十幅幔子做帳幕。這些幔子要用搓的細麻和藍色、紫色、朱紅色紗織成，並且以刺繡的手藝繡上基路伯。
EXOD|26|2|每幅幔子要長二十八肘，每幅幔子寬四肘，全部的幔子尺寸都要一樣。
EXOD|26|3|這五幅幔子要彼此相連；那五幅也彼此相連。
EXOD|26|4|在這一組相連幔子的末幅邊上要縫藍色的鈕環；在另一組相連幔子的末幅邊上也要照樣做。
EXOD|26|5|這幅幔子上要縫五十個鈕環，另一組相連幔子的末幅上也縫五十個鈕環，環環相對。
EXOD|26|6|要做五十個金鉤，用鉤子使幔子彼此相連，成為一個帳幕。
EXOD|26|7|「你要用山羊毛織十一幅幔子來作帳幕的罩棚。
EXOD|26|8|每幅幔子要長三十肘，每幅幔子寬四肘；十一幅幔子的尺寸都要一樣。
EXOD|26|9|要把五幅幔子連成一幅，又把六幅幔子連成一幅，這第六幅幔子要在罩棚的前面摺上去。
EXOD|26|10|在這一組相連幔子的末幅邊上要縫五十個鈕環；在另一組相連幔子的末幅邊上也縫五十個鈕環。
EXOD|26|11|要做五十個銅鉤，鉤在鈕環中，使罩棚相連成為一個。
EXOD|26|12|罩棚幔子餘下垂著的，那餘下的半幅要垂在帳幕的背面。
EXOD|26|13|罩棚的幔子兩旁所餘下的，這邊一肘，那邊一肘，要垂在帳幕的兩邊，蓋住帳幕。
EXOD|26|14|要用染紅的公羊皮做罩棚的蓋，再用精美皮料做外層的蓋。
EXOD|26|15|「你要用金合歡木做豎立帳幕的木板，
EXOD|26|16|木板要長十肘，每塊板寬一肘半，
EXOD|26|17|每塊板有兩個榫頭可以彼此銜接。帳幕一切的板都要這樣做。
EXOD|26|18|你要做帳幕的木板：南面，就是面向南方的那一邊，要做二十塊板。
EXOD|26|19|在這二十塊板底下要做四十個帶卯眼的銀座；兩個卯眼接連這塊板上的兩個榫頭，另外兩個卯眼接連那塊板上的兩個榫頭。
EXOD|26|20|帳幕的第二邊，就是北面，也要做二十塊板，
EXOD|26|21|和四十個帶卯眼的銀座；這塊板底下有兩個卯眼，那塊板底下也有兩個卯眼。
EXOD|26|22|帳幕的後面，就是西面，要做六塊板。
EXOD|26|23|帳幕後面的角落要做兩塊板。
EXOD|26|24|下端的板是成雙的，上端要連在一起，直到頂端的第一個環子；兩塊板都要這樣，做成兩個角落。
EXOD|26|25|一共有八塊板和十六個帶卯眼的銀座；這塊板底下有兩個卯眼，那塊板底下也有兩個卯眼。
EXOD|26|26|「你要用金合歡木做橫木：為帳幕這面的板做五根橫木，
EXOD|26|27|為帳幕那面的板做五根橫木，又為帳幕後面，就是朝西的板做五根橫木。
EXOD|26|28|板腰間的橫木，要從一頭通到另一頭。
EXOD|26|29|板要包上金子，又要做板上的金環來套橫木；橫木也要包上金子。
EXOD|26|30|要照著在山上所指示你的樣式，把帳幕豎立起來。
EXOD|26|31|「你要用藍色、紫色、朱紅色紗，和搓的細麻織幔子，以刺繡的手藝繡上基路伯。
EXOD|26|32|要把幔子掛在四根包金的金合歡木柱子上，柱子有金鉤，並且安在四個帶卯眼的銀座上。
EXOD|26|33|要把幔子垂掛在鉤子上，把法櫃抬進幔子內；這幔子要將聖所和至聖所隔開。
EXOD|26|34|又要把櫃蓋安在至聖所內的法櫃上，
EXOD|26|35|把供桌安在幔子的外面，供桌在北面，燈臺在帳幕的南面，和供桌相對。
EXOD|26|36|「你要用藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝為帳幕織門簾。
EXOD|26|37|要用金合歡木為簾子做五根柱子，包上金子。柱子有金鉤，又為柱子鑄造五個帶卯眼的銅座。」
EXOD|27|1|「你要用金合歡木做祭壇，長五肘，寬五肘，這壇是正方形的，高三肘。
EXOD|27|2|要在壇的四角做四個翹角，與壇接連一塊；要把壇包上銅。
EXOD|27|3|要做桶子來盛壇上的灰，又要做鏟子、盤子、肉叉和火盆；壇上一切的器具都要用銅做。
EXOD|27|4|要為壇做一個銅網，在網的四角做四個銅環，
EXOD|27|5|把網安在壇四圍的邊的下面，使網垂到壇的半腰。
EXOD|27|6|又要用金合歡木為壇做槓，包上銅。
EXOD|27|7|這槓要穿過壇兩旁的環子，用來抬壇。
EXOD|27|8|要用板做壇，壇的中心是空的，都照著在山上所指示你的樣式做。」
EXOD|27|9|「你要做帳幕的院子。南面，就是面向南方的那一邊，要用搓的細麻做院子的帷幔，長一百肘，
EXOD|27|10|院子要有二十根柱子，二十個帶卯眼的銅座。要用銀做柱子的鉤和箍。
EXOD|27|11|北面的長度也一樣，帷幔長一百肘，要有二十根柱子，二十個帶卯眼的銅座。要用銀做柱子的鉤和箍。
EXOD|27|12|院子的西面有帷幔，寬五十肘，帷幔要有十根柱子，十個帶卯眼的座。
EXOD|27|13|院子的東面，就是面向東方的那一邊，寬五十肘。
EXOD|27|14|一邊的帷幔有十五肘，要有三根柱子，三個帶卯眼的座。
EXOD|27|15|另一邊的帷幔也有十五肘，要有三根柱子，三個帶卯眼的座。
EXOD|27|16|院子的門要有二十肘長的簾子，用藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝織成；要有四根柱子，四個帶卯眼的座。
EXOD|27|17|院子四圍一切的柱子都要用銀子箍著，要用銀做柱子的鉤子，用銅做帶卯眼的座。
EXOD|27|18|院子要長一百肘，寬五十肘 ，高五肘。要用搓的細麻做帷幔，用銅做帶卯眼的座。
EXOD|27|19|帳幕中各樣用途的器具，以及帳幕一切的橛子和院子裏一切的橛子，都要用銅做。」
EXOD|27|20|「你要吩咐 以色列 人，把搗成的純橄欖油拿來給你，用以點燈，使燈經常點著；
EXOD|27|21|在會幕中法櫃前的幔子外， 亞倫 和他的兒子要從晚上到早晨，在耶和華面前照管這燈。這要成為 以色列 人世世代代永遠的定例。」
EXOD|28|1|「你要從 以色列 人中，叫你的哥哥 亞倫 和他的兒子 拿答 、 亞比戶 、 以利亞撒 、 以他瑪 一同親近你，作事奉我的祭司。
EXOD|28|2|你要為你哥哥 亞倫 做聖衣，以示尊嚴和華美。
EXOD|28|3|要吩咐一切心中有智慧的，就是我用智慧的靈所充滿的人，為 亞倫 做衣服，使他分別為聖，作事奉我的祭司。
EXOD|28|4|所要做的是胸袋、以弗得、外袍、織成的內袍、禮冠和腰帶。他們要為你哥哥 亞倫 和他的兒子做聖衣，使他們作祭司事奉我。
EXOD|28|5|要用金色、藍色、紫色、朱紅色紗，和細麻去縫製。
EXOD|28|6|「他們要用金色、藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝做以弗得。
EXOD|28|7|以弗得當有兩條肩帶，接上兩端，使它相連。
EXOD|28|8|以弗得的精緻帶子，要以一樣的手藝，用金色、藍色、紫色、朱紅色紗，和搓的細麻縫製，與以弗得接連在一起。
EXOD|28|9|要取兩塊紅瑪瑙，在上面刻 以色列 兒子的名字：
EXOD|28|10|六個名字在一塊寶石上，六個名字在另一塊寶石上，都按照他們出生的次序。
EXOD|28|11|要以雕刻寶石的手藝，如同刻印章，把 以色列 兒子的名字刻在這兩塊寶石上，並把寶石鑲在金槽裏。
EXOD|28|12|要把這兩塊寶石安在以弗得的兩條肩帶上，為 以色列 人作紀念石。 亞倫 要在耶和華面前把他們的名字帶在兩肩上，作為紀念。
EXOD|28|13|要用金子做兩個槽，
EXOD|28|14|再用純金打兩條鏈子，像編成的繩子一樣，把這編成的金鏈扣在槽上。」
EXOD|28|15|「你要以刺繡的手藝做一個決斷的胸袋，和做以弗得的方法一樣，用金色、藍色、紫色、朱紅色紗，和搓的細麻縫製。
EXOD|28|16|胸袋是正方形的，疊成兩層，長一虎口，寬一虎口。
EXOD|28|17|要在上面鑲四行寶石：第一行是紅寶石、紅璧璽、紅玉；
EXOD|28|18|第二行是綠寶石、藍寶石、金剛石；
EXOD|28|19|第三行是紫瑪瑙、白瑪瑙、紫晶；
EXOD|28|20|第四行是水蒼玉、紅瑪瑙、碧玉。這些都要鑲在金槽中。
EXOD|28|21|這些寶石要有 以色列 十二個兒子的名字，如同刻印章，每一顆有自己的名字，代表十二個支派。
EXOD|28|22|要在胸袋上用純金打鏈子，像編成的繩子一樣。
EXOD|28|23|要為胸袋做兩個金環，把這兩個環安在胸袋的兩端。
EXOD|28|24|要把那兩條編成的金鏈繫在胸袋兩端的兩個環上。
EXOD|28|25|又要把鏈子的另外兩端扣在兩個槽上，安在以弗得前面的肩帶上。
EXOD|28|26|要做兩個金環，安在胸袋的兩端，在以弗得裏面的邊上。
EXOD|28|27|再做兩個金環，安在以弗得前面兩條肩帶的下邊，靠近接縫處，在以弗得精緻帶子的上面。
EXOD|28|28|要用藍色的帶子把胸袋的環與以弗得的環繫住，使胸袋綁在以弗得的精緻帶子上，不致鬆脫。
EXOD|28|29|亞倫 進聖所的時候，要把刻著 以色列 兒子名字的決斷胸袋帶著，放在心上，在耶和華面前常作紀念。
EXOD|28|30|又要將烏陵和土明 放在決斷胸袋裏； 亞倫 進到耶和華面前的時候，要放在心上。這樣， 亞倫 在耶和華面前要把 以色列 人的決斷胸袋常常帶著，放在心上。」
EXOD|28|31|「你要做以弗得的外袍，顏色全是藍的。
EXOD|28|32|袍上方的中間要留一個領口，領口周圍的領邊要以手藝編織而成，好像鎧甲的領口，免得破裂。
EXOD|28|33|袍子下襬，就是下襬的周圍要用藍色、紫色、朱紅色紗做石榴，周圍的石榴中間要有金鈴鐺：
EXOD|28|34|一個金鈴鐺一個石榴，一個金鈴鐺一個石榴，在袍子下襬的周圍。
EXOD|28|35|亞倫 供職的時候要穿這袍。他進入聖所到耶和華面前，以及出來的時候，袍上的鈴聲必被聽見，使他不至於死。
EXOD|28|36|「你要用純金做一面牌，如同刻印章，在上面刻『歸耶和華為聖』。
EXOD|28|37|要用藍色的帶子把牌繫在禮冠上，在禮冠的正前面。
EXOD|28|38|這牌必在 亞倫 的額上， 亞倫 要擔當干犯聖物的罪孽；這聖物是 以色列 人在一切聖禮物上所分別為聖的。這牌要常在他的額上，使他們可以在耶和華面前蒙悅納。
EXOD|28|39|要用細麻編織內袍，用細麻做禮冠，又以刺繡的手藝做腰帶。
EXOD|28|40|「你要為 亞倫 的兒子做內袍、腰帶、頭巾，以示尊嚴和華美。
EXOD|28|41|要把這些給你哥哥 亞倫 和他的兒子穿戴，又要膏他們，授予聖職，使他們分別為聖，作事奉我的祭司。
EXOD|28|42|要用細麻布給他們做褲子來遮掩下體，從腰間直到大腿。
EXOD|28|43|亞倫 和他兒子進入會幕，或接近祭壇，在聖所供職的時候要穿上褲子，免得擔當罪孽而死。這要成為 亞倫 和他後裔永遠的定例。」
EXOD|29|1|「這是你使他們分別為聖，作事奉我的祭司時要做的事：取一頭公牛犢，兩隻無殘疾的公綿羊，
EXOD|29|2|無酵餅、用油調和的無酵餅，和抹油的無酵薄餅；這些餅都要用細麥麵做成。
EXOD|29|3|這些餅要裝在一個籃子裏，用籃子帶來，又把公牛和兩隻公綿羊牽來。
EXOD|29|4|要帶 亞倫 和他兒子到會幕的門口，用水洗他們。
EXOD|29|5|要拿服裝，給 亞倫 穿上內袍和以弗得的外袍，以及以弗得，又帶上胸袋，束上以弗得精緻的帶子。
EXOD|29|6|要把禮冠戴在他頭上，將聖冕加在禮冠上，
EXOD|29|7|把膏油倒在他頭上膏他。
EXOD|29|8|要帶他的兒子來，給他們穿上內袍。
EXOD|29|9|要給 亞倫 和他的兒子束上腰帶，裹上頭巾，他們就憑永遠的定例得祭司的職分。又要授聖職給 亞倫 和他的兒子。
EXOD|29|10|「你要把公牛牽到會幕前， 亞倫 和他的兒子要按手在公牛的頭上。
EXOD|29|11|你要在耶和華面前，在會幕的門口宰這公牛。
EXOD|29|12|要取些公牛的血，用指頭抹在祭壇的四個翹角上，把其餘的血全倒在壇的底座上。
EXOD|29|13|要把所有包著內臟的脂肪、肝上的網油、兩個腎和腎上的脂肪，都燒在壇上。
EXOD|29|14|只是公牛的肉、皮、糞都要在營外用火焚燒；這牛是贖罪祭。
EXOD|29|15|「你要牽一隻公綿羊來， 亞倫 和他兒子要按手在這羊的頭上。
EXOD|29|16|你要宰這羊，把血灑在祭壇的周圍。
EXOD|29|17|再把羊切成肉塊，洗淨內臟和腿，連肉塊和頭放在一處。
EXOD|29|18|要把全羊燒在壇上。這是獻給耶和華的燔祭，是獻給耶和華馨香的火祭。」
EXOD|29|19|「你要把第二隻公綿羊牽來， 亞倫 和他兒子要按手在這羊的頭上。
EXOD|29|20|你要宰這羊，取些血抹在 亞倫 的右耳垂和他兒子的右耳垂上，又抹在他們右手的大拇指和右腳的大腳趾上，然後把其餘的血灑在壇的周圍。
EXOD|29|21|你要取些膏油和壇上的血，彈在 亞倫 和他的衣服上，以及他兒子和他們的衣服上； 亞倫 和他的衣服，他兒子和他們的衣服都成為聖了。
EXOD|29|22|「你要取這羊的脂肪，肥尾巴、包著內臟的脂肪、肝上的網油、兩個腎、腎上的脂肪和右腿，這是聖職禮所獻的公綿羊；
EXOD|29|23|再從耶和華面前那裝無酵餅的籃子中取一個餅、一個油餅和一個薄餅，
EXOD|29|24|把它們都放在 亞倫 的手和他兒子的手上，在耶和華面前搖一搖，作為搖祭。
EXOD|29|25|然後，你要從他們手中接過來，放在燔祭上，一起燒在壇上，作為耶和華面前馨香之氣；這是獻給耶和華的火祭。
EXOD|29|26|「你要取 亞倫 聖職禮所獻公綿羊的胸，在耶和華面前搖一搖，作為搖祭；這份就是你的。
EXOD|29|27|那搖祭的胸和舉祭的腿，就是聖職禮獻公綿羊時所搖的、所舉的，你要使它們分別為聖，是歸給 亞倫 和他兒子的。
EXOD|29|28|這是 亞倫 和他子孫憑永遠的定例從 以色列 人中所應得的；因為這是舉祭，是從 以色列 人的平安祭中取出，作為獻給耶和華的舉祭。
EXOD|29|29|「 亞倫 的聖衣要傳給他的子孫，使他們在受膏和承接聖職的時候穿上。
EXOD|29|30|他的子孫接續他當祭司的，每逢進入會幕在聖所供職的時候，要穿這聖衣七天。
EXOD|29|31|「你要拿聖職禮所獻的公綿羊，在聖處煮牠的肉。
EXOD|29|32|亞倫 和他兒子要在會幕的門口吃這羊的肉和籃子裏的餅。
EXOD|29|33|他們要吃那些用來贖罪之物，好承接聖職，使他們分別為聖。外人不可吃，因為這是聖物。
EXOD|29|34|那聖職禮所獻的肉或餅，若有剩餘留到早晨，就要把剩下的用火燒了，不可再吃，因為這是聖物。
EXOD|29|35|「你要這樣照我一切所吩咐的，向 亞倫 和他兒子行授聖職禮七天。
EXOD|29|36|為了贖罪，每天要獻一頭公牛為贖罪祭。你要為祭壇贖罪，使壇潔淨，並要用膏抹壇，使壇成為聖。
EXOD|29|37|要為壇贖罪七天，使壇成為聖，壇就成為至聖。凡觸摸壇的都成為聖。」
EXOD|29|38|「這是你要獻在壇上的：每天不可間斷地獻兩隻一歲的羔羊；
EXOD|29|39|早晨獻第一隻羔羊，黃昏獻第二隻羔羊。
EXOD|29|40|獻第一隻羔羊時，要同時獻上十分之一伊法細麵，調和四分之一欣搗成的油，再獻四分之一欣酒作澆酒祭。
EXOD|29|41|黃昏你獻第二隻羔羊，要照早晨的素祭和同獻的澆酒祭獻上，作為獻給耶和華馨香的火祭。
EXOD|29|42|這要在耶和華面前，在會幕的門口，作為你們世世代代經常獻的燔祭。我要在那裏與你們 相會，和你說話。
EXOD|29|43|我要在那裏與 以色列 人相會，會幕就要因我的榮耀成為聖。
EXOD|29|44|我要使會幕和祭壇分別為聖，也要使 亞倫 和他的兒子分別為聖，作事奉我的祭司。
EXOD|29|45|我要住在 以色列 人中，作他們的上帝。
EXOD|29|46|他們必知道我是耶和華－他們的上帝，是將他們從 埃及 地領出來的，為要住在他們中間。我是耶和華－他們的上帝 。」
EXOD|30|1|「你要用金合歡木做一座燒香的壇，
EXOD|30|2|長一肘，寬一肘，這壇是正方形的，高二肘。壇的四個翹角與壇接連一塊。
EXOD|30|3|要把壇的上面與壇的四圍，以及壇的四個翹角包上純金；又要在壇的四圍鑲上金邊。
EXOD|30|4|要在壇的兩個對側，金邊下面做兩個金環，用來穿槓抬壇。
EXOD|30|5|要用金合歡木做槓，包上金子。
EXOD|30|6|要把壇放在法櫃前的幔子外，對著法櫃上的櫃蓋，就是我與你相會的地方。
EXOD|30|7|亞倫 要在壇上燒芬芳的香；每早晨整理燈的時候，他都要燒這香。
EXOD|30|8|黃昏點燈的時候， 亞倫 也要燒這香。這是你們世世代代在耶和華面前常燒的香。
EXOD|30|9|在這壇上不可燒別樣的香，不可獻燔祭、素祭，也不可獻澆酒祭。
EXOD|30|10|亞倫 每年一次要為壇的四個翹角贖罪。他每年一次要用贖罪祭的血為壇贖罪，作為世世代代的定例。這壇在耶和華面前是至聖的。」
EXOD|30|11|耶和華吩咐 摩西 說：
EXOD|30|12|「你數點 以色列 人，計算人頭時，被數的每一個人要把他生命的贖價獻給耶和華，免得災殃在數點中臨到他們。
EXOD|30|13|每一個被數的人要按照聖所的舍客勒，付半舍客勒，一舍客勒是二十季拉；這半舍客勒是獻給耶和華的禮物。
EXOD|30|14|每一個被數的人，就是二十歲以上的，要將這禮物獻給耶和華。
EXOD|30|15|富有的不必多付，貧窮的也不可少出，各人都要獻半舍客勒給耶和華，作你們生命的贖價。
EXOD|30|16|你要向 以色列 人收這贖罪的銀子，用在會幕的事工。這要在耶和華面前為 以色列 人作紀念，作你們生命的贖價。」
EXOD|30|17|耶和華吩咐 摩西 說：
EXOD|30|18|「你要用銅做洗濯盆和盆座，用來洗濯。要將盆放在會幕和祭壇的中間，盆裏盛水。
EXOD|30|19|亞倫 和他的兒子要用這盆洗手洗腳。
EXOD|30|20|他們進會幕，或是走近壇前供職，獻火祭給耶和華的時候，必須用水洗濯，免得死亡；
EXOD|30|21|他們要洗手洗腳，免得死亡。這是 亞倫 和他的後裔世世代代永遠的定例。」
EXOD|30|22|耶和華吩咐 摩西 說：
EXOD|30|23|「你要取上等的香料，就是五百舍客勒流質的沒藥、二百五十香肉桂、二百五十香菖蒲，
EXOD|30|24|和五百桂皮，都按照聖所的舍客勒；再取一欣橄欖油，
EXOD|30|25|以做香的方法調和製成聖膏油，它就成為聖膏油。
EXOD|30|26|要用這膏油抹會幕和法櫃，
EXOD|30|27|供桌和供桌的一切器具，燈臺和燈臺的器具 ，以及香壇、
EXOD|30|28|燔祭壇和壇的一切器具，洗濯盆和盆座。
EXOD|30|29|你要使這些分別為聖，成為至聖；凡觸摸它們的都成為聖。
EXOD|30|30|要膏 亞倫 和他的兒子，使他們分別為聖，作事奉我的祭司。
EXOD|30|31|你要吩咐 以色列 人說：『你們要世世代代以這油為我的聖膏油。
EXOD|30|32|不可把這油倒在別人身上，也不可用配製這膏油的方法製成同樣的膏油。這膏油是聖的，你們要以它為聖。
EXOD|30|33|凡調和與此類似的膏油，或將它膏在別人身上的，這人要從百姓中剪除。』」
EXOD|30|34|耶和華吩咐 摩西 說：「你要取香料，就是拿他弗、施喜列、喜利比拿，這些香料再加純乳香，每樣都要相同的分量。
EXOD|30|35|你要用這些加上鹽，以配製香料的方法，製成純淨又神聖的香。
EXOD|30|36|要取一點這香，搗成細的粉，放在會幕中的法櫃前，就是我和你相會的地方。你們要以這香為至聖。
EXOD|30|37|你們不可用這配製的方法為自己做香；要以這香為聖，歸於耶和華。
EXOD|30|38|為要聞香味而配製同樣的香的，這人要從百姓中剪除。」
EXOD|31|1|耶和華吩咐 摩西 說：
EXOD|31|2|「你看，我已經題名召 猶大 支派中 戶珥 的孫子， 烏利 的兒子 比撒列 。
EXOD|31|3|我以上帝的靈充滿他，使他有智慧，有聰明，有知識，能做各樣的工，
EXOD|31|4|能設計圖案，用金、銀、銅製造各物，
EXOD|31|5|又能雕刻鑲嵌用的寶石，雕刻木頭，做各樣的工。
EXOD|31|6|看哪，我委派 但 支派中 亞希撒抹 的兒子 亞何利亞伯 與他同工。凡心裏有智慧的，我更要賜給他們智慧的心，能做我所吩咐你的一切，
EXOD|31|7|就是會幕、法櫃和其上的櫃蓋、會幕中一切的器具、
EXOD|31|8|供桌和供桌的器具、純金的燈臺和燈臺的一切器具、香壇、
EXOD|31|9|燔祭壇和壇的一切器具、洗濯盆與盆座、
EXOD|31|10|供祭司職分用的精緻禮服， 亞倫 祭司的聖衣和他兒子的衣服，
EXOD|31|11|以及膏油和聖所用的芬芳的香。他們都要照我所吩咐的一切去做。」
EXOD|31|12|耶和華對 摩西 說：
EXOD|31|13|「你要吩咐 以色列 人說：『你們務要守我的安息日，因為這是你我之間世世代代的記號，叫你們知道我是耶和華，是使你們分別為聖的。
EXOD|31|14|你們要守安息日，以它為聖日。凡干犯這日的，必被處死；凡在這日做工的，那人必從百姓中剪除。
EXOD|31|15|六日要做工，但第七日是向耶和華守完全安息的安息聖日。凡在安息日做工的，必被處死。』
EXOD|31|16|以色列 人要守安息日，世世代代守安息日為永遠的約。
EXOD|31|17|這是我和 以色列 人之間永遠的記號，因為六日之內耶和華造天地，第七日就安息舒暢。」
EXOD|31|18|耶和華在 西奈山 和 摩西 說完了話，就把兩塊法版交給他，是上帝用指頭寫的石版。
EXOD|32|1|百姓見 摩西 遲遲不下山，就聚集到 亞倫 那裏，對他說：「起來！為我們造神明，在我們前面引路，因為領我們出 埃及 地的那個 摩西 ，我們不知道他遭遇了甚麼事。」
EXOD|32|2|亞倫 對他們說：「你們去摘下你們妻子、兒女耳上的金環，拿來給我。」
EXOD|32|3|眾百姓就摘下他們耳上的金環，拿來給 亞倫 。
EXOD|32|4|亞倫 從他們手裏接過來，用模子塑造它，把它鑄成一頭牛犢。他們就說：「 以色列 啊，這是領你出 埃及 地的神明！」
EXOD|32|5|亞倫 看見，就在牛犢面前築壇。 亞倫 宣告說：「明日要向耶和華守節。」
EXOD|32|6|次日清早，百姓起來獻燔祭和平安祭，就坐下吃喝，起來玩樂。
EXOD|32|7|耶和華吩咐 摩西 ：「下去吧，因為你從 埃及 領上來的百姓已經敗壞了。
EXOD|32|8|他們這麼快偏離了我所吩咐的道，為自己鑄了一頭牛犢，向它跪拜，向它獻祭，說：『 以色列 啊，這就是領你出 埃及 地的神明。』」
EXOD|32|9|耶和華對 摩西 說：「我看這百姓，看哪，他們真是硬著頸項的百姓。
EXOD|32|10|現在，你且由著我，我要向他們發烈怒，滅絕他們，但我要使你成為大國。」
EXOD|32|11|摩西 就懇求耶和華－他的上帝，說：「耶和華啊，你為甚麼向你的百姓發烈怒呢？這百姓是你用大能大力的手從 埃及 地領出來的！
EXOD|32|12|為甚麼讓 埃及 人說：『他領他們出去，是要降災禍給他們，在山中把他們殺了，將他們從地上除滅』呢？求你回心轉意，不發你的烈怒，不降災禍給你的百姓。
EXOD|32|13|求你記念你的僕人 亞伯拉罕 、 以撒 、 以色列 。你曾向他們指著自己起誓說：『我必使你們的後裔像天上的星那樣多，並且我要將所應許的這全地賜給你們的後裔，讓他們永遠承受為業。』」
EXOD|32|14|於是耶和華改變心意，不把所說的災禍降給他的百姓。
EXOD|32|15|摩西 轉身下山，手裏拿著兩塊法版。這版的兩面都寫著字，正面背面都有字。
EXOD|32|16|版是上帝的工作，字是上帝寫的字，刻在版上。
EXOD|32|17|約書亞 一聽見百姓呼喊的聲音，就對 摩西 說：「在營裏有戰爭的聲音。」
EXOD|32|18|摩西 說：「這不是打勝仗的聲音，也不是打敗仗的聲音，我聽見的是歌唱的聲音。」
EXOD|32|19|摩西 走近營前，看見牛犢，又看見人在跳舞，就發烈怒，把兩塊版從手中扔到山下摔碎了。
EXOD|32|20|他將他們所鑄的牛犢用火焚燒，磨得粉碎，撒在水面上，叫 以色列 人喝。
EXOD|32|21|摩西 對 亞倫 說：「這百姓向你做了甚麼呢？你竟使他們陷入大罪中！」
EXOD|32|22|亞倫 說：「求我主不要發烈怒。你知道這百姓，他們是向惡的。
EXOD|32|23|他們對我說：『你為我們造神明，在我們前面引路，因為領我們出 埃及 地的那個 摩西 ，我們不知道他遭遇了甚麼事。』
EXOD|32|24|我對他們說：『凡有金環的可以摘下來』，他們就給了我。我把金環扔在火中，這牛犢就出來了。」
EXOD|32|25|摩西 見百姓放肆，因 亞倫 縱容他們，使這事成了敵人的笑柄，
EXOD|32|26|就站在營門前，說：「凡屬耶和華的人，都到我這裏來！」於是 利未 人都聚集到他那裏。
EXOD|32|27|他對他們說：「耶和華－ 以色列 的上帝這樣說：『你們各人把刀佩在腰間，從這門到那門，來回走遍全營，各人要殺自己的弟兄、鄰舍和親人。』」
EXOD|32|28|利未 人遵照 摩西 的話做了。那一天百姓中倒下的約有三千人。
EXOD|32|29|摩西 說：「今天你們要奉獻自己 來事奉耶和華，因為各人犧牲自己的兒子和弟兄，使耶和華今天賜福給你們。」
EXOD|32|30|第二天， 摩西 對百姓說：「你們犯了大罪。我如今要上耶和華那裏去，或許可以為你們贖罪。」
EXOD|32|31|摩西 回到耶和華那裏，說：「唉！這百姓犯了大罪，為自己造了金的神明。
EXOD|32|32|現在，求你赦免他們的罪；不然，就把我從你所寫的冊上除名。」
EXOD|32|33|耶和華對 摩西 說：「誰得罪我，我就把他從我的冊上除去。
EXOD|32|34|現在你去，領這百姓往我所告訴你的地方去，看哪，我的使者必在你的前面引路。到了該懲罰的時候，我必懲罰他們的罪。」
EXOD|32|35|耶和華降災與百姓，因為他們和 亞倫 一起造了牛犢。
EXOD|33|1|耶和華吩咐 摩西 說：「去，離開這裏，你和你從 埃及 地領出來的百姓要上到我起誓應許給 亞伯拉罕 、 以撒 和 雅各 之地去；我曾對他們說：『我要將這地賜給你的後裔』。
EXOD|33|2|我要差遣使者在你前面，把 迦南 人、 亞摩利 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人趕出
EXOD|33|3|那流奶與蜜之地。但我不與你們上去，因為你們是硬著頸項的百姓，免得我在路上把你們滅絕。」
EXOD|33|4|百姓一聽見這壞的信息，他們就悲哀，沒有人佩戴首飾。
EXOD|33|5|耶和華對 摩西 說：「你對 以色列 人說：『你們是硬著頸項的百姓，我若在你們中間一起上去，只一瞬間，就必把你們滅絕。現在把你們身上的首飾摘下來，我好知道該怎樣處置你們。』」
EXOD|33|6|以色列 人離開 何烈山 以後，就把身上的首飾全都摘下來。
EXOD|33|7|摩西 拿一個帳棚支搭在營外，離營有一段距離，他稱這帳棚為會幕。凡求問耶和華的，就到營外的會幕那裏去。
EXOD|33|8|當 摩西 出營到會幕去的時候，百姓就都起來，各人站在自己帳棚的門口，望著 摩西 ，直到他進了會幕。
EXOD|33|9|摩西 進會幕的時候，雲柱就降下來，停在會幕的門前，耶和華就與 摩西 說話。
EXOD|33|10|眾百姓看見雲柱停在會幕的門前，就都起來，各人在自己帳棚的門口下拜。
EXOD|33|11|耶和華與 摩西 面對面說話，好像人與朋友說話。 摩西 回到營裏去，他的年輕助手 嫩 的兒子 約書亞 卻沒有離開會幕。
EXOD|33|12|摩西 對耶和華說：「看，你曾對我說：『將這百姓領上去』；卻沒有讓我知道你要差派誰與我同去。你還說：『我按你的名認識你，你也在我眼前蒙了恩。』
EXOD|33|13|我如今若在你眼前蒙恩，求你將你的道指示我，使我可以認識你，並在你眼前蒙恩。求你顧念這國是你的子民。」
EXOD|33|14|耶和華說：「我必親自去，讓你安心。」
EXOD|33|15|摩西 說：「你若不親自去，就不要把我們從這裏領上去。
EXOD|33|16|現在，人如何得知我和你的百姓在你眼前蒙恩呢？豈不是因為你與我們同去，使我和你的百姓與地面上的萬民有分別嗎？」
EXOD|33|17|耶和華對 摩西 說：「你所說的這件事，我也會去做，因為你在我眼前蒙了恩，並且我按你的名認識你。」
EXOD|33|18|摩西 說：「求你顯出你的榮耀給我看。」
EXOD|33|19|耶和華說：「我要顯示我一切的美善，在你面前經過，並要在你面前宣告耶和華的名。我要恩待誰就恩待誰，要憐憫誰就憐憫誰。」
EXOD|33|20|他又說：「只是你不能看見我的面，因為沒有人看見我還可以存活。」
EXOD|33|21|耶和華說：「看哪，靠近我這裏有個地方，你可以站在這磐石上。
EXOD|33|22|當我的榮耀經過的時候，我必將你放在磐石縫裏，用我的手掌遮掩你，等我過去，
EXOD|33|23|然後我要將我的手掌收回，你就可以看見我的背，卻看不到我的面。」
EXOD|34|1|耶和華對 摩西 說：「你要鑿出兩塊石版，和先前的一樣；我要把你摔碎的那版上先前所寫的字，寫在這版上。
EXOD|34|2|明日早晨，你要預備好了，上 西奈山 ，在山頂那裏站在我面前。
EXOD|34|3|誰也不可和你上去，整座山都不可見到人，也不可有羊群牛群在山下吃草。」
EXOD|34|4|摩西 就鑿出兩塊石版，和先前的一樣。他清晨起來，遵照耶和華吩咐他的，上 西奈山 去，手裏拿著兩塊石版。
EXOD|34|5|耶和華在雲中降臨，與 摩西 一同站在那裏，宣告耶和華的名。
EXOD|34|6|耶和華在他面前經過，宣告： 「耶和華，耶和華， 有憐憫，有恩惠的上帝， 不輕易發怒， 且有豐盛的慈愛和信實，
EXOD|34|7|為千代的人存留慈愛， 赦免罪孽、過犯和罪惡， 萬不以有罪的為無罪， 必懲罰人的罪， 自父及子，直到三、四代。」
EXOD|34|8|摩西 急忙俯伏在地敬拜，
EXOD|34|9|說：「主啊，我若在你眼前蒙恩，求主在我們中間同行。雖然這是硬著頸項的百姓，求你赦免我們的罪孽和罪惡，接納我們為你的產業。」
EXOD|34|10|耶和華說：「看哪，我要立約，要在你眾百姓面前行奇妙的事，是在全地萬國中未曾做過的。你周圍的萬民要看見我藉著你所行，耶和華可畏懼的作為。
EXOD|34|11|「我今天所吩咐你的，你要謹守。看哪，我要從你面前趕出 亞摩利 人、 迦南 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人。
EXOD|34|12|你要謹慎，不可與你所要去那地的居民立約，免得他們成為你中間的圈套。
EXOD|34|13|你要拆毀他們的祭壇，打碎他們的柱像，砍斷他們的 亞舍拉 。
EXOD|34|14|不可敬拜別神，因為耶和華是忌邪 的上帝，他的名是忌邪者。
EXOD|34|15|你不可與那地的居民立約，因為他們隨從自己的神明行淫；祭他們神明的時候，有人邀請你參加，你就會吃他的祭物。
EXOD|34|16|你為你兒子娶他們的女兒為妻，他們的女兒因著隨從她們的神明行淫，就引誘你的兒子也隨從她們的神明行淫。
EXOD|34|17|「不可為自己鑄造神像。
EXOD|34|18|「你要守除酵節，照我所吩咐你的，在亞筆月內所定的日期吃無酵餅七天，因為你是在亞筆月內出了 埃及 。
EXOD|34|19|「凡頭生的都是我的；無論是牛是羊，一切頭生的公的牲畜都要分別出來 。
EXOD|34|20|頭生的驢可以用羔羊代贖。若不贖牠，就要打斷牠的頸項。凡頭生的兒子都要贖出來。沒有人可以空手來朝見我。
EXOD|34|21|「六日你要做工，第七日要安息，即使在耕種或收割的時候也要安息。
EXOD|34|22|在收割初熟麥子的時候要守七七節，又要在年底守收藏節。
EXOD|34|23|你所有的男丁要一年三次朝見主耶和華－ 以色列 的上帝。
EXOD|34|24|我要從你面前趕走列國，擴張你的疆界。你一年三次上去朝見耶和華－你上帝的時候，必沒有人貪圖你的地。
EXOD|34|25|「不可將我祭牲的血和有酵之物一同獻上。逾越節的祭牲也不可留到早晨。
EXOD|34|26|土地裏上好的初熟之物要奉到耶和華－你上帝的殿。不可用母山羊的奶來煮牠的小山羊。」
EXOD|34|27|耶和華對 摩西 說：「你要將這些話寫上，因為我按這話與你和 以色列 人立約。」
EXOD|34|28|摩西 在耶和華那裏四十晝夜，不吃飯不喝水。他把這約的話，那十條誡命 ，寫在版上。
EXOD|34|29|摩西 下 西奈山 。 摩西 從山上下來的時候，手裏拿著兩塊法版。 摩西 不知道自己臉上的皮膚因耶和華和他說話而發光。
EXOD|34|30|亞倫 和 以色列 眾人看見 摩西 ，看哪，他臉上的皮膚發光，他們就怕靠近他。
EXOD|34|31|摩西 叫他們來， 亞倫 和會眾的官長回到他那裏， 摩西 就跟他們說話。
EXOD|34|32|隨後 以色列 眾人都近前來，他就把耶和華在 西奈山 與他所說的一切話都吩咐他們。
EXOD|34|33|摩西 跟他們說完了話，就用面紗蒙上臉。
EXOD|34|34|但 摩西 進到耶和華面前與他說話的時候，就把面紗揭下，直到出來。 摩西 出來，將所吩咐他的話告訴 以色列 人。
EXOD|34|35|以色列 人看見 摩西 的臉，他臉上的皮膚發光。 摩西 就用面紗蒙上臉，直到他進去與耶和華說話才揭下。
EXOD|35|1|摩西 召集 以色列 全會眾，對他們說：「這是耶和華吩咐你們遵行的事：
EXOD|35|2|六日要做工，第七日你們要奉為向耶和華守完全安息的安息聖日。凡在這日做工的，要被處死。
EXOD|35|3|在安息日這一天，不可在你們一切的住處生火。」
EXOD|35|4|摩西 對 以色列 全會眾說：「這是耶和華所吩咐的話，說：
EXOD|35|5|要從你們當中拿禮物獻給耶和華；凡甘心樂意的，可以把耶和華的禮物拿來，就是金、銀、銅，
EXOD|35|6|藍色、紫色、朱紅色紗，細麻，山羊毛，
EXOD|35|7|染紅的公羊皮，精美的皮料，金合歡木，
EXOD|35|8|點燈的油，做膏油的香料、做香的香料，
EXOD|35|9|紅瑪瑙與寶石，可以鑲嵌在以弗得和胸袋上。」
EXOD|35|10|「你們當中凡心裏有智慧的都要來，製造一切耶和華所吩咐的，
EXOD|35|11|就是帳幕、帳幕的罩棚、帳幕的蓋、鉤子、豎板、橫木、柱子和帶卯眼的座，
EXOD|35|12|櫃子、櫃子的槓、櫃蓋和遮掩的幔子，
EXOD|35|13|供桌、供桌的槓、供桌一切的器具和供餅，
EXOD|35|14|燈臺、燈臺的器具、燈和點燈的油，
EXOD|35|15|香壇、壇的槓、膏油和芬芳的香，帳幕門口的門簾，
EXOD|35|16|燔祭壇、壇的銅網、壇的槓和壇的一切器具，洗濯盆和盆座，
EXOD|35|17|院子的帷幔、柱子、帶卯眼的座和院子的門簾，
EXOD|35|18|帳幕的橛子、院子的橛子和繩子，
EXOD|35|19|以及聖所事奉用的精緻禮服， 亞倫 祭司的聖衣和他兒子的衣服，供祭司職分用。」
EXOD|35|20|以色列 全會眾從 摩西 的面前出去。
EXOD|35|21|凡心受感動，靈被驅策的，都帶耶和華的禮物來，為要造會幕和其中一切的器具，以及縫製聖衣。
EXOD|35|22|凡甘心樂意的，連男帶女都來了，各將金器，就是胸針、耳環、打印的戒指，和項鏈帶來，搖著金器的搖祭獻給耶和華。
EXOD|35|23|凡有藍色、紫色、朱紅色紗、細麻、山羊毛、染紅的公羊皮、精美皮料的，都拿了來；
EXOD|35|24|凡願意獻銀和銅作禮物的，都拿禮物來獻給耶和華；凡有金合歡木可做各種用途的也都拿了來。
EXOD|35|25|凡心中有智慧，可以親手紡織的婦女，也把所紡的藍色、紫色、朱紅色紗，和細麻都拿了來。
EXOD|35|26|凡有智慧，心裏受感動的婦女都來紡山羊毛。
EXOD|35|27|眾官長把紅瑪瑙和寶石，可以鑲嵌在以弗得與胸袋上的，都拿了來，
EXOD|35|28|又拿做香，做膏油，和點燈所需的香料和油來。
EXOD|35|29|以色列 人，無論男女，凡心裏受感動的，都帶甘心祭來獻給耶和華，為要做耶和華藉 摩西 所吩咐的一切工。
EXOD|35|30|摩西 對 以色列 人說：「看， 猶大 支派中 戶珥 的孫子， 烏利 的兒子 比撒列 ，耶和華已經題名召他，
EXOD|35|31|又以上帝的靈充滿他，使他有智慧、聰明、知識，能做各樣的工，
EXOD|35|32|能設計圖案，用金、銀、銅製造各物，
EXOD|35|33|又能雕刻鑲嵌用的寶石，雕刻木頭，做各樣精巧的工。
EXOD|35|34|耶和華又賜給他和 但 支派中， 亞希撒抹 的兒子 亞何利亞伯 能教導人的心。
EXOD|35|35|耶和華使他們的心滿有智慧，能做各樣的工，無論是雕刻的工，圖案設計的工，用藍色、紫色、朱紅色紗，和細麻作刺繡的工，以及編織的工，他們都能勝任，也能設計圖案。」
EXOD|36|1|比撒列 和 亞何利亞伯 ，以及一切心裏有智慧，蒙耶和華賜智慧和聰明，懂得做聖所各樣用途之工的人，都照耶和華所吩咐的去做。
EXOD|36|2|摩西 把 比撒列 和 亞何利亞伯 ，以及那些蒙耶和華賜他心裏有智慧，心受感動願意前來做工的人都召來。
EXOD|36|3|這些人就從 摩西 收了 以色列 人為建造聖所，以及聖所各用途之工而奉獻的禮物。每天早晨，百姓繼續把甘心祭拿來。
EXOD|36|4|凡有智慧能做聖所一切工的人，都各自離開他們原本的工作前來，
EXOD|36|5|對 摩西 說：「百姓送來的禮物很多，已經超過耶和華吩咐建造之工所需要的了。」
EXOD|36|6|摩西 吩咐，他們就在營中傳令說：「無論男女，不必再為聖所的禮物做任何的工。」這樣才使百姓停止，不再拿禮物來，
EXOD|36|7|他們所有的材料已經足夠整個工程之用，而且有餘。
EXOD|36|8|做工的人當中，凡心裏有智慧的，用十幅幔子做帳幕，幔子是用搓的細麻和藍色、紫色、朱紅色紗織成的，並且以刺繡的手藝繡上基路伯。
EXOD|36|9|每幅幔子長二十八肘，每幅幔子寬四肘，全部的幔子都是一樣的尺寸。
EXOD|36|10|他使這五幅幔子彼此相連，又使那五幅幔子彼此相連。
EXOD|36|11|他在這一組相連幔子的末幅邊上縫了藍色的鈕環；在另一組相連幔子的末幅邊上也照樣做。
EXOD|36|12|他在這幅幔子上縫五十個鈕環，在另一組相連幔子的末幅上也縫五十個鈕環，環環相對。
EXOD|36|13|他又做了五十個金鉤，用鉤子使幔子彼此相連，成為一個帳幕。
EXOD|36|14|他用山羊毛織十一幅幔子，作為帳幕上的罩棚。
EXOD|36|15|每幅幔子長三十肘，每幅幔子寬四肘；十一幅幔子都是一樣的尺寸。
EXOD|36|16|他把五幅幔子連成一幅，又把六幅幔子連成一幅。
EXOD|36|17|他在這一組相連幔子的末幅邊上縫了五十個鈕環；在另一組相連幔子的末幅邊上也縫了五十個鈕環。
EXOD|36|18|他又做五十個銅鉤，使罩棚相連成為一個。
EXOD|36|19|他用染紅的公羊皮做罩棚的蓋，再用精美皮料做外層的蓋。
EXOD|36|20|他用金合歡木做豎立帳幕的木板，
EXOD|36|21|木板長十肘，每塊板寬一肘半，
EXOD|36|22|每塊板有兩個榫頭可以彼此銜接。帳幕一切的板都是這樣做。
EXOD|36|23|他做帳幕的木板：南面，就是面向南方的那一邊，做二十塊板，
EXOD|36|24|在這二十塊板底下做了四十個帶卯眼的銀座：兩個卯眼接連這塊板上的兩個榫頭，另外兩個卯眼接連那塊板上的兩個榫頭。
EXOD|36|25|他在帳幕的第二邊，就是北面，也做二十塊板，
EXOD|36|26|和四十個帶卯眼的銀座；這塊板底下有兩個卯眼，那塊板底下也有兩個卯眼。
EXOD|36|27|他在帳幕的後面，就是西面，做六塊板，
EXOD|36|28|在帳幕後面的角落做兩塊板。
EXOD|36|29|下端的板是成雙的，上端連在一起，直到頂端的第一個環子；兩塊板都是這樣，做成兩個角落。
EXOD|36|30|一共有八塊板和十六個帶卯眼的銀座，每塊板底下有兩個卯眼。
EXOD|36|31|他用金合歡木做橫木：為帳幕這面的板做五根橫木，
EXOD|36|32|為帳幕那面的板做五根橫木，又為帳幕後面，就是朝西的板做五根橫木，
EXOD|36|33|他做了板腰間的橫木，從一頭通到另一頭。
EXOD|36|34|他將板包上金子，又做板上的金環來套橫木；橫木也包上金子。
EXOD|36|35|他用藍色、紫色、朱紅色紗，和搓的細麻織幔子，以刺繡的手藝繡上基路伯。
EXOD|36|36|他又用金合歡木為幔子做四根柱子，包上金子，柱子有金鉤，又為柱子鑄了四個帶卯眼的銀座。
EXOD|36|37|他用藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝為帳幕織門簾，
EXOD|36|38|又為簾子做五根柱子和柱子的鉤子，把柱頂和柱子的箍包上金子。柱子有五個帶卯眼的銅座。
EXOD|37|1|比撒列 用金合歡木做一個櫃子，長二肘半，寬一肘半，高一肘半。
EXOD|37|2|裏裏外外包上金子，四圍鑲上金邊。
EXOD|37|3|他又鑄了四個金環，安在櫃子的四腳上；這邊兩個環，那邊兩個環。
EXOD|37|4|他用金合歡木做了兩根槓，包上金子，
EXOD|37|5|又把槓穿過櫃旁的環，以便抬櫃。
EXOD|37|6|他用純金做了一個櫃蓋，長二肘半，寬一肘半，
EXOD|37|7|他造兩個用金子錘出的基路伯，從櫃蓋的兩端錘出它們。
EXOD|37|8|這端一個基路伯，那端一個基路伯；從櫃蓋的兩端錘出兩個基路伯。
EXOD|37|9|二基路伯的翅膀向上張開，用翅膀遮住櫃蓋，臉彼此相對；基路伯的臉朝向櫃蓋。
EXOD|37|10|他用金合歡木做了一張供桌，長二肘，寬一肘，高一肘半，
EXOD|37|11|把它包上純金，四圍鑲上金邊。
EXOD|37|12|供桌的四圍各做了一掌寬的邊緣，邊緣鑲上金邊。
EXOD|37|13|他又鑄了四個金環，把環安在四個桌腳的四角上。
EXOD|37|14|環靠近邊緣，以便穿槓抬供桌。
EXOD|37|15|他用金合歡木做了兩根槓，包上金子，用來抬供桌。
EXOD|37|16|他又用純金做了桌上的器具，就是盤、碟，以及澆酒祭的杯和壺。
EXOD|37|17|他造一座用純金錘出的燈臺；燈臺的座、幹、杯、花萼和花瓣，都和燈臺接連一塊。
EXOD|37|18|燈臺兩旁伸出六根枝子：這邊三根，那邊三根。
EXOD|37|19|這邊的枝子上有三個杯，形狀像杏花，有花萼有花瓣；那邊的枝子上也有三個杯，形狀像杏花，有花萼有花瓣。從燈臺伸出來的六根枝子都是如此。
EXOD|37|20|燈臺本身有四個杯，形狀像杏花，有花萼有花瓣。
EXOD|37|21|燈臺的第一對枝子下面有花萼，燈臺的第二對枝子下面有花萼，燈臺的第三對枝子下面也有花萼；燈臺伸出的六根枝子都是如此。
EXOD|37|22|花萼和枝子都和燈臺接連一塊，全是從一塊純金錘出來的。
EXOD|37|23|他用純金做燈臺的七盞燈，以及燈剪和燈盤。
EXOD|37|24|他用一他連得的純金做燈臺和燈臺的一切器具。
EXOD|37|25|他用金合歡木做香壇，長一肘，寬一肘，這壇是正方形的，高二肘。壇的四個翹角與壇接連一塊。
EXOD|37|26|他把壇的上面與壇的四圍，以及壇的四個翹角包上純金，又在壇的四圍鑲上金邊。
EXOD|37|27|他在壇的兩個對側，金邊下面做了兩個金環，用來穿槓抬壇。
EXOD|37|28|他又用金合歡木做槓，包上金子。
EXOD|37|29|他按配製香料的方法製成聖膏油和芬芳的純香。
EXOD|38|1|他用金合歡木做燔祭壇，長五肘，寬五肘，是正方形的，高三肘。
EXOD|38|2|在壇的四角做四個翹角，與壇接連一塊，把壇包上銅。
EXOD|38|3|他做壇的一切器具，就是桶子、鏟子、盤子、肉叉和火盆；這一切器具都是用銅做的。
EXOD|38|4|他又為壇做一個銅網，安在壇四圍的邊的下面，垂到壇的半腰。
EXOD|38|5|他在銅網的四角上鑄了四個環，用來穿槓。
EXOD|38|6|他用金合歡木做槓，包上銅，
EXOD|38|7|把槓穿過壇兩旁的環子，用來抬壇。他用板做壇，壇的中心是空的。
EXOD|38|8|他用銅做洗濯盆和盆座，是用會幕門前事奉之婦人的銅鏡做的。
EXOD|38|9|他又做院子，在南面，就是面向南方的那一邊，用搓的細麻做院子的帷幔，一百肘。
EXOD|38|10|帷幔有二十根柱子，二十個帶卯眼的銅座；柱子的鉤和箍都是銀的。
EXOD|38|11|北面的帷幔一百肘。帷幔有二十根柱子，二十個帶卯眼的銅座；柱子的鉤和箍都是銀的。
EXOD|38|12|西面的帷幔五十肘。帷幔有十根柱子，十個帶卯眼的座；柱子的鉤和箍都是銀的。
EXOD|38|13|院子的東面，就是面向東方的那一邊，五十肘。
EXOD|38|14|一邊的帷幔有十五肘，有三根柱子，三個帶卯眼的座。
EXOD|38|15|另一邊也一樣，院子門口左右的帷幔也有十五肘，有三根柱子，三個帶卯眼的座。
EXOD|38|16|院子四面的帷幔都是用搓的細麻做的。
EXOD|38|17|柱子帶卯眼的座是銅的，柱子的鉤和箍是銀的，柱頂是用銀包的。院子一切的柱子都是用銀子箍著的。
EXOD|38|18|院子的門簾是以刺繡的手藝，用藍色、紫色、朱紅色紗，和搓的細麻織的，長二十肘，寬也就是高五肘，與院子帷幔的高度相同。
EXOD|38|19|門簾有四根柱子，四個帶卯眼的銅座；柱子上的鉤和箍是銀的，柱頂是用銀包的。
EXOD|38|20|帳幕一切的橛子和院子四圍的橛子都是銅的。
EXOD|38|21|這是帳幕，就是法櫃帳幕中物件的總數，是照 摩西 的吩咐， 亞倫 祭司的兒子 以他瑪 經手， 利未 人數點的。
EXOD|38|22|凡耶和華吩咐 摩西 的，都是由 猶大 支派中 戶珥 的孫子， 烏利 的兒子 比撒列 去做的；
EXOD|38|23|與他同工的有 但 支派中 亞希撒抹 的兒子 亞何利亞伯 ；他是雕刻師，也是設計師，又是用藍色、紫色、朱紅色紗，和細麻的刺繡師。
EXOD|38|24|為聖所一切工作用的金子，就是所奉獻的金子，按聖所的舍客勒，一共是二十九他連得，七百三十舍客勒。
EXOD|38|25|會中被數的人所獻的銀子，按聖所的舍客勒，一共是一百他連得，一千七百七十五舍客勒。
EXOD|38|26|凡曾被數的，就是二十歲以上的人，共有六十萬三千五百五十人。按聖所的舍客勒，每人半舍客勒，就是一比加。
EXOD|38|27|一百他連得銀子是用來鑄造聖所帶卯眼的座和幔子下帶卯眼的座；用一百他連得鑄造一百個帶卯眼的座，每個帶卯眼的座一他連得。
EXOD|38|28|一千七百七十五舍客勒是用來鑄造柱子的鉤，包柱頂，以及箍著柱子。
EXOD|38|29|所奉獻的銅共有七十他連得，二千四百舍客勒。
EXOD|38|30|這些銅是用來做會幕門口帶卯眼的座，銅壇、壇的銅網和壇的一切器具，
EXOD|38|31|院子四圍帶卯眼的座和院子門口帶卯眼的座，以及帳幕一切的橛子和院子四圍所有的橛子。
EXOD|39|1|他們用藍色、紫色、朱紅色紗縫製精緻的禮服，在聖所用以供職；他們為 亞倫 做聖衣，是照耶和華所吩咐 摩西 的。
EXOD|39|2|以弗得是用金色、藍色、紫色、朱紅色紗，和搓的細麻做的。
EXOD|39|3|他們把金子錘成薄片，剪成細線，與藍色、紫色、朱紅色紗，以刺繡的手藝織在一起。
EXOD|39|4|他們又為以弗得做兩條相連的肩帶，接連在以弗得的兩端。
EXOD|39|5|以弗得的精緻帶子以一樣的手藝，用金色、藍色、紫色、朱紅色紗，和搓的細麻縫製，與以弗得接連在一起，是照耶和華所吩咐 摩西 的。
EXOD|39|6|他們琢出兩塊紅瑪瑙，鑲在金槽裏，如同刻印章，刻上 以色列 眾子的名字。
EXOD|39|7|他把這兩塊寶石安在以弗得的兩條肩帶上，為 以色列 人作紀念石，是照耶和華所吩咐 摩西 的。
EXOD|39|8|胸袋是以刺繡的手藝，如同以弗得的做法，用金色、藍色、紫色、朱紅色紗，和搓的細麻縫製。
EXOD|39|9|胸袋是正方形的，他們把它做成兩層，這兩層各長一虎口，寬一虎口。
EXOD|39|10|他們在上面鑲四行寶石：第一行是紅寶石、紅璧璽、紅玉；
EXOD|39|11|第二行是綠寶石、藍寶石、金剛石；
EXOD|39|12|第三行是紫瑪瑙、白瑪瑙、紫晶；
EXOD|39|13|第四行是水蒼玉、紅瑪瑙、碧玉。這些都鑲在金槽中。
EXOD|39|14|這些寶石有 以色列 十二個兒子的名字，如同刻印章，每一顆有自己的名字，代表十二個支派。
EXOD|39|15|他們在胸袋上用純金打鏈子，像編成的繩子一樣。
EXOD|39|16|他們又做了兩個金槽和兩個金環，把這兩個環安在胸袋的兩端。
EXOD|39|17|他們把那兩條編成的金鏈繫在胸袋兩端的兩個環上，
EXOD|39|18|又把鏈子的另外兩端扣在兩個槽上，安在以弗得前面的肩帶上。
EXOD|39|19|他們做了兩個金環，安在胸袋的兩端，在以弗得裏面的邊上，
EXOD|39|20|又做兩個金環，安在以弗得前面兩條肩帶的下邊，靠近接縫處，在精緻帶子的上面。
EXOD|39|21|他們用藍色的帶子把胸袋的環與以弗得的環繫住，使胸袋綁在以弗得精緻的帶子上，不致鬆脫，是照耶和華所吩咐 摩西 的。
EXOD|39|22|以弗得的外袍是以編織的手藝做的，顏色全是藍的。
EXOD|39|23|袍上方的中間留了一個領口，領口的周圍織出領邊，好像鎧甲的領口，免得破裂。
EXOD|39|24|他們在袍子下襬用藍色、紫色、朱紅色紗，和搓的細麻 做石榴，
EXOD|39|25|又用純金鑄了鈴鐺，把鈴鐺釘在石榴中間，袍子下襬周圍的石榴中間：
EXOD|39|26|一個鈴鐺一個石榴，一個鈴鐺一個石榴，在袍子下襬的周圍，用以供職，是照耶和華所吩咐 摩西 的。
EXOD|39|27|他們用編織的工為 亞倫 和他的兒子做細麻布內袍、
EXOD|39|28|細麻布禮冠、細麻布精緻頭巾，和搓的細麻布褲子，
EXOD|39|29|又用藍色、紫色、朱紅色紗，和搓的細麻，以刺繡的手藝做腰帶，是照耶和華所吩咐 摩西 的。
EXOD|39|30|他們用純金做一面聖冠上的牌，如同刻印章，在上面寫著「歸耶和華為聖」，
EXOD|39|31|又用藍色的帶子把牌繫在禮冠上，是照耶和華所吩咐 摩西 的。
EXOD|39|32|會幕的帳幕一切的工程就這樣做完了。凡耶和華所吩咐 摩西 的， 以色列 人都照樣做了。
EXOD|39|33|他們把帳幕運到 摩西 那裏，帳幕和帳幕的一切器具，就是鉤、板、橫木、柱子、帶卯眼的座，
EXOD|39|34|染紅公羊皮的蓋、精美皮料的蓋、遮掩的幔子，
EXOD|39|35|法櫃、櫃的槓、櫃蓋，
EXOD|39|36|供桌、供桌的一切器具、供餅，
EXOD|39|37|純金的燈臺、擺列的燈、燈臺的一切器具、點燈的油，
EXOD|39|38|金壇、膏油、芬芳的香、帳幕的門簾，
EXOD|39|39|銅壇、壇的銅網、壇的槓、壇的一切器具，洗濯盆和盆座，
EXOD|39|40|院子的帷幔、柱子、帶卯眼的座、院子的門簾、繩子、橛子，帳幕，就是會幕使用的一切器具，
EXOD|39|41|以及聖所事奉用的精緻禮服， 亞倫 祭司的聖衣和他兒子的衣服，供祭司職分用。
EXOD|39|42|這一切工作都是 以色列 人照耶和華所吩咐 摩西 做的。
EXOD|39|43|摩西 看見這一切的工，看哪，耶和華怎樣吩咐，他們就照樣做了， 摩西 就為他們祝福。
EXOD|40|1|耶和華吩咐 摩西 說：
EXOD|40|2|「正月初一，你要立起會幕的帳幕，
EXOD|40|3|把法櫃安放在裏面，用幔子將櫃遮掩。
EXOD|40|4|把供桌搬進去，擺設桌上的器具。又把燈臺搬進去，點上燈。
EXOD|40|5|把金香壇安在法櫃前，掛上帳幕的門簾。
EXOD|40|6|把燔祭壇安在會幕的帳幕門前。
EXOD|40|7|把洗濯盆安在會幕和壇的中間，在盆裏盛水。
EXOD|40|8|又要在院子周圍支起帷幔，把院子的門簾掛上。
EXOD|40|9|你要用膏油抹帳幕和其中所有的，使帳幕和一切器具分別為聖，就都成為聖。
EXOD|40|10|又要抹燔祭壇和壇的一切器具，使壇分別為聖，壇就成為至聖。
EXOD|40|11|要抹洗濯盆和盆座，使盆分別為聖。
EXOD|40|12|你要帶 亞倫 和他兒子到會幕門口，用水洗身。
EXOD|40|13|要給 亞倫 穿上聖衣，又膏他，使他分別為聖，作事奉我的祭司。
EXOD|40|14|又要帶他的兒子來，給他們穿上內袍。
EXOD|40|15|你怎樣膏他們的父親，也要照樣膏他們，使他們成為事奉我的祭司。他們受了膏，就必世世代代永遠得祭司的職分。」
EXOD|40|16|摩西 這樣做了；耶和華怎樣吩咐 摩西 ，他就照樣做了。
EXOD|40|17|第二年正月初一，帳幕就立起來。
EXOD|40|18|摩西 支起帳幕，安上帶卯眼的座，安上板，穿上橫木，立起柱子。
EXOD|40|19|他在帳幕的上面搭上罩棚，把罩棚外層的蓋子蓋在其上，是照著耶和華所吩咐他的。
EXOD|40|20|他把法版放在櫃裏，把槓穿在櫃的兩旁，把櫃蓋安在櫃上。
EXOD|40|21|把櫃抬進帳幕，掛上遮掩櫃的幔子，把法櫃遮蓋了，是照耶和華所吩咐 摩西 的。
EXOD|40|22|他把供桌安在會幕內，在帳幕的北邊，幔子的外面。
EXOD|40|23|把餅擺設在供桌上，在耶和華面前，是照耶和華所吩咐 摩西 的。
EXOD|40|24|他把燈臺安在會幕內，在帳幕的南邊，供桌的對面，
EXOD|40|25|並在耶和華面前點燈，是照耶和華所吩咐 摩西 的。
EXOD|40|26|他把金壇安在會幕內，幔子的前面，
EXOD|40|27|又在壇上燒芬芳的香，是照耶和華所吩咐 摩西 的。
EXOD|40|28|他又掛上帳幕的門簾。
EXOD|40|29|在會幕的帳幕門口安設燔祭壇，把燔祭和素祭獻在壇上，是照耶和華所吩咐 摩西 的。
EXOD|40|30|他又把洗濯盆安在會幕和祭壇的中間，盆裏盛水，以便洗濯。
EXOD|40|31|摩西 和 亞倫 ，以及 亞倫 的兒子用這盆洗手洗腳。
EXOD|40|32|他們進會幕或走近壇的時候，就都洗濯，是照耶和華所吩咐 摩西 的。
EXOD|40|33|他在帳幕和祭壇的四圍支起院子的帷幔，把院子的門簾掛上。這樣， 摩西 就做完了工。
EXOD|40|34|那時，雲彩遮蓋會幕，耶和華的榮光充滿了帳幕。
EXOD|40|35|摩西 不能進會幕，因為雲彩停在其上，耶和華的榮光充滿了帳幕。
EXOD|40|36|每逢雲彩從帳幕升上去， 以色列 人就起程前行；
EXOD|40|37|雲彩若不升上去，他們就不起程，直等到雲彩升上去。
EXOD|40|38|在他們所行的路上，在 以色列 全家的眼前，白天，耶和華的雲彩在帳幕上，黑夜，有火在雲彩中。
