JOHN|1|1|Споконвіку було Слово, а Слово в Бога було, і Бог було Слово.
JOHN|1|2|Воно в Бога було споконвіку.
JOHN|1|3|Усе через Нього повстало, і ніщо, що повстало, не повстало без Нього.
JOHN|1|4|І життя було в Нім, а життя було Світлом людей.
JOHN|1|5|А Світло у темряві світить, і темрява не обгорнула його.
JOHN|1|6|Був один чоловік, що від Бога був посланий, йому ймення Іван.
JOHN|1|7|Він прийшов на свідоцтво, щоб засвідчити про Світло, щоб повірили всі через нього.
JOHN|1|8|Він тим Світлом не був, але свідчити мав він про Світло.
JOHN|1|9|Світлом правдивим був Той, Хто просвічує кожну людину, що приходить на світ.
JOHN|1|10|Воно в світі було, і світ через Нього повстав, але світ не пізнав Його.
JOHN|1|11|До свого Воно прибуло, та свої відцурались Його.
JOHN|1|12|А всім, що Його прийняли, їм владу дало дітьми Божими стати, тим, що вірять у Ймення Його,
JOHN|1|13|що не з крови, ані з пожадливости тіла, ані з пожадливости мужа, але народились від Бога.
JOHN|1|14|І Слово сталося тілом, і перебувало між нами, повне благодаті та правди, і ми бачили славу Його, славу як Однородженого від Отця.
JOHN|1|15|Іван свідчить про Нього, і кликав, говорячи: Це був Той, що про Нього казав я: Той, Хто прийде за мною, існував передо мною, бо був перше, ніж я.
JOHN|1|16|А з Його повноти ми одержали всі, а то благодать на благодать.
JOHN|1|17|Закон бо через Мойсея був даний, а благодать та правда з'явилися через Ісуса Христа.
JOHN|1|18|Ніхто Бога ніколи не бачив, Однороджений Син, що в лоні Отця, Той Сам виявив був.
JOHN|1|19|А це ось свідоцтво Іванове, як юдеї послали були з Єрусалиму священиків та Левитів, щоб спитали його: Хто ти такий?
JOHN|1|20|І він визнав, і не зрікся, а визнав: Я не Христос.
JOHN|1|21|І запитали його: А хто ж? Чи Ілля? І відказує: Ні! Чи пророк? І дав відповідь: Ні!
JOHN|1|22|Сказали ж йому: Хто ж ти такий? щоб дати відповідь тим, хто послав нас. Що ти кажеш про себе самого?
JOHN|1|23|Відказав: Я голос того, хто кличе: В пустині рівняйте дорогу Господню, як Ісая пророк заповів.
JOHN|1|24|Посланці ж із фарисеїв були.
JOHN|1|25|І вони запитали його та сказали йому: Для чого ж ти христиш, коли ти не Христос, ні Ілля, ні пророк?
JOHN|1|26|Відповів їм Іван, промовляючи: Я водою хрищу, а між вами стоїть, що Його ви не знаєте.
JOHN|1|27|Він Той, Хто за мною йде, Хто до мене був, Кому розв'язати ремінця від узуття Його я негідний.
JOHN|1|28|Це в Віфанії діялося, на тім боці Йордану, де христив був Іван.
JOHN|1|29|Наступного дня Іван бачить Ісуса, що до нього йде, та й каже: Оце Агнець Божий, що на Себе гріх світу бере!
JOHN|1|30|Це Той, що про Нього казав я: За мною йде Муж, що передо мною Він був, бо був перше, ніж я.
JOHN|1|31|І не знав я Його; та для того прийшов я, христивши водою, щоб Ізраїлеві Він з'явився.
JOHN|1|32|І свідчив Іван, промовляючи: Бачив я Духа, що сходив, як голуб, із неба, та зоставався на Ньому.
JOHN|1|33|І не знав я Його, але Той, Хто христити водою послав мене, мені оповів: Над Ким Духа побачиш, що сходить і зостається на Ньому, це Той, Хто христитиме Духом Святим.
JOHN|1|34|І я бачив, і засвідчив, що Він Божий Син!
JOHN|1|35|Наступного дня стояв знову Іван та двоє з учнів його.
JOHN|1|36|І, поглянувши на Ісуса, що проходив, Він сказав: Ото Агнець Божий!
JOHN|1|37|І почули два учні, як він говорив, та й пішли за Ісусом.
JOHN|1|38|А Ісус обернувся й побачив, що вони йшли за Ним, та й каже до них: Чого ви шукаєте? А вони відказали Йому: Равві перекладене це визначає: Учителю, де Ти живеш?
JOHN|1|39|Він говорить до них: Ходіть і побачте! Ті пішли та й побачили, де Він жив, і в Нього той день перебули. Було ж коло години десятої.
JOHN|1|40|А один із тих двох, що чули від Івана та йшли вслід за Ним, був Андрій, брат Симона Петра.
JOHN|1|41|Він знайшов перше Симона, брата свого, та й говорить до нього: Знайшли ми Месію, що визначає: Христос.
JOHN|1|42|І привів він його до Ісуса. На нього ж споглянувши, промовив Ісус: Ти Симон, син Йонин; будеш званий ти Кифа, що визначає: скеля.
JOHN|1|43|Наступного дня захотів Він піти в Галілею. І знайшов Він Пилипа та й каже йому: Іди за Мною!
JOHN|1|44|А Пилип із Віфсаїди походив, із міста Андрія й Петра.
JOHN|1|45|Пилип Нафанаїла знаходить та й каже йому: Ми знайшли Того, що про Нього писав був Мойсей у Законі й Пророки, Ісуса, сина Йосипового, із Назарету.
JOHN|1|46|І сказав йому Нафанаїл: Та хіба ж може бути з Назарету що добре? Пилип йому каже: Прийди та побач.
JOHN|1|47|Ісус, угледівши Нафанаїла, що до Нього йде, говорить про нього: Ото справді ізраїльтянин, що немає в нім підступу!
JOHN|1|48|Говорить Йому Нафанаїл: Звідки знаєш мене? Ісус відповів і до нього сказав: Я бачив тебе ще давніш, ніж Пилип тебе кликав, як під фіґовим деревом був ти.
JOHN|1|49|Відповів Йому Нафанаїл: Учителю, Ти Син Божий, Ти Цар Ізраїлів!
JOHN|1|50|Ісус відповів і до нього сказав: Через те віриш ти, що сказав Я тобі, що під фіґовим деревом бачив тебе? Більш від цього побачиш!
JOHN|1|51|І Він каже йому: Поправді, поправді кажу вам: Відтепер ви побачите небо відкрите та Анголів Божих, що на Людського Сина підіймаються та спускаються.
JOHN|2|1|А третього дня весілля справляли в Кані Галілейській, і була там Ісусова мати.
JOHN|2|2|На весілля запрошений був теж Ісус та учні Його.
JOHN|2|3|Як забракло ж вина, то мати Ісусова каже до Нього: Не мають вина!
JOHN|2|4|Ісус же відказує їй: Що тобі, жоно, до Мене? Не прийшла ще година Моя!
JOHN|2|5|А мати Його до слуг каже: Зробіть усе те, що Він вам скаже!
JOHN|2|6|Було тут шість камінних посудин на воду, що стояли для очищення юдейського, що відер по дві чи по три вміщали.
JOHN|2|7|Ісус каже до слуг: Наповніть водою посудини. І їх поналивали вщерть.
JOHN|2|8|І Він каже до них: Тепер зачерпніть, і занесіть до весільного старости. І занесли.
JOHN|2|9|Як весільний же староста скуштував воду, що сталась вином, а він не знав, звідки воно, знали ж слуги, що води наливали, то староста кличе тоді молодого
JOHN|2|10|та й каже йому: Кожна людина подає перше добре вино, а як понапиваються, тоді гірше; а ти добре вино аж на досі зберіг...
JOHN|2|11|Такий початок чудам зробив Ісус у Кані Галілейській, і виявив славу Свою. І ввірували в Нього учні Його.
JOHN|2|12|Після цього відправивсь Він Сам, і мати Його, і брати Його, і Його учні до Капернауму, і там перебули небагато днів.
JOHN|2|13|А зближалася Пасха юдейська, і до Єрусалиму подався Ісус.
JOHN|2|14|І знайшов Він, що продавали у храмі волів, і овець, і голубів, та сиділи міняльники.
JOHN|2|15|І, зробивши бича з мотузків, Він вигнав із храму всіх, вівці й воли, а міняльникам гроші розсипав, і поперевертав їм столи.
JOHN|2|16|І сказав продавцям голубів: Заберіть оце звідси, і не робіть із дому Отця Мого дому торгового!
JOHN|2|17|Тоді учні Його згадали, що написано: Ревність до дому Твого з'їдає Мене!
JOHN|2|18|І обізвались юдеї й сказали Йому: Яке нам знамено покажеш, що Ти можеш робити таке?
JOHN|2|19|Ісус відповів і промовив до них: Зруйнуйте цей храм, і за три дні Я поставлю його!
JOHN|2|20|Відказали ж юдеї: Сорок шість літ будувався цей храм, а Ти за три дні поставиш його?
JOHN|2|21|А Він говорив про храм тіла Свого.
JOHN|2|22|Коли ж Він із мертвих воскрес, то учні Його згадали, що Він говорив це, і ввірували в Писання та в слово, що сказав був Ісус.
JOHN|2|23|А як в Єрусалимі Він був у свято Пасхи, то багато-хто ввірували в Його Ймення, побачивши чуда Його, що чинив.
JOHN|2|24|Але Сам Ісус їм не звірявся, бо Сам знав усіх,
JOHN|2|25|і потреби не мав, щоб хто свідчив Йому про людину, бо знав Сам, що в людині було.
JOHN|3|1|Був один чоловік із фарисеїв Никодим на ім'я, начальник юдейський.
JOHN|3|2|Він до Нього прийшов уночі, та й промовив Йому: Учителю, знаємо ми, що прийшов Ти від Бога, як Учитель, бо не може ніхто таких чуд учинити, які чиниш Ти, коли Бог із ним не буде.
JOHN|3|3|Ісус відповів і до нього сказав: Поправді, поправді кажу Я тобі: Коли хто не народиться згори, то не може побачити Божого Царства.
JOHN|3|4|Никодим Йому каже: Як може людина родитися, бувши старою? Хіба може вона ввійти до утроби своїй матері знову й родитись?
JOHN|3|5|Ісус відповів: Поправді, поправді кажу Я тобі: Коли хто не родиться з води й Духа, той не може ввійти в Царство Боже.
JOHN|3|6|Що вродилося з тіла є тіло, що ж уродилося з Духа є дух.
JOHN|3|7|Не дивуйся тому, що сказав Я тобі: Вам необхідно родитись згори.
JOHN|3|8|Дух дихає, де хоче, і його голос ти чуєш, та не відаєш, звідкіля він приходить, і куди він іде. Так буває і з кожним, хто від Духа народжений.
JOHN|3|9|Відповів Никодим і до Нього сказав: Як це статися може?
JOHN|3|10|Ісус відповів і до нього сказав: Ти учитель ізраїльський, то чи ж цього не знаєш?
JOHN|3|11|Поправді, поправді кажу Я тобі: Ми говоримо те, що ми знаємо, а свідчимо про те, що ми бачили, але свідчення нашого ви не приймаєте.
JOHN|3|12|Коли Я говорив вам про земне, та не вірите ви, то як же повірите ви, коли Я говоритиму вам про небесне?
JOHN|3|13|І не сходив на небо ніхто, тільки Той, Хто з неба зійшов, Людський Син, що на небі.
JOHN|3|14|І, як Мойсей підніс змія в пустині, так мусить піднесений бути й Син Людський,
JOHN|3|15|щоб кожен, хто вірує в Нього, мав вічне життя.
JOHN|3|16|Так бо Бог полюбив світ, що дав Сина Свого Однородженого, щоб кожен, хто вірує в Нього, не згинув, але мав життя вічне.
JOHN|3|17|Бо Бог не послав Свого Сина на світ, щоб Він світ засудив, але щоб через Нього світ спасся.
JOHN|3|18|Хто вірує в Нього, не буде засуджений; хто ж не вірує, той вже засуджений, що не повірив в Ім'я Однородженого Сина Божого.
JOHN|3|19|Суд же такий, що світло на світ прибуло, люди ж темряву більш полюбили, як світло, лихі бо були їхні вчинки!
JOHN|3|20|Бо кожен, хто робить лихе, ненавидить світло, і не приходить до світла, щоб не зганено вчинків його.
JOHN|3|21|А хто робить за правдою, той до світла йде, щоб діла його виявились, бо зроблені в Бозі вони.
JOHN|3|22|По цьому прийшов Ісус та учні Його до країни Юдейської, і з ними Він там проживав та христив.
JOHN|3|23|А Іван теж христив в Еноні поблизу Салиму, бо було там багато води; і приходили люди й христились,
JOHN|3|24|бо Іван до в'язниці не був ще посаджений.
JOHN|3|25|І зчинилось змагання Іванових учнів з юдеями про очищення.
JOHN|3|26|І прийшли до Івана вони та й сказали йому: Учителю, Той, Хто був із тобою по той бік Йордану, про Якого ти свідчив, ото христить і Він, і до Нього всі йдуть.
JOHN|3|27|Іван відповів і сказав: Людина нічого приймати не може, як їй з неба не дасться.
JOHN|3|28|Ви самі мені свідчите, що я говорив: я не Христос, але посланий я перед Ним.
JOHN|3|29|Хто має заручену, той молодий. А дружко молодого, що стоїть і його слухає, дуже тішиться з голосу молодого. Така радість моя оце здійснилась!
JOHN|3|30|Він має рости, я ж маліти.
JOHN|3|31|Хто зверху приходить, Той над усіма. Хто походить із землі, то той земний, і говорить поземному. Хто приходить із неба, Той над усіма,
JOHN|3|32|і що бачив і чув, те Він свідчить, та свідоцтва Його не приймає ніхто.
JOHN|3|33|Хто ж прийняв свідоцтво Його, той ствердив тим, що Бог правдивий.
JOHN|3|34|Бо Кого Бог послав, Той Божі слова промовляє, бо Духа дає Бог без міри.
JOHN|3|35|Отець любить Сина, і дав усе в Його руку.
JOHN|3|36|Хто вірує в Сина, той має вічне життя; а хто в Сина не вірує, той життя не побачить а гнів Божий на нім перебуває.
JOHN|4|1|Як Господь же довідався, що почули фарисеї, що Ісус учнів більше збирає та христить, як Іван,
JOHN|4|2|хоч Ісус не христив Сам, а учні Його,
JOHN|4|3|Він покинув Юдею та знову пішов у Галілею.
JOHN|4|4|І потрібно було Самарію Йому переходити.
JOHN|4|5|Отож, прибуває Він до самарійського міста, що зветься Сіхар, недалеко від поля, яке Яків був дав своєму синові Йосипові.
JOHN|4|6|Там же була Яковова криниця. І Ісус, дорогою зморений, сів отак край криниці. Було коло години десь шостої.
JOHN|4|7|Надходить ось жінка одна з Самарії набрати води. Ісус каже до неї: Дай напитись Мені!
JOHN|4|8|Бо учні Його відійшли були в місто, щоб купити поживи.
JOHN|4|9|Тоді каже Йому самарянка: Як же Ти, юдеянин бувши, та просиш напитись від мене, самарянки? Бо юдеї не сходяться із самарянами.
JOHN|4|10|Ісус відповів і промовив до неї: Коли б знала ти Божий дар, і Хто Той, Хто говорить тобі: Дай напитись Мені, ти б у Нього просила, і Він тобі дав би живої води.
JOHN|4|11|Каже жінка до Нього: І черпака в Тебе, Пане, нема, а криниця глибока, звідки ж маєш Ти воду живу?
JOHN|4|12|Чи Ти більший за нашого отця Якова, що нам дав цю криницю, і він сам із неї пив, і сини його, і худоба його?
JOHN|4|13|Ісус відповів і сказав їй: Кожен, хто воду цю п'є, буде прагнути знову.
JOHN|4|14|А хто питиме воду, що Я йому дам, прагнути не буде повік, бо вода, що Я йому дам, стане в нім джерелом тієї води, що тече в життя вічне.
JOHN|4|15|Каже жінка до Нього: Дай мені, Пане, цієї води, щоб я пити не хотіла, і сюди не приходила брати.
JOHN|4|16|Говорить до неї Ісус: Іди, поклич чоловіка свого та й вертайся сюди.
JOHN|4|17|Жінка відповіла та й сказала: Чоловіка не маю... Відказав їй Ісус: Ти добре сказала: Чоловіка не маю.
JOHN|4|18|Бо п'ятьох чоловіків ти мала, а той, кого маєш тепер, не муж він тобі. Це ти правду сказала.
JOHN|4|19|Каже жінка до Нього: Бачу, Пане, що Пророк Ти.
JOHN|4|20|Отці наші вклонялися Богу на цій ось горі, а ви твердите, що в Єрусалимі те місце, де потрібно вклонятись.
JOHN|4|21|Ісус промовляє до неї: Повір, жінко, Мені, що надходить година, коли ні на горі цій, ані в Єрусалимі вклонятись Отцеві не будете ви.
JOHN|4|22|Ви вклоняєтесь тому, чого ви не знаєте, ми вклоняємось тому, що знаємо, бо спасіння від юдеїв.
JOHN|4|23|Але наступає година, і тепер вона є, коли богомільці правдиві вклонятися будуть Отцеві в дусі та в правді, бо Отець Собі прагне таких богомільців.
JOHN|4|24|Бог є Дух, і ті, що Йому вклоняються, повинні в дусі та в правді вклонятись.
JOHN|4|25|Відказує жінка Йому: Я знаю, що прийде Месія, що зветься Христос, як Він прийде, то все розповість нам.
JOHN|4|26|Промовляє до неї Ісус: Це Я, що розмовляю з тобою...
JOHN|4|27|І тоді надійшли Його учні, і дивувались, що з жінкою Він розмовляв. Проте жаден із них не спитав: Чого хочеш? або: Про що з нею говориш?
JOHN|4|28|Покинула жінка тоді водоноса свого, і побігла до міста, та й людям говорить:
JOHN|4|29|Ходіть но, побачте Того Чоловіка, що сказав мені все, що я вчинила. Чи Він не Христос?
JOHN|4|30|І вони повиходили з міста, і до Нього прийшли.
JOHN|4|31|Тим часом же учні просили Його та й казали: Учителю, їж!
JOHN|4|32|А Він їм відказав: Я маю поживу на їдження, якої не знаєте ви.
JOHN|4|33|Питали тоді один одного учні: Хіба хто приніс Йому їсти?
JOHN|4|34|Ісус каже до них: Пожива Моя чинити волю Того, Хто послав Мене, і справу Його довершити.
JOHN|4|35|Чи не кажете ви: Ще чотири от місяці, і настануть жнива? А Я вам кажу: Підійміть свої очі, та гляньте на ниви, як для жнив уже пополовіли вони!
JOHN|4|36|А хто жне, той заплату бере, та збирає врожай в життя вічне, щоб хто сіє й хто жне разом раділи.
JOHN|4|37|Бо про це поговірка правдива: Хто інший сіє, а хто інший жне.
JOHN|4|38|Я вас жати послав, де ви не працювали: працювали інші, ви ж до їхньої праці ввійшли.
JOHN|4|39|З того ж міста багато-хто із самарян в Нього ввірували через слово жінки, що свідчила: Він сказав мені все, що я вчинила була!
JOHN|4|40|А коли самаряни до Нього прийшли, то благали Його, щоб у них позостався. І Він перебув там два дні.
JOHN|4|41|Значно ж більш вони ввірували через слово Його.
JOHN|4|42|А до жінки казали вони: Не за слово твоє ми вже віруємо, самі бо ми чули й пізнали, що справді Спаситель Він світу!
JOHN|4|43|Як минуло ж два дні, Він ізвідти пішов в Галілею.
JOHN|4|44|Сам бо свідчив Ісус, що не має пошани пророк у вітчизні своїй.
JOHN|4|45|А коли Він прийшов в Галілею, Його прийняли галілеяни, побачивши все, що вчинив Він в Єрусалимі на святі, бо ходили на свято й вони.
JOHN|4|46|Тоді знову прийшов Ісус у Кану Галілейську, де перемінив був Він воду на вино. І був там один царедворець, що син його хворів у Капернаумі.
JOHN|4|47|Він, почувши, що Ісус із Юдеї прибув в Галілею, до Нього прийшов і благав Його, щоб пішов і сина йому вздоровив, бо мав той умерти.
JOHN|4|48|Ісус же промовив до нього: Як знамен тих та чуд не побачите, не ввіруєте!
JOHN|4|49|Царедворець говорить до Нього: Піди, Господи, поки не вмерла дитина моя!
JOHN|4|50|Промовляє до нього Ісус: Іди, син твій живе! І повірив той слову, що до нього промовив Ісус, і пішов.
JOHN|4|51|А коли ще в дорозі він був, то раби його перестріли його й сповістили, говорячи: Син твій живе.
JOHN|4|52|А він їх запитав про годину, о котрій стало легше йому. Вони ж відказали до нього: Учора о сьомій годині гарячка покинула його.
JOHN|4|53|Зрозумів тоді батько, що була то година, о котрій до нього промовив Ісус: Син твій живе. І ввірував сам і ввесь його дім.
JOHN|4|54|Це знов друге знамено Ісус учинив, як вернувся до Галілеї з Юдеї.
JOHN|5|1|Після того юдейське Свято було, і до Єрусалиму Ісус відійшов.
JOHN|5|2|А в Єрусалимі, біля брами Овечої, є купальня, Віфесда по-єврейському зветься, що мала п'ять ґанків.
JOHN|5|3|У них лежало багато слабих, сліпих, кривих, сухих, що чекали, щоб воду порушено.
JOHN|5|4|Бо Ангол Господній часами спускавсь до купальні, і порушував воду, і хто перший улазив, як воду порушено, той здоровим ставав, хоч би яку мав хворобу.
JOHN|5|5|А був там один чоловік, що тридцять і вісім років був недужим.
JOHN|5|6|Як Ісус його вгледів, що лежить, та, відаючи, що багато він часу слабує, говорить до нього: Хочеш бути здоровим?
JOHN|5|7|Відповів Йому хворий: Пане, я не маю людини, щоб вона, як порушено воду, до купальні всадила мене. А коли я приходжу, то передо мною вже інший улазить.
JOHN|5|8|Говорить до нього Ісус: Уставай, візьми ложе своє та й ходи!
JOHN|5|9|І зараз одужав оцей чоловік, і взяв ложе своє та й ходив. Того ж дня субота була,
JOHN|5|10|тому то сказали юдеї вздоровленому: Є субота, і не годиться тобі брати ложа свого.
JOHN|5|11|А він відповів їм: Хто мене вздоровив, Той до мене сказав: Візьми ложе своє та й ходи.
JOHN|5|12|А вони запитали його: Хто Той Чоловік, що до тебе сказав: Візьми ложе своє та й ходи?
JOHN|5|13|Та не знав уздоровлений, Хто то Він, бо Ісус ухиливсь від народу, що був на тім місці.
JOHN|5|14|Після того Ісус стрів у храмі його, та й промовив до нього: Ось видужав ти. Не гріши ж уже більше, щоб не сталось тобі чого гіршого!
JOHN|5|15|Чоловік же пішов і юдеям звістив, що Той, Хто вздоровив його, то Ісус.
JOHN|5|16|І тому зачали юдеї переслідувати Ісуса, що таке Він чинив у суботу.
JOHN|5|17|А Ісус відповів їм: Отець Мій працює аж досі, працюю і Я.
JOHN|5|18|І тому то юдеї ще більш намагалися вбити Його, що не тільки суботу порушував Він, але й Бога Отцем Своїм звав, тим роблячись Богові рівним.
JOHN|5|19|Відповів же Ісус і сказав їм: Поправді, поправді кажу вам: Син нічого робити не може Сам від Себе, тільки те, що Він бачить, що робить Отець; бо що робить Він, те так само й Син робить.
JOHN|5|20|Бо Отець любить Сина, і показує все, що Сам робить, Йому. І покаже Йому діла більші від цих, щоб ви дивувались.
JOHN|5|21|Бо як мертвих Отець воскрешає й оживлює, так і Син, кого хоче, оживлює.
JOHN|5|22|Бо Отець і не судить нікого, а ввесь суд віддав Синові,
JOHN|5|23|щоб усі шанували і Сина, як шанують Отця. Хто не шанує Сина, не шанує Отця, що послав Його.
JOHN|5|24|Поправді, поправді кажу вам: Хто слухає слова Мого, і вірує в Того, Хто послав Мене, життя вічне той має, і на суд не приходить, але перейшов він від смерти в життя.
JOHN|5|25|Поправді, поправді кажу вам: Наступає година, і тепер уже є, коли голос Божого Сина почують померлі, а ті, що почують, оживуть.
JOHN|5|26|Бо як має Отець життя Сам у Собі, так і Синові дав життя мати в Самому Собі.
JOHN|5|27|І Він дав Йому силу чинити і суд, бо Він Людський Син.
JOHN|5|28|Не дивуйтесь цьому, бо надходить година, коли всі, хто в гробах, Його голос почують,
JOHN|5|29|і повиходять ті, що чинили добро, на воскресення життя, а котрі зло чинили, на воскресення Суду.
JOHN|5|30|Я нічого не можу робити Сам від Себе. Як Я чую, суджу, і Мій суд справедливий, не шукаю бо волі Своєї, але волі Отця, що послав Мене.
JOHN|5|31|Коли свідчу про Себе Я Сам, то свідоцтво Моє неправдиве.
JOHN|5|32|Є Інший, Хто свідчить про Мене, і Я знаю, що правдиве свідоцтво, яким свідчить про Мене.
JOHN|5|33|Ви послали були до Івана, і він свідчив про правду.
JOHN|5|34|Та Я не від людини свідоцтва приймаю, але це говорю, щоб були ви спасені.
JOHN|5|35|Він світильником був, що горів і світив, та ви тільки хвилю хотіли потішитись світлом його.
JOHN|5|36|Але Я маю свідчення більше за Іванове, бо ті справи, що Отець Мені дав, щоб Я виконав їх, ті справи, що Я їх чиню, самі свідчать про Мене, що Отець Мене послав!
JOHN|5|37|Та й Отець, що послав Мене, Сам засвідчив про Мене; але ви ані голосу Його не чули ніколи, ані виду Його не бачили.
JOHN|5|38|Навіть слова Його ви не маєте, щоб у вас перебувало, бо не вірите в Того, Кого Він послав.
JOHN|5|39|Дослідіть но Писання, бо ви думаєте, що в них маєте вічне життя, вони ж свідчать про Мене!
JOHN|5|40|Та до Мене прийти ви не хочете, щоб мати життя.
JOHN|5|41|Від людей не приймаю Я слави,
JOHN|5|42|але вас Я пізнав, що любови до Бога в собі ви не маєте.
JOHN|5|43|Я прийшов у Ймення Свого Отця, та Мене не приймаєте ви. Коли ж прийде інший у ймення своє, того приймете ви.
JOHN|5|44|Як ви можете вірувати, коли славу один від одного приймаєте, а слави тієї, що від Бога Єдиного, не прагнете ви?
JOHN|5|45|Не думайте, що Я перед Отцем буду вас винуватити, є, хто вас винуватити буде, Мойсей, що на нього надієтесь ви!
JOHN|5|46|Коли б ви Мойсеєві вірили, то й Мені б ви повірили, бо про Мене писав він.
JOHN|5|47|Якщо писанням його ви не вірите, то як віри поймете словам Моїм?
JOHN|6|1|Після того Ісус перейшов на той бік Галілейського чи Тіверіядського моря.
JOHN|6|2|А за Ним ішла безліч народу, бо бачили чуда Його, що чинив над недужими.
JOHN|6|3|Ісус же на гору зійшов, і сидів там зо Своїми учнями.
JOHN|6|4|Наближалася ж Пасха, свято юдейське.
JOHN|6|5|А Ісус, звівши очі Свої та побачивши, яка безліч народу до Нього йде, говорить Пилипові: Де ми купимо хліба, щоб вони поживились?
JOHN|6|6|Він же це говорив, його випробовуючи, бо знав Сам, що Він має робити.
JOHN|6|7|Пилип Йому відповідь дав: І за двісті динаріїв їм хліба не стане, щоб кожен із них бодай трохи дістав.
JOHN|6|8|Говорить до Нього Андрій, один з учнів Його, брат Симона Петра:
JOHN|6|9|Є тут хлопчина один, що має п'ять ячних хлібів та дві рибі, але що то на безліч таку!
JOHN|6|10|А Ісус відказав: Скажіть людям сідати! А була на тім місці велика трава. І засіло чоловіка числом із п'ять тисяч.
JOHN|6|11|А Ісус узяв хліби, і, подяку вчинивши, роздав тим, хто сидів. Так само і з риб, скільки хотіли вони.
JOHN|6|12|І, як наїлись вони, Він говорить до учнів Своїх: Позбирайте куски позосталі, щоб ніщо не загинуло.
JOHN|6|13|І зібрали вони. І дванадцять повних кошів наклали кусків, що лишились їдцям із п'яти ячних хлібів.
JOHN|6|14|А люди, що бачили чудо, яке Ісус учинив, гомоніли: Це Той справді Пророк, що повинен прибути на світ!
JOHN|6|15|Спостерігши ж Ісус, що вони мають замір прийти та забрати Його, щоб настановити царем, знов на гору пішов Сам один.
JOHN|6|16|А як вечір настав, то зійшли Його учні над море.
JOHN|6|17|І, ввійшовши до човна, на другий бік моря вони попливли, до Капернауму. І темрява вже наступила була, а Ісус ще до них не приходив.
JOHN|6|18|Від великого ж вітру, що віяв, хвилювалося море.
JOHN|6|19|Як вони ж пропливли стадій із двадцять п'ять або з тридцять, то Ісуса побачили, що йде Він по морю, і до човна зближається, і їх страх обгорнув...
JOHN|6|20|Він же каже до них: Це Я, не лякайтесь!
JOHN|6|21|І хотіли вони взяти до човна Його; та човен зараз пристав до землі, до якої пливли.
JOHN|6|22|А наступного дня той народ, що на тім боці моря стояв, побачив, що там іншого човна, крім одного того, що до нього ввійшли були учні Його, не було, і що до човна не входив Ісус із Своїми учнями, але відпливли самі учні.
JOHN|6|23|А тим часом із Тіверіяди припливли човни інші близько до місця того, де вони їли хліб, як Господь учинив був подяку.
JOHN|6|24|Отож, як побачили люди, що Ісуса та учнів Його там нема, то в човни посідали самі й прибули до Капернауму, і шукали Ісуса.
JOHN|6|25|І, на тім боці моря знайшовши Його, сказали Йому: Коли Ти прибув сюди, Учителю?
JOHN|6|26|Відповів їм Ісус і сказав: Поправді, поправді кажу вам: Мене не тому ви шукаєте, що бачили чуда, а що їли з хлібів і наситились.
JOHN|6|27|Пильнуйте не про поживу, що гине, але про поживу, що зостається на вічне життя, яку дасть нам Син Людський, бо відзначив Його Бог Отець.
JOHN|6|28|Сказали ж до Нього вони: Що ми маємо почати, щоб робити діла Божі?
JOHN|6|29|Ісус відповів і сказав їм: Оце діло Боже, щоб у Того ви вірували, Кого Він послав.
JOHN|6|30|А вони відказали Йому: Яке ж знамено Ти чиниш, щоб побачили ми й поняли Тобі віри? Що Ти робиш?
JOHN|6|31|Наші отці їли манну в пустині, як написано: Хліб із неба їм дав на поживу.
JOHN|6|32|А Ісус їм сказав: Поправді, поправді кажу вам: Не Мойсей хліб із неба вам дав, Мій Отець дає вам хліб правдивий із неба.
JOHN|6|33|Бо хліб Божий є Той, Хто сходить із неба й дає життя світові.
JOHN|6|34|А вони відказали до Нього: Давай, Господи, хліба такого нам завжди!
JOHN|6|35|Ісус же сказав їм: Я хліб життя. Хто до Мене приходить, не голодуватиме він, а хто вірує в Мене, ніколи не прагнутиме.
JOHN|6|36|Але Я вам сказав, що Мене хоч ви й бачили, та не віруєте.
JOHN|6|37|Усе прийде до Мене, що Отець дає Мені, а того, хто до Мене приходить, Я не вижену геть.
JOHN|6|38|Бо Я з неба зійшов не на те, щоб волю чинити Свою, але волю Того, Хто послав Мене.
JOHN|6|39|Оце ж воля Того, Хто послав Мене, щоб з усього, що дав Мені Він, Я нічого не стратив, але воскресив те останнього дня.
JOHN|6|40|Оце ж воля Мого Отця, щоб усякий, хто Сина бачить та вірує в Нього, мав вічне життя, і того воскрешу Я останнього дня.
JOHN|6|41|Тоді стали юдеї ремствувати на Нього, що сказав: Я той хліб, що з неба зійшов.
JOHN|6|42|І казали вони: хіба Він не Ісус, син Йосипів, що ми знаємо батька та матір Його? Як же Він каже: Я з неба зійшов?
JOHN|6|43|А Ісус відповів і промовив до них: Не ремствуйте ви між собою!
JOHN|6|44|Ніхто бо не може до Мене прийти, як Отець, що послав Мене, не притягне його, і того воскрешу Я останнього дня.
JOHN|6|45|У Пророків написано: І всі будуть від Бога навчені. Кожен, хто від Бога почув і навчився, приходить до Мене.
JOHN|6|46|Це не значить, щоб хтось Отця бачив, тільки Той Отця бачив, Хто походить від Бога.
JOHN|6|47|Поправді, поправді кажу Вам: Хто вірує в Мене, життя вічне той має.
JOHN|6|48|Я хліб життя!
JOHN|6|49|Отці ваші в пустині їли манну, і померли.
JOHN|6|50|То є хліб, Який сходить із неба, щоб не вмер, хто Його споживає.
JOHN|6|51|Я хліб живий, що з неба зійшов: коли хто споживатиме хліб цей, той повік буде жити. А хліб, що дам Я, то є тіло Моє, яке Я за життя світові дам.
JOHN|6|52|Тоді між собою змагатися стали юдеї, говорячи: Як же Він може дати нам тіла спожити?
JOHN|6|53|І сказав їм Ісус: Поправді, поправді кажу вам: Якщо ви споживати не будете тіла Сина Людського й пити не будете крови Його, то в собі ви не будете мати життя.
JOHN|6|54|Хто тіло Моє споживає та кров Мою п'є, той має вічне життя, і того воскрешу Я останнього дня.
JOHN|6|55|Бо тіло Моє то правдиво пожива, Моя ж кров то правдиво пиття.
JOHN|6|56|Хто тіло Моє споживає та кров Мою п'є, той в Мені перебуває, а Я в ньому.
JOHN|6|57|Як Живий Отець послав Мене, і живу Я Отцем, так і той, хто Мене споживає, і він житиме Мною.
JOHN|6|58|То є хліб, що з неба зійшов. Не як ваші отці їли манну й померли, хто цей хліб споживає, той жити буде повік!
JOHN|6|59|Оце Він говорив, коли в Капернаумі навчав у синагозі.
JOHN|6|60|А багато-хто з учнів Його, як почули оце, гомоніли: Жорстока це мова! Хто слухати може її?
JOHN|6|61|А Ісус, Сам у Собі знавши це, що учні Його на те ремствують, промовив до них: Чи оце вас спокушує?
JOHN|6|62|А що ж, як побачите Людського Сина, що сходить туди, де перше Він був?
JOHN|6|63|То дух, що оживлює, тіло ж не помагає нічого. Слова, що їх Я говорив вам, то дух і життя.
JOHN|6|64|Але є дехто з вас, хто не вірує. Бо Ісус знав спочатку, хто ті, хто не вірує, і хто видасть Його.
JOHN|6|65|І сказав Він: Я тому й говорив вам, що до Мене прибути не може ніхто, як не буде йому від Отця дане те.
JOHN|6|66|Із того часу відпали багато-хто з учнів Його, і не ходили вже з Ним.
JOHN|6|67|І сказав Ісус Дванадцятьом: Чи не хочете й ви відійти?
JOHN|6|68|Відповів Йому Симон Петро: До кого ми підемо, Господи? Ти маєш слова життя вічного.
JOHN|6|69|Ми ж увірували та пізнали, що Ти Христос, Син Бога Живого!
JOHN|6|70|Відповів їм Ісус: Чи не Дванадцятьох Я вас вибрав? Та один із вас диявол...
JOHN|6|71|Це сказав Він про Юду, сина Симонового, Іскаріота. Бо цей мав Його видати, хоч він був один із Дванадцятьох.
JOHN|7|1|Після цього Ісус ходив по Галілеї, не хотів бо ходити по Юдеї, бо юдеї шукали нагоди, щоб убити Його.
JOHN|7|2|А надходило свято юдейське Кучки.
JOHN|7|3|І сказали до Нього брати Його: Піди звідси, і йди до Юдеї, щоб і учні Твої побачили вчинки Твої, що Ти робиш.
JOHN|7|4|Тайкома бо не робить нічого ніхто, але сам прагне бути відомий. Коли Ти таке чиниш, то з'яви Себе світові.
JOHN|7|5|Бо не вірували в Нього навіть брати Його!
JOHN|7|6|А Ісус промовляє до них: Не настав ще Мій час, але завжди готовий час ваш.
JOHN|7|7|Вас ненавидіти світ не може, а Мене він ненавидить, бо Я свідчу про нього, що діла його злі.
JOHN|7|8|Ідіть на це свято, Я ж іще не піду на це свято, бо не виповнився ще Мій час.
JOHN|7|9|Це сказавши до них, Він зоставсь у Галілеї.
JOHN|7|10|Коли ж вийшли на свято брати Його, тоді й Сам Він пішов, не відкрито, але ніби потай.
JOHN|7|11|А юдеї за свята шукали Його та питали: Де Він?
JOHN|7|12|І поголоска велика про Нього в народі була. Одні говорили: Він добрий, а інші казали: Ні, Він зводить з дороги народ...
JOHN|7|13|Та відкрито про Нього ніхто не казав, бо боялись юдеїв.
JOHN|7|14|У половині вже свята Ісус у храм увійшов і навчав.
JOHN|7|15|І дивувались юдеї й казали: Як Він знає Писання, не вчившись?
JOHN|7|16|Відповів їм Ісус і сказав: Наука Моя не Моя, а Того, Хто послав Мене.
JOHN|7|17|Коли хоче хто волю чинити Його, той довідається про науку, чи від Бога вона, чи від Себе Самого кажу Я.
JOHN|7|18|Хто говорить від себе самого, той власної слави шукає, а Хто слави шукає Того, Хто послав Його, Той правдивий, і в Ньому неправди нема.
JOHN|7|19|Чи ж Закона вам дав не Мойсей? Та ніхто з вас Закона того не виконує. Нащо хочете вбити Мене?
JOHN|7|20|Народ відповів: Чи Ти демона маєш? Хто Тебе хоче вбити?
JOHN|7|21|Ісус відповів і сказав їм: Одне діло зробив Я, і всі ви дивуєтесь.
JOHN|7|22|Через це Мойсей дав обрізання вам, не тому, що воно від Мойсея, але від отців, та ви й у суботу обрізуєте чоловіка.
JOHN|7|23|Коли ж чоловік у суботу приймає обрізання, щоб Закону Мойсеєвого не порушити, чого ж ремствуєте ви на Мене, що Я всю людину в суботу вздоровив?
JOHN|7|24|Не судіть за обличчям, але суд справедливий чиніть!
JOHN|7|25|Дехто ж з єрусалимлян казали: Хіба це не Той, що Його шукають убити?
JOHN|7|26|Бо говорить відкрито ось Він, і нічого не кажуть Йому. Чи то справді дізналися старші, що Він дійсно Христос?
JOHN|7|27|Та ми знаєм Цього, звідки Він. Про Христа ж, коли прийде, ніхто знати не буде, звідки Він.
JOHN|7|28|І скликнув у храмі Ісус, навчаючи й кажучи: І Мене знаєте ви, і знаєте, звідки Я. А Я не прийшов Сам від Себе; правдивий же Той, Хто послав Мене, що Його ви не знаєте.
JOHN|7|29|Я знаю Його, Я бо від Нього, і послав Мене Він!
JOHN|7|30|Тож шукали вони, щоб схопити Його, та ніхто не наклав рук на Нього, бо то ще не настала година Його.
JOHN|7|31|А багато з народу в Нього ввірували та казали: Коли прийде Христос, чи ж Він чуда чинитиме більші, як чинить Оцей?
JOHN|7|32|Фарисеї прочули такі поголоски про Нього в народі. Тоді первосвященики та фарисеї послали свою службу, щоб схопити Його.
JOHN|7|33|Ісус же сказав: Ще недовго побуду Я з вами, та й до Того піду, Хто послав Мене.
JOHN|7|34|Ви будете шукати Мене, і не знайдете; а туди, де Я є, ви прибути не можете...
JOHN|7|35|Тоді говорили юдеї між собою: Куди це Він хоче йти, що не знайдемо Його? Чи не хоче йти до виселенців між греки, та й греків навчати?
JOHN|7|36|Що за слово, яке Він сказав: Ви будете шукати Мене, і не знайдете; а туди, де Я є, ви прибути не можете?
JOHN|7|37|А останнього великого дня свята Ісус стояв і кликав, говорячи: Коли прагне хто з вас нехай прийде до Мене та й п'є!
JOHN|7|38|Хто вірує в Мене, як каже Писання, то ріки живої води потечуть із утроби його.
JOHN|7|39|Це ж сказав Він про Духа, що мали прийняти Його, хто ввірував у Нього. Не було бо ще Духа на них, не був бо Ісус ще прославлений.
JOHN|7|40|А багато з народу, почувши слова ті, казали: Він справді пророк!
JOHN|7|41|Інші казали: Він Христос. А ще інші казали: Хіба прийде Христос із Галілеї?
JOHN|7|42|Чи ж не каже Писання, що Христос прийде з роду Давидового, і з села Віфлеєму, звідкіля був Давид?
JOHN|7|43|Так повстала незгода в народі з-за Нього.
JOHN|7|44|А декотрі з них мали замір схопити Його, та ніхто не поклав рук на Нього.
JOHN|7|45|І вернулася служба до первосвящеників та фарисеїв, а ті їх запитали: Чому не привели ви Його?
JOHN|7|46|Відказала та служба: Чоловік ще ніколи так не промовляв, як Оцей Чоловік...
JOHN|7|47|А їм відповіли фарисеї: Чи й вас із дороги не зведено?
JOHN|7|48|Хіба хто з старших або з фарисеїв увірував у Нього?
JOHN|7|49|Та проклятий народ, що не знає Закону!
JOHN|7|50|Говорить до них Никодим, що приходив до Нього вночі, і що був один із них:
JOHN|7|51|Хіба судить Закон наш людину, як перше її не вислухає, і не дізнається, що вона робить?
JOHN|7|52|Йому відповіли та сказали вони: Чи й ти не з Галілеї? Досліди та побач, що не прийде Пророк із Галілеї.
JOHN|7|53|І до дому свого пішов кожен.
JOHN|8|1|Ісус же на гору Оливну пішов.
JOHN|8|2|А над ранком прийшов знов у храм, і всі люди збігались до Нього. А Він сів і навчав їх.
JOHN|8|3|І ось книжники та фарисеї приводять до Нього в перелюбі схоплену жінку, і посередині ставлять її,
JOHN|8|4|та й говорять Йому: Оцю жінку, Учителю, зловлено на гарячому вчинку перелюбу...
JOHN|8|5|Мойсей же в Законі звелів нам таких побивати камінням. А Ти що говориш?
JOHN|8|6|Це ж казали вони, Його спокушуючи, та щоб мати на Нього оскарження. А Ісус, нахилившись додолу, по землі писав пальцем...
JOHN|8|7|А коли ті не переставали питати Його, Він підвівся й промовив до них: Хто з вас без гріха, нехай перший на неї той каменем кине!...
JOHN|8|8|І Він знов нахилився додолу, і писав по землі...
JOHN|8|9|А вони, це почувши й сумлінням докорені, стали один по одному виходити, почавши з найстарших та аж до останніх. І зоставсь Сам Ісус і та жінка, що стояла всередині...
JOHN|8|10|І підвівся Ісус, і нікого, крім жінки, не бачивши, промовив до неї: Де ж ті, жінко, що тебе оскаржали? Чи ніхто тебе не засудив?
JOHN|8|11|А вона відказала: Ніхто, Господи... І сказав їй Ісус: Не засуджую й Я тебе. Іди собі, але більш не гріши!
JOHN|8|12|І знову Ісус промовляв до них, кажучи: Я Світло для світу. Хто йде вслід за Мною, не буде ходити у темряві той, але матиме світло життя.
JOHN|8|13|Фарисеї ж Йому відказали: Ти Сам свідчиш про Себе, тим свідоцтво Твоє неправдиве.
JOHN|8|14|Відповів і сказав їм Ісус: Хоч і свідчу про Себе Я Сам, та правдиве свідоцтво Моє, бо Я знаю, звідкіля Я прийшов і куди Я йду. Ви ж не відаєте, відкіля Я приходжу, і куди Я йду.
JOHN|8|15|Ви за тілом судите, Я не суджу нікого.
JOHN|8|16|А коли Я суджу, то правдивий Мій суд, бо не Сам Я, а Я та Отець, що послав Він Мене!
JOHN|8|17|Та й у вашім Законі написано, що свідчення двох чоловіків правдиве.
JOHN|8|18|Я Сам свідчу про Себе Самого, і свідчить про Мене Отець, що послав Він Мене.
JOHN|8|19|І сказали до Нього вони: Де Отець Твій? Ісус відповів: Не знаєте ви ні Мене, ні Мого Отця. Якби знали Мене, то й Отця Мого знали б.
JOHN|8|20|Ці слова Він казав при скарбниці, у храмі навчаючи. І ніхто не схопив Його, бо то ще не настала година Його...
JOHN|8|21|І сказав Він їм знову: Я відходжу, ви ж шукати Мене будете, і помрете в гріху своїм. Куди Я йду, туди ви прибути не можете...
JOHN|8|22|А юдеї казали: Чи не вб'є Він Сам Себе, коли каже: Куди Я йду, туди ви прибути не можете?
JOHN|8|23|І сказав Він до них: Ви від долу, Я звисока, і ви зо світу цього, Я не з цього світу.
JOHN|8|24|Тому Я сказав вам, що помрете в своїх гріхах. Бо коли не ввіруєте, що то Я, то помрете в своїх гріхах.
JOHN|8|25|А вони запитали Його: Хто Ти такий? І Ісус відказав їм: Той, Хто спочатку, як і говорю Я до вас.
JOHN|8|26|Я маю багато про вас говорити й судити; правдивий же Той, Хто послав Мене, і Я світові те говорю, що від Нього почув.
JOHN|8|27|Але не зрозуміли вони, що то Він про Отця говорив їм.
JOHN|8|28|Тож Ісус їм сказав: Коли ви підіймете Людського Сина, тоді зрозумієте, що то Я, і що Сам Я від Себе нічого не дію, але те говорю, як Отець Мій Мене був навчив.
JOHN|8|29|А Той, Хто послав Мене, перебуває зо Мною; Отець не зоставив Самого Мене, бо Я завжди чиню, що Йому до вподоби.
JOHN|8|30|Коли Він говорив це, то багато-хто в Нього увірували.
JOHN|8|31|Тож промовив Ісус до юдеїв, що в Нього ввірували: Як у слові Моїм позостанетеся, тоді справді Моїми учнями будете,
JOHN|8|32|і пізнаєте правду, а правда вас вільними зробить!
JOHN|8|33|Вони відказали Йому: Авраамів ми рід, і нічиїми невільниками не були ми ніколи. То як же Ти кажеш: Ви станете вільні?
JOHN|8|34|Відповів їм Ісус: Поправді, поправді кажу вам, що кожен, хто чинить гріх, той раб гріха.
JOHN|8|35|І не зостається раб у домі повік, але Син зостається повік.
JOHN|8|36|Коли Син отже зробить вас вільними, то справді ви будете вільні.
JOHN|8|37|Знаю Я, що ви рід Авраамів, але хочете смерть заподіяти Мені, бо наука Моя не вміщається в вас.
JOHN|8|38|Я те говорю, що Я бачив в Отця, та й ви робите те, що ви бачили в батька свого.
JOHN|8|39|Сказали вони Йому в відповідь: Наш отець Авраам. Відказав їм Ісус: Коли б ви Авраамові діти були, то чинили б діла Авраамові.
JOHN|8|40|А тепер ось ви хочете вбити Мене, Чоловіка, що вам казав правду, яку чув Я від Бога. Цього Авраам не робив.
JOHN|8|41|Ви робите діла батька свого. Вони ж відказали Йому: Не родилися ми від перелюбу, одного ми маєм Отця то Бога.
JOHN|8|42|А Ісус їм сказав: Якби Бог був Отець ваш, ви б любили Мене, бо від Бога Я вийшов і прийшов, не від Себе ж Самого прийшов Я, а Мене Він послав.
JOHN|8|43|Чому мови Моєї ви не розумієте? Бо не можете чути ви слова Мого.
JOHN|8|44|Ваш батько диявол, і пожадливості батька свого ви виконувати хочете. Він був душогуб споконвіку, і в правді не встояв, бо правди нема в нім. Як говорить неправду, то говорить зо свого, бо він неправдомовець і батько неправді.
JOHN|8|45|А Мені ви не вірите, бо Я правду кажу.
JOHN|8|46|Хто з вас може Мені докорити за гріх? Коли ж правду кажу, чом Мені ви не вірите?
JOHN|8|47|Хто від Бога, той слухає Божі слова; через те ви не слухаєте, що ви не від Бога.
JOHN|8|48|Відізвались юдеї й сказали Йому: Чи ж не добре ми кажемо, що Ти самарянин і демона маєш?
JOHN|8|49|Ісус відповів: Не маю Я демона, та шаную Свого Отця, ви ж Мене зневажаєте.
JOHN|8|50|Не шукаю ж Я власної слави, є Такий, Хто шукає та судить.
JOHN|8|51|Поправді, поправді кажу вам: Хто слово Моє берегтиме, не побачить той смерти повік!
JOHN|8|52|І сказали до Нього юдеї: Тепер ми дізнались, що демона маєш: умер Авраам і пророки, а Ти кажеш: Хто науку Мою берегтиме, не скуштує той смерти повік.
JOHN|8|53|Чи ж Ти більший, аніж отець наш Авраам, що помер? Та повмирали й пророки. Ким Ти робиш Самого Себе?
JOHN|8|54|Ісус відповів: Як Я славлю Самого Себе, то ніщо Моя слава. Мене прославляє Отець Мій, про Якого ви кажете, що Він Бог ваш.
JOHN|8|55|І ви не пізнали Його, а Я знаю Його. А коли Я скажу, що не знаю Його, буду неправдомовець, подібний до вас. Та Я знаю Його, і слово Його зберігаю.
JOHN|8|56|Отець ваш Авраам прагнув із радістю, щоб побачити день Мій, і він бачив, і тішився.
JOHN|8|57|А юдеї ж до Нього сказали: Ти й п'ятидесяти років не маєш іще, і Авраама Ти бачив?
JOHN|8|58|Ісус їм відказав: Поправді, поправді кажу вам: Перш, ніж був Авраам, Я є.
JOHN|8|59|І схопили каміння вони, щоб кинути на Нього. Та сховався Ісус, і з храму пішов.
JOHN|9|1|А коли Він проходив, побачив чоловіка, що сліпим був з народження.
JOHN|9|2|І спитали Його учні Його, говорячи: Учителю, хто згрішив: чи він сам, чи батьки його, що сліпим він родився?
JOHN|9|3|Ісус відповів: Не згрішив ані він, ні батьки його, а щоб діла Божі з'явились на ньому.
JOHN|9|4|Ми мусимо виконувати діла Того, Хто послав Мене, аж поки є день. Надходить он ніч, коли жаден нічого не зможе виконувати.
JOHN|9|5|Доки Я в світі, Я Світло для світу.
JOHN|9|6|Промовивши це, Він сплюнув на землю, і з слини грязиво зробив, і очі сліпому помазав грязивом,
JOHN|9|7|і до нього промовив: Піди, умийся в ставку Сілоам визначає це Посланий. Тож пішов той і вмився, і вернувся видющим...
JOHN|9|8|А сусіди та ті, що бачили перше його, як був він сліпий, говорили: Чи ж не той це, що сидів та просив?
JOHN|9|9|Говорили одні, що це він, а інші казали: Ні, подібний до нього. А він відказав: Це я!
JOHN|9|10|І питали його: Як же очі відкрились тобі?
JOHN|9|11|А той оповідав: Чоловік, що Його звуть Ісусом, грязиво зробив, і очі помазав мені, і до мене сказав: Піди в Сілоам та й умийся. Я ж пішов та й умився, і став бачити.
JOHN|9|12|І сказали до нього: Де Він? Відказує той: Я не знаю.
JOHN|9|13|Ведуть тоді до фарисеїв того, що був перше незрячий.
JOHN|9|14|А була то субота, як грязиво Ісус учинив і відкрив йому очі.
JOHN|9|15|І знов запитали його й фарисеї, як видющим він став. А він розповів їм: Грязиво поклав Він на очі мені, а я вмився, та й бачу.
JOHN|9|16|Тоді деякі з фарисеїв казали: Не від Бога Оцей Чоловік, бо суботи не держить. А інші казали: Як же чуда такі може грішна людина чинити? І незгода між ними була.
JOHN|9|17|Тому знову говорять сліпому: Що ти кажеш про Нього, коли очі відкрив Він тобі? А той відказав: Він Пророк!
JOHN|9|18|Юдеї проте йому не повірили, що незрячим він був і прозрів, аж поки не покликано батьків того прозрілого.
JOHN|9|19|І запитали їх, кажучи: Чи ваш оце син, про якого ви кажете, ніби родився сліпим? Як же він тепер бачить?
JOHN|9|20|А батьки його відповіли та сказали: Ми знаєм, що цей то наш син, і що він народився сліпим.
JOHN|9|21|Але як тепер бачить, не знаємо, або хто йому очі відкрив, ми не відаємо. Поспитайте його, він дорослий, хай сам скаже про себе...
JOHN|9|22|Таке говорили батьки його, бо боялись юдеїв: юдеї бо вже були змовились, як хто за Христа Його визнає, щоб той був відлучений від синагоги.
JOHN|9|23|Ось тому говорили батьки його: Він дорослий, його поспитайте.
JOHN|9|24|І покликали вдруге того чоловіка, що був сліпим, і сказали йому: Віддай хвалу Богові. Ми знаємо, що грішний Отой Чоловік.
JOHN|9|25|Але він відповів: Чи Він грішний не знаю. Одне тільки знаю, що я був сліпим, а тепер бачу!...
JOHN|9|26|І спитали його: Що тобі Він зробив? Як відкрив тобі очі?
JOHN|9|27|Відповів він до них: Я вже вам говорив, та не слухали ви. Що бажаєте знову почути? Може й ви Його учнями хочете стати?
JOHN|9|28|А вони його вилаяли та й сказали: То ти Його учень, а ми учні Мойсеєві.
JOHN|9|29|Ми знаємо, що Бог говорив до Мойсея, звідки ж узявся Оцей, ми не відаємо.
JOHN|9|30|Відповів чоловік і сказав їм: То ж воно й дивно, що не знаєте ви, звідки Він, а Він мені очі відкрив!
JOHN|9|31|Та ми знаємо, що грішників Бог не послухає; хто ж богобійний, і виконує волю Його, того слухає Він.
JOHN|9|32|Відвіку не чувано, щоб хто очі відкрив був сліпому з народження.
JOHN|9|33|Коли б не від Бога був Цей, Він нічого не міг би чинити.
JOHN|9|34|Вони відповіли та й сказали йому: Ти ввесь у гріхах народився, і чи тобі нас учити? І геть його вигнали.
JOHN|9|35|Дізнався Ісус, що вони того вигнали геть, і, знайшовши його, запитав: Чи віруєш ти в Сина Божого?
JOHN|9|36|Відповів той, говорячи: Хто ж то, Пане, Такий, щоб я вірував у Нього?
JOHN|9|37|Промовив до нього Ісус: І ти бачив Його, і Той, Хто говорить з тобою то Він!...
JOHN|9|38|А він відказав: Я вірую, Господи! І вклонився Йому.
JOHN|9|39|І промовив Ісус: На суд Я прийшов у цей світ, щоб бачили темні, а видющі щоб стали незрячі.
JOHN|9|40|І почули це деякі з тих фарисеїв, що були з Ним, та й сказали Йому: Чи ж і ми невидющі?
JOHN|9|41|Відказав їм Ісус: Якби ви невидющі були, то не мали б гріха; а тепер ви говорите: Бачимо, то й ваш гріх зостається при вас!
JOHN|10|1|Поправді, поправді кажу вам: Хто не входить дверима в кошару, але перелазить деінде, той злодій і розбійник.
JOHN|10|2|А хто входить дверима, той вівцям пастух.
JOHN|10|3|Воротар відчиняє йому, і його голосу слухають вівці; і свої вівці він кличе по йменню, і випроваджує їх.
JOHN|10|4|А як вижене всі свої вівці, він іде перед ними, і вівці слідом за ним ідуть, бо знають голос його.
JOHN|10|5|За чужим же не підуть вони, а будуть утікати від нього, бо не знають вони чужого голосу.
JOHN|10|6|Оцю притчу повів їм Ісус, але не зрозуміли вони, про що їм говорив.
JOHN|10|7|І знову промовив Ісус: Поправді, поправді кажу вам, що Я двері вівцям.
JOHN|10|8|Усі, скільки їх перше Мене приходило, то злодії й розбійники, але вівці не слухали їх.
JOHN|10|9|Я двері: коли через Мене хто ввійде, спасеться, і той ввійде та вийде, і пасовисько знайде.
JOHN|10|10|Злодій тільки на те закрадається, щоб красти й убивати та нищити. Я прийшов, щоб ви мали життя, і подостатком щоб мали.
JOHN|10|11|Я Пастир Добрий! Пастир добрий кладе життя власне за вівці.
JOHN|10|12|А наймит, і той, хто не вівчар, кому вівці не свої, коли бачить, що вовк наближається, то кидає вівці й тікає, а вовк їх хапає й полошить.
JOHN|10|13|А наймит утікає тому, що він наймит, і не дбає про вівці.
JOHN|10|14|Я Пастир Добрий, і знаю Своїх, і Свої Мене знають.
JOHN|10|15|Як Отець Мене знає, так і Я Отця знаю, і власне життя Я за вівці кладу.
JOHN|10|16|Також маю Я інших овець, які не з цієї кошари, Я повинен і їх припровадити. І Мій голос почують вони, і буде отара одна й Один Пастир!
JOHN|10|17|Через те Отець любить Мене, що Я власне життя віддаю, щоб ізнову прийняти його.
JOHN|10|18|Ніхто в Мене його не бере, але Я Сам від Себе кладу його. Маю владу віддати його, і маю владу прийняти його знову, Я цю заповідь взяв від Свого Отця.
JOHN|10|19|З-за цих слів між юдеями знову незгода знялася.
JOHN|10|20|І багато-хто з них говорили: Він демона має, і несамовитий. Чого слухаєте ви Його?
JOHN|10|21|Інші казали: Ці слова не того, хто демона має. Хіба демон може очі сліпим відкривати?...
JOHN|10|22|Було тоді свято Відновлення в Єрусалимі. Стояла зима.
JOHN|10|23|А Ісус у храмі ходив, у Соломоновім ґанку.
JOHN|10|24|Юдеї тоді обступили Його та й казали Йому: Доки будеш тримати в непевності нас? Якщо Ти Христос, то відкрито скажи нам!
JOHN|10|25|Відповів їм Ісус: Я вам був сказав, та не вірите ви. Ті діла, що чиню їх у Ймення Свого Отця, вони свідчать про Мене.
JOHN|10|26|Та не вірите ви, не з Моїх бо овець ви.
JOHN|10|27|Мого голосу слухають вівці Мої, і знаю Я їх, і за Мною слідком вони йдуть.
JOHN|10|28|І Я життя вічне даю їм, і вони не загинуть повік, і ніхто їх не вихопить із Моєї руки.
JOHN|10|29|Мій Отець, що дав їх Мені, Він більший за всіх, і вихопити ніхто їх не може Отцеві з руки.
JOHN|10|30|Я й Отець Ми одне!
JOHN|10|31|Знов каміння схопили юдеї, щоб укаменувати Його.
JOHN|10|32|Відповів їм Ісус: Від Отця показав Я вам добрих учинків багато, за котрий же з тих учинків хочете Мене каменувати?
JOHN|10|33|Юдеї Йому відказали: Не за добрий учинок хочемо Тебе вкаменувати, а за богозневагу, бо Ти, бувши людиною, за Бога Себе видаєш...
JOHN|10|34|Відповів їм Ісус: Хіба не написано в вашім Законі: Я сказав: ви боги?
JOHN|10|35|Коли тих Він богами назвав, що до них слово Боже було, а Писання не може порушене бути,
JOHN|10|36|то Тому, що Отець освятив і послав Його в світ, закидаєте ви: Зневажаєш Ти Бога, через те, що сказав Я: Я Син Божий?
JOHN|10|37|Коли Я не чиню діл Свого Отця, то не вірте Мені.
JOHN|10|38|А коли Я чиню, то хоч ви Мені віри й не ймете, повірте ділам, щоб пізнали й повірили ви, що Отець у Мені, а Я ув Отці!
JOHN|10|39|Тоді знову шукали вони, щоб схопити Його, але вийшов із рук їхніх Він.
JOHN|10|40|І Він знову на той бік Йордану пішов, на те місце, де Іван найперше христив, та й там перебував.
JOHN|10|41|І багато до Нього приходили та говорили, що хоч жадного чуда Іван не вчинив, але все, що про Нього Іван говорив, правдиве було.
JOHN|10|42|І багато-хто ввірували в Нього там.
JOHN|11|1|Був же хворий один, Лазар у Віфанії, із села Марії й сестри її Марти.
JOHN|11|2|А Марія, що брат її Лазар був хворий, була та, що помазала Господа миром, і волоссям своїм Йому ноги обтерла.
JOHN|11|3|Тоді сестри послали до Нього, говорячи: Ось нездужає, Господи, той, що кохаєш його!...
JOHN|11|4|Як почув же Ісус, то промовив: Не на смерть ця недуга, а на Божу славу, щоб Син Божий прославився нею.
JOHN|11|5|А Ісус любив Марту, і сестру її, і Лазаря.
JOHN|11|6|А коли Він почув, що нездужає той, то зостався два дні на тім місці, де був.
JOHN|11|7|Після ж того говорить до учнів: Ходімо знову в Юдею.
JOHN|11|8|Йому учні сказали: Учителю, таж допіру юдеї хотіли камінням побити Тебе, а Ти знов туди підеш?
JOHN|11|9|Ісус відповів: Хіба дня не дванадцять годин? Як хто ходить за дня, не спіткнеться, цьогосвітнє бо світло він бачить.
JOHN|11|10|А хто ходить нічної пори, той спіткнеться, бо немає в нім світла.
JOHN|11|11|Оце Він сказав, а по тому говорить до них: Друг наш Лазар заснув, та піду розбудити Його.
JOHN|11|12|А учні сказали Йому: Як заснув, то він, Господи, видужає.
JOHN|11|13|Та про смерть його мовив Ісус, вони ж думали, що про сонний спочинок Він каже.
JOHN|11|14|Тоді просто сказав їм Ісус: Умер Лазар.
JOHN|11|15|І Я тішусь за вас, що там Я не був, щоб повірили ви. Та ходімо до нього.
JOHN|11|16|Сказав же Хома, називаний Близнюк, до співучнів: Ходімо й ми, щоб із Ним повмирати.
JOHN|11|17|Як прибув же Ісус, то знайшов, що чотири вже дні той у гробі.
JOHN|11|18|А Віфанія поблизу Єрусалиму була, яких стадій з п'ятнадцять.
JOHN|11|19|І багато з юдеїв до Марти й Марії прийшли, щоб за брата розважити їх.
JOHN|11|20|Тоді Марта, почувши, що надходить Ісус, побігла зустріти Його, Марія ж удома сиділа.
JOHN|11|21|І Марта сказала Ісусові: Коли б, Господи, був Ти отут, то не вмер би мій брат...
JOHN|11|22|Та й тепер, знаю я, що чого тільки в Бога попросиш, то дасть Тобі Бог!
JOHN|11|23|Промовляє до неї Ісус: Воскресне твій брат!
JOHN|11|24|Відказує Марта Йому: Знаю, що в воскресення останнього дня він воскресне.
JOHN|11|25|Промовив до неї Ісус: Я воскресення й життя. Хто вірує в Мене, хоч і вмре, буде жити.
JOHN|11|26|І кожен, хто живе та хто вірує в Мене, повіки не вмре. Чи ти віруєш в це?
JOHN|11|27|Вона каже Йому: Так, Господи! Я вірую, що Ти Христос, Син Божий, що має прийти на цей світ.
JOHN|11|28|І промовивши це, відійшла, та й покликала нишком Марію, сестру свою, кажучи: Учитель тут, і Він кличе тебе!
JOHN|11|29|А та, як зачула, квапливо встала й до Нього пішла.
JOHN|11|30|А Ісус не ввійшов був іще до села, а знаходивсь на місці, де Марта зустріла Його.
JOHN|11|31|Юдеї тоді, що були з нею в домі й її розважали, як побачили, що Марія квапливо встала й побігла, подалися за нею, гадаючи, що до гробу пішла вона, плакати там.
JOHN|11|32|Як Марія ж прийшла туди, де був Ісус, і Його вгледіла, то припала до ніг Йому та й говорила до Нього: Коли б, Господи, був Ти отут, то не вмер би мій брат!
JOHN|11|33|А Ісус, як побачив, що плаче вона, і плачуть юдеї, що з нею прийшли, то в дусі розжалобився та й зворушився Сам,
JOHN|11|34|і сказав: Де його ви поклали? Говорять Йому: Іди, Господи, та подивися!
JOHN|11|35|І закапали сльози Ісусові...
JOHN|11|36|А юдеї казали: Дивись, як кохав Він його!
JOHN|11|37|А з них дехто сказали: Чи не міг же зробити Отой, Хто очі сліпому відкрив, щоб і цей не помер?
JOHN|11|38|Ісус же розжалобивсь знову в Собі, і до гробу прийшов. Була ж то печера, і камінь на ній налягав.
JOHN|11|39|Промовляє Ісус: Відваліть цього каменя! Сестра вмерлого Марта говорить до Нього: Уже, Господи, чути, бо чотири вже дні він у гробі...
JOHN|11|40|Ісус каже до неї: Чи тобі не казав Я, що як будеш ти вірувати, славу Божу побачиш?
JOHN|11|41|І зняли тоді каменя. А Ісус ізвів очі до неба й промовив: Отче, дяку приношу Тобі, що Мене Ти почув.
JOHN|11|42|Та Я знаю, що Ти завжди почуєш Мене, але ради народу, що довкола стоїть, Я сказав, щоб увірували, що послав Ти Мене.
JOHN|11|43|І, промовивши це, Він скричав гучним голосом: Лазарю, вийди сюди!
JOHN|11|44|І вийшов померлий, по руках і ногах обв'язаний пасами, а обличчя у нього було перев'язане хусткою... Ісус каже до них: Розв'яжіть його та й пустіть, щоб ходив...
JOHN|11|45|І багато з юдеїв, що посходилися до Марії, та бачили те, що Він учинив, у Нього ввірували.
JOHN|11|46|А деякі з них пішли до фарисеїв, і їм розповіли, що Ісус учинив.
JOHN|11|47|Тоді первосвященики та фарисеї скликали раду й казали: Що маємо робити, бо Цей Чоловік пребагато чуд чинить?
JOHN|11|48|Якщо так позоставимо Його, то всі в Нього ввірують, і прийдуть римляни, та й візьмуть нам і Край, і народ!
JOHN|11|49|А один із них, Кайяфа, що був первосвящеником року того, промовив до них: Ви нічого не знаєте,
JOHN|11|50|і не поміркуєте, що краще для вас, щоб один чоловік прийняв смерть за людей, аніж щоб увесь народ мав загинути!
JOHN|11|51|А того не сказав сам від себе, але, первосвящеником бувши в тім році, пророкував, що Ісус за народ мав умерти,
JOHN|11|52|і не лише за народ, але й щоб сполучити в одне розпорошених Божих дітей.
JOHN|11|53|Отож, від того дня вони змовилися, щоб убити Його.
JOHN|11|54|І тому не ходив більш Ісус між юдеями явно, але звідти вдавсь до околиць поближче пустині, до міста, що зветься Єфрем, і тут залишався з Своїми учнями.
JOHN|11|55|Наближалася ж Пасха юдейська, і багато-хто з Краю вдались перед Пасхою в Єрусалим, щоб очистити себе.
JOHN|11|56|І шукали Ісуса вони, а в храмі стоявши, гомоніли один до одного: А як вам здається? Хіба Він не прийде на свято?
JOHN|11|57|А первосвященики та фарисеї наказа дали: як дізнається хто, де Він перебуватиме, нехай донесе, щоб схопити Його.
JOHN|12|1|Ісус же за шість день до Пасхи прибув до Віфанії, де жив Лазар, що його воскресив Ісус із мертвих.
JOHN|12|2|І для Нього вечерю там справили, а Марта прислуговувала. Був же й Лазар одним із тих, що до столу з Ним сіли.
JOHN|12|3|А Марія взяла літру мира, з найдорожчого нарду пахучого, і намастила Ісусові ноги, і волоссям своїм Йому ноги обтерла... І пахощі мира наповнили дім!
JOHN|12|4|І говорить один з Його учнів, Юда Іскаріотський, що мав Його видати:
JOHN|12|5|Чому мира оцього за триста динарів не продано, та й не роздано вбогим?
JOHN|12|6|А це він сказав не тому, що про вбогих журився, а тому, що був злодій: він мав скриньку на гроші, і крав те, що вкидали.
JOHN|12|7|І промовив Ісус: Позостав її ти, це вона на день похорону заховала Мені...
JOHN|12|8|Бо вбогих ви маєте завжди з собою, а Мене не постійно ви маєте!
JOHN|12|9|А натовп великий юдеїв довідався, що Він там, та й поприходили не з-за Ісуса Самого, але щоб побачити й Лазаря, що його воскресив Він із мертвих.
JOHN|12|10|А первосвященики змовилися, щоб і Лазареві смерть заподіяти,
JOHN|12|11|бо багато з юдеїв з-за нього відходили, та в Ісуса ввірували.
JOHN|12|12|А другого дня, коли безліч народу, що зібрався на свято, прочула, що до Єрусалиму надходить Ісус,
JOHN|12|13|то взяли вони пальмове віття, і вийшли назустріч Йому та й кричали: Осанна! Благословенний, хто йде у Господнє Ім'я! Цар Ізраїлів!
JOHN|12|14|Ісус же, знайшовши осля, сів на нього, як написано:
JOHN|12|15|Не бійся, дочко Сіонська! Ото Цар твій іде, сидячи на ослі молодому!
JOHN|12|16|А учні Його спочатку того не зрозуміли були, але, як прославивсь Ісус, то згадали тоді, що про Нього було так написано, і що цеє вчинили Йому.
JOHN|12|17|Тоді свідчив народ, який був із Ним, що Він викликав Лазаря з гробу, і воскресив його з мертвих.
JOHN|12|18|Через це й зустрів натовп Його, бо почув, що Він учинив таке чудо.
JOHN|12|19|Фарисеї тоді між собою казали: Ви бачите, що нічого не вдієте: ось пішов увесь світ услід за Ним!
JOHN|12|20|А між тими, що в свято прийшли поклонитись, були й деякі геллени.
JOHN|12|21|І вони підійшли до Пилипа, що з Віфсаїди Галілейської, і просили його та казали: Ми хочемо, пане, побачити Ісуса.
JOHN|12|22|Іде Пилип та Андрієві каже; іде Андрій і Пилип та Ісусові розповідають.
JOHN|12|23|Ісус же їм відповідає, говорячи: Надійшла година, щоб Син Людський прославивсь.
JOHN|12|24|Поправді, поправді кажу вам: коли зерно пшеничне, як у землю впаде, не помре, то одне зостається; як умре ж, плід рясний принесе.
JOHN|12|25|Хто кохає душу свою, той погубить її; хто ж ненавидить душу свою на цім світі, збереже її в вічне життя.
JOHN|12|26|Як хто служить Мені, хай іде той за Мною, і де Я, там буде й слуга Мій. Як хто служить Мені, того пошанує Отець.
JOHN|12|27|Затривожена зараз душа Моя. І що Я повім? Заступи Мене, Отче, від цієї години! Та на те Я й прийшов на годину оцю...
JOHN|12|28|Прослав, Отче, Ім'я Своє! Залунав тоді голос із неба: І прославив, і знову прославлю!
JOHN|12|29|А народ, що стояв і почув, говорив: Загреміло! Інші казали: Це Ангол Йому говорив!
JOHN|12|30|Ісус відповів і сказав: Не для Мене цей голос лунав, а для вас.
JOHN|12|31|Тепер суд цьому світові. Князь світу цього буде вигнаний звідси тепер.
JOHN|12|32|І, як буду піднесений з землі, то до Себе Я всіх притягну.
JOHN|12|33|А Він це говорив, щоб зазначити, якою то смертю Він має померти.
JOHN|12|34|А народ відповів Йому: Ми чули з Закону, що Христос перебуває повік, то чого ж Ти говориш, що Людському Сину потрібно піднесеному бути? Хто такий Цей Син Людський?
JOHN|12|35|І сказав їм Ісус: Короткий ще час світло з вами. Ходіть, поки маєте світло, щоб вас темрява не обгорнула. А хто в темряві ходить, не знає, куди він іде...
JOHN|12|36|Аж доки ви маєте світло, то віруйте в світло, щоб синами світла ви стали. Промовивши це, Ісус відійшов, і сховався від них.
JOHN|12|37|І хоч Він стільки чуд перед ними вчинив був, та в Нього вони не ввірували,
JOHN|12|38|щоб справдилось слово пророка Ісаї, який провіщав: Хто повірив тому, що ми, Господи, чули, а Господнє рамено кому об'явилось?
JOHN|12|39|Тому не могли вони вірити, що знову Ісая прорік:
JOHN|12|40|Засліпив їхні очі, і скам'янив їхнє серце, щоб очима не бачили, ані серцем щоб не зрозуміли, і не навернулись, щоб Я їх уздоровив!
JOHN|12|41|Це Ісая сказав, коли бачив славу Його, і про Нього звіщав.
JOHN|12|42|Проте багато-хто навіть із старших у Нього ввірували, та не признавались через фарисеїв, щоб не вигнано їх із синагоги.
JOHN|12|43|Бо любили вони славу людську більше, аніж славу Божу.
JOHN|12|44|А Ісус підняв голос, та й промовляв: Хто вірує в Мене, не в Мене він вірує, але в Того, Хто послав Мене.
JOHN|12|45|А хто бачить Мене, той бачить Того, хто послав Мене.
JOHN|12|46|Я, Світло, на світ прийшов, щоб кожен, хто вірує в Мене, у темряві не зоставався.
JOHN|12|47|Коли б же хто слів Моїх слухав та не вірував, Я того не суджу, бо Я не прийшов світ судити, але щоб спасти світ.
JOHN|12|48|Хто цурається Мене, і Моїх слів не приймає, той має для себе суддю: те слово, що Я говорив, останнього дня воно буде судити його!
JOHN|12|49|Бо від Себе Я не говорив, а Отець, що послав Мене, то Він Мені заповідь дав, що Я маю казати та що говорити.
JOHN|12|50|І відаю Я, що Його ота заповідь то вічне життя. Тож що Я говорю, то так говорю, як Отець Мені розповідав.
JOHN|13|1|Перед святом же Пасхи Ісус, знавши, що настала година Йому перейти до Отця з цього світу, полюбивши Своїх, що на світі були, до кінця полюбив їх.
JOHN|13|2|Під час же вечері, як диявол уже був укинув у серце синові Симона Юді Іскаріотському, щоб він видав Його,
JOHN|13|3|то Ісус, знавши те, що Отець віддав все Йому в руки, і що від Бога прийшов Він, і до Бога відходить,
JOHN|13|4|устає від вечері, і здіймає одежу, бере рушника й підперізується.
JOHN|13|5|Потому налив Він води до вмивальниці, та й зачав обмивати ноги учням, і витирати рушником, що ним був підперезаний.
JOHN|13|6|І підходить до Симона Петра, а той каже Йому: Ти, Господи, митимеш ноги мені?
JOHN|13|7|Ісус відказав і промовив йому: Що Я роблю, ти не знаєш тепер, але опісля зрозумієш.
JOHN|13|8|Говорить до Нього Петро: Ти повік мені ніг не обмиєш! Ісус відповів йому: Коли Я не вмию тебе, ти не матимеш частки зо Мною.
JOHN|13|9|До Нього проказує Симон Петро: Господи, не самі мої ноги, а й руки та голову!
JOHN|13|10|Ісус каже йому: Хто обмитий, тільки ноги обмити потребує, бо він чистий увесь. І ви чисті, та не всі.
JOHN|13|11|Бо Він знав Свого зрадника, тому то сказав: Ви чисті не всі.
JOHN|13|12|Коли ж пообмивав їхні ноги, і одежу Свою Він надів, засів знову за стіл і промовив до них: Чи знаєте ви, що Я зробив вам?
JOHN|13|13|Ви Мене називаєте: Учитель і Господь, і добре ви кажете, бо Я є.
JOHN|13|14|А коли обмив ноги вам Я, Господь і Вчитель, то повинні й ви один одному ноги вмивати.
JOHN|13|15|Бо то Я вам приклада дав, щоб і ви те чинили, як Я вам учинив.
JOHN|13|16|Поправді, поправді кажу вам: Раб не більший за пана свого, посланець же не більший від того, хто вислав його.
JOHN|13|17|Коли знаєте це, то блаженні ви, якщо таке чините!
JOHN|13|18|Не про всіх вас кажу. Знаю Я, кого вибрав, але щоб збулося Писання: Хто хліб споживає зо Мною, підняв той на Мене п'яту свою!
JOHN|13|19|Уже тепер вам кажу, перше ніж те настане, щоб як станеться, ви ввірували, що то Я.
JOHN|13|20|Поправді, поправді кажу вам: Хто приймає Мого посланця, той приймає Мене; хто ж приймає Мене, той приймає Того, Хто послав Мене!
JOHN|13|21|Промовивши це, затривожився духом Ісус, і освідчив, говорячи: Поправді, поправді кажу вам, що один із вас видасть Мене!...
JOHN|13|22|І озиралися учні один на одного, непевними бувши, про кого Він каже.
JOHN|13|23|При столі, при Ісусовім лоні, був один з Його учнів, якого любив Ісус.
JOHN|13|24|От цьому кивнув Симон Петро та й шепнув: Запитай, хто б то був, що про нього Він каже?
JOHN|13|25|І, пригорнувшись до лоня Ісусового, той говорить до Нього: Хто це, Господи?
JOHN|13|26|Ісус же відказує: Це той, кому, умочивши, подам Я куска. І, вмочивши куска, подав синові Симона, Юді Іскаріотському!...
JOHN|13|27|За тим же куском тоді в нього ввійшов сатана. А Ісус йому каже: Що ти робиш роби швидше...
JOHN|13|28|Але жаден із тих, хто був при столі, того не зрозумів, до чого сказав Він йому.
JOHN|13|29|А тому, що тримав Юда скриньку на гроші, то деякі думали, ніби каже до нього Ісус: Купи, що потрібно на свято для нас, або щоб убогим подав що.
JOHN|13|30|А той, узявши кусок хліба, зараз вийшов. Була ж ніч.
JOHN|13|31|Тоді, як він вийшов, промовляє Ісус: Тепер ось прославивсь Син Людський, і в Ньому прославився Бог.
JOHN|13|32|Коли в Ньому прославився Бог, то і Його Бог прославить у Собі, і зараз прославить Його!
JOHN|13|33|Мої дітоньки, не довго вже бути Мені з вами! Ви шукати Мене будете, але як сказав Я юдеям: Куди Я йду, туди ви прибути не можете, те й вам говорю Я тепер.
JOHN|13|34|Нову заповідь Я вам даю: Любіть один одного! Як Я вас полюбив, так любіть один одного й ви!
JOHN|13|35|По тому пізнають усі, що ви учні Мої, як будете мати любов між собою.
JOHN|13|36|А Симон Петро Йому каже: Куди, Господи, ідеш Ти? Ісус відповів: Куди Я йду, туди ти тепер іти за Мною не можеш, але потім ти підеш за Мною.
JOHN|13|37|Говорить до Нього Петро: Чому, Господи, іти за Тобою тепер я не можу? За Тебе я душу свою покладу!
JOHN|13|38|Ісус відповідає: За Мене покладеш ти душу свою? Поправді, поправді кажу Я тобі: Півень не заспіває, як ти тричі зречешся Мене...
JOHN|14|1|Нехай серце вам не тривожиться! Віруйте в Бога, і в Мене віруйте!
JOHN|14|2|Багато осель у домі Мого Отця; а коли б то не так, то сказав би Я вам, що йду приготувати місце для вас?
JOHN|14|3|А коли відійду й приготую вам місце, Я знову прийду й заберу вас до Себе, щоб де Я були й ви.
JOHN|14|4|А куди Я йду дорогу ви знаєте.
JOHN|14|5|Говорить до Нього Хома: Ми не знаємо, Господи, куди йдеш; як же можемо знати дорогу?
JOHN|14|6|Промовляє до нього Ісус: Я дорога, і правда, і життя. До Отця не приходить ніхто, якщо не через Мене.
JOHN|14|7|Коли б то були ви пізнали Мене, ви пізнали були б і Мого Отця. Відтепер Його знаєте ви, і Його бачили.
JOHN|14|8|Говорить до Нього Пилип: Господи, покажи нам Отця, і вистачить нам!
JOHN|14|9|Промовляє до нього Ісус: Стільки часу Я з вами, ти ж не знаєш, Пилипе, Мене? Хто бачив Мене, той бачив Отця, то як же ти кажеш: Покажи нам Отця?
JOHN|14|10|Чи не віруєш ти, що Я в Отці, а Отець у Мені? Слова, що Я вам говорю, говорю не від Себе, а Отець, що в Мені перебуває, Той чинить діла ті.
JOHN|14|11|Повірте Мені, що Я в Отці, а Отець у Мені! Коли ж ні, то повірте за вчинки самі.
JOHN|14|12|Поправді, поправді кажу вам: Хто вірує в Мене, той учинить діла, які чиню Я, і ще більші від них він учинить, бо Я йду до Отця.
JOHN|14|13|І коли що просити ви будете в Імення Моє, те вчиню, щоб у Сині прославивсь Отець.
JOHN|14|14|Коли будете в Мене просити чого в Моє Ймення, то вчиню.
JOHN|14|15|Якщо Ви Мене любите, Мої заповіді зберігайте!
JOHN|14|16|І вблагаю Отця Я, і Втішителя іншого дасть вам, щоб із вами повік перебував,
JOHN|14|17|Духа правди, що Його світ прийняти не може, бо не бачить Його та не знає Його. Його знаєте ви, бо при вас перебуває, і в вас буде Він.
JOHN|14|18|Я не кину вас сиротами, Я прибуду до вас!
JOHN|14|19|Ще недовго, і вже світ Мене не побачить, але ви Мене бачити будете, бо живу Я і ви жити будете!
JOHN|14|20|Того дня пізнаєте ви, що в Своїм Я Отці, а ви в Мені, і Я в вас.
JOHN|14|21|Хто заповіді Мої має та їх зберігає, той любить Мене. А хто любить Мене, то полюбить його Мій Отець, і Я полюблю Його, і об'явлюсь йому Сам.
JOHN|14|22|Запитує Юда, не Іскаріотський, Його: Що то, Господи, що Ти нам об'явитися маєш, а не світові?
JOHN|14|23|Ісус відповів і до нього сказав: Як хто любить Мене, той слово Моє берегтиме, і Отець Мій полюбить його, і Ми прийдемо до нього, і оселю закладемо в нього.
JOHN|14|24|Хто не любить Мене, той не береже Моїх слів. А слово, що чуєте ви, не Моє, а Отця, що послав Мене.
JOHN|14|25|Говорив це Я вам, бувши з вами.
JOHN|14|26|Утішитель же, Дух Святий, що Його Отець пошле в Ім'я Моє, Той навчить вас усього, і пригадає вам усе, що Я вам говорив.
JOHN|14|27|Зоставляю вам мир, мир Свій вам даю! Я даю вам не так, як дає світ. Серце ваше нехай не тривожиться, ані не лякається!
JOHN|14|28|Чули ви, що Я вам говорив: Я відходжу, і вернуся до вас. Якби ви любили Мене, то ви б тішилися, що Я йду до Отця, бо більший за Мене Отець.
JOHN|14|29|І тепер Я сказав вам, передніше, ніж сталося, щоб ви вірували, коли станеться.
JOHN|14|30|Небагато вже Я говоритиму з вами, бо надходить князь світу цього, а в Мені він нічого не має,
JOHN|14|31|та щоб світ зрозумів, що люблю Я Отця, і як Отець наказав Мені, так роблю. Уставайте, ходім звідсіля!
JOHN|15|1|Я правдива Виноградина, а Отець Мій Виноградар.
JOHN|15|2|Усяку галузку в Мене, що плоду не приносить, Він відтинає, але всяку, що плід родить, обчищає її, щоб рясніше родила.
JOHN|15|3|Через Слово, що Я вам говорив, ви вже чисті.
JOHN|15|4|Перебувайте в Мені, а Я в вас! Як та вітка не може вродити плоду сама з себе, коли не позостанеться на виноградині, так і ви, як в Мені перебувати не будете.
JOHN|15|5|Я Виноградина, ви галуззя! Хто в Мені перебуває, а Я в ньому, той рясно зароджує, бо без Мене нічого чинити не можете ви.
JOHN|15|6|Коли хто перебувати не буде в Мені, той буде відкинений геть, як галузка, і всохне. І громадять їх, і кладуть на огонь, і згорять.
JOHN|15|7|Коли ж у Мені перебувати ви будете, а слова Мої позостануться в вас, то просіть, чого хочете, і станеться вам!
JOHN|15|8|Отець Мій прославиться в тому, якщо рясно зародите й будете учні Мої.
JOHN|15|9|Як Отець полюбив Мене, так і Я полюбив вас. Перебувайте в любові Моїй!
JOHN|15|10|Якщо будете ви зберігати Мої заповіді, то в любові Моїй перебуватимете, як і Я зберіг Заповіді Свого Отця, і перебуваю в любові Його.
JOHN|15|11|Це Я вам говорив, щоб радість Моя була в вас, і щоб повна була ваша радість!
JOHN|15|12|Оце Моя заповідь, щоб любили один одного ви, як Я вас полюбив!
JOHN|15|13|Ніхто більшої любови не має над ту, як хто свою душу поклав би за друзів своїх.
JOHN|15|14|Ви друзі Мої, якщо чините все, що Я вам заповідую.
JOHN|15|15|Я вже більше не буду рабами вас звати, бо не відає раб, що пан його чинить. А вас назвав друзями Я, бо Я вам об'явив усе те, що почув від Мого Отця.
JOHN|15|16|Не ви Мене вибрали, але Я вибрав вас, і вас настановив, щоб ішли ви й приносили плід, і щоб плід ваш зостався, щоб дав вам Отець, чого тільки попросите в Імення Моє.
JOHN|15|17|Це Я вам заповідую, щоб любили один одного ви!
JOHN|15|18|Коли вас світ ненавидить, знайте, що Мене він зненавидів перше, як вас.
JOHN|15|19|Коли б ви зо світу були, то своє світ любив би. А що ви не зо світу, але Я вас зо світу обрав, тому світ вас ненавидить.
JOHN|15|20|Пригадайте те слово, яке Я вам сказав: Раб не більший за пана свого. Як Мене переслідували, то й вас переслідувати будуть; як слово Моє зберігали, берегтимуть і ваше.
JOHN|15|21|Але все це робитимуть вам за Ім'я Моє, бо не знають Того, хто послав Мене.
JOHN|15|22|Коли б Я не прийшов і до них не казав, то не мали б гріха, а тепер вимовки не мають вони за свій гріх.
JOHN|15|23|Хто Мене ненавидить, і Мого Отця той ненавидить.
JOHN|15|24|Коли б Я серед них не вчинив був тих діл, яких не чинив ніхто інший, то не мали б гріха. Та тепер вони бачили, і зненавиділи і Мене, і Мого Отця.
JOHN|15|25|Та щоб справдилось слово, що в їхнім Законі написане: Мене безпідставно зненавиділи!
JOHN|15|26|А коли Втішитель прибуде, що Його від Отця Я пошлю вам, Той Дух правди, що походить від Отця, Він засвідчить про Мене.
JOHN|15|27|Та засвідчте і ви, бо ви від початку зо Мною.
JOHN|16|1|Оце Я сказав вам, щоб ви не спокусились.
JOHN|16|2|Вас виженуть із синагог. Прийде навіть година, коли кожен, хто вам смерть заподіє, то думатиме, ніби службу приносить він Богові!
JOHN|16|3|А це вам учинять, бо вони не пізнали Отця, ні Мене.
JOHN|16|4|Але Я це сказав вам, щоб згадали про те, про що говорив був Я вам, як настане година. Цього вам не казав Я спочатку, бо з вами Я був.
JOHN|16|5|Тепер же до Того Я йду, Хто послав Мене, і ніхто з вас Мене не питає: Куди йдеш?
JOHN|16|6|Та від того, що це Я сказав вам, серце ваше наповнилось смутком.
JOHN|16|7|Та Я правду кажу вам: Краще для вас, щоб пішов Я, бо як Я не піду, Утішитель не прийде до вас. А коли Я піду, то пошлю вам Його.
JOHN|16|8|А як прийде, Він світові виявить про гріх, і про правду, і про суд:
JOHN|16|9|тож про гріх, що не вірують у Мене;
JOHN|16|10|а про правду, що Я до Отця Свого йду, і Мене не побачите вже;
JOHN|16|11|а про суд, що засуджений князь цього світу.
JOHN|16|12|Я ще маю багато сказати вам, та тепер ви не можете знести.
JOHN|16|13|А коли прийде Він, Той Дух правди, Він вас попровадить до цілої правди, бо не буде казати Сам від Себе, а що тільки почує, казатиме, і що має настати, звістить вам.
JOHN|16|14|Він прославить Мене, бо Він візьме з Мого та й вам сповістить.
JOHN|16|15|Усе, що має Отець, то Моє; через те Я й сказав, що Він візьме з Мого та й вам сповістить.
JOHN|16|16|Незабаром, і Мене вже не будете бачити, і знов незабаром і Мене ви побачите, бо Я йду до Отця.
JOHN|16|17|А деякі з учнів Його говорили один до одного: Що таке, що сказав Він до нас: Незабаром, і Мене вже не будете бачити, і знов незабаром і Мене ви побачите, та: Я йду до Отця?...
JOHN|16|18|Гомоніли також: Що таке, що говорить: Незабаром? Про що каже, не знаємо...
JOHN|16|19|Ісус же пізнав, що хочуть поспитати Його, і сказав їм: Чи про це між собою міркуєте ви, що сказав Я: Незабаром, і вже Мене бачити не будете ви, і знов незабаром і Мене ви побачите?
JOHN|16|20|Поправді, поправді кажу вам, що ви будете плакати та голосити, а світ буде радіти. Сумувати ви будете, але сум ваш обернеться в радість!
JOHN|16|21|Журиться жінка, що родить, бо настала година її. Як дитинку ж породить вона, то вже не пам'ятає терпіння з-за радощів, що людина зродилась на світ...
JOHN|16|22|Так сумуєте й ви ось тепер, та побачу вас знову, і серце ваше радітиме, і ніхто радости вашої вам не відійме!
JOHN|16|23|Ні про що ж того дня ви Мене не спитаєте. Поправді, поправді кажу вам: Чого тільки попросите ви від Отця в Моє Ймення, Він дасть вам.
JOHN|16|24|Не просили ви досі нічого в Ім'я Моє. Просіть і отримаєте, щоб повна була ваша радість.
JOHN|16|25|Оце все Я в притчах до вас говорив. Настає година, коли притчами Я вже не буду до вас промовляти, але явно звіщу про Отця вам.
JOHN|16|26|Того дня ви проситимете в Моє Ймення, і Я вам не кажу, що вблагаю Отця Я за вас,
JOHN|16|27|бо Отець любить Сам вас за те, що ви полюбили Мене та й увірували, що Я вийшов від Бога.
JOHN|16|28|Від Отця вийшов Я, і на світ Я прийшов. І знов покидаю Я світ та й іду до Отця.
JOHN|16|29|Його учні відказують: Ось тепер Ти говориш відкрито, і жадної притчі не кажеш.
JOHN|16|30|Тепер відаємо ми, що Ти знаєш усе, і потреби не маєш, щоб Тебе хто питав. Тому віруємо, що Ти вийшов від Бога!
JOHN|16|31|Ісус їм відповів: Тепер віруєте?
JOHN|16|32|Ото настає година, і вже настала, що ви розпорошитесь кожен у власне своє, а Мене ви Самого покинете... Та не Сам Я, бо зо Мною Отець!
JOHN|16|33|Це Я вам розповів, щоб мали ви мир у Мені. Страждання зазнаєте в світі, але будьте відважні: Я світ переміг!
JOHN|17|1|По мові оцій Ісус очі Свої звів до неба й промовив: Прийшла, Отче, година, прослав Сина Свого, щоб і Син Твій прославив Тебе,
JOHN|17|2|бо Ти дав Йому владу над тілом усяким, щоб Він дав життя вічне всім їм, яких дав Ти Йому.
JOHN|17|3|Життя ж вічне це те, щоб пізнали Тебе, єдиного Бога правдивого, та Ісуса Христа, що послав Ти Його.
JOHN|17|4|Я прославив Тебе на землі, довершив Я те діло, що Ти дав Мені виконати.
JOHN|17|5|І тепер прослав, Отче, Мене Сам у Себе тією славою, яку в Тебе Я мав, поки світ не постав.
JOHN|17|6|Я Ім'я Твоє виявив людям, що Мені Ти із світу їх дав. Твоїми були вони, і Ти дав їх Мені, і вони зберегли Твоє слово.
JOHN|17|7|Тепер пізнали вони, що все те, що Ти Мені дав, від Тебе походить,
JOHN|17|8|бо слова, що дав Ти Мені, Я їм передав, і вони прийняли й зрозуміли правдиво, що Я вийшов від Тебе, і ввірували, що послав Ти Мене.
JOHN|17|9|Я благаю за них. Не за світ Я благаю, а за тих, кого дав Ти Мені, Твої бо вони!
JOHN|17|10|Усе бо Моє то Твоє, а Твоє то Моє, і прославивсь Я в них.
JOHN|17|11|І не на світі вже Я, а вони ще на світі, а Я йду до Тебе. Святий Отче, заховай в Ім'я Своє їх, яких дав Ти Мені, щоб як Ми, єдине були!
JOHN|17|12|Коли з ними на світі Я був, Я беріг їх у Ймення Твоє, тих, що дав Ти Мені, і зберіг, і ніхто з них не згинув, крім призначеного на загибіль, щоб збулося Писання.
JOHN|17|13|Тепер же до Тебе Я йду, але це говорю Я на світі, щоб мали вони в собі радість Мою досконалу.
JOHN|17|14|Я їм дав Твоє слово, але світ їх зненавидів, бо вони не від світу, як і Я не від світу.
JOHN|17|15|Не благаю, щоб Ти їх зо світу забрав, але щоб зберіг їх від злого.
JOHN|17|16|Не від світу вони, як і Я не від світу.
JOHN|17|17|Освяти Ти їх правдою! Твоє слово то правда.
JOHN|17|18|Як на світ Ти послав Мене, так і Я на світ послав їх.
JOHN|17|19|А за них Я посвячую в жертву Самого Себе, щоб освячені правдою стали й вони.
JOHN|17|20|Та не тільки за них Я благаю, а й за тих, що ради їхнього слова ввірують у Мене,
JOHN|17|21|щоб були всі одно: як Ти, Отче, в Мені, а Я у Тобі, щоб одно були в Нас і вони, щоб увірував світ, що Мене Ти послав.
JOHN|17|22|А ту славу, що дав Ти Мені, Я їм передав, щоб єдине були, як єдине і Ми.
JOHN|17|23|Я у них, а Ти у Мені, щоб були досконалі в одно, і щоб пізнав світ, що послав Мене Ти, і що їх полюбив Ти, як Мене полюбив.
JOHN|17|24|Бажаю Я, Отче, щоб і ті, кого дав Ти Мені, там зо Мною були, де знаходжуся Я, щоб бачили славу Мою, яку дав Ти Мені, бо Ти полюбив Мене перше закладин світу.
JOHN|17|25|Отче Праведний! Хоча не пізнав Тебе світ, та пізнав Тебе Я. І пізнали вони, що послав Мене Ти.
JOHN|17|26|Я ж Ім'я Твоє їм об'явив й об'являтиму, щоб любов, що Ти нею Мене полюбив, була в них, а Я в них!...
JOHN|18|1|Промовивши це, Ісус вийшов із учнями Своїми на той бік потоку Кедрону, де був сад, до якого ввійшов Він та учні Його.
JOHN|18|2|Але й Юда, що видав Його, знав те місце, бо там часто збирались Ісус й Його учні.
JOHN|18|3|Отож Юда, узявши відділ війська та службу від первосвящеників і фарисеїв, приходить туди із смолоскипами, та з ліхтарями, та з зброєю.
JOHN|18|4|А Ісус, усе відавши, що з Ним статися має, виходить та й каже до них: Кого ви шукаєте?
JOHN|18|5|Йому відповіли: Ісуса Назарянина. Він говорить до них: Це Я... А стояв із ними й Юда, що видав Його.
JOHN|18|6|І як тільки сказав їм: Це Я, вони подалися назад, та й на землю попадали...
JOHN|18|7|І Він знов запитав їх: Кого ви шукаєте? Вони ж відказали: Ісуса Назарянина.
JOHN|18|8|Ісус відповів: Я сказав вам, що це Я... Отож, як Мене ви шукаєте, то дайте оцим відійти,
JOHN|18|9|щоб збулося те слово, що Він був сказав: Я не втратив нікого із тих, кого дав Ти Мені.
JOHN|18|10|Тоді Симон Петро, меча мавши, його вихопив, і рубонув раба первосвященика, і відтяв праве вухо йому. А рабу на ім'я було Малх.
JOHN|18|11|Та промовив Ісус до Петра: Всунь у піхви меча! Чи ж не мав би Я пити ту чашу, що Отець дав Мені?
JOHN|18|12|Відділ же війська та тисяцький і служба юдейська схопили Ісуса, і зв'язали Його,
JOHN|18|13|і повели Його перше до Анни, бо тестем доводивсь Кайяфі, що первосвящеником був того року.
JOHN|18|14|Це ж був той Кайяфа, що порадив юдеям, що ліпше померти людині одній за народ.
JOHN|18|15|А Симон Петро й інший учень ішли за Ісусом слідом. Той же учень відомий був первосвященикові, і ввійшов у двір первосвящеників із Ісусом.
JOHN|18|16|А Петро за ворітьми стояв. Тоді вийшов той учень, що відомий був первосвященикові, і сказав воротарці, і впровадив Петра.
JOHN|18|17|І питає Петра воротарка служниця: Ти хіба не з учнів Цього Чоловіка? Той відказує: Ні!
JOHN|18|18|А раби й служба, розклавши огонь, стояли та й грілися, бо був холод. І Петро стояв із ними та грівся.
JOHN|18|19|А первосвященик спитався Ісуса про учнів Його, і про науку Його.
JOHN|18|20|Ісус Йому відповідь дав: Я світові явно казав. Я постійно навчав у синагозі й у храмі, куди всі юдеї збираються, а таємно нічого Я не говорив.
JOHN|18|21|Чого ти питаєш Мене? Поспитайся тих, що чули, що Я їм говорив. Отже, знають вони, про що Я говорив.
JOHN|18|22|А як Він це сказав, то один із присутньої там служби вдарив Ісуса в щоку, говорячи: То так відповідаєш первосвященикові?
JOHN|18|23|Ісус йому відповідь дав: Якщо зле Я сказав, покажи, що то зле; коли ж добре, за що Мене б'єш?
JOHN|18|24|І відіслав Його Анна зв'язаним первосвященикові Кайяфі.
JOHN|18|25|А Симон Петро стояв, гріючись. І сказали до нього: Чи й ти не з учнів Його? Він відрікся й сказав: Ні!
JOHN|18|26|Говорить один із рабів первосвященика, родич тому, що йому Петро вухо відтяв: Чи тебе я не бачив у саду з Ним?
JOHN|18|27|І знову відрікся Петро, і заспівав півень хвилі тієї...
JOHN|18|28|А Ісуса ведуть від Кайяфи в преторій. Був же ранок. Та вони не ввійшли до преторія, щоб не опоганитись, а щоб їсти пасху.
JOHN|18|29|Тоді вийшов Пилат назовні до них і сказав: Яку скаргу приносите ви на Цього Чоловіка?
JOHN|18|30|Вони відповіли та й сказали йому: Коли б Цей злочинцем не був, ми б Його тобі не видавали.
JOHN|18|31|А Пилат їм сказав: Візьміть Його, та й за вашим Законом судіть Його. Юдеї сказали йому: Нам не вільно нікого вбивати,
JOHN|18|32|щоб збулося Ісусове слово, що його Він прорік, зазначаючи, якою то смертю Він має померти.
JOHN|18|33|Тоді знову Пилат увійшов у преторій, і покликав Ісуса, і до Нього сказав: Чи Ти Цар Юдейський?
JOHN|18|34|Ісус відповів: Чи від себе самого питаєш ти це, чи то інші тобі говорили про Мене?
JOHN|18|35|Пилат відповів: Чи ж юдеянин я? Твій народ та первосвященики мені Тебе видали. Що таке Ти вчинив?
JOHN|18|36|Ісус відповів: Моє Царство не із світу цього. Якби із цього світу було Моє Царство, то служба Моя воювала б, щоб не виданий був Я юдеям. Та тепер Моє Царство не звідси...
JOHN|18|37|Сказав же до Нього Пилат: Так Ти Цар? Ісус відповів: Сам ти кажеш, що Цар Я. Я на те народився, і на те прийшов у світ, щоб засвідчити правду. І кожен, хто з правди, той чує Мій голос.
JOHN|18|38|Говорить до Нього Пилат: Що є правда? І сказавши оце, до юдеїв знов вийшов, та й каже до них: Не знаходжу Я в Ньому провини ніякої.
JOHN|18|39|Та ви маєте звичай, щоб я випустив вам одного на Пасху. Чи хочете отже, відпущу вам Царя Юдейського?
JOHN|18|40|Та знову вони зняли крик, вимагаючи: Не Його, а Варавву! А Варавва був злочинець.
JOHN|19|1|От тоді взяв Ісуса Пилат, та й звелів збичувати Його.
JOHN|19|2|Вояки ж, сплівши з терну вінка, Йому поклали на голову, та багряницю наділи на Нього,
JOHN|19|3|і приступали до Нього й казали: Радій, Царю Юдейський! І били по щоках Його...
JOHN|19|4|Тоді вийшов назовні ізнову Пилат та й говорить до них: Ось Його я виводжу назовні до вас, щоб ви переконались, що провини ніякої в Нім не знаходжу.
JOHN|19|5|І вийшов назовні Ісус, у терновім вінку та в багрянім плащі. А Пилат до них каже: Оце Чоловік!
JOHN|19|6|Як зобачили ж Його первосвященики й служба, то закричали, говорячи: Розіпни, розіпни! Пилат каже до них: То візьміть Його ви й розіпніть, бо провини я в Нім не знаходжу!
JOHN|19|7|Відказали юдеї йому: Ми маємо Закона, а за Законом Він мусить умерти, бо за Божого Сина Себе видавав!
JOHN|19|8|Як зачув же Пилат оце слово, налякався ще більш,
JOHN|19|9|і вернувся в преторій ізнову, і питає Ісуса: Звідки Ти? Та Ісус йому відповіді не подав.
JOHN|19|10|І каже до Нього Пилат: Не говориш до мене? Хіба ж Ти не знаєш, що маю я владу розп'ясти Тебе, і маю владу Тебе відпустити?
JOHN|19|11|Ісус відповів: Надо Мною ти жадної влади не мав би, коли б тобі зверху не дано було; тому більший гріх має той, хто Мене тобі видав...
JOHN|19|12|Після цього Пилат намагався пустити Його, та юдеї кричали, говорячи: Якщо Його пустиш, то не кесарів приятель ти! Усякий, хто себе за царя видає, противиться кесареві.
JOHN|19|13|Як зачув же Пилат оце слово, то вивів назовні Ісуса, і засів на суддеве сидіння, на місці, що зветься літостротон, по-гебрейському ж гаввата.
JOHN|19|14|Був то ж день Приготовлення Пасхи, година була близько шостої. І він каже юдеям: Ось ваш Цар!
JOHN|19|15|Та вони закричали: Геть, геть із Ним! Розіпни Його! Пилат каже до них: Царя вашого маю розп'ясти? Первосвященики відповіли: Ми не маєм царя, окрім кесаря!
JOHN|19|16|Ось тоді він їм видав Його, щоб розп'ясти... І взяли Ісуса й повели...
JOHN|19|17|І, нісши Свого хреста, Він вийшов на місце, Череповищем зване, по-гебрейському Голгофа.
JOHN|19|18|Там Його розп'яли, а з Ним разом двох інших, з одного та з другого боку, а Ісуса всередині.
JOHN|19|19|А Пилат написав і написа, та й умістив на хресті. Було ж там написано: Ісус Назарянин, Цар Юдейський.
JOHN|19|20|І багато з юдеїв читали цього написа, бо те місце, де Ісус був розп'ятий, було близько від міста. А було по-гебрейському, по-грецькому й по-римському написано.
JOHN|19|21|Тож сказали Пилатові юдейські первосвященики: Не пиши: Цар Юдейський, але що Він Сам говорив: Я Цар Юдейський.
JOHN|19|22|Пилат відповів: Що я написав написав!
JOHN|19|23|Розп'явши ж Ісуса, вояки взяли одіж Його, та й поділили на чотири частині, по частині для кожного вояка, теж і хітона. А хітон був не шитий, а витканий цілий відверху.
JOHN|19|24|Тож сказали один до одного: Не будемо дерти його, але жереба киньмо на нього, кому припаде. Щоб збулося Писання: Поділили одежу Мою між собою, і метнули про шату Мою жеребка. Вояки ж це й зробили...
JOHN|19|25|Під хрестом же Ісуса стояли Його мати, і сестра Його матері, Марія Клеопова, і Марія Магдалина.
JOHN|19|26|Як побачив Ісус матір та учня, що стояв тут, якого любив, то каже до матері: Оце, жоно, твій син!
JOHN|19|27|Потім каже до учня: Оце мати твоя! І з тієї години той учень узяв її до себе.
JOHN|19|28|Потім, знавши Ісус, що вже все довершилось, щоб збулося Писання, проказує: Прагну!
JOHN|19|29|Тут стояла посудина, повна оцту. Вояки ж, губку оцтом наповнивши, і на тростину її настромивши, піднесли до уст Його.
JOHN|19|30|А коли Ісус оцту прийняв, то промовив: Звершилось!... І, голову схиливши, віддав Свого духа...
JOHN|19|31|Був же день Приготовлення, тож юдеї, щоб тіла на хресті не зосталися в суботу, був бо Великдень тієї суботи просили Пилата зламати голінки розп'ятим, і зняти.
JOHN|19|32|Тож прийшли вояки й поламали голінки першому й другому, що розп'ятий з Ним був.
JOHN|19|33|Коли ж підійшли до Ісуса й побачили, що Він уже вмер, то голінок Йому не зламали,
JOHN|19|34|та один з вояків списом бока Йому проколов, і зараз витекла звідти кров та вода.
JOHN|19|35|І самовидець засвідчив, і правдиве свідоцтво його; і він знає, що правду говорить, щоб повірили й ви.
JOHN|19|36|о це сталось тому, щоб збулося Писання: Йому кості ламати не будуть!
JOHN|19|37|І знов друге Писання говорить: Дивитися будуть на Того, Кого прокололи.
JOHN|19|38|Потім Йосип із Аріматеї, що був учень Ісуса, але потайний, бо боявся юдеїв, став просити Пилата, щоб тіло Ісусове взяти. І дозволив Пилат. Тож прийшов він, і взяв тіло Ісусове.
JOHN|19|39|Прибув також і Никодим, що давніше приходив вночі до Ісуса, і смирну приніс, із алоєм помішану, щось літрів із сто.
JOHN|19|40|Отож, узяли вони тіло Ісусове, та й обгорнули його плащаницею із пахощами, як є звичай ховати в юдеїв.
JOHN|19|41|На тім місці, де Він був розп'ятий, знаходився сад, а в саду новий гріб, що в ньому ніколи ніхто не лежав.
JOHN|19|42|Тож отут, з-за юдейського дня Приготовлення вони поклали Ісуса, бо поблизу був гріб.
JOHN|20|1|А дня першого в тижні, рано вранці, як ще темно було, прийшла Марія Магдалина до гробу, та й бачить, що камінь від гробу відвалений.
JOHN|20|2|Тож біжить вона та й прибуває до Симона Петра, та до другого учня, що Ісус його любив, та й каже до них: Взяли Господа з гробу, і ми не знаємо, де поклали Його!
JOHN|20|3|Тоді вийшов Петро й другий учень, і до гробу пішли.
JOHN|20|4|Вони ж бігли обидва укупі, але другий той учень попереду біг, хутчіш від Петра, і перший до гробу прибув.
JOHN|20|5|І, нахилившися, бачить лежить плащаниця... Але він не ввійшов.
JOHN|20|6|Прибуває і Симон Петро, що слідком за ним біг, і входить до гробу, і плащаницю оглядає, що лежала,
JOHN|20|7|і хустка, що була на Його голові, лежить не з плащаницею, але осторонь, згорнена, в іншому місці...
JOHN|20|8|Тоді ж увійшов й інший учень, що перший до гробу прибув, і побачив, і ввірував.
JOHN|20|9|Бо ще не розуміли з Писання вони, що Він має воскреснути з мертвих.
JOHN|20|10|І учні вернулися знову до себе.
JOHN|20|11|А Марія стояла при гробі назовні та й плакала. Плачучи, нахилилась до гробу.
JOHN|20|12|І бачить два Анголи, що в білім сиділи, один у головах, а другий у ніг, де лежало Ісусове тіло...
JOHN|20|13|І говорять до неї вони: Чого плачеш ти, жінко? Та відказує їм: Узяли мого Господа, і я не знаю, де Його поклали...
JOHN|20|14|І, сказавши оце, обернулась назад, і бачить Ісуса, що стояв, та вона не пізнала, що то Ісус...
JOHN|20|15|Промовляє до неї Ісус: Чого плачеш ти, жінко? Кого ти шукаєш? Вона ж, думаючи, що то садівник, говорить до Нього: Якщо, пане, узяв ти Його, то скажи мені, де поклав ти Його, і Його я візьму!
JOHN|20|16|Ісус мовить до неї: Маріє! А вона обернулася та по-єврейському каже Йому: Раббуні! цебто: Учителю мій!
JOHN|20|17|Говорить до неї Ісус: Не торкайся до Мене, бо Я ще не зійшов до Отця. Але йди до братів Моїх та їм розповіж: Я йду до Свого Отця й Отця вашого, і до Бога Мого й Бога вашого!
JOHN|20|18|Іде Марія Магдалина, та й учням звіщає, що бачила Господа, і Він це їй сказав...
JOHN|20|19|Того ж дня дня першого в тижні, коли вечір настав, а двері, де учні зібрались були, були замкнені, бо боялись юдеїв, з'явився Ісус, і став посередині, та й промовляє до них: Мир вам!
JOHN|20|20|І, сказавши оце, показав Він їм руки та бока. А учні зраділи, побачивши Господа.
JOHN|20|21|Тоді знову сказав їм Ісус: Мир вам! Як Отець послав Мене, і Я вас посилаю!
JOHN|20|22|Сказавши оце, Він дихнув, і говорить до них: Прийміть Духа Святого!
JOHN|20|23|Кому гріхи простите, простяться їм, а кому затримаєте, то затримаються!
JOHN|20|24|А Хома, один з Дванадцятьох, званий Близнюк, із ними не був, як приходив Ісус.
JOHN|20|25|Інші ж учні сказали йому: Ми бачили Господа!... А він відказав їм: Коли на руках Його знаку відцвяшного я не побачу, і пальця свого не вкладу до відцвяшної рани, і своєї руки не вкладу до боку Його, не ввірую!
JOHN|20|26|За вісім же день знов удома були Його учні, а з ними й Хома. І, як замкнені двері були, прийшов Ісус, і став посередині та й проказав: Мир вам!
JOHN|20|27|Потім каже Хомі: Простягни свого пальця сюди, та на руки Мої подивись. Простягни й свою руку, і вклади до боку Мого. І не будь ти невіруючий, але віруючий!
JOHN|20|28|А Хома відповів і сказав Йому: Господь мій і Бог мій!
JOHN|20|29|Промовляє до нього Ісус: Тому ввірував ти, що побачив Мене? Блаженні, що не бачили й увірували!
JOHN|20|30|Багато ж і інших ознак учинив був Ісус у присутності учнів Своїх, що в книзі оцій не записані.
JOHN|20|31|Це ж написано, щоб ви ввірували, що Ісус є Христос, Божий Син, і щоб, віруючи, життя мали в Ім'я Його!
JOHN|21|1|Після цього з'явивсь Ісус знов Своїм учням над морем Тіверіядським. А з'явився отак.
JOHN|21|2|Укупі були Симон Петро, і Хома, званий Близнюк, і Нафанаїл, із Кани Галілейської, і обидва сини Зеведеєві, і двоє інших із учнів Його.
JOHN|21|3|Говорить їм Симон Петро: Піду риби вловити. Вони кажуть до нього: І ми підемо з тобою. І пішли вони, і всіли до човна. Та ночі тієї нічого вони не вловили.
JOHN|21|4|А як ранок настав, то Ісус став над берегом, але учні не знали, що то був Ісус.
JOHN|21|5|Ісус тоді каже до них: Чи не маєте, діти, якоїсь поживи? Ні, вони відказали.
JOHN|21|6|А Він їм сказав: Закиньте невода праворуч від човна, то й знайдете! Вони кинули, і вже не могли його витягнути із-за безлічі риби...
JOHN|21|7|Тоді учень, якого любив був Ісус, говорить Петрові: Це ж Господь!... А Симон Петро, як зачув, що Господь то, накинув на себе одежину, бо він був нагий, та й кинувся в море...
JOHN|21|8|Інші ж учні, що були недалеко від берега якихсь ліктів із двісті припливли човником, тягнучи невода з рибою.
JOHN|21|9|А коли вони вийшли на землю, то бачать розложений жар, а на нім рибу й хліб.
JOHN|21|10|Ісус каже до них: Принесіть тієї риби, що оце ви вловили!
JOHN|21|11|Пішов Симон Петро та й на землю витягнув невода, повного риби великої, сто п'ятдесят три. І хоч стільки було її, не продерся проте невід.
JOHN|21|12|Ісус каже до учнів: Ідіть, снідайте! А з учнів ніхто не наважився спитати Його: Хто Ти такий? Бо знали вони, що Господь то...
JOHN|21|13|Тож підходить Ісус, бере хліб і дає їм, так само ж і рибу.
JOHN|21|14|Це вже втретє з'явився Ісус Своїм учням, як із мертвих воскрес.
JOHN|21|15|Як вони вже поснідали, то Ісус промовляє до Симона Петра: Симоне, сину Йонин, чи ти любиш мене більше цих? Той каже Йому: Так, Господи, відаєш Ти, що кохаю Тебе! Промовляє йому: Паси ягнята Мої!
JOHN|21|16|І говорить йому Він удруге: Симоне, сину Йонин, чи ти любиш Мене? Той каже Йому: Так, Господи, відаєш Ти, що кохаю Тебе! Промовляє йому: Паси вівці Мої!
JOHN|21|17|Утретє Він каже йому: Симоне, сину Йонин, чи кохаєш Мене? Засмутився Петро, що спитав його втретє: Чи кохаєш Мене? І він каже Йому: Ти все відаєш, Господи, відаєш Ти, що кохаю Тебе! Промовляє до нього Ісус: Паси вівці Мої!
JOHN|21|18|Поправді, поправді кажу Я тобі: Коли був ти молодший, то ти сам підперізувався, і ходив, куди ти бажав. А коли постарієш, свої руки простягнеш, і інший тебе підпереже, і поведе, куди не захочеш...
JOHN|21|19|А оце Він сказав, щоб зазначити, якою то смертю той Бога прославить. Сказавши таке, Він говорить йому: Іди за Мною!
JOHN|21|20|Обернувся Петро, та й ось бачить, що за ним слідкома йде той учень, якого любив Ісус, який на вечері до лоня Йому був схилився й спитав: Хто, Господи, видасть Тебе?
JOHN|21|21|Петро, як побачив того, говорить Ісусові: Господи, цей же що?
JOHN|21|22|Промовляє до нього Ісус: Якщо Я схотів, щоб він позостався, аж поки прийду, що до того тобі? Ти йди за Мною!
JOHN|21|23|І це слово рознеслось було між братами, що той учень не вмре. Проте Ісус не сказав йому, що не вмре, а: Якщо Я схотів, щоб він позостався, аж поки прийду, що до того тобі?
JOHN|21|24|Це той учень, що свідчить про це, що й оце написав. І знаємо ми, що правдиве свідоцтво його!
JOHN|21|25|Багато є й іншого, що Ісус учинив. Але думаю, що коли б написати про все те зокрема про кожне, то й сам світ не вмістив би написаних книг! Амінь.
