EZRA|1|1|In anno primo Cyri regis Persarum, ut compleretur verbum Domini ex ore Ieremiae, suscitavit Dominus spiritum Cyri regis Persarum, qui emisit edictum in omni regno suo etiam per scripturam dicens:
EZRA|1|2|" Haec dicit Cyrus rex Persarum: Omnia regna terrae dedit mihi Dominus, Deus caeli, et ipse praecepit mihi, ut aedificarem ei domum in Ierusalem, quae est in Iudaea.
EZRA|1|3|Quis ex vobis est de omni populo eius? Sit Dominus Deus suus cum eo, et ascendat in Ierusalem, quae est in Iudaea, et aedificet domum Domini, Dei Israel; ipse est Deus, qui est in Ierusalem.
EZRA|1|4|Et omnes reliqui in cunctis locis, ubicumque habitant, adiuventur a viris de loco suo, argento et auro et substantia et pecore sicut et oblationibus spontaneis pro templo Dei, quod est in Ierusalem ".
EZRA|1|5|Et surrexerunt principes familiarum de Iuda et Beniamin et sacerdotes et Levitae et omnis, cuius Deus suscitavit spiritum, ut ascenderent ad aedificandum templum Domini, quod erat in Ierusalem.
EZRA|1|6|Universique, qui erant in circuitu, confortaverunt manus eorum cum vasis argenteis et aureis, substantia, pecore et pensitationibus, praeter oblationes spontaneas.
EZRA|1|7|Rex quoque Cyrus protulit vasa templi Domini, quae tulerat Nabuchodonosor de Ierusalem et posuerat ea in templo dei sui;
EZRA|1|8|protulit autem ea Cyrus rex Persarum per manum Mithridatis praepositi thesauri, qui enumeravit ea Sasabassar principi Iudae.
EZRA|1|9|Et hic est numerus eorum: phialae aureae triginta, phialae argenteae mille, cultri viginti novem, scyphi aurei triginta,
EZRA|1|10|scyphi quoque argentei quadringenti decem, vasa alia plurima; 11 omnia vasa aurea et argentea quinque milia quadringenta. Universa tulit Sasabassar cum his, qui ascendebant de transmigratione Babylonis in Ierusalem.
EZRA|2|1|Hi sunt autem provinciae filii, qui ascenderunt de captivitate migrantium, quos transtulerat Nabuchodonosor rex Babylonis in Babylonem, et reversi sunt in Ierusalem et Iudam, unusquisque in civitatem suam.
EZRA|2|2|Qui venerunt cum Zorobabel, Iesua, Nehemias, Saraia, Rahelaia, Mardochaeus, Belsan, Mesphar, Beguai, Rehum, Baana.Numerus virorum populi Israel:
EZRA|2|3|filii Pharos duo milia centum septuaginta duo;
EZRA|2|4|filii Saphatia trecenti septuaginta duo;
EZRA|2|5|filii Area septingenti septuaginta quinque;
EZRA|2|6|filii Phahathmoab, hi sunt filii Iesua et Ioab, duo milia octingenti duodecim;
EZRA|2|7|filii Elam mille ducenti quinquaginta quattuor;
EZRA|2|8|filii Zethua nongenti quadraginta quinque;
EZRA|2|9|filii Zachai septingenti sexaginta;
EZRA|2|10|filii Bani sescenti quadraginta duo;
EZRA|2|11|filii Bebai sescenti viginti tres;
EZRA|2|12|filii Azgad mille ducenti viginti duo;
EZRA|2|13|filii Adonicam sescenti sexaginta sex;
EZRA|2|14|filii Beguai duo milia quinquaginta sex;
EZRA|2|15|filii Adin quadringenti quinquaginta quattuor;
EZRA|2|16|filii Ater, qui erant ex Ezechia, nonaginta octo;
EZRA|2|17|filii Besai trecenti viginti tres;
EZRA|2|18|filii Iora centum duodecim;
EZRA|2|19|filii Hasum ducenti viginti tres;
EZRA|2|20|filii Gebbar nonaginta quinque;
EZRA|2|21|filii Bethlehem centum viginti tres;
EZRA|2|22|viri Netopha quinquaginta sex;
EZRA|2|23|viri Anathoth centum viginti octo;
EZRA|2|24|filii Azmaveth quadraginta duo;
EZRA|2|25|filii Cariathiarim, Cephira et Beroth septingenti quadraginta tres;
EZRA|2|26|filii Rama et Gabaa sescenti viginti unus;
EZRA|2|27|viri Machmas centum viginti duo;
EZRA|2|28|viri Bethel et Hai ducenti viginti tres;
EZRA|2|29|filii Nabo quinquaginta duo;
EZRA|2|30|filii Megbis centum quinquaginta sex;
EZRA|2|31|filii Elam alterius mille ducenti quinquaginta quattuor;
EZRA|2|32|filii Harim trecenti viginti;
EZRA|2|33|filii Lod, Hadid et Ono septingenti viginti quinque;
EZRA|2|34|filii Iericho trecenti quadraginta quinque;
EZRA|2|35|filii Senaa tria milia sescenti triginta.
EZRA|2|36|Sacerdotes: filii Iedaia de domo Iesua nongenti septuaginta tres,
EZRA|2|37|filii Emmer mille quinquaginta duo,
EZRA|2|38|filii Phassur mille ducenti quadraginta septem,
EZRA|2|39|filii Harim mille decem et septem.
EZRA|2|40|Levitae: filii Iesua, hi sunt filii Cadmihel, Bennui, Odoviae, septuaginta quattuor.
EZRA|2|41|Cantores: filii Asaph centum viginti octo.
EZRA|2|42|Ianitores: filii Sellum, filii Ater, filii Telmon, filii Accub, filii Hatita, filii Sobai: universi centum triginta novem.
EZRA|2|43|Oblati: filii Siha, filii Hasupha, filii Tabbaoth,
EZRA|2|44|filii Ceros, filii Siaa, filii Phadon,
EZRA|2|45|filii Lebana, filii Hagaba, filii Accub,
EZRA|2|46|filii Hagab, filii Semlai, filii Hanan,
EZRA|2|47|filii Giddel, filii Gaher, filii Raaia,
EZRA|2|48|filii Rasin, filii Necoda, filii Gazam,
EZRA|2|49|filii Oza, filii Phasea, filii Besai,
EZRA|2|50|filii Asena, filii Meunitarum, filii Nephusorum,
EZRA|2|51|filii Bacbuc, filii Hacupha, filii Harhur,
EZRA|2|52|filii Basluth, filii Mahida, filii Harsa,
EZRA|2|53|filii Bercos, filii Sisara, filii Thema,
EZRA|2|54|filii Nasia, filii Hatipha.
EZRA|2|55|Filii servorum Salomonis: filii Sotai, filii Sophereth, filii Pheruda,
EZRA|2|56|filii Iaala, filii Darcon, filii Giddel,
EZRA|2|57|filii Saphatia, filii Hatil, filii Phochereth Hassebaim, filii Ami.
EZRA|2|58|Omnes oblati et filii servorum Salomonis trecenti nonaginta duo.
EZRA|2|59|Et hi, qui ascenderunt de Thelmela, Thelharsa, Cherub et Addon et Emmer et non potuerunt indicare domum patrum suorum et semen suum, utrum ex Israel essent:
EZRA|2|60|filii Dalaia, filii Tobia, filii Necoda, sescenti quinquaginta duo.
EZRA|2|61|Et de filiis sacerdotum: filii Hobia, filii Accos, filii Berzellai, qui accepit de filiabus Berzellai Galaaditis uxorem et vocatus est nomine eorum.
EZRA|2|62|Hi quaesierunt tabulas genealogiae suae et non invenerunt; et eiecti sunt de sacerdotio.
EZRA|2|63|Et dixit praepositus eis, ut non comederent de sanctificatis sanctuarii, donec surgeret sacerdos pro Urim et Tummim.
EZRA|2|64|Omnis multitudo simul quadraginta duo milia trecenti sexaginta,
EZRA|2|65|exceptis servis eorum et ancillis, qui erant septem milia trecenti triginta septem, insuper et cantores atque cantatrices ducenti.
EZRA|2|66|Equi eorum septingenti triginta sex, muli eorum ducenti quadraginta quinque,
EZRA|2|67|cameli eorum quadringenti triginta quinque, asini eorum sex milia septingenti viginti.
EZRA|2|68|Nonnulli autem de principibus familiarum, cum ingrederentur templum domini, quod est in Ierusalem, sponte obtulerunt in domum Dei ad exstruendam eam in loco suo.
EZRA|2|69|Se cundum vires suas dederunt in aerarium operis auri solidos sexaginta milia et mille, argenti minas quinque milia et vestes sacerdotales centum.
EZRA|2|70|Habitaverunt ergo ibi sacerdotes et Levitae et quidam de populo; cantores autem et ianitores et oblati in urbibus suis, universusque Israel in civitatibus suis.
EZRA|3|1|Iamque venerat mensis septi mus, et erant filii Israel in civita tibus suis. Congregatus est ergo populus quasi vir unus in Ierusalem.
EZRA|3|2|Et surrexit Iesua filius Iosedec et fratres eius sacerdotes et Zorobabel filius Salathiel et fratres eius et aedificaverunt altare Dei Israel, ut offerrent in eo holocautomata, sicut scriptum est in lege Moysi viri Dei.
EZRA|3|3|Collocaverunt autem altare super bases suas, deterrentibus eos per circuitum populis terrarum, et obtulerunt super illud holocaustum Domino mane et vespere.
EZRA|3|4|Feceruntque sollemnitatem Tabernaculorum, sicut scriptum est, et holocaustum diebus singulis per ordinem, secundum praeceptum pro singulis diebus;
EZRA|3|5|et praeter holocaustum sempiternum illa etiam pro calendis et universis sollemnitatibus, quae erant consecratae Domino, et pro omnibus, quae ultro offerebantur Domino.
EZRA|3|6|A primo die mensis septimi coeperunt offerre holocaustum Domino; porro templum Dei nondum fundatum erat.
EZRA|3|7|Dederunt autem pecunias latomis et fabris, cibum quoque et potum et oleum Sidoniis Tyriisque, ut deferrent ligna cedrina de Libano ad mare Ioppe, iuxta quod concesserat Cyrus rex Persarum eis.
EZRA|3|8|Anno autem secundo adventus eorum ad templum Dei in Ierusalem mense secundo, coeperunt Zorobabel filius Salathiel et Iesua filius Iosedec et reliqui de fratribus eorum sacerdotes et Levitae et omnes, qui venerant de captivitate in Ierusalem, et constituerunt Levitas a viginti annis et supra, ut dirigerent opus templi Domini.
EZRA|3|9|Stetitque Iesua et filii eius et fratres eius, Cadmihel, Bennui et Odovia quasi vir unus, ut dirigerent eos, qui faciebant opus in templo Dei; itemque filii Henadad et filii eorum et fratres eorum Levitae.
EZRA|3|10|Fundato igitur ab aedificatoribus templo Domini, steterunt sacerdotes in ornatu suo cum tubis, et Levitae filii Asaph in cymbalis, ut laudarent Deum iuxta mandatum David regis Israel.
EZRA|3|11|Et concinebant in hymnis et gratiarum actione Domino: " Quoniam bonus, quoniam in aeternum misericordia eius " super Israel. Omnis quoque populus vociferabatur clamore magno in laudando Dominum, eo quod fundatum esset templum Domini.
EZRA|3|12|Plurimi etiam senes de sacerdotibus et Levitis et principibus familiarum, qui viderant oculis suis prius templum in loco suo, flebant voce magna; et multi vociferantes in laetitia elevabant vocem.
EZRA|3|13|Nec poterat quisquam agnoscere vocem clamoris laetantium et vocem fletus populi, quoniam populus vociferabatur clamore magno, et strepitus audiebatur procul.
EZRA|4|1|Audierunt autem hostes Iudae et Beniamin, quia filii captivita tis aedificarent templum Domino, Deo Israel,
EZRA|4|2|et accedentes ad Zorobabel et ad principes familiarum dixerunt eis: " Aedificemus vobiscum, quia ita ut vos quaerimus Deum vestrum et immolavimus victimas a diebus Asarhaddon regis Assyriae, qui adduxit nos huc ".
EZRA|4|3|Et dixit eis Zorobabel et Iesua et reliqui principes familiarum Israel: Non est vobis et nobis, ut aedificemus domum Deo nostro, sed nos ipsi soli aedificabimus Domino, Deo Israel, sicut praecepit nobis Cyrus rex Persarum ".
EZRA|4|4|Factum est igitur, ut populus terrae impediret manus populi Iudae et turbaret eos in aedificando.
EZRA|4|5|Conduxerunt autem adversus eos consiliatores, ut destruerent consilium eorum omnibus diebus Cyri regis Persarum et usque ad regnum Darii regis Persarum.
EZRA|4|6|In regno autem Asueri, in principio regni eius, scripserunt accusationem adversus habitatores Iudae et Ierusalem.
EZRA|4|7|Et in diebus Artaxerxis scripsit Beselam, Mithridates et Tabel et reliqui, qui erant in consilio eorum, ad Artaxerxem regem Persarum; scriptura autem accusationis erat scripta litteris Syriacis et composita sermone Syro.
EZRA|4|8|Rehum praefectus et Samsai scriba scripserunt epistulam unam de Ierusalem Artaxerxi regi huiuscemodi:
EZRA|4|9|" Rehum praefectus et Samsai scriba et reliqui socii eorum, iudices et duces, magistratus Persae, Erchuaei, Babylonii, Susanechaei, hoc est Elamitae,
EZRA|4|10|et ceteri de gentibus, quas transtulit Asenaphar magnus et gloriosus et habitare fecit in civitatibus Samariae et in reliquis regionibus trans flumen in pace ".
EZRA|4|11|Hoc est exemplar epistulae, quam miserunt ad eum: Artaxerxi regi, servi tui, viri, qui sunt trans fluvium. Igitur
EZRA|4|12|notum sit regi quia Iudaei, qui ascenderunt a te ad nos, venerunt in Ierusalem civitatem rebellem et pessimam, quam aedificant, exstruentes muros eius, fundamenta iam componentes.
EZRA|4|13|Nunc notum sit regi quia, si civitas illa aedificata fuerit, et muri eius instaurati, tributum et annonam et vectigal non dabunt, et ad ultimum regibus noxa erit.
EZRA|4|14|Nos autem, memores salis, quod in palatio comedimus, et quia laesiones regis videre nefas ducimus, idcirco misimus et nuntiavimus regi,
EZRA|4|15|ut recenseas in libris historiarum patrum tuorum, et invenies in his historiis et scies quoniam urbs illa urbs rebellis est et nocens regibus et provinciis, et seditiones concitantur in ea ex diebus antiquis; quam ob rem et civitas ipsa destructa est.
EZRA|4|16|Nuntiamus nos regi quoniam, si civitas illa aedificata fuerit, et muri ipsius instaurati, possessionem trans fluvium non habebis ".
EZRA|4|17|Verbum misit rex ad Rehum praefectum et Samsai scribam et ad reliquos, qui erant in consilio eorum, qui habitabant in Samaria et in regione trans fluvium: " Pax. Nunc igitur scriptura,
EZRA|4|18|quam misistis ad nos, manifeste lecta est coram me.
EZRA|4|19|Et a me praeceptum est, et recensuerunt inveneruntque quoniam civitas illa a diebus antiquis adversum reges rebellabat, et rebelliones et seditiones concitabantur in ea;
EZRA|4|20|nam et reges fortissimi fuerunt in Ierusalem, qui et dominati sunt omni regioni, quae trans fluvium est, tributum quoque et annonam et vectigal accipiebant.
EZRA|4|21|Nunc ergo praecipite, ut desistant isti homines, et urbs illa non aedificetur, donec forte a me iussum fuerit.
EZRA|4|22|Videte, ne negligenter hoc impleatis, et paulatim crescat malum contra reges ".
EZRA|4|23|Itaque exemplum edicti Artaxerxis regis lectum est coram Rehum praefectum et Samsai scriba et consiliariis eorum; et abierunt festini in Ierusalem ad Iudaeos et prohibuerunt eos in brachio et robore.
EZRA|4|24|Tunc intermissum est opus domus Domini in Ierusalem et non fiebat usque ad annum secundum regni Darii regis Persarum.
EZRA|5|1|Prophetae autem Aggaeus et Zacharias filius Addo propheta verunt ad Iudaeos, qui erant in Iudaea et Ierusalem, in nomine Dei Israel, quod erat super eos.
EZRA|5|2|Tunc surrexerunt Zorobabel filius Salathiel et Iesua filius Iosedec et coeperunt aedificare templum Dei in Ierusalem; prophetae autem Dei adiuvabant eos.
EZRA|5|3|In ipso autem tempore venit ad eos Thathanai, qui erat dux trans flumen, et Stharbuzanai et consiliarii eorum, sicque dixerunt eis: " Quis dedit vobis potestatem, ut domum hanc aedificaretis et materiam istam praepararetis?
EZRA|5|4|Quae sunt nomina hominum auctorum aedificationis illius? ".
EZRA|5|5|Oculus autem Dei eorum factus est super senes Iudaeorum, et non obstiterunt eis, usque dum res ad Darium referretur, et tunc sententia de hac re redderetur.
EZRA|5|6|Exemplar epistulae, quam misit Thathanai dux regionis trans flumen et Stharbuzanai et consiliatores eius et duces, qui erant trans flumen, ad Darium regem.
EZRA|5|7|Sermo, quem miserant ei, sic scriptus erat: Dario regi pax omnis.
EZRA|5|8|Notum sit regi isse nos ad Iudaeam provinciam, ad domum Dei magni, quae aedificatur lapide quadrato, et ligna ponuntur in parietibus; opusque illud diligenter exstruitur et crescit in manibus eorum.
EZRA|5|9|Interrogavimus ergo senes illos et ita diximus eis: "Quis dedit vobis potestatem, ut domum hanc aedificaretis et materiam istam praepararetis?".
EZRA|5|10|Sed et nomina eorum quaesivimus ab eis, ut nuntiaremus tibi, scripsimusque nomina eorum virorum, qui sunt principes in eis.
EZRA|5|11|Huiuscemodi autem sermonem responderunt nobis dicentes: "Nos sumus servi Dei caeli et terrae et aedificamus templum, quod erat exstructum ante hos annos multos, quodque rex Israel magnus aedificaverat et exstruxerat.
EZRA|5|12|Postquam autem ad iracundiam provocaverunt patres nostri Deum caeli, tradidit eos in manus Nabuchodonosor regis Babylonis Chaldaei, qui domum hanc destruxit et populum eius transtulit in Babylonem.
EZRA|5|13|Anno autem primo Cyri regis Babylonis, Cyrus rex proposuit edictum, ut domus Dei haec aedificaretur.
EZRA|5|14|Nam et vasa templi Dei aurea et argentea, quae Nabuchodonosor tulerat de templo, quod erat in Ierusalem, et asportaverat ea in templum Babylonis, protulit Cyrus rex de templo Babylonis, et data sunt viro cuidam nomine Sasabassar, quem et principem constituit,
EZRA|5|15|dixitque ei: 'Haec vasa tolle et vade et pone ea in templo, quod est in Ierusalem, et domus Dei aedificetur in loco suo'.
EZRA|5|16|Tunc itaque Sasabassar ille venit et posuit fundamenta templi Dei in Ierusalem, et ex eo tempore usque nunc aedificatur et necdum completum est".
EZRA|5|17|Nunc ergo, si videtur regi bonum, recenseat in aerario regis, quod est in Babylone, utrumnam a Cyro rege potestas data fuerit, ut aedificaretur domus Dei in Ierusalem, et voluntatem regis super hac re mittat ad nos ".
EZRA|6|1|Tunc Darius rex praecepit, et recensuerunt in tabulis aerarii, quod est in Babylone,
EZRA|6|2|et inventum est in Ecbatanis, quod est castrum in Medena provincia, volumen unum, et sic scriptus erat in eo commentarius:
EZRA|6|3|" Anno primo Cyri regis, Cyrus rex decrevit de domo Dei, quae est in Ierusalem: Aedificetur domus, ubi immolent et sacrificent; altitudo eius cubitorum sexaginta et latitudo eius cubitorum sexaginta,
EZRA|6|4|ordines de lapidibus quadratis tres et ordo de lignis unus; sumptus autem de domo regis dabuntur.
EZRA|6|5|Sed et vasa templi Dei aurea et argentea, quae Nabuchodonosor tulerat de templo Ierusalem et attulerat in Babylonem, reddantur et referantur in templum, quod est in Ierusalem, in locum suum, in templo Dei.
EZRA|6|6|Nunc ergo, Thathanai dux regionis, quae est trans flumen, Stharbuzanai et consiliarii eius et duces, qui estis trans flumen, procul recedite ab illo loco,
EZRA|6|7|dimittite fieri templum Dei illud; dux Iudaeorum et seniores eorum aedificent domum Dei illam in loco suo.
EZRA|6|8|Sed et a me praeceptum est quomodo agere debeatis cum senioribus Iudaeorum illis, qui aedificant domum Dei illam: ut de arca regis, id est de tributis, quae dantur de regione trans flumen, studiose sumptus dentur viris illis sine intermissione.
EZRA|6|9|Et si quid necesse fuerit, sive vituli et arietes et agni in holocaustum Deo caeli, sive frumentum, sal, vinum et oleum, secundum ordinationem sacerdotum, qui sunt in Ierusalem, detur eis per singulos dies sine neglegentia.
EZRA|6|10|Et offerant oblationes suaves Deo caeli orentque pro vita regis et filiorum eius.
EZRA|6|11|A me ergo positum est decretum, ut omnis homo, qui hanc mutaverit iussionem, tollatur lignum de domo ipsius et erigatur et configatur in eo; domus autem eius ponatur in sterquilinium.
EZRA|6|12|Deus autem, qui habitare fecit nomen suum ibi, dissipet omnia regna et populum, qui extenderit manum suam, ut contemnat et dissipet domum Dei illam, quae est in Ierusalem. Ego Darius statui decretum, quod studiose impleri volo ".
EZRA|6|13|Igitur Thathanai dux regionis trans flumen et duces et consiliarii eius, secundum quod praeceperat Darius rex, sic diligenter exsecuti sunt.
EZRA|6|14|Seniores autem Iudaeorum prosperabantur in aedificatione iuxta prophetiam Aggaei prophetae et Zachariae filii Addo et perfecerunt aedificationem, iubente Deo Israel et iubente Cyro et Dario et Artaxerxe regibus Persarum,
EZRA|6|15|et compleverunt domum Dei istam die tertia mensis Adar, qui est annus sextus regni Darii regis.
EZRA|6|16|Fecerunt autem filii Israel, sacerdotes et Levitae et reliqui filiorum transmigrationis dedicationem domus Dei illius in gaudio.
EZRA|6|17|Et obtulerunt in dedicationem domus Dei illius boves centum, arietes ducentos, agnos quadringentos, hircos caprarum pro peccato totius Israel duodecim, iuxta numerum tribuum Israel.
EZRA|6|18|Et statuerunt sacerdotes in ordinibus suis et Levitas in vicibus suis in ministerium Dei in Ierusalem, sicut scriptum est in libro Moysi.
EZRA|6|19|Fecerunt autem filii Israel transmigrationis Pascha quarta decima die mensis primi.
EZRA|6|20|Levitae universi se purificaverunt; purificati autem cuncti immolaverunt Pascha universis filiis transmigrationis et fratribus suis sacerdotibus et sibi.
EZRA|6|21|Et comederunt filii Israel, qui reversi fuerant de transmigratione, et omnes, qui a coinquinatione gentium terrae transierunt ad eos, ut quaererent Dominum, Deum Israel.
EZRA|6|22|Et fecerunt sollemnitatem Azymorum septem diebus in laetitia, quoniam laetificaverat eos Dominus et converterat cor regis Assyriae ad eos, ut adiuvaret manus eorum in opere domus Domini, Dei Israel.
EZRA|7|1|Post haec autem in regno Arta xerxis regis Persarum, Esdras fi lius Saraiae filii Azariae filii Helciae
EZRA|7|2|filii Sellum filii Sadoc filii Achitob
EZRA|7|3|filii Amariae filii Azariae filii Meraioth
EZRA|7|4|filii Zaraiae filii Ozi filii Bocci
EZRA|7|5|filii Abisue filii Phinees filii Eleazar filii Aaron summi sacerdotis,
EZRA|7|6|ipse Esdras ascendit de Babylone et ipse scriba velox in lege Moysi, quam dedit Dominus, Deus Israel. Cumque manus Domini Dei eius esset super eum, dedit ei rex omnem petitionem eius.
EZRA|7|7|Et ascenderunt de filiis Israel et de filiis sacerdotum et de filiis Levitarum et de cantoribus et de ianitoribus et de oblatis in Ierusalem, anno septimo Artaxerxis regis.
EZRA|7|8|Venit in Ierusalem mense quinto, ipse est annus septimus regis.
EZRA|7|9|In primo die mensis primi coepit ascendere de Babylone et in primo die mensis quinti venit in Ierusalem, iuxta manum Dei sui bonam super se.
EZRA|7|10|Esdras enim applicavit cor suum, ut investigaret et impleret legem Domini et faceret et doceret in Israel praeceptum et iudicium.
EZRA|7|11|Hoc est autem exemplar epistulae, quam dedit rex Artaxerxes Esdrae sacerdoti, scribae erudito in mandatis Domini et praeceptis eius in Israel.
EZRA|7|12|" Artaxerxes rex regum Esdrae sacerdoti, scribae legis Dei caeli, salutem.
EZRA|7|13|A me decretum est, ut cuicumque placuerit in regno meo de populo Israel et de sacerdotibus eius et de Levitis ire in Ierusalem, tecum vadat.
EZRA|7|14|A facie enim regis et septem consiliatorum eius missus es, ut visites Iudaeam et Ierusalem secundum legem Dei tui, quae est in manu tua,
EZRA|7|15|et ut feras argentum et aurum, quod rex et consiliatores eius sponte obtulerunt Deo Israel, cuius in Ierusalem tabernaculum est.
EZRA|7|16|Et omne argentum et aurum, quodcumque inveneris in universa provincia Babylonis simul cum oblationibus sponte oblatis a populo et a sacerdotibus pro domo Dei sui, quae est in Ierusalem,
EZRA|7|17|igitur studiose eme de hac pecunia boves, arietes, agnos et oblationes et libamina eorum et offer ea super altare templi Dei vestri, quod est in Ierusalem.
EZRA|7|18|Sed et, si quid tibi et fratribus tuis placuerit de reliquo argento et auro ut faciatis iuxta voluntatem Dei vestri, facite.
EZRA|7|19|Vasa quoque, quae dantur tibi in ministerium domus Dei tui, trade in conspectu Dei in Ierusalem.
EZRA|7|20|Sed et cetera, quibus opus fuerit in domum Dei tui, quantumcumque necesse est ut expendas, dabitur ab aerario regis.
EZRA|7|21|Et ego Artaxerxes rex statui atque decrevi omnibus custodibus arcae publicae, qui sunt trans flumen, ut quodcumque petierit a vobis Esdras sacerdos, scriba legis Dei caeli, absque mora detis
EZRA|7|22|usque ad argenti talenta centum et usque ad frumenti coros centum et usque ad vini batos centum et usque ad batos olei centum; sal vero absque mensura.
EZRA|7|23|Omne, quod requirit Deus caeli, tribuatur diligenter in domo Dei caeli, ne forte irascatur contra regnum regis et filiorum eius.
EZRA|7|24|Vobis quoque notum facimus de universis sacerdotibus et Levitis et cantoribus et ianitoribus, oblatis et ministris domus Dei huius, ut tributum et annonas et vectigal non habeatis potestatem imponendi super eos.
EZRA|7|25|Tu autem, Esdra, secundum sapientiam Dei tui, quae est in manu tua, constitue praesides et iudices, ut iudicent omni populo, qui est trans flumen, his videlicet, qui noverunt legem Dei tui; sed et imperitos docete.
EZRA|7|26|Et omnis, qui non fecerit legem Dei tui et legem regis diligenter, iudicium erit de eo, sive in mortem sive in exsilium sive in damnum substantiae eius vel certe in carcerem ".
EZRA|7|27|Benedictus Dominus, Deus patrum nostrorum, qui dedit hoc in corde regis, ut glorificaret domum Domini, quae est in Ierusalem,
EZRA|7|28|et in me inclinavit misericordiam regis et consiliariorum eius et cunctorum principum eius potentium. Et ego confortatus manu Domini Dei mei, quae erat in me, congregavi de Israel principes, qui ascenderent mecum.
EZRA|8|1|Hi sunt ergo principes familiarum et genealogia eorum, qui ascenderunt mecum in regno Artaxerxis regis de Babylone:
EZRA|8|2|De filiis Phinees, Gersom. De filiis Ithamar, Daniel. De filiis David, Hattus filius Secheniae.
EZRA|8|3|De filiis Pharos, Zacharias; et cum eo numerati sunt viri centum quinquaginta.
EZRA|8|4|De filiis Phahathmoab, Elioenai filius Zaraiae, et cum eo ducenti viri.
EZRA|8|5|De filiis Zethua, Sechenia filius Iahaziel, et cum eo trecenti viri.
EZRA|8|6|De filiis Adin, Ebed filius Ionathan, et cum eo quinquaginta viri.
EZRA|8|7|De filiis Elam, Iesaias filius Athaliae, et cum eo septuaginta viri.
EZRA|8|8|De filiis Saphatiae, Zabadia filius Michael, et cum eo octoginta viri.
EZRA|8|9|De filiis Ioab, Abdia filius Iahiel, et cum eo ducenti decem et octo viri.
EZRA|8|10|De filiis Bani, Selomith filius Iosphiae, et cum eo centum sexaginta viri.
EZRA|8|11|De filiis Bebai, Zacharias filius Bebai, et cum eo viginti octo viri.
EZRA|8|12|De filiis Azgad, Iohanan filius Eccetan, et cum eo centum et decem viri.
EZRA|8|13|De filiis Adonicam ascenderunt iuniores, et haec nomina eorum: Eliphalet et Iehiel et Semeias, et cum eis sexaginta viri.
EZRA|8|14|De filiis Beguai, Uthai filius Zabud, et cum eis septuaginta viri.
EZRA|8|15|Congregavi autem eos ad fluvium, qui decurrit ad Ahava, et mansimus ibi tribus diebus. Recensui populum et sacerdotes; de filiis autem Levi non inveni ibi.
EZRA|8|16|Itaque misi Eliezer et Ariel et Semeiam et Ioiarib et Elnathan et Nathan et Zachariam et Mosollam principes sapientes.
EZRA|8|17|Et misi eos ad Eddo, qui est primus in Chasphiae loco, et posui in ore eorum verba, quae loquerentur ad Eddo et fratres eius, ut adducerent nobis ministros domus Dei nostri.
EZRA|8|18|Et adduxerunt nobis per manum Dei nostri bonam super nos virum doctissimum de filiis Moholi filii Levi filii Israel nomine Serebiam et filios eius et fratres eius decem et octo
EZRA|8|19|et Hasabiam et cum eo Iesaiam de filiis Merari filiosque eius et fratres eius viginti
EZRA|8|20|et de oblatis, quos dederant David et principes ad ministeria Levitarum, ducentos viginti viros; omnes hi suis nominibus recensiti sunt.
EZRA|8|21|Et praedicavi ibi ieiunium iuxta fluvium Ahava, ut affligeremur coram Deo nostro et peteremus ab eo iter prosperum nobis et filiis nostris universaeque substantiae nostrae.
EZRA|8|22|Erubui enim petere a rege praesidium et equites, qui defenderent nos ab inimico in via, quia dixeramus regi: " Manus Dei nostri est super omnes, qui quaerunt eum in bonitate, et potentia eius et fortitudo eius super omnes, qui derelinquunt eum ".
EZRA|8|23|Ieiunavimus autem et rogavimus Deum nostrum per hoc, et evenit nobis prospere.
EZRA|8|24|Et separavi de principibus sacerdotum duodecim, Serebiam et Hasabiam et cum eis de fratribus eorum decem,
EZRA|8|25|appendique eis argentum et aurum et vasa: tributum domus Dei nostri, quod obtulerat rex et consiliatores eius et principes eius universusque Israel eorum, qui ibi inveniebantur.
EZRA|8|26|Et appendi in manibus eorum argenti talenta sescenta quinquaginta et vasa argentea centum, quae habebant talenta duo, auri centum talenta,
EZRA|8|27|et crateres aureos viginti, qui habebant solidos millenos, et vasa aeris fulgentis optimi duo pretiosa ut aurum.
EZRA|8|28|Et dixi eis: " Vos sancti Domini, et vasa sancta et argentum et aurum consecrata Domino, Deo patrum nostrorum;
EZRA|8|29|vigilate et custodite, donec appendatis coram principibus sacerdotum et Levitarum et ducibus familiarum Israel in Ierusalem, in habitaculis domus Domini ".
EZRA|8|30|Susceperunt autem sacerdotes et Levitae pondus argenti et auri et vasorum, ut deferrent Ierusalem in domum Dei nostri.
EZRA|8|31|Promovimus ergo a flumine Ahava duodecimo die mensis primi, ut pergeremus Ierusalem; et manus Dei nostri fuit super nos et liberavit nos de manu inimici et insidiatoris in via,
EZRA|8|32|et venimus Ierusalem et mansimus ibi tribus diebus.
EZRA|8|33|Die autem quarta appensum est argentum et aurum et vasa in domo Dei nostri per manum Meremoth filii Uriae sacerdotis et cum eo Eleazar filius Phinees cumque eis Iozabad filius Iesua et Noadia filius Bennui Levitae,
EZRA|8|34|iuxta numerum et pondus omnia; descriptumque est omne pondus. In tempore illo,
EZRA|8|35|qui venerant de captivitate, filii transmigrationis, obtulerunt holocautomata Deo Israel, vitulos duodecim pro omni populo Israel, arietes nonaginta sex, agnos septuaginta septem, hircos pro peccato duodecim: omnia in holocaustum Domino.
EZRA|8|36|Dederunt autem edicta regis satrapis regis et ducibus trans flumen et sublevaverunt populum et domum Dei.
EZRA|9|1|Postquam autem haec completa sunt, accesserunt ad me princi pes dicentes: " Non est separatus populus Israel, sacerdotes et Levitae a populis terrarum et abominationibus eorum, Chananaei videlicet et Hetthaei et Pherezaei et Iebusaei et Ammonitarum et Moabitarum et Aegyptiorum et Amorraeorum.
EZRA|9|2|Tulerunt enim de filiabus eorum sibi et filiis suis et commiscuerunt semen sanctum cum populis terrarum; manus etiam principum et magistratuum fuit in transgressione hac prima ".
EZRA|9|3|Cumque audissem sermonem istum, scidi vestimentum meum et pallium et evelli capillos capitis mei et barbae et sedi maerens.
EZRA|9|4|Convenerunt autem ad me omnes, qui timebant verba Dei Israel pro transgressione eorum, qui de captivitate venerant; et ego sedebam tristis usque ad sacrificium vespertinum.
EZRA|9|5|Et in sacrificio vespertino surrexi de afflictione mea et, scisso vestimento et pallio, curvavi genua mea et expandi manus meas ad Dominum Deum meum.
EZRA|9|6|Et dixi: " Deus meus, confundor et erubesco levare faciem meam ad te, quoniam iniquitates nostrae multiplicatae sunt super caput nostrum, et delicta nostra creverunt usque ad caelum
EZRA|9|7|a diebus patrum nostrorum. Peccavimus graviter usque ad diem hanc, et propter iniquitates nostras traditi sumus, ipsi et reges nostri et sacerdotes nostri, in manum regum terrarum et in gladium et in captivitatem et in rapinam et in confusionem vultus sicut et die hac.
EZRA|9|8|Et nunc ad momentum invenimus gratiam apud Dominum Deum nostrum, ut servaret nobis reliquias et figeret nobis tentorium in loco sancto eius et illuminaret oculos nostros Deus noster et daret nobis solacium modicum in servitute nostra.
EZRA|9|9|Quia servi sumus, et in servitute nostra non dereliquit nos Deus noster, sed inclinavit super nos misericordiam regum Persarum, ut darent nobis solacium, et erigeretur domus Dei nostri, et instaurarentur ruinae eius, et dedit nobis refugium in Iuda et Ierusalem.
EZRA|9|10|Et nunc quid dicemus, Deus noster, post haec? Dereliquimus mandata tua,
EZRA|9|11|quae praecepisti in manu servorum tuorum prophetarum dicens: "Terra, ad quam vos ingredimini, ut possideatis eam, terra immunda est, iuxta immunditiam populorum terrarum et abominationem eorum, qui repleverunt eam a fine usque ad finem coinquinatione sua.
EZRA|9|12|Nunc ergo filias vestras ne detis filiis eorum et filias eorum ne accipiatis filiis vestris et non quaeratis pacem eorum et prosperitatem eorum usque in aeternum, ut confortemini et comedatis, quae bona sunt terrae, et heredes habeatis filios vestros usque in saeculum".
EZRA|9|13|Et post omnia, quae venerunt super nos in operibus nostris pessimis et in delicto nostro magno, quia tu, Deus noster, non iudicasti secundum iniquitates nostras et dedisti nobis salutem, sicut est hodie,
EZRA|9|14|numquid amplius irrita faciemus mandata tua et matrimonia iungemus cum populis abominationum istarum? Numquid iratus es nobis usque ad consummationem, ut non essent reliquiae et salus?
EZRA|9|15|Domine, Deus Israel, tua clementia superstites sumus sicut die hac! Ecce coram te sumus in delicto nostro; non enim stari potest coram te propter hoc ".
EZRA|10|1|Dum ergo oraret Esdras et imploraret flens et prostratus ante templum Dei, collectus est ad eum de Israel coetus grandis nimis virorum et mulierum et puerorum; et flevit populus fletu multo.
EZRA|10|2|Et respondit Sechenias filius Iehiel de filiis Elam et dixit Esdrae: " Nos praevaricati sumus in Deum nostrum et duximus uxores alienigenas de populis terrae. Nunc autem spes est in Israel super hoc:
EZRA|10|3|percutiamus foedus cum Domino Deo nostro, ut proiciamus universas uxores et eos, qui de his nati sunt, iuxta voluntatem Domini et eorum, qui timent praeceptum Domini Dei nostri, et secundum legem fiat.
EZRA|10|4|Surge, tuum est decernere, nosque erimus tecum; confortare et fac ".
EZRA|10|5|Surrexit ergo Esdras et fecit principes sacerdotum et Levitarum et omnem Israel iurare, ut facerent secundum verbum hoc, et iuraverunt.
EZRA|10|6|Et surrexit Esdras ante domum Dei et abiit ad cubiculum Iohanan filii Eliasib et pernoctavit ibi; panem non comedit et aquam non bibit, lugebat enim transgressionem eorum, qui venerant de captivitate.
EZRA|10|7|Et missa est vox in Iuda et in Ierusalem omnibus filiis transmigrationis, ut congregarentur in Ierusalem;
EZRA|10|8|et omnis, qui non venerit in tribus diebus iuxta consilium principum et seniorum, auferetur universa substantia eius, et ipse abicietur de coetu transmigrationis.
EZRA|10|9|Convenerunt igitur omnes viri Iudae et Beniamin in Ierusalem tribus diebus, ipse est mensis nonus vicesimo die mensis, et sedit omnis populus in platea domus Dei, trementes pro peccato et pluviis.
EZRA|10|10|Et surrexit Esdras sacerdos et dixit ad eos: " Vos transgressi estis et duxistis uxores alienigenas, ut adderetis super delictum Israel.
EZRA|10|11|Et nunc date confessionem Domino, Deo patrum vestrorum, et facite placitum eius et separamini a populis terrae et ab uxoribus alienigenis ".
EZRA|10|12|Et respondit universa multitudo dixitque voce magna: " Iuxta verbum tuum ad nos, sic fiat.
EZRA|10|13|Verumtamen quia populus multus est et tempus pluviae, et non sustinemus stare foris, et opus non est diei unius vel duorum - multi quippe peccavimus in sermone isto -
EZRA|10|14|constituantur principes in universa multitudine; et omnes in civitatibus nostris, qui duxerunt uxores alienigenas, veniant in temporibus statutis, et cum his seniores per civitatem et civitatem et iudices eius, donec avertatur ira Dei nostri a nobis super peccato hoc ".
EZRA|10|15|Tantummodo Ionathan filius Asael et Iaasia filius Thecue steterunt contra hoc, et Mosollam et Sabethai Levites adiuverunt eos.
EZRA|10|16|Feceruntque sic filii transmigrationis. Et elegit Esdras sacerdos viros principes familiarum iuxta domus patrum eorum, omnes autem per nomina eorum, et sederunt in die primo mensis decimi, ut quaererent rem.
EZRA|10|17|Et absolverunt causam cunctorum, qui duxerant uxores alienigenas, intra diem primam mensis primi.
EZRA|10|18|Et inventi sunt de filiis sacerdotum, qui duxerant uxores alienigenas. De filiis Iesua filii Iosedec et de fratribus eius: Maasia et Eliezer et Iarib et Godolia;
EZRA|10|19|et dederunt manus suas, ut eicerent uxores suas et pro delicto suo arietem offerrent.
EZRA|10|20|Et de filiis Emmer: Hanani et Zabadia.
EZRA|10|21|Et de filiis Harim: Maasia et Elia et Semeia et Iehiel et Ozias.
EZRA|10|22|Et de filiis Phassur: Elioenai, Maasia, Ismael, Nathanael, Iozabad et Elasa.
EZRA|10|23|Et de filiis Levitarum: Iozabad et Semei et Celaia, ipse est Celita, Phethahia, Iuda et Eliezer.
EZRA|10|24|Et de cantoribus: Eliasib. Et de ianitoribus: Sellum et Telem et Uri.
EZRA|10|25|Et ex Israel de filiis Pharos: Remia et Iezia et Melchia et Miamin et Eleazar et Melchia et Banaia.
EZRA|10|26|Et de filiis Elam: Matthania, Zacharias et Iehiel et Abdi et Ierimoth et Elia.
EZRA|10|27|Et de filiis Zethua: Elioenai, Eliasib, Matthania et Ierimoth et Zabad et Aziza.
EZRA|10|28|Et de filiis Bebai: Iohanan, Hanania, Zabbai, Athalai.
EZRA|10|29|Et de filiis Beguai: Mosollam et Melluch et Adaia, Iasub et Saal et Ramoth.
EZRA|10|30|Et de filiis Phahathmoab: Edna et Chalal, Banaias et Maasias, Matthanias, Beseleel, Bennui et Manasse.
EZRA|10|31|Et de filiis Harim: Eliezer, Iesia, Melchias, Semeias, Simeon,
EZRA|10|32|Beniamin, Melluch, Samarias.
EZRA|10|33|Et de filiis Hasum: Matthanai, Matthatha, Zabad, Eliphalet, Iermai, Manasse, Semei.
EZRA|10|34|De filiis Bani: Maaddi, Amram et Ioel,
EZRA|10|35|Banaia et Badaias, Cheliau,
EZRA|10|36|Vania, Meremoth et Eliasib,
EZRA|10|37|Matthanias, Matthanai et Iasi.
EZRA|10|38|Et de filiis Bennui: Semei
EZRA|10|39|et Selemias et Nathan et Adaias
EZRA|10|40|et Mechnedebai, Sisai, Sarai,
EZRA|10|41|Azareel et Selemias, Samaria,
EZRA|10|42|Sellum, Amaria, Ioseph.
EZRA|10|43|De filiis Nabo: Iehiel, Matthathias, Zabad, Zabina, Ieddu et Ioel et Banaia.
EZRA|10|44|Omnes hi acceperant uxores alienigenas et dimiserunt uxores et filios.
