1PET|1|1|Petrus apostolus Iesu Christi electis advenis dispersionis Pon ti, Galatiae, Cappadociae, Asiae et Bithyniae,
1PET|1|2|secundum praescientiam Dei Patris, in sanctificatione Spiritus, in oboedientiam et aspersionem sanguinis Iesu Christi: gratia vobis et pax multiplicetur.
1PET|1|3|Benedictus Deus et Pater Domini nostri Iesu Christi, qui secundum magnam misericordiam suam regeneravit nos in spem vivam per resurrectionem Iesu Christi ex mortuis,
1PET|1|4|in hereditatem incorruptibilem et incontaminatam et immarcescibilem, conservatam in caelis propter vos,
1PET|1|5|qui in virtute Dei custodimini per fidem in salutem, paratam revelari in tempore novissimo.
1PET|1|6|In quo exsultatis, modicum nunc si oportet contristati in variis tentationibus,
1PET|1|7|ut probatio vestrae fidei multo pretiosior auro, quod perit, per ignem quidem probato, inveniatur in laudem et gloriam et honorem in revelatione Iesu Christi.
1PET|1|8|Quem cum non videritis, diligitis; in quem nunc non videntes, credentes autem, exsultatis laetitia inenarrabili et glorificata,
1PET|1|9|reportantes finem fidei vestrae salutem animarum.
1PET|1|10|De qua salute exquisierunt atque scrutati sunt prophetae, qui de futura in vos gratia prophetaverunt,
1PET|1|11|scrutantes in quod vel quale tempus significaret, qui erat in eis Spiritus Christi, praenuntians eas, quae in Christo sunt, passiones et posteriores glorias;
1PET|1|12|quibus revelatum est quia non sibi ipsis, vobis autem ministrabant ea, quae nunc nuntiata sunt vobis per eos, qui evangelizaverunt vos, Spiritu Sancto misso de caelo, in quae desiderant angeli prospicere.
1PET|1|13|Propter quod succincti lumbos mentis vestrae, sobrii, perfecte sperate in eam, quae offertur vobis, gratiam in revelatione Iesu Christi.
1PET|1|14|Quasi filii oboedientiae, non configurati prioribus in ignorantia vestra desideriis,
1PET|1|15|sed secundum eum, qui vocavit vos, sanctum, et ipsi sancti in omni conversatione sitis,
1PET|1|16|quoniam scriptum est: " Sancti eritis, quia ego sanctus sum ".
1PET|1|17|Et si Patrem invocatis eum, qui sine acceptione personarum iudicat secundum uniuscuiusque opus, in timore incolatus vestri tempore conversamini,
1PET|1|18|scientes quod non corruptibilibus argento vel auro redempti estis de vana vestra conversatione a patribus tradita,
1PET|1|19|sed pretioso sanguine quasi Agni incontaminati et immaculati Christi,
1PET|1|20|praecogniti quidem ante constitutionem mundi, manifestati autem novissimis temporibus propter vos,
1PET|1|21|qui per ipsum fideles estis in Deum, qui suscitavit eum a mortuis et dedit ei gloriam, ut fides vestra et spes esset in Deum.
1PET|1|22|Animas vestras castificantes in oboedientia veritatis ad fraternitatis amorem non fictum, ex corde invicem diligite attentius,
1PET|1|23|renati non ex semine corruptibili sed incorruptibili per verbum Dei vivum et permanens:
1PET|1|24|quiaomnis caro ut fenum,et omnis gloria eius tamquam flos feni.Exaruit fenum, et flos decidit;
1PET|1|25|verbum autem Domini manet in aeternum.Hoc est autem verbum, quod evangelizatum est in vos.
1PET|2|1|Deponentes igitur omnem ma litiam et omnem dolum et simu lationes et invidias et omnes detractiones,
1PET|2|2|sicut modo geniti infantes, rationale sine dolo lac concupiscite, ut in eo crescatis in salutem,
1PET|2|3|si gustastis quoniam dulcis Dominus.
1PET|2|4|Ad quem accedentes, lapidem vivum, ab hominibus quidem reprobatum, coram Deo autem electum, pretiosum,
1PET|2|5|et ipsi tamquam lapides vivi aedificamini domus spiritalis in sacerdotium sanctum offerre spiritales hostias acceptabiles Deo per Iesum Christum.
1PET|2|6|Propter quod continet Scriptura: Ecce pono in Sion lapidem angularem, electum, pretiosum;et, qui credit in eo, non confundetur ".
1PET|2|7|Vobis igitur honor credentibus; non credentibus autem Lapis, quem reprobaverunt aedificantes, hic factus est in caput anguli "
1PET|2|8|et " lapis offensionis et petra scandali "; qui offendunt verbo non credentes, in quod et positi sunt.
1PET|2|9|Vos autem genus electum, regale sacerdotium, gens sancta, populus in acquisitionem, ut virtutes annuntietis eius, qui de tenebris vos vocavit in admirabile lumen suum:
1PET|2|10|qui aliquando non populus, nunc autem populus Dei; qui non consecuti misericordiam, nunc autem misericordiam consecuti.
1PET|2|11|Carissimi, obsecro tamquam advenas et peregrinos abstinere vos a carnalibus desideriis, quae militant adversus animam;
1PET|2|12|conversationem vestram inter gentes habentes bonam, ut in eo, quod detrectant de vobis tamquam de malefactoribus, ex bonis operibus considerantes glorificent Deum in die visitationis.
1PET|2|13|Subiecti estote omni humanae creaturae propter Dominum: sive regi quasi praecellenti
1PET|2|14|sive ducibus tamquam ab eo missis ad vindictam malefactorum, laudem vero bonorum;
1PET|2|15|quia sic est voluntas Dei, ut benefacientes obmutescere faciatis imprudentium hominum ignorantiam,
1PET|2|16|quasi liberi, et non quasi velamen habentes malitiae libertatem, sed sicut servi Dei.
1PET|2|17|Omnes honorate, fraternitatem diligite, Deum timete, regem honorificate.
1PET|2|18|Servi, subditi estote in omni timore dominis, non tantum bonis et modestis sed etiam pravis.
1PET|2|19|Haec est enim gratia, si propter conscientiam Dei sustinet quis tristitias, patiens iniuste.
1PET|2|20|Quae enim gloria est, si peccantes et colaphizati sustinetis? Sed si benefacientes et patientes sustinetis, haec est gratia apud Deum.
1PET|2|21|In hoc enim vocati estis, quiaet Christus passus est pro vobis,vobis relinquens exemplum,ut sequamini vestigia eius:
1PET|2|22|qui peccatum non fecit,nec inventus est dolus in ore ipsius;
1PET|2|23|qui cum malediceretur, non remaledicebat;cum pateretur, non comminabatur, commendabat autem iuste iudicanti;
1PET|2|24|qui peccata nostra ipse pertulitin corpore suo super lignum,ut peccatis mortui iustitiae viveremus;cuius livore sanati estis.
1PET|2|25|Eratis enim sicut oves errantes,sed conversi estis nunc ad pastorem et episcopum animarum vestrarum.
1PET|3|1|Similiter mulieres subditae sint suis viris, ut et si qui non cre dunt verbo, per mulierum conversationem sine verbo lucrifiant,
1PET|3|2|considerantes castam in timore conversationem vestram;
1PET|3|3|quarum sit non extrinsecus capillaturae aut circumdationis auri aut indumenti vestimentorum cultus,
1PET|3|4|sed qui absconditus cordis est homo, in incorruptibilitate mitis et quieti spiritus, qui est in conspectu Dei locuples.
1PET|3|5|Sic enim aliquando et sanctae mulieres sperantes in Deo ornabant se subiectae propriis viris,
1PET|3|6|sicut Sara oboediebat Abrahae dominum eum vocans: cuius estis filiae benefacientes et non timentes ullam perturbationem.
1PET|3|7|Viri similiter cohabitantes secundum scientiam quasi infirmiori vaso muliebri impertientes honorem, tamquam et coheredibus gratiae vitae, uti ne impediantur orationes vestrae.
1PET|3|8|In fine autem omnes unanimes, compatientes, fraternitatis amatores, misericordes, humiles,
1PET|3|9|non reddentes malum pro malo vel maledictum pro maledicto, sed e contrario benedicentes, quia in hoc vocati estis, ut benedictionem hereditate accipiatis.
1PET|3|10|" Qui enim vult vitam diligereet videre dies bonos,coerceat linguam suam a malo,
1PET|3|11|et labia eius ne loquantur dolum;declinet autem a malo et faciat bonum,inquirat pacem et persequatur eam.
1PET|3|12|Quia oculi Domini super iustos,et aures eius in preces eorum;vultus autem Domini super facientes mala ".
1PET|3|13|Et quis est qui vobis noceat, si boni aemulatores fueritis?
1PET|3|14|Sed et si patimini propter iustitiam, beati! Timorem autem eorum ne timueritis et non conturbemini,
1PET|3|15|Dominum autem Christum sanctificate in cordibus vestris, parati semper ad defensionem omni poscenti vos rationem de ea, quae in vobis est spe;
1PET|3|16|sed cum mansuetudine et timore, conscientiam habentes bonam, ut in quo de vobis detrectatur, confundantur, qui calumniantur vestram bonam in Christo conversationem.
1PET|3|17|Melius est enim benefacientes, si velit voluntas Dei, pati quam malefacientes.
1PET|3|18|Quia et Christus semel pro peccatis passus est, iustus pro iniustis, ut vos adduceret ad Deum, mortificatus quidem carne, vivificatus autem Spiritu:
1PET|3|19|in quo et his, qui in carcere erant, spiritibus adveniens praedicavit,
1PET|3|20|qui increduli fuerant aliquando, quando exspectabat Dei patientia in diebus Noe, cum fabricaretur arca, in qua pauci, id est octo animae, salvae factae sunt per aquam.
1PET|3|21|Cuius antitypum, baptisma, et vos nunc salvos facit, non carnis depositio sordium sed conscientiae bonae rogatio in Deum, per resurrectionem Iesu Christi,
1PET|3|22|qui est in dextera Dei, profectus in caelum, subiectis sibi angelis et potestatibus et virtutibus.
1PET|4|1|Christo igitur passo in carne, et vos eadem cogitatione armami ni, quia, qui passus est carne, desiit a peccato;
1PET|4|2|ut iam non hominum concupiscentiis sed voluntate Dei, quod reliquum est in carne vivat temporis.
1PET|4|3|Sufficit enim praeteritum tempus ad voluntatem gentium consummandam, vobis, qui ambulastis in luxuriis, concupiscentiis, vinolentiis, comissationibus, potationibus et illicitis idolorum cultibus.
1PET|4|4|In quo mirantur non concurrentibus vobis in eandem luxuriae effusionem, blasphemantes;
1PET|4|5|qui reddent rationem ei, qui paratus est iudicare vivos et mortuos.
1PET|4|6|Propter hoc enim et mortuis evangelizatum est, ut iudicentur quidem secundum homines carne, vivant autem secundum Deum Spiritu.
1PET|4|7|Omnium autem finis appropinquavit. Estote itaque prudentes et vigilate in orationibus.
1PET|4|8|Ante omnia mutuam in vosmetipsos caritatem continuam habentes, quia caritas operit multitudinem peccatorum;
1PET|4|9|hospitales invicem sine murmuratione;
1PET|4|10|unusquisque, sicut accepit donationem, in alterutrum illam administrantes, sicut boni dispensatores multiformis gratiae Dei.
1PET|4|11|Si quis loquitur, quasi sermones Dei; si quis ministrat, tamquam ex virtute, quam largitur Deus, ut in omnibus glorificetur Deus per Iesum Christum: cui est gloria et imperium in saecula saeculorum. Amen.
1PET|4|12|Carissimi, nolite mirari in fervore, qui ad tentationem vobis fit, quasi novi aliquid vobis contingat,
1PET|4|13|sed, quemadmodum communicatis Christi passionibus, gaudete, ut et in revelatione gloriae eius gaudeatis exsultantes.
1PET|4|14|Si exprobramini in nomine Christi, beati, quoniam Spiritus gloriae et Dei super vos requiescit.
1PET|4|15|Nemo enim vestrum patiatur quasi homicida aut fur aut maleficus aut alienorum speculator;
1PET|4|16|si autem ut christianus, non erubescat, glorificet autem Deum in isto nomine.
1PET|4|17|Quoniam tempus est, ut incipiat iudicium a domo Dei; si autem primum a nobis, qui finis eorum, qui non credunt Dei evangelio?
1PET|4|18|" Et si iustus vix salvatur,impius et peccator ubi parebit? ".
1PET|4|19|Itaque et hi, qui patiuntur secundum voluntatem Dei, fideli Creatori commendent animas suas in benefacto.
1PET|5|1|Seniores ergo, qui in vobis sunt, obsecro, consenior et testis Chri sti passionum, qui et eius, quae in futuro revelanda est, gloriae communicator:
1PET|5|2|Pascite, qui est in vobis, gregem Dei, providentes non coacto sed spontanee secundum Deum, neque turpis lucri gratia sed voluntarie,
1PET|5|3|neque ut dominantes in cleris sed formae facti gregis.
1PET|5|4|Et cum apparuerit Princeps pastorum, percipietis immarcescibilem gloriae coro nam.
1PET|5|5|Similiter, adulescentes, subditi estote senioribus. Omnes autem invicem humilitatem induite, quiaDeus superbis resistit,humilibus autem dat gratiam.
1PET|5|6|Humiliamini igitur sub potenti manu Dei, ut vos exaltet in tempore,
1PET|5|7|omnem sollicitudinem vestram proicientes in eum, quoniam ipsi cura est de vobis.
1PET|5|8|Sobrii estote, vigilate. Adversarius vester Diabolus tamquam leo rugiens circuit quaerens quem devoret.
1PET|5|9|Cui resistite fortes fide, scientes eadem passionum ei, quae in mundo est, vestrae fraternitati fieri.
1PET|5|10|Deus autem omnis gratiae, qui vocavit vos in aeternam suam gloriam in Christo Iesu, modicum passos ipse perficiet, confirmabit, solidabit, fundabit.
1PET|5|11|Ipsi imperium in saecula saeculorum. Amen.
1PET|5|12|Per Silvanum vobis fidelem fratrem, ut arbitror, breviter scripsi, obsecrans et contestans hanc esse veram gratiam Dei; in qua state.
1PET|5|13|Salutat vos, quae est in Babylone, coelecta et Marcus filius meus.
1PET|5|14|Salutate invicem in osculo caritatis.Pax vobis omnibus, qui estis in Christo.
