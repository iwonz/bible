PROV|1|1|大卫 的儿子， 以色列 王 所罗门 的箴言：
PROV|1|2|要使人懂得智慧和训诲， 明白通达的言语，
PROV|1|3|使人领受明智的训诲， 就是公义、公平和正直，
PROV|1|4|使愚蒙人灵巧， 使年轻人有知识，有智谋。
PROV|1|5|智慧人听见，增长学问， 聪明人得着智谋，
PROV|1|6|明白箴言和譬喻， 懂得智慧人的言词和谜语。
PROV|1|7|敬畏耶和华是知识的开端； 愚妄人藐视智慧和训诲。
PROV|1|8|我儿啊，要听你父亲的训诲， 不可离弃你母亲的教诲；
PROV|1|9|因为这要作你头上恩惠的华冠， 作你颈上的项链。
PROV|1|10|我儿啊，罪人若引诱你， 你不可随从。
PROV|1|11|他们若说：“你与我们同去， 我们要埋伏杀人流血， 无故地潜藏，杀害无辜；
PROV|1|12|我们好像阴间，把他们活活吞下， 囫囵吞下，如吞下那下到地府的人；
PROV|1|13|我们必得各样宝物， 将所夺来的装满房屋；
PROV|1|14|你来与我们同伙， 共用一个钱囊。”
PROV|1|15|我儿啊，不要与他们走同一道路， 禁止你的脚走他们的路径。
PROV|1|16|因为他们的脚奔跑行恶， 他们急速杀人流血。
PROV|1|17|在飞鸟眼前张设网罗， 一定会徒劳无功；
PROV|1|18|同样，他们埋伏，是自流己血， 他们潜藏，是自害己命。
PROV|1|19|凡靠暴力敛财的，所行之路都是如此， 这种念头必夺去自己的生命。
PROV|1|20|智慧 在街市上呼喊， 在广场上高声呐喊，
PROV|1|21|在热闹街头呼叫， 在城门口，在城中，发出言语，说：
PROV|1|22|“你们无知的人喜爱无知， 傲慢人喜欢傲慢， 愚昧人恨恶知识， 要到几时呢？
PROV|1|23|你们当因我的责备回转， 我要将我的灵浇灌你们， 将我的话指示你们。
PROV|1|24|因为我呼唤，你们不听， 我招手，无人理会。
PROV|1|25|你们忽视我一切的劝戒， 拒听我的责备。
PROV|1|26|你们遭难，我就发笑； 惊恐临到你们， 惊恐如狂风来临， 灾难好像暴风来到， 急难痛苦临到你们身上， 我必嗤笑。
PROV|1|27|
PROV|1|28|那时，他们就会呼求我，我却不回答， 恳切寻求我，却寻不见。
PROV|1|29|因为他们恨恶知识， 选择不敬畏耶和华，
PROV|1|30|不听我的劝戒， 藐视我一切的责备，
PROV|1|31|所以他们要自食其果， 饱胀在自己的计谋中。
PROV|1|32|愚蒙人背道，害死自己， 愚昧人安逸，自取灭亡。
PROV|1|33|惟听从我的，必安然居住， 得享宁静，不怕灾祸。”
PROV|2|1|我儿啊，你若领受我的言语， 珍藏我的命令，
PROV|2|2|留心听智慧， 专心求聪明；
PROV|2|3|你若呼求明理， 扬声求聪明，
PROV|2|4|寻找她，如寻找银子， 搜寻她，如搜寻宝藏，
PROV|2|5|你就懂得敬畏耶和华， 得以认识上帝。
PROV|2|6|因为耶和华赏赐智慧， 知识和聪明都由他口而出。
PROV|2|7|他为正直人珍藏健全的知识， 给行为纯正的人作盾牌，
PROV|2|8|为要保护公正的路， 庇护虔诚人的道。
PROV|2|9|那时，你就明白公义、公平、 正直，和一切完善的道路。
PROV|2|10|因为智慧要进入你的心， 知识要使你内心欢愉。
PROV|2|11|智谋要庇护你， 聪明必保护你，
PROV|2|12|救你脱离恶人的道， 脱离言谈乖谬的人。
PROV|2|13|他们离弃正直的路， 行走黑暗的道，
PROV|2|14|喜欢作恶， 喜爱恶人的错谬。
PROV|2|15|他们的路歪曲， 他们偏离中道。
PROV|2|16|智慧要救你远离陌生女子， 远离那油嘴滑舌的外邦女子。
PROV|2|17|她离弃年轻时的配偶， 忘了自己神圣的盟约。
PROV|2|18|她的家陷入死亡， 她的路偏向阴魂。
PROV|2|19|凡到她那里去的，不得回转， 也得不到生命的路。
PROV|2|20|智慧使你行善人的道， 守义人的路。
PROV|2|21|正直人必在地上居住， 完全人必在其上存留；
PROV|2|22|惟恶人要从地上剪除， 奸诈人要被拔出。
PROV|3|1|我儿啊，不要忘记我的教诲， 你的心要谨守我的命令，
PROV|3|2|因为它们 必加给你长久的日子， 生命的年数与平安。
PROV|3|3|不可使慈爱和诚信离开你， 要系在你颈项上，刻在你心版上。
PROV|3|4|这样，你必在上帝和世人眼前 蒙恩惠，有美好的见识。
PROV|3|5|你要专心仰赖耶和华， 不可倚靠自己的聪明，
PROV|3|6|在你一切所行的路上都要认定他， 他必使你的道路平直。
PROV|3|7|不要自以为有智慧； 要敬畏耶和华，远离恶事。
PROV|3|8|这便医治你的肉体 ， 滋润你的百骨。
PROV|3|9|你要以财物 和一切初熟的土产尊崇耶和华，
PROV|3|10|这样，你的仓库必充满有余， 你的酒池有新酒盈溢。
PROV|3|11|我儿啊，不可轻看耶和华的管教， 也不可厌烦他的责备，
PROV|3|12|因为耶和华所爱的，他必责备， 正如父亲责备所喜爱的儿子。
PROV|3|13|得智慧，得聪明的， 这人有福了。
PROV|3|14|因为智慧的获利胜过银子， 所得的盈余强如金子，
PROV|3|15|比宝石 更宝贵， 你一切所喜爱的，都不足与其比较。
PROV|3|16|她的右手有长寿， 左手有富贵。
PROV|3|17|她的道是安乐， 她的路全是平安。
PROV|3|18|她给持守她的人作生命树， 谨守她的必定蒙福。
PROV|3|19|耶和华以智慧奠立地基， 以聪明铺设诸天，
PROV|3|20|以知识使深渊裂开， 使天空滴下甘露。
PROV|3|21|我儿啊，要谨守健全的知识和智谋， 不可使它们偏离你的眼目。
PROV|3|22|这样，它们必使你的生命有活力， 又作你颈项的美饰。
PROV|3|23|那时，你就坦然行路， 不致跌倒。
PROV|3|24|你躺下，必不惧怕； 你躺卧，睡得香甜。
PROV|3|25|忽然来的惊恐，你不要害怕； 恶人遭毁灭，也不要恐惧，
PROV|3|26|因为耶和华是你的倚靠， 他必保护你的脚不陷入罗网。
PROV|3|27|你的手若有行善的力量， 不可推辞，要施与那应得的人。
PROV|3|28|你若手头方便， 不可对邻舍说： “去吧，明天再来，我必给你。”
PROV|3|29|你的邻舍既在你附近安居， 不可设计害他。
PROV|3|30|人若未曾加害你， 不可无故与他相争。
PROV|3|31|不可嫉妒残暴的人， 不可选择他的任何道路。
PROV|3|32|因为走偏方向的人是耶和华所憎恶的； 正直人为他所亲密。
PROV|3|33|耶和华诅咒恶人的家； 义人的居所他却赐福。
PROV|3|34|他讥诮那爱讥诮的人； 但赐恩给谦卑的人。
PROV|3|35|智慧人必承受尊荣； 愚昧人高升却是羞辱。
PROV|4|1|孩子们，要听父亲的训诲， 留心明白道理。
PROV|4|2|因我给你们好的教导， 不可离弃我的教诲。
PROV|4|3|当我在父亲面前还是小孩， 是母亲独一娇儿的时候，
PROV|4|4|他教导我说：“你的心要持守我的话， 遵守我的命令，你就会存活。
PROV|4|5|要获得智慧，要获得聪明， 不可忘记， 也不可偏离我口中的言语。
PROV|4|6|不可离弃智慧，智慧就庇护你， 要爱她，她就保护你。
PROV|4|7|智慧为首，所以要获得智慧， 要用你一切所有的换取聪明。
PROV|4|8|高举智慧，她就使你升高， 拥抱智慧，她就使你尊荣。
PROV|4|9|她必将恩惠的华冠加在你头上， 把荣冕赐给你。”
PROV|4|10|我儿啊，要听，要领受我的言语， 你就必延年益寿。
PROV|4|11|我已指教你走智慧的道， 引导你行正直的路。
PROV|4|12|你行走，脚步没有阻碍； 你奔跑，也不致跌倒。
PROV|4|13|要持定训诲，不可放松； 要谨守它，因为它是你的生命。
PROV|4|14|不可行恶人的路， 不要走坏人的道；
PROV|4|15|要躲避，不可经过， 要转离而去。
PROV|4|16|他们若不行恶，难以成眠， 不使人跌倒，就睡卧不安；
PROV|4|17|因为他们以邪恶当饼吃， 以暴力当酒喝。
PROV|4|18|但义人的路好像黎明的光， 越照越明，直到正午。
PROV|4|19|恶人的道幽暗， 自己不知因何跌倒。
PROV|4|20|我儿啊，要留心听我的话， 侧耳听我的言语，
PROV|4|21|不可使它们偏离你的眼目， 要存记在你心中。
PROV|4|22|因为找到它们的，就找到生命， 得到全身的医治。
PROV|4|23|你要保守你心，胜过保守一切， 因为生命的泉源由心发出。
PROV|4|24|要离开歪曲的口， 转离偏邪的嘴唇。
PROV|4|25|你的两眼要向前看， 你的双目 直视前方。
PROV|4|26|要修平 你脚下的路， 你一切的道就必稳固。
PROV|4|27|不可偏左偏右， 你的脚要离开邪恶。
PROV|5|1|我儿啊，要留心听我的智慧， 侧耳听我的聪明，
PROV|5|2|为要使你谨守智谋， 嘴唇保护知识。
PROV|5|3|因为陌生女子的嘴唇滴下蜂蜜， 她的口比油更滑，
PROV|5|4|后来却苦似茵蔯， 锐利如两刃的剑。
PROV|5|5|她的脚坠落死亡， 她的脚步踏入阴间，
PROV|5|6|她无法找到生命的道路， 她的路变迁不定，自己却不知道。
PROV|5|7|孩子们，现在要听从我， 不可离弃我口中的言语。
PROV|5|8|你所行的道要远离她， 不可靠近她家的门口，
PROV|5|9|免得将你的尊荣给别人， 将你的岁月给残忍的人；
PROV|5|10|免得陌生人满得你的财富， 你劳苦所得的归入外邦人的家。
PROV|5|11|在你人生终结，你皮肉和身体衰残时， 你必唉声叹气，
PROV|5|12|说：“我为何恨恶管教， 心里轻看责备呢？
PROV|5|13|我不听从教师的话， 也没有侧耳听那教导我的。
PROV|5|14|在聚集的会众中， 我几乎坠入深渊。”
PROV|5|15|你要喝自己池中的水， 饮自己井里的活水。
PROV|5|16|你的泉源岂可溢流在外？ 你的河水岂可流到街上？
PROV|5|17|让它们惟独归你， 不可与陌生人同享。
PROV|5|18|要使你的泉源蒙福， 要喜爱你年轻时的妻子。
PROV|5|19|她如可爱的母鹿，如优美的母羊， 愿她的胸怀使你时时满足， 愿你常常迷恋她的爱情。
PROV|5|20|我儿啊，你为何迷恋陌生女子？ 为何拥抱外邦女子的胸怀？
PROV|5|21|因为人所行的道都在耶和华眼前， 他察验 人一切的路。
PROV|5|22|恶人被自己的罪孽抓住， 被自己罪恶的绳索缠绕。
PROV|5|23|他因不受管教而死亡， 因极度愚昧而走迷。
PROV|6|1|我儿啊，你若为朋友担保， 替陌生人击掌，
PROV|6|2|你就被口中的言语套住， 被嘴里的言语抓住。
PROV|6|3|我儿啊，你既落在朋友手中，当这样行才可救自己： 你要谦卑自己，去恳求你的朋友。
PROV|6|4|不要让你的眼睛睡觉， 不可容你的眼皮打盹。
PROV|6|5|要救自己，如羚羊脱离猎人的手， 如鸟脱离捕鸟人的手。
PROV|6|6|懒惰人哪， 你去察看蚂蚁的动作，就可得智慧。
PROV|6|7|蚂蚁没有领袖， 没有官长，没有君王，
PROV|6|8|尚且在夏天预备食物， 在收割时储存粮食。
PROV|6|9|懒惰人哪，你要睡到几时呢？ 你什么时候才睡醒呢？
PROV|6|10|再睡片时，打盹片时， 抱着双臂躺卧片时，
PROV|6|11|你的贫穷就如盗贼来到， 你的贫乏仿佛拿盾牌的人来临。
PROV|6|12|无赖的恶徒 行事全凭歪曲的口，
PROV|6|13|他眨眼传神， 以脚示意，用指点划，
PROV|6|14|存心乖谬， 常设恶谋，散播纷争。
PROV|6|15|所以，灾难必突然临到他， 他必顷刻被毁，无从医治。
PROV|6|16|耶和华所恨恶的有六样， 他心所憎恶的共有七样：
PROV|6|17|就是高傲的眼，撒谎的舌， 杀害无辜的手，
PROV|6|18|图谋恶计的心， 飞奔行恶的脚，
PROV|6|19|口吐谎言的假证人， 并在弟兄间散播纷争的人。
PROV|6|20|我儿啊，要遵守你父亲的命令， 不可离弃你母亲的教诲。
PROV|6|21|要常挂在你心上， 系在你颈项上。
PROV|6|22|你行走，她必引导你， 你躺卧，她必保护你， 你睡醒，她必与你谈论。
PROV|6|23|因为诫命是灯，教诲是光， 管教的责备是生命的道，
PROV|6|24|要保护你远离邪恶的妇女， 远离外邦女子谄媚的舌头。
PROV|6|25|你不要因她的美色而动心， 也不要被她的眼皮勾引。
PROV|6|26|因为连最后一块饼都会被妓女拿走 ； 有夫之妇会猎取宝贵的生命。
PROV|6|27|人若兜火在怀中， 他的衣服岂能不烧着呢？
PROV|6|28|人若走在火炭上， 他的脚岂能不烫伤呢？
PROV|6|29|与邻舍之妻同寝的，也是如此， 凡亲近她的，难免受罚。
PROV|6|30|贼因饥饿偷窃充饥， 人不藐视他，
PROV|6|31|但若被抓到，要赔偿七倍， 他必赔上家中一切财物。
PROV|6|32|与妇人行奸淫的，便是无知， 做这事的，必毁了自己。
PROV|6|33|他必受损伤和羞辱， 他的羞耻不得消除。
PROV|6|34|丈夫因嫉恨发怒， 报仇的时候绝不留情。
PROV|6|35|他不接受任何赔偿， 你送许多礼物，他也不肯和解。
PROV|7|1|我儿啊，要遵守我的言语， 存记我的命令。
PROV|7|2|遵守我的命令就得存活， 谨守我的教诲，好像保护眼中的瞳人。
PROV|7|3|要系在你指头上， 刻在你心版上。
PROV|7|4|对智慧说“你是我的姊妹”， 称呼聪明为亲人，
PROV|7|5|她就保护你远离陌生女子， 远离油嘴滑舌的外邦女子。
PROV|7|6|我曾在我房屋的窗户内， 透过窗格子往外观看，
PROV|7|7|看见在愚蒙人中， 注意到孩儿中有一个无知的青年，
PROV|7|8|从街上经过，靠近她的巷口， 直往她家的路去，
PROV|7|9|在黄昏，在傍晚， 在半夜，黑暗之中。
PROV|7|10|看哪，有一个女子来迎接他， 是妓女的打扮，有诡诈的心思。
PROV|7|11|她喧嚷，不守约束， 她的脚在家里留不住，
PROV|7|12|有时在街市，有时在广场， 或在各巷口等候。
PROV|7|13|她拉住那青年吻他， 厚着脸皮对他说：
PROV|7|14|“我已献了平安祭， 今日我还了所许的愿。
PROV|7|15|因此，我出来迎接你， 渴望见你的面，我总算找到你了！
PROV|7|16|我已在床上铺好被单， 是 埃及 麻织的花纹布，
PROV|7|17|又用没药、沉香、桂皮 薰了我的床。
PROV|7|18|你来，让我们饱享爱情，直到早晨， 让我们彼此亲爱欢乐。
PROV|7|19|因为我丈夫不在家， 出门远行，
PROV|7|20|他手带钱囊， 要到月圆才回家。”
PROV|7|21|这女子用许多巧言引诱他， 用谄媚的嘴唇催逼他。
PROV|7|22|青年立刻跟随她，好像牛去被宰杀， 又像愚妄人带着脚镣去受刑，
PROV|7|23|直到箭穿进他的肝，如同雀鸟急投罗网， 却不知会赔上自己的生命。
PROV|7|24|孩子们，现在要听从我， 要留心听我口中的言语。
PROV|7|25|你的心不可偏向她的道， 不要误入她的迷途。
PROV|7|26|因为她击倒许多人， 无数的人被她杀戮 。
PROV|7|27|她的家是在阴间之路， 下到死亡之宫。
PROV|8|1|智慧岂不呼唤？ 聪明岂不扬声？
PROV|8|2|她站立在十字路口， 在道路旁高处的顶上，
PROV|8|3|在城门旁，城门口， 入口处，她呼喊：
PROV|8|4|“人哪，我呼唤你们， 我向世人扬声。
PROV|8|5|愚蒙人哪，你们要学习灵巧， 愚昧人哪，你们的心要明辨。
PROV|8|6|你们当听，因我要说尊贵的事， 我要张开嘴唇讲正直的事。
PROV|8|7|我的口要发出真理， 我的嘴唇憎恶邪恶。
PROV|8|8|我口中的言语都是公义， 并无奸诈和歪曲。
PROV|8|9|聪明人看为正确， 有知识的，都以为正直。
PROV|8|10|你们当领受我的训诲，胜过领受银子， 宁得知识，强如得上选的金子。
PROV|8|11|“因为智慧比宝石更美， 一切可喜爱的都不足与其比较。
PROV|8|12|我－智慧以灵巧为居所， 又寻得知识和智谋。
PROV|8|13|敬畏耶和华就是恨恶邪恶； 我恨恶骄傲、狂妄、恶道，和乖谬的口。
PROV|8|14|我有策略和健全的知识， 我聪明，又有能力。
PROV|8|15|君王藉我治国， 王子藉我定公平，
PROV|8|16|王公贵族，所有公义的审判官， 都藉我掌权 。
PROV|8|17|爱我的，我也爱他， 恳切寻求我的，必寻见。
PROV|8|18|财富和尊荣在我， 恒久的财宝和繁荣 也在我。
PROV|8|19|我的果实胜过金子，强如纯金， 我的出产超乎上选的银子。
PROV|8|20|我在公义的道上走， 在公平的路中行，
PROV|8|21|使爱我的承受财产， 充满他们的库房。
PROV|8|22|“耶和华在造化的起头， 在太初创造万物之先，就有 了我。
PROV|8|23|从亘古，从太初， 未有大地以前，我已被立。
PROV|8|24|没有深渊， 没有大水的泉源，我已出生。
PROV|8|25|大山未曾奠定， 小山未有之先，我已出生。
PROV|8|26|那时，他还没有创造大地和田野， 并世上头一撮尘土。
PROV|8|27|他立高天，我在那里， 他在渊面的周围划出圆圈，
PROV|8|28|上使穹苍坚硬， 下使渊源稳固，
PROV|8|29|为沧海定出范围，使水不越过界限， 奠定大地的根基。
PROV|8|30|那时，我在他旁边为工程师， 天天充满喜乐，时时在他面前欢笑，
PROV|8|31|在他的全地欢笑， 喜爱住在人世间。
PROV|8|32|“孩子们，现在要听从我， 谨守我道的有福了。
PROV|8|33|要听训诲，得智慧， 不可弃绝。
PROV|8|34|听从我，天天在我门口守望， 在我门框旁等候的，那人有福了。
PROV|8|35|因为寻得我的，就寻得生命， 他必蒙耶和华的恩惠。
PROV|8|36|得罪我的，害了自己的生命， 凡恨恶我的，喜爱死亡。”
PROV|9|1|智慧建造房屋， 凿成七根柱子，
PROV|9|2|宰杀牲畜，调好美酒， 又摆设筵席，
PROV|9|3|派遣女仆出去， 自己在城中至高处呼唤：
PROV|9|4|“谁是愚蒙的人，让他转到这里来！” 又对那无知的人说：
PROV|9|5|“你们来，吃我的饼， 喝我调的酒。
PROV|9|6|你们要离弃愚蒙，就得存活， 并要走明智的道路。”
PROV|9|7|纠正傲慢人的，必招羞辱， 责备恶人的，必被侮辱。
PROV|9|8|不要责备傲慢人，免得他恨你； 要责备智慧人，他必爱你。
PROV|9|9|教导智慧人，他就越有智慧， 指示义人，他就增长学问。
PROV|9|10|敬畏耶和华是智慧的开端， 认识至圣者便是聪明。
PROV|9|11|藉着我，你的日子必增多， 你生命的年数也必加添。
PROV|9|12|你若有智慧，是自己有智慧； 你若傲慢，就自己承担。
PROV|9|13|愚昧的女子喧嚷， 她是愚蒙，一无所知。
PROV|9|14|她坐在自己家门口， 在城中高处的座位上，
PROV|9|15|呼唤过路的， 向那些在路上直走的人说：
PROV|9|16|“谁是愚蒙的人，让他转到这里来！” 又对那无知的人说：
PROV|9|17|“偷来的水是甜的， 暗藏的饼是美的。”
PROV|9|18|人却不知有阴魂在她那里， 她召唤的人是在阴间的深处。
PROV|10|1|所罗门的箴言： 智慧之子使父亲喜乐； 愚昧之子使母亲担忧。
PROV|10|2|不义之财毫无益处； 惟有公义能救人脱离死亡。
PROV|10|3|耶和华不使义人捱饿； 恶人所欲的，耶和华必拒绝。
PROV|10|4|手懒的，必致穷乏； 手勤的，却要富足。
PROV|10|5|夏天储存的，是智慧之子； 收割时沉睡的，是蒙羞之子。
PROV|10|6|福祉临到义人头上； 恶人的口藏匿残暴。
PROV|10|7|义人的称号带来祝福； 恶人的名字必然败坏。
PROV|10|8|智慧的心，领受诫命； 愚妄的嘴唇，必致倾倒。
PROV|10|9|行正直路的，步步安稳； 走弯曲道的，必致败露。
PROV|10|10|挤眉弄眼的，使人忧患； 愚妄的嘴唇，必致倾倒。
PROV|10|11|义人的口是生命的泉源； 恶人的口藏匿残暴。
PROV|10|12|恨能挑启争端； 爱能遮掩一切过错。
PROV|10|13|聪明人嘴里有智慧； 无知的人背上受刑杖。
PROV|10|14|智慧人积存知识； 愚妄人的口速致败坏。
PROV|10|15|有钱人的财物是他坚固的城； 贫寒人的贫乏使他败坏。
PROV|10|16|义人的报酬带来生命； 恶人的所得用来犯罪。
PROV|10|17|遵守训诲的，行在生命道上； 离弃责备的，走迷了路。
PROV|10|18|隐藏怨恨的，有说谎的嘴唇； 口出毁谤的，是愚昧人。
PROV|10|19|多言多语难免有过； 节制嘴唇是有智慧。
PROV|10|20|义人的舌如上选的银子； 恶人的心所值无几。
PROV|10|21|义人的嘴唇牧养多人； 愚妄人因无知而死亡。
PROV|10|22|耶和华所赐的福使人富足， 并不加上忧虑。
PROV|10|23|愚昧人以行恶为乐； 聪明人以智慧为乐。
PROV|10|24|恶人所怕的，必临到他； 义人的心愿，必蒙应允。
PROV|10|25|暴风一过，恶人归于无有； 义人却有永久的根基。
PROV|10|26|懒惰人使那差他的人， 如醋倒牙，如烟薰目。
PROV|10|27|敬畏耶和华使人长寿； 恶人的年岁必减少。
PROV|10|28|义人的盼望带来喜乐； 恶人的指望必致灭没。
PROV|10|29|耶和华的道是正直人的保障； 却成了作恶人的败坏。
PROV|10|30|义人永不动摇； 恶人不得住在地上。
PROV|10|31|义人的口结出智慧； 乖谬的舌必被割断。
PROV|10|32|义人的嘴唇懂得令人喜悦； 恶人的口只知乖谬。
PROV|11|1|诡诈的天平为耶和华所憎恶； 公平的法码为他所喜悦。
PROV|11|2|骄傲来，羞耻也来； 谦逊人却有智慧。
PROV|11|3|正直人的纯正必引导自己； 奸诈人的邪恶必毁灭自己。
PROV|11|4|遭怒的日子钱财无益； 惟有公义能救人脱离死亡。
PROV|11|5|完全人的义修平自己的路； 但恶人必因自己的恶跌倒。
PROV|11|6|正直人的义必拯救自己； 奸诈人必被自己的欲望缠住。
PROV|11|7|恶人一死，他的指望就灭绝； 罪人的盼望也必灭绝。
PROV|11|8|义人得脱离患难， 有恶人来代替他。
PROV|11|9|不虔敬的人用口败坏邻舍； 义人却因知识得救。
PROV|11|10|义人享福，全城喜乐； 恶人灭亡，人人欢呼。
PROV|11|11|因正直人的祝福，城必升高； 因邪恶人的口，它必倾覆。
PROV|11|12|藐视邻舍的，便是无知； 聪明人却静默不言。
PROV|11|13|到处传话的，泄漏机密； 内心老实的，保守秘密。
PROV|11|14|无智谋，民就败落； 谋士多，就必得胜。
PROV|11|15|为陌生人担保的，必受亏损； 恨恶击掌的，却得安稳。
PROV|11|16|恩慈的妇女得尊荣； 强壮的男子得财富。
PROV|11|17|仁慈的人善待自己； 残忍的人扰害己身。
PROV|11|18|恶人做事，得虚幻的报酬； 撒公义种子的，得实在的报偿。
PROV|11|19|真正行义的，必得生命； 追求邪恶的，必致死亡。
PROV|11|20|心中歪曲的，为耶和华所憎恶； 行为正直的，为他所喜悦。
PROV|11|21|击掌保证，恶人难免受罚； 义人的后裔必得拯救。
PROV|11|22|妇女美貌而无见识， 如同金环戴在猪鼻上。
PROV|11|23|义人的心愿尽是好的； 恶人的指望却带来愤怒。
PROV|11|24|有施舍的，钱财增添； 吝惜过度，反致穷乏。
PROV|11|25|慷慨待人，必然丰裕； 滋润人的，连自己也得滋润。
PROV|11|26|屯粮不卖的，百姓必诅咒他； 愿意出售的，祝福临到头上。
PROV|11|27|恳切求善的，就求得恩宠； 但那求恶的，恶必临到他。
PROV|11|28|倚靠财富的，自己必跌倒； 义人必兴旺如绿叶。
PROV|11|29|扰害己家的，必承受虚空 ； 愚妄人作心中有智慧者的仆人。
PROV|11|30|义人的果实是生命树； 智慧人必能得人。
PROV|11|31|看哪，义人在地上尚且受报， 何况恶人和罪人呢？
PROV|12|1|喜爱管教的，就是喜爱知识； 恨恶责备的，却像畜牲。
PROV|12|2|善人蒙耶和华的恩宠； 设诡计的，耶和华必定罪。
PROV|12|3|人靠恶行不能坚立； 义人的根必不动摇。
PROV|12|4|才德的妻子是丈夫的冠冕； 蒙羞的妇人使丈夫骨头朽烂。
PROV|12|5|义人的思念是公平； 恶人的计谋是诡诈。
PROV|12|6|恶人的言论埋伏流人的血； 正直人的口却拯救人。
PROV|12|7|恶人倾覆，归于无有； 义人的家却屹立不倒。
PROV|12|8|人按自己的智慧得称赞； 心中偏邪的，必被藐视。
PROV|12|9|被人藐视，但有自己仆人 的， 胜过妄自尊大，却缺乏食物。
PROV|12|10|义人顾惜他牲畜的命； 恶人的怜悯也是残忍。
PROV|12|11|耕种自己田地的，必得饱食； 追求虚浮的，却是无知。
PROV|12|12|恶人想得坏人的猎物； 义人的根结出果实。
PROV|12|13|嘴唇的过错是恶人的圈套； 但义人必脱离患难。
PROV|12|14|人因口所结的果实，必饱得美福； 人手所做的，必归到自己身上。
PROV|12|15|愚妄人所行的，在自己眼中看为正直； 惟智慧人从善如流。
PROV|12|16|愚妄人的恼怒立时显露； 通达人却能忍辱。
PROV|12|17|说出真话的，显明公义； 作假见证的，显出诡诈。
PROV|12|18|说话浮躁，犹如刺刀； 智慧人的舌头却能医治。
PROV|12|19|诚实的嘴唇永远坚立； 说谎的舌头只存片时。
PROV|12|20|图谋恶事的，心存诡诈； 劝人和睦的，便得喜乐。
PROV|12|21|义人不遭灾害； 恶人满受祸患。
PROV|12|22|说谎的嘴唇，为耶和华所憎恶； 行事诚实，为他所喜悦。
PROV|12|23|通达人隐藏知识； 愚昧人的心彰显愚昧。
PROV|12|24|殷勤人的手必掌权； 懒惰的人必服苦役。
PROV|12|25|人心忧虑，就必沉重； 一句良言，使心欢乐。
PROV|12|26|义人引导他的邻舍 ； 恶人的道叫人迷失。
PROV|12|27|懒惰的人不烤猎物； 殷勤的人却得宝贵的财物。
PROV|12|28|在公义的路上有生命； 在其道上并无死亡。
PROV|13|1|智慧之子听父亲的训诲； 傲慢人不听责备。
PROV|13|2|人因口所结的果实，必享美福； 奸诈人却意图残暴。
PROV|13|3|谨慎守口的，得保生命； 大张嘴唇的，必致败亡。
PROV|13|4|懒惰的人奢求，却无所得； 殷勤的人必然丰裕。
PROV|13|5|义人恨恶谎言； 恶人可憎可耻。
PROV|13|6|行为纯正的，有公义保护； 犯罪的，被罪恶倾覆。
PROV|13|7|假冒富足的，一无所有； 装作穷乏的，多有财物。
PROV|13|8|财富可作人的生命赎价； 穷乏人却听不见威吓的话。
PROV|13|9|义人的光使人欢喜 ； 恶人的灯要熄灭。
PROV|13|10|骄傲挑启纷争； 听劝言却有智慧。
PROV|13|11|不劳而获之财 必减少； 逐渐积蓄的必增多。
PROV|13|12|盼望迟延，令人心忧； 愿望实现，就是得到生命树。
PROV|13|13|藐视训言的，自取灭亡； 敬畏诫命的，必得善报。
PROV|13|14|智慧人的教诲是生命的泉源， 使人避开死亡的圈套。
PROV|13|15|美好的见识使人得宠； 奸诈人的道路恒久奸诈 。
PROV|13|16|通达人都凭知识行事； 愚昧人张扬自己的愚昧。
PROV|13|17|邪恶的使者必陷入祸患； 忠信的使臣带来医治。
PROV|13|18|弃绝管教的，必贫穷受辱； 领受责备的，必享尊荣。
PROV|13|19|愿望实现，心觉甘甜； 远离恶事，为愚昧人所憎恶。
PROV|13|20|与智慧人同行的，必得智慧； 和愚昧人作伴的，必受亏损。
PROV|13|21|祸患追赶罪人； 义人却得善报。
PROV|13|22|善人给子孙遗留产业； 罪人积财却归义人。
PROV|13|23|穷乏人开垦的地虽多产粮食， 却因不公而被夺走。
PROV|13|24|不忍用杖打儿子的，是恨恶他； 疼爱儿子的，勤加管教。
PROV|13|25|义人吃喝食欲满足； 恶人肚腹却是缺乏。
PROV|14|1|妇人的智慧建立家室； 愚昧却亲手拆毁它 。
PROV|14|2|行事正直的，敬畏耶和华； 偏离正路的，却藐视他。
PROV|14|3|在愚妄人的口中有骄傲的杖； 智慧人的嘴唇必保护自己。
PROV|14|4|没有牛，槽就空空； 土产丰盛却凭牛的力气。
PROV|14|5|诚实的证人不说谎； 虚假的证人口吐谎言。
PROV|14|6|傲慢人枉寻智慧； 聪明人易得知识。
PROV|14|7|不要到愚昧人面前， 你无法从他嘴唇里知道知识。
PROV|14|8|通达人的智慧使他认清自己的道路； 愚昧人的愚昧却是自欺。
PROV|14|9|愚妄人嘲笑赎愆祭 ； 但正直人蒙悦纳。
PROV|14|10|心中的苦楚，只有自己知道； 心里的喜乐，陌生人无法分享。
PROV|14|11|恶人的房屋必倒塌； 正直人的帐棚必兴旺。
PROV|14|12|有一条路，人以为正， 至终成为死亡之路。
PROV|14|13|人在喜笑中，心也会忧愁； 快乐的终点就是愁苦。
PROV|14|14|心中背道的，必满尝其果； 善人必从自己的行为得到回报。
PROV|14|15|无知的人什么话都信； 通达人谨慎自己的脚步。
PROV|14|16|智慧人有所惧怕，就远离恶事； 愚昧人却狂傲自恃。
PROV|14|17|轻易发怒的，行事愚昧； 擅长诡计的，被人恨恶。
PROV|14|18|愚蒙人承受愚昧为产业； 通达人得知识为冠冕。
PROV|14|19|坏人在善人面前俯伏； 恶人在义人门口也是如此。
PROV|14|20|穷乏人，连邻舍也恨他； 有钱人，爱他的人众多。
PROV|14|21|藐视邻舍的，这人有罪； 施恩给困苦人的，这人有福。
PROV|14|22|谋恶的，岂非走入迷途？ 谋善的，有慈爱和诚实。
PROV|14|23|任何勤劳总有收获； 仅耍嘴皮必致穷乏。
PROV|14|24|智慧人的冠冕是富有智慧； 愚昧人的愚昧终究是愚昧。
PROV|14|25|诚实作证，救人性命； 口吐谎言是诡诈。
PROV|14|26|敬畏耶和华的，大有倚靠； 他的儿女也有避难所。
PROV|14|27|敬畏耶和华是生命的泉源， 使人离开死亡的圈套。
PROV|14|28|君王的荣耀在乎民多； 没有百姓，王就衰败。
PROV|14|29|不轻易发怒的，大有聪明； 性情暴躁的，大显愚昧。
PROV|14|30|平静的心使肉体有生气； 嫉妒使骨头朽烂。
PROV|14|31|欺压贫寒人的，是蔑视造他的主； 怜悯贫穷人的，是尊敬主。
PROV|14|32|恶人因所行的恶必被推倒； 义人临死 ，有所投靠。
PROV|14|33|智慧安居在聪明人的心中， 在愚昧人的心中却不认识 。
PROV|14|34|公义使邦国高举； 罪恶是百姓的羞辱。
PROV|14|35|君王的恩宠临到智慧的臣仆； 但其愤怒临到蒙羞的臣仆。
PROV|15|1|回答柔和，使怒消退； 言语粗暴，触动怒气。
PROV|15|2|智慧人的舌善发知识； 愚昧人的口吐出愚昧。
PROV|15|3|耶和华的眼目无处不在， 恶人善人，他都鉴察。
PROV|15|4|温良的舌是生命树； 邪恶的舌使人心碎。
PROV|15|5|愚妄人藐视父亲的管教； 领受责备，使人精明。
PROV|15|6|义人家中多有财富； 恶人获利反受扰害。
PROV|15|7|智慧人的嘴传扬知识； 愚昧人的心并非如此。
PROV|15|8|恶人献祭，为耶和华所憎恶； 正直人祈祷，为他所喜悦。
PROV|15|9|恶人的道路，为耶和华所憎恶； 追求公义的，为他所喜爱。
PROV|15|10|背弃正路的，必受严刑； 恨恶责备的，必致死亡。
PROV|15|11|阴间和冥府 尚且在耶和华面前， 何况世人的心呢？
PROV|15|12|傲慢人不爱受责备， 也不去接近智慧人。
PROV|15|13|心中喜乐，面有喜色； 心里忧愁，灵就忧伤。
PROV|15|14|聪明人的心追求知识； 愚昧人的口吞吃愚昧。
PROV|15|15|困苦人的日子都是愁苦； 心中欢畅的，常享宴席。
PROV|15|16|财宝稀少，敬畏耶和华， 强如财宝众多，烦乱不安。
PROV|15|17|有爱，吃素菜， 强如相恨，吃肥牛。
PROV|15|18|暴怒的人挑启争端； 忍怒的人止息纷争。
PROV|15|19|懒惰人的道像荆棘的篱笆； 正直人的路是平坦大道。
PROV|15|20|智慧之子使父亲喜乐； 愚昧的人藐视母亲。
PROV|15|21|无知的人以愚昧为乐； 聪明的人按正直而行。
PROV|15|22|不先商议，所谋无效； 谋士众多，所谋得成。
PROV|15|23|口善应对，自觉喜乐； 话合其时，何等美好。
PROV|15|24|生命之道使智慧人上升， 使他远离底下的阴间。
PROV|15|25|耶和华必拆毁骄傲人的家， 却要立定寡妇的地界。
PROV|15|26|恶谋为耶和华所憎恶； 良言却是纯净的。
PROV|15|27|暴力敛财的，扰害己家； 恨恶贿赂的，必得存活。
PROV|15|28|义人的心思量应答； 恶人的口吐出恶言。
PROV|15|29|耶和华远离恶人， 却听义人的祈祷。
PROV|15|30|眼睛发光，使心喜乐； 好的信息，滋润骨头。
PROV|15|31|耳听使人得生命的责备， 必居住在智慧人之中。
PROV|15|32|弃绝管教的，轻看自己的生命； 领受责备的，却得智慧的心。
PROV|15|33|敬畏耶和华是智慧的训诲； 要得尊荣，先有谦卑。
PROV|16|1|心中的筹谋在乎人， 舌头的应对出于耶和华。
PROV|16|2|人一切所行的，在自己眼中看为纯洁， 惟有耶和华衡量人的内心。
PROV|16|3|你所做的，要交托耶和华， 你所谋的，就必坚立。
PROV|16|4|耶和华造万物各适其用， 就是恶人也为祸患的日子所造。
PROV|16|5|凡心里骄傲的，为耶和华所憎恶； 击掌保证，他难免受罚。
PROV|16|6|因慈爱和信实，罪孽得赎； 敬畏耶和华的，远离恶事。
PROV|16|7|人所行的若蒙耶和华喜悦， 耶和华也使仇敌与他和好。
PROV|16|8|少获利，行事公义， 强如多获利，行事不义。
PROV|16|9|人心筹算自己的道路； 惟耶和华指引他的脚步。
PROV|16|10|王的嘴唇有圣言， 审判之时，他的口必不差错。
PROV|16|11|公道的秤和天平属耶和华， 囊中一切的法码是他所定。
PROV|16|12|作恶，为王所憎恶， 因国位是靠公义坚立。
PROV|16|13|公义的嘴唇，王喜悦， 说正直话的，他喜爱。
PROV|16|14|王的震怒是死亡的使者， 但智慧人能平息王怒。
PROV|16|15|王脸上的光使人有生命， 他的恩惠好像云带来的春雨。
PROV|16|16|得智慧胜过得金子， 选聪明强如选银子。
PROV|16|17|正直人的道远离恶事， 谨守己路的，保全性命。
PROV|16|18|骄傲在败坏以先， 内心高傲在跌倒之前。
PROV|16|19|心里谦卑与困苦人来往， 强如与骄傲人同分战利品。
PROV|16|20|留心训言的 ，必得福乐； 倚靠耶和华的，这人有福。
PROV|16|21|心中有智慧的，必称为聪明人； 嘴唇的甜言，增长人的学问。
PROV|16|22|人有智慧就有生命的泉源； 愚妄人必受愚妄的惩戒。
PROV|16|23|智慧人的心使他的口谨慎， 又使他的嘴唇增长学问。
PROV|16|24|良言如同蜂巢， 使心甘甜，使骨得医治。
PROV|16|25|有一条路，人以为正， 至终却成为死亡之路。
PROV|16|26|劳力的人为自己劳力， 因为他的口腹催逼他。
PROV|16|27|匪徒图谋奸恶， 嘴唇上的言语仿佛烧焦的火。
PROV|16|28|乖谬的人散播纷争， 造谣的离间密友。
PROV|16|29|残暴的人引诱邻舍， 领他走不好的道路。
PROV|16|30|紧闭双目的，图谋乖谬； 紧咬嘴唇的，成就恶事。
PROV|16|31|白发是荣耀的冠冕， 行在公义道上的，必能得着。
PROV|16|32|不轻易发怒的，胜过勇士； 控制自己脾气的，强如取城。
PROV|16|33|人虽可掷签在膝上， 定事却由耶和华。
PROV|17|1|一块干饼，大家相安； 胜过宴席满屋，大家相争。
PROV|17|2|明智的仆人必管辖蒙羞的儿子， 并在兄弟中同分产业。
PROV|17|3|鼎为炼银，炉为炼金， 惟有耶和华熬炼人心。
PROV|17|4|行恶的，留心听恶毒的嘴唇； 说谎的，侧耳听邪恶的舌头。
PROV|17|5|讥笑穷乏人的，是蔑视造他的主； 幸灾乐祸的，难免受罚。
PROV|17|6|子孙为老人的冠冕； 父母是儿女的荣耀。
PROV|17|7|愚顽人说美言并不相宜， 君子说谎言也不合宜。
PROV|17|8|贿赂在馈赠者的眼中看为玉石， 随处运转都得顺利。
PROV|17|9|包容过错的，寻求友爱； 喋喋不休的，离间密友。
PROV|17|10|一句责备的话深入聪明人的心， 强如打愚昧人一百下。
PROV|17|11|恶人只寻求背叛， 残忍的使者必奉差攻击他。
PROV|17|12|宁可遇见失丧小熊的母熊， 也不愿遇见正行愚昧的愚昧人。
PROV|17|13|以恶报善的， 祸患必不离他的家。
PROV|17|14|纷争掀起，如同缺口的水； 因此，争端尚未爆发就当制止。
PROV|17|15|定恶人为义的，定义人为有罪的， 都为耶和华所憎恶。
PROV|17|16|愚昧人既无知， 为何手拿银钱去买智慧呢？
PROV|17|17|朋友时常亲爱， 弟兄为患难而生。
PROV|17|18|在邻舍面前击掌担保的， 是无知的人。
PROV|17|19|喜爱争吵的，是喜爱过犯； 门盖得高的，自取败坏。
PROV|17|20|心中歪曲的，得不着福乐； 舌头颠倒是非的，陷在祸患中。
PROV|17|21|生愚昧之子的，自己必愁苦； 愚顽人的父亲毫无喜乐。
PROV|17|22|喜乐的心能治好疾病； 忧伤的灵使骨头枯干。
PROV|17|23|恶人暗中受贿赂， 以致弯曲公正的路。
PROV|17|24|聪明人面前有智慧； 愚昧人眼望地的尽头。
PROV|17|25|愚昧的儿子使父亲愁烦， 使那生他的母亲忧苦。
PROV|17|26|刑罚义人实为不善， 责打正直的君子也不宜。
PROV|17|27|节制言语的，有见识； 性情温良的人，有聪明。
PROV|17|28|愚妄人若静默不言，可算为智慧， 闭上嘴唇也可算为聪明。
PROV|18|1|孤僻的人只顾自己的心愿 ， 他鄙视一切健全的知识。
PROV|18|2|愚昧人不喜爱聪明， 只喜爱表达自己的心意。
PROV|18|3|邪恶来，藐视跟着来； 羞耻到，辱骂同时到。
PROV|18|4|人的口所讲的话如同深水， 智慧之泉如涌流的河水。
PROV|18|5|偏袒恶人的情面，是不好的。 审判时使义人受屈，也是不善。
PROV|18|6|愚昧人的嘴唇挑起争端， 一开口就招鞭打。
PROV|18|7|愚昧人的口自取败坏， 他的嘴唇是自己生命的圈套。
PROV|18|8|造谣者的话如同美食， 深入人的肚腹。
PROV|18|9|做工懈怠的， 是破坏者的兄弟。
PROV|18|10|耶和华的名是坚固台， 义人奔入就得安稳。
PROV|18|11|有钱人的财物是他坚固的城， 在他幻想中，犹如高墙。
PROV|18|12|败坏之先，人心骄傲； 要得尊荣，先有谦卑。
PROV|18|13|未听完就回话的， 就是他的愚昧和羞辱。
PROV|18|14|人的心灵忍耐疾病； 心灵忧伤，谁能承当呢？
PROV|18|15|聪明人的心得知识； 智慧人的耳求知识。
PROV|18|16|人的礼物为他开路， 引他到高位的人面前。
PROV|18|17|先诉情由的，似乎有理； 另一人来到，就察出实情。
PROV|18|18|掣签能止息纷争， 也能化解双方激烈的争辩。
PROV|18|19|被冒犯的弟兄 强如难以攻下的坚城； 纷争如同城堡的门闩。
PROV|18|20|人的肚腹必因口所结的果实饱足； 他必因嘴唇所出的感到满足。
PROV|18|21|生死在舌头的掌握之下， 喜爱弄舌的，必吃它所结的果实。
PROV|18|22|得着妻子的，得着好处， 他是蒙了耶和华的恩惠。
PROV|18|23|穷乏人说哀求的话； 有钱人却用威吓的话回答。
PROV|18|24|朋友太多的人，必受损害 ； 但有一知己比兄弟更亲密。
PROV|19|1|行为纯正的穷乏人 胜过嘴唇歪曲的愚昧人。
PROV|19|2|热心而无见识，实为不善； 脚步急快的，易入歧途。
PROV|19|3|人因愚昧自毁前途， 他的心却埋怨耶和华。
PROV|19|4|财富使朋友增多； 贫寒人连仅有的朋友也离弃他。
PROV|19|5|作假见证的，难免受罚； 口吐谎言的，不能逃脱。
PROV|19|6|有权贵的，许多人求他赏脸； 爱送礼的，人都作他的朋友。
PROV|19|7|穷乏人连兄弟都恨他， 何况朋友，更是远离他！ 他用言语追随，他们却不在。
PROV|19|8|得着智慧的，爱惜生命； 持守聪明的，寻得好处。
PROV|19|9|作假见证的，难免受罚； 口吐谎言的，必定灭亡。
PROV|19|10|愚昧人奢华度日并不相宜， 仆人管辖王子，也不应该。
PROV|19|11|人有见识就不轻易发怒， 宽恕人的过失便是自己的荣耀。
PROV|19|12|王的愤怒好像狮子吼叫； 他的恩惠却如草上的甘露。
PROV|19|13|愚昧的儿子是父亲的祸患， 妻子的争吵如雨连连滴漏。
PROV|19|14|房屋钱财是祖宗所遗留的； 惟有贤慧的妻是耶和华所赐的。
PROV|19|15|懒惰使人沉睡， 懈怠的人必捱饿。
PROV|19|16|遵守诫命的，保全生命； 轻忽己路的，必致死亡。
PROV|19|17|怜悯贫寒人的，就是借给耶和华， 他的报偿，耶和华必归还他。
PROV|19|18|趁还有指望，管教你的儿子， 不可执意摧毁他。
PROV|19|19|暴怒的人必受惩罚， 你若救他，必须再救。
PROV|19|20|要听劝言，接受训诲， 使你终久有智慧。
PROV|19|21|人心多有计谋； 惟有耶和华的筹算才能成就。
PROV|19|22|仁慈的人令人喜爱 ， 穷乏人强如说谎言的。
PROV|19|23|敬畏耶和华的，得着生命， 他必饱足安居，不遭祸患。
PROV|19|24|懒惰人把手埋入盘里， 连缩回送进口中也不肯。
PROV|19|25|责打傲慢人，能使无知的人变精明； 责备聪明人，他就明白知识。
PROV|19|26|虐待父亲、驱逐母亲的， 是蒙羞致辱之子。
PROV|19|27|我儿啊，停止听 那叫你偏离知识言语的教导 。
PROV|19|28|卑劣的见证嘲笑公平， 恶人的口吞下罪孽。
PROV|19|29|刑罚是为傲慢人预备的， 鞭打则是为愚昧人的背预备的。
PROV|20|1|酒能使人傲慢，烈酒使人喧嚷， 凡沉溺其中的，都无智慧。
PROV|20|2|王的威吓如狮子吼叫， 激怒他的是自害己命。
PROV|20|3|止息纷争是人的尊荣， 愚妄人争闹不休。
PROV|20|4|懒惰人因冬寒不去耕种， 到收割时，他去寻找，一无所得。
PROV|20|5|人心中的筹算如同深水， 惟聪明人才能汲引出来。
PROV|20|6|很多人声称自己忠信， 但诚信的人谁能遇着呢？
PROV|20|7|义人行为纯正， 他后代的子孙有福了！
PROV|20|8|王坐在审判的位上， 以眼目驱散一切邪恶。
PROV|20|9|谁能说：“我已经洁净了我的心， 脱净了我的罪？”
PROV|20|10|两样的法码和两样的伊法 ， 都为耶和华所憎恶。
PROV|20|11|孩童的行动或纯洁，或正直， 都以行为显明自己。
PROV|20|12|能听的耳，能看的眼， 二者都为耶和华所造。
PROV|20|13|不要贪睡，免致贫穷； 眼要睁开，就可吃饱。
PROV|20|14|买东西的说：“不好，不好！” 及至离去，他却自夸。
PROV|20|15|有金子和许多宝石， 惟知识的嘴唇是贵重的珍宝。
PROV|20|16|谁为陌生人担保，就拿谁的衣服； 谁为外邦人作保，谁就要承当。
PROV|20|17|靠谎言而得的食物，令人愉悦； 到后来，他的口必充满碎石。
PROV|20|18|计谋凭筹算立定， 打仗要凭智谋。
PROV|20|19|到处传话的，泄漏机密； 口无遮拦的，不可与他结交。
PROV|20|20|咒骂父母的， 他的灯必熄灭，在漆黑中。
PROV|20|21|起初很快得来的产业， 终久却不是福。
PROV|20|22|你不要说：“我要以恶报恶”； 要等候耶和华，他必拯救你。
PROV|20|23|两样的法码为耶和华所憎恶， 诡诈的天平也为不善。
PROV|20|24|人的脚步为耶和华所定， 人岂能明白自己的道路呢？
PROV|20|25|人冒失地声称：“这是神圣的！” 许愿之后才细想，就是自陷圈套。
PROV|20|26|智慧的王驱散恶人， 用轮子滚过他们。
PROV|20|27|人的灵是耶和华的灯， 鉴察人的内心深处。
PROV|20|28|慈爱和诚实庇护君王， 他的王位因慈爱而立稳。
PROV|20|29|强壮是青年的荣耀； 白发为老人的尊荣。
PROV|20|30|鞭伤除净邪恶， 责打可洁净人心深处。
PROV|21|1|王的心在耶和华手中像河水， 他能使它随意流转。
PROV|21|2|人一切所行的，在自己眼中看为正直， 惟有耶和华衡量人心。
PROV|21|3|行公义和公平 比献祭更蒙耶和华悦纳。
PROV|21|4|眼高心傲，就是恶人的灯， 都是罪。
PROV|21|5|殷勤筹划的，足致丰裕； 行事急躁的，必致缺乏。
PROV|21|6|用诡诈之舌所得的财富 如被吹散的雾气，趋向灭亡 。
PROV|21|7|恶人的残暴必扫去自己， 因他们不肯按公平行事。
PROV|21|8|有罪的人其路弯曲； 纯洁的人行为正直。
PROV|21|9|宁可住在房顶的一角， 也不与好争吵的妇人同住。
PROV|21|10|恶人的心渴想邪恶， 他的眼并不怜悯邻舍。
PROV|21|11|傲慢人受惩罚，愚蒙人可得智慧； 智慧人受训诲，便得知识。
PROV|21|12|公义的上帝 鉴察恶人的家， 他倾覆恶人，以致灭亡。
PROV|21|13|塞耳不听贫寒人哀求的， 他自己呼求，也不蒙应允。
PROV|21|14|暗中送的礼物挽回怒气， 怀里的贿赂能止息暴怒。
PROV|21|15|秉公行义使义人喜乐， 却使作恶的人败坏。
PROV|21|16|人偏离智慧的路， 必与阴魂为伍 。
PROV|21|17|爱宴乐的，必致穷乏； 贪爱酒和油的，必不富足。
PROV|21|18|恶人作义人的赎价， 奸诈人代替正直人。
PROV|21|19|宁可住在旷野之地， 也不与争吵易怒的妇人同住。
PROV|21|20|智慧人的居所积蓄宝物与膏油 ； 愚昧人却挥霍一空。
PROV|21|21|追求公义慈爱的， 就寻得生命、公义 和尊荣。
PROV|21|22|智慧人爬上勇士的城墙， 摧毁他所倚靠的堡垒。
PROV|21|23|谨守口和舌的， 就保护自己免受灾难。
PROV|21|24|心骄气傲的人名叫傲慢， 他行事出于狂妄骄傲。
PROV|21|25|懒惰人的欲望害死自己， 因为他的手不肯做工；
PROV|21|26|有人终日贪得无餍， 义人却施舍而不吝惜。
PROV|21|27|恶人献的祭是可憎的， 何况他存恶意来献呢？
PROV|21|28|不实的见证必消灭； 惟聆听真情的，他的证词有力。
PROV|21|29|恶人脸无羞耻； 正直人行事坚定 。
PROV|21|30|没有人能以智慧、聪明、 谋略抵挡耶和华。
PROV|21|31|马是为打仗之日预备的； 得胜却在于耶和华。
PROV|22|1|美名胜过大财， 宏恩强如金银。
PROV|22|2|有钱人与穷乏人相遇 ， 他们都为耶和华所造。
PROV|22|3|通达人见祸就藏躲； 愚蒙人却前往受害。
PROV|22|4|敬畏耶和华心存谦卑， 就得财富、尊荣、生命为赏赐。
PROV|22|5|歪曲的人路上有荆棘和罗网， 保护自己生命的，必要远离。
PROV|22|6|教养孩童走当行的道， 就是到老他也不偏离。
PROV|22|7|有钱人管辖穷乏人， 欠债的是债主的仆人。
PROV|22|8|撒不义种子的必收割灾祸， 他逞怒的杖也必废掉。
PROV|22|9|眼目仁慈的必蒙福， 因他将食物分给贫寒人。
PROV|22|10|赶出傲慢人，争端就消除， 纷争和羞辱也必止息。
PROV|22|11|喜爱清心，嘴唇有恩言的， 王必与他为友。
PROV|22|12|耶和华的眼目保护知识， 却毁坏奸诈人的言语。
PROV|22|13|懒惰人说：“外面有狮子， 我在街上必被杀害。”
PROV|22|14|陌生女子的口是深坑， 耶和华所憎恶的，必陷在其中。
PROV|22|15|愚昧迷住孩童的心， 用管教的杖可以远远赶除。
PROV|22|16|欺压贫寒人为要利己的， 并送礼给有钱人的，都必缺乏。
PROV|22|17|你要侧耳听智慧人的言语 ， 留心领会我的知识。
PROV|22|18|你若心中存记， 嘴唇也准备就绪，这是美的。
PROV|22|19|我今日特地指教你， 为要使你倚靠耶和华。
PROV|22|20|谋略和知识的美事 ， 我岂没有写给你吗？
PROV|22|21|要使你明白真情实理， 好将实情回覆那差你来的人。
PROV|22|22|不可因人贫寒就抢夺他， 也不可在城门口欺压困苦人，
PROV|22|23|因耶和华必为他们辩护， 也必夺取那抢夺者的命。
PROV|22|24|不可结交好生气的人， 也不可与暴怒的人来往，
PROV|22|25|恐怕你效法他的行为， 自己就陷在圈套里。
PROV|22|26|不要为人击掌担保， 也不要为债务作保。
PROV|22|27|你若没有什么可偿还， 何必使人夺去你睡卧的床呢？
PROV|22|28|祖先所立的地界， 你不可挪移。
PROV|22|29|你看见办事殷勤的人吗？ 他必侍立在君王面前， 不在平庸的人面前。
PROV|23|1|你若与长官坐席， 要留意在你面前的是谁。
PROV|23|2|你若是胃口大的人， 就当拿刀放在喉咙上。
PROV|23|3|不可贪恋长官的美食， 因为那是欺哄人的食物。
PROV|23|4|不要劳碌求富， 要有聪明来节制。
PROV|23|5|你定睛在财富，它就消失， 因为它必长翅膀，如鹰向天飞去。
PROV|23|6|守财奴 的饭，你不要吃， 也不要贪恋他的美味；
PROV|23|7|因为他的心怎样算计 ， 他为人就是这样。 他虽对你说：请吃，请喝， 他的心却与你相背。
PROV|23|8|你所吃的那点食物必吐出来， 你恭维的话语也必落空。
PROV|23|9|不要说话给愚昧人听， 因他必藐视你智慧的言语。
PROV|23|10|不可挪移古时的地界， 也不可侵占孤儿的田地，
PROV|23|11|因他们的救赎者 大有能力， 他必向你为他们辩护。
PROV|23|12|你要留心领受训诲， 侧耳听从知识的言语。
PROV|23|13|不可不管教孩童， 因为你用杖打他，他不会死。
PROV|23|14|你用杖打他， 就可以救他的性命免下阴间。
PROV|23|15|我儿啊，你若心存智慧， 我的心就甚欢喜。
PROV|23|16|你的嘴唇若说正直话， 我的心肠也必快乐。
PROV|23|17|你的心不要羡慕罪人， 却要羡慕常常敬畏耶和华的人，
PROV|23|18|因为你必有前途， 你的指望也不致断绝。
PROV|23|19|我儿啊，你当听，当存智慧， 好在正道上引导你的心。
PROV|23|20|不可与好饮酒的人在一起， 也不要跟贪吃肉的人来往，
PROV|23|21|因为贪食好酒的，必致贫穷， 爱睡觉的，必穿破烂衣服。
PROV|23|22|你要听从生你的父亲； 不可因母亲年老而轻看她。
PROV|23|23|你当获得真理，不可出卖， 智慧、训诲和聪明也是一样。
PROV|23|24|义人的父亲必大大快乐， 生智慧儿子的，必因他欢喜。
PROV|23|25|愿你的父母欢喜， 愿那生你的母亲快乐。
PROV|23|26|我儿啊，要将你的心归我， 你的眼目也要喜爱 我的道路。
PROV|23|27|妓女是深坑， 外邦女子是窄井。
PROV|23|28|她像强盗埋伏， 她使奸诈的人增多。
PROV|23|29|谁有祸患？谁有灾难？ 谁有纷争？谁有焦虑？ 谁无故受伤？谁的眼目红赤？
PROV|23|30|就是那流连饮酒的人， 常去寻找调和的酒。
PROV|23|31|酒发红，在杯中闪烁时， 你不可观看； 虽下咽舒畅， 终究它必咬你如蛇，刺你如毒蛇。
PROV|23|32|
PROV|23|33|你的眼睛必看见怪异的事， 你的心必发出乖谬的话。
PROV|23|34|你必像躺在深海中， 或卧在桅杆顶上，
PROV|23|35|说：“人击打我，但我未受伤， 重击我，我不觉得。 我几时清醒， 还要再去寻酒。”
PROV|24|1|你不要嫉妒恶人， 也不要渴望与他们相处，
PROV|24|2|因为他们的心图谋暴行， 他们的嘴唇谈论奸恶。
PROV|24|3|房屋因智慧建造， 因聪明立稳；
PROV|24|4|又因知识， 屋内充满各样美好宝贵的财物。
PROV|24|5|有智慧的勇士大有能力， 有知识的人力上加力。
PROV|24|6|你去打仗，要凭智谋； 谋士众多，就必得胜。
PROV|24|7|对愚妄人，智慧高不可及， 所以他在城门不敢开口。
PROV|24|8|图谋行恶的， 必称为奸诈人。
PROV|24|9|愚妄人的筹划尽是罪恶， 傲慢者为人所憎恶。
PROV|24|10|在患难时你若灰心， 你的力量就微小。
PROV|24|11|人被拉到死亡，你要解救； 人将被杀，你须拦阻。
PROV|24|12|你若说：“看哪，这事我们不知道”， 那衡量人心的岂不明白吗？ 保护你性命的岂不知道吗？ 他岂不按各人所做的报应各人吗？
PROV|24|13|我儿啊，你要吃蜜，因为它是美好的， 要让甘甜的蜜滴入你的口。
PROV|24|14|你要知道，智慧对你的生命正像如此。 你若找着，必有前途， 你的指望也不致断绝。
PROV|24|15|你这恶人，不可埋伏攻击义人的家， 也不可毁坏他安居之所。
PROV|24|16|因为义人虽七次跌倒，仍必兴起； 恶人却被祸患倾倒。
PROV|24|17|你的仇敌跌倒，你不要欢喜， 他倾倒，你的心不要快乐；
PROV|24|18|恐怕耶和华看见就不喜悦， 将怒气从仇敌身上转过来。
PROV|24|19|不要为作恶的心怀不平， 也不要嫉妒恶人，
PROV|24|20|因为坏人没有前途， 恶人的灯也必熄灭。
PROV|24|21|我儿啊，你要敬畏耶和华与君王， 不可结交反覆无常的人，
PROV|24|22|因为他们的灾难必忽然兴起。 谁能知道耶和华与君王所施行的毁灭呢？
PROV|24|23|以下也是智慧人的箴言： 审判时看人情面是不好的。
PROV|24|24|对恶人说“你是义人”的， 万民必诅咒，万族必恼恨。
PROV|24|25|责备恶人的，必得喜悦， 美好的福分也必临到他。
PROV|24|26|应对合宜的， 犹如与人亲吻。
PROV|24|27|你要在外面预备材料， 在田间为自己准备齐全， 然后才建造你的房屋。
PROV|24|28|不可无故作证反对邻舍， 也不可用嘴唇欺骗人。
PROV|24|29|不可说：“人怎样待我，我也怎样待他， 我必照他所做的报复他。”
PROV|24|30|我经过懒惰人的田地， 走过无知人的葡萄园，
PROV|24|31|看哪，它长满了荆棘， 荨麻盖地面， 石墙也坍塌了。
PROV|24|32|我看见就留心思想， 我看着就领受训诲。
PROV|24|33|再睡片时，打盹片时， 抱着双臂躺卧片时，
PROV|24|34|你的贫穷就如盗贼来到， 你的贫乏仿佛拿盾牌的人来临。
PROV|25|1|以下也是 所罗门 的箴言，是 犹大 王 希西家 的人所誊录的。
PROV|25|2|隐藏事情是上帝的荣耀； 查明事情乃君王的荣耀。
PROV|25|3|天之高，地之深， 君王之心测不透。
PROV|25|4|除去银子的渣滓， 银匠就做出器皿来。
PROV|25|5|除去王面前的恶人， 国位就靠公义坚立。
PROV|25|6|不可在君王面前妄自尊大， 也不要站在大人的位上。
PROV|25|7|宁可让人家说“请你上到这里来”， 强如在你觐见的贵人面前令你退下。
PROV|25|8|不要冒失出去与人争讼 ， 免得你的邻舍羞辱你， 最后你就不知怎么做。
PROV|25|9|要与邻舍争辩你的案情， 不可泄漏他人的隐密，
PROV|25|10|恐怕听见的人责骂你， 你就难以摆脱臭名。
PROV|25|11|一句话说得合宜， 就如金苹果在银网子里
PROV|25|12|智慧人的劝戒在顺从的人耳中， 好像金环和金首饰。
PROV|25|13|忠信的使者对那差他的人， 就如收割时有冰雪的凉气， 使主人的心舒畅。
PROV|25|14|人空夸礼物而不肯赠送， 就好像有风有云却无雨。
PROV|25|15|恒常的忍耐可以劝服君王， 柔和的舌头能折断骨头。
PROV|25|16|你得了蜜，吃够就好， 免得过饱就吐出来。
PROV|25|17|你的脚要少进邻舍的家， 免得他厌烦你，恨恶你。
PROV|25|18|作假见证陷害邻舍的， 就是大锤，是利刀，是快箭。
PROV|25|19|患难时倚靠奸诈的人， 好像牙齿断裂，又如脚脱臼。
PROV|25|20|对伤心的人唱歌， 就如冷天脱他的衣服， 又如在碱上倒醋 。
PROV|25|21|你的仇敌若饿了，就给他饭吃， 若渴了，就给他水喝；
PROV|25|22|因为你这样做，就是把炭火堆在他的头上， 耶和华必回报你。
PROV|25|23|正如北风生雨， 毁谤的舌头也生怒容。
PROV|25|24|宁可住在房顶的一角， 也不与好争吵的妇人同住。
PROV|25|25|有好消息从遥远的地方来， 就如凉水滋润口渴的人。
PROV|25|26|义人在恶人面前退缩， 好像搅浑之泉，污染之井。
PROV|25|27|吃蜜过多是不好的， 自求荣耀也是一样。
PROV|25|28|人不克制自己的心， 就像毁坏的城没有墙。
PROV|26|1|愚昧人得尊荣不相宜， 正如夏天落雪，收割时下雨。
PROV|26|2|诅咒不会无故临到 ， 正如麻雀掠过，燕子翻飞。
PROV|26|3|鞭子是为打马，辔头是为勒驴， 刑杖正是为打愚昧人的背。
PROV|26|4|不要照愚昧人的愚昧话回答他， 免得你与他一样。
PROV|26|5|要照愚昧人的愚昧话回答他， 免得他自以为有智慧。
PROV|26|6|藉愚昧人的手寄信的， 就像砍断双脚，喝下残暴。
PROV|26|7|箴言在愚昧人的口中， 正如瘸子的脚悬空无用。
PROV|26|8|将尊荣给愚昧人的， 就像石头绑在弹弓上。
PROV|26|9|箴言在愚昧人的口中， 好像荆棘刺入醉汉的手。
PROV|26|10|雇愚昧人的，与雇过路人的， 就像弓箭手射伤任何人。
PROV|26|11|愚昧人重复做愚昧之事， 就如狗转过来吃自己所吐的。
PROV|26|12|你看见自以为有智慧的人吗？ 愚昧人比他更有指望。
PROV|26|13|懒惰人说：“道路有猛狮， 街上有壮狮。”
PROV|26|14|懒惰人在床上， 就像门在轴心上转动一样。
PROV|26|15|懒惰人把手埋入盘里， 就是送进口中也觉得累。
PROV|26|16|懒惰人眼看自己 比七个善于应对的人更有智慧。
PROV|26|17|过路时卷入与己无关的纷争， 好像人揪住狗耳一般。
PROV|26|18|人欺骗邻舍，却说 “我只是开玩笑而已”， 他就像疯狂的人抛掷致死的火把和利箭。
PROV|26|19|
PROV|26|20|火缺了柴就必熄灭； 无人造谣，纷争就止息。
PROV|26|21|好争吵的人煽动争端， 就如余火加炭，火上加柴一样。
PROV|26|22|造谣者的话如同美食， 深入人的肚腹。
PROV|26|23|火热的 嘴唇，邪恶的心， 好像银渣包在瓦器上。
PROV|26|24|仇敌用嘴唇掩饰， 心里却藏着诡诈；
PROV|26|25|他用甜言蜜语，你不能相信他， 因为他心中有七样可憎恶的事。
PROV|26|26|他虽用诡诈掩饰怨恨， 他的邪恶必在集会中显露。
PROV|26|27|挖陷坑的，自己必陷在其中； 滚石头的，石头反滚在他身上。
PROV|26|28|虚谎的舌憎恨他所压伤的人； 谄媚的口败坏人的事。
PROV|27|1|不要为明天自夸， 因为你不知道每天会发生何事。
PROV|27|2|要让陌生人夸奖你，不可用口自夸； 让外邦人称赞你，不可用嘴唇称赞自己。
PROV|27|3|石头沉，沙土重， 愚妄人的恼怒比这两样更沉重。
PROV|27|4|愤怒为残忍，怒气像狂澜， 惟有嫉妒，谁能挡得住呢？
PROV|27|5|当面的责备 胜过隐藏的爱情。
PROV|27|6|朋友加的伤痕出于忠诚； 敌人的亲吻却是多余。
PROV|27|7|人吃饱了，厌恶蜂房的蜜； 人饥饿了，一切苦物都觉甘甜。
PROV|27|8|人离故乡漂泊， 就像雀鸟离窝四处飞翔。
PROV|27|9|膏油与香料使人心喜悦， 朋友诚心的劝勉也是如此甘美。
PROV|27|10|你的朋友和父亲的朋友， 你都不可离弃。 你遭难时，不要上兄弟的家去； 相近的邻舍强如远方的兄弟。
PROV|27|11|我儿啊，你要做智慧人，好叫我的心欢喜， 使我可以回答那辱骂我的人。
PROV|27|12|通达人见祸就藏躲； 愚蒙人却前往受害。
PROV|27|13|谁为陌生人担保，就拿谁的衣服； 谁为外邦女子作保，谁就要承当。
PROV|27|14|清晨起来大声给朋友祝福的， 就算是诅咒他。
PROV|27|15|下雨天连连滴漏， 好争吵的妇人就像这样；
PROV|27|16|拦阻她的，就是拦阻风， 又像用右手抓油。
PROV|27|17|以铁磨铁，越磨越利， 朋友当面琢磨，也是如此。
PROV|27|18|看守无花果树的，必吃树上的果子； 敬奉主人的，必得尊荣。
PROV|27|19|水中照脸，彼此相符； 人心相映，也是如此。
PROV|27|20|阴间和冥府 永不满足， 人的眼目也是如此。
PROV|27|21|鼎为炼银，炉为炼金， 口中的称赞也试炼人。
PROV|27|22|用杵把愚妄人与谷粒一同捣在臼中， 他的愚昧还是离不了他。
PROV|27|23|你要详细知道你羊群的景况， 留心照顾你的牛群，
PROV|27|24|因为财富不能永留， 冠冕岂能存到万代？
PROV|27|25|青草除去，嫩草长出， 山上的菜蔬也被采收。
PROV|27|26|绵羊可以做衣服， 公山羊可作田地的价值，
PROV|27|27|并有母山羊奶够你吃， 够你养家和女仆的生活。
PROV|28|1|恶人虽无人追赶也逃跑； 义人却胆壮像狮子。
PROV|28|2|地上因有罪过，君王就多更换； 因聪明和有见识的人，国必长存。
PROV|28|3|穷乏人欺压贫寒人， 好像暴雨扫过，不留粮食。
PROV|28|4|离弃律法的，夸奖恶人； 遵守律法的，却与恶人相争。
PROV|28|5|恶人不明白公义； 惟有寻求耶和华的，无不明白。
PROV|28|6|行为纯正的穷乏人 胜过行事歪曲的有钱人。
PROV|28|7|谨守教诲的，是聪明之子； 与贪食者为伍的，却羞辱其父。
PROV|28|8|人以厚利增加财富， 是给那怜悯贫寒人的积财。
PROV|28|9|转耳不听教诲的， 他的祈祷也可憎。
PROV|28|10|诱惑正直人行恶道的，必掉在自己的坑里； 惟有完全人必承受福分。
PROV|28|11|有钱人自以为有智慧， 但聪明的贫寒人能看穿他。
PROV|28|12|义人高升，有大荣耀； 恶人兴起，人就躲藏。
PROV|28|13|遮掩自己过犯的，必不顺利； 承认且离弃过犯的，必蒙怜悯。
PROV|28|14|常存敬畏的，这人有福了； 心里刚硬的，必陷在祸患里。
PROV|28|15|邪恶的君王压制贫民， 好像吼叫的狮子，又如觅食的熊。
PROV|28|16|无知的君王多行暴虐； 恨恶非分之财的，必年长日久。
PROV|28|17|背负流人血之罪的，必逃跑直到地府； 愿无人帮助他！
PROV|28|18|行为正直的，必蒙拯救； 行事弯曲的，立时跌倒。
PROV|28|19|耕种自己田地的，粮食充足； 追求虚浮的，穷困潦倒。
PROV|28|20|诚实人必多得福； 想要急速发财的，难免受罚。
PROV|28|21|看人情面是不好的； 却有人因一块饼而犯法。
PROV|28|22|守财奴 想要急速发财， 却不知穷乏必临到他身上。
PROV|28|23|责备人的，后来蒙人喜悦， 多于那用舌头谄媚人的。
PROV|28|24|抢夺父母竟说“这不是罪过”， 此人与毁灭者同类。
PROV|28|25|心中贪婪的，挑起争端； 倚靠耶和华的，必得丰裕。
PROV|28|26|心中自以为是的，就是愚昧人； 凭智慧行事的，必蒙拯救。
PROV|28|27|赒济穷乏人的，不致缺乏； 遮眼不看的，多受诅咒。
PROV|28|28|恶人兴起，人就躲藏； 恶人败亡，义人必增多。
PROV|29|1|人屡次受责罚，仍然硬着颈项， 他必顷刻被毁，无从医治。
PROV|29|2|义人增多，民就喜乐； 恶人掌权，民就叹息。
PROV|29|3|爱慕智慧的，使父亲喜乐； 结交妓女的，却浪费钱财。
PROV|29|4|王藉公平，使国坚定； 强索贡物的，使它毁坏。
PROV|29|5|谄媚邻舍的， 就是设网罗绊他的脚。
PROV|29|6|恶人犯罪，自陷圈套； 惟独义人欢呼喜乐。
PROV|29|7|义人关注贫寒人的案情； 恶人不明了这种知识。
PROV|29|8|傲慢人煽动全城； 智慧人止息众怒。
PROV|29|9|智慧人与愚妄人有争讼， 或怒或笑，总不得安宁。
PROV|29|10|好流人血的，恨恶完全人， 正直人却顾惜 他的性命。
PROV|29|11|愚昧人怒气全发； 智慧人自我平息。
PROV|29|12|君王若听谎言， 他一切臣仆都是奸恶。
PROV|29|13|穷乏人和欺压者相遇 ， 耶和华使他们的眼目明亮。
PROV|29|14|君王凭诚信判断贫寒人， 他的国位必永远坚立。
PROV|29|15|杖打和责备能增加智慧； 任性的少年使母亲羞愧。
PROV|29|16|恶人多，过犯也加多， 义人必看见他们败亡。
PROV|29|17|管教你的儿子，他就使你得安宁， 也使你心里喜乐。
PROV|29|18|没有异象 ，民就放肆； 惟遵守律法的，便为有福。
PROV|29|19|仆人不能靠言语受教； 他即使明白，也不回应。
PROV|29|20|你见过言语急躁的人吗？ 愚昧人比他更有指望。
PROV|29|21|人将仆人从小娇养， 至终必带来忧伤 。
PROV|29|22|好生气的人挑起争端， 暴怒的人多多犯错。
PROV|29|23|人的高傲使自己蒙羞； 心里谦逊的，必得尊荣。
PROV|29|24|与盗贼分赃的，是恨恶自己的性命； 他虽听见发誓的声音，也不告诉人。
PROV|29|25|惧怕人的，陷入圈套； 惟有倚靠耶和华的，必得安稳。
PROV|29|26|求王恩的人多； 人获公正来自耶和华。
PROV|29|27|不义之人，义人憎恶； 行事正直的，恶人憎恶。
PROV|30|1|雅基 的儿子、 玛撒 人 亚古珥 的言语 ，是这人对 以铁 和 乌甲 说的。
PROV|30|2|我比众人更像畜牲， 也没有人的聪明。
PROV|30|3|我没有学好智慧， 也不认识至圣者。
PROV|30|4|谁升天又降下来？ 谁聚风在手掌中？ 谁包水在衣服里？ 谁立定地的四极？ 他名叫什么？ 他儿子名叫什么？ 你知道吗？
PROV|30|5|上帝的言语句句都是炼净的， 投靠他的，他便作他们的盾牌。
PROV|30|6|你不可加添他的言语， 恐怕他责备你，你就显为说谎的。
PROV|30|7|我求你两件事， 在我未死之先，不要拒绝我：
PROV|30|8|求你使虚假和谎言远离我， 使我不贫穷也不富足， 赐给我需用的饮食。
PROV|30|9|免得我饱足了，就不认你，说： “耶和华是谁呢？” 又恐怕我贫穷就偷窃， 以致亵渎我上帝的名。
PROV|30|10|不要向主人谗害他的仆人， 恐怕他诅咒你，你便算为有罪。
PROV|30|11|有一类人，诅咒父亲， 不给母亲祝福。
PROV|30|12|有一类人，自以为纯洁， 却没有洗净自己的污秽。
PROV|30|13|有一类人，眼目何其高傲， 眼皮也是高举。
PROV|30|14|有一类人，牙如剑，齿如刀， 要吞灭地上的困苦人和世间的贫穷人。
PROV|30|15|水蛭有两个女儿： “给呀，给呀。” 有三样不知足的， 不说“够了”的有四样：
PROV|30|16|阴间和不生育的子宫， 吸水不足的地，还有不说“够了”的火。
PROV|30|17|嘲笑父亲、藐视而不听从母亲的， 谷中的乌鸦必啄他的眼睛，小鹰也必吃它。
PROV|30|18|我所测不透的奇妙有三样， 我所不知道的有四样：
PROV|30|19|就是鹰在空中飞的道， 蛇在磐石上爬的道， 船在海中行的道， 男与女交合的道。
PROV|30|20|淫妇的道是这样， 她吃了，把嘴一擦就说： “我没有行恶。”
PROV|30|21|使地震动的有三样， 地承担不起的有四样：
PROV|30|22|就是仆人作王， 愚顽人吃得饱足，
PROV|30|23|令人憎恶的女子出嫁， 婢女取代她的女主人。
PROV|30|24|地上有四样东西虽小，却甚聪明：
PROV|30|25|蚂蚁是无力之类， 却在夏天预备粮食。
PROV|30|26|石獾并非强壮之类， 却在岩石中造房子。
PROV|30|27|蝗虫没有君王， 却分队而出。
PROV|30|28|壁虎你用手就可抓住， 它却住在王宫。
PROV|30|29|脚步威武的有三样， 行走威武的有四样：
PROV|30|30|狮子－百兽中最勇猛的、 无论遇见什么绝不退缩，
PROV|30|31|猎狗，公山羊， 和有整排士兵的君王。
PROV|30|32|你若行事愚顽，自高自傲， 或是设计恶谋，就当用手捂口。
PROV|30|33|搅动牛奶必成乳酪， 扭鼻子必出血， 照样，激发烈怒必挑起争端。
PROV|31|1|玛撒 王 利慕伊勒 的言语，就是他母亲教导他的 。
PROV|31|2|我儿，怎么了？ 我腹中生的儿，怎么了？ 我许愿而得的儿，怎么了？
PROV|31|3|不要将你的精力给妇女， 也不要有败坏君王的行为。
PROV|31|4|利慕伊勒 啊，君王不宜，君王不宜喝酒， 王子寻找烈酒也不相宜；
PROV|31|5|恐怕喝了就忘记所颁的法令， 颠倒所有困苦人的是非。
PROV|31|6|可以把烈酒给将亡的人喝， 把酒给心里愁苦的人喝，
PROV|31|7|让他喝了，就忘记他的贫穷， 不再记得他的苦楚。
PROV|31|8|你当为不能自辩的人 开口， 为所有孤独无助者伸冤。
PROV|31|9|你当开口按公义判断， 当为困苦和贫穷的人辩护。
PROV|31|10|才德的妇人谁能得着呢？ 她的价值远胜过宝石。
PROV|31|11|她丈夫心里信赖她， 必不缺少利益；
PROV|31|12|她终其一生， 使丈夫有益无损。
PROV|31|13|她寻找羊毛和麻， 欢喜用手做工。
PROV|31|14|她好像商船， 从远方运来粮食，
PROV|31|15|未到黎明她就起来， 把食物分给家中的人， 将当做的工分派女仆。
PROV|31|16|她想得田地，就去买来， 用手中的成果栽葡萄园。
PROV|31|17|她以能力束腰， 使膀臂有力。
PROV|31|18|她觉得自己获利不错， 她的灯终夜不灭。
PROV|31|19|她伸手拿卷线杆， 她的手掌把住纺车。
PROV|31|20|她张手赒济困苦人， 伸手帮助贫穷人。
PROV|31|21|她不因下雪为家里的人担心， 因为全家都穿上朱红衣服。
PROV|31|22|她为自己制作被单， 她的衣服是细麻和紫色布做的。
PROV|31|23|她丈夫在城门口与本地的长老同坐， 为人所认识。
PROV|31|24|她做细麻布衣裳来卖， 又将腰带卖给商家。
PROV|31|25|能力和威仪是她的衣服， 她想到日后的景况就喜笑。
PROV|31|26|她开口就发智慧， 她舌上有仁慈的教诲。
PROV|31|27|她管理家务， 并不吃闲饭。
PROV|31|28|她的儿女起来称她有福， 她的丈夫也称赞她：
PROV|31|29|“才德的女子很多， 惟独你超过一切。”
PROV|31|30|魅力是虚假的，美貌是虚浮的； 惟敬畏耶和华的妇女必得称赞。
PROV|31|31|她手中的成果你们要赏给她， 愿她的工作在城门口荣耀她。
