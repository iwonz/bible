TITUS|1|1|Paulus servus Dei, apostolus autem Iesu Christi secundum fi dem electorum Dei et agnitionem veritatis, quae secundum pietatem est
TITUS|1|2|in spem vitae aeternae, quam promisit, qui non mentitur, Deus ante tempora saecularia;
TITUS|1|3|manifestavit autem temporibus suis verbum suum in praedicatione, quae credita est mihi secundum praeceptum salvatoris nostri Dei,
TITUS|1|4|Tito germano filio secundum communem fidem: gratia et pax a Deo Patre et Christo Iesu salvatore nostro.
TITUS|1|5|Huius rei gratia reliqui te Cretae, ut ea, quae desunt, corrigas et constituas per civitates presbyteros, sicut ego tibi disposui,
TITUS|1|6|si quis sine crimine est, unius uxoris vir, filios habens fideles, non in accusatione luxuriae aut non subiectos.
TITUS|1|7|Oportet enim episcopum sine crimine esse sicut Dei dispensatorem, non superbum, non iracundum, non vinolentum, non percussorem, non turpis lucri cupidum,
TITUS|1|8|sed hospitalem, benignum, sobrium, iustum, sanctum, continentem,
TITUS|1|9|amplectentem eum, qui secundum doctrinam est, fidelem sermonem, ut potens sit et exhortari in doctrina sana et eos, qui contradicunt, arguere.
TITUS|1|10|Sunt enim multi et non subiecti, vaniloqui et seductores, maxime qui de circumcisione sunt,
TITUS|1|11|quibus oportet silentium imponere, quia universas domos subvertunt docentes, quae non oportet, turpis lucri gratia.
TITUS|1|12|Dixit quidam ex illis, proprius ipsorum propheta: " Cretenses semper mendaces, malae bestiae, ventres pigri ".
TITUS|1|13|Testimonium hoc verum est. Quam ob causam increpa illos dure, ut sani sint in fide,
TITUS|1|14|non intendentes Iudaicis fabulis et mandatis hominum aversantium veritatem.
TITUS|1|15|Omnia munda mundis; coinquinatis autem et infidelibus nihil mundum, sed inquinatae sunt eorum et mens et conscientia.
TITUS|1|16|Confitentur se nosse Deum, factis autem negant, cum sunt abominati et inoboedientes et ad omne opus bonum reprobi.
TITUS|2|1|Tu autem loquere, quae decent sanam doctrinam.
TITUS|2|2|Senes, ut sobrii sint, pudici, prudentes, sani fide, dilectione, patientia.
TITUS|2|3|Anus similiter in habitu sanctae, non criminatrices, non vino multo deditae, bene docentes,
TITUS|2|4|ut prudentiam doceant adulescentulas, ut viros suos ament, filios diligant,
TITUS|2|5|prudentes sint, castae, domus curam habentes, benignae, subditae suis viris, ut non blasphemetur verbum Dei.
TITUS|2|6|Iuvenes similiter hortare, ut sobrii sint.
TITUS|2|7|In omnibus teipsum praebens exemplum bonorum operum, in doctrina integritatem, gravitatem,
TITUS|2|8|in verbo sano irreprehensibilem, ut is, qui ex adverso est, vereatur, nihil habens malum dicere de nobis.
TITUS|2|9|Servos dominis suis subditos esse in omnibus, placentes esse, non contradicentes,
TITUS|2|10|non fraudantes, sed omnem fidem bonam ostendentes, ut doctrinam salutaris nostri Dei ornent in omnibus.
TITUS|2|11|Apparuit enim gratia Dei salutaris omnibus hominibus
TITUS|2|12|erudiens nos, ut abnegantes impietatem et saecularia desideria sobrie et iuste et pie vivamus in hoc saeculo,
TITUS|2|13|exspectantes beatam spem et adventum gloriae magni Dei et salvatoris nostri Iesu Christi;
TITUS|2|14|qui dedit semetipsum pro nobis, ut nos redimeret ab omni iniquitate et mundaret sibi populum peculiarem, sectatorem bonorum operum.
TITUS|2|15|Haec loquere et exhortare et argue cum omni imperio. Nemo te contemnat!
TITUS|3|1|Admone illos principibus, pote statibus subditos esse, dicto oboedire, ad omne opus bonum paratos esse,
TITUS|3|2|neminem blasphemare, non litigiosos esse, modestos, omnem ostendentes mansuetudinem ad omnes homines.
TITUS|3|3|Eramus enim et nos aliquando insipientes, inoboedientes, errantes, servientes concupiscentiis et voluptatibus variis, in malitia et invidia agentes, odibiles, odientes invicem.
TITUS|3|4|Cum autem benignitas et humanitas apparuit salvatoris nostri Dei,
TITUS|3|5|non ex operibus iustitiae, quae fecimus nos, sed secundum suam misericordiam salvos nos fecit per lavacrum regenerationis et renovationis Spiritus Sancti,
TITUS|3|6|quem effudit super nos abunde per Iesum Christum salvatorem nostrum,
TITUS|3|7|ut iustificati gratia ipsius heredes simus secundum spem vitae aeternae.
TITUS|3|8|Fidelis sermo, et volo te de his confirmare, ut curent bonis operibus praeesse, qui crediderunt Deo. Haec sunt bona et utilia hominibus;
TITUS|3|9|stultas autem quaestiones et genealogias et contentiones et pugnas circa legem devita, sunt enim inutiles et vanae.
TITUS|3|10|Haereticum hominem post unam et secundam correptionem devita,
TITUS|3|11|sciens quia subversus est, qui eiusmodi est, et delinquit, proprio iudicio condemnatus.
TITUS|3|12|Cum misero ad te Artemam aut Tychicum, festina ad me venire Nicopolim; ibi enim statui hiemare.
TITUS|3|13|Zenam legis peritum et Apollo sollicite instrue, ut nihil illis desit.
TITUS|3|14|Discant autem et nostri bonis operibus praeesse ad usus necessarios, ut non sint infructuosi.
TITUS|3|15|Salutant te, qui mecum sunt, omnes. Saluta, qui nos amant in fide.Gratia cum omnibus vobis.
