OBAD|1|1|The vision of Obadiah. This is what the Sovereign LORD says about Edom- We have heard a message from the LORD: An envoy was sent to the nations to say, "Rise, and let us go against her for battle"-
OBAD|1|2|"See, I will make you small among the nations; you will be utterly despised.
OBAD|1|3|The pride of your heart has deceived you, you who live in the clefts of the rocks and make your home on the heights, you who say to yourself, 'Who can bring me down to the ground?'
OBAD|1|4|Though you soar like the eagle and make your nest among the stars, from there I will bring you down," declares the LORD.
OBAD|1|5|"If thieves came to you, if robbers in the night- Oh, what a disaster awaits you- would they not steal only as much as they wanted? If grape pickers came to you, would they not leave a few grapes?
OBAD|1|6|But how Esau will be ransacked, his hidden treasures pillaged!
OBAD|1|7|All your allies will force you to the border; your friends will deceive and overpower you; those who eat your bread will set a trap for you, but you will not detect it.
OBAD|1|8|"In that day," declares the LORD, "will I not destroy the wise men of Edom, men of understanding in the mountains of Esau?
OBAD|1|9|Your warriors, O Teman, will be terrified, and everyone in Esau's mountains will be cut down in the slaughter.
OBAD|1|10|Because of the violence against your brother Jacob, you will be covered with shame; you will be destroyed forever.
OBAD|1|11|On the day you stood aloof while strangers carried off his wealth and foreigners entered his gates and cast lots for Jerusalem, you were like one of them.
OBAD|1|12|You should not look down on your brother in the day of his misfortune, nor rejoice over the people of Judah in the day of their destruction, nor boast so much in the day of their trouble.
OBAD|1|13|You should not march through the gates of my people in the day of their disaster, nor look down on them in their calamity in the day of their disaster, nor seize their wealth in the day of their disaster.
OBAD|1|14|You should not wait at the crossroads to cut down their fugitives, nor hand over their survivors in the day of their trouble.
OBAD|1|15|"The day of the LORD is near for all nations. As you have done, it will be done to you; your deeds will return upon your own head.
OBAD|1|16|Just as you drank on my holy hill, so all the nations will drink continually; they will drink and drink and be as if they had never been.
OBAD|1|17|But on Mount Zion will be deliverance; it will be holy, and the house of Jacob will possess its inheritance.
OBAD|1|18|The house of Jacob will be a fire and the house of Joseph a flame; the house of Esau will be stubble, and they will set it on fire and consume it. There will be no survivors from the house of Esau." The LORD has spoken.
OBAD|1|19|People from the Negev will occupy the mountains of Esau, and people from the foothills will possess the land of the Philistines. They will occupy the fields of Ephraim and Samaria, and Benjamin will possess Gilead.
OBAD|1|20|This company of Israelite exiles who are in Canaan will possess the land as far as Zarephath; the exiles from Jerusalem who are in Sepharad will possess the towns of the Negev.
OBAD|1|21|Deliverers will go up on Mount Zion to govern the mountains of Esau. And the kingdom will be the LORD's.
