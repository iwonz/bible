2PET|1|1|Симон Петр, раб и Апостол Иисуса Христа, принявшим с нами равно драгоценную веру по правде Бога нашего и Спасителя Иисуса Христа:
2PET|1|2|благодать и мир вам да умножится в познании Бога и Христа Иисуса, Господа нашего.
2PET|1|3|Как от Божественной силы Его даровано нам все потребное для жизни и благочестия, через познание Призвавшего нас славою и благостию,
2PET|1|4|которыми дарованы нам великие и драгоценные обетования, дабы вы через них соделались причастниками Божеского естества, удалившись от господствующего в мире растления похотью:
2PET|1|5|то вы, прилагая к сему все старание, покажите в вере вашей добродетель, в добродетели рассудительность,
2PET|1|6|в рассудительности воздержание, в воздержании терпение, в терпении благочестие,
2PET|1|7|в благочестии братолюбие, в братолюбии любовь.
2PET|1|8|Если это в вас есть и умножается, то вы не останетесь без успеха и плода в познании Господа нашего Иисуса Христа.
2PET|1|9|А в ком нет сего, тот слеп, закрыл глаза, забыл об очищении прежних грехов своих.
2PET|1|10|Посему, братия, более и более старайтесь делать твердым ваше звание и избрание; так поступая, никогда не преткнетесь,
2PET|1|11|ибо так откроется вам свободный вход в вечное Царство Господа нашего и Спасителя Иисуса Христа.
2PET|1|12|Для того я никогда не перестану напоминать вам о сем, хотя вы то и знаете, и утверждены в настоящей истине.
2PET|1|13|Справедливым же почитаю, доколе нахожусь в этой [телесной] храмине, возбуждать вас напоминанием,
2PET|1|14|зная, что скоро должен оставить храмину мою, как и Господь наш Иисус Христос открыл мне.
2PET|1|15|Буду же стараться, чтобы вы и после моего отшествия всегда приводили это на память.
2PET|1|16|Ибо мы возвестили вам силу и пришествие Господа нашего Иисуса Христа, не хитросплетенным басням последуя, но быв очевидцами Его величия.
2PET|1|17|Ибо Он принял от Бога Отца честь и славу, когда от велелепной славы принесся к Нему такой глас: Сей есть Сын Мой возлюбленный, в Котором Мое благоволение.
2PET|1|18|И этот глас, принесшийся с небес, мы слышали, будучи с Ним на святой горе.
2PET|1|19|И притом мы имеем вернейшее пророческое слово; и вы хорошо делаете, что обращаетесь к нему, как к светильнику, сияющему в темном месте, доколе не начнет рассветать день и не взойдет утренняя звезда в сердцах ваших,
2PET|1|20|зная прежде всего то, что никакого пророчества в Писании нельзя разрешить самому собою.
2PET|1|21|Ибо никогда пророчество не было произносимо по воле человеческой, но изрекали его святые Божии человеки, будучи движимы Духом Святым.
2PET|2|1|Были и лжепророки в народе, как и у вас будут лжеучители, которые введут пагубные ереси и, отвергаясь искупившего их Господа, навлекут сами на себя скорую погибель.
2PET|2|2|И многие последуют их разврату, и через них путь истины будет в поношении.
2PET|2|3|И из любостяжания будут уловлять вас льстивыми словами; суд им давно готов, и погибель их не дремлет.
2PET|2|4|Ибо, если Бог ангелов согрешивших не пощадил, но, связав узами адского мрака, предал блюсти на суд для наказания;
2PET|2|5|и если не пощадил первого мира, но в восьми душах сохранил семейство Ноя, проповедника правды, когда навел потоп на мир нечестивых;
2PET|2|6|и если города Содомские и Гоморрские, осудив на истребление, превратил в пепел, показав пример будущим нечестивцам,
2PET|2|7|а праведного Лота, утомленного обращением между людьми неистово развратными, избавил
2PET|2|8|(ибо сей праведник, живя между ними, ежедневно мучился в праведной душе, видя и слыша дела беззаконные) –
2PET|2|9|то, конечно, знает Господь, как избавлять благочестивых от искушения, а беззаконников соблюдать ко дню суда, для наказания,
2PET|2|10|а наипаче тех, которые идут вслед скверных похотей плоти, презирают начальства, дерзки, своевольны и не страшатся злословить высших,
2PET|2|11|тогда как и Ангелы, превосходя их крепостью и силою, не произносят на них пред Господом укоризненного суда.
2PET|2|12|Они, как бессловесные животные, водимые природою, рожденные на уловление и истребление, злословя то, чего не понимают, в растлении своем истребятся.
2PET|2|13|Они получат возмездие за беззаконие, ибо они полагают удовольствие во вседневной роскоши; срамники и осквернители, они наслаждаются обманами своими, пиршествуя с вами.
2PET|2|14|Глаза у них исполнены любострастия и непрестанного греха; они прельщают неутвержденные души; сердце их приучено к любостяжанию: это сыны проклятия.
2PET|2|15|Оставив прямой путь, они заблудились, идя по следам Валаама, сына Восорова, который возлюбил мзду неправедную,
2PET|2|16|но был обличен в своем беззаконии: бессловесная ослица, проговорив человеческим голосом, остановила безумие пророка.
2PET|2|17|Это безводные источники, облака и мглы, гонимые бурею: им приготовлен мрак вечной тьмы.
2PET|2|18|Ибо, произнося надутое пустословие, они уловляют в плотские похоти и разврат тех, которые едва отстали от находящихся в заблуждении.
2PET|2|19|Обещают им свободу, будучи сами рабы тления; ибо, кто кем побежден, тот тому и раб.
2PET|2|20|Ибо если, избегнув скверн мира чрез познание Господа и Спасителя нашего Иисуса Христа, опять запутываются в них и побеждаются ими, то последнее бывает для таковых хуже первого.
2PET|2|21|Лучше бы им не познать пути правды, нежели, познав, возвратиться назад от преданной им святой заповеди.
2PET|2|22|Но с ними случается по верной пословице: пес возвращается на свою блевотину, и: вымытая свинья [идет] валяться в грязи.
2PET|3|1|Это уже второе послание пишу к вам, возлюбленные; в них напоминанием возбуждаю ваш чистый смысл,
2PET|3|2|чтобы вы помнили слова, прежде реченные святыми пророками, и заповедь Господа и Спасителя, преданную Апостолами вашими.
2PET|3|3|Прежде всего знайте, что в последние дни явятся наглые ругатели, поступающие по собственным своим похотям
2PET|3|4|и говорящие: где обетование пришествия Его? Ибо с тех пор, как стали умирать отцы, от начала творения, все остается так же.
2PET|3|5|Думающие так не знают, что вначале словом Божиим небеса и земля составлены из воды и водою:
2PET|3|6|потому тогдашний мир погиб, быв потоплен водою.
2PET|3|7|А нынешние небеса и земля, содержимые тем же Словом, сберегаются огню на день суда и погибели нечестивых человеков.
2PET|3|8|Одно то не должно быть сокрыто от вас, возлюбленные, что у Господа один день, как тысяча лет, и тысяча лет, как один день.
2PET|3|9|Не медлит Господь [исполнением] обетования, как некоторые почитают то медлением; но долготерпит нас, не желая, чтобы кто погиб, но чтобы все пришли к покаянию.
2PET|3|10|Придет же день Господень, как тать ночью, и тогда небеса с шумом прейдут, стихии же, разгоревшись, разрушатся, земля и все дела на ней сгорят.
2PET|3|11|Если так все это разрушится, то какими должно быть в святой жизни и благочестии вам,
2PET|3|12|ожидающим и желающим пришествия дня Божия, в который воспламененные небеса разрушатся и разгоревшиеся стихии растают?
2PET|3|13|Впрочем мы, по обетованию Его, ожидаем нового неба и новой земли, на которых обитает правда.
2PET|3|14|Итак, возлюбленные, ожидая сего, потщитесь явиться пред Ним неоскверненными и непорочными в мире;
2PET|3|15|и долготерпение Господа нашего почитайте спасением, как и возлюбленный брат наш Павел, по данной ему премудрости, написал вам,
2PET|3|16|как он говорит об этом и во всех посланиях, в которых есть нечто неудобовразумительное, что невежды и неутвержденные, к собственной своей погибели, превращают, как и прочие Писания.
2PET|3|17|Итак вы, возлюбленные, будучи предварены о сем, берегитесь, чтобы вам не увлечься заблуждением беззаконников и не отпасть от своего утверждения,
2PET|3|18|но возрастайте в благодати и познании Господа нашего и Спасителя Иисуса Христа. Ему слава и ныне и в день вечный. Аминь.
