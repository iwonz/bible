GAL|1|1|Paul, an apostle--sent not from men nor by man, but by Jesus Christ and God the Father, who raised him from the dead--
GAL|1|2|and all the brothers with me, To the churches in Galatia:
GAL|1|3|Grace and peace to you from God our Father and the Lord Jesus Christ,
GAL|1|4|who gave himself for our sins to rescue us from the present evil age, according to the will of our God and Father,
GAL|1|5|to whom be glory for ever and ever. Amen.
GAL|1|6|I am astonished that you are so quickly deserting the one who called you by the grace of Christ and are turning to a different gospel--
GAL|1|7|which is really no gospel at all. Evidently some people are throwing you into confusion and are trying to pervert the gospel of Christ.
GAL|1|8|But even if we or an angel from heaven should preach a gospel other than the one we preached to you, let him be eternally condemned!
GAL|1|9|As we have already said, so now I say again: If anybody is preaching to you a gospel other than what you accepted, let him be eternally condemned!
GAL|1|10|Am I now trying to win the approval of men, or of God? Or am I trying to please men? If I were still trying to please men, I would not be a servant of Christ.
GAL|1|11|I want you to know, brothers, that the gospel I preached is not something that man made up.
GAL|1|12|I did not receive it from any man, nor was I taught it; rather, I received it by revelation from Jesus Christ.
GAL|1|13|For you have heard of my previous way of life in Judaism, how intensely I persecuted the church of God and tried to destroy it.
GAL|1|14|I was advancing in Judaism beyond many Jews of my own age and was extremely zealous for the traditions of my fathers.
GAL|1|15|But when God, who set me apart from birth and called me by his grace, was pleased
GAL|1|16|to reveal his Son in me so that I might preach him among the Gentiles, I did not consult any man,
GAL|1|17|nor did I go up to Jerusalem to see those who were apostles before I was, but I went immediately into Arabia and later returned to Damascus.
GAL|1|18|Then after three years, I went up to Jerusalem to get acquainted with Peter and stayed with him fifteen days.
GAL|1|19|I saw none of the other apostles--only James, the Lord's brother.
GAL|1|20|I assure you before God that what I am writing you is no lie.
GAL|1|21|Later I went to Syria and Cilicia.
GAL|1|22|I was personally unknown to the churches of Judea that are in Christ.
GAL|1|23|They only heard the report: "The man who formerly persecuted us is now preaching the faith he once tried to destroy."
GAL|1|24|And they praised God because of me.
GAL|2|1|Fourteen years later I went up again to Jerusalem, this time with Barnabas. I took Titus along also.
GAL|2|2|I went in response to a revelation and set before them the gospel that I preach among the Gentiles. But I did this privately to those who seemed to be leaders, for fear that I was running or had run my race in vain.
GAL|2|3|Yet not even Titus, who was with me, was compelled to be circumcised, even though he was a Greek.
GAL|2|4|This matter arose because some false brothers had infiltrated our ranks to spy on the freedom we have in Christ Jesus and to make us slaves.
GAL|2|5|We did not give in to them for a moment, so that the truth of the gospel might remain with you.
GAL|2|6|As for those who seemed to be important--whatever they were makes no difference to me; God does not judge by external appearance--those men added nothing to my message.
GAL|2|7|On the contrary, they saw that I had been entrusted with the task of preaching the gospel to the Gentiles, just as Peter had been to the Jews.
GAL|2|8|For God, who was at work in the ministry of Peter as an apostle to the Jews, was also at work in my ministry as an apostle to the Gentiles.
GAL|2|9|James, Peter and John, those reputed to be pillars, gave me and Barnabas the right hand of fellowship when they recognized the grace given to me. They agreed that we should go to the Gentiles, and they to the Jews.
GAL|2|10|All they asked was that we should continue to remember the poor, the very thing I was eager to do.
GAL|2|11|When Peter came to Antioch, I opposed him to his face, because he was clearly in the wrong.
GAL|2|12|Before certain men came from James, he used to eat with the Gentiles. But when they arrived, he began to draw back and separate himself from the Gentiles because he was afraid of those who belonged to the circumcision group.
GAL|2|13|The other Jews joined him in his hypocrisy, so that by their hypocrisy even Barnabas was led astray.
GAL|2|14|When I saw that they were not acting in line with the truth of the gospel, I said to Peter in front of them all, "You are a Jew, yet you live like a Gentile and not like a Jew. How is it, then, that you force Gentiles to follow Jewish customs?
GAL|2|15|"We who are Jews by birth and not 'Gentile sinners'
GAL|2|16|know that a man is not justified by observing the law, but by faith in Jesus Christ. So we, too, have put our faith in Christ Jesus that we may be justified by faith in Christ and not by observing the law, because by observing the law no one will be justified.
GAL|2|17|"If, while we seek to be justified in Christ, it becomes evident that we ourselves are sinners, does that mean that Christ promotes sin? Absolutely not!
GAL|2|18|If I rebuild what I destroyed, I prove that I am a lawbreaker.
GAL|2|19|For through the law I died to the law so that I might live for God.
GAL|2|20|I have been crucified with Christ and I no longer live, but Christ lives in me. The life I live in the body, I live by faith in the Son of God, who loved me and gave himself for me.
GAL|2|21|I do not set aside the grace of God, for if righteousness could be gained through the law, Christ died for nothing!"
GAL|3|1|You foolish Galatians! Who has bewitched you? Before your very eyes Jesus Christ was clearly portrayed as crucified.
GAL|3|2|I would like to learn just one thing from you: Did you receive the Spirit by observing the law, or by believing what you heard?
GAL|3|3|Are you so foolish? After beginning with the Spirit, are you now trying to attain your goal by human effort?
GAL|3|4|Have you suffered so much for nothing--if it really was for nothing?
GAL|3|5|Does God give you his Spirit and work miracles among you because you observe the law, or because you believe what you heard?
GAL|3|6|Consider Abraham: "He believed God, and it was credited to him as righteousness."
GAL|3|7|Understand, then, that those who believe are children of Abraham.
GAL|3|8|The Scripture foresaw that God would justify the Gentiles by faith, and announced the gospel in advance to Abraham: "All nations will be blessed through you."
GAL|3|9|So those who have faith are blessed along with Abraham, the man of faith.
GAL|3|10|All who rely on observing the law are under a curse, for it is written: "Cursed is everyone who does not continue to do everything written in the Book of the Law."
GAL|3|11|Clearly no one is justified before God by the law, because, "The righteous will live by faith."
GAL|3|12|The law is not based on faith; on the contrary, "The man who does these things will live by them."
GAL|3|13|Christ redeemed us from the curse of the law by becoming a curse for us, for it is written: "Cursed is everyone who is hung on a tree."
GAL|3|14|He redeemed us in order that the blessing given to Abraham might come to the Gentiles through Christ Jesus, so that by faith we might receive the promise of the Spirit.
GAL|3|15|Brothers, let me take an example from everyday life. Just as no one can set aside or add to a human covenant that has been duly established, so it is in this case.
GAL|3|16|The promises were spoken to Abraham and to his seed. The Scripture does not say "and to seeds," meaning many people, but "and to your seed," meaning one person, who is Christ.
GAL|3|17|What I mean is this: The law, introduced 430 years later, does not set aside the covenant previously established by God and thus do away with the promise.
GAL|3|18|For if the inheritance depends on the law, then it no longer depends on a promise; but God in his grace gave it to Abraham through a promise.
GAL|3|19|What, then, was the purpose of the law? It was added because of transgressions until the Seed to whom the promise referred had come. The law was put into effect through angels by a mediator.
GAL|3|20|A mediator, however, does not represent just one party; but God is one.
GAL|3|21|Is the law, therefore, opposed to the promises of God? Absolutely not! For if a law had been given that could impart life, then righteousness would certainly have come by the law.
GAL|3|22|But the Scripture declares that the whole world is a prisoner of sin, so that what was promised, being given through faith in Jesus Christ, might be given to those who believe.
GAL|3|23|Before this faith came, we were held prisoners by the law, locked up until faith should be revealed.
GAL|3|24|So the law was put in charge to lead us to Christ that we might be justified by faith.
GAL|3|25|Now that faith has come, we are no longer under the supervision of the law.
GAL|3|26|You are all sons of God through faith in Christ Jesus,
GAL|3|27|for all of you who were baptized into Christ have clothed yourselves with Christ.
GAL|3|28|There is neither Jew nor Greek, slave nor free, male nor female, for you are all one in Christ Jesus.
GAL|3|29|If you belong to Christ, then you are Abraham's seed, and heirs according to the promise.
GAL|4|1|What I am saying is that as long as the heir is a child, he is no different from a slave, although he owns the whole estate.
GAL|4|2|He is subject to guardians and trustees until the time set by his father.
GAL|4|3|So also, when we were children, we were in slavery under the basic principles of the world.
GAL|4|4|But when the time had fully come, God sent his Son, born of a woman, born under law,
GAL|4|5|to redeem those under law, that we might receive the full rights of sons.
GAL|4|6|Because you are sons, God sent the Spirit of his Son into our hearts, the Spirit who calls out, "Abba, Father."
GAL|4|7|So you are no longer a slave, but a son; and since you are a son, God has made you also an heir.
GAL|4|8|Formerly, when you did not know God, you were slaves to those who by nature are not gods.
GAL|4|9|But now that you know God--or rather are known by God--how is it that you are turning back to those weak and miserable principles? Do you wish to be enslaved by them all over again?
GAL|4|10|You are observing special days and months and seasons and years!
GAL|4|11|I fear for you, that somehow I have wasted my efforts on you.
GAL|4|12|I plead with you, brothers, become like me, for I became like you. You have done me no wrong.
GAL|4|13|As you know, it was because of an illness that I first preached the gospel to you.
GAL|4|14|Even though my illness was a trial to you, you did not treat me with contempt or scorn. Instead, you welcomed me as if I were an angel of God, as if I were Christ Jesus himself.
GAL|4|15|What has happened to all your joy? I can testify that, if you could have done so, you would have torn out your eyes and given them to me.
GAL|4|16|Have I now become your enemy by telling you the truth?
GAL|4|17|Those people are zealous to win you over, but for no good. What they want is to alienate you from us, so that you may be zealous for them.
GAL|4|18|It is fine to be zealous, provided the purpose is good, and to be so always and not just when I am with you.
GAL|4|19|My dear children, for whom I am again in the pains of childbirth until Christ is formed in you,
GAL|4|20|how I wish I could be with you now and change my tone, because I am perplexed about you!
GAL|4|21|Tell me, you who want to be under the law, are you not aware of what the law says?
GAL|4|22|For it is written that Abraham had two sons, one by the slave woman and the other by the free woman.
GAL|4|23|His son by the slave woman was born in the ordinary way; but his son by the free woman was born as the result of a promise.
GAL|4|24|These things may be taken figuratively, for the women represent two covenants. One covenant is from Mount Sinai and bears children who are to be slaves: This is Hagar.
GAL|4|25|Now Hagar stands for Mount Sinai in Arabia and corresponds to the present city of Jerusalem, because she is in slavery with her children.
GAL|4|26|But the Jerusalem that is above is free, and she is our mother.
GAL|4|27|For it is written: "Be glad, O barren woman, who bears no children; break forth and cry aloud, you who have no labor pains; because more are the children of the desolate woman than of her who has a husband."
GAL|4|28|Now you, brothers, like Isaac, are children of promise.
GAL|4|29|At that time the son born in the ordinary way persecuted the son born by the power of the Spirit. It is the same now.
GAL|4|30|But what does the Scripture say? "Get rid of the slave woman and her son, for the slave woman's son will never share in the inheritance with the free woman's son."
GAL|4|31|Therefore, brothers, we are not children of the slave woman, but of the free woman.
GAL|5|1|It is for freedom that Christ has set us free. Stand firm, then, and do not let yourselves be burdened again by a yoke of slavery.
GAL|5|2|Mark my words! I, Paul, tell you that if you let yourselves be circumcised, Christ will be of no value to you at all.
GAL|5|3|Again I declare to every man who lets himself be circumcised that he is obligated to obey the whole law.
GAL|5|4|You who are trying to be justified by law have been alienated from Christ; you have fallen away from grace.
GAL|5|5|But by faith we eagerly await through the Spirit the righteousness for which we hope.
GAL|5|6|For in Christ Jesus neither circumcision nor uncircumcision has any value. The only thing that counts is faith expressing itself through love.
GAL|5|7|You were running a good race. Who cut in on you and kept you from obeying the truth?
GAL|5|8|That kind of persuasion does not come from the one who calls you.
GAL|5|9|"A little yeast works through the whole batch of dough."
GAL|5|10|I am confident in the Lord that you will take no other view. The one who is throwing you into confusion will pay the penalty, whoever he may be.
GAL|5|11|Brothers, if I am still preaching circumcision, why am I still being persecuted? In that case the offense of the cross has been abolished.
GAL|5|12|As for those agitators, I wish they would go the whole way and emasculate themselves!
GAL|5|13|You, my brothers, were called to be free. But do not use your freedom to indulge the sinful nature; rather, serve one another in love.
GAL|5|14|The entire law is summed up in a single command: "Love your neighbor as yourself."
GAL|5|15|If you keep on biting and devouring each other, watch out or you will be destroyed by each other.
GAL|5|16|So I say, live by the Spirit, and you will not gratify the desires of the sinful nature.
GAL|5|17|For the sinful nature desires what is contrary to the Spirit, and the Spirit what is contrary to the sinful nature. They are in conflict with each other, so that you do not do what you want.
GAL|5|18|But if you are led by the Spirit, you are not under law.
GAL|5|19|The acts of the sinful nature are obvious: sexual immorality, impurity and debauchery;
GAL|5|20|idolatry and witchcraft; hatred, discord, jealousy, fits of rage, selfish ambition, dissensions, factions
GAL|5|21|and envy; drunkenness, orgies, and the like. I warn you, as I did before, that those who live like this will not inherit the kingdom of God.
GAL|5|22|But the fruit of the Spirit is love, joy, peace, patience, kindness, goodness, faithfulness,
GAL|5|23|gentleness and self-control. Against such things there is no law.
GAL|5|24|Those who belong to Christ Jesus have crucified the sinful nature with its passions and desires.
GAL|5|25|Since we live by the Spirit, let us keep in step with the Spirit.
GAL|5|26|Let us not become conceited, provoking and envying each other.
GAL|6|1|Brothers, if someone is caught in a sin, you who are spiritual should restore him gently. But watch yourself, or you also may be tempted.
GAL|6|2|Carry each other's burdens, and in this way you will fulfill the law of Christ.
GAL|6|3|If anyone thinks he is something when he is nothing, he deceives himself.
GAL|6|4|Each one should test his own actions. Then he can take pride in himself, without comparing himself to somebody else,
GAL|6|5|for each one should carry his own load.
GAL|6|6|Anyone who receives instruction in the word must share all good things with his instructor.
GAL|6|7|Do not be deceived: God cannot be mocked. A man reaps what he sows.
GAL|6|8|The one who sows to please his sinful nature, from that nature will reap destruction; the one who sows to please the Spirit, from the Spirit will reap eternal life.
GAL|6|9|Let us not become weary in doing good, for at the proper time we will reap a harvest if we do not give up.
GAL|6|10|Therefore, as we have opportunity, let us do good to all people, especially to those who belong to the family of believers.
GAL|6|11|See what large letters I use as I write to you with my own hand!
GAL|6|12|Those who want to make a good impression outwardly are trying to compel you to be circumcised. The only reason they do this is to avoid being persecuted for the cross of Christ.
GAL|6|13|Not even those who are circumcised obey the law, yet they want you to be circumcised that they may boast about your flesh.
GAL|6|14|May I never boast except in the cross of our Lord Jesus Christ, through which the world has been crucified to me, and I to the world.
GAL|6|15|Neither circumcision nor uncircumcision means anything; what counts is a new creation.
GAL|6|16|Peace and mercy to all who follow this rule, even to the Israel of God.
GAL|6|17|Finally, let no one cause me trouble, for I bear on my body the marks of Jesus.
GAL|6|18|The grace of our Lord Jesus Christ be with your spirit, brothers. Amen.
