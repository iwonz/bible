LUKE|1|1|Inasmuch as many have undertaken to compile a narrative of the things that have been accomplished among us,
LUKE|1|2|just as those who from the beginning were eyewitnesses and ministers of the word have delivered them to us,
LUKE|1|3|it seemed good to me also, having followed all things closely for some time past, to write an orderly account for you, most excellent Theophilus,
LUKE|1|4|that you may have certainty concerning the things you have been taught.
LUKE|1|5|In the days of Herod, king of Judea, there was a priest named Zechariah, of the division of Abijah. And he had a wife from the daughters of Aaron, and her name was Elizabeth.
LUKE|1|6|And they were both righteous before God, walking blamelessly in all the commandments and statutes of the Lord.
LUKE|1|7|But they had no child, because Elizabeth was barren, and both were advanced in years.
LUKE|1|8|Now while he was serving as priest before God when his division was on duty,
LUKE|1|9|according to the custom of the priesthood, he was chosen by lot to enter the temple of the Lord and burn incense.
LUKE|1|10|And the whole multitude of the people were praying outside at the hour of incense.
LUKE|1|11|And there appeared to him an angel of the Lord standing on the right side of the altar of incense.
LUKE|1|12|And Zechariah was troubled when he saw him, and fear fell upon him.
LUKE|1|13|But the angel said to him, "Do not be afraid, Zechariah, for your prayer has been heard, and your wife Elizabeth will bear you a son, and you shall call his name John.
LUKE|1|14|And you will have joy and gladness, and many will rejoice at his birth,
LUKE|1|15|for he will be great before the Lord. And he must not drink wine or strong drink, and he will be filled with the Holy Spirit, even from his mother's womb.
LUKE|1|16|And he will turn many of the children of Israel to the Lord their God,
LUKE|1|17|and he will go before him in the spirit and power of Elijah, to turn the hearts of the fathers to the children, and the disobedient to the wisdom of the just, to make ready for the Lord a people prepared."
LUKE|1|18|And Zechariah said to the angel, "How shall I know this? For I am an old man, and my wife is advanced in years."
LUKE|1|19|And the angel answered him, "I am Gabriel, who stands in the presence of God, and I was sent to speak to you and to bring you this good news.
LUKE|1|20|And behold, you will be silent and unable to speak until the day that these things take place, because you did not believe my words, which will be fulfilled in their time."
LUKE|1|21|And the people were waiting for Zechariah, and they were wondering at his delay in the temple.
LUKE|1|22|And when he came out, he was unable to speak to them, and they realized that he had seen a vision in the temple. And he kept making signs to them and remained mute.
LUKE|1|23|And when his time of service was ended, he went to his home.
LUKE|1|24|After these days his wife Elizabeth conceived, and for five months she kept herself hidden, saying,
LUKE|1|25|"Thus the Lord has done for me in the days when he looked on me, to take away my reproach among people."
LUKE|1|26|In the sixth month the angel Gabriel was sent from God to a city of Galilee named Nazareth,
LUKE|1|27|to a virgin betrothed to a man whose name was Joseph, of the house of David. And the virgin's name was Mary.
LUKE|1|28|And he came to her and said, "Greetings, O favored one, the Lord is with you!"
LUKE|1|29|But she was greatly troubled at the saying, and tried to discern what sort of greeting this might be.
LUKE|1|30|And the angel said to her, "Do not be afraid, Mary, for you have found favor with God.
LUKE|1|31|And behold, you will conceive in your womb and bear a son, and you shall call his name Jesus.
LUKE|1|32|He will be great and will be called the Son of the Most High. And the Lord God will give to him the throne of his father David,
LUKE|1|33|and he will reign over the house of Jacob forever, and of his kingdom there will be no end."
LUKE|1|34|And Mary said to the angel, "How will this be, since I am a virgin?"
LUKE|1|35|And the angel answered her, "The Holy Spirit will come upon you, and the power of the Most High will overshadow you; therefore the child to be born will be called holy- the Son of God.
LUKE|1|36|And behold, your relative Elizabeth in her old age has also conceived a son, and this is the sixth month with her who was called barren.
LUKE|1|37|For nothing will be impossible with God."
LUKE|1|38|And Mary said, "Behold, I am the servant of the Lord; let it be to me according to your word." And the angel departed from her.
LUKE|1|39|In those days Mary arose and went with haste into the hill country, to a town in Judah,
LUKE|1|40|and she entered the house of Zechariah and greeted Elizabeth.
LUKE|1|41|And when Elizabeth heard the greeting of Mary, the baby leaped in her womb. And Elizabeth was filled with the Holy Spirit,
LUKE|1|42|and she exclaimed with a loud cry, "Blessed are you among women, and blessed is the fruit of your womb!
LUKE|1|43|And why is this granted to me that the mother of my Lord should come to me?
LUKE|1|44|For behold, when the sound of your greeting came to my ears, the baby in my womb leaped for joy.
LUKE|1|45|And blessed is she who believed that there would be a fulfillment of what was spoken to her from the Lord."
LUKE|1|46|And Mary said, "My soul magnifies the Lord,
LUKE|1|47|and my spirit rejoices in God my Savior,
LUKE|1|48|for he has looked on the humble estate of his servant. For behold, from now on all generations will call me blessed;
LUKE|1|49|for he who is mighty has done great things for me, and holy is his name.
LUKE|1|50|And his mercy is for those who fear him from generation to generation.
LUKE|1|51|He has shown strength with his arm; he has scattered the proud in the thoughts of their hearts;
LUKE|1|52|he has brought down the mighty from their thrones and exalted those of humble estate;
LUKE|1|53|he has filled the hungry with good things, and the rich he has sent empty away.
LUKE|1|54|He has helped his servant Israel, in remembrance of his mercy,
LUKE|1|55|as he spoke to our fathers, to Abraham and to his offspring forever."
LUKE|1|56|And Mary remained with her about three months and returned to her home.
LUKE|1|57|Now the time came for Elizabeth to give birth, and she bore a son.
LUKE|1|58|And her neighbors and relatives heard that the Lord had shown great mercy to her, and they rejoiced with her.
LUKE|1|59|And on the eighth day they came to circumcise the child. And they would have called him Zechariah after his father,
LUKE|1|60|but his mother answered, "No; he shall be called John."
LUKE|1|61|And they said to her, "None of your relatives is called by this name."
LUKE|1|62|And they made signs to his father, inquiring what he wanted him to be called.
LUKE|1|63|And he asked for a writing tablet and wrote, "His name is John." And they all wondered.
LUKE|1|64|And immediately his mouth was opened and his tongue loosed, and he spoke, blessing God.
LUKE|1|65|And fear came on all their neighbors. And all these things were talked about through all the hill country of Judea,
LUKE|1|66|and all who heard them laid them up in their hearts, saying, "What then will this child be?" For the hand of the Lord was with him.
LUKE|1|67|And his father Zechariah was filled with the Holy Spirit and prophesied, saying,
LUKE|1|68|"Blessed be the Lord God of Israel, for he has visited and redeemed his people
LUKE|1|69|and has raised up a horn of salvation for us in the house of his servant David,
LUKE|1|70|as he spoke by the mouth of his holy prophets from of old,
LUKE|1|71|that we should be saved from our enemies and from the hand of all who hate us;
LUKE|1|72|to show the mercy promised to our fathers and to remember his holy covenant,
LUKE|1|73|the oath that he swore to our father Abraham, to grant us
LUKE|1|74|that we, being delivered from the hand of our enemies, might serve him without fear,
LUKE|1|75|in holiness and righteousness before him all our days.
LUKE|1|76|And you, child, will be called the prophet of the Most High; for you will go before the Lord to prepare his ways,
LUKE|1|77|to give knowledge of salvation to his people in the forgiveness of their sins,
LUKE|1|78|because of the tender mercy of our God, whereby the sunrise shall visit us from on high
LUKE|1|79|to give light to those who sit in darkness and in the shadow of death, to guide our feet into the way of peace."
LUKE|1|80|And the child grew and became strong in spirit, and he was in the wilderness until the day of his public appearance to Israel.
LUKE|2|1|In those days a decree went out from Caesar Augustus that all the world should be registered.
LUKE|2|2|This was the first registration when Quirinius was governor of Syria.
LUKE|2|3|And all went to be registered, each to his own town.
LUKE|2|4|And Joseph also went up from Galilee, from the town of Nazareth, to Judea, to the city of David, which is called Bethlehem, because he was of the house and lineage of David,
LUKE|2|5|to be registered with Mary, his betrothed, who was with child.
LUKE|2|6|And while they were there, the time came for her to give birth.
LUKE|2|7|And she gave birth to her firstborn son and wrapped him in swaddling cloths and laid him in a manger, because there was no place for them in the inn.
LUKE|2|8|And in the same region there were shepherds out in the field, keeping watch over their flock by night.
LUKE|2|9|And an angel of the Lord appeared to them, and the glory of the Lord shone around them, and they were filled with fear.
LUKE|2|10|And the angel said to them, "Fear not, for behold, I bring you good news of a great joy that will be for all the people.
LUKE|2|11|For unto you is born this day in the city of David a Savior, who is Christ the Lord.
LUKE|2|12|And this will be a sign for you: you will find a baby wrapped in swaddling cloths and lying in a manger."
LUKE|2|13|And suddenly there was with the angel a multitude of the heavenly host praising God and saying,
LUKE|2|14|"Glory to God in the highest, and on earth peace among those with whom he is pleased!"
LUKE|2|15|When the angels went away from them into heaven, the shepherds said to one another, "Let us go over to Bethlehem and see this thing that has happened, which the Lord has made known to us."
LUKE|2|16|And they went with haste and found Mary and Joseph, and the baby lying in a manger.
LUKE|2|17|And when they saw it, they made known the saying that had been told them concerning this child.
LUKE|2|18|And all who heard it wondered at what the shepherds told them.
LUKE|2|19|But Mary treasured up all these things, pondering them in her heart.
LUKE|2|20|And the shepherds returned, glorifying and praising God for all they had heard and seen, as it had been told them.
LUKE|2|21|And at the end of eight days, when he was circumcised, he was called Jesus, the name given by the angel before he was conceived in the womb.
LUKE|2|22|And when the time came for their purification according to the Law of Moses, they brought him up to Jerusalem to present him to the Lord
LUKE|2|23|(as it is written in the Law of the Lord, "Every male who first opens the womb shall be called holy to the Lord")
LUKE|2|24|and to offer a sacrifice according to what is said in the Law of the Lord, "a pair of turtledoves, or two young pigeons."
LUKE|2|25|Now there was a man in Jerusalem, whose name was Simeon, and this man was righteous and devout, waiting for the consolation of Israel, and the Holy Spirit was upon him.
LUKE|2|26|And it had been revealed to him by the Holy Spirit that he would not see death before he had seen the Lord's Christ.
LUKE|2|27|And he came in the Spirit into the temple, and when the parents brought in the child Jesus, to do for him according to the custom of the Law,
LUKE|2|28|he took him up in his arms and blessed God and said,
LUKE|2|29|"Lord, now you are letting your servant depart in peace, according to your word;
LUKE|2|30|for my eyes have seen your salvation
LUKE|2|31|that you have prepared in the presence of all peoples,
LUKE|2|32|a light for revelation to the Gentiles, and for glory to your people Israel."
LUKE|2|33|And his father and his mother marveled at what was said about him.
LUKE|2|34|And Simeon blessed them and said to Mary his mother, "Behold, this child is appointed for the fall and rising of many in Israel, and for a sign that is opposed
LUKE|2|35|(and a sword will pierce through your own soul also), so that thoughts from many hearts may be revealed."
LUKE|2|36|And there was a prophetess, Anna, the daughter of Phanuel, of the tribe of Asher. She was advanced in years, having lived with her husband seven years from when she was a virgin,
LUKE|2|37|and then as a widow until she was eighty-four. She did not depart from the temple, worshiping with fasting and prayer night and day.
LUKE|2|38|And coming up at that very hour she began to give thanks to God and to speak of him to all who were waiting for the redemption of Jerusalem.
LUKE|2|39|And when they had performed everything according to the Law of the Lord, they returned into Galilee, to their own town of Nazareth.
LUKE|2|40|And the child grew and became strong, filled with wisdom. And the favor of God was upon him.
LUKE|2|41|Now his parents went to Jerusalem every year at the Feast of the Passover.
LUKE|2|42|And when he was twelve years old, they went up according to custom.
LUKE|2|43|And when the feast was ended, as they were returning, the boy Jesus stayed behind in Jerusalem. His parents did not know it,
LUKE|2|44|but supposing him to be in the group they went a day's journey, but then they began to search for him among their relatives and acquaintances,
LUKE|2|45|and when they did not find him, they returned to Jerusalem, searching for him.
LUKE|2|46|After three days they found him in the temple, sitting among the teachers, listening to them and asking them questions.
LUKE|2|47|And all who heard him were amazed at his understanding and his answers.
LUKE|2|48|And when his parents saw him, they were astonished. And his mother said to him, "Son, why have you treated us so? Behold, your father and I have been searching for you in great distress."
LUKE|2|49|And he said to them, "Why were you looking for me? Did you not know that I must be in my Father's house?"
LUKE|2|50|And they did not understand the saying that he spoke to them.
LUKE|2|51|And he went down with them and came to Nazareth and was submissive to them. And his mother treasured up all these things in her heart.
LUKE|2|52|And Jesus increased in wisdom and in stature and in favor with God and man.
LUKE|3|1|In the fifteenth year of the reign of Tiberius Caesar, Pontius Pilate being governor of Judea, and Herod being tetrarch of Galilee, and his brother Philip tetrarch of the region of Ituraea and Trachonitis, and Lysanias tetrarch of Abilene,
LUKE|3|2|during the high priesthood of Annas and Caiaphas, the word of God came to John the son of Zechariah in the wilderness.
LUKE|3|3|And he went into all the region around the Jordan, proclaiming a baptism of repentance for the forgiveness of sins.
LUKE|3|4|As it is written in the book of the words of Isaiah the prophet, "The voice of one crying in the wilderness: Prepare the way of the Lord, make his paths straight.
LUKE|3|5|Every valley shall be filled, and every mountain and hill shall be made low, and the crooked shall become straight, and the rough places shall become level ways,
LUKE|3|6|and all flesh shall see the salvation of God."
LUKE|3|7|He said therefore to the crowds that came out to be baptized by him, "You brood of vipers! Who warned you to flee from the wrath to come?
LUKE|3|8|Bear fruits in keeping with repentance. And do not begin to say to yourselves, 'We have Abraham as our father.' For I tell you, God is able from these stones to raise up children for Abraham.
LUKE|3|9|Even now the axe is laid to the root of the trees. Every tree therefore that does not bear good fruit is cut down and thrown into the fire."
LUKE|3|10|And the crowds asked him, "What then shall we do?"
LUKE|3|11|And he answered them, "Whoever has two tunics is to share with him who has none, and whoever has food is to do likewise."
LUKE|3|12|Tax collectors also came to be baptized and said to him, "Teacher, what shall we do?"
LUKE|3|13|And he said to them, "Collect no more than you are authorized to do."
LUKE|3|14|Soldiers also asked him, "And we, what shall we do?" And he said to them, "Do not extort money from anyone by threats or by false accusation, and be content with your wages."
LUKE|3|15|As the people were in expectation, and all were questioning in their hearts concerning John, whether he might be the Christ,
LUKE|3|16|John answered them all, saying, "I baptize you with water, but he who is mightier than I is coming, the strap of whose sandals I am not worthy to untie. He will baptize you with the Holy Spirit and with fire.
LUKE|3|17|His winnowing fork is in his hand, to clear his threshing floor and to gather the wheat into his barn, but the chaff he will burn with unquenchable fire."
LUKE|3|18|So with many other exhortations he preached good news to the people.
LUKE|3|19|But Herod the tetrarch, who had been reproved by him for Herodias, his brother's wife, and for all the evil things that Herod had done,
LUKE|3|20|added this to them all, that he locked up John in prison.
LUKE|3|21|Now when all the people were baptized, and when Jesus also had been baptized and was praying, the heavens were opened,
LUKE|3|22|and the Holy Spirit descended on him in bodily form, like a dove; and a voice came from heaven, "You are my beloved Son; with you I am well pleased."
LUKE|3|23|Jesus, when he began his ministry, was about thirty years of age, being the son (as was supposed) of Joseph, the son of Heli,
LUKE|3|24|the son of Matthat, the son of Levi, the son of Melchi, the son of Jannai, the son of Joseph,
LUKE|3|25|the son of Mattathias, the son of Amos, the son of Nahum, the son of Esli, the son of Naggai,
LUKE|3|26|the son of Maath, the son of Mattathias, the son of Semein, the son of Josech, the son of Joda,
LUKE|3|27|the son of Joanan, the son of Rhesa, the son of Zerubbabel, the son of Shealtiel, the son of Neri,
LUKE|3|28|the son of Melchi, the son of Addi, the son of Cosam, the son of Elmadam, the son of Er,
LUKE|3|29|the son of Joshua, the son of Eliezer, the son of Jorim, the son of Matthat, the son of Levi,
LUKE|3|30|the son of Simeon, the son of Judah, the son of Joseph, the son of Jonam, the son of Eliakim,
LUKE|3|31|the son of Melea, the son of Menna, the son of Mattatha, the son of Nathan, the son of David,
LUKE|3|32|the son of Jesse, the son of Obed, the son of Boaz, the son of Sala, the son of Nahshon,
LUKE|3|33|the son of Amminadab, the son of Admin, the son of Arni, the son of Hezron, the son of Perez, the son of Judah,
LUKE|3|34|the son of Jacob, the son of Isaac, the son of Abraham, the son of Terah, the son of Nahor,
LUKE|3|35|the son of Serug, the son of Reu, the son of Peleg, the son of Eber, the son of Shelah,
LUKE|3|36|the son of Cainan, the son of Arphaxad, the son of Shem, the son of Noah, the son of Lamech,
LUKE|3|37|the son of Methuselah, the son of Enoch, the son of Jared, the son of Mahalaleel, the son of Cainan,
LUKE|3|38|the son of Enos, the son of Seth, the son of Adam, the son of God.
LUKE|4|1|And Jesus, full of the Holy Spirit, returned from the Jordan and was led by the Spirit in the wilderness
LUKE|4|2|for forty days, being tempted by the devil. And he ate nothing during those days. And when they were ended, he was hungry.
LUKE|4|3|The devil said to him, "If you are the Son of God, command this stone to become bread."
LUKE|4|4|And Jesus answered him, "It is written, 'Man shall not live by bread alone.'"
LUKE|4|5|And the devil took him up and showed him all the kingdoms of the world in a moment of time,
LUKE|4|6|and said to him, "To you I will give all this authority and their glory, for it has been delivered to me, and I give it to whom I will.
LUKE|4|7|If you, then, will worship me, it will all be yours."
LUKE|4|8|And Jesus answered him, "It is written, "' You shall worship the Lord your God, and him only shall you serve.'"
LUKE|4|9|And he took him to Jerusalem and set him on the pinnacle of the temple and said to him, "If you are the Son of God, throw yourself down from here,
LUKE|4|10|for it is written, "' He will command his angels concerning you, to guard you,'
LUKE|4|11|and "'On their hands they will bear you up, lest you strike your foot against a stone.'"
LUKE|4|12|And Jesus answered him, "It is said, 'You shall not put the Lord your God to the test.'"
LUKE|4|13|And when the devil had ended every temptation, he departed from him until an opportune time.
LUKE|4|14|And Jesus returned in the power of the Spirit to Galilee, and a report about him went out through all the surrounding country.
LUKE|4|15|And he taught in their synagogues, being glorified by all.
LUKE|4|16|And he came to Nazareth, where he had been brought up. And as was his custom, he went to the synagogue on the Sabbath day, and he stood up to read.
LUKE|4|17|And the scroll of the prophet Isaiah was given to him. He unrolled the scroll and found the place where it was written,
LUKE|4|18|"The Spirit of the Lord is upon me, because he has anointed me to proclaim good news to the poor. He has sent me to proclaim liberty to the captives and recovering of sight to the blind, to set at liberty those who are oppressed,
LUKE|4|19|to proclaim the year of the Lord's favor."
LUKE|4|20|And he rolled up the scroll and gave it back to the attendant and sat down. And the eyes of all in the synagogue were fixed on him.
LUKE|4|21|And he began to say to them, "Today this Scripture has been fulfilled in your hearing."
LUKE|4|22|And all spoke well of him and marveled at the gracious words that were coming from his mouth. And they said, "Is not this Joseph's son?"
LUKE|4|23|And he said to them, "Doubtless you will quote to me this proverb, 'Physician, heal yourself.' What we have heard you did at Capernaum, do here in your hometown as well."
LUKE|4|24|And he said, "Truly, I say to you, no prophet is acceptable in his hometown.
LUKE|4|25|But in truth, I tell you, there were many widows in Israel in the days of Elijah, when the heavens were shut up three years and six months, and a great famine came over all the land,
LUKE|4|26|and Elijah was sent to none of them but only to Zarephath, in the land of Sidon, to a woman who was a widow.
LUKE|4|27|And there were many lepers in Israel in the time of the prophet Elisha, and none of them was cleansed, but only Naaman the Syrian."
LUKE|4|28|When they heard these things, all in the synagogue were filled with wrath.
LUKE|4|29|And they rose up and drove him out of the town and brought him to the brow of the hill on which their town was built, so that they could throw him down the cliff.
LUKE|4|30|But passing through their midst, he went away.
LUKE|4|31|And he went down to Capernaum, a city of Galilee. And he was teaching them on the Sabbath,
LUKE|4|32|and they were astonished at his teaching, for his word possessed authority.
LUKE|4|33|And in the synagogue there was a man who had the spirit of an unclean demon, and he cried out with a loud voice,
LUKE|4|34|"Ha! What have you to do with us, Jesus of Nazareth? Have you come to destroy us? I know who you are- the Holy One of God."
LUKE|4|35|But Jesus rebuked him, saying, "Be silent and come out of him!" And when the demon had thrown him down in their midst, he came out of him, having done him no harm.
LUKE|4|36|And they were all amazed and said to one another, "What is this word? For with authority and power he commands the unclean spirits, and they come out!"
LUKE|4|37|And reports about him went out into every place in the surrounding region.
LUKE|4|38|And he arose and left the synagogue and entered Simon's house. Now Simon's mother-in-law was ill with a high fever, and they appealed to him on her behalf.
LUKE|4|39|And he stood over her and rebuked the fever, and it left her, and immediately she rose and began to serve them.
LUKE|4|40|Now when the sun was setting, all those who had any who were sick with various diseases brought them to him, and he laid his hands on every one of them and healed them.
LUKE|4|41|And demons also came out of many, crying, "You are the Son of God!" But he rebuked them and would not allow them to speak, because they knew that he was the Christ.
LUKE|4|42|And when it was day, he departed and went into a desolate place. And the people sought him and came to him, and would have kept him from leaving them,
LUKE|4|43|but he said to them, "I must preach the good news of the kingdom of God to the other towns as well; for I was sent for this purpose."
LUKE|4|44|And he was preaching in the synagogues of Judea.
LUKE|5|1|On one occasion, while the crowd was pressing in on him to hear the word of God, he was standing by the lake of Gennesaret,
LUKE|5|2|and he saw two boats by the lake, but the fishermen had gone out of them and were washing their nets.
LUKE|5|3|Getting into one of the boats, which was Simon's, he asked him to put out a little from the land. And he sat down and taught the people from the boat.
LUKE|5|4|And when he had finished speaking, he said to Simon, "Put out into the deep and let down your nets for a catch."
LUKE|5|5|And Simon answered, "Master, we toiled all night and took nothing! But at your word I will let down the nets."
LUKE|5|6|And when they had done this, they enclosed a large number of fish, and their nets were breaking.
LUKE|5|7|They signaled to their partners in the other boat to come and help them. And they came and filled both the boats, so that they began to sink.
LUKE|5|8|But when Simon Peter saw it, he fell down at Jesus' knees, saying, "Depart from me, for I am a sinful man, O Lord."
LUKE|5|9|For he and all who were with him were astonished at the catch of fish that they had taken,
LUKE|5|10|and so also were James and John, sons of Zebedee, who were partners with Simon. And Jesus said to Simon, "Do not be afraid; from now on you will be catching men."
LUKE|5|11|And when they had brought their boats to land, they left everything and followed him.
LUKE|5|12|While he was in one of the cities, there came a man full of leprosy. And when he saw Jesus, he fell on his face and begged him, "Lord, if you will, you can make me clean."
LUKE|5|13|And Jesus stretched out his hand and touched him, saying, "I will; be clean." And immediately the leprosy left him.
LUKE|5|14|And he charged him to tell no one, but "go and show yourself to the priest, and make an offering for your cleansing, as Moses commanded, for a proof to them."
LUKE|5|15|But now even more the report about him went abroad, and great crowds gathered to hear him and to be healed of their infirmities.
LUKE|5|16|But he would withdraw to desolate places and pray.
LUKE|5|17|On one of those days, as he was teaching, Pharisees and teachers of the law were sitting there, who had come from every village of Galilee and Judea and from Jerusalem. And the power of the Lord was with him to heal.
LUKE|5|18|And behold, some men were bringing on a bed a man who was paralyzed, and they were seeking to bring him in and lay him before Jesus,
LUKE|5|19|but finding no way to bring him in, because of the crowd, they went up on the roof and let him down with his bed through the tiles into the midst before Jesus.
LUKE|5|20|And when he saw their faith, he said, "Man, your sins are forgiven you."
LUKE|5|21|And the scribes and the Pharisees began to question, saying, "Who is this who speaks blasphemies? Who can forgive sins but God alone?"
LUKE|5|22|When Jesus perceived their thoughts, he answered them, "Why do you question in your hearts?
LUKE|5|23|Which is easier, to say, 'Your sins are forgiven you,' or to say, 'Rise and walk'?
LUKE|5|24|But that you may know that the Son of Man has authority on earth to forgive sins"- he said to the man who was paralyzed- "I say to you, rise, pick up your bed and go home."
LUKE|5|25|And immediately he rose up before them and picked up what he had been lying on and went home, glorifying God.
LUKE|5|26|And amazement seized them all, and they glorified God and were filled with awe, saying, "We have seen extraordinary things today."
LUKE|5|27|After this he went out and saw a tax collector named Levi, sitting at the tax booth. And he said to him, "Follow me."
LUKE|5|28|And leaving everything, he rose and followed him.
LUKE|5|29|And Levi made him a great feast in his house, and there was a large company of tax collectors and others reclining at table with them.
LUKE|5|30|And the Pharisees and their scribes grumbled at his disciples, saying, "Why do you eat and drink with tax collectors and sinners?"
LUKE|5|31|And Jesus answered them, "Those who are well have no need of a physician, but those who are sick.
LUKE|5|32|I have not come to call the righteous but sinners to repentance."
LUKE|5|33|And they said to him, "The disciples of John fast often and offer prayers, and so do the disciples of the Pharisees, but yours eat and drink."
LUKE|5|34|And Jesus said to them, "Can you make wedding guests fast while the bridegroom is with them?
LUKE|5|35|The days will come when the bridegroom is taken away from them, and then they will fast in those days."
LUKE|5|36|He also told them a parable: "No one tears a piece from a new garment and puts it on an old garment. If he does, he will tear the new, and the piece from the new will not match the old.
LUKE|5|37|And no one puts new wine into old wineskins. If he does, the new wine will burst the skins and it will be spilled, and the skins will be destroyed.
LUKE|5|38|But new wine must be put into fresh wineskins.
LUKE|5|39|And no one after drinking old wine desires new, for he says, 'The old is good.'"
LUKE|6|1|On a Sabbath, while he was going through the grainfields, his disciples plucked and ate some heads of grain, rubbing them in their hands.
LUKE|6|2|But some of the Pharisees said, "Why are you doing what is not lawful to do on the Sabbath?"
LUKE|6|3|And Jesus answered them, "Have you not read what David did when he was hungry, he and those who were with him:
LUKE|6|4|how he entered the house of God and took and ate the bread of the Presence, which is not lawful for any but the priests to eat, and also gave it to those with him?"
LUKE|6|5|And he said to them, "The Son of Man is lord of the Sabbath."
LUKE|6|6|On another Sabbath, he entered the synagogue and was teaching, and a man was there whose right hand was withered.
LUKE|6|7|And the scribes and the Pharisees watched him, to see whether he would heal on the Sabbath, so that they might find a reason to accuse him.
LUKE|6|8|But he knew their thoughts, and he said to the man with the withered hand, "Come and stand here." And he rose and stood there.
LUKE|6|9|And Jesus said to them, "I ask you, is it lawful on the Sabbath to do good or to do harm, to save life or to destroy it?"
LUKE|6|10|And after looking around at them all he said to him, "Stretch out your hand." And he did so, and his hand was restored.
LUKE|6|11|But they were filled with fury and discussed with one another what they might do to Jesus.
LUKE|6|12|In these days he went out to the mountain to pray, and all night he continued in prayer to God.
LUKE|6|13|And when day came, he called his disciples and chose from them twelve, whom he named apostles:
LUKE|6|14|Simon, whom he named Peter, and Andrew his brother, and James and John, and Philip, and Bartholomew,
LUKE|6|15|and Matthew, and Thomas, and James the son of Alphaeus, and Simon who was called the Zealot,
LUKE|6|16|and Judas the son of James, and Judas Iscariot, who became a traitor.
LUKE|6|17|And he came down with them and stood on a level place, with a great crowd of his disciples and a great multitude of people from all Judea and Jerusalem and the seacoast of Tyre and Sidon,
LUKE|6|18|who came to hear him and to be healed of their diseases. And those who were troubled with unclean spirits were cured.
LUKE|6|19|And all the crowd sought to touch him, for power came out from him and healed them all.
LUKE|6|20|And he lifted up his eyes on his disciples, and said: "Blessed are you who are poor, for yours is the kingdom of God.
LUKE|6|21|"Blessed are you who are hungry now, for you shall be satisfied. "Blessed are you who weep now, for you shall laugh.
LUKE|6|22|"Blessed are you when people hate you and when they exclude you and revile you and spurn your name as evil, on account of the Son of Man!
LUKE|6|23|Rejoice in that day, and leap for joy, for behold, your reward is great in heaven; for so their fathers did to the prophets.
LUKE|6|24|"But woe to you who are rich, for you have received your consolation.
LUKE|6|25|"Woe to you who are full now, for you shall be hungry. "Woe to you who laugh now, for you shall mourn and weep.
LUKE|6|26|"Woe to you, when all people speak well of you, for so their fathers did to the false prophets.
LUKE|6|27|"But I say to you who hear, Love your enemies, do good to those who hate you,
LUKE|6|28|bless those who curse you, pray for those who abuse you.
LUKE|6|29|To one who strikes you on the cheek, offer the other also, and from one who takes away your cloak do not withhold your tunic either.
LUKE|6|30|Give to everyone who begs from you, and from one who takes away your goods do not demand them back.
LUKE|6|31|And as you wish that others would do to you, do so to them.
LUKE|6|32|"If you love those who love you, what benefit is that to you? For even sinners love those who love them.
LUKE|6|33|And if you do good to those who do good to you, what benefit is that to you? For even sinners do the same.
LUKE|6|34|And if you lend to those from whom you expect to receive, what credit is that to you? Even sinners lend to sinners, to get back the same amount.
LUKE|6|35|But love your enemies, and do good, and lend, expecting nothing in return, and your reward will be great, and you will be sons of the Most High, for he is kind to the ungrateful and the evil.
LUKE|6|36|Be merciful, even as your Father is merciful.
LUKE|6|37|"Judge not, and you will not be judged; condemn not, and you will not be condemned; forgive, and you will be forgiven;
LUKE|6|38|give, and it will be given to you. Good measure, pressed down, shaken together, running over, will be put into your lap. For with the measure you use it will be measured back to you."
LUKE|6|39|He also told them a parable: "Can a blind man lead a blind man? Will they not both fall into a pit?
LUKE|6|40|A disciple is not above his teacher, but everyone when he is fully trained will be like his teacher.
LUKE|6|41|Why do you see the speck that is in your brother's eye, but do not notice the log that is in your own eye?
LUKE|6|42|How can you say to your brother, 'Brother, let me take out the speck that is in your eye,' when you yourself do not see the log that is in your own eye? You hypocrite, first take the log out of your own eye, and then you will see clearly to take out the speck that is in your brother's eye.
LUKE|6|43|"For no good tree bears bad fruit, nor again does a bad tree bear good fruit,
LUKE|6|44|for each tree is known by its own fruit. For figs are not gathered from thornbushes, nor are grapes picked from a bramble bush.
LUKE|6|45|The good person out of the good treasure of his heart produces good, and the evil person out of his evil treasure produces evil, for out of the abundance of the heart his mouth speaks.
LUKE|6|46|"Why do you call me 'Lord, Lord,' and not do what I tell you?
LUKE|6|47|Everyone who comes to me and hears my words and does them, I will show you what he is like:
LUKE|6|48|he is like a man building a house, who dug deep and laid the foundation on the rock. And when a flood arose, the stream broke against that house and could not shake it, because it had been well built.
LUKE|6|49|But the one who hears and does not do them is like a man who built a house on the ground without a foundation. When the stream broke against it, immediately it fell, and the ruin of that house was great."
LUKE|7|1|After he had finished all his sayings in the hearing of the people, he entered Capernaum.
LUKE|7|2|Now a centurion had a servant who was sick and at the point of death, who was highly valued by him.
LUKE|7|3|When the centurion heard about Jesus, he sent to him elders of the Jews, asking him to come and heal his servant.
LUKE|7|4|And when they came to Jesus, they pleaded with him earnestly, saying, "He is worthy to have you do this for him,
LUKE|7|5|for he loves our nation, and he is the one who built us our synagogue."
LUKE|7|6|And Jesus went with them. When he was not far from the house, the centurion sent friends, saying to him, "Lord, do not trouble yourself, for I am not worthy to have you come under my roof.
LUKE|7|7|Therefore I did not presume to come to you. But say the word, and let my servant be healed.
LUKE|7|8|For I too am a man set under authority, with soldiers under me: and I say to one, 'Go,' and he goes; and to another, 'Come,' and he comes; and to my servant, 'Do this,' and he does it."
LUKE|7|9|When Jesus heard these things, he marveled at him, and turning to the crowd that followed him, said, "I tell you, not even in Israel have I found such faith."
LUKE|7|10|And when those who had been sent returned to the house, they found the servant well.
LUKE|7|11|Soon afterward he went to a town called Nain, and his disciples and a great crowd went with him.
LUKE|7|12|As he drew near to the gate of the town, behold, a man who had died was being carried out, the only son of his mother, and she was a widow, and a considerable crowd from the town was with her.
LUKE|7|13|And when the Lord saw her, he had compassion on her and said to her, "Do not weep."
LUKE|7|14|Then he came up and touched the bier, and the bearers stood still. And he said, "Young man, I say to you, arise."
LUKE|7|15|And the dead man sat up and began to speak, and Jesus gave him to his mother.
LUKE|7|16|Fear seized them all, and they glorified God, saying, "A great prophet has arisen among us!" and "God has visited his people!"
LUKE|7|17|And this report about him spread through the whole of Judea and all the surrounding country.
LUKE|7|18|The disciples of John reported all these things to him. And John,
LUKE|7|19|calling two of his disciples to him, sent them to the Lord, saying, "Are you the one who is to come, or shall we look for another?"
LUKE|7|20|And when the men had come to him, they said, "John the Baptist has sent us to you, saying, 'Are you the one who is to come, or shall we look for another?'"
LUKE|7|21|In that hour he healed many people of diseases and plagues and evil spirits, and on many who were blind he bestowed sight.
LUKE|7|22|And he answered them, "Go and tell John what you have seen and heard: the blind receive their sight, the lame walk, lepers are cleansed, and the deaf hear, the dead are raised up, the poor have good news preached to them.
LUKE|7|23|And blessed is the one who is not offended by me."
LUKE|7|24|When John's messengers had gone, Jesus began to speak to the crowds concerning John: "What did you go out into the wilderness to see? A reed shaken by the wind?
LUKE|7|25|What then did you go out to see? A man dressed in soft clothing? Behold, those who are dressed in splendid clothing and live in luxury are in kings' courts.
LUKE|7|26|What then did you go out to see? A prophet? Yes, I tell you, and more than a prophet.
LUKE|7|27|This is he of whom it is written, "' Behold, I send my messenger before your face, who will prepare your way before you.'
LUKE|7|28|I tell you, among those born of women none is greater than John. Yet the one who is least in the kingdom of God is greater than he."
LUKE|7|29|(When all the people heard this, and the tax collectors too, they declared God just, having been baptized with the baptism of John,
LUKE|7|30|but the Pharisees and the lawyers rejected the purpose of God for themselves, not having been baptized by him.)
LUKE|7|31|"To what then shall I compare the people of this generation, and what are they like?
LUKE|7|32|They are like children sitting in the marketplace and calling to one another, "' We played the flute for you, and you did not dance; we sang a dirge, and you did not weep.'
LUKE|7|33|For John the Baptist has come eating no bread and drinking no wine, and you say, 'He has a demon.'
LUKE|7|34|The Son of Man has come eating and drinking, and you say, 'Look at him! A glutton and a drunkard, a friend of tax collectors and sinners!'
LUKE|7|35|Yet wisdom is justified by all her children."
LUKE|7|36|One of the Pharisees asked him to eat with him, and he went into the Pharisee's house and took his place at the table.
LUKE|7|37|And behold, a woman of the city, who was a sinner, when she learned that he was reclining at table in the Pharisee's house, brought an alabaster flask of ointment,
LUKE|7|38|and standing behind him at his feet, weeping, she began to wet his feet with her tears and wiped them with the hair of her head and kissed his feet and anointed them with the ointment.
LUKE|7|39|Now when the Pharisee who had invited him saw this, he said to himself, "If this man were a prophet, he would have known who and what sort of woman this is who is touching him, for she is a sinner."
LUKE|7|40|And Jesus answering said to him, "Simon, I have something to say to you." And he answered, "Say it, Teacher."
LUKE|7|41|"A certain moneylender had two debtors. One owed five hundred denarii, and the other fifty.
LUKE|7|42|When they could not pay, he cancelled the debt of both. Now which of them will love him more?"
LUKE|7|43|Simon answered, "The one, I suppose, for whom he cancelled the larger debt." And he said to him, "You have judged rightly."
LUKE|7|44|Then turning toward the woman he said to Simon, "Do you see this woman? I entered your house; you gave me no water for my feet, but she has wet my feet with her tears and wiped them with her hair.
LUKE|7|45|You gave me no kiss, but from the time I came in she has not ceased to kiss my feet.
LUKE|7|46|You did not anoint my head with oil, but she has anointed my feet with ointment.
LUKE|7|47|Therefore I tell you, her sins, which are many, are forgiven- for she loved much. But he who is forgiven little, loves little."
LUKE|7|48|And he said to her, "Your sins are forgiven."
LUKE|7|49|Then those who were at table with him began to say among themselves, "Who is this, who even forgives sins?"
LUKE|7|50|And he said to the woman, "Your faith has saved you; go in peace."
LUKE|8|1|Soon afterward he went on through cities and villages, proclaiming and bringing the good news of the kingdom of God. And the twelve were with him,
LUKE|8|2|and also some women who had been healed of evil spirits and infirmities: Mary, called Magdalene, from whom seven demons had gone out,
LUKE|8|3|and Joanna, the wife of Chuza, Herod's household manager, and Susanna, and many others, who provided for them out of their means.
LUKE|8|4|And when a great crowd was gathering and people from town after town came to him, he said in a parable:
LUKE|8|5|"A sower went out to sow his seed. And as he sowed, some fell along the path and was trampled underfoot, and the birds of the air devoured it.
LUKE|8|6|And some fell on the rock, and as it grew up, it withered away, because it had no moisture.
LUKE|8|7|And some fell among thorns, and the thorns grew up with it and choked it.
LUKE|8|8|And some fell into good soil and grew and yielded a hundredfold." As he said these things, he called out, "He who has ears to hear, let him hear."
LUKE|8|9|And when his disciples asked him what this parable meant,
LUKE|8|10|he said, "To you it has been given to know the secrets of the kingdom of God, but for others they are in parables, so that 'seeing they may not see, and hearing they may not understand.'
LUKE|8|11|Now the parable is this: The seed is the word of God.
LUKE|8|12|The ones along the path are those who have heard. Then the devil comes and takes away the word from their hearts, so that they may not believe and be saved.
LUKE|8|13|And the ones on the rock are those who, when they hear the word, receive it with joy. But these have no root; they believe for a while, and in time of testing fall away.
LUKE|8|14|And as for what fell among the thorns, they are those who hear, but as they go on their way they are choked by the cares and riches and pleasures of life, and their fruit does not mature.
LUKE|8|15|As for that in the good soil, they are those who, hearing the word, hold it fast in an honest and good heart, and bear fruit with patience.
LUKE|8|16|"No one after lighting a lamp covers it with a jar or puts it under a bed, but puts it on a stand, so that those who enter may see the light.
LUKE|8|17|For nothing is hidden that will not be made manifest, nor is anything secret that will not be known and come to light.
LUKE|8|18|Take care then how you hear, for to the one who has, more will be given, and from the one who has not, even what he thinks that he has will be taken away."
LUKE|8|19|Then his mother and his brothers came to him, but they could not reach him because of the crowd.
LUKE|8|20|And he was told, "Your mother and your brothers are standing outside, desiring to see you."
LUKE|8|21|But he answered them, "My mother and my brothers are those who hear the word of God and do it."
LUKE|8|22|One day he got into a boat with his disciples, and he said to them, "Let us go across to the other side of the lake." So they set out,
LUKE|8|23|and as they sailed he fell asleep. And a windstorm came down on the lake, and they were filling with water and were in danger.
LUKE|8|24|And they went and woke him, saying, "Master, Master, we are perishing!" And he awoke and rebuked the wind and the raging waves, and they ceased, and there was a calm.
LUKE|8|25|He said to them, "Where is your faith?" And they were afraid, and they marveled, saying to one another, "Who then is this, that he commands even winds and water, and they obey him?"
LUKE|8|26|Then they sailed to the country of the Gerasenes, which is opposite Galilee.
LUKE|8|27|When Jesus had stepped out on land, there met him a man from the city who had demons. For a long time he had worn no clothes, and he had not lived in a house but among the tombs.
LUKE|8|28|When he saw Jesus, he cried out and fell down before him and said with a loud voice, "What have you to do with me, Jesus, Son of the Most High God? I beg you, do not torment me."
LUKE|8|29|For he had commanded the unclean spirit to come out of the man. (For many a time it had seized him. He was kept under guard and bound with chains and shackles, but he would break the bonds and be driven by the demon into the desert.)
LUKE|8|30|Jesus then asked him, "What is your name?" And he said, "Legion," for many demons had entered him.
LUKE|8|31|And they begged him not to command them to depart into the abyss.
LUKE|8|32|Now a large herd of pigs was feeding there on the hillside, and they begged him to let them enter these. So he gave them permission.
LUKE|8|33|Then the demons came out of the man and entered the pigs, and the herd rushed down the steep bank into the lake and were drowned.
LUKE|8|34|When the herdsmen saw what had happened, they fled and told it in the city and in the country.
LUKE|8|35|Then people went out to see what had happened, and they came to Jesus and found the man from whom the demons had gone, sitting at the feet of Jesus, clothed and in his right mind, and they were afraid.
LUKE|8|36|And those who had seen it told them how the demon-possessed man had been healed.
LUKE|8|37|Then all the people of the surrounding country of the Gerasenes asked him to depart from them, for they were seized with great fear. So he got into the boat and returned.
LUKE|8|38|The man from whom the demons had gone begged that he might be with him, but Jesus sent him away, saying,
LUKE|8|39|"Return to your home, and declare how much God has done for you." And he went away, proclaiming throughout the whole city how much Jesus had done for him.
LUKE|8|40|Now when Jesus returned, the crowd welcomed him, for they were all waiting for him.
LUKE|8|41|And there came a man named Jairus, who was a ruler of the synagogue. And falling at Jesus' feet, he implored him to come to his house,
LUKE|8|42|for he had an only daughter, about twelve years of age, and she was dying. As Jesus went, the people pressed around him.
LUKE|8|43|And there was a woman who had had a discharge of blood for twelve years, and though she had spent all her living on physicians, she could not be healed by anyone.
LUKE|8|44|She came up behind him and touched the fringe of his garment, and immediately her discharge of blood ceased.
LUKE|8|45|And Jesus said, "Who was it that touched me?" When all denied it, Peter said, "Master, the crowds surround you and are pressing in on you!"
LUKE|8|46|But Jesus said, "Someone touched me, for I perceive that power has gone out from me."
LUKE|8|47|And when the woman saw that she was not hidden, she came trembling, and falling down before him declared in the presence of all the people why she had touched him, and how she had been immediately healed.
LUKE|8|48|And he said to her, "Daughter, your faith has made you well; go in peace."
LUKE|8|49|While he was still speaking, someone from the ruler's house came and said, "Your daughter is dead; do not trouble the Teacher any more."
LUKE|8|50|But Jesus on hearing this answered him, "Do not fear; only believe, and she will be well."
LUKE|8|51|And when he came to the house, he allowed no one to enter with him, except Peter and John and James, and the father and mother of the child.
LUKE|8|52|And all were weeping and mourning for her, but he said, "Do not weep, for she is not dead but sleeping."
LUKE|8|53|And they laughed at him, knowing that she was dead.
LUKE|8|54|But taking her by the hand he called, saying, "Child, arise."
LUKE|8|55|And her spirit returned, and she got up at once. And he directed that something should be given her to eat.
LUKE|8|56|And her parents were amazed, but he charged them to tell no one what had happened.
LUKE|9|1|And he called the twelve together and gave them power and authority over all demons and to cure diseases,
LUKE|9|2|and he sent them out to proclaim the kingdom of God and to heal.
LUKE|9|3|And he said to them, "Take nothing for your journey, no staff, nor bag, nor bread, nor money; and do not have two tunics.
LUKE|9|4|And whatever house you enter, stay there, and from there depart.
LUKE|9|5|And wherever they do not receive you, when you leave that town shake off the dust from your feet as a testimony against them."
LUKE|9|6|And they departed and went through the villages, preaching the gospel and healing everywhere.
LUKE|9|7|Now Herod the tetrarch heard about all that was happening, and he was perplexed, because it was said by some that John had been raised from the dead,
LUKE|9|8|by some that Elijah had appeared, and by others that one of the prophets of old had risen.
LUKE|9|9|Herod said, "John I beheaded, but who is this about whom I hear such things?" And he sought to see him.
LUKE|9|10|On their return the apostles told him all that they had done. And he took them and withdrew apart to a town called Bethsaida.
LUKE|9|11|When the crowds learned it, they followed him, and he welcomed them and spoke to them of the kingdom of God and cured those who had need of healing.
LUKE|9|12|Now the day began to wear away, and the twelve came and said to him, "Send the crowd away to go into the surrounding villages and countryside to find lodging and get provisions, for we are here in a desolate place."
LUKE|9|13|But he said to them, "You give them something to eat." They said, "We have no more than five loaves and two fish- unless we are to go and buy food for all these people."
LUKE|9|14|For there were about five thousand men. And he said to his disciples, "Have them sit down in groups of about fifty each."
LUKE|9|15|And they did so, and had them all sit down.
LUKE|9|16|And taking the five loaves and the two fish, he looked up to heaven and said a blessing over them. Then he broke the loaves and gave them to the disciples to set before the crowd.
LUKE|9|17|And they all ate and were satisfied. And what was left over was picked up, twelve baskets of broken pieces.
LUKE|9|18|Now it happened that as he was praying alone, the disciples were with him. And he asked them, "Who do the crowds say that I am?"
LUKE|9|19|And they answered, "John the Baptist. But others say, Elijah, and others, that one of the prophets of old has risen."
LUKE|9|20|Then he said to them, "But who do you say that I am?" And Peter answered, "The Christ of God."
LUKE|9|21|And he strictly charged and commanded them to tell this to no one,
LUKE|9|22|saying, "The Son of Man must suffer many things and be rejected by the elders and chief priests and scribes, and be killed, and on the third day be raised."
LUKE|9|23|And he said to all, "If anyone would come after me, let him deny himself and take up his cross daily and follow me.
LUKE|9|24|For whoever would save his life will lose it, but whoever loses his life for my sake will save it.
LUKE|9|25|For what does it profit a man if he gains the whole world and loses or forfeits himself?
LUKE|9|26|For whoever is ashamed of me and of my words, of him will the Son of Man be ashamed when he comes in his glory and the glory of the Father and of the holy angels.
LUKE|9|27|But I tell you truly, there are some standing here who will not taste death until they see the kingdom of God."
LUKE|9|28|Now about eight days after these sayings he took with him Peter and John and James and went up on the mountain to pray.
LUKE|9|29|And as he was praying, the appearance of his face was altered, and his clothing became dazzling white.
LUKE|9|30|And behold, two men were talking with him, Moses and Elijah,
LUKE|9|31|who appeared in glory and spoke of his departure, which he was about to accomplish at Jerusalem.
LUKE|9|32|Now Peter and those who were with him were heavy with sleep, but when they became fully awake they saw his glory and the two men who stood with him.
LUKE|9|33|And as the men were parting from him, Peter said to Jesus, "Master, it is good that we are here. Let us make three tents, one for you and one for Moses and one for Elijah"- not knowing what he said.
LUKE|9|34|As he was saying these things, a cloud came and overshadowed them, and they were afraid as they entered the cloud.
LUKE|9|35|And a voice came out of the cloud, saying, "This is my Son, my Chosen One; listen to him!"
LUKE|9|36|And when the voice had spoken, Jesus was found alone. And they kept silent and told no one in those days anything of what they had seen.
LUKE|9|37|On the next day, when they had come down from the mountain, a great crowd met him.
LUKE|9|38|And behold, a man from the crowd cried out, "Teacher, I beg you to look at my son, for he is my only child.
LUKE|9|39|And behold, a spirit seizes him, and he suddenly cries out. It convulses him so that he foams at the mouth; and shatters him, and will hardly leave him.
LUKE|9|40|And I begged your disciples to cast it out, but they could not."
LUKE|9|41|Jesus answered, "O faithless and twisted generation, how long am I to be with you and bear with you? Bring your son here."
LUKE|9|42|While he was coming, the demon threw him to the ground and convulsed him. But Jesus rebuked the unclean spirit and healed the boy, and gave him back to his father.
LUKE|9|43|And all were astonished at the majesty of God. But while they were all marveling at everything he was doing, Jesus said to his disciples,
LUKE|9|44|"Let these words sink into your ears: The Son of Man is about to be delivered into the hands of men."
LUKE|9|45|But they did not understand this saying, and it was concealed from them, so that they might not perceive it. And they were afraid to ask him about this saying.
LUKE|9|46|An argument arose among them as to which of them was the greatest.
LUKE|9|47|But Jesus, knowing the reasoning of their hearts, took a child and put him by his side
LUKE|9|48|and said to them, "Whoever receives this child in my name receives me, and whoever receives me receives him who sent me. For he who is least among you all is the one who is great."
LUKE|9|49|John answered, "Master, we saw someone casting out demons in your name, and we tried to stop him, because he does not follow with us."
LUKE|9|50|But Jesus said to him, "Do not stop him, for the one who is not against you is for you."
LUKE|9|51|When the days drew near for him to be taken up, he set his face to go to Jerusalem.
LUKE|9|52|And he sent messengers ahead of him, who went and entered a village of the Samaritans, to make preparations for him.
LUKE|9|53|But the people did not receive him, because his face was set toward Jerusalem.
LUKE|9|54|And when his disciples James and John saw it, they said, "Lord, do you want us to tell fire to come down from heaven and consume them?"
LUKE|9|55|But he turned and rebuked them.
LUKE|9|56|And they went on to another village.
LUKE|9|57|As they were going along the road, someone said to him, "I will follow you wherever you go."
LUKE|9|58|And Jesus said to him, "Foxes have holes, and birds of the air have nests, but the Son of Man has nowhere to lay his head."
LUKE|9|59|To another he said, "Follow me." But he said, "Lord, let me first go and bury my father."
LUKE|9|60|And Jesus said to him, "Leave the dead to bury their own dead. But as for you, go and proclaim the kingdom of God."
LUKE|9|61|Yet another said, "I will follow you, Lord, but let me first say farewell to those at my home."
LUKE|9|62|Jesus said to him, "No one who puts his hand to the plow and looks back is fit for the kingdom of God."
LUKE|10|1|After this the Lord appointed seventy-two others and sent them on ahead of him, two by two, into every town and place where he himself was about to go.
LUKE|10|2|And he said to them, "The harvest is plentiful, but the laborers are few. Therefore pray earnestly to the Lord of the harvest to send out laborers into his harvest.
LUKE|10|3|Go your way; behold, I am sending you out as lambs in the midst of wolves.
LUKE|10|4|Carry no moneybag, no knapsack, no sandals, and greet no one on the road.
LUKE|10|5|Whatever house you enter, first say, 'Peace be to this house!'
LUKE|10|6|And if a son of peace is there, your peace will rest upon him. But if not, it will return to you.
LUKE|10|7|And remain in the same house, eating and drinking what they provide, for the laborer deserves his wages. Do not go from house to house.
LUKE|10|8|Whenever you enter a town and they receive you, eat what is set before you.
LUKE|10|9|Heal the sick in it and say to them, 'The kingdom of God has come near to you.'
LUKE|10|10|But whenever you enter a town and they do not receive you, go into its streets and say,
LUKE|10|11|'Even the dust of your town that clings to our feet we wipe off against you. Nevertheless know this, that the kingdom of God has come near.'
LUKE|10|12|I tell you, it will be more bearable on that day for Sodom than for that town.
LUKE|10|13|"Woe to you, Chorazin! Woe to you, Bethsaida! For if the mighty works done in you had been done in Tyre and Sidon, they would have repented long ago, sitting in sackcloth and ashes.
LUKE|10|14|But it will be more bearable in the judgment for Tyre and Sidon than for you.
LUKE|10|15|And you, Capernaum, will you be exalted to heaven? You shall be brought down to Hades.
LUKE|10|16|"The one who hears you hears me, and the one who rejects you rejects me, and the one who rejects me rejects him who sent me."
LUKE|10|17|The seventy-two returned with joy, saying, "Lord, even the demons are subject to us in your name!"
LUKE|10|18|And he said to them, "I saw Satan fall like lightning from heaven.
LUKE|10|19|Behold, I have given you authority to tread on serpents and scorpions, and over all the power of the enemy, and nothing shall hurt you.
LUKE|10|20|Nevertheless, do not rejoice in this, that the spirits are subject to you, but rejoice that your names are written in heaven."
LUKE|10|21|In that same hour he rejoiced in the Holy Spirit and said, "I thank you, Father, Lord of heaven and earth, that you have hidden these things from the wise and understanding and revealed them to little children; yes, Father, for such was your gracious will.
LUKE|10|22|All things have been handed over to me by my Father, and no one knows who the Son is except the Father, or who the Father is except the Son and anyone to whom the Son chooses to reveal him."
LUKE|10|23|Then turning to the disciples he said privately, "Blessed are the eyes that see what you see!
LUKE|10|24|For I tell you that many prophets and kings desired to see what you see, and did not see it, and to hear what you hear, and did not hear it."
LUKE|10|25|And behold, a lawyer stood up to put him to the test, saying, "Teacher, what shall I do to inherit eternal life?"
LUKE|10|26|He said to him, "What is written in the Law? How do you read it?"
LUKE|10|27|And he answered, "You shall love the Lord your God with all your heart and with all your soul and with all your strength and with all your mind, and your neighbor as yourself."
LUKE|10|28|And he said to him, "You have answered correctly; do this, and you will live."
LUKE|10|29|But he, desiring to justify himself, said to Jesus, "And who is my neighbor?"
LUKE|10|30|Jesus replied, "A man was going down from Jerusalem to Jericho, and he fell among robbers, who stripped him and beat him and departed, leaving him half dead.
LUKE|10|31|Now by chance a priest was going down that road, and when he saw him he passed by on the other side.
LUKE|10|32|So likewise a Levite, when he came to the place and saw him, passed by on the other side.
LUKE|10|33|But a Samaritan, as he journeyed, came to where he was, and when he saw him, he had compassion.
LUKE|10|34|He went to him and bound up his wounds, pouring on oil and wine. Then he set him on his own animal and brought him to an inn and took care of him.
LUKE|10|35|And the next day he took out two denarii and gave them to the innkeeper, saying, 'Take care of him, and whatever more you spend, I will repay you when I come back.'
LUKE|10|36|Which of these three, do you think, proved to be a neighbor to the man who fell among the robbers?"
LUKE|10|37|He said, "The one who showed him mercy." And Jesus said to him, "You go, and do likewise."
LUKE|10|38|Now as they went on their way, Jesus entered a village. And a woman named Martha welcomed him into her house.
LUKE|10|39|And she had a sister called Mary, who sat at the Lord's feet and listened to his teaching.
LUKE|10|40|But Martha was distracted with much serving. And she went up to him and said, "Lord, do you not care that my sister has left me to serve alone? Tell her then to help me."
LUKE|10|41|But the Lord answered her, "Martha, Martha, you are anxious and troubled about many things,
LUKE|10|42|but one thing is necessary. Mary has chosen the good portion, which will not be taken away from her."
LUKE|11|1|Now Jesus was praying in a certain place, and when he finished, one of his disciples said to him, "Lord, teach us to pray, as John taught his disciples."
LUKE|11|2|And he said to them, "When you pray, say: "Father, hallowed be your name. Your kingdom come.
LUKE|11|3|Give us each day our daily bread,
LUKE|11|4|and forgive us our sins, for we ourselves forgive everyone who is indebted to us. And lead us not into temptation."
LUKE|11|5|And he said to them, "Which of you who has a friend will go to him at midnight and say to him, 'Friend, lend me three loaves,
LUKE|11|6|for a friend of mine has arrived on a journey, and I have nothing to set before him';
LUKE|11|7|and he will answer from within, 'Do not bother me; the door is now shut, and my children are with me in bed. I cannot get up and give you anything'?
LUKE|11|8|I tell you, though he will not get up and give him anything because he is his friend, yet because of his impudence he will rise and give him whatever he needs.
LUKE|11|9|And I tell you, ask, and it will be given to you; seek, and you will find; knock, and it will be opened to you.
LUKE|11|10|For everyone who asks receives, and the one who seeks finds, and to the one who knocks it will be opened.
LUKE|11|11|What father among you, if his son asks for a fish, will instead of a fish give him a serpent;
LUKE|11|12|or if he asks for an egg, will give him a scorpion?
LUKE|11|13|If you then, who are evil, know how to give good gifts to your children, how much more will the heavenly Father give the Holy Spirit to those who ask him!"
LUKE|11|14|Now he was casting out a demon that was mute. When the demon had gone out, the mute man spoke, and the people marveled.
LUKE|11|15|But some of them said, "He casts out demons by Beelzebul, the prince of demons,"
LUKE|11|16|while others, to test him, kept seeking from him a sign from heaven.
LUKE|11|17|But he, knowing their thoughts, said to them, "Every kingdom divided against itself is laid waste, and a divided household falls.
LUKE|11|18|And if Satan also is divided against himself, how will his kingdom stand? For you say that I cast out demons by Beelzebul.
LUKE|11|19|And if I cast out demons by Beelzebul, by whom do your sons cast them out? Therefore they will be your judges.
LUKE|11|20|But if it is by the finger of God that I cast out demons, then the kingdom of God has come upon you.
LUKE|11|21|When a strong man, fully armed, guards his own palace, his goods are safe;
LUKE|11|22|but when one stronger than he attacks him and overcomes him, he takes away his armor in which he trusted and divides his spoil.
LUKE|11|23|Whoever is not with me is against me, and whoever does not gather with me scatters.
LUKE|11|24|"When the unclean spirit has gone out of a person, it passes through waterless places seeking rest, and finding none it says, 'I will return to my house from which I came.'
LUKE|11|25|And when it comes, it finds the house swept and put in order.
LUKE|11|26|Then it goes and brings seven other spirits more evil than itself, and they enter and dwell there. And the last state of that person is worse than the first."
LUKE|11|27|As he said these things, a woman in the crowd raised her voice and said to him, "Blessed is the womb that bore you, and the breasts at which you nursed!"
LUKE|11|28|But he said, "Blessed rather are those who hear the word of God and keep it!"
LUKE|11|29|When the crowds were increasing, he began to say, "This generation is an evil generation. It seeks for a sign, but no sign will be given to it except the sign of Jonah.
LUKE|11|30|For as Jonah became a sign to the people of Nineveh, so will the Son of Man be to this generation.
LUKE|11|31|The queen of the South will rise up at the judgment with the men of this generation and condemn them, for she came from the ends of the earth to hear the wisdom of Solomon, and behold, something greater than Solomon is here.
LUKE|11|32|The men of Nineveh will rise up at the judgment with this generation and condemn it, for they repented at the preaching of Jonah, and behold, something greater than Jonah is here.
LUKE|11|33|"No one after lighting a lamp puts it in a cellar or under a basket, but on a stand, so that those who enter may see the light.
LUKE|11|34|Your eye is the lamp of your body. When your eye is healthy, your whole body is full of light, but when it is bad, your body is full of darkness.
LUKE|11|35|Therefore be careful lest the light in you be darkness.
LUKE|11|36|If then your whole body is full of light, having no part dark, it will be wholly bright, as when a lamp with its rays gives you light."
LUKE|11|37|While Jesus was speaking, a Pharisee asked him to dine with him, so he went in and reclined at table.
LUKE|11|38|The Pharisee was astonished to see that he did not first wash before dinner.
LUKE|11|39|And the Lord said to him, "Now you Pharisees cleanse the outside of the cup and of the dish, but inside you are full of greed and wickedness.
LUKE|11|40|You fools! Did not he who made the outside make the inside also?
LUKE|11|41|But give as alms those things that are within, and behold, everything is clean for you.
LUKE|11|42|"But woe to you Pharisees! For you tithe mint and rue and every herb, and neglect justice and the love of God. These you ought to have done, without neglecting the others.
LUKE|11|43|Woe to you Pharisees! For you love the best seat in the synagogues and greetings in the marketplaces.
LUKE|11|44|Woe to you! For you are like unmarked graves, and people walk over them without knowing it."
LUKE|11|45|One of the lawyers answered him, "Teacher, in saying these things you insult us also."
LUKE|11|46|And he said, "Woe to you lawyers also! For you load people with burdens hard to bear, and you yourselves do not touch the burdens with one of your fingers.
LUKE|11|47|Woe to you! For you build the tombs of the prophets whom your fathers killed.
LUKE|11|48|So you are witnesses and you consent to the deeds of your fathers, for they killed them, and you build their tombs.
LUKE|11|49|Therefore also the Wisdom of God said, 'I will send them prophets and apostles, some of whom they will kill and persecute,'
LUKE|11|50|so that the blood of all the prophets, shed from the foundation of the world, may be charged against this generation,
LUKE|11|51|from the blood of Abel to the blood of Zechariah, who perished between the altar and the sanctuary. Yes, I tell you, it will be required of this generation.
LUKE|11|52|Woe to you lawyers! For you have taken away the key of knowledge. You did not enter yourselves, and you hindered those who were entering."
LUKE|11|53|As he went away from there, the scribes and the Pharisees began to press him hard and to provoke him to speak about many things,
LUKE|11|54|lying in wait for him, to catch him in something he might say.
LUKE|12|1|In the meantime, when so many thousands of the people had gathered together that they were trampling one another, he began to say to his disciples first, "Beware of the leaven of the Pharisees, which is hypocrisy.
LUKE|12|2|Nothing is covered up that will not be revealed, or hidden that will not be known.
LUKE|12|3|Therefore whatever you have said in the dark shall be heard in the light, and what you have whispered in private rooms shall be proclaimed on the housetops.
LUKE|12|4|"I tell you, my friends, do not fear those who kill the body, and after that have nothing more that they can do.
LUKE|12|5|But I will warn you whom to fear: fear him who, after he has killed, has authority to cast into hell. Yes, I tell you, fear him!
LUKE|12|6|Are not five sparrows sold for two pennies? And not one of them is forgotten before God.
LUKE|12|7|Why, even the hairs of your head are all numbered. Fear not; you are of more value than many sparrows.
LUKE|12|8|"And I tell you, everyone who acknowledges me before men, the Son of Man also will acknowledge before the angels of God,
LUKE|12|9|but the one who denies me before men will be denied before the angels of God.
LUKE|12|10|And everyone who speaks a word against the Son of Man will be forgiven, but the one who blasphemes against the Holy Spirit will not be forgiven.
LUKE|12|11|And when they bring you before the synagogues and the rulers and the authorities, do not be anxious about how you should defend yourself or what you should say,
LUKE|12|12|for the Holy Spirit will teach you in that very hour what you ought to say."
LUKE|12|13|Someone in the crowd said to him, "Teacher, tell my brother to divide the inheritance with me."
LUKE|12|14|But he said to him, "Man, who made me a judge or arbitrator over you?"
LUKE|12|15|And he said to them, "Take care, and be on your guard against all covetousness, for one's life does not consist in the abundance of his possessions."
LUKE|12|16|And he told them a parable, saying, "The land of a rich man produced plentifully,
LUKE|12|17|and he thought to himself, 'What shall I do, for I have nowhere to store my crops?'
LUKE|12|18|And he said, 'I will do this: I will tear down my barns and build larger ones, and there I will store all my grain and my goods.
LUKE|12|19|And I will say to my soul, Soul, you have ample goods laid up for many years; relax, eat, drink, be merry.'
LUKE|12|20|But God said to him, 'Fool! This night your soul is required of you, and the things you have prepared, whose will they be?'
LUKE|12|21|So is the one who lays up treasure for himself and is not rich toward God."
LUKE|12|22|And he said to his disciples, "Therefore I tell you, do not be anxious about your life, what you will eat, nor about your body, what you will put on.
LUKE|12|23|For life is more than food, and the body more than clothing.
LUKE|12|24|Consider the ravens: they neither sow nor reap, they have neither storehouse nor barn, and yet God feeds them. Of how much more value are you than the birds!
LUKE|12|25|And which of you by being anxious can add a single hour to his span of life?
LUKE|12|26|If then you are not able to do as small a thing as that, why are you anxious about the rest?
LUKE|12|27|Consider the lilies, how they grow: they neither toil nor spin, yet I tell you, even Solomon in all his glory was not arrayed like one of these.
LUKE|12|28|But if God so clothes the grass, which is alive in the field today, and tomorrow is thrown into the oven, how much more will he clothe you, O you of little faith!
LUKE|12|29|And do not seek what you are to eat and what you are to drink, nor be worried.
LUKE|12|30|For all the nations of the world seek after these things, and your Father knows that you need them.
LUKE|12|31|Instead, seek his kingdom, and these things will be added to you.
LUKE|12|32|"Fear not, little flock, for it is your Father's good pleasure to give you the kingdom.
LUKE|12|33|Sell your possessions, and give to the needy. Provide yourselves with moneybags that do not grow old, with a treasure in the heavens that does not fail, where no thief approaches and no moth destroys.
LUKE|12|34|For where your treasure is, there will your heart be also.
LUKE|12|35|"Stay dressed for action and keep your lamps burning,
LUKE|12|36|and be like men who are waiting for their master to come home from the wedding feast, so that they may open the door to him at once when he comes and knocks.
LUKE|12|37|Blessed are those servants whom the master finds awake when he comes. Truly, I say to you, he will dress himself for service and have them recline at table, and he will come and serve them.
LUKE|12|38|If he comes in the second watch, or in the third, and finds them awake, blessed are those servants!
LUKE|12|39|But know this, that if the master of the house had known at what hour the thief was coming, he would not have left his house to be broken into.
LUKE|12|40|You also must be ready, for the Son of Man is coming at an hour you do not expect."
LUKE|12|41|Peter said, "Lord, are you telling this parable for us or for all?"
LUKE|12|42|And the Lord said, "Who then is the faithful and wise manager, whom his master will set over his household, to give them their portion of food at the proper time?
LUKE|12|43|Blessed is that servant whom his master will find so doing when he comes.
LUKE|12|44|Truly, I say to you, he will set him over all his possessions.
LUKE|12|45|But if that servant says to himself, 'My master is delayed in coming,' and begins to beat the male and female servants, and to eat and drink and get drunk,
LUKE|12|46|the master of that servant will come on a day when he does not expect him and at an hour he does not know, and will cut him in pieces and put him with the unfaithful.
LUKE|12|47|And that servant who knew his master's will but did not get ready or act according to his will, will receive a severe beating.
LUKE|12|48|But the one who did not know, and did what deserved a beating, will receive a light beating. Everyone to whom much was given, of him much will be required, and from him to whom they entrusted much, they will demand the more.
LUKE|12|49|"I came to cast fire on the earth, and would that it were already kindled!
LUKE|12|50|I have a baptism to be baptized with, and how great is my distress until it is accomplished!
LUKE|12|51|Do you think that I have come to give peace on earth? No, I tell you, but rather division.
LUKE|12|52|For from now on in one house there will be five divided, three against two and two against three.
LUKE|12|53|They will be divided, father against son and son against father, mother against daughter and daughter against mother, mother-in-law against her daughter-in-law and daughter-in-law against mother-in-law."
LUKE|12|54|He also said to the crowds, "When you see a cloud rising in the west, you say at once, 'A shower is coming.' And so it happens.
LUKE|12|55|And when you see the south wind blowing, you say, 'There will be scorching heat,' and it happens.
LUKE|12|56|You hypocrites! You know how to interpret the appearance of earth and sky, but why do you not know how to interpret the present time?
LUKE|12|57|"And why do you not judge for yourselves what is right?
LUKE|12|58|As you go with your accuser before the magistrate, make an effort to settle with him on the way, lest he drag you to the judge, and the judge hand you over to the officer, and the officer put you in prison.
LUKE|12|59|I tell you, you will never get out until you have paid the very last penny."
LUKE|13|1|There were some present at that very time who told him about the Galileans whose blood Pilate had mingled with their sacrifices.
LUKE|13|2|And he answered them, "Do you think that these Galileans were worse sinners than all the other Galileans, because they suffered in this way?
LUKE|13|3|No, I tell you; but unless you repent, you will all likewise perish.
LUKE|13|4|Or those eighteen on whom the tower in Siloam fell and killed them: do you think that they were worse offenders than all the others who lived in Jerusalem?
LUKE|13|5|No, I tell you; but unless you repent, you will all likewise perish."
LUKE|13|6|And he told this parable: "A man had a fig tree planted in his vineyard, and he came seeking fruit on it and found none.
LUKE|13|7|And he said to the vinedresser, 'Look, for three years now I have come seeking fruit on this fig tree, and I find none. Cut it down. Why should it use up the ground?'
LUKE|13|8|And he answered him, 'Sir, let it alone this year also, until I dig around it and put on manure.
LUKE|13|9|Then if it should bear fruit next year, well and good; but if not, you can cut it down.'"
LUKE|13|10|Now he was teaching in one of the synagogues on the Sabbath.
LUKE|13|11|And there was a woman who had had a disabling spirit for eighteen years. She was bent over and could not fully straighten herself.
LUKE|13|12|When Jesus saw her, he called her over and said to her, "Woman, you are freed from your disability."
LUKE|13|13|And he laid his hands on her, and immediately she was made straight, and she glorified God.
LUKE|13|14|But the ruler of the synagogue, indignant because Jesus had healed on the Sabbath, said to the people, "There are six days in which work ought to be done. Come on those days and be healed, and not on the Sabbath day."
LUKE|13|15|Then the Lord answered him, "You hypocrites! Does not each of you on the Sabbath untie his ox or his donkey from the manger and lead it away to water it?
LUKE|13|16|And ought not this woman, a daughter of Abraham whom Satan bound for eighteen years, be loosed from this bond on the Sabbath day?"
LUKE|13|17|As he said these things, all his adversaries were put to shame, and all the people rejoiced at all the glorious things that were done by him.
LUKE|13|18|He said therefore, "What is the kingdom of God like? And to what shall I compare it?
LUKE|13|19|It is like a grain of mustard seed that a man took and sowed in his garden, and it grew and became a tree, and the birds of the air made nests in its branches."
LUKE|13|20|And again he said, "To what shall I compare the kingdom of God?
LUKE|13|21|It is like leaven that a woman took and hid in three measures of flour, until it was all leavened."
LUKE|13|22|He went on his way through towns and villages, teaching and journeying toward Jerusalem.
LUKE|13|23|And someone said to him, "Lord, will those who are saved be few?" And he said to them,
LUKE|13|24|"Strive to enter through the narrow door. For many, I tell you, will seek to enter and will not be able.
LUKE|13|25|When once the master of the house has risen and shut the door, and you begin to stand outside and to knock at the door, saying, 'Lord, open to us,' then he will answer you, 'I do not know where you come from.'
LUKE|13|26|Then you will begin to say, 'We ate and drank in your presence, and you taught in our streets.'
LUKE|13|27|But he will say, 'I tell you, I do not know where you come from. Depart from me, all you workers of evil!'
LUKE|13|28|In that place there will be weeping and gnashing of teeth, when you see Abraham and Isaac and Jacob and all the prophets in the kingdom of God but you yourselves cast out.
LUKE|13|29|And people will come from east and west, and from north and south, and recline at table in the kingdom of God.
LUKE|13|30|And behold, some are last who will be first, and some are first who will be last."
LUKE|13|31|At that very hour some Pharisees came and said to him, "Get away from here, for Herod wants to kill you."
LUKE|13|32|And he said to them, "Go and tell that fox, 'Behold, I cast out demons and perform cures today and tomorrow, and the third day I finish my course.
LUKE|13|33|Nevertheless, I must go on my way today and tomorrow and the day following, for it cannot be that a prophet should perish away from Jerusalem.'
LUKE|13|34|O Jerusalem, Jerusalem, the city that kills the prophets and stones those who are sent to it! How often would I have gathered your children together as a hen gathers her brood under her wings, and you would not!
LUKE|13|35|Behold, your house is forsaken. And I tell you, you will not see me until you say, 'Blessed is he who comes in the name of the Lord!'"
LUKE|14|1|One Sabbath, when he went to dine at the house of a ruler of the Pharisees, they were watching him carefully.
LUKE|14|2|And behold, there was a man before him who had dropsy.
LUKE|14|3|And Jesus responded to the lawyers and Pharisees, saying, "Is it lawful to heal on the Sabbath, or not?"
LUKE|14|4|But they remained silent. Then he took him and healed him and sent him away.
LUKE|14|5|And he said to them, "Which of you, having a son or an ox that has fallen into a well on a Sabbath day, will not immediately pull him out?"
LUKE|14|6|And they could not reply to these things.
LUKE|14|7|Now he told a parable to those who were invited, when he noticed how they chose the places of honor, saying to them,
LUKE|14|8|"When you are invited by someone to a wedding feast, do not sit down in a place of honor, lest someone more distinguished than you be invited by him,
LUKE|14|9|and he who invited you both will come and say to you, 'Give your place to this person,' and then you will begin with shame to take the lowest place.
LUKE|14|10|But when you are invited, go and sit in the lowest place, so that when your host comes he may say to you, 'Friend, move up higher.' Then you will be honored in the presence of all who sit at table with you.
LUKE|14|11|For everyone who exalts himself will be humbled, and he who humbles himself will be exalted."
LUKE|14|12|He said also to the man who had invited him, "When you give a dinner or a banquet, do not invite your friends or your brothers or your relatives or rich neighbors, lest they also invite you in return and you be repaid.
LUKE|14|13|But when you give a feast, invite the poor, the crippled, the lame, the blind,
LUKE|14|14|and you will be blessed, because they cannot repay you. You will be repaid at the resurrection of the just."
LUKE|14|15|When one of those who reclined at table with him heard these things, he said to him, "Blessed is everyone who will eat bread in the kingdom of God!"
LUKE|14|16|But he said to him, "A man once gave a great banquet and invited many.
LUKE|14|17|And at the time for the banquet he sent his servant to say to those who had been invited, 'Come, for everything is now ready.'
LUKE|14|18|But they all alike began to make excuses. The first said to him, 'I have bought a field, and I must go out and see it. Please have me excused.'
LUKE|14|19|And another said, 'I have bought five yoke of oxen, and I go to examine them. Please have me excused.'
LUKE|14|20|And another said, 'I have married a wife, and therefore I cannot come.'
LUKE|14|21|So the servant came and reported these things to his master. Then the master of the house became angry and said to his servant, 'Go out quickly to the streets and lanes of the city, and bring in the poor and crippled and blind and lame.'
LUKE|14|22|And the servant said, 'Sir, what you commanded has been done, and still there is room.'
LUKE|14|23|And the master said to the servant, 'Go out to the highways and hedges and compel people to come in, that my house may be filled.
LUKE|14|24|For I tell you, none of those men who were invited shall taste my banquet.'"
LUKE|14|25|Now great crowds accompanied him, and he turned and said to them,
LUKE|14|26|"If anyone comes to me and does not hate his own father and mother and wife and children and brothers and sisters, yes, and even his own life, he cannot be my disciple.
LUKE|14|27|Whoever does not bear his own cross and come after me cannot be my disciple.
LUKE|14|28|For which of you, desiring to build a tower, does not first sit down and count the cost, whether he has enough to complete it?
LUKE|14|29|Otherwise, when he has laid a foundation and is not able to finish, all who see it begin to mock him,
LUKE|14|30|saying, 'This man began to build and was not able to finish.'
LUKE|14|31|Or what king, going out to encounter another king in war, will not sit down first and deliberate whether he is able with ten thousand to meet him who comes against him with twenty thousand?
LUKE|14|32|And if not, while the other is yet a great way off, he sends a delegation and asks for terms of peace.
LUKE|14|33|So therefore, any one of you who does not renounce all that he has cannot be my disciple.
LUKE|14|34|"Salt is good, but if salt has lost its taste, how shall its saltiness be restored?
LUKE|14|35|It is of no use either for the soil or for the manure pile. It is thrown away. He who has ears to hear, let him hear."
LUKE|15|1|Now the tax collectors and sinners were all drawing near to hear him.
LUKE|15|2|And the Pharisees and the scribes grumbled, saying, "This man receives sinners and eats with them."
LUKE|15|3|So he told them this parable:
LUKE|15|4|"What man of you, having a hundred sheep, if he has lost one of them, does not leave the ninety-nine in the open country, and go after the one that is lost, until he finds it?
LUKE|15|5|And when he has found it, he lays it on his shoulders, rejoicing.
LUKE|15|6|And when he comes home, he calls together his friends and his neighbors, saying to them, 'Rejoice with me, for I have found my sheep that was lost.'
LUKE|15|7|Just so, I tell you, there will be more joy in heaven over one sinner who repents than over ninety-nine righteous persons who need no repentance.
LUKE|15|8|"Or what woman, having ten silver coins, if she loses one coin, does not light a lamp and sweep the house and seek diligently until she finds it?
LUKE|15|9|And when she has found it, she calls together her friends and neighbors, saying, 'Rejoice with me, for I have found the coin that I had lost.'
LUKE|15|10|Just so, I tell you, there is joy before the angels of God over one sinner who repents."
LUKE|15|11|And he said, "There was a man who had two sons.
LUKE|15|12|And the younger of them said to his father, 'Father, give me the share of property that is coming to me.' And he divided his property between them.
LUKE|15|13|Not many days later, the younger son gathered all he had and took a journey into a far country, and there he squandered his property in reckless living.
LUKE|15|14|And when he had spent everything, a severe famine arose in that country, and he began to be in need.
LUKE|15|15|So he went and hired himself out to one of the citizens of that country, who sent him into his fields to feed pigs.
LUKE|15|16|And he was longing to be fed with the pods that the pigs ate, and no one gave him anything.
LUKE|15|17|"But when he came to himself, he said, 'How many of my father's hired servants have more than enough bread, but I perish here with hunger!
LUKE|15|18|I will arise and go to my father, and I will say to him, "Father, I have sinned against heaven and before you.
LUKE|15|19|I am no longer worthy to be called your son. Treat me as one of your hired servants."'
LUKE|15|20|And he arose and came to his father. But while he was still a long way off, his father saw him and felt compassion, and ran and embraced him and kissed him.
LUKE|15|21|And the son said to him, 'Father, I have sinned against heaven and before you. I am no longer worthy to be called your son.'
LUKE|15|22|But the father said to his servants, 'Bring quickly the best robe, and put it on him, and put a ring on his hand, and shoes on his feet.
LUKE|15|23|And bring the fattened calf and kill it, and let us eat and celebrate.
LUKE|15|24|For this my son was dead, and is alive again; he was lost, and is found.' And they began to celebrate.
LUKE|15|25|"Now his older son was in the field, and as he came and drew near to the house, he heard music and dancing.
LUKE|15|26|And he called one of the servants and asked what these things meant.
LUKE|15|27|And he said to him, 'Your brother has come, and your father has killed the fattened calf, because he has received him back safe and sound.'
LUKE|15|28|But he was angry and refused to go in. His father came out and entreated him,
LUKE|15|29|but he answered his father, 'Look, these many years I have served you, and I never disobeyed your command, yet you never gave me a young goat, that I might celebrate with my friends.
LUKE|15|30|But when this son of yours came, who has devoured your property with prostitutes, you killed the fattened calf for him!'
LUKE|15|31|And he said to him, 'Son, you are always with me, and all that is mine is yours.
LUKE|15|32|It was fitting to celebrate and be glad, for this your brother was dead, and is alive; he was lost, and is found.'"
LUKE|16|1|He also said to the disciples, "There was a rich man who had a manager, and charges were brought to him that this man was wasting his possessions.
LUKE|16|2|And he called him and said to him, 'What is this that I hear about you? Turn in the account of your management, for you can no longer be manager.'
LUKE|16|3|And the manager said to himself, 'What shall I do, since my master is taking the management away from me? I am not strong enough to dig, and I am ashamed to beg.
LUKE|16|4|I have decided what to do, so that when I am removed from management, people may receive me into their houses.'
LUKE|16|5|So, summoning his master's debtors one by one, he said to the first, 'How much do you owe my master?'
LUKE|16|6|He said, 'A hundred measures of oil.' He said to him, 'Take your bill, and sit down quickly and write fifty.'
LUKE|16|7|Then he said to another, 'And how much do you owe?' He said, 'A hundred measures of wheat.' He said to him, 'Take your bill, and write eighty.'
LUKE|16|8|The master commended the dishonest manager for his shrewdness. For the sons of this world are more shrewd in dealing with their own generation than the sons of light.
LUKE|16|9|And I tell you, make friends for yourselves by means of unrighteous wealth, so that when it fails they may receive you into the eternal dwellings.
LUKE|16|10|"One who is faithful in a very little is also faithful in much, and one who is dishonest in a very little is also dishonest in much.
LUKE|16|11|If then you have not been faithful in the unrighteous wealth, who will entrust to you the true riches?
LUKE|16|12|And if you have not been faithful in that which is another's, who will give you that which is your own?
LUKE|16|13|No servant can serve two masters, for either he will hate the one and love the other, or he will be devoted to the one and despise the other. You cannot serve God and money."
LUKE|16|14|The Pharisees, who were lovers of money, heard all these things, and they ridiculed him.
LUKE|16|15|And he said to them, "You are those who justify yourselves before men, but God knows your hearts. For what is exalted among men is an abomination in the sight of God.
LUKE|16|16|"The Law and the Prophets were until John; since then the good news of the kingdom of God is preached, and everyone forces his way into it.
LUKE|16|17|But it is easier for heaven and earth to pass away than for one dot of the Law to become void.
LUKE|16|18|"Everyone who divorces his wife and marries another commits adultery, and he who marries a woman divorced from her husband commits adultery.
LUKE|16|19|"There was a rich man who was clothed in purple and fine linen and who feasted sumptuously every day.
LUKE|16|20|And at his gate was laid a poor man named Lazarus, covered with sores,
LUKE|16|21|who desired to be fed with what fell from the rich man's table. Moreover, even the dogs came and licked his sores.
LUKE|16|22|The poor man died and was carried by the angels to Abraham's side. The rich man also died and was buried,
LUKE|16|23|and in Hades, being in torment, he lifted up his eyes and saw Abraham far off and Lazarus at his side.
LUKE|16|24|And he called out, 'Father Abraham, have mercy on me, and send Lazarus to dip the end of his finger in water and cool my tongue, for I am in anguish in this flame.'
LUKE|16|25|But Abraham said, 'Child, remember that you in your lifetime received your good things, and Lazarus in like manner bad things; but now he is comforted here, and you are in anguish.
LUKE|16|26|And besides all this, between us and you a great chasm has been fixed, in order that those who would pass from here to you may not be able, and none may cross from there to us.'
LUKE|16|27|And he said, 'Then I beg you, father, to send him to my father's house-
LUKE|16|28|for I have five brothers- so that he may warn them, lest they also come into this place of torment.'
LUKE|16|29|But Abraham said, 'They have Moses and the Prophets; let them hear them.'
LUKE|16|30|And he said, 'No, father Abraham, but if someone goes to them from the dead, they will repent.'
LUKE|16|31|He said to him, 'If they do not hear Moses and the Prophets, neither will they be convinced if someone should rise from the dead.'"
LUKE|17|1|And he said to his disciples, "Temptations to sin are sure to come, but woe to the one through whom they come!
LUKE|17|2|It would be better for him if a millstone were hung around his neck and he were cast into the sea than that he should cause one of these little ones to sin.
LUKE|17|3|Pay attention to yourselves! If your brother sins, rebuke him, and if he repents, forgive him,
LUKE|17|4|and if he sins against you seven times in the day, and turns to you seven times, saying, 'I repent,' you must forgive him."
LUKE|17|5|The apostles said to the Lord, "Increase our faith!"
LUKE|17|6|And the Lord said, "If you had faith like a grain of mustard seed, you could say to this mulberry tree, 'Be uprooted and planted in the sea,' and it would obey you.
LUKE|17|7|"Will any one of you who has a servant plowing or keeping sheep say to him when he has come in from the field, 'Come at once and sit down at table'?
LUKE|17|8|Will he not rather say to him, 'Prepare supper for me, and dress properly, and serve me while I eat and drink, and afterward you will eat and drink'?
LUKE|17|9|Does he thank the servant because he did what was commanded?
LUKE|17|10|So you also, when you have done all that you were commanded, say, 'We are unworthy servants; we have only done what was our duty.'"
LUKE|17|11|On the way to Jerusalem he was passing along between Samaria and Galilee.
LUKE|17|12|And as he entered a village, he was met by ten lepers, who stood at a distance
LUKE|17|13|and lifted up their voices, saying, "Jesus, Master, have mercy on us."
LUKE|17|14|When he saw them he said to them, "Go and show yourselves to the priests." And as they went they were cleansed.
LUKE|17|15|Then one of them, when he saw that he was healed, turned back, praising God with a loud voice;
LUKE|17|16|and he fell on his face at Jesus' feet, giving him thanks. Now he was a Samaritan.
LUKE|17|17|Then Jesus answered, "Were not ten cleansed? Where are the nine?
LUKE|17|18|Was no one found to return and give praise to God except this foreigner?"
LUKE|17|19|And he said to him, "Rise and go your way; your faith has made you well."
LUKE|17|20|Being asked by the Pharisees when the kingdom of God would come, he answered them, "The kingdom of God is not coming with signs to be observed,
LUKE|17|21|nor will they say, 'Look, here it is!' or 'There!' for behold, the kingdom of God is in the midst of you."
LUKE|17|22|And he said to the disciples, "The days are coming when you will desire to see one of the days of the Son of Man, and you will not see it.
LUKE|17|23|And they will say to you, 'Look, there!' or 'Look, here!' Do not go out or follow them.
LUKE|17|24|For as the lightning flashes and lights up the sky from one side to the other, so will the Son of Man be in his day.
LUKE|17|25|But first he must suffer many things and be rejected by this generation.
LUKE|17|26|Just as it was in the days of Noah, so will it be in the days of the Son of Man.
LUKE|17|27|They were eating and drinking and marrying and being given in marriage, until the day when Noah entered the ark, and the flood came and destroyed them all.
LUKE|17|28|Likewise, just as it was in the days of Lot- they were eating and drinking, buying and selling, planting and building,
LUKE|17|29|but on the day when Lot went out from Sodom, fire and sulfur rained from heaven and destroyed them all-
LUKE|17|30|so will it be on the day when the Son of Man is revealed.
LUKE|17|31|On that day, let the one who is on the housetop, with his goods in the house, not come down to take them away, and likewise let the one who is in the field not turn back.
LUKE|17|32|Remember Lot's wife.
LUKE|17|33|Whoever seeks to preserve his life will lose it, but whoever loses his life will keep it.
LUKE|17|34|I tell you, in that night there will be two in one bed. One will be taken and the other left.
LUKE|17|35|There will be two women grinding together. One will be taken and the other left."
LUKE|17|36|***
LUKE|17|37|And they said to him, "Where, Lord?" He said to them, "Where the corpse is, there the vultures will gather."
LUKE|18|1|And he told them a parable to the effect that they ought always to pray and not lose heart.
LUKE|18|2|He said, "In a certain city there was a judge who neither feared God nor respected man.
LUKE|18|3|And there was a widow in that city who kept coming to him and saying, 'Give me justice against my adversary.'
LUKE|18|4|For a while he refused, but afterward he said to himself, 'Though I neither fear God nor respect man,
LUKE|18|5|yet because this widow keeps bothering me, I will give her justice, so that she will not beat me down by her continual coming.'"
LUKE|18|6|And the Lord said, "Hear what the unrighteous judge says.
LUKE|18|7|And will not God give justice to his elect, who cry to him day and night? Will he delay long over them?
LUKE|18|8|I tell you, he will give justice to them speedily. Nevertheless, when the Son of Man comes, will he find faith on earth?"
LUKE|18|9|He also told this parable to some who trusted in themselves that they were righteous, and treated others with contempt:
LUKE|18|10|"Two men went up into the temple to pray, one a Pharisee and the other a tax collector.
LUKE|18|11|The Pharisee, standing by himself, prayed thus: 'God, I thank you that I am not like other men, extortioners, unjust, adulterers, or even like this tax collector.
LUKE|18|12|I fast twice a week; I give tithes of all that I get.'
LUKE|18|13|But the tax collector, standing far off, would not even lift up his eyes to heaven, but beat his breast, saying, 'God, be merciful to me, a sinner!'
LUKE|18|14|I tell you, this man went down to his house justified, rather than the other. For everyone who exalts himself will be humbled, but the one who humbles himself will be exalted."
LUKE|18|15|Now they were bringing even infants to him that he might touch them. And when the disciples saw it, they rebuked them.
LUKE|18|16|But Jesus called them to him, saying, "Let the children come to me, and do not hinder them, for to such belongs the kingdom of God.
LUKE|18|17|Truly, I say to you, whoever does not receive the kingdom of God like a child shall not enter it."
LUKE|18|18|And a ruler asked him, "Good Teacher, what must I do to inherit eternal life?"
LUKE|18|19|And Jesus said to him, "Why do you call me good? No one is good except God alone.
LUKE|18|20|You know the commandments: 'Do not commit adultery, Do not murder, Do not steal, Do not bear false witness, Honor your father and mother.'"
LUKE|18|21|And he said, "All these I have kept from my youth."
LUKE|18|22|When Jesus heard this, he said to him, "One thing you still lack. Sell all that you have and distribute to the poor, and you will have treasure in heaven; and come, follow me."
LUKE|18|23|But when he heard these things, he became very sad, for he was extremely rich.
LUKE|18|24|Jesus, looking at him with sadness, said, "How difficult it is for those who have wealth to enter the kingdom of God!
LUKE|18|25|For it is easier for a camel to go through the eye of a needle than for a rich person to enter the kingdom of God."
LUKE|18|26|Those who heard it said, "Then who can be saved?"
LUKE|18|27|But he said, "What is impossible with men is possible with God."
LUKE|18|28|And Peter said, "See, we have left our homes and followed you."
LUKE|18|29|And he said to them, "Truly, I say to you, there is no one who has left house or wife or brothers or parents or children, for the sake of the kingdom of God,
LUKE|18|30|who will not receive many times more in this time, and in the age to come eternal life."
LUKE|18|31|And taking the twelve, he said to them, "See, we are going up to Jerusalem, and everything that is written about the Son of Man by the prophets will be accomplished.
LUKE|18|32|For he will be delivered over to the Gentiles and will be mocked and shamefully treated and spit upon.
LUKE|18|33|And after flogging him, they will kill him, and on the third day he will rise."
LUKE|18|34|But they understood none of these things. This saying was hidden from them, and they did not grasp what was said.
LUKE|18|35|As he drew near to Jericho, a blind man was sitting by the roadside begging.
LUKE|18|36|And hearing a crowd going by, he inquired what this meant.
LUKE|18|37|They told him, "Jesus of Nazareth is passing by."
LUKE|18|38|And he cried out, "Jesus, Son of David, have mercy on me!"
LUKE|18|39|And those who were in front rebuked him, telling him to be silent. But he cried out all the more, "Son of David, have mercy on me!"
LUKE|18|40|And Jesus stopped and commanded him to be brought to him. And when he came near, he asked him,
LUKE|18|41|"What do you want me to do for you?" He said, "Lord, let me recover my sight."
LUKE|18|42|And Jesus said to him, "Recover your sight; your faith has made you well."
LUKE|18|43|And immediately he recovered his sight and followed him, glorifying God. And all the people, when they saw it, gave praise to God.
LUKE|19|1|He entered Jericho and was passing through.
LUKE|19|2|And there was a man named Zacchaeus. He was a chief tax collector and was rich.
LUKE|19|3|And he was seeking to see who Jesus was, but on account of the crowd he could not, because he was small of stature.
LUKE|19|4|So he ran on ahead and climbed up into a sycamore tree to see him, for he was about to pass that way.
LUKE|19|5|And when Jesus came to the place, he looked up and said to him, "Zacchaeus, hurry and come down, for I must stay at your house today."
LUKE|19|6|So he hurried and came down and received him joyfully.
LUKE|19|7|And when they saw it, they all grumbled, "He has gone in to be the guest of a man who is a sinner."
LUKE|19|8|And Zacchaeus stood and said to the Lord, "Behold, Lord, the half of my goods I give to the poor. And if I have defrauded anyone of anything, I restore it fourfold."
LUKE|19|9|And Jesus said to him, "Today salvation has come to this house, since he also is a son of Abraham.
LUKE|19|10|For the Son of Man came to seek and to save the lost."
LUKE|19|11|As they heard these things, he proceeded to tell a parable, because he was near to Jerusalem, and because they supposed that the kingdom of God was to appear immediately.
LUKE|19|12|He said therefore, "A nobleman went into a far country to receive for himself a kingdom and then return.
LUKE|19|13|Calling ten of his servants, he gave them ten minas, and said to them, 'Engage in business until I come.'
LUKE|19|14|But his citizens hated him and sent a delegation after him, saying, 'We do not want this man to reign over us.'
LUKE|19|15|When he returned, having received the kingdom, he ordered these servants to whom he had given the money to be called to him, that he might know what they had gained by doing business.
LUKE|19|16|The first came before him, saying, 'Lord, your mina has made ten minas more.'
LUKE|19|17|And he said to him, 'Well done, good servant! Because you have been faithful in a very little, you shall have authority over ten cities.'
LUKE|19|18|And the second came, saying, 'Lord, your mina has made five minas.'
LUKE|19|19|And he said to him, 'And you are to be over five cities.'
LUKE|19|20|Then another came, saying, 'Lord, here is your mina, which I kept laid away in a handkerchief;
LUKE|19|21|for I was afraid of you, because you are a severe man. You take what you did not deposit, and reap what you did not sow.'
LUKE|19|22|He said to him, 'I will condemn you with your own words, you wicked servant! You knew that I was a severe man, taking what I did not deposit and reaping what I did not sow?
LUKE|19|23|Why then did you not put my money in the bank, and at my coming I might have collected it with interest?'
LUKE|19|24|And he said to those who stood by, 'Take the mina from him, and give it to the one who has the ten minas.'
LUKE|19|25|And they said to him, 'Lord, he has ten minas!'
LUKE|19|26|'I tell you that to everyone who has, more will be given, but from the one who has not, even what he has will be taken away.
LUKE|19|27|But as for these enemies of mine, who did not want me to reign over them, bring them here and slaughter them before me.'"
LUKE|19|28|And when he had said these things, he went on ahead, going up to Jerusalem.
LUKE|19|29|When he drew near to Bethphage and Bethany, at the mount that is called Olivet, he sent two of the disciples,
LUKE|19|30|saying, "Go into the village in front of you, where on entering you will find a colt tied, on which no one has ever yet sat. Untie it and bring it here.
LUKE|19|31|If anyone asks you, 'Why are you untying it?' you shall say this: 'The Lord has need of it.'"
LUKE|19|32|So those who were sent went away and found it just as he had told them.
LUKE|19|33|And as they were untying the colt, its owners said to them, "Why are you untying the colt?"
LUKE|19|34|And they said, "The Lord has need of it."
LUKE|19|35|And they brought it to Jesus, and throwing their cloaks on the colt, they set Jesus on it.
LUKE|19|36|And as he rode along, they spread their cloaks on the road.
LUKE|19|37|As he was drawing near- already on the way down the Mount of Olives- the whole multitude of his disciples began to rejoice and praise God with a loud voice for all the mighty works that they had seen,
LUKE|19|38|saying, "Blessed is the King who comes in the name of the Lord! Peace in heaven and glory in the highest!"
LUKE|19|39|And some of the Pharisees in the crowd said to him, "Teacher, rebuke your disciples."
LUKE|19|40|He answered, "I tell you, if these were silent, the very stones would cry out."
LUKE|19|41|And when he drew near and saw the city, he wept over it,
LUKE|19|42|saying, "Would that you, even you, had known on this day the things that make for peace! But now they are hidden from your eyes.
LUKE|19|43|For the days will come upon you, when your enemies will set up a barricade around you and surround you and hem you in on every side
LUKE|19|44|and tear you down to the ground, you and your children within you. And they will not leave one stone upon another in you, because you did not know the time of your visitation."
LUKE|19|45|And he entered the temple and began to drive out those who sold,
LUKE|19|46|saying to them, "It is written, 'My house shall be a house of prayer,' but you have made it a den of robbers."
LUKE|19|47|And he was teaching daily in the temple. The chief priests and the scribes and the principal men of the people were seeking to destroy him,
LUKE|19|48|but they did not find anything they could do, for all the people were hanging on his words.
LUKE|20|1|One day, as Jesus was teaching the people in the temple and preaching the gospel, the chief priests and the scribes with the elders came up
LUKE|20|2|and said to him, "Tell us by what authority you do these things, or who it is that gave you this authority."
LUKE|20|3|He answered them, "I also will ask you a question. Now tell me,
LUKE|20|4|Was the baptism of John from heaven or from man?"
LUKE|20|5|And they discussed it with one another, saying, "If we say, 'From heaven,' he will say, 'Why did you not believe him?'
LUKE|20|6|But if we say, 'From man,' all the people will stone us to death, for they are convinced that John was a prophet."
LUKE|20|7|So they answered that they did not know where it came from.
LUKE|20|8|And Jesus said to them, "Neither will I tell you by what authority I do these things."
LUKE|20|9|And he began to tell the people this parable: "A man planted a vineyard and let it out to tenants and went into another country for a long while.
LUKE|20|10|When the time came, he sent a servant to the tenants, so that they would give him some of the fruit of the vineyard. But the tenants beat him and sent him away empty-handed.
LUKE|20|11|And he sent another servant. But they also beat and treated him shamefully, and sent him away empty-handed.
LUKE|20|12|And he sent yet a third. This one also they wounded and cast out.
LUKE|20|13|Then the owner of the vineyard said, 'What shall I do? I will send my beloved son; perhaps they will respect him.'
LUKE|20|14|But when the tenants saw him, they said to themselves, 'This is the heir. Let us kill him, so that the inheritance may be ours.'
LUKE|20|15|And they threw him out of the vineyard and killed him. What then will the owner of the vineyard do to them?
LUKE|20|16|He will come and destroy those tenants and give the vineyard to others." When they heard this, they said, "Surely not!"
LUKE|20|17|But he looked directly at them and said, "What then is this that is written: "' The stone that the builders rejected has become the cornerstone'?
LUKE|20|18|Everyone who falls on that stone will be broken to pieces, and when it falls on anyone, it will crush him."
LUKE|20|19|The scribes and the chief priests sought to lay hands on him at that very hour, for they perceived that he had told this parable against them, but they feared the people.
LUKE|20|20|So they watched him and sent spies, who pretended to be sincere, that they might catch him in something he said, so as to deliver him up to the authority and jurisdiction of the governor.
LUKE|20|21|So they asked him, "Teacher, we know that you speak and teach rightly, and show no partiality, but truly teach the way of God.
LUKE|20|22|Is it lawful for us to give tribute to Caesar, or not?"
LUKE|20|23|But he perceived their craftiness, and said to them,
LUKE|20|24|"Show me a denarius. Whose likeness and inscription does it have?" They said, "Caesar's."
LUKE|20|25|He said to them, "Then render to Caesar the things that are Caesar's, and to God the things that are God's."
LUKE|20|26|And they were not able in the presence of the people to catch him in what he said, but marveling at his answer they became silent.
LUKE|20|27|There came to him some Sadducees, those who deny that there is a resurrection,
LUKE|20|28|and they asked him a question, saying, "Teacher, Moses wrote for us that if a man's brother dies, having a wife but no children, the man must take the widow and raise up offspring for his brother.
LUKE|20|29|Now there were seven brothers. The first took a wife, and died without children.
LUKE|20|30|And the second
LUKE|20|31|and the third took her, and likewise all seven left no children and died.
LUKE|20|32|Afterward the woman also died.
LUKE|20|33|In the resurrection, therefore, whose wife will the woman be? For the seven had her as wife."
LUKE|20|34|And Jesus said to them, "The sons of this age marry and are given in marriage,
LUKE|20|35|but those who are considered worthy to attain to that age and to the resurrection from the dead neither marry nor are given in marriage,
LUKE|20|36|for they cannot die anymore, because they are equal to angels and are sons of God, being sons of the resurrection.
LUKE|20|37|But that the dead are raised, even Moses showed, in the passage about the bush, where he calls the Lord the God of Abraham and the God of Isaac and the God of Jacob.
LUKE|20|38|Now he is not God of the dead, but of the living, for all live to him."
LUKE|20|39|Then some of the scribes answered, "Teacher, you have spoken well."
LUKE|20|40|For they no longer dared to ask him any question.
LUKE|20|41|But he said to them, "How can they say that the Christ is David's son?
LUKE|20|42|For David himself says in the Book of Psalms, "' The Lord said to my Lord, Sit at my right hand,
LUKE|20|43|until I make your enemies your footstool.'
LUKE|20|44|David thus calls him Lord, so how is he his son?"
LUKE|20|45|And in the hearing of all the people he said to his disciples,
LUKE|20|46|"Beware of the scribes, who like to walk around in long robes, and love greetings in the marketplaces and the best seats in the synagogues and the places of honor at feasts,
LUKE|20|47|who devour widows' houses and for a pretense make long prayers. They will receive the greater condemnation."
LUKE|21|1|Jesus looked up and saw the rich putting their gifts into the offering box,
LUKE|21|2|and he saw a poor widow put in two small copper coins.
LUKE|21|3|And he said, "Truly, I tell you, this poor widow has put in more than all of them.
LUKE|21|4|For they all contributed out of their abundance, but she out of her poverty put in all she had to live on."
LUKE|21|5|And while some were speaking of the temple, how it was adorned with noble stones and offerings, he said,
LUKE|21|6|"As for these things that you see, the days will come when there will not be left here one stone upon another that will not be thrown down."
LUKE|21|7|And they asked him, "Teacher, when will these things be, and what will be the sign when these things are about to take place?"
LUKE|21|8|And he said, "See that you are not led astray. For many will come in my name, saying, 'I am he!' and, 'The time is at hand!' Do not go after them.
LUKE|21|9|And when you hear of wars and tumults, do not be terrified, for these things must first take place, but the end will not be at once."
LUKE|21|10|Then he said to them, "Nation will rise against nation, and kingdom against kingdom.
LUKE|21|11|There will be great earthquakes, and in various places famines and pestilences. And there will be terrors and great signs from heaven.
LUKE|21|12|But before all this they will lay their hands on you and persecute you, delivering you up to the synagogues and prisons, and you will be brought before kings and governors for my name's sake.
LUKE|21|13|This will be your opportunity to bear witness.
LUKE|21|14|Settle it therefore in your minds not to meditate beforehand how to answer,
LUKE|21|15|for I will give you a mouth and wisdom, which none of your adversaries will be able to withstand or contradict.
LUKE|21|16|You will be delivered up even by parents and brothers and relatives and friends, and some of you they will put to death.
LUKE|21|17|You will be hated by all for my name's sake.
LUKE|21|18|But not a hair of your head will perish.
LUKE|21|19|By your endurance you will gain your lives.
LUKE|21|20|"But when you see Jerusalem surrounded by armies, then know that its desolation has come near.
LUKE|21|21|Then let those who are in Judea flee to the mountains, and let those who are inside the city depart, and let not those who are out in the country enter it,
LUKE|21|22|for these are days of vengeance, to fulfill all that is written.
LUKE|21|23|Alas for women who are pregnant and for those who are nursing infants in those days! For there will be great distress upon the earth and wrath against this people.
LUKE|21|24|They will fall by the edge of the sword and be led captive among all nations, and Jerusalem will be trampled underfoot by the Gentiles, until the times of the Gentiles are fulfilled.
LUKE|21|25|"And there will be signs in sun and moon and stars, and on the earth distress of nations in perplexity because of the roaring of the sea and the waves,
LUKE|21|26|people fainting with fear and with foreboding of what is coming on the world. For the powers of the heavens will be shaken.
LUKE|21|27|And then they will see the Son of Man coming in a cloud with power and great glory.
LUKE|21|28|Now when these things begin to take place, straighten up and raise your heads, because your redemption is drawing near."
LUKE|21|29|And he told them a parable: "Look at the fig tree, and all the trees.
LUKE|21|30|As soon as they come out in leaf, you see for yourselves and know that the summer is already near.
LUKE|21|31|So also, when you see these things taking place, you know that the kingdom of God is near.
LUKE|21|32|Truly, I say to you, this generation will not pass away until all has taken place.
LUKE|21|33|Heaven and earth will pass away, but my words will not pass away.
LUKE|21|34|"But watch yourselves lest your hearts be weighed down with dissipation and drunkenness and cares of this life, and that day come upon you suddenly like a trap.
LUKE|21|35|For it will come upon all who dwell on the face of the whole earth.
LUKE|21|36|But stay awake at all times, praying that you may have strength to escape all these things that are going to take place, and to stand before the Son of Man."
LUKE|21|37|And every day he was teaching in the temple, but at night he went out and lodged on the mount called Olivet.
LUKE|21|38|And early in the morning all the people came to him in the temple to hear him.
LUKE|22|1|Now the Feast of Unleavened Bread drew near, which is called the Passover.
LUKE|22|2|And the chief priests and the scribes were seeking how to put him to death, for they feared the people.
LUKE|22|3|Then Satan entered into Judas called Iscariot, who was of the number of the twelve.
LUKE|22|4|He went away and conferred with the chief priests and officers how he might betray him to them.
LUKE|22|5|And they were glad, and agreed to give him money.
LUKE|22|6|So he consented and sought an opportunity to betray him to them in the absence of a crowd.
LUKE|22|7|Then came the day of Unleavened Bread, on which the Passover lamb had to be sacrificed.
LUKE|22|8|So Jesus sent Peter and John, saying, "Go and prepare the Passover for us, that we may eat it."
LUKE|22|9|They said to him, "Where will you have us prepare it?"
LUKE|22|10|He said to them, "Behold, when you have entered the city, a man carrying a jar of water will meet you. Follow him into the house that he enters
LUKE|22|11|and tell the master of the house, 'The Teacher says to you, Where is the guest room, where I may eat the Passover with my disciples?'
LUKE|22|12|And he will show you a large upper room furnished; prepare it there."
LUKE|22|13|And they went and found it just as he had told them, and they prepared the Passover.
LUKE|22|14|And when the hour came, he reclined at table, and the apostles with him.
LUKE|22|15|And he said to them, "I have earnestly desired to eat this Passover with you before I suffer.
LUKE|22|16|For I tell you I will not eat it until it is fulfilled in the kingdom of God."
LUKE|22|17|And he took a cup, and when he had given thanks he said, "Take this, and divide it among yourselves.
LUKE|22|18|For I tell you that from now on I will not drink of the fruit of the vine until the kingdom of God comes."
LUKE|22|19|And he took bread, and when he had given thanks, he broke it and gave it to them, saying, "This is my body, which is given for you. Do this in remembrance of me."
LUKE|22|20|And likewise the cup after they had eaten, saying, "This cup that is poured out for you is the new covenant in my blood.
LUKE|22|21|But behold, the hand of him who betrays me is with me on the table.
LUKE|22|22|For the Son of Man goes as it has been determined, but woe to that man by whom he is betrayed!"
LUKE|22|23|And they began to question one another, which of them it could be who was going to do this.
LUKE|22|24|A dispute also arose among them, as to which of them was to be regarded as the greatest.
LUKE|22|25|And he said to them, "The kings of the Gentiles exercise lordship over them, and those in authority over them are called benefactors.
LUKE|22|26|But not so with you. Rather, let the greatest among you become as the youngest, and the leader as one who serves.
LUKE|22|27|For who is the greater, one who reclines at table or one who serves? Is it not the one who reclines at table? But I am among you as the one who serves.
LUKE|22|28|"You are those who have stayed with me in my trials,
LUKE|22|29|and I assign to you, as my Father assigned to me, a kingdom,
LUKE|22|30|that you may eat and drink at my table in my kingdom and sit on thrones judging the twelve tribes of Israel.
LUKE|22|31|"Simon, Simon, behold, Satan demanded to have you, that he might sift you like wheat,
LUKE|22|32|but I have prayed for you that your faith may not fail. And when you have turned again, strengthen your brothers."
LUKE|22|33|Peter said to him, "Lord, I am ready to go with you both to prison and to death."
LUKE|22|34|Jesus said, "I tell you, Peter, the rooster will not crow this day, until you deny three times that you know me."
LUKE|22|35|And he said to them, "When I sent you out with no moneybag or knapsack or sandals, did you lack anything?" They said, "Nothing."
LUKE|22|36|He said to them, "But now let the one who has a moneybag take it, and likewise a knapsack. And let the one who has no sword sell his cloak and buy one.
LUKE|22|37|For I tell you that this Scripture must be fulfilled in me: 'And he was numbered with the transgressors.' For what is written about me has its fulfillment."
LUKE|22|38|And they said, "Look, Lord, here are two swords." And he said to them, "It is enough."
LUKE|22|39|And he came out and went, as was his custom, to the Mount of Olives, and the disciples followed him.
LUKE|22|40|And when he came to the place, he said to them, "Pray that you may not enter into temptation."
LUKE|22|41|And he withdrew from them about a stone's throw, and knelt down and prayed,
LUKE|22|42|saying, "Father, if you are willing, remove this cup from me. Nevertheless, not my will, but yours, be done."
LUKE|22|43|And there appeared to him an angel from heaven, strengthening him.
LUKE|22|44|And being in an agony he prayed more earnestly; and his sweat became like great drops of blood falling down to the ground.
LUKE|22|45|And when he rose from prayer, he came to the disciples and found them sleeping for sorrow,
LUKE|22|46|and he said to them, "Why are you sleeping? Rise and pray that you may not enter into temptation."
LUKE|22|47|While he was still speaking, there came a crowd, and the man called Judas, one of the twelve, was leading them. He drew near to Jesus to kiss him,
LUKE|22|48|but Jesus said to him, "Judas, would you betray the Son of Man with a kiss?"
LUKE|22|49|And when those who were around him saw what would follow, they said, "Lord, shall we strike with the sword?"
LUKE|22|50|And one of them struck the servant of the high priest and cut off his right ear.
LUKE|22|51|But Jesus said, "No more of this!" And he touched his ear and healed him.
LUKE|22|52|Then Jesus said to the chief priests and officers of the temple and elders, who had come out against him, "Have you come out as against a robber, with swords and clubs?
LUKE|22|53|When I was with you day after day in the temple, you did not lay hands on me. But this is your hour, and the power of darkness."
LUKE|22|54|Then they seized him and led him away, bringing him into the high priest's house, and Peter was following at a distance.
LUKE|22|55|And when they had kindled a fire in the middle of the courtyard and sat down together, Peter sat down among them.
LUKE|22|56|Then a servant girl, seeing him as he sat in the light and looking closely at him, said, "This man also was with him."
LUKE|22|57|But he denied it, saying, "Woman, I do not know him."
LUKE|22|58|And a little later someone else saw him and said, "You also are one of them." But Peter said, "Man, I am not."
LUKE|22|59|And after an interval of about an hour still another insisted, saying, "Certainly this man also was with him, for he too is a Galilean."
LUKE|22|60|But Peter said, "Man, I do not know what you are talking about." And immediately, while he was still speaking, the rooster crowed.
LUKE|22|61|And the Lord turned and looked at Peter. And Peter remembered the saying of the Lord, how he had said to him, "Before the rooster crows today, you will deny me three times."
LUKE|22|62|And he went out and wept bitterly.
LUKE|22|63|Now the men who were holding Jesus in custody were mocking him as they beat him.
LUKE|22|64|They also blindfolded him and kept asking him, "Prophesy! Who is it that struck you?"
LUKE|22|65|And they said many other things against him, blaspheming him.
LUKE|22|66|When day came, the assembly of the elders of the people gathered together, both chief priests and scribes. And they led him away to their council, and they said,
LUKE|22|67|"If you are the Christ, tell us." But he said to them, "If I tell you, you will not believe,
LUKE|22|68|and if I ask you, you will not answer.
LUKE|22|69|But from now on the Son of Man shall be seated at the right hand of the power of God."
LUKE|22|70|So they all said, "Are you the Son of God, then?" And he said to them, "You say that I am."
LUKE|22|71|Then they said, "What further testimony do we need? We have heard it ourselves from his own lips."
LUKE|23|1|Then the whole company of them arose and brought him before Pilate.
LUKE|23|2|And they began to accuse him, saying, "We found this man misleading our nation and forbidding us to give tribute to Caesar, and saying that he himself is Christ, a king."
LUKE|23|3|And Pilate asked him, "Are you the King of the Jews?" And he answered him, "You have said so."
LUKE|23|4|Then Pilate said to the chief priests and the crowds, "I find no guilt in this man."
LUKE|23|5|But they were urgent, saying, "He stirs up the people, teaching throughout all Judea, from Galilee even to this place."
LUKE|23|6|When Pilate heard this, he asked whether the man was a Galilean.
LUKE|23|7|And when he learned that he belonged to Herod's jurisdiction, he sent him over to Herod, who was himself in Jerusalem at that time.
LUKE|23|8|When Herod saw Jesus, he was very glad, for he had long desired to see him, because he had heard about him, and he was hoping to see some sign done by him.
LUKE|23|9|So he questioned him at some length, but he made no answer.
LUKE|23|10|The chief priests and the scribes stood by, vehemently accusing him.
LUKE|23|11|And Herod with his soldiers treated him with contempt and mocked him. Then, arraying him in splendid clothing, he sent him back to Pilate.
LUKE|23|12|And Herod and Pilate became friends with each other that very day, for before this they had been at enmity with each other.
LUKE|23|13|Pilate then called together the chief priests and the rulers and the people,
LUKE|23|14|and said to them, "You brought me this man as one who was misleading the people. And after examining him before you, behold, I did not find this man guilty of any of your charges against him.
LUKE|23|15|Neither did Herod, for he sent him back to us. Look, nothing deserving death has been done by him.
LUKE|23|16|I will therefore punish and release him."
LUKE|23|17|***
LUKE|23|18|But they all cried out together, "Away with this man, and release to us Barabbas"-
LUKE|23|19|a man who had been thrown into prison for an insurrection started in the city and for murder.
LUKE|23|20|Pilate addressed them once more, desiring to release Jesus,
LUKE|23|21|but they kept shouting, "Crucify, crucify him!"
LUKE|23|22|A third time he said to them, "Why, what evil has he done? I have found in him no guilt deserving death. I will therefore punish and release him."
LUKE|23|23|But they were urgent, demanding with loud cries that he should be crucified. And their voices prevailed.
LUKE|23|24|So Pilate decided that their demand should be granted.
LUKE|23|25|He released the man who had been thrown into prison for insurrection and murder, for whom they asked, but he delivered Jesus over to their will.
LUKE|23|26|And as they led him away, they seized one Simon of Cyrene, who was coming in from the country, and laid on him the cross, to carry it behind Jesus.
LUKE|23|27|And there followed him a great multitude of the people and of women who were mourning and lamenting for him.
LUKE|23|28|But turning to them Jesus said, "Daughters of Jerusalem, do not weep for me, but weep for yourselves and for your children.
LUKE|23|29|For behold, the days are coming when they will say, 'Blessed are the barren and the wombs that never bore and the breasts that never nursed!'
LUKE|23|30|Then they will begin to say to the mountains, 'Fall on us,' and to the hills, 'Cover us.'
LUKE|23|31|For if they do these things when the wood is green, what will happen when it is dry?"
LUKE|23|32|Two others, who were criminals, were led away to be put to death with him.
LUKE|23|33|And when they came to the place that is called The Skull, there they crucified him, and the criminals, one on his right and one on his left.
LUKE|23|34|And Jesus said, "Father, forgive them, for they know not what they do." And they cast lots to divide his garments.
LUKE|23|35|And the people stood by, watching, but the rulers scoffed at him, saying, "He saved others; let him save himself, if he is the Christ of God, his Chosen One!"
LUKE|23|36|The soldiers also mocked him, coming up and offering him sour wine
LUKE|23|37|and saying, "If you are the King of the Jews, save yourself!"
LUKE|23|38|There was also an inscription over him, "This is the King of the Jews."
LUKE|23|39|One of the criminals who were hanged railed at him, saying, "Are you not the Christ? Save yourself and us!"
LUKE|23|40|But the other rebuked him, saying, "Do you not fear God, since you are under the same sentence of condemnation?
LUKE|23|41|And we indeed justly, for we are receiving the due reward of our deeds; but this man has done nothing wrong."
LUKE|23|42|And he said, "Jesus, remember me when you come into your kingdom."
LUKE|23|43|And he said to him, "Truly, I say to you, today you will be with me in Paradise."
LUKE|23|44|It was now about the sixth hour, and there was darkness over the whole land until the ninth hour,
LUKE|23|45|while the sun's light failed. And the curtain of the temple was torn in two.
LUKE|23|46|Then Jesus, calling out with a loud voice, said, "Father, into your hands I commit my spirit!" And having said this he breathed his last.
LUKE|23|47|Now when the centurion saw what had taken place, he praised God, saying, "Certainly this man was innocent!"
LUKE|23|48|And all the crowds that had assembled for this spectacle, when they saw what had taken place, returned home beating their breasts.
LUKE|23|49|And all his acquaintances and the women who had followed him from Galilee stood at a distance watching these things.
LUKE|23|50|Now there was a man named Joseph, from the Jewish town of Arimathea. He was a member of the council, a good and righteous man,
LUKE|23|51|who had not consented to their decision and action; and he was looking for the kingdom of God.
LUKE|23|52|This man went to Pilate and asked for the body of Jesus.
LUKE|23|53|Then he took it down and wrapped it in a linen shroud and laid him in a tomb cut in stone, where no one had ever yet been laid.
LUKE|23|54|It was the day of Preparation, and the Sabbath was beginning.
LUKE|23|55|The women who had come with him from Galilee followed and saw the tomb and how his body was laid.
LUKE|23|56|Then they returned and prepared spices and ointments. On the Sabbath they rested according to the commandment.
LUKE|24|1|But on the first day of the week, at early dawn, they went to the tomb, taking the spices they had prepared.
LUKE|24|2|And they found the stone rolled away from the tomb,
LUKE|24|3|but when they went in they did not find the body of the Lord Jesus.
LUKE|24|4|While they were perplexed about this, behold, two men stood by them in dazzling apparel.
LUKE|24|5|And as they were frightened and bowed their faces to the ground, the men said to them, "Why do you seek the living among the dead?
LUKE|24|6|He is not here, but has risen. Remember how he told you, while he was still in Galilee,
LUKE|24|7|that the Son of Man must be delivered into the hands of sinful men and be crucified and on the third day rise."
LUKE|24|8|And they remembered his words,
LUKE|24|9|and returning from the tomb they told all these things to the eleven and to all the rest.
LUKE|24|10|Now it was Mary Magdalene and Joanna and Mary the mother of James and the other women with them who told these things to the apostles,
LUKE|24|11|but these words seemed to them an idle tale, and they did not believe them.
LUKE|24|12|But Peter rose and ran to the tomb; stooping and looking in, he saw the linen cloths by themselves; and he went home marveling at what had happened.
LUKE|24|13|That very day two of them were going to a village named Emmaus, about seven miles from Jerusalem,
LUKE|24|14|and they were talking with each other about all these things that had happened.
LUKE|24|15|While they were talking and discussing together, Jesus himself drew near and went with them.
LUKE|24|16|But their eyes were kept from recognizing him.
LUKE|24|17|And he said to them, "What is this conversation that you are holding with each other as you walk?" And they stood still, looking sad.
LUKE|24|18|Then one of them, named Cleopas, answered him, "Are you the only visitor to Jerusalem who does not know the things that have happened there in these days?"
LUKE|24|19|And he said to them, "What things?" And they said to him, "Concerning Jesus of Nazareth, a man who was a prophet mighty in deed and word before God and all the people,
LUKE|24|20|and how our chief priests and rulers delivered him up to be condemned to death, and crucified him.
LUKE|24|21|But we had hoped that he was the one to redeem Israel. Yes, and besides all this, it is now the third day since these things happened.
LUKE|24|22|Moreover, some women of our company amazed us. They were at the tomb early in the morning,
LUKE|24|23|and when they did not find his body, they came back saying that they had even seen a vision of angels, who said that he was alive.
LUKE|24|24|Some of those who were with us went to the tomb and found it just as the women had said, but him they did not see."
LUKE|24|25|And he said to them, "O foolish ones, and slow of heart to believe all that the prophets have spoken!
LUKE|24|26|Was it not necessary that the Christ should suffer these things and enter into his glory?"
LUKE|24|27|And beginning with Moses and all the Prophets, he interpreted to them in all the Scriptures the things concerning himself.
LUKE|24|28|So they drew near to the village to which they were going. He acted as if he were going farther,
LUKE|24|29|but they urged him strongly, saying, "Stay with us, for it is toward evening and the day is now far spent." So he went in to stay with them.
LUKE|24|30|When he was at table with them, he took the bread and blessed and broke it and gave it to them.
LUKE|24|31|And their eyes were opened, and they recognized him. And he vanished from their sight.
LUKE|24|32|They said to each other, "Did not our hearts burn within us while he talked to us on the road, while he opened to us the Scriptures?"
LUKE|24|33|And they rose that same hour and returned to Jerusalem. And they found the eleven and those who were with them gathered together,
LUKE|24|34|saying, "The Lord has risen indeed, and has appeared to Simon!"
LUKE|24|35|Then they told what had happened on the road, and how he was known to them in the breaking of the bread.
LUKE|24|36|As they were talking about these things, Jesus himself stood among them, and said to them, "Peace to you!"
LUKE|24|37|But they were startled and frightened and thought they saw a spirit.
LUKE|24|38|And he said to them, "Why are you troubled, and why do doubts arise in your hearts?
LUKE|24|39|See my hands and my feet, that it is I myself. Touch me, and see. For a spirit does not have flesh and bones as you see that I have."
LUKE|24|40|And when he had said this, he showed them his hands and his feet.
LUKE|24|41|And while they still disbelieved for joy and were marveling, he said to them, "Have you anything here to eat?"
LUKE|24|42|They gave him a piece of broiled fish,
LUKE|24|43|and he took it and ate before them.
LUKE|24|44|Then he said to them, "These are my words that I spoke to you while I was still with you, that everything written about me in the Law of Moses and the Prophets and the Psalms must be fulfilled."
LUKE|24|45|Then he opened their minds to understand the Scriptures,
LUKE|24|46|and said to them, "Thus it is written, that the Christ should suffer and on the third day rise from the dead,
LUKE|24|47|and that repentance and forgiveness of sins should be proclaimed in his name to all nations, beginning from Jerusalem.
LUKE|24|48|You are witnesses of these things.
LUKE|24|49|And behold, I am sending the promise of my Father upon you. But stay in the city until you are clothed with power from on high."
LUKE|24|50|Then he led them out as far as Bethany, and lifting up his hands he blessed them.
LUKE|24|51|While he blessed them, he parted from them and was carried up into heaven.
LUKE|24|52|And they worshiped him and returned to Jerusalem with great joy,
LUKE|24|53|and were continually in the temple blessing God.
