GEN|1|1|起初，上帝创造天地。
GEN|1|2|地是空虚混沌，深渊上面一片黑暗；上帝的灵 运行在水面上。
GEN|1|3|上帝说：“要有光”，就有了光。
GEN|1|4|上帝看光是好的，于是上帝就把光和暗分开。
GEN|1|5|上帝称光为“昼”，称暗为“夜”。有晚上，有早晨，这是第一日。
GEN|1|6|上帝说：“众水之间要有穹苍，把水和水分开。”
GEN|1|7|上帝就造了穹苍，把穹苍以下的水和穹苍以上的水分开。事就这样成了。
GEN|1|8|上帝称穹苍为“天”。有晚上，有早晨，这是第二日。
GEN|1|9|上帝说：“天下面的水要聚集在一处，使干地露出来。”事就这样成了。
GEN|1|10|上帝称干地为“地”，称聚集在一起的水为“海”。上帝看为好的。
GEN|1|11|上帝说：“地要长出植物，就是含种子的五谷菜蔬，和会结果子、果子里有种子的树，在地上各从其类。”事就这样成了。
GEN|1|12|于是地长出了植物：含种子的五谷菜蔬，各从其类；会结果子、果子里有种子的树，各从其类。上帝看为好的。
GEN|1|13|有晚上，有早晨，这是第三日。
GEN|1|14|上帝说：“天上要有光体来分昼夜，让它们作记号，定季节、日子、年份，
GEN|1|15|它们要在天空发光，照在地上。”事就这样成了。
GEN|1|16|于是上帝造了两个大光体，大的管昼，小的管夜，又造了星辰。
GEN|1|17|上帝把这些光体摆列在天空，照在地上，
GEN|1|18|管理昼夜，分别光暗。上帝看为好的。
GEN|1|19|有晚上，有早晨，这是第四日。
GEN|1|20|上帝说：“水要滋生众多有生命之物；要有鸟飞在地面以上，天空之中。”
GEN|1|21|上帝就创造了大鱼和在水里滋生的各样活动的生物，各从其类，以及各样有翅膀的鸟，各从其类。上帝看为好的。
GEN|1|22|上帝就赐福给这一切，说：“要繁殖增多，充满在海的水里；飞鸟也要在地上增多。”
GEN|1|23|有晚上，有早晨，这是第五日。
GEN|1|24|上帝说：“地要生出有生命之物，各从其类，就是牲畜、爬行动物、地上的走兽，各从其类。”事就这样成了。
GEN|1|25|于是上帝造了地上的走兽，各从其类；牲畜，各从其类；和地上一切的爬行动物，各从其类。上帝看为好的。
GEN|1|26|上帝说：“我们要照着我们的形像，按着我们的样式造人，使他们管理海里的鱼、天空的鸟、地上的牲畜和全地，以及地上爬的一切爬行动物。”
GEN|1|27|上帝就照着他的形像创造人，照着上帝的形像创造他们 ；他创造了他们，有男有女。
GEN|1|28|上帝赐福给他们，上帝对他们说：“要生养众多，遍满这地，治理它；要管理海里的鱼、天空的鸟和地上各样活动的生物。”
GEN|1|29|上帝说：“看哪，我把全地一切含种子的五谷菜蔬和一切会结果子、果子里有种子的树，都赐给你们；这些都可作食物。
GEN|1|30|至于地上一切的走兽、天空一切的飞鸟，并一切在地上爬行的，有生命的动物，我把绿色植物赐给它们作食物。”事就这样成了。
GEN|1|31|上帝看一切所造的，看哪，都非常好。有晚上，有早晨，这是第六日。
GEN|2|1|天和地，以及万象都完成了。
GEN|2|2|到第七日，上帝已经完成了造物之工，就在第七日安息了，歇了他所做一切的工。
GEN|2|3|上帝赐福给第七日，将它分别为圣，因为在这日，上帝安息了，歇了他所做一切创造的工。
GEN|2|4|这就是天地创造的来历。 在耶和华上帝造地和天的时候，
GEN|2|5|地上还没有田野的草木，田间的菜蔬还没有长出来，因为耶和华上帝还没有降雨在地上，也没有人耕种土地。
GEN|2|6|但是，有雾气从地上腾，滋润整个土地的表面。
GEN|2|7|耶和华上帝用地上的尘土造人，将生命之气吹进他的鼻孔，这人就成了有灵的活人 。
GEN|2|8|耶和华上帝在东方的 伊甸 栽了一个园子，把所造的人安置在那里。
GEN|2|9|耶和华上帝使各样的树从土地里长出来，可以悦人的眼目，好作食物。园子当中有生命树和知善恶的树 。
GEN|2|10|有一条河从 伊甸 流出来，滋润那园子，从那里分成四个源头：
GEN|2|11|第一条名叫 比逊 ，它环绕 哈腓拉 全地，在那里有金子。
GEN|2|12|那地的金子很好，在那里也有珍珠 和红玛瑙。
GEN|2|13|第二条河名叫 基训 ，它环绕 古实 全地。
GEN|2|14|第三条河名叫 底格里斯 ，它流到 亚述 的东边。第四条河就是 幼发拉底 。
GEN|2|15|耶和华上帝把那人安置在 伊甸园 ，让他耕耘看管。
GEN|2|16|耶和华上帝吩咐那人说：“园中各样树上所出的，你可以随意吃，
GEN|2|17|只是知善恶的树所出的，你不可吃，因为你吃它的日子必定死！”
GEN|2|18|耶和华上帝说：“那人单独一个不好，我要为他造一个配偶帮助他。”
GEN|2|19|耶和华上帝用泥土造了野地各样的走兽和天空各样的飞鸟，都带到那人面前，看他叫什么。那人怎样叫各样的动物，那就是它的名字。
GEN|2|20|那人就给一切牲畜、天空的飞鸟和野地各样的走兽都起了名。只是 亚当 没有找到配偶帮助他。
GEN|2|21|耶和华上帝使他沉睡，他就睡了；于是取下他的一根肋骨，又在原处把肉合起来。
GEN|2|22|耶和华上帝就用那人身上所取的肋骨造了一个女人，带她到那人面前。
GEN|2|23|那人说： “这正是我骨中的骨， 肉中的肉， 可以称她为女人， 因为她是从男人身上取出来的。”
GEN|2|24|因此，人要离开父母，与妻子结合，二人成为一体。
GEN|2|25|当时夫妻二人赤身露体，并不觉得羞耻。
GEN|3|1|耶和华上帝所造的，惟有蛇比田野一切的走兽更狡猾。蛇对女人说：“上帝岂是真说，你们不可吃园中任何树上所出的吗？”
GEN|3|2|女人对蛇说：“园中树上的果子，我们都可以吃；
GEN|3|3|只是园子中间那棵树的果子，上帝曾说：‘你们不可吃，也不可摸，免得你们死。’”
GEN|3|4|蛇对女人说：“你们不一定死；
GEN|3|5|因为上帝知道，你们吃的日子眼睛就开了，你们就像上帝一样知道善恶。”
GEN|3|6|于是女人见那棵树好作食物，又悦人的眼目，那树令人喜爱，能使人有智慧，她就摘下果子吃了，又给了与她一起的丈夫，他也吃了。
GEN|3|7|他们二人的眼睛就开了，知道自己赤身露体，就编织无花果树的叶子，为自己做成裙子。
GEN|3|8|天起了凉风，那人和他妻子听见耶和华上帝在园中来回行走的声音，就藏在园里的树木中，躲避耶和华上帝的面。
GEN|3|9|耶和华上帝呼唤那人，对他说：“你在哪里？”
GEN|3|10|他说：“我在园中听见你的声音，我就害怕；因为我赤身露体，我就藏了起来。”
GEN|3|11|耶和华上帝说：“谁告诉你，你是赤身露体呢？莫非你吃了那树上所出的，就是我吩咐你不可吃的吗？”
GEN|3|12|那人说：“你赐给我、与我一起的女人，是她把那树上所出的给我，我就吃了。”
GEN|3|13|耶和华上帝对女人说：“你怎么会做这种事呢？”女人说：“那蛇引诱我，我就吃了。”
GEN|3|14|耶和华上帝对蛇说： “你既做了这事，就必受诅咒， 比一切的牲畜和野兽更重。 你必用肚子行走， 终生吃土。
GEN|3|15|我要使你和女人彼此为仇， 你的后裔和女人的后裔也彼此为仇。 他要伤你的头， 你要伤他的脚跟。 ”
GEN|3|16|又对女人说： “我必多多加增你怀胎的痛苦， 你生儿女时必多受痛苦。 你必恋慕你丈夫， 他必管辖你。”
GEN|3|17|又对 亚当 说： “你既听从你妻子的话， 吃了那树上所出的， 就是我吩咐你不可吃的， 土地必因你的缘故受诅咒； 你必终生劳苦才能从土地得吃的。
GEN|3|18|土地必给你长出荆棘和蒺藜来； 你也要吃田间的五谷菜蔬。
GEN|3|19|你必汗流满面才有食物可吃， 直到你归了土地， 因为你是从土地而出的。 你本是尘土，仍要归回尘土。”
GEN|3|20|那人给他妻子起名叫 夏娃 ，因为她是众生之母 。
GEN|3|21|耶和华上帝用兽皮做衣服给 亚当 和他的妻子穿。
GEN|3|22|耶和华上帝说：“看哪，那人已经像我们中间的一个，知道善恶，现在恐怕他又伸手摘生命树所出的来吃，就永远活着。”
GEN|3|23|耶和华上帝就驱逐他出 伊甸园 ，使他耕种土地，他原是从土地里被取出来的。
GEN|3|24|耶和华上帝把那人赶出去，就在 伊甸园 东边安设基路伯和发出火焰转动的剑，把守生命树的道路。
GEN|4|1|那人和他妻子 夏娃 同房， 夏娃 就怀孕，生了 该隐 ，她说：“我靠耶和华得了一个男的。”
GEN|4|2|她又生了 该隐 的弟弟 亚伯 。 亚伯 是牧羊的； 该隐 是耕地的。
GEN|4|3|过了一些日子， 该隐 拿地里的出产为供物献给耶和华；
GEN|4|4|亚伯 也把他羊群中头生的和羊的脂肪献上。耶和华看中了 亚伯 和他的供物，
GEN|4|5|却看不中 该隐 和他的供物。 该隐 就非常生气，沉下脸来。
GEN|4|6|耶和华对 该隐 说：“你为什么生气呢？你为什么沉下脸来呢？
GEN|4|7|你若做得对，岂不仰起头来吗？你若做得不对，罪就伏在门前。它想要控制你，你却要制伏它。”
GEN|4|8|该隐 与他弟弟 亚伯 说话 。 二人正在田间时， 该隐 起来攻击他弟弟 亚伯 ，把他杀了。
GEN|4|9|耶和华对 该隐 说：“你弟弟 亚伯 在哪里？”他说：“我不知道！我岂是看守我弟弟的吗？”
GEN|4|10|耶和华说：“你做了什么事呢？你弟弟血的声音从地里向我哀号。
GEN|4|11|现在你必从这地受诅咒，这地开了口，从你手里接受你弟弟的血。
GEN|4|12|你耕种土地，它不再给你效力；你必流离飘荡在地上。”
GEN|4|13|该隐 对耶和华说：“我的惩罚太重，过于我所能承当的。
GEN|4|14|看哪，今日你赶我离开这块土地，不能见你的面；我必流离飘荡在地上，凡遇见我的必杀我。”
GEN|4|15|耶和华对他说：“既然如此 ，凡杀 该隐 的，必遭报七倍。”耶和华就给 该隐 立一个记号，免得人遇见他就杀他。
GEN|4|16|于是 该隐 离开了耶和华的面，去住在 伊甸 东边 挪得 之地。
GEN|4|17|该隐 与妻子同房，她就怀孕，生了 以诺 。 该隐 建造一座城，就照他儿子的名字称那城为 以诺 。
GEN|4|18|以诺 生 以拿 ， 以拿 生 米户雅利 ， 米户雅利 生 玛土撒利 ， 玛土撒利 生 拉麦 。
GEN|4|19|拉麦 娶了两个妻子：一个名叫 亚大 ，一个名叫 洗拉 。
GEN|4|20|亚大 生 雅八 ； 雅八 是住帐棚、牧养牲畜之人的祖师。
GEN|4|21|雅八 的兄弟名叫 犹八 ；他是所有弹琴吹箫之人的祖师。
GEN|4|22|洗拉 又生了 土八．该隐 ；他是打造各样铜器铁器的工匠。 土八．该隐 的妹妹是 拿玛 。
GEN|4|23|拉麦 对他两个妻子说： 亚大 、 洗拉 啊，听我的声音； 拉麦 的妻子啊，侧耳听我的言语： 大人伤我，我把他杀了； 小孩损我，我把他害了 。
GEN|4|24|若杀 该隐 ，遭报七倍， 杀 拉麦 的，必遭报七十七倍。
GEN|4|25|亚当 又与妻子同房，她就生了一个儿子，给他起名叫 塞特 ，说：“上帝给我立了另一个子嗣代替 亚伯 ，因为 该隐 杀了他。”
GEN|4|26|塞特 也生了一个儿子，起名叫 以挪士 。那时候，人开始求告耶和华的名。
GEN|5|1|这是 亚当 后代的家谱。当上帝造人的日子，他照着自己的样式造人。
GEN|5|2|他造男造女。在他们被造的日子，上帝赐福给他们，称他们为人。
GEN|5|3|亚当 活到一百三十岁，生了一个儿子，形像样式和自己相似，就给他起名叫 塞特 。
GEN|5|4|亚当 生 塞特 之后，又活了八百年，并且生儿育女。
GEN|5|5|亚当 共活了九百三十年，就死了。
GEN|5|6|塞特 活到一百零五岁，生了 以挪士 。
GEN|5|7|塞特 生 以挪士 之后，又活了八百零七年，并且生儿育女。
GEN|5|8|塞特 共活了九百一十二年，就死了。
GEN|5|9|以挪士 活到九十岁，生了 该南 。
GEN|5|10|以挪士 生 该南 之后，又活了八百一十五年，并且生儿育女。
GEN|5|11|以挪士 共活了九百零五年，就死了。
GEN|5|12|该南 活到七十岁，生了 玛勒列 。
GEN|5|13|该南 生 玛勒列 之后，又活了八百四十年，并且生儿育女。
GEN|5|14|该南 共活了九百一十年，就死了。
GEN|5|15|玛勒列 活到六十五岁，生了 雅列 。
GEN|5|16|玛勒列 生 雅列 之后，又活了八百三十年，并且生儿育女。
GEN|5|17|玛勒列 共活了八百九十五年，就死了。
GEN|5|18|雅列 活到一百六十二岁，生了 以诺 。
GEN|5|19|雅列 生 以诺 之后，又活了八百年，并且生儿育女。
GEN|5|20|雅列 共活了九百六十二年，就死了。
GEN|5|21|以诺 活到六十五岁，生了 玛土撒拉 。
GEN|5|22|以诺 生 玛土撒拉 之后，与上帝同行三百年，并且生儿育女。
GEN|5|23|以诺 共活了三百六十五年。
GEN|5|24|以诺 与上帝同行，上帝把他接去，他就不在了。
GEN|5|25|玛土撒拉 活到一百八十七岁，生了 拉麦 。
GEN|5|26|玛土撒拉 生 拉麦 之后，又活了七百八十二年，并且生儿育女。
GEN|5|27|玛土撒拉 共活了九百六十九年，就死了。
GEN|5|28|拉麦 活到一百八十二岁，生了一个儿子，
GEN|5|29|给他起名叫 挪亚 ，说：“在耶和华所诅咒的地上，这个儿子必使我们从工作和手中的劳苦得到安慰。”
GEN|5|30|拉麦 生 挪亚 之后，又活了五百九十五年，并且生儿育女。
GEN|5|31|拉麦 共活了七百七十七年，就死了。
GEN|5|32|挪亚 活到五百岁，生了 闪 、 含 和 雅弗 。
GEN|6|1|当人开始在地面上增多、又生女儿的时候，
GEN|6|2|上帝的儿子们看见人的女子美貌，就随意挑选，娶来为妻。
GEN|6|3|耶和华说：“人既属乎血气，我的灵就不永远住在他里面；然而他的年岁还可到一百二十年。”
GEN|6|4|那时候有巨人在地上，后来也有；上帝的儿子们和人的女子们交合，生了孩子。那些人就是古代的勇士，有名的人物。
GEN|6|5|耶和华见人在地上罪大恶极，终日心里所想的尽都是恶事，
GEN|6|6|耶和华就因造人在地上感到遗憾，心中忧伤。
GEN|6|7|耶和华说：“我要把所造的人和走兽，爬行动物，以及天空的飞鸟，都从地面上除灭，因为我造了他们感到遗憾。”
GEN|6|8|只有 挪亚 在耶和华眼前蒙恩。
GEN|6|9|这是 挪亚 的后代。 挪亚 是个义人，在他的世代中是个完全人。 挪亚 与上帝同行。
GEN|6|10|挪亚 生了三个儿子，就是 闪 、 含 和 雅弗 。
GEN|6|11|这地在上帝面前败坏了，地上充满了暴力。
GEN|6|12|上帝观看这地，看哪，它败坏了，因为凡血肉之躯在地上的行为都败坏了。
GEN|6|13|上帝对 挪亚 说：“在我面前，凡血肉之躯的结局已经临到，因着他们，地上充满了暴力。看哪，我要把他们和这地一起毁灭。
GEN|6|14|你要为自己用歌斐木造一艘方舟，并在方舟内造房间，内外都要抹上沥青。
GEN|6|15|方舟的造法是这样：要长三百肘，宽五十肘，高三十肘。
GEN|6|16|方舟上面要造天窗，向上一肘。方舟的门要开在旁边。方舟要分上、中、下三层。
GEN|6|17|看哪，我要使洪水泛滥在地上，毁灭天下凡有生命气息的血肉之躯，地上的一切都要灭亡。
GEN|6|18|但我要与你立约；你同你的儿子、妻子和媳妇都要进入方舟。
GEN|6|19|凡有血肉的动物，每样一对，一公一母，你要带进方舟，好跟你一起保全生命。
GEN|6|20|飞鸟各从其类，牲畜各从其类，地上的爬行动物各从其类，每样一对，都要到你那里，好保全生命。
GEN|6|21|你要拿各样可吃的食物，储存在你那里，作你和它们的粮食。”
GEN|6|22|挪亚 就去做了；凡上帝吩咐他的，他都照样去做。
GEN|7|1|耶和华对 挪亚 说：“你和你的全家都要进入方舟，因为在这世代中，我看你在我面前是个义人。
GEN|7|2|凡洁净的牲畜，你要各取七公七母；不洁净的牲畜，你要各取一公一母；
GEN|7|3|天空的飞鸟也要各取七公七母，为了要留种，活在全地面上。
GEN|7|4|因为再过七天，我要降雨在地上四十昼夜，把我所造的一切生物从地面上除灭。”
GEN|7|5|挪亚 就遵照耶和华吩咐他的去做。
GEN|7|6|当洪水 在地上泛滥的时候， 挪亚 已六百岁。
GEN|7|7|挪亚 同他的儿子、妻子和媳妇都进入方舟，躲避洪水。
GEN|7|8|洁净的牲畜和不洁净的牲畜，飞鸟及所有爬行在土地上的，
GEN|7|9|都一对一对，有公有母，到 挪亚 那里，进入方舟，正如上帝所吩咐 挪亚 的。
GEN|7|10|过了七天，洪水泛滥在地上。
GEN|7|11|挪亚 六百岁那一年的二月十七日，就在那一天，大深渊的泉源都裂开，天上的窗户也敞开了，
GEN|7|12|四十昼夜有大雨降在地上。
GEN|7|13|正在那日， 挪亚 和他的儿子 闪 、 含 、 雅弗 ，以及 挪亚 的妻子和三个媳妇，都一同进入方舟。
GEN|7|14|他们和一切走兽，各从其类；一切牲畜，各从其类；地上爬的一切爬行动物，各从其类；一切的鸟，就是一切有翅膀的飞禽，各从其类；
GEN|7|15|凡有生命气息的血肉之躯，都一对一对到 挪亚 那里，进入方舟。
GEN|7|16|凡有血肉的，都一公一母进入方舟，正如上帝所吩咐 挪亚 的。耶和华就把他关在方舟里。
GEN|7|17|洪水在地上泛滥四十天，水往上涨，使方舟浮起，方舟就从地上漂起来。
GEN|7|18|水势汹涌，在地上大大上涨，方舟在水面上漂荡。
GEN|7|19|水势在地上极其浩大，普天下所有的高山都淹没了。
GEN|7|20|水势汹涌，比山高出十五肘 ，山岭都淹没了。
GEN|7|21|凡有血肉在地上行动的，就是飞鸟、牲畜、走兽和地上成群的群聚动物，以及所有的人，都死了。
GEN|7|22|在干地上凡鼻孔里有生命气息的都死了。
GEN|7|23|耶和华除灭了地面上各类的生物，包括人和牲畜、爬行动物，以及天空的飞鸟；他们就都从地上除灭了，只剩下 挪亚 和那些与他同在方舟里的。
GEN|7|24|水势汹涌，在地上共一百五十天。
GEN|8|1|上帝记念 挪亚 和 挪亚 方舟里的一切走兽牲畜。上帝使风吹地，水势渐落。
GEN|8|2|深渊的泉源和天上的窗户都关闭了，雨不再从天降下。
GEN|8|3|水从地上逐渐消退。过了一百五十天，水就退了。
GEN|8|4|七月十七日，方舟停在 亚拉腊山 上。
GEN|8|5|水继续退去，直到十月；十月初一，山顶都露出来了。
GEN|8|6|过了四十天， 挪亚 打开他所造的方舟的窗户，
GEN|8|7|放出一只乌鸦。那乌鸦飞来飞去，直到地上的水都干了。
GEN|8|8|他又从他那里放出一只鸽子，要看水从地面上退了没有。
GEN|8|9|但全地面都是水，鸽子找不到落脚之地，就回到方舟 挪亚 那里。 挪亚 伸手接了鸽子，把它带进方舟。
GEN|8|10|挪亚 又另外等了七天，再把鸽子从方舟放出去。
GEN|8|11|到了晚上，鸽子回到他那里，看哪，嘴里有一片刚啄下来的橄榄叶， 挪亚 就知道水已经从地上退了。
GEN|8|12|他又另外等了七天，再放出鸽子，这次鸽子不再回到他那里了。
GEN|8|13|当 挪亚 六百零一岁，正月初一的时候，地上的水都干了。 挪亚 打开方舟的盖观看，看哪，地面干了。
GEN|8|14|到了二月二十七日，地就都干了。
GEN|8|15|上帝对 挪亚 说：
GEN|8|16|“你同你的妻子、儿子、媳妇都要出方舟。
GEN|8|17|凡与你一起有血肉的生物，就是飞鸟、牲畜和地上爬的一切爬行动物，都要带出来。 它们要在地上滋生，繁殖增多。”
GEN|8|18|于是 挪亚 同他的儿子、妻子、媳妇都出来了。
GEN|8|19|一切走兽、爬行动物和飞鸟，地上所有的动物，各从其类，也都出了方舟。
GEN|8|20|挪亚 为耶和华筑了一座坛，拿各种洁净的牲畜和各种洁净的飞鸟，献在坛上为燔祭。
GEN|8|21|耶和华闻了那馨香之气，耶和华心里说：“我不再因人的缘故诅咒土地，因为人从幼年就心里怀着恶念；我也不再照我曾做的毁灭一切生物了。
GEN|8|22|地还存在的时候，撒种、收割、寒暑、冬夏、昼夜都永不止息。”
GEN|9|1|上帝赐福给 挪亚 和他的儿子，对他们说：“你们要生养众多，遍满这地。
GEN|9|2|地上一切的走兽、天空一切的飞鸟、所有爬行在土地上的和海里一切的鱼都必怕你们，畏惧你们，它们都要交在你们手里。
GEN|9|3|凡活的动物都可作你们的食物。这一切我都赐给你们，如同绿色的菜蔬一样。
GEN|9|4|只是带着生命的肉，就是带着血的，你们不可吃。
GEN|9|5|流你们血、害你们命的，我必向他追讨；我要向一切走兽追讨，向人和向人的弟兄追讨人命。
GEN|9|6|凡流人血的，他的血也必被人所流，因为上帝造人，是照自己的形像造的。
GEN|9|7|你们要生养众多，在地上繁衍昌盛。”
GEN|9|8|上帝对 挪亚 和同他一起的儿子说：
GEN|9|9|“看哪，我要与你们和你们后裔立我的约，
GEN|9|10|包括和你们一起所有的生物，就是飞鸟、牲畜、地上一切的走兽，凡从方舟里出来地上一切的生物。
GEN|9|11|我与你们立我的约：凡有血肉的，不再被洪水灭绝，也不再有洪水毁坏这地了。”
GEN|9|12|上帝说：“这是我与你们，以及和你们一起的一切生物所立之约的记号，直到万代：
GEN|9|13|我把彩虹放在云中，这就是我与地立约的记号了。
GEN|9|14|我使云遮地的时候，会有彩虹出现在云中，
GEN|9|15|我就记念我与你们，以及各样有血肉的生物所立的约：不再有洪水泛滥去毁灭一切有血肉的了。
GEN|9|16|彩虹出现在云中，我看见了，就要记念上帝与地上一切有血肉的生物所立的永约。”
GEN|9|17|上帝对 挪亚 说：“这就是我与地上一切有血肉的立约的记号。”
GEN|9|18|挪亚 的儿子，从方舟出来的，有 闪 、 含 和 雅弗 。 含 是 迦南 的父亲。
GEN|9|19|这是 挪亚 的三个儿子，他们的后裔散布全地。
GEN|9|20|挪亚 是农夫，是他开始栽葡萄园的。
GEN|9|21|他喝了一些酒就醉了，在他的帐棚里赤着身子。
GEN|9|22|迦南 的父亲 含 看见他父亲赤身，就到外面告诉他的两个兄弟。
GEN|9|23|于是 闪 和 雅弗 拿了外衣搭在二人肩上，倒退着进去，遮盖父亲的赤身；他们背着脸，看不见父亲的赤身。
GEN|9|24|挪亚 酒醒以后，知道小儿子向他所做的事，
GEN|9|25|就说： “ 迦南 当受诅咒， 必给他弟兄作奴仆的奴仆。”
GEN|9|26|又说： “耶和华— 闪 的上帝是应当称颂的！ 愿 迦南 作 闪 的奴仆。
GEN|9|27|愿上帝使 雅弗 扩张， 愿他住在 闪 的帐棚里； 愿 迦南 作他的奴仆。”
GEN|9|28|洪水以后， 挪亚 又活了三百五十年。
GEN|9|29|挪亚 共活了九百五十年，就死了。
GEN|10|1|这是 挪亚 的儿子 闪 、 含 、 雅弗 的后代。洪水以后，他们都生了儿子。
GEN|10|2|雅弗 的儿子是 歌篾 、 玛各 、 玛代 、 雅完 、 土巴 、 米设 、 提拉 。
GEN|10|3|歌篾 的儿子是 亚实基拿 、 利法 、 陀迦玛 。
GEN|10|4|雅完 的儿子是 以利沙 、 他施 、 基提 、 罗单 人 。
GEN|10|5|从这些人中有沿海国家的人散居各处，有自己的土地，各有各的语言、宗族、国家。
GEN|10|6|含 的儿子是 古实 、 麦西 、 弗 、 迦南 。
GEN|10|7|古实 的儿子是 西巴 、 哈腓拉 、 撒弗他 、 拉玛 、 撒弗提迦 。 拉玛 的儿子是 示巴 、 底但 。
GEN|10|8|古实 又生 宁录 ，他是地上第一个勇士。
GEN|10|9|他在耶和华面前是个英勇的猎人，所以有话说：“像 宁录 在耶和华面前是个英勇的猎人。”
GEN|10|10|他王国的开始是在 巴别 、 以力 、 亚甲 、 甲尼 ，都在 示拿 地。
GEN|10|11|他从那地出来往 亚述 去，建造了 尼尼微 、 利河伯 、 迦拉 ，
GEN|10|12|以及 尼尼微 和 迦拉 之间的 利鲜 ，那是座大城。
GEN|10|13|麦西 生 路低 人、 亚拿米 人、 利哈比 人、 拿弗土希 人、
GEN|10|14|帕斯鲁细 人、 迦斯路希 人、 迦斐托 人； 非利士 人是从 迦斐托 人 出来的。
GEN|10|15|迦南 生了长子 西顿 ，又生 赫
GEN|10|16|和 耶布斯 人、 亚摩利 人、 革迦撒 人、
GEN|10|17|希未 人、 亚基 人、 西尼 人、
GEN|10|18|亚瓦底 人、 洗玛利 人、 哈马 人，后来 迦南 的家族散开了。
GEN|10|19|迦南 的疆界是从 西顿 到 基拉耳 ，直到 迦萨 ，又到 所多玛 、 蛾摩拉 、 押玛 、 洗扁 ，直到 拉沙 。
GEN|10|20|这就是 含 的后裔，各有自己的宗族、语言、土地和国家。
GEN|10|21|闪 也生了儿子，他是 雅弗 的哥哥 ，是 希伯 人的祖先。
GEN|10|22|闪 的儿子是 以拦 、 亚述 、 亚法撒 、 路德 、 亚兰 。
GEN|10|23|亚兰 的儿子是 乌斯 、 户勒 、 基帖 、 玛施 。
GEN|10|24|亚法撒 生 沙拉 ， 沙拉 生 希伯 。
GEN|10|25|希伯 生了两个儿子，一个名叫 法勒 ，因为那时人分地居住； 法勒 的兄弟名叫 约坍 。
GEN|10|26|约坍 生 亚摩答 、 沙列 、 哈萨玛非 、 耶拉 、
GEN|10|27|哈多兰 、 乌萨 、 德拉 、
GEN|10|28|俄巴路 、 亚比玛利 、 示巴 、
GEN|10|29|阿斐 、 哈腓拉 、 约巴 ，这些都是 约坍 的儿子。
GEN|10|30|他们所住的地方是从 米沙 直到 西发 ，到东边的山。
GEN|10|31|这就是 闪 的后裔，各有自己的宗族、语言、土地和国家。
GEN|10|32|这些是 挪亚 儿子的宗族，按着他们的后代立国。洪水以后，邦国就从他们散布在地上。
GEN|11|1|那时，全地只有一种语言，都说一样的话。
GEN|11|2|他们向东迁移的时候，在 示拿 地找到一片平原，就住在那里。
GEN|11|3|他们彼此商量说：“来，让我们来做砖，把砖烧透了。”他们就拿砖当石头，又拿柏油当泥浆。
GEN|11|4|他们说：“来，让我们建造一座城和一座塔，塔顶通天。我们要为自己立名，免得我们分散在全地面上。”
GEN|11|5|耶和华降临，要看世人所建造的城和塔。
GEN|11|6|耶和华说：“看哪，他们成了同一个民族，都有一样的语言。这只是他们开始做的事，现在他们想要做的任何事，就没有什么可拦阻他们了。
GEN|11|7|来，我们下去，在那里变乱他们的语言，使他们彼此语言不通。”
GEN|11|8|于是耶和华使他们从那里分散在全地面上；他们就停止建造那城了。
GEN|11|9|因为耶和华在那里变乱了全地的语言，把人从那里分散在全地面上，所以那城名叫 巴别 。
GEN|11|10|这是 闪 的后代。洪水以后二年， 闪 一百岁生了 亚法撒 。
GEN|11|11|闪 生 亚法撒 之后又活了五百年，并且生儿育女。
GEN|11|12|亚法撒 活到三十五岁，生了 沙拉 。
GEN|11|13|亚法撒 生 沙拉 之后又活了四百零三年，并且生儿育女。
GEN|11|14|沙拉 活到三十岁，生了 希伯 。
GEN|11|15|沙拉 生 希伯 之后又活了四百零三年，并且生儿育女。
GEN|11|16|希伯 活到三十四岁，生了 法勒 。
GEN|11|17|希伯 生 法勒 之后又活了四百三十年，并且生儿育女。
GEN|11|18|法勒 活到三十岁，生了 拉吴 。
GEN|11|19|法勒 生 拉吴 之后又活了二百零九年，并且生儿育女。
GEN|11|20|拉吴 活到三十二岁，生了 西鹿 。
GEN|11|21|拉吴 生 西鹿 之后又活了二百零七年，并且生儿育女。
GEN|11|22|西鹿 活到三十岁，生了 拿鹤 。
GEN|11|23|西鹿 生 拿鹤 之后又活了二百年，并且生儿育女。
GEN|11|24|拿鹤 活到二十九岁，生了 他拉 。
GEN|11|25|拿鹤 生 他拉 之后又活了一百一十九年，并且生儿育女。
GEN|11|26|他拉 活到七十岁，生了 亚伯兰 、 拿鹤 和 哈兰 。
GEN|11|27|这是 他拉 的后代。 他拉 生 亚伯兰 、 拿鹤 和 哈兰 ； 哈兰 生 罗得 。
GEN|11|28|哈兰 死在他父亲 他拉 的面前，死在他的出生地 迦勒底 的 吾珥 。
GEN|11|29|亚伯兰 、 拿鹤 各娶了妻。 亚伯兰 的妻子名叫 撒莱 ， 拿鹤 的妻子名叫 密迦 ，是 哈兰 的女儿。 哈兰 是 密迦 和 亦迦 的父亲。
GEN|11|30|撒莱 不生育，没有孩子。
GEN|11|31|他拉 带着他儿子 亚伯兰 和他孙子， 哈兰 的儿子 罗得 ，以及他的媳妇， 亚伯兰 的妻子 撒莱 ，一同出了 迦勒底 的 吾珥 ，要往 迦南 地去；他们来到 哈兰 ，就住在那里。
GEN|11|32|他拉 共活了二百零五年，就死在 哈兰 。
GEN|12|1|耶和华对 亚伯兰 说：“你要离开本地、本族、父家，往我所要指示你的地去。
GEN|12|2|我必使你成为大国，我必赐福给你，使你的名为大；你要使别人得福 。
GEN|12|3|为你祝福的，我必赐福给他；诅咒你的，我必诅咒他。地上的万族都必因你得福。”
GEN|12|4|亚伯兰 就遵照耶和华的吩咐去了； 罗得 也和他同去。 亚伯兰 离开 哈兰 的时候年七十五岁。
GEN|12|5|亚伯兰 带着他妻子 撒莱 和侄儿 罗得 ，以及他们在 哈兰 积蓄的财物、获得的人口，往 迦南 地去。他们就来到了 迦南 地。
GEN|12|6|亚伯兰 经过那地，直到 示剑 地方， 摩利 橡树那里；当时 迦南 人住在那地。
GEN|12|7|耶和华向 亚伯兰 显现，说：“我要把这地赐给你的后裔。” 亚伯兰 就在那里为向他显现的耶和华筑了一座坛。
GEN|12|8|从那里他又迁到 伯特利 东边的山，支搭帐棚；西边是 伯特利 ，东边是 艾 。他在那里又为耶和华筑了一座坛，求告耶和华的名。
GEN|12|9|后来 亚伯兰 渐渐迁往 尼革夫 去。
GEN|12|10|那地遭遇饥荒。 亚伯兰 因那地的饥荒严重，就下到 埃及 ，要在那里寄居。
GEN|12|11|将近 埃及 ，他对妻子 撒莱 说：“看哪，我知道你是美貌的女人。
GEN|12|12|埃及 人看见你会说：‘这是他的妻子’，他们就会杀我，却让你活着。
GEN|12|13|所以，请你说你是我的妹妹，使我可以因你得平安，我的性命也因你存活。”
GEN|12|14|亚伯兰 到达 埃及 时， 埃及 人看见那女人极其美貌。
GEN|12|15|法老的臣仆看见了她，就在法老面前称赞她。那女人就被带进法老的宫中。
GEN|12|16|法老就因她厚待 亚伯兰 ，给了 亚伯兰 许多牛、羊、公驴、奴仆、婢女、母驴、骆驼。
GEN|12|17|耶和华因 亚伯兰 妻子 撒莱 的缘故，降大灾击打法老和他的全家。
GEN|12|18|法老召了 亚伯兰 来，说：“你向我做的是什么事呢？为什么没有告诉我她是你的妻子？
GEN|12|19|为什么说‘她是我的妹妹’，以致我把她接来要作我的妻子呢？现在 ，看哪，你的妻子在这里，带她走吧！”
GEN|12|20|于是法老吩咐人把 亚伯兰 和他妻子，以及他一切所有的都送走了。
GEN|13|1|亚伯兰 带着他的妻子与 罗得 ，以及一切所有的，从 埃及 上 尼革夫 去。
GEN|13|2|亚伯兰 的牲畜和金银极多。
GEN|13|3|他从 尼革夫 渐渐往 伯特利 去，到了 伯特利 和 艾 的中间，当初他支搭帐棚的地方，
GEN|13|4|也是他起先筑坛的地方。 亚伯兰 在那里求告耶和华的名。
GEN|13|5|与 亚伯兰 同行的 罗得 也有牛群、羊群、帐棚。
GEN|13|6|那地容不下他们住在一起；因为他们的财物非常多，使他们不能同住一起。
GEN|13|7|当时， 迦南 人与 比利洗 人在那地居住。 亚伯兰 的牧人和 罗得 的牧人之间起了争端。
GEN|13|8|亚伯兰 就对 罗得 说：“你我不可以相争，你的牧人和我的牧人也不可以相争，因为我们是一家人。
GEN|13|9|遍地不都在你眼前吗？请你离开我吧！你向左，我就向右；你向右，我就向左。”
GEN|13|10|罗得 举目，看见 约旦河 整个平原，直到 琐珥 ，都是水源充足之地。在耶和华未毁灭 所多玛 、 蛾摩拉 以前，那地好像耶和华的园子，又像 埃及 地。
GEN|13|11|于是 罗得 选择了 约旦河 整个平原。 罗得 往东迁移，他们就彼此分开了。
GEN|13|12|亚伯兰 住在 迦南 地； 罗得 住在平原的城镇，他渐渐迁移帐棚，直到 所多玛 。
GEN|13|13|所多玛 人在耶和华面前罪大恶极。
GEN|13|14|罗得 离开 亚伯兰 以后，耶和华对 亚伯兰 说：“你要从你所在的地方，举目向东西南北观看；
GEN|13|15|你所看见一切的地，我都要把它赐给你和你的后裔，直到永远。
GEN|13|16|我要使你的后裔好像地上的尘沙，人若能数地上的尘沙，才能数你的后裔。
GEN|13|17|你起来，纵横走遍这地，因为我必把这地赐给你。”
GEN|13|18|亚伯兰 就迁移帐棚，来到 希伯仑 ， 幔利 的橡树那里居住，在那里为耶和华筑了一座坛。
GEN|14|1|当 暗拉非 作 示拿 王， 亚略 作 以拉撒 王， 基大老玛 作 以拦 王， 提达 作 戈印 王的时候，
GEN|14|2|他们攻打 所多玛 王 比拉 、 蛾摩拉 王 比沙 、 押玛 王 示纳 、 洗扁 王 善以别 和 比拉 王， 比拉 就是 琐珥 。
GEN|14|3|这些王都会合在 西订谷 ， 西订谷 就是 盐海 。
GEN|14|4|他们已经服事 基大老玛 十二年，第十三年就背叛了。
GEN|14|5|第十四年， 基大老玛 和与他结盟的王都来了，在 亚特律．加宁 击败 利乏音 人，在 哈麦 击败 苏西 人，在 沙微．基列亭 击败 以米 人，
GEN|14|6|在 何利 人的 西珥山 击败 何利 人，一直到靠近旷野的 伊勒．巴兰 。
GEN|14|7|他们转回，来到 安．密巴 ，就是 加低斯 ，击败了 亚玛力 全地的人，以及住在 哈洗逊．他玛 的 亚摩利 人。
GEN|14|8|于是 所多玛 王、 蛾摩拉 王、 押玛 王、 洗扁 王和 比拉 王， 比拉 就是 琐珥 ，都出来，在 西订谷 摆阵，与他们交战，
GEN|14|9|就是与 以拦 王 基大老玛 、 戈印 王 提达 、 示拿 王 暗拉非 、 以拉撒 王 亚略 交战；这就是四王对五王之战。
GEN|14|10|西订谷 有许多柏油坑。 所多玛 王和 蛾摩拉 王逃跑，掉在坑里，其余的人都往山上逃跑。
GEN|14|11|四王就把 所多玛 和 蛾摩拉 所有的财物和所有的粮食都掳掠去了；
GEN|14|12|他们也把 亚伯兰 的侄儿 罗得 和 罗得 的财物都掳掠去了。当时 罗得 住在 所多玛 。
GEN|14|13|有一个逃脱的人来告诉 希伯来 人 亚伯兰 ； 亚伯兰 正住在 亚摩利 人 幔利 的橡树那里。 幔利 、 以实各 和 亚乃 都是弟兄，曾与 亚伯兰 结盟。
GEN|14|14|亚伯兰 听见他侄儿 被掳去，就把三百一十八个生在他家中、受过训练的壮丁全都出动 去追，一直到 但 。
GEN|14|15|在夜间，他和他的仆人分队击败了敌人，并且追杀他们，直到 大马士革 北边的 何把 。
GEN|14|16|他把一切被掳掠的财物夺回，也把他侄儿 罗得 和他的财物，以及人和妇女都夺回来。
GEN|14|17|亚伯兰 击败 基大老玛 和与他结盟的王回来的时候， 所多玛 王出来，在 沙微谷 迎接他， 沙微谷 就是 王的谷 。
GEN|14|18|又有 撒冷 王 麦基洗德 带着饼和酒出来；他是至高上帝的祭司。
GEN|14|19|他为 亚伯兰 祝福，说： “愿至高的上帝、 天地的主赐福给 亚伯兰 ！
GEN|14|20|至高的上帝把敌人交在你手里， 他是应当称颂的！” 亚伯兰 就把所有的拿出十分之一给他。
GEN|14|21|所多玛 王对 亚伯兰 说：“你把人还给我，财物你自己拿去吧！”
GEN|14|22|亚伯兰 对 所多玛 王说：“我指着耶和华—至高的上帝、天地的主起誓：
GEN|14|23|凡是你的东西，就是一根线、一条鞋带，我都不拿，免得你说：‘是我使 亚伯兰 富足！’
GEN|14|24|我什么都不要，只是仆人所吃的，以及与我同去的 亚乃 、 以实各 、 幔利 所应得的份，让他们拿去吧！”
GEN|15|1|这些事以后，耶和华的话在异象中临到 亚伯兰 ，说：“ 亚伯兰 哪，不要惧怕！我是你的盾牌，你必得丰富的赏赐。”
GEN|15|2|亚伯兰 说：“主耶和华啊，我还没有儿子，你能赐我什么呢？承受我家业的是 大马士革 人 以利以谢 。”
GEN|15|3|亚伯兰 又说：“看哪，你没有给我后嗣。你看，那生在我家中的人要继承我。”
GEN|15|4|看哪，耶和华的话又临到他，说：“这人不会继承你，你本身所生的才会继承你。”
GEN|15|5|于是耶和华带他到外面，说：“你向天观看，去数星星，你能数得清吗？”又对他说：“你的后裔将要如此。”
GEN|15|6|亚伯兰 信耶和华，耶和华就以此算他为义。
GEN|15|7|耶和华又对他说：“我是耶和华，曾领你出 迦勒底 的 吾珥 ，为要把这地赐你为业。”
GEN|15|8|亚伯兰 说：“主耶和华啊，我怎能知道我必得这地为业呢？”
GEN|15|9|耶和华对他说：“你为我取一头三岁的母牛犊，一只三岁的母山羊，一只三岁的公绵羊，一只斑鸠和一只雏鸽。”
GEN|15|10|亚伯兰 就把这些都取来，每样从中间劈成两半，一半对着另一半排列，只有鸟没有劈开。
GEN|15|11|当鸷鸟下来，落在这些尸体上时， 亚伯兰 就把它们赶走了。
GEN|15|12|日落的时候， 亚伯兰 沉睡了。看哪，有大而可怕的黑暗落在他身上。
GEN|15|13|耶和华对 亚伯兰 说：“你要确实知道，你的后裔必寄居在别人的地，服事那地的人；那地的人要虐待他们四百年。
GEN|15|14|但我要惩罚他们所服事的那国，以后他们必带着许多财物从那里出来。
GEN|15|15|至于你，你要平平安安归到你祖先那里，必享长寿，被人埋葬。
GEN|15|16|到了第四代，他们必回到这里，因为 亚摩利 人的罪恶到现在还没有满盈。”
GEN|15|17|日落天黑的时候，看哪，有冒烟的炉和烧着的火把从那些肉块中经过。
GEN|15|18|在那日，耶和华与 亚伯兰 立约，说：“我已赐给你的后裔这一片地，从 埃及河 直到 大河 ， 幼发拉底河 ，
GEN|15|19|就是 基尼 人、 基尼洗 人、 甲摩尼 人、
GEN|15|20|赫 人、 比利洗 人、 利乏音 人、
GEN|15|21|亚摩利 人、 迦南 人、 革迦撒 人、 耶布斯 人的地。”
GEN|16|1|亚伯兰 的妻子 撒莱 没有为他生孩子。 撒莱 有一个婢女，是 埃及 人，名叫 夏甲 。
GEN|16|2|撒莱 对 亚伯兰 说：“看哪，耶和华使我不能生育。你来和我的婢女同房，也许我可以从她得孩子 。” 亚伯兰 听从了 撒莱 的话。
GEN|16|3|于是 亚伯兰 的妻子 撒莱 把她的婢女， 埃及 人 夏甲 ，给了丈夫为妾；那时 亚伯兰 在 迦南 已经住了十年。
GEN|16|4|亚伯兰 与 夏甲 同房， 夏甲 就怀了孕。她看见自己有孕，就轻视她的女主人。
GEN|16|5|撒莱 对 亚伯兰 说：“我因你受了委屈。我把我的婢女放在你怀中，她见自己怀了孕，就轻视我。愿耶和华在你我之间判断。”
GEN|16|6|亚伯兰 对 撒莱 说：“看哪，婢女在你手里，你可以照你看为好的对待她。”于是， 撒莱 虐待她，她就从 撒莱 面前逃走了。
GEN|16|7|耶和华的使者在旷野的水泉旁，在 书珥 路上的水泉旁遇见 夏甲 ，
GEN|16|8|对她说：“ 撒莱 的婢女 夏甲 ，你从哪里来？要到哪里去？”她说：“我从我的女主人 撒莱 面前逃出来。”
GEN|16|9|耶和华的使者对她说：“你要回到你的女主人那里，屈服在她手下。”
GEN|16|10|耶和华的使者对她说： “我必使你的后裔极其繁多， 多到不可胜数。”
GEN|16|11|耶和华的使者又对她说： “看哪，你已怀孕， 要生一个儿子。 你要给他起名叫 以实玛利 ， 因为耶和华听见了你的苦楚。
GEN|16|12|他为人必像野驴。 他的手要攻打人， 人的手也要攻打他； 他必常与他的众弟兄作对 。”
GEN|16|13|夏甲 就称那向她说话的耶和华为“你是看见 的上帝”，因为她说：“他看见了我之后，我还能在这里看见他吗？”
GEN|16|14|所以这井名叫 庇耳．拉海．莱 ，看哪，它位于 加低斯 和 巴列 的中间。
GEN|16|15|后来 夏甲 为 亚伯兰 生了一个儿子； 亚伯兰 给 夏甲 生的儿子起名叫 以实玛利 。
GEN|16|16|夏甲 为 亚伯兰 生 以实玛利 的时候， 亚伯兰 年八十六岁。
GEN|17|1|亚伯兰 九十九岁时，耶和华向他显现，对他说：“我是全能的上帝。你当在我面前行走，作完全的人，
GEN|17|2|我要与你立约，使你的后裔极其繁多。”
GEN|17|3|亚伯兰 脸伏于地；上帝又对他说：
GEN|17|4|“看哪，这就是我与你立的约，你要成为多国的父。
GEN|17|5|从今以后，你的名字不再叫 亚伯兰 ，要叫 亚伯拉罕 ，因为我已经立你作多国之父。
GEN|17|6|我必使你生养极其繁多；国度要从你而立，君王要从你而出。
GEN|17|7|我要与你，以及你世世代代的后裔坚立我的约，成为永远的约，是要作你和你后裔的上帝。
GEN|17|8|我要把你现在寄居的地，就是 迦南 全地，赐给你和你的后裔永远为业；我也必作他们的上帝。”
GEN|17|9|上帝又对 亚伯拉罕 说：“你和你的后裔一定要世世代代遵守我的约。
GEN|17|10|这就是我与你，以及你的后裔所立的约，是你们所当遵守的，你们所有的男子都要受割礼。
GEN|17|11|你们要割去肉体的包皮，这是我与你们立约的记号。
GEN|17|12|你们世世代代的男子，无论是在家里生的，或是用银子从外人买来而不是你后裔生的，都要在生下来的第八日受割礼。
GEN|17|13|你家里生的和你用银子买的，都必须受割礼。这样，我的约就在你们肉体上成为永远的约。
GEN|17|14|不受割礼的男子都必从民中剪除，因他违背了我的约。”
GEN|17|15|上帝又对 亚伯拉罕 说：“至于你的妻子 撒莱 ，不可再叫她 撒莱 ，她的名要叫 撒拉 。
GEN|17|16|我必赐福给她，也要从她赐一个儿子给你。我必赐福给 撒拉 ，她要兴起多国；必有百姓的君王从她而出。”
GEN|17|17|亚伯拉罕 就脸伏于地窃笑，心里想：“一百岁的人还能有孩子吗？ 撒拉 已经九十岁了，还能生育吗？”
GEN|17|18|亚伯拉罕 对上帝说：“但愿 以实玛利 活在你面前。”
GEN|17|19|上帝说：“不！你妻子 撒拉 必为你生一个儿子，你要给他起名叫 以撒 。我要与他坚立我的约，成为他后裔永远的约。
GEN|17|20|至于 以实玛利 ，我已听见你了：看哪，我必赐福给他，使他兴旺，极其繁多。他必生十二个族长，我要使他成为大国。
GEN|17|21|到明年所定的时候， 撒拉 必为你生 以撒 ，我要与他坚立我的约。”
GEN|17|22|上帝和 亚伯拉罕 说完了话，就离开他上升去了。
GEN|17|23|在那一天， 亚伯拉罕 遵照上帝所说的，给他的儿子 以实玛利 和家里所有的男丁，无论是在家里生的，或是用银子买来的，都行了割礼 。
GEN|17|24|亚伯拉罕 受割礼时，年九十九岁。
GEN|17|25|他儿子 以实玛利 受割礼时，年十三岁。
GEN|17|26|在那一天， 亚伯拉罕 和他儿子 以实玛利 一同受了割礼。
GEN|17|27|家里所有的男人，无论是在家里生的，或是用银子从外人买来的，也都一同受了割礼。
GEN|18|1|耶和华在 幔利 橡树那里向 亚伯拉罕 显现。天正热的时候， 亚伯拉罕 坐在帐棚门口。
GEN|18|2|他举目观看，看哪，有三个人站在他附近。他一看见，就从帐棚门口跑去迎接他们，俯伏在地，
GEN|18|3|说：“我主，我若在你眼前蒙恩，请不要离开你的仆人走过去。
GEN|18|4|容我拿点水来，请你们洗脚，在树下休息。
GEN|18|5|既然你们来到仆人这里了，我再拿点饼来，让你们恢复心力，然后再走。”他们说：“就照你说的去做吧。”
GEN|18|6|亚伯拉罕 急忙进帐棚到 撒拉 那里，说：“你赶快拿三细亚细面，揉面做饼。”
GEN|18|7|亚伯拉罕 又跑到牛群里，牵了一头又嫩又好的牛犊来，交给仆人，仆人就急忙去预备。
GEN|18|8|亚伯拉罕 取了乳酪和奶，以及预备好了的牛犊来，摆在他们面前，自己在树下站在旁边，他们就吃了。
GEN|18|9|他们对 亚伯拉罕 说：“你妻子 撒拉 在哪里？”他说：“看哪，在帐棚里。”
GEN|18|10|有一位说：“明年这时候 ，我一定会回到你这里。看哪，你的妻子 撒拉 会生一个儿子。” 撒拉 在那人后面的帐棚门口也听见了。
GEN|18|11|亚伯拉罕 和 撒拉 都年纪老迈， 撒拉 的月经已停了。
GEN|18|12|撒拉 心里窃笑，说：“我已衰老，我的主也老了，怎能有这喜事呢？”
GEN|18|13|耶和华对 亚伯拉罕 说：“ 撒拉 为什么窃笑，说：‘我已年老，果真能生育吗？’
GEN|18|14|耶和华岂有难成的事吗？到了所定的时候，我必回到你这里。明年这时候， 撒拉 会生一个儿子。”
GEN|18|15|撒拉 因为害怕，就不承认，说：“我没有笑。”那人说：“不，你的确笑了。”
GEN|18|16|三人从那里起程，面向 所多玛 观望， 亚伯拉罕 与他们同行，要送他们一程。
GEN|18|17|耶和华说：“我所要做的事岂可瞒着 亚伯拉罕 呢？
GEN|18|18|亚伯拉罕 必要成为强大的国；地上的万国都必因他得福。
GEN|18|19|我拣选他 ，为要叫他命令他的子孙和后代家属遵行耶和华的道，秉公行义，使耶和华所应许 亚伯拉罕 的话都实现了。”
GEN|18|20|耶和华说：“ 所多玛 和 蛾摩拉 罪恶极其严重，控告他们的声音很大。
GEN|18|21|我要下去察看他们所做的，是否真的像那达到我这里的声音一样；如果不是，我也要知道。”
GEN|18|22|二人转身离开那里，往 所多玛 去；但 亚伯拉罕 仍然站在耶和华面前。
GEN|18|23|亚伯拉罕 近前来，说：“你真的要把义人和恶人一同剿灭吗？
GEN|18|24|假若那城里有五十个义人，你真的还要剿灭，不因城里这五十个义人饶了那地方吗？
GEN|18|25|你绝不会做这样的事，把义人与恶人一同杀了，使义人与恶人一样。你绝不会这样！审判全地的主岂不做公平的事吗？”
GEN|18|26|耶和华说：“我若在 所多玛城 里找到五十个义人，我就为他们的缘故饶恕那整个地方。”
GEN|18|27|亚伯拉罕 回答说：“看哪，我虽只是尘土灰烬，还敢向主说话。
GEN|18|28|假若这五十个义人少了五个，你就因为少了五个而毁灭全城吗？”他说：“我在那里若找到四十五个，就不毁灭。”
GEN|18|29|亚伯拉罕 又对他说：“假若在那里找到四十个呢？”他说：“为这四十个的缘故，我也不做。”
GEN|18|30|亚伯拉罕 说：“求主不要生气，容我说，假若在那里找到三十个呢？”他说：“我在那里若找到三十个，我也不做。”
GEN|18|31|亚伯拉罕 说：“看哪，我还敢向主说，假若在那里找到二十个呢？”他说：“为这二十个的缘故，我也不毁灭。”
GEN|18|32|亚伯拉罕 说：“求主不要生气，我再说一次，假若在那里找到十个呢？”他说：“为这十个的缘故，我也不毁灭。”
GEN|18|33|耶和华与 亚伯拉罕 说完了话就走了； 亚伯拉罕 也回到自己的地方去了。
GEN|19|1|两个天使在傍晚到了 所多玛 ， 罗得 正坐在 所多玛 的城门口。 罗得 一看见，就起身迎接他们，脸伏于地下拜，
GEN|19|2|说：“看哪，我主，请你们转到仆人家里过夜，洗你们的脚，清早起来再上路。”他们说：“不！我们要在广场上过夜。”
GEN|19|3|罗得 恳切地请他们，他们就转向他，进到他屋里。 罗得 为他们预备宴席，烤无酵饼，他们就吃了。
GEN|19|4|他们还没有躺下， 所多玛城 的人，连老带少所有的人，个个都来围住那屋子。
GEN|19|5|他们呼叫 罗得 ，对他说：“今天晚上到你这里来的人在哪里？把他们带出来，让我们亲近他们。”
GEN|19|6|罗得 出了门，把身后的门关上，到众人那里，
GEN|19|7|说：“我的弟兄们，请你们不要做这恶事。
GEN|19|8|看哪，我有两个女儿，还没有亲近过男人，让我领她们出来给你们，就照你们看为好的对待她们吧！只是这两个人既然到我舍下，请不要向他们做这事。”
GEN|19|9|众人说：“站到一边去吧！”又说：“这个人来寄居，还想扮审判官呢！现在我们要害你比害他们更厉害。”众人就往前冲向 罗得 ，要攻破大门。
GEN|19|10|那两个人伸出手来，把 罗得 拉进屋子他们那里，就关上门。
GEN|19|11|他们击打门外的人，无论老少，都眼睛迷糊，找门找得很烦躁。
GEN|19|12|那两个人对 罗得 说：“你这里还有什么人吗？无论是女婿，是儿女，这城中所有属你的人，你都要把他们从这地方带出去。
GEN|19|13|我们要毁灭这地方，因为控告城内百姓的声音在耶和华面前非常大，耶和华派我们来毁灭这城。”
GEN|19|14|罗得 出去，告诉娶了 他女儿的女婿们说：“起来，离开这地方，因为耶和华要毁灭这城。”他的女婿们却以为他说的是笑话。
GEN|19|15|天亮了，天使催逼 罗得 说：“起来！带着你的妻子和你这里的两个女儿出去，免得你因这城的罪孽同被剿灭。”
GEN|19|16|但 罗得 迟延不走。二人因为耶和华怜悯 罗得 ，就拉着他的手和他妻子的手，以及他两个女儿的手，把他们领出来，安置在城外；
GEN|19|17|领他们出来以后，就说：“逃命吧！不可回头看，也不可在平原站住。要往山上逃跑，免得你被剿灭。”
GEN|19|18|罗得 对他们说：“我主啊，不要这样！
GEN|19|19|看哪，你仆人已经在你眼前蒙恩，你又向我大施慈爱，救我的性命。但是我不能逃到山上去，恐怕这灾祸追上我，我就死了。
GEN|19|20|看哪，这城又近又小，比较容易逃到那里。这不是一座小城吗？求你容我逃到那里，使我的性命可以存活。”
GEN|19|21|天使对他说：“看哪，这事我也应允你，不倾覆你所说的这城。
GEN|19|22|你要赶快逃到那城，因为你还没有到那里，我不能做什么。”因此那城名叫 琐珥 。
GEN|19|23|罗得 到了 琐珥 ，太阳已经升出地面。
GEN|19|24|当时，耶和华把硫磺与火，从天上耶和华那里降与 所多玛 和 蛾摩拉 ，
GEN|19|25|把那些城和全平原，城里所有的居民和土地上生长的，都毁灭了。
GEN|19|26|罗得 的妻子在他后边回头一看，就变成了一根盐柱。
GEN|19|27|亚伯拉罕 清早起来，到了他先前站在耶和华面前的地方，
GEN|19|28|面向 所多玛 和 蛾摩拉 ，以及平原全地观望。他观看，看哪，那地有浓烟上腾，好像烧窑的浓烟。
GEN|19|29|当上帝毁灭平原诸城的时候，他记念 亚伯拉罕 ；在倾覆 罗得 所住之城的时候，就把 罗得 从倾覆中带出来。
GEN|19|30|罗得 因为怕住在 琐珥 ，就同他两个女儿从 琐珥 上去，住在山上。他和两个女儿住在一个洞里。
GEN|19|31|大女儿对小女儿说：“我们的父亲老了，这地又没有男人可以照世上的礼俗来与我们结合。
GEN|19|32|来！我们叫父亲喝酒，然后与他同寝。这样，我们可以从我们的父亲存留后裔。”
GEN|19|33|于是，那晚她们叫父亲喝酒，大女儿就进去和她父亲同寝；她几时躺下，几时起来，父亲都不知道。
GEN|19|34|第二天，大女儿对小女儿说：“看哪，我昨夜与父亲同寝。今晚我们再叫他喝酒，你进去与他同寝。这样，我们可以从父亲存留后裔。”
GEN|19|35|于是，那晚她们又叫父亲喝酒，小女儿起来与她父亲同寝；她几时躺下，几时起来，父亲都不知道。
GEN|19|36|这样， 罗得 的两个女儿都从她们的父亲怀了孕。
GEN|19|37|大女儿生了儿子，给他起名叫 摩押 ，就是现今 摩押 人的始祖。
GEN|19|38|小女儿也生了儿子，给他起名叫 便．亚米 ，就是现今 亚扪 人的始祖。
GEN|20|1|亚伯拉罕 从那里往 尼革夫 迁移，寄居在 加低斯 和 书珥 之间的 基拉耳 。
GEN|20|2|亚伯拉罕 称他的妻子 撒拉 为妹妹。 基拉耳 王 亚比米勒 派人把 撒拉 带走。
GEN|20|3|夜间，上帝在梦中来到 亚比米勒 那里，对他说：“看哪，你要死了，因为你带来的女人，她是有丈夫的女子！”
GEN|20|4|亚比米勒 还未亲近 撒拉 ；他说：“主啊，连公义的国，你也要毁灭吗？
GEN|20|5|那人岂不是自己对我说‘她是我妹妹’吗？连这女人自己也说：‘他是我哥哥。’我做这事是心正手洁的。”
GEN|20|6|上帝在梦中对他说：“我也知道你做这事是心中正直的；是我拦阻了你，免得你得罪我。所以我不让你侵犯她。
GEN|20|7|现在你当把这人的妻子归还给他；因为他是先知，他要为你祷告，使你存活。你若不归还，你当知道，你和你所有的人都必定死。”
GEN|20|8|亚比米勒 清早起来，叫了他的众臣仆来，把这一切事说给他们听，他们就很害怕。
GEN|20|9|亚比米勒 召了 亚伯拉罕 来，对他说：“你怎么向我这样做呢？我什么事得罪你，你竟使我和我的国陷在大罪中呢？你对我做了不该做的事了！”
GEN|20|10|亚比米勒 对 亚伯拉罕 说：“你看见什么才做这事呢？”
GEN|20|11|亚伯拉罕 说：“我以为这地方的人根本不敬畏上帝，必为我妻子的缘故杀我。
GEN|20|12|况且她也真是我的妹妹；她与我是同父异母的，后来作了我的妻子。
GEN|20|13|当上帝叫我离开父家、飘流在外的时候，我对她说：我们无论走到什么地方，你要对人说：‘他是我哥哥’，这就是你以慈爱待我了。”
GEN|20|14|亚比米勒 把牛、羊、奴仆、婢女送给 亚伯拉罕 ，也把他的妻子 撒拉 归还给他。
GEN|20|15|亚比米勒 说：“看哪，我的地都在你面前，你看为好的地方就居住吧。”
GEN|20|16|他对 撒拉 说：“看哪，我给你哥哥一千银子。看哪，这要在你全家人面前遮羞 ，向众人证实你是清白的。”
GEN|20|17|亚伯拉罕 向上帝祷告，上帝就医好 亚比米勒 和他的妻子，以及他的使女们，他们就能生育。
GEN|20|18|因耶和华为 亚伯拉罕 的妻子 撒拉 的缘故，已经使 亚比米勒 家中的妇人不能怀孕。
GEN|21|1|耶和华照着他所说的眷顾 撒拉 ，耶和华实现了他对 撒拉 的应许。
GEN|21|2|亚伯拉罕 年老，到上帝对他说的那所定的时候， 撒拉 怀了孕，给他生了一个儿子。
GEN|21|3|亚伯拉罕 给 撒拉 所生的儿子起名叫 以撒 。
GEN|21|4|以撒 出生后第八日， 亚伯拉罕 遵照上帝所吩咐的，为 以撒 行割礼。
GEN|21|5|他儿子 以撒 出生的时候， 亚伯拉罕 年一百岁。
GEN|21|6|撒拉 说：“上帝使我欢笑，凡听见的人必与我一同欢笑”，
GEN|21|7|又说：“谁能预先对 亚伯拉罕 说， 撒拉 要乳养孩子呢？因为在他年老的时候，我为他生了一个儿子。”
GEN|21|8|孩子渐渐长大，就断了奶。 以撒 断奶的那一天， 亚伯拉罕 摆设丰盛的宴席。
GEN|21|9|那时， 撒拉 看见 埃及 人 夏甲 为 亚伯拉罕 所生的儿子戏笑，
GEN|21|10|就对 亚伯拉罕 说：“你把这使女和她儿子赶出去！因为这使女的儿子不可与我的儿子 以撒 一同承受产业。”
GEN|21|11|亚伯拉罕 为这事非常忧愁，因为关乎他的儿子。
GEN|21|12|上帝对 亚伯拉罕 说：“你不必为这孩子和你的使女忧愁。 撒拉 对你说的话，你都要听从；因为从 以撒 生的，才要称为你的后裔。
GEN|21|13|至于使女的儿子，我也必使他成为一国，因为他是你的后裔。”
GEN|21|14|亚伯拉罕 清早起来，拿饼和一皮袋水，给了 夏甲 ，搭在她肩上，把她和孩子一起送走。 夏甲 就走了，但她却在 别是巴 的旷野流浪。
GEN|21|15|皮袋的水用完了， 夏甲 就把孩子放在一棵小树下，
GEN|21|16|自己走开约有一箭之远，相对而坐，说：“我不忍心看见孩子死”。她就坐在对面，放声大哭。
GEN|21|17|上帝听见孩子的声音，上帝的使者就从天上呼叫 夏甲 说：“ 夏甲 ，你为何这样呢？不要害怕，上帝已经听见孩子在那里的声音了。
GEN|21|18|起来！把孩子扶起来，用你的手握住他，因我必使他成为大国。”
GEN|21|19|上帝开了 夏甲 的眼睛，她就看见一口水井。她就去，把皮袋装满了水，给孩子喝。
GEN|21|20|上帝与这孩子同在，他就渐渐长大，住在旷野，成了一个弓箭手。
GEN|21|21|他住在 巴兰 的旷野；他母亲从 埃及 地为他娶了一个妻子。
GEN|21|22|那时候， 亚比米勒 和他的将军 非各 对 亚伯拉罕 说：“凡你所做的事，上帝都与你同在。
GEN|21|23|我愿你如今在这里指着上帝对我起誓，不要亏待我和我的儿子，以及我的子孙。我怎样忠诚待你，你也要照样忠诚待我和你所寄居的这地。”
GEN|21|24|亚伯拉罕 说：“我愿意起誓。”
GEN|21|25|先前， 亚比米勒 的仆人霸占了一口水井， 亚伯拉罕 为这事责备 亚比米勒 。
GEN|21|26|亚比米勒 说：“我不知道谁做了这事，你也没有告诉我，我到今日才听到。”
GEN|21|27|亚伯拉罕 把羊和牛给了 亚比米勒 ，二人就彼此立约。
GEN|21|28|亚伯拉罕 把七只小母羊另放在一处。
GEN|21|29|亚比米勒 对 亚伯拉罕 说：“你把这七只小母羊另放一处是什么意思呢？”
GEN|21|30|他说：“你要从我手里接受这七只小母羊，作我挖了这口井的证据。”
GEN|21|31|所以他给那地方起名叫 别是巴 ，因为他们二人在那里起了誓。
GEN|21|32|他们在 别是巴 立了约， 亚比米勒 就和他的将军 非各 起身回 非利士 人的地去了。
GEN|21|33|亚伯拉罕 就在 别是巴 种了一棵柳树，在那里求告耶和华—永恒上帝的名。
GEN|21|34|亚伯拉罕 在 非利士 人的地寄居了许多日子。
GEN|22|1|这些事以后，上帝考验 亚伯拉罕 ，对他说：“ 亚伯拉罕 ！”他说：“我在这里。”
GEN|22|2|上帝说：“你要带你的儿子，就是你所爱的独子 以撒 ，往 摩利亚 地去，在我指示你的一座山上，把他献为燔祭。”
GEN|22|3|亚伯拉罕 清早起来，预备了驴，带着跟他一起的两个仆人和他儿子 以撒 ，劈好了燔祭的柴，就起身往上帝指示他的地方去了。
GEN|22|4|到了第三日， 亚伯拉罕 举目遥望那地方。
GEN|22|5|亚伯拉罕 对他的仆人说：“你们和驴留在这里，我和孩子要去那里敬拜，然后回到你们这里来。”
GEN|22|6|亚伯拉罕 把燔祭的柴放在他儿子 以撒 身上，自己手里拿着火与刀；于是二人同行。
GEN|22|7|以撒 对他父亲 亚伯拉罕 说：“我父啊！” 亚伯拉罕 说：“我儿，我在这里。” 以撒 说：“看哪，火与柴都有了，但燔祭的羔羊在哪里呢？”
GEN|22|8|亚伯拉罕 说：“我儿，上帝必自己预备燔祭的羔羊。”于是二人同行。
GEN|22|9|他们到了上帝指示他的地方， 亚伯拉罕 在那里筑坛，把柴摆好，绑了他儿子 以撒 ，放在坛的柴上。
GEN|22|10|亚伯拉罕 就伸手拿刀，要杀他的儿子。
GEN|22|11|耶和华的使者从天上呼唤他说：“ 亚伯拉罕 ！ 亚伯拉罕 ！”他说：“我在这里。”
GEN|22|12|天使说：“不可在这孩子身上下手！一点也不可伤害他！现在我知道你是敬畏上帝的人了，因为你没有把你的儿子，就是你的独子，留下不给我。”
GEN|22|13|亚伯拉罕 举目观看，看哪，一只公绵羊两角缠在灌木丛中。 亚伯拉罕 就去牵了那只公绵羊，献为燔祭，代替他的儿子。
GEN|22|14|亚伯拉罕 给那地方起名叫“耶和华以勒” 。直到今日人还说：“在耶和华的山上必有预备。”
GEN|22|15|耶和华的使者第二次从天上呼唤 亚伯拉罕 ，
GEN|22|16|说：“耶和华说：‘你既行了这事，没有留下你的儿子，就是你的独子，我指着自己起誓：
GEN|22|17|我必多多赐福给你，我必使你的后裔大大增多，如同天上的星、海边的沙。你的后裔必得仇敌的城门，
GEN|22|18|并且地上的万国都必因你的后裔得福，因为你听从了我的话。’”
GEN|22|19|于是 亚伯拉罕 回到他仆人那里。他们一同起身，往 别是巴 去， 亚伯拉罕 就住在 别是巴 。
GEN|22|20|这些事以后，有人告诉 亚伯拉罕 说：“看哪， 密迦 也为你兄弟 拿鹤 生了几个儿子：
GEN|22|21|长子 乌斯 、他的兄弟 布斯 、 亚兰 的父亲 基摩利 、
GEN|22|22|基薛 、 哈琐 、 必达 、 益拉 和 彼土利 。”
GEN|22|23|彼土利 生 利百加 。这八个人都是 密迦 为 亚伯拉罕 的兄弟 拿鹤 生的。
GEN|22|24|拿鹤 的妾名叫 流玛 ，她也生了 提八 、 迦含 、 他辖 和 玛迦 。
GEN|23|1|撒拉 享寿一百二十七岁，这是 撒拉 一生的岁数 。
GEN|23|2|撒拉 死在 迦南 地的 基列．亚巴 ，就是 希伯仑 。 亚伯拉罕 来哀悼 撒拉 ，为她哭泣。
GEN|23|3|然后， 亚伯拉罕 起来，离开死人面前，对 赫 人说：
GEN|23|4|“我在你们中间是外人，是寄居的。请给我你们那里的一块坟地，我好埋葬我的亡妻，使她不在我的面前。”
GEN|23|5|赫 人回答 亚伯拉罕 说：
GEN|23|6|“我主请听。你在我们中间是一位尊贵的王子，只管在我们最好的坟地里埋葬你的死人；我们没有一人会拒绝你在他的坟地里埋葬你的死人。”
GEN|23|7|于是， 亚伯拉罕 起来，向当地的百姓 赫 人下拜，
GEN|23|8|对他们说：“你们若愿意让我埋葬我的亡妻，使她不在我面前，就请听我，为我求 琐辖 的儿子 以弗仑 ，
GEN|23|9|把他田地尽头的 麦比拉洞 卖给我。他可以按照足价卖给我，作为我在你们中间的坟地。”
GEN|23|10|那时， 以弗仑 正坐在 赫 人中间。 赫 人 以弗仑 就回答 亚伯拉罕 ，说给所有出入城门的 赫 人听：
GEN|23|11|“不，我主请听。我要把这块田送给你，连田间的洞也送给你，在我同族的人眼前都给你，让你埋葬你的死人。”
GEN|23|12|亚伯拉罕 就在当地的百姓面前下拜，
GEN|23|13|对 以弗仑 说，也给当地百姓听：“你若应允，请你听我。我要把田的价钱给你，请你收下，我就在那里埋葬我的死人。”
GEN|23|14|以弗仑 回答 亚伯拉罕 说：
GEN|23|15|“我主请听。四百舍客勒银子的地，在你我中间算什么呢？只管埋葬你的死人吧！”
GEN|23|16|亚伯拉罕 听从了 以弗仑 。 亚伯拉罕 就照着他说给 赫 人听的，把买卖通用的银子，秤了四百舍客勒银子给 以弗仑 。
GEN|23|17|于是， 以弗仑 把那块位于 幔利 对面的 麦比拉 田，和其中的洞，以及田间周围的树木都成交了，
GEN|23|18|在所有出入城门的 赫 人眼前，卖给 亚伯拉罕 作为他的产业。
GEN|23|19|后来， 亚伯拉罕 把他妻子 撒拉 安葬在 迦南 地 幔利 对面的 麦比拉 田间的洞里， 幔利 就是 希伯仑 。
GEN|23|20|从此，那块田和田间的洞就从 赫 人移交给 亚伯拉罕 作坟地的产业。
GEN|24|1|亚伯拉罕 年纪老迈，耶和华在一切事上都赐福给他。
GEN|24|2|亚伯拉罕 对他家中管理他一切产业最老的仆人说：“把你的手放在我大腿底下。
GEN|24|3|我要叫你指着耶和华—天和地的上帝起誓，不要为我儿子娶我所居住的 迦南 地的女子为妻。
GEN|24|4|你要往我的本地本族去，为我的儿子 以撒 娶妻。”
GEN|24|5|仆人对他说：“如果那女子不肯跟我来到这地，我必须把你的儿子带回到你出来的地方吗？”
GEN|24|6|亚伯拉罕 对他说：“你要谨慎，不可带我儿子回那里去。
GEN|24|7|耶和华—天上的上帝曾带领我离开父家和本族的地，对我说话，向我起誓说：‘我要将这地赐给你的后裔。’他要差遣使者在你面前，你就可以从那里为我儿子娶妻。
GEN|24|8|倘若那女子不肯跟你来，我叫你起的誓就与你无关了，只是你不可带我的儿子回到那里去。”
GEN|24|9|仆人就把手放在他主人 亚伯拉罕 的大腿底下，为这事向他起誓。
GEN|24|10|那仆人从他主人的骆驼中取了十匹骆驼，他手中也带着他主人各样的贵重物品离开 ，起身往 美索不达米亚 去，到了 拿鹤 的城。
GEN|24|11|傍晚时，众女子出来打水，他就让骆驼跪在城外的水井旁。
GEN|24|12|他说：“耶和华—我主人 亚伯拉罕 的上帝啊，求你施恩给我的主人 亚伯拉罕 ，让我今日就遇见吧！
GEN|24|13|看哪，我站在井旁，城内居民的女子们正出来打水。
GEN|24|14|我向哪一个少女说：‘请你放下水瓶来，给我水喝’，她若说：‘请喝！我也给你的骆驼喝’，愿她作你所选定给你仆人 以撒 的妻。这样，我就知道你施恩给我的主人了。”
GEN|24|15|话还没说完，看哪， 利百加 肩头上扛着水瓶出来。 利百加 是 彼土利 所生的； 彼土利 是 亚伯拉罕 的兄弟 拿鹤 妻子 密迦 的儿子。
GEN|24|16|那少女容貌极其美丽，是未曾与人亲近的童女。她下到井旁，打满了瓶子的水，就上来。
GEN|24|17|仆人跑上前去迎着她，说：“请你让我喝你瓶子里的一点水。”
GEN|24|18|少女说：“我主请喝！”就急忙拿下瓶子托在手上，给他喝水。
GEN|24|19|那少女给他喝足了，又说：“我也为你的骆驼打水，直到骆驼喝足了。”
GEN|24|20|她就急忙把瓶子里的水倒在槽里，又跑到井旁打水，为所有的骆驼打了水。
GEN|24|21|那人定睛看着少女，一句话也不说，要知道耶和华是否使他的道路亨通。
GEN|24|22|骆驼喝足了，那人就拿出一个比加 重的金环，一对十舍客勒重的金手镯，
GEN|24|23|说：“请告诉我，你是谁的女儿？你父亲家里有没有地方可以让我们过夜？”
GEN|24|24|少女说：“我是 密迦 为 拿鹤 生的儿子 彼土利 的女儿。”
GEN|24|25|又说：“我们家里有充足的干草和饲料，也有住宿的地方。”
GEN|24|26|那人就低头向耶和华敬拜，
GEN|24|27|说：“耶和华—我主人 亚伯拉罕 的上帝是应当称颂的，因他不断以慈爱信实待我主人。至于我，耶和华一路引领我，直到我主人的兄弟家里。”
GEN|24|28|那少女跑去，把这些话告诉她母亲家里的人。
GEN|24|29|利百加 有一个哥哥，名叫 拉班 ， 拉班 就跑到外面井旁那人那里。
GEN|24|30|当他看见金环和戴在他妹妹手上的金镯，又听见他妹妹 利百加 说的话：“那人如此对我说”，他就来到那人面前，看哪，他还站在井旁的骆驼旁边，
GEN|24|31|就对他说：“你这蒙耶和华赐福的人，请进来吧！为什么站在外面？我已经收拾了房屋，也为骆驼预备了地方。”
GEN|24|32|那人就进了 拉班 的家。 拉班 卸了骆驼，用饲料喂它们，拿水给那人和随从他的人洗脚，
GEN|24|33|把食物摆在他面前，请他吃。他却说：“我不吃，等我把我的事情说完了再吃。” 拉班 说：“请说。”
GEN|24|34|他说：“我是 亚伯拉罕 的仆人。
GEN|24|35|耶和华大大地赐福给我主人，使他发达，赐给他羊群、牛群、金银、奴仆、婢女、骆驼和驴。
GEN|24|36|我主人的妻子 撒拉 年老的时候为我主人生了一个儿子；我主人把他一切所有的都给了他。
GEN|24|37|我主人叫我起誓说：‘不要为我儿子娶我所居住的 迦南 地的女子为妻。
GEN|24|38|你要往我父家、我本族那里去，为我的儿子娶妻。’
GEN|24|39|我对我主人说：‘恐怕那女子不肯跟我来。’
GEN|24|40|他就说：‘我所事奉的耶和华必要差遣他的使者与你同去，使你的道路亨通，你就可以在我父家、我本族那里，为我的儿子娶妻。
GEN|24|41|只要你到了我本族那里，我叫你起的誓就与你无关。他们若不把女子交给你，我叫你起的誓也与你无关。’
GEN|24|42|“我今日到了井旁，就说：‘耶和华—我主人 亚伯拉罕 的上帝啊，愿你使我所行的道路亨通。
GEN|24|43|看哪，我站在井旁，对哪一个出来打水的女子说：请你让我喝你瓶子里的一点水，
GEN|24|44|她若说：你只管喝，我也为你的骆驼打水；愿那女子作耶和华给我主人儿子所选定的妻子。’
GEN|24|45|“我心里的话还没有说完，看哪， 利百加 肩头上扛着水瓶出来，下到井旁打水。我对她说：‘请你给我水喝。’
GEN|24|46|她就急忙从肩头上拿下瓶子来，说：‘请喝！我也给你的骆驼喝。’我就喝了；她也给我的骆驼喝了。
GEN|24|47|我问她说：‘你是谁的女儿？’她说：‘我是 彼土利 的女儿， 彼土利 是 密迦 和 拿鹤 生的儿子。’我就把环子戴在她鼻子上，把镯子戴在她双手上。
GEN|24|48|然后我低头向耶和华敬拜，称颂耶和华—我主人 亚伯拉罕 的上帝，因为他引导我走合适的道路，使我得着我主人兄弟的孙女，给我主人的儿子为妻。
GEN|24|49|现在你们若愿以慈爱诚信待我主人，就告诉我；若不然，也告诉我，使我可以或向左，或向右。”
GEN|24|50|拉班 和 彼土利 回答说：“这事既然出于耶和华，我们不能向你说好说歹。
GEN|24|51|看哪， 利百加 就在你面前，可以将她带去，遵照耶和华所说的，给你主人的儿子为妻。”
GEN|24|52|亚伯拉罕 的仆人听见他们这些话，就向耶和华俯伏在地。
GEN|24|53|仆人拿出金器、银器和衣服送给 利百加 ，又将贵重的物品送给她哥哥和她母亲。
GEN|24|54|然后，仆人和随从的人才吃喝，并且住了一夜。早晨起来，仆人说：“请让我回我主人那里去吧。”
GEN|24|55|利百加 的哥哥和母亲说：“让她同我们再住几天，也许十天，然后她可以去。”
GEN|24|56|仆人对他们说：“耶和华既然使我道路亨通，你们就不要耽误我，请让我走，回我主人那里去吧！”
GEN|24|57|他们说：“我们把她叫来问问她 。”
GEN|24|58|他们就叫了 利百加 来，对她说：“你和这人同去吗？”她说：“我去。”
GEN|24|59|于是他们送他们的妹妹 利百加 和她的奶妈，同 亚伯拉罕 的仆人，以及随从他的人走了。
GEN|24|60|他们就为 利百加 祝福，对她说： “我们的妹妹啊， 愿你作千万人的母亲！ 愿你的后裔得着仇敌的城门！”
GEN|24|61|利百加 和她的女仆们起来，骑上骆驼，跟着那人去。仆人就带着 利百加 走了。
GEN|24|62|那时， 以撒 住在 尼革夫 。他刚从 庇耳．拉海．莱 回来。
GEN|24|63|傍晚时， 以撒 出来，到田间默想。他举目一看，看哪，来了一队骆驼。
GEN|24|64|利百加 举目看见 以撒 ，就急忙下了骆驼，
GEN|24|65|对那仆人说：“这从田间走来迎接我们的人是谁？”仆人说：“他是我的主人。” 利百加 就拿面纱盖住自己。
GEN|24|66|仆人把他所做的一切事都告诉 以撒 。
GEN|24|67|以撒 就领 利百加 进了母亲 撒拉 的帐棚，娶了她为妻，并且爱她。 以撒 自从母亲离世以后，这才得了安慰。
GEN|25|1|亚伯拉罕 再娶了一个妻子，名叫 基土拉 。
GEN|25|2|她为他生了 心兰 、 约珊 、 米但 、 米甸 、 伊施巴 和 书亚 。
GEN|25|3|约珊 生了 示巴 和 底但 。 底但 的子孙是 亚书利 族、 利都是 族和 利乌米 族。
GEN|25|4|米甸 的儿子是 以法 、 以弗 、 哈诺 、 亚比大 和 以勒大 。这些都是 基土拉 的子孙。
GEN|25|5|亚伯拉罕 把他一切所有的都给了 以撒 。
GEN|25|6|至于 亚伯拉罕 妾的儿子， 亚伯拉罕 趁着自己还活着的时候把财物分给他们，打发他们离开他的儿子 以撒 ，往东方去，直到东方之地。
GEN|25|7|这是 亚伯拉罕 一生的年日，他活了一百七十五年。
GEN|25|8|亚伯拉罕 寿高年迈，安享天年，息劳而终，归到他祖先 那里。
GEN|25|9|他两个儿子 以撒 、 以实玛利 把他安葬在 麦比拉 洞里。这洞在 幔利 的对面、 赫 人 琐辖 的儿子 以弗仑 的田中，
GEN|25|10|就是 亚伯拉罕 向 赫 人买的那块田。 亚伯拉罕 和他妻子 撒拉 都葬在那里。
GEN|25|11|亚伯拉罕 死了以后，上帝赐福给他的儿子 以撒 。 以撒 住在 庇耳．拉海．莱 附近。
GEN|25|12|这是 撒拉 的婢女、 埃及 人 夏甲 为 亚伯拉罕 生的儿子 以实玛利 的后代。
GEN|25|13|以实玛利 儿子们的名字，按着他们后代的名字如下： 以实玛利 的长子 尼拜约 ，又有 基达 、 亚德别 、 米比衫 、
GEN|25|14|米施玛 、 度玛 、 玛撒 、
GEN|25|15|哈大 、 提玛 、 伊突 、 拿非施 ，和 基底玛 。
GEN|25|16|这些都是 以实玛利 的儿子们。他们的村庄和营寨按着他们命名；他们作了十二族的族长。
GEN|25|17|以实玛利 一生的岁数是一百三十七岁，断气而死，归到他祖先那里。
GEN|25|18|他的子孙住在 哈腓拉 ，直到 埃及 东边的 书珥 ，向着 亚述 ，在他众弟兄的对面安顿下来 。
GEN|25|19|这是 亚伯拉罕 的儿子 以撒 的后代。 亚伯拉罕 生 以撒 。
GEN|25|20|以撒 四十岁时娶 利百加 为妻。 利百加 是 巴旦．亚兰 地的 亚兰 人 彼土利 的女儿，是 亚兰 人 拉班 的妹妹。
GEN|25|21|以撒 因他妻子不生育，就为她祈求耶和华。耶和华应允他的祈求，他的妻子 利百加 就怀了孕。
GEN|25|22|胎儿们在她腹中彼此相争，她就说：“若是如此，我为什么会这样呢 ？”她就去求问耶和华。
GEN|25|23|耶和华对她说： 两国在你腹中； 两族要从你身上分立。 这族必强于那族； 将来大的要服侍小的。
GEN|25|24|到了生产的日期，看哪，腹中是对双胞胎。
GEN|25|25|先出生的身体带红，浑身有毛，好像皮衣；他们就给他起名叫 以扫 。
GEN|25|26|随后， 以扫 的弟弟也出生，他的手抓住 以扫 的脚跟，因此给他起名叫 雅各 。两个儿子出生时， 以撒 六十岁。
GEN|25|27|两个孩子渐渐长大， 以扫 善于打猎，常在田野； 雅各 为人安静，常住在帐棚里。
GEN|25|28|以撒 爱 以扫 ，因为常吃他的野味； 利百加 却爱 雅各 。
GEN|25|29|有一天， 雅各 熬了汤， 以扫 从田野回来，疲惫不堪。
GEN|25|30|以扫 对 雅各 说：“我累死了，请你让我吃这红的，这红的汤吧！”因此 以扫 又叫 以东 。
GEN|25|31|雅各 说：“你今日把长子的名分卖给我吧。”
GEN|25|32|以扫 说：“看哪，我快要死了，这长子的名分对我有什么用呢？”
GEN|25|33|雅各 说：“你今日对我起誓吧。” 以扫 就向他起誓，把长子的名分卖给了 雅各 。
GEN|25|34|于是 雅各 把饼和豆汤给了 以扫 ， 以扫 吃喝以后，起来走了。这样， 以扫 轻看他长子的名分。
GEN|26|1|那地有了饥荒，不是 亚伯拉罕 的时候曾有过的那次饥荒， 以撒 就到 基拉耳 ， 非利士 人的王 亚比米勒 那里去。
GEN|26|2|耶和华向 以撒 显现，说：“你不要下 埃及 去，要住在我所指示你的地。
GEN|26|3|你要寄居在这地，我必与你同在，赐福给你，因为我要将这一切的地都赐给你和你的后裔。我必坚定我向你父亲 亚伯拉罕 所起的誓。
GEN|26|4|我要使你的后裔增多，好像天上的星，又要将这一切的地赐给你的后裔，并且地上的万国都必因你的后裔得福，
GEN|26|5|因为 亚伯拉罕 听从我的话，遵守我的吩咐、诫令、律例和教导。”
GEN|26|6|于是， 以撒 住在 基拉耳 。
GEN|26|7|那地方的人问起他的妻子，他就说：“她是我的妹妹。”原来他害怕说“我的妻子”。他想：“或许这地方的人会因 利百加 杀我，因为她容貌美丽。”
GEN|26|8|他在那里住了一段很长的日子。有一天， 非利士 人的王 亚比米勒 从窗户往外观看，看哪， 以撒 在抚爱他的妻子 利百加 。
GEN|26|9|亚比米勒 召 以撒 来，说：“看哪，她实在是你的妻子，你怎么说‘她是我的妹妹’呢？” 以撒 对他说：“因为我想，恐怕我会因她而死。”
GEN|26|10|亚比米勒 说：“你向我们做的是什么事呢？百姓中有一个人几乎要和你的妻子同寝，你就把我们陷在罪中了。”
GEN|26|11|于是 亚比米勒 命令众百姓说：“凡侵犯这个人，或他妻子的，必要把他处死。”
GEN|26|12|以撒 在那地耕种，那一年有百倍的收成。耶和华赐福给他，
GEN|26|13|他就发达，日渐昌盛，成了大富翁。
GEN|26|14|他有羊群牛群，又有许多仆人， 非利士 人就嫉妒他。
GEN|26|15|他父亲 亚伯拉罕 在世的时候，他父亲的仆人所挖的井， 非利士 人全都塞住，填满了土。
GEN|26|16|亚比米勒 对 以撒 说：“你离开我们去吧，因为你比我们强盛得多。”
GEN|26|17|以撒 就离开那里，在 基拉耳谷 支搭帐棚，住在那里。
GEN|26|18|他父亲 亚伯拉罕 在世的时候所挖的水井，在 亚伯拉罕 死后，都被 非利士 人塞住了， 以撒 就重新把井挖出来，仍照他父亲所取的名为它们命名。
GEN|26|19|以撒 的仆人在谷中挖井，就在那里得了一口活水井。
GEN|26|20|基拉耳 的牧人与 以撒 的牧人相争，说：“这水是我们的。” 以撒 就给那井起名叫 埃色 ，因为他们和他相争。
GEN|26|21|以撒 的仆人又挖了一口井，他们又为这井相争， 以撒 就给这井起名叫 西提拿 。
GEN|26|22|以撒 离开那里，又挖了一口井，他们不再为这井相争了，他就给那井起名叫 利河伯 。他说：“耶和华现在给我们宽阔之地，我们必在这地兴旺。”
GEN|26|23|以撒 从那里上 别是巴 去。
GEN|26|24|当夜耶和华向他显现，说：“我是你父亲 亚伯拉罕 的上帝。不要惧怕，因为我与你同在，要赐福给你，也要为我仆人 亚伯拉罕 的缘故，使你的后裔增多。”
GEN|26|25|以撒 就在那里筑了一座坛，求告耶和华的名，并且在那里支搭帐棚；他的仆人就在那里挖了一口井。
GEN|26|26|亚比米勒 同他的顾问 亚户撒 和他军队的元帅 非各 ，从 基拉耳 来到 以撒 那里。
GEN|26|27|以撒 对他们说：“你们既然恨我，赶我离开你们，为什么又到我这里来呢？”
GEN|26|28|他们说：“我们明明看见耶和华与你同在；因此就说，让我们双方彼此起誓，我们跟你立约，
GEN|26|29|使你不加害我们，正如我们未曾侵犯你，素来善待你，并且送你平平安安地走。你是蒙耶和华赐福的！”
GEN|26|30|以撒 为他们摆设宴席，他们就一起吃喝。
GEN|26|31|他们清早起来，彼此起誓。 以撒 送他们走，他们就平平安安地离开他去了。
GEN|26|32|那一天， 以撒 的仆人来，把挖井的消息告诉他，说：“我们得到水了。”
GEN|26|33|他就给那井起名叫 示巴 ，因此那城名叫 别是巴 ，直到今日。
GEN|26|34|以扫 四十岁的时候娶了 赫 人 比利 的女儿 犹滴 ，和 赫 人 以伦 的女儿 巴实抹 为妻。
GEN|26|35|她们使 以撒 和 利百加 心里愁烦。
GEN|27|1|以撒 年老，眼睛昏花，不能看见，就叫他大儿子 以扫 来，对他说：“我儿。” 以扫 对他说：“我在这里。”
GEN|27|2|他说：“看哪，我老了，不知道哪一天死。
GEN|27|3|现在拿你打猎的工具，就是箭囊和弓，到田野去为我打猎，
GEN|27|4|照我所爱的做成美味，拿来给我吃，好让我在未死之前为你祝福。”
GEN|27|5|以撒 对他儿子 以扫 说话的时候， 利百加 听见了。 以扫 往田野去打猎，要把猎物带回来。
GEN|27|6|利百加 就对她儿子 雅各 说：“看哪，我听见你父亲对你哥哥 以扫 说：
GEN|27|7|‘你去把猎物带回来，做成美味给我吃，让我在未死之前，在耶和华面前为你祝福。’
GEN|27|8|现在，我儿，你要听我的话，照我所吩咐你的，
GEN|27|9|到羊群里去，从那里牵两只肥美的小山羊来给我，我就照你父亲所爱的，把它们做成美味给他。
GEN|27|10|然后，你拿到你父亲那里给他吃，好让他在未死之前为你祝福。”
GEN|27|11|雅各 对他母亲 利百加 说：“看哪，我哥哥 以扫 浑身都有毛，我身上却是光滑的；
GEN|27|12|倘若父亲摸着我，我在他眼中就是骗子了。这样，我就自招诅咒，而不是祝福。”
GEN|27|13|他母亲对他说：“我儿，你所受的诅咒临到我身上吧！你只管听我的话，去牵小山羊来给我。”
GEN|27|14|他就去牵来，交给他母亲。他母亲就照他父亲所爱的，做成美味。
GEN|27|15|利百加 把大儿子 以扫 在家里最好的衣服给她小儿子 雅各 穿，
GEN|27|16|又用小山羊的皮包在 雅各 的手上和颈项光滑的地方，
GEN|27|17|就把所做的美味和饼交在她儿子 雅各 的手里。
GEN|27|18|雅各 来到他父亲那里，说：“我的父亲！”他说：“我在这里。我儿，你是谁？”
GEN|27|19|雅各 对他父亲说：“我是你的长子 以扫 。我已照你吩咐我的做了。请起来坐着，吃我的野味，你好为我祝福。”
GEN|27|20|以撒 对他儿子说：“我儿，你怎么这样快就找到了呢？”他说：“因为这是耶和华—你的上帝使我遇见的。”
GEN|27|21|以撒 对 雅各 说：“我儿，靠近一点，让我摸摸你，你真的是我的儿子 以扫 吗？”
GEN|27|22|雅各 就靠近他父亲 以撒 。 以撒 摸着他，说：“声音是 雅各 的声音，手却是 以扫 的手。”
GEN|27|23|以撒 认不出他来，因为他手上有毛，像他哥哥 以扫 的手一样。于是， 以撒 就为他祝福。
GEN|27|24|以撒 说：“你真的是我儿子 以扫 吗？”他说：“我是。”
GEN|27|25|以撒 说：“拿给我，让我吃我儿子的野味，我好为你祝福。” 雅各 拿给他，他就吃了，又拿酒给他，他也喝了。
GEN|27|26|他父亲 以撒 对他说：“我儿，靠近一点来亲我！”
GEN|27|27|他就近前亲吻父亲。他父亲一闻他衣服上的香气，就为他祝福，说： “看，我儿的香气 好像耶和华赐福之田地的香气。
GEN|27|28|愿上帝赐你天上的甘露， 地上的肥土， 和丰富的五谷新酒。
GEN|27|29|愿万民事奉你， 万族向你下拜。 愿你作你弟兄的主， 你母亲的儿子向你下拜。 诅咒你的，愿他受诅咒； 祝福你的，愿他蒙祝福。”
GEN|27|30|以撒 为 雅各 祝福完毕， 雅各 才从他父亲那里出来，他哥哥 以扫 正打猎回来。
GEN|27|31|以扫 也做了美味，拿来给他父亲，对他父亲说：“父亲，请起来，吃你儿子的野味，你好为我祝福。”
GEN|27|32|他父亲 以撒 对他说：“你是谁？”他说：“我是你的儿子，你的长子 以扫 。”
GEN|27|33|以撒 就大大战兢，说：“那么，是谁打了猎物拿来给我呢？你未来之前我已经吃了，也为他祝福了，他将来就必蒙福。”
GEN|27|34|以扫 听了他父亲的话，就大声痛哭，对他父亲说：“我父啊，求你也为我祝福！”
GEN|27|35|以撒 说：“你弟弟已经用诡计来把你的福分夺去了。”
GEN|27|36|以扫 说：“他名叫 雅各 ，岂不是这样吗？他欺骗了我两次：他先前夺了我长子的名分，看哪，他现在又夺了我的福分。” 以扫 又说：“你没有留下给我的祝福吗？”
GEN|27|37|以撒 回答 以扫 说：“看哪，我已立他作你的主，使他的弟兄都给他作仆人，并赐他五谷新酒可以养生。我儿，那么，现在我还能为你做什么呢？”
GEN|27|38|以扫 对他父亲说：“我父啊，你只有一个祝福吗？我父啊，求你也为我祝福！” 以扫 就放声而哭。
GEN|27|39|他父亲 以撒 回答说： “看哪，你所住的地方必缺乏肥沃的土地， 缺乏天上的甘露 。
GEN|27|40|你必倚靠刀剑度日， 又必服侍你的兄弟； 到你强盛的时候， 必从你颈项上挣开他的轭。
GEN|27|41|以扫 因他父亲给 雅各 的祝福，就怨恨 雅各 ，心里说：“为我父亲居丧的时候近了，到那时候，我要杀我的弟弟 雅各 。”
GEN|27|42|有人把 利百加 大儿子 以扫 的话告诉 利百加 ，她就派人去，叫了她小儿子 雅各 来，对他说：“看哪，你哥哥 以扫 想要杀你来泄恨。
GEN|27|43|现在，我儿，听我的话，起来，逃往 哈兰 ，到我哥哥 拉班 那里去，
GEN|27|44|同他住一段日子，直等到你哥哥的怒气消了。
GEN|27|45|等到你哥哥向你消了怒气，忘了你向他所做的事，我就派人去，把你从那里带回来。我何必在一天之内丧失你们二人呢？”
GEN|27|46|利百加 对 以撒 说：“我因这 赫 人的女子活得不耐烦了；倘若 雅各 也从本地女子中娶像这样的 赫 人女子为妻，我为什么要活着呢？”
GEN|28|1|以撒 叫了 雅各 来，为他祝福，并吩咐他说：“你不要娶 迦南 的女子为妻。
GEN|28|2|你起身往 巴旦．亚兰 去，到你外祖父 彼土利 的家，从你舅父 拉班 的女儿中娶一位作你的妻子。
GEN|28|3|愿全能的上帝赐福给你，使你生养众多，成为许多民族，
GEN|28|4|将应许 亚伯拉罕 的福赐给你和你的后裔，使你承受你所寄居的地为业，就是上帝赐给 亚伯拉罕 的地。”
GEN|28|5|以撒 送 雅各 走了， 雅各 就往 巴旦．亚兰 去，到 亚兰 人 彼土利 的儿子 拉班 那里， 拉班 是 利百加 的哥哥， 利百加 是 雅各 和 以扫 的母亲。
GEN|28|6|以扫 见 以撒 已经为 雅各 祝福，而且送他往 巴旦．亚兰 去，在那里娶妻，并且见 以撒 祝福 雅各 的时候吩咐他说：“不要娶 迦南 的女子为妻”，
GEN|28|7|又见 雅各 听从父母的话往 巴旦．亚兰 去了，
GEN|28|8|以扫 就看出他父亲 以撒 看 迦南 女子不顺眼。
GEN|28|9|于是他往 以实玛利 那里去，在两个妻子之外， 又娶了 玛哈拉 为妻，她是 亚伯拉罕 儿子 以实玛利 的女儿，是 尼拜约 的妹妹。
GEN|28|10|雅各 离开 别是巴 ，往 哈兰 去。
GEN|28|11|到了一个地方，因为已经日落，就在那里过夜。他拾起那地方的一块石头枕在头下，就躺在那地方。
GEN|28|12|他做梦，看哪，一个梯子立在地上，梯子的顶端直伸到天；看哪，上帝的使者在梯子上，上去下来。
GEN|28|13|看哪，耶和华站在梯子上面 ，说：“我是耶和华—你祖父 亚伯拉罕 的上帝， 以撒 的上帝。你现在躺卧之地，我要将它赐给你和你的后裔。
GEN|28|14|你的后裔必像地上的尘沙，必向东西南北开展；地上万族必因你和你的后裔得福。
GEN|28|15|看哪，我必与你同在，无论你往哪里去，我必保佑你，领你归回这地。我总不离弃你，直到我实现了对你所说的话。”
GEN|28|16|雅各 睡醒了，说：“耶和华真的在这里，我竟不知道！”
GEN|28|17|他就惧怕，说：“这地方何等可畏！这不是别的，是上帝的殿，是天的门。”
GEN|28|18|雅各 清早起来，拿起枕在头下的石头，立作柱子，浇油在上面。
GEN|28|19|他给那地方起名叫 伯特利 ；那地方原先名叫 路斯 。
GEN|28|20|雅各 许愿说：“上帝若与我同在，在我所行的路上保佑我，给我食物吃，衣服穿，
GEN|28|21|使我平平安安回到我父亲的家，我就必以耶和华为我的上帝。
GEN|28|22|我所立为柱子的这块石头必作上帝的殿；凡你所赐给我的，我必将十分之一献给你。”
GEN|29|1|雅各 起行，到了东方人之地。
GEN|29|2|他观看，看哪，田间有一口井，看哪，有三群羊卧在井旁；因为人都取那井里的水给羊喝。井口上的那块石头很大。
GEN|29|3|羊群都在那里聚集，人就把石头移开井口，取水给羊喝，然后又把石头放回井口原处。
GEN|29|4|雅各 对他们说：“弟兄们，你们从哪里来？”他们说：“我们是从 哈兰 来的。”
GEN|29|5|他对他们说：“你们认识 拿鹤 的孙子 拉班 吗？”他们说：“我们认识。”
GEN|29|6|雅各 对他们说：“他平安吗？”他们说：“平安。看哪，他女儿 拉结 和羊一起来了。”
GEN|29|7|雅各 说：“看哪，日正当中，不是牲畜聚集的时候。你们取水给羊喝，再去牧放吧！”
GEN|29|8|他们说：“我们不能这样，必须等所有的羊群聚集，人把石头移开井口，我们才可以取水给羊喝。”
GEN|29|9|雅各 正和他们说话的时候， 拉结 和她父亲的羊来了，因为她是牧羊的。
GEN|29|10|雅各 看见他舅父 拉班 的女儿 拉结 和舅父 拉班 的羊群，就上前把石头移开井口，取水给舅父 拉班 的羊喝。
GEN|29|11|雅各 亲了 拉结 ，就放声大哭。
GEN|29|12|雅各 告诉 拉结 ，自己是她父亲的亲戚 ，是 利百加 的儿子。 拉结 就跑去告诉她父亲。
GEN|29|13|拉班 听见外甥 雅各 的消息，就跑去迎接他，抱着他，亲他，带他到自己的家。 雅各 把这一切的事告诉 拉班 。
GEN|29|14|拉班 对他说：“你实在是我的骨肉。” 雅各 就和他同住了一个月。
GEN|29|15|拉班 对 雅各 说：“虽然你是我的亲戚，怎么可以让你白白服事我呢？告诉我，你要什么作工资呢？”
GEN|29|16|拉班 有两个女儿，大的名叫 利亚 ，小的名叫 拉结 。
GEN|29|17|利亚 的双眼无神， 拉结 却长得美貌秀丽。
GEN|29|18|雅各 爱 拉结 ，就说：“我愿为你的小女儿 拉结 服事你七年。”
GEN|29|19|拉班 说：“我把她给你，胜过给别人，你与我同住吧！”
GEN|29|20|雅各 就为 拉结 服事了七年；他因为爱 拉结 ，就看这七年如同几天。
GEN|29|21|雅各 对 拉班 说：“日期已经满了，请把我的妻子给我，我好与她同房。”
GEN|29|22|拉班 就摆设宴席，请了当地所有的人。
GEN|29|23|到了晚上， 拉班 带女儿 利亚 来送给 雅各 ， 雅各 就与她同房。
GEN|29|24|拉班 也把自己的婢女 悉帕 给女儿 利亚 作婢女。
GEN|29|25|到了早晨，看哪，她是 利亚 ， 雅各 对 拉班 说：“你向我做的是什么事呢？我服事你，不是为 拉结 吗？你为什么欺骗我呢？”
GEN|29|26|拉班 说：“大女儿还没有给人就先把小女儿给人，我们这地方没有这样的规矩。
GEN|29|27|你先为这个满了七日，我们就把那个也给你，不过你要另外再服事我七年。”
GEN|29|28|雅各 就这样做了。满了 利亚 的七日， 拉班 就把女儿 拉结 给 雅各 为妻。
GEN|29|29|拉班 又把自己的婢女 辟拉 给女儿 拉结 作婢女。
GEN|29|30|雅各 也与 拉结 同房，并且爱 拉结 胜过爱 利亚 ，于是他又服事了 拉班 七年。
GEN|29|31|耶和华见 利亚 失宠 ，就使她生育， 拉结 却不生育。
GEN|29|32|利亚 怀孕生子，给他起名叫 吕便 ，因为她说：“耶和华看见我的苦情，如今我的丈夫必爱我。”
GEN|29|33|她又怀孕生子，给他起名叫 西缅 ，说：“耶和华因为听见我失宠，所以又赐给我这个儿子。”
GEN|29|34|她又怀孕生子，说：“我给丈夫生了三个儿子，现在，这次他必亲近我了。”因此， 雅各 给他起名叫 利未 。
GEN|29|35|她又怀孕生子，说：“这次我要赞美耶和华。”因此给他起名叫 犹大 。于是她停了生育。
GEN|30|1|拉结 见自己不给 雅各 生孩子，就嫉妒她姊姊，对 雅各 说：“你给我孩子，不然，让我死了吧。”
GEN|30|2|雅各 对 拉结 生气，说：“是我代替上帝使你生不出孩子的吗？”
GEN|30|3|拉结 说：“看哪，我的使女 辟拉 在这里，你可以与她同房，使她生子归在我膝下，我也可以藉着她得孩子 。”
GEN|30|4|拉结 就把她的婢女 辟拉 给丈夫为妾， 雅各 与她同房。
GEN|30|5|辟拉 怀孕，为 雅各 生了一个儿子。
GEN|30|6|拉结 给他起名叫 但 ，说：“上帝为我伸冤，也听了我的声音，赐给我一个儿子。”
GEN|30|7|拉结 的婢女 辟拉 又怀孕，为 雅各 生了第二个儿子。
GEN|30|8|拉结 给他起名叫 拿弗他利 ，说：“我与我姊姊大大较力，并且得胜了。”
GEN|30|9|利亚 见自己停了生育，就把她的婢女 悉帕 给 雅各 为妾。
GEN|30|10|利亚 的婢女 悉帕 为 雅各 生了一个儿子。
GEN|30|11|利亚 给他起名叫 迦得 ，说：“真是幸运！”
GEN|30|12|利亚 的婢女 悉帕 又为 雅各 生了第二个儿子。
GEN|30|13|利亚 给他起名叫 亚设 ，说：“我真有福啊，众女子都要称我有福。”
GEN|30|14|收割麦子的时候， 吕便 到田里去，找到曼陀罗草 ，就拿给他的母亲 利亚 。 拉结 对 利亚 说：“请你给我一些你儿子的曼陀罗草吧。”
GEN|30|15|利亚 对她说：“你夺走了我的丈夫还是小事吗？你还要夺取我儿子的曼陀罗草吗？” 拉结 说：“今夜他可以与你同寝，来交换你儿子的曼陀罗草。”
GEN|30|16|到了晚上， 雅各 从田里回来， 利亚 出来迎接他，说：“你要与我同寝，因为我真的用我儿子的曼陀罗草把你雇下了。”那一夜， 雅各 就与她同寝。
GEN|30|17|上帝应允了 利亚 ，她就怀孕，为 雅各 生了第五个儿子。
GEN|30|18|利亚 给他起名叫 以萨迦 ，说：“上帝给了我工价，因为我把婢女给了我的丈夫。”
GEN|30|19|利亚 又怀孕，为 雅各 生了第六个儿子。
GEN|30|20|利亚 给他起名叫 西布伦 ，说：“上帝赐给我厚礼了；这次，我丈夫必看重我，因为我为他生了六个儿子。”
GEN|30|21|后来她又生了一个女儿，给她起名叫 底拿 。
GEN|30|22|上帝顾念 拉结 ，应允她，使她能生育。
GEN|30|23|拉结 怀孕生子，说：“上帝除去了我的羞耻。”
GEN|30|24|拉结 就给他起名叫 约瑟 ，说：“愿耶和华再增添一个儿子给我。”
GEN|30|25|拉结 生 约瑟 之后， 雅各 对 拉班 说：“请让我走，回到我的本乡本土去。
GEN|30|26|请你把我服事你所得的妻子和孩子给我，让我走吧！我怎样服事你，你都知道。”
GEN|30|27|拉班 对他说：“愿你看得起我，因我占卜得知，耶和华赐福给我是因你的缘故。”
GEN|30|28|又说：“请为我定你的工资，我就给你。”
GEN|30|29|雅各 对他说：“我怎样服事你，你的牲畜在我这里变得怎样，你都知道。
GEN|30|30|我未来以前，你拥有的很少，现在却已大量增加，因为耶和华随着我的脚步赐福给你。现在，我到什么时候才可以成家立业呢？”
GEN|30|31|拉班 说：“我该给你什么呢？” 雅各 说：“你什么也不必给我，只要你为我做这件事，我就继续牧放你的羊群。
GEN|30|32|今天我要走遍你的羊群，把绵羊中凡有点的、有斑的，和小绵羊中凡是黑色的羊；以及山羊中凡有斑的、有点的，都从那里挑出来，作为我的工资。
GEN|30|33|以后你来当面查看我的工资，任何我这里的山羊不是有点有斑的，小绵羊不是黑色的，就算是我偷的。这就可以证明我是正直的。”
GEN|30|34|拉班 说：“看哪，就照你所说的做吧。”
GEN|30|35|当日， 拉班 把有纹的、有斑的公山羊，一切有点的、有斑的、有少许白色 的母山羊，以及小绵羊中所有黑色的 ，都挑出来，交在他儿子们的手里，
GEN|30|36|又使自己和 雅各 相隔三天的路程。 雅各 就牧放 拉班 其余的羊。
GEN|30|37|雅各 拿杨树、杏树、枫树的嫩枝，把皮剥出白色的条纹，使枝子露出白色来。
GEN|30|38|他把剥了皮的枝子对着羊群，插在羊喝水的水沟和水槽里。羊来喝水的时候，它们彼此交配。
GEN|30|39|羊对着枝子交配，就生下有纹的、有点的、有斑的来。
GEN|30|40|雅各 把小绵羊分出来，让羊对着 拉班 羊群中有纹的和所有黑色的。于是他把自己的羊群分开，不叫它们和 拉班 的羊混在一起。
GEN|30|41|当肥壮的羊交配的时候， 雅各 就把枝子插在水沟里，使羊对着枝子交配。
GEN|30|42|可是当瘦弱的羊交配的时候，他就不插枝子。这样，瘦弱的就归 拉班 ，肥壮的就归 雅各 。
GEN|30|43|于是这人极其发达，拥有许多的羊群、奴仆、婢女、骆驼和驴。
GEN|31|1|雅各 听见 拉班 儿子们的话，说：“ 雅各 把我们父亲所有的都夺去了！他从我们父亲所拥有的获得这一切的财富。”
GEN|31|2|雅各 见 拉班 的脸色，看哪，待他不如从前了。
GEN|31|3|耶和华对 雅各 说：“你要回你祖先之地，到你本族那里去，我必与你同在。”
GEN|31|4|雅各 就派人叫 拉结 和 利亚 到田野他的羊群那里去，
GEN|31|5|对她们说：“我看你们父亲待我的脸色不如从前了，但我父亲的上帝向来与我同在。
GEN|31|6|你们也知道，我尽了全力服事你们的父亲。
GEN|31|7|可是你们的父亲欺骗我，十次更改我的工资，但上帝不容许他害我。
GEN|31|8|他若说：‘有点的归给你作工资’，羊群所生的都是有点的；他若说：‘有纹的归给你作工资’，羊群所生的都是有纹的。
GEN|31|9|这样，上帝把你们父亲的牲畜拿来赐给我了。
GEN|31|10|“羊群交配的时候，我在梦中举目一看，看哪，跳母羊的公羊都是有纹的、有点的、有花斑的。
GEN|31|11|上帝的使者在梦中呼叫我说：‘ 雅各 。’我说：‘我在这里。’
GEN|31|12|他说：‘你举目观看，跳母羊的公羊都是有纹的、有点的、有花斑的。 拉班 向你所做的一切，我都看见了。
GEN|31|13|我是 伯特利 的上帝；你曾在那里用油膏过柱子，向我许过愿。现在你起来，离开这地，回你本族之地去吧！’”
GEN|31|14|拉结 和 利亚 回答 雅各 说：“在我们父亲家里还有我们可分得的产业吗？
GEN|31|15|我们不是被他看作外人吗？因为他卖了我们，还吞吃了我们的银钱。
GEN|31|16|上帝从我们父亲所拿走的一切财物，都是我们和我们孩子的。现在，凡上帝所吩咐你的，你只管去做吧！”
GEN|31|17|雅各 起来，叫他的孩子和妻子都骑上骆驼，
GEN|31|18|又赶着他一切的牲畜和他所得的一切财物，就是他在 巴旦．亚兰 所得的，他拥有的牲畜 ，往 迦南 地他父亲 以撒 那里去了。
GEN|31|19|当时 拉班 去剪羊毛， 拉结 偷了他父亲家中的神像。
GEN|31|20|雅各 瞒住 亚兰 人 拉班 ，不通知他就逃走了。
GEN|31|21|雅各 带着他所有的逃走了；他起程，渡过 大河 ，面向着 基列山 。
GEN|31|22|到第三天，有人告诉 拉班 ， 雅各 逃跑了。
GEN|31|23|拉班 带着他的弟兄们去追他，追了七天，就在 基列山 追上了。
GEN|31|24|夜间，上帝来到 亚兰 人 拉班 那里，在梦中对他说：“你要小心，不可对 雅各 说好说歹。”
GEN|31|25|拉班 追上 雅各 。 雅各 在山上支搭帐棚； 拉班 和他的弟兄们也在 基列山 上支搭帐棚。
GEN|31|26|拉班 对 雅各 说：“你做的是什么事呢？你瞒着我把我的女儿们带走，好像用刀剑掳去一般。
GEN|31|27|你为什么暗暗地逃跑，瞒着我，不通知我一声，叫我可以欢乐、唱歌、击鼓、弹琴送你回去呢？
GEN|31|28|为什么不容许我与外孙和女儿吻别呢？你现在所做的真是愚蠢！
GEN|31|29|我的手本有能力害你，只是你父亲的上帝昨夜对我说：‘你要小心，不可对 雅各 说好说歹。’
GEN|31|30|现在你既然这么想念你的父家，不得不去，为什么又偷了我的神明呢？”
GEN|31|31|雅各 回答 拉班 说：“因为我害怕，我想，恐怕你把你的女儿从我这里夺走。
GEN|31|32|至于你的神明，你若在谁那里搜出来，就不让谁活。当着我们弟兄面前，你认一认在我这里有什么东西是你的，你就拿去吧。”原来 雅各 并不知道 拉结 偷了神明。
GEN|31|33|拉班 进了 雅各 、 利亚 ，以及两个使女的帐棚，却没有找到，就从 利亚 的帐棚出来，进入 拉结 的帐棚。
GEN|31|34|拉结 拿了神像，藏在骆驼的鞍子里，自己坐在上面。 拉班 搜遍了那帐棚，并没有找到。
GEN|31|35|拉结 对她父亲说：“请我主不要生气，因为我恰有月事，不能在你面前起来。” 拉班 搜寻，却找不到神像。
GEN|31|36|于是 雅各 发怒，斥责 拉班 。 雅各 对 拉班 说：“我有什么过犯，有什么罪恶，你竟这样火速地追我？
GEN|31|37|你搜遍了我一切的物件，你找到什么呢？可以放在你我弟兄面前，叫他们在我们两个之间评评理。
GEN|31|38|我在你那里这二十年，你的母绵羊、母山羊没有掉过胎。你羊群中的公绵羊，我没有吃过；
GEN|31|39|被野兽撕裂的，我没有带来给你，是我自己赔偿的。无论是白日被偷的，或是黑夜被偷的，你都从我手中索取。
GEN|31|40|我常常白日受尽炎热，黑夜受尽寒霜，不得合眼入睡。
GEN|31|41|我这二十年在你家里，为你两个女儿服事了你十四年，为你的羊群服事了你六年，你却十次更改我的工资。
GEN|31|42|若不是我父亲 以撒 所敬畏的上帝，就是 亚伯拉罕 的上帝与我同在，你如今必定打发我空手而去。上帝看见我的苦情和我手的辛劳，就在昨夜责备了你。”
GEN|31|43|拉班 回答 雅各 说：“这两个女儿是我的女儿，这些孩子是我的孩子，这些羊群也都是我的羊群；凡你所看见的都是我的。我的女儿和她们所生的孩子，我今日还能对他们做什么呢？
GEN|31|44|现在，来吧！让我和你立约，作你我之间的证据。”
GEN|31|45|雅各 就拿一块石头立作柱子，
GEN|31|46|对弟兄们说：“大家来堆积石头。”他们拿石头堆成一堆，于是在那里，在石堆旁边吃喝。
GEN|31|47|拉班 称那石堆为 伊迦尔．撒哈杜他 ， 雅各 却称那石堆为 迦累得 。
GEN|31|48|拉班 说：“今日这石堆成为你我之间的证据。”因此这地方名叫 迦累得 ，
GEN|31|49|又叫 米斯巴 ，因为他说：“我们彼此离别以后，愿耶和华在你我中间鉴察 。
GEN|31|50|你若苦待我的女儿，或在我的女儿以外另娶妻，虽没有人在场，你看，有上帝在你我中间作证。”
GEN|31|51|拉班 又对 雅各 说：“看哪，这石堆，看哪，这柱子，是我在你我中间所立的。
GEN|31|52|这石堆是证据，这柱子也是证据。我必不越过这石堆去害你；你也不可越过这石堆和柱子来害我。
GEN|31|53|愿 亚伯拉罕 的上帝和 拿鹤 的上帝，就是他们父亲的上帝 ，在你我中间判断。” 雅各 就指着他父亲 以撒 所敬畏的上帝起誓，
GEN|31|54|又在山上献祭，请弟兄们来吃饭。他们吃了饭，就在山上过夜。
GEN|31|55|拉班 清早起来，与他外孙和女儿亲吻，为他们祝福，就回到自己的地方去了。
GEN|32|1|雅各 继续行路，上帝的使者遇见他。
GEN|32|2|雅各 看见他们就说：“这是上帝的军营。”于是给那地方起名叫 玛哈念 。
GEN|32|3|雅各 派使者在他前面到 西珥 地，就是 以东 地他哥哥 以扫 那里。
GEN|32|4|他吩咐他们说：“你们要对我主 以扫 说：‘你的仆人 雅各 这样说：我在 拉班 那里寄居，延迟到如今。
GEN|32|5|我有牛、驴、羊群、奴仆、婢女，现在派人来报告我主，为了要在你眼前蒙恩。’”
GEN|32|6|使者回到 雅各 那里，说：“我们到了你哥哥 以扫 那里。他正迎着你来，并且有四百人和他一起。”
GEN|32|7|雅各 就很惧怕，而且愁烦。他把跟他同行的人和羊群、牛群、骆驼分成两队，
GEN|32|8|说：“ 以扫 若来击杀其中一队，剩下的另一队还可以逃脱。”
GEN|32|9|雅各 说：“耶和华—我祖父 亚伯拉罕 的上帝，我父亲 以撒 的上帝啊，你曾对我说：‘回你本地本族去，我要厚待你。’
GEN|32|10|你向仆人所施的一切慈爱和信实，我一点也不配得。我先前只用我的一根杖过这 约旦河 ，如今我却成了两队。
GEN|32|11|求你救我脱离我哥哥的手，脱离 以扫 的手，因为我怕他来杀我，连母亲和儿女都不放过。
GEN|32|12|你曾说：‘我必定厚待你，使你的后裔如同海边的沙，多得不可胜数。’”
GEN|32|13|当夜， 雅各 在那里住宿，就从他手中所拥有的拿礼物要送给他哥哥 以扫 ，
GEN|32|14|就是二百只母山羊、二十只公山羊、二百只母绵羊、二十只公绵羊、
GEN|32|15|三十匹哺乳的母骆驼和它们的小骆驼、四十头母牛、十头公牛、二十匹母驴和十匹公驴。
GEN|32|16|他把每种牲畜各分一群，交在仆人手中，对仆人说：“你们要在我的前头过去，使群和群之间保持一段距离”。
GEN|32|17|他又吩咐领头的人说：“我哥哥 以扫 遇见你的时候，问你说：‘你是谁的人？要往哪里去？你前面这些是谁的？’
GEN|32|18|你就说：‘是你仆人 雅各 的，是送给我主 以扫 的礼物。看哪，他自己也在我们后面。’”
GEN|32|19|他又吩咐第二、第三和所有赶畜群的人说：“你们遇见 以扫 的时候要照这样的话对他说，
GEN|32|20|你们还要说：‘看哪，你仆人 雅各 在我们后面。’”因 雅各 说：“我藉着在我前面送去的礼物给他面子，然后再见他的面，或许他会宽容我。”
GEN|32|21|于是礼物在他前面过去了；那夜， 雅各 在营中住宿。
GEN|32|22|他夜间起来，带着两个妻子，两个婢女和十一个孩子，过了 雅博 渡口。
GEN|32|23|他带着他们，送他们过河，他所有的一切也都过去，
GEN|32|24|只剩下 雅各 一人。有一个人来和他摔跤，直到黎明。
GEN|32|25|那人见自己胜不过他，就摸了他的大腿窝一下。 雅各 的大腿窝就在和那人摔跤的时候扭了。
GEN|32|26|那人说：“天快亮了，让我走吧！” 雅各 说：“你不给我祝福，我就不让你走。”
GEN|32|27|那人说：“你叫什么名字？”他说：“ 雅各 。”
GEN|32|28|那人说：“你的名字不要再叫 雅各 ，要叫 以色列 ，因为你与上帝和人较力，都得胜了。”
GEN|32|29|雅各 问他说：“请告诉我你的名字。”那人说：“何必问我的名字呢？”于是他在那里为 雅各 祝福。
GEN|32|30|雅各 就给那地方起名叫 毗努伊勒 ，说：“我面对面见了上帝，我的性命仍得保全。”
GEN|32|31|太阳刚出来的时候， 雅各 经过 毗努伊勒 ，他的大腿就瘸了。
GEN|32|32|因此， 以色列 人不吃大腿窝的筋，直到今日，因为那人摸了 雅各 大腿窝的筋。
GEN|33|1|雅各 举目观看，看哪， 以扫 来了，有四百人和他一起。 雅各 就把孩子们分开交给 利亚 、 拉结 和两个婢女。
GEN|33|2|他叫两个婢女和她们的孩子走在前头， 利亚 和她的孩子跟在后面，而 拉结 和 约瑟 在最后。
GEN|33|3|他自己却走到他们前面，一连七次俯伏在地才挨近他哥哥。
GEN|33|4|以扫 跑来迎接他，将他抱住，伏在他的颈项上亲他，他们都哭了。
GEN|33|5|以扫 举目看见妇人和孩子，就说：“这些和你一起的是谁呢？” 雅各 说：“这些孩子是上帝施恩给你仆人的。”
GEN|33|6|于是两个婢女和她们的孩子前来下拜，
GEN|33|7|利亚 和她的孩子也前来下拜，随后 约瑟 和 拉结 也前来下拜。
GEN|33|8|以扫 说：“我所遇见的这些畜群是什么意思呢？” 雅各 说：“是为了要在我主眼前蒙恩。”
GEN|33|9|以扫 说：“弟弟啊，我的已经够了，你的你自己留着吧！”
GEN|33|10|雅各 说：“不，我若在你眼前蒙恩，就请你从我手里收下这礼物；因为我见了你的面，如同见了上帝的面，并且你也宽容了我。
GEN|33|11|请你收下我带来给你的礼物，因为上帝恩待我，使我一切都充足。” 雅各 再三求他，他才收下。
GEN|33|12|以扫 说：“让我们起身前行，我和你一起走吧。”
GEN|33|13|雅各 对他说：“我主知道孩子们还年幼娇嫩，我的牛羊也正在哺乳中，只要催赶一天，群羊都会死了。
GEN|33|14|请我主在仆人前面先走，我要按着在我面前的牲畜和孩子的步伐慢慢前进，直走到 西珥 我主那里。”
GEN|33|15|以扫 说：“让我把跟随我的人留几个在你这里。” 雅各 说：“何必这样呢？只要能在我主眼前蒙恩就够了。”
GEN|33|16|于是， 以扫 当日起行，回 西珥 去了。
GEN|33|17|雅各 就往 疏割 去，在那里为自己盖房屋，又为牲畜搭棚，因此那地方叫 疏割 。
GEN|33|18|雅各 从 巴旦．亚兰 平安地回到 迦南 地的 示剑城 ，他在城的前面支搭帐棚。
GEN|33|19|他用一百可锡塔 从 示剑 的父亲 哈抹 的众子手中买了搭帐棚的那块地。
GEN|33|20|雅各 在那里筑了一座坛，起名叫 伊利．伊罗伊．以色列 。
GEN|34|1|利亚 给 雅各 所生的女儿 底拿 出去，要探望那地的女子们。
GEN|34|2|那地的族长 希未 人 哈抹 的儿子 示剑 看见她，就拉住她，与她同寝，玷辱了她。
GEN|34|3|示剑 的心喜欢 雅各 的女儿 底拿 ，爱上这少女，甜言蜜语地安慰她。
GEN|34|4|示剑 对他父亲 哈抹 说：“求你为我聘这女孩为妻。”
GEN|34|5|雅各 听见 示剑 污辱了他的女儿 底拿 。那时他的儿子们正和牲畜在田野， 雅各 就沉默，等他们回来。
GEN|34|6|示剑 的父亲 哈抹 出来，到 雅各 那里，要和他讲话。
GEN|34|7|雅各 的儿子们听见这事，就从田野回来，人人悲愤，十分恼怒，因 示剑 在 以色列 中做了丑事，与 雅各 的女儿同寝，这本是不该做的事。
GEN|34|8|哈抹 和他们谈话，说：“我儿子 示剑 的心喜欢你们家的女儿，请你们把她嫁给我的儿子。
GEN|34|9|你们与我们彼此结亲；你们可以把你们家的女儿嫁给我们，也可以娶我们家的女儿。
GEN|34|10|你们与我们同住吧！这地都在你们面前，只管在这里居住，做买卖，置产业。”
GEN|34|11|示剑 对女子的父亲和兄弟们说：“愿你们看得起我，你们向我要什么，我必给你们，
GEN|34|12|无论向我要多贵重的聘金和礼物，我必照你们所说的给你们，只要你们将这少女嫁给我。”
GEN|34|13|雅各 的儿子们因 示剑 污辱了他们的妹妹 底拿 ，就用诡诈的话回答 示剑 和他父亲 哈抹 ，
GEN|34|14|对他们说：“我们不能做这样的事，把我们的妹妹嫁给没有受割礼的人为妻，因为那是我们的羞耻。
GEN|34|15|惟有一个条件，我们才答应你们，就是你们所有的男丁都要受割礼，和我们一样，
GEN|34|16|我们就把我们家的女儿嫁给你们，也娶你们家的女儿；我们就与你们同住，大家成为一族人。
GEN|34|17|倘若你们不听从我们受割礼，我们就带我们家的女儿走了。”
GEN|34|18|这些话在 哈抹 和他儿子 示剑 的眼中看为美。
GEN|34|19|那年轻人毫不迟延做这事，因为他爱上了 雅各 的女儿；他在他父亲家中也是最受人尊重的。
GEN|34|20|哈抹 和他儿子 示剑 到他们的城门口，对城里的人讲说：
GEN|34|21|“这些人对我们友善，不如允许他们在这地居住，做买卖；看哪，这地宽阔，足以容纳他们。我们可以娶他们家的女儿，也可以把我们家的女儿嫁给他们。
GEN|34|22|惟有一个条件，这些人才答应和我们同住，成为一族人，就是我们中间所有的男丁都要受割礼，和他们一样。
GEN|34|23|他们的牲畜、财物和一切的牲口岂不都归给我们吗？只要答应他们，他们就与我们同住。”
GEN|34|24|凡从城门出入的人都听从了 哈抹 和他儿子 示剑 的话。于是，凡从城门出入的男丁都受了割礼。
GEN|34|25|到第三天，他们正疼痛的时候， 雅各 的两个儿子，就是 底拿 的哥哥 西缅 和 利未 ，各拿刀剑，不动声色地来到城中，把所有的男丁都杀了，
GEN|34|26|又用刀杀了 哈抹 和他儿子 示剑 ，把 底拿 从 示剑 家里带走，就离开了。
GEN|34|27|雅各 的儿子们因为他们的妹妹受污辱，就来到被杀的人那里，洗劫那城，
GEN|34|28|夺走了他们的羊群、牛群和驴，以及城里和田间所有的；
GEN|34|29|又俘掳抢劫他们一切的财物、孩童、妇女，以及房屋中所有的。
GEN|34|30|雅各 对 西缅 和 利未 说：“你们连累了我，使我在这地的居民中，就是在 迦南 人和 比利洗 人中坏了名声。我的人丁稀少，他们必聚集来击杀我，我和全家的人都要被灭绝。”
GEN|34|31|他们却说：“他岂可待我们的妹妹如同妓女呢？”
GEN|35|1|上帝对 雅各 说：“起来！上 伯特利 去，住在那里。在那里筑一座坛给上帝，就是你逃避你哥哥 以扫 的时候向你显现的上帝。”
GEN|35|2|雅各 就对他家中的人，以及所有和他一起的人说：“除掉你们中间外邦的神明，要自洁，更换衣服。
GEN|35|3|我们要起来，上 伯特利 去，在那里我要筑一座坛给上帝，就是在我遭难的日子应允我，在我行走的路上与我同在的上帝。”
GEN|35|4|他们就把手中所有外邦的神明和自己耳朵上的环子交给 雅各 ； 雅各 把它们埋在 示剑 那里的橡树下。
GEN|35|5|他们起行。上帝使周围城镇的人都惊恐，就不追赶 雅各 的儿子们了。
GEN|35|6|于是 雅各 和所有与他一起的人到了 迦南 地的 路斯 ，就是 伯特利 。
GEN|35|7|他在那里筑了一座坛，给那地方起名叫 伊勒．伯特利 ，因为他逃避他哥哥的时候，上帝曾在那里向他显现。
GEN|35|8|利百加 的奶妈 底波拉 死了，葬在 伯特利 下边的橡树下；那棵树名叫 亚伦．巴古 。
GEN|35|9|雅各 从 巴旦．亚兰 回来，上帝又向他显现，赐福给他。
GEN|35|10|上帝对他说：“你的名原是 雅各 ，从今以后不要再叫 雅各 ，你的名要叫 以色列 。”于是，上帝就叫他的名为 以色列 。
GEN|35|11|上帝又对他说：“我是全能的上帝；你要生养众多，将来有一国和许多的国从你而来，又有许多君王从你生出 。
GEN|35|12|至于我赐给 亚伯拉罕 和 以撒 的地，我必赐给你；我必赐这地给你的后裔。”
GEN|35|13|上帝就从与 雅各 说话的那地方升上去了。
GEN|35|14|雅各 就在上帝与他说话的地方立了一根柱子，就是石柱，在它上面献浇酒祭，又浇油。
GEN|35|15|雅各 就给上帝与他说话的那地方起名叫 伯特利 。
GEN|35|16|他们从 伯特利 起行，到 以法他 还有一段路程， 拉结 生产，生得十分艰难。
GEN|35|17|她生得十分艰难的时候，接生婆对她说：“不要怕，你又要有一个儿子了。”
GEN|35|18|她快要死，还有一口气的时候，就给她儿子起名叫 便．俄尼 ；他父亲却给他起名叫 便雅悯 。
GEN|35|19|拉结 死了，葬在往 以法他 的路旁； 以法他 就是 伯利恒 。
GEN|35|20|雅各 在她的坟上立了一块碑，就是 拉结 的墓碑，到今日还在。
GEN|35|21|以色列 起行，在 以得台 的那一边支搭帐棚。
GEN|35|22|以色列 住在那地的时候， 吕便 去与他父亲的妾 辟拉 同寝， 以色列 也听见了这件事 。 雅各 共有十二个儿子。
GEN|35|23|利亚 的儿子是 雅各 的长子 吕便 ，还有 西缅 、 利未 、 犹大 、 以萨迦 、 西布伦 。
GEN|35|24|拉结 的儿子是 约瑟 、 便雅悯 。
GEN|35|25|拉结 的婢女 辟拉 的儿子是 但 、 拿弗他利 。
GEN|35|26|利亚 的婢女 悉帕 的儿子是 迦得 、 亚设 。这是 雅各 在 巴旦．亚兰 所生的儿子。
GEN|35|27|雅各 来到他父亲 以撒 那里，到了 幔利 ， 基列．亚巴 ，就是 希伯仑 ，是 亚伯拉罕 和 以撒 寄居的地方。
GEN|35|28|以撒 共活了一百八十年。
GEN|35|29|以撒 年纪老迈，安享天年，息劳而终，归到他祖先 那里。他两个儿子 以扫 和 雅各 把他安葬了。
GEN|36|1|这是 以扫 的后代， 以扫 就是 以东 。
GEN|36|2|以扫 娶 迦南 的女子为妻，就是 赫 人 以伦 的女儿 亚大 和 希未 人 祭便 的孙女， 亚拿 的女儿 阿何利巴玛 ，
GEN|36|3|又娶了 以实玛利 的女儿， 尼拜约 的妹妹 巴实抹 。
GEN|36|4|亚大 为 以扫 生了 以利法 ； 巴实抹 生了 流珥 ；
GEN|36|5|阿何利巴玛 生了 耶乌施 、 雅兰 、 可拉 。这些都是 以扫 的儿子，是在 迦南 地生的。
GEN|36|6|以扫 带着他的妻子、儿女和家中所有的人，以及他的牛羊、牲畜和一切财物，就是他在 迦南 地所得的，往别处去，离开了他的兄弟 雅各 。
GEN|36|7|因为他们拥有的很多，不能住在一起。因为牲畜的缘故，寄居的地方容不下他们。
GEN|36|8|于是 以扫 住在 西珥山 ； 以扫 就是 以东 。
GEN|36|9|这是 以扫 的后代，他是 西珥山 里 以东 人的始祖。
GEN|36|10|以扫 子孙的名字如下： 以扫 的妻子 亚大 生 以利法 ； 以扫 的妻子 巴实抹 生 流珥 。
GEN|36|11|以利法 的儿子是 提幔 、 阿抹 、 洗玻 、 迦坦 、 基纳斯 。
GEN|36|12|亭纳 是 以扫 儿子 以利法 的妾，她为 以利法 生了 亚玛力 。这是 以扫 的妻子 亚大 的子孙。
GEN|36|13|流珥 的儿子是 拿哈 、 谢拉 、 沙玛 、 米撒 。这是 以扫 妻子 巴实抹 的子孙。
GEN|36|14|以扫 的妻子 阿何利巴玛 是 祭便 的孙女， 亚拿 的女儿。她为 以扫 生了 耶乌施 、 雅兰 、 可拉 。
GEN|36|15|这是 以扫 子孙中作族长的： 以扫 的长子 以利法 的子孙中，有 提幔 族长、 阿抹 族长、 洗玻 族长、 基纳斯 族长、
GEN|36|16|可拉 族长、 迦坦 族长、 亚玛力 族长。这是在 以东 地，从 以利法 所出的族长，是 亚大 的子孙。
GEN|36|17|以扫 的儿子 流珥 的子孙中，有 拿哈 族长、 谢拉 族长、 沙玛 族长、 米撒 族长。这是在 以东 地，从 流珥 所出的族长，是 以扫 妻子 巴实抹 的子孙。
GEN|36|18|以扫 的妻子 阿何利巴玛 的子孙中，有 耶乌施 族长、 雅兰 族长、 可拉 族长。这是从 以扫 的妻子， 亚拿 的女儿 阿何利巴玛 的子孙中所出的族长。
GEN|36|19|以上的族长都是 以扫 的子孙； 以扫 就是 以东 。
GEN|36|20|这是那地原来的居民， 何利 人 西珥 的子孙： 罗坍 、 朔巴 、 祭便 、 亚拿 、
GEN|36|21|底顺 、 以察 、 底珊 。这是在 以东 地，从 何利 人 西珥 子孙中所出的族长。
GEN|36|22|罗坍 的儿子是 何利 、 希幔 ， 罗坍 的妹妹是 亭纳 。
GEN|36|23|朔巴 的儿子是 亚勒文 、 玛拿辖 、 以巴录 、 示玻 、 阿南 。
GEN|36|24|祭便 的儿子是 爱亚 、 亚拿 ，当时在旷野牧放他父亲 祭便 的驴，发现温泉的就是这 亚拿 。
GEN|36|25|亚拿 的儿子是 底顺 ， 亚拿 的女儿是 阿何利巴玛 。
GEN|36|26|底顺 的儿子是 欣但 、 伊是班 、 益兰 、 基兰 。
GEN|36|27|以察 的儿子是 辟罕 、 撒番 、 亚干 。
GEN|36|28|底珊 的儿子是 乌斯 、 亚兰 。
GEN|36|29|这是从 何利 人所出的族长： 罗坍 族长、 朔巴 族长、 祭便 族长、 亚拿 族长、
GEN|36|30|底顺 族长、 以察 族长、 底珊 族长。这是从 何利 人所出的族长，都在 西珥 地，按着族长 来分。
GEN|36|31|以色列 未有君王治理之前，这些是在 以东 地作王的。
GEN|36|32|比珥 的儿子 比拉 在 以东 作王，他的城名叫 亭哈巴 。
GEN|36|33|比拉 死了， 波斯拉 人 谢拉 的儿子 约巴 接续他作王。
GEN|36|34|约巴 死了， 提幔 人之地的 户珊 接续他作王。
GEN|36|35|户珊 死了， 比达 的儿子 哈达 接续他作王， 哈达 曾在 摩押 地击败 米甸 人，他的城名叫 亚未得 。
GEN|36|36|哈达 死了， 玛士利加 人 桑拉 接续他作王。
GEN|36|37|桑拉 死了， 大河 边的 利河伯 人 扫罗 接续他作王。
GEN|36|38|扫罗 死了， 亚革波 的儿子 巴勒．哈南 接续他作王。
GEN|36|39|亚革波 的儿子 巴勒．哈南 死了， 哈达尔 接续他作王，他的城名叫 巴乌 。他的妻子名叫 米希她别 ，是 米．萨合 的孙女， 玛特列 的女儿。
GEN|36|40|这些是 以扫 的族长，按着他们的宗族、住处和名字： 亭纳 族长、 亚勒瓦 族长、 耶帖 族长、
GEN|36|41|阿何利巴玛 族长、 以拉 族长、 比嫩 族长、
GEN|36|42|基纳斯 族长、 提幔 族长、 米比萨 族长、
GEN|36|43|玛基叠 族长、 以兰 族长。这些是 以东 人在所得为业的地上，按着他们住处的族长。 以扫 是 以东 人的始祖。
GEN|37|1|雅各 住在 迦南 地，就是他父亲寄居的地。
GEN|37|2|这是 雅各 的事迹。 约瑟 十七岁与他哥哥们一同牧羊。他是个少年，与他父亲的妾 辟拉 和 悉帕 的儿子们常在一起。 约瑟 把他们的恶行报给父亲。
GEN|37|3|以色列 爱 约瑟 过于其他的儿子，因为 约瑟 是他年老生的；他给 约瑟 做了一件长袍 。
GEN|37|4|哥哥们见父亲爱 约瑟 过于他们，就恨 约瑟 ，不与他说友善的话。
GEN|37|5|约瑟 做了一个梦，告诉他哥哥们，他们就更加恨他。
GEN|37|6|约瑟 对他们说：“请听我做的这个梦：
GEN|37|7|看哪，我们在田里捆禾稼；看哪，我的捆起来站着；看哪，你们的捆围着我的捆下拜。”
GEN|37|8|他的哥哥们对他说：“难道你真的要作我们的王吗？难道你真的要统治我们吗？”他们就因他的梦和他的话更加恨他。
GEN|37|9|后来他又做了另一个梦，告诉他哥哥们说：“看哪，我又做了一个梦；看哪，太阳、月亮和十一颗星都向我下拜。”
GEN|37|10|约瑟 告诉他父亲和哥哥们，他父亲就责备他说：“你做的这是什么梦！难道我和你母亲、你的兄弟真的要俯伏在地，来向你下拜吗？”
GEN|37|11|他的哥哥们都嫉妒他，他父亲却把这事存在心里。
GEN|37|12|约瑟 的哥哥们到 示剑 去放他们父亲的羊。
GEN|37|13|以色列 对 约瑟 说：“你哥哥们不是在 示剑 放羊吗？来，我派你到他们那里去。” 约瑟 对他说：“我在这里。”
GEN|37|14|以色列 对他说：“你去看看你哥哥们是否平安，羊群是否平安，再回来告诉我。”于是他派 约瑟 出 希伯仑谷 ， 约瑟 就往 示剑 去了。
GEN|37|15|有人遇见他，看哪，他在田野走迷了路。那人问他说：“你找什么？”
GEN|37|16|他说：“我找我的哥哥们，请告诉我，他们在哪里放羊。”
GEN|37|17|那人说：“他们已经离开这里走了，我听见他们说：‘我们往 多坍 去。’” 约瑟 就去追哥哥们，在 多坍 找到了他们。
GEN|37|18|他们远远看见他，趁他还没有走近他们，就图谋要杀死他。
GEN|37|19|他们彼此说：“看哪！那做梦的来了。
GEN|37|20|现在，来吧！我们把他杀了，丢在一个坑里，就说有恶兽把他吃了。我们且看他的梦将来怎么样。”
GEN|37|21|吕便 听见了，要救 约瑟 脱离他们的手，说：“我们不可害他的性命”；
GEN|37|22|吕便 又对他们说：“不可流他的血，可以把他丢在这旷野的坑里，不可下手害他。” 吕便 要救他脱离他们的手，把他还给他父亲。
GEN|37|23|约瑟 到了他哥哥们那里，他们就剥去他的外衣，就是他身上那件长袍。
GEN|37|24|他们抓住他，把他丢在坑里。那坑是空的，里头没有水。
GEN|37|25|他们坐下吃饭，举目观看，看哪，有一群 以实玛利 人从 基列 来，用骆驼驮着香料、乳香、没药，要带下 埃及 去。
GEN|37|26|犹大 对他的兄弟们说：“我们杀我们的弟弟，遮掩他的血有什么好处呢？
GEN|37|27|来，我们把他卖给 以实玛利 人，不要下手害他，因为他是我们的弟弟，我们的骨肉。”他的兄弟们就听从了他。
GEN|37|28|那时，有些 米甸 的商人从那里经过，就把 约瑟 从坑里拉上来。他们以二十块银子把 约瑟 卖给 以实玛利 人，他们就把 约瑟 带到 埃及 去了。
GEN|37|29|吕便 回到坑旁，看哪， 约瑟 不在坑里，就撕裂自己的衣服，
GEN|37|30|回到他兄弟们那里，说：“孩子不在了。我往哪里去才好呢？”
GEN|37|31|于是，他们宰了一只公山羊，拿了 约瑟 的那件外衣染上了血，
GEN|37|32|派人把长袍送到他们的父亲那里，说：“我们发现这个， 请认一认，是不是你儿子的外衣？”
GEN|37|33|他认出来，就说：“这是我儿子的外衣，恶兽把他吃了， 约瑟 一定被撕碎了！”
GEN|37|34|雅各 就撕裂衣服，腰间围上麻布，为他儿子哀伤了多日。
GEN|37|35|他的儿女都起来安慰他，他却不肯受安慰，说：“我必哀伤着下阴间，到我儿子那里。” 约瑟 的父亲就为他哀哭。
GEN|37|36|米甸 人把 约瑟 卖到 埃及 ，给法老的官员，就是护卫长 波提乏 。
GEN|38|1|那时， 犹大 离开他兄弟们下去，到一个名叫 希拉 的 亚杜兰 人的家附近支搭帐棚。
GEN|38|2|犹大 在那里看见一个名叫 拔．书亚 的 迦南 女子，就娶她为妻，与她同房，
GEN|38|3|她就怀孕生了儿子， 犹大 给他起名叫 珥 。
GEN|38|4|她又怀孕生了儿子，给他起名叫 俄南 。
GEN|38|5|她又再生了儿子，给他起名叫 示拉 。她生 示拉 的时候， 犹大 正在 基悉 。
GEN|38|6|犹大 为长子 珥 娶妻，名叫 她玛 。
GEN|38|7|犹大 的长子 珥 在耶和华眼中看为恶，耶和华就杀死了他。
GEN|38|8|犹大 对 俄南 说：“你当与你哥哥的妻子同房，向她尽你的本分，为你哥哥生子立后。”
GEN|38|9|俄南 知道如果与嫂嫂同房，所生的孩子不属于自己，就泄在地上，不为哥哥生子立后。
GEN|38|10|俄南 所做的在耶和华眼中看为恶，耶和华也杀死了他。
GEN|38|11|犹大 对他媳妇 她玛 说：“你去住在你父亲家里守寡，等我儿子 示拉 长大。”因为他说：“恐怕 示拉 也像两个哥哥一样死去。” 她玛 就去，住在她父亲家里。
GEN|38|12|过了一段很长的日子， 犹大 的妻子， 书亚 的女儿死了。 犹大 受到了安慰，就和他朋友 亚杜兰 人 希拉 上 亭拿 去，到他的剪羊毛的人那里。
GEN|38|13|有人告诉 她玛 说：“看哪，你的公公上 亭拿 剪羊毛去了。”
GEN|38|14|她玛 见 示拉 已经长大，却还没有娶她为妻，就脱去她寡妇的衣裳，用面纱蒙着，盖住自己，坐在往 亭拿 的路上， 伊拿印 城门口。
GEN|38|15|犹大 看见她，以为是妓女，因为她蒙着脸。
GEN|38|16|犹大 就转到路边她那里，说：“来吧！让我与你同寝。”他并不知道她就是他的媳妇。 她玛 说：“你要与我同寝，把什么给我呢？”
GEN|38|17|犹大 说：“我从羊群里取一只小山羊，派人送来给你。” 她玛 说：“在未送之前，你能给我一个信物吗？”
GEN|38|18|他说：“我给你什么信物呢？” 她玛 说：“你的印、你的带子 和你手里的杖。”于是 犹大 给了她，与她同寝，她就从 犹大 怀了孕。
GEN|38|19|她玛 起来走了，除去面纱，照常穿上寡妇的衣裳。
GEN|38|20|犹大 托他朋友 亚杜兰 人送一只小山羊去，要从那女人手里取回信物，却找不到她。
GEN|38|21|他问那地方的人说：“ 伊拿印 路旁的神庙娼妓在哪里？”他们说：“这里没有神庙娼妓。”
GEN|38|22|他回到 犹大 那里说：“我找不到她，并且那地方的人说：‘这里没有神庙娼妓。’”
GEN|38|23|犹大 说：“让她拿去吧，免得我们被人讥笑。看哪，我把这小山羊送去了，可是你找不到她。”
GEN|38|24|大约过了三个月，有人告诉 犹大 说：“你的媳妇 她玛 行淫，并且，看哪，她因行淫而怀了孕。” 犹大 说：“拉她出来，把她烧了！”
GEN|38|25|她玛 被拉出来的时候，就派人到她公公那里，对他说：“这些东西是谁的，我就是从谁怀了孕。”她又说：“请你认一认，这印、这带子和这杖是谁的？”
GEN|38|26|犹大 承认说：“她比我更有理，因为我没有把她给我的儿子 示拉 。” 犹大 再也不跟她同寝。
GEN|38|27|她玛 生产的时候到了，看哪，腹里怀的是双胞胎。
GEN|38|28|生产的时候，一个孩子伸出手来；接生婆拿红线绑在他手上，说：“这是头生的。”
GEN|38|29|这孩子把手收回去，看哪，他哥哥生出来了；接生婆说：“你竟然为自己冲出一个裂缝！”于是，他的名字叫 法勒斯 。
GEN|38|30|后来，那手上有红线的兄弟也生出来，他的名字叫 谢拉 。
GEN|39|1|约瑟 被带下 埃及 去。有一个 埃及 人 波提乏 ，是法老的官员，是护卫长，他从那些带 约瑟 下来的 以实玛利 人手中把 约瑟 买了去。
GEN|39|2|约瑟 在他 埃及 主人的家中，耶和华与他同在，他是一个通达的人。
GEN|39|3|他主人见耶和华与他同在，又见耶和华使他手里所办的事都顺利，
GEN|39|4|约瑟 就在主人眼前蒙恩，伺候他主人，主人派他管理家务，把一切所有的都交在他手里。
GEN|39|5|自从主人派 约瑟 管理家务和他一切所有的，耶和华就因 约瑟 的缘故赐福给那 埃及 人的家；凡家里和田间一切所有的，都蒙耶和华赐福。
GEN|39|6|波提乏 把他一切所有的都交在 约瑟 手中，除了自己所吃的食物，其他的事一概不知。 约瑟 英俊健美。
GEN|39|7|这些事以后， 约瑟 主人的妻子以目送情给 约瑟 ，说：“你与我同寝吧！”
GEN|39|8|约瑟 拒绝，对他主人的妻子说：“看哪，一切家务我主人一概不知，他把所有的都交在我手里。
GEN|39|9|在这家里没有人比我更大，除你以外，他也没有留下一样不交给我，因为你是他的妻子。我怎能行这么大的恶，得罪上帝呢？”
GEN|39|10|她天天这样对 约瑟 说， 约瑟 却不听从她，不与她同寝，也不和她在一起。
GEN|39|11|有一天， 约瑟 进屋里去办事，家里没有一个人在那屋子里，
GEN|39|12|妇人就拉住他的衣服，说：“你与我同寝吧！” 约瑟 把衣服留在她手里，逃出外面去了。
GEN|39|13|妇人看见 约瑟 把衣服留在她手里逃到外面，
GEN|39|14|就叫了家里的人来，对他们说：“看，他带了一个 希伯来 人到我们这里戏弄我们。他到我这里来，要与我同寝，我就大声喊叫。
GEN|39|15|他听见我放声大喊，就把他的衣服留在我这里，逃出外面去了。”
GEN|39|16|妇人把 约瑟 的衣服放在身边，直到他主人回家，
GEN|39|17|就用这样的话对他说：“你带到我们这里来的那 希伯来 仆人进来要调戏我，
GEN|39|18|我放声大喊，他就把衣服留在我身边，逃到外面。”
GEN|39|19|主人听见他妻子对他说的话，说：“你的仆人就是这样对待我”，就非常生气。
GEN|39|20|约瑟 的主人把他抓起来，关在监狱里，就是王的囚犯被关的地方。于是 约瑟 在那里坐牢。
GEN|39|21|但耶和华与 约瑟 同在，向他施恩，使他在监狱长的眼前蒙恩。
GEN|39|22|监狱长就把监狱里所有的囚犯都交在 约瑟 手下；在那里的一切事都由他处理。
GEN|39|23|任何交在 约瑟 手中的事，监狱长一概不察，因为耶和华与 约瑟 同在，耶和华使他所做的都顺利。
GEN|40|1|这些事以后， 埃及 王的司酒长和司膳长得罪了他们的主 埃及 王。
GEN|40|2|法老就对司酒长和司膳长两个官员发怒，
GEN|40|3|把他们关在护卫长府内的监狱里，就是 约瑟 被囚的地方。
GEN|40|4|护卫长把他们交给 约瑟 ， 约瑟 就伺候他们。他们被关了一段日子。
GEN|40|5|关在监狱里的这两个人，就是 埃及 王的司酒长和司膳长，在同一个晚上各自做了一个梦，每个梦都有自己的解释。
GEN|40|6|到了早晨， 约瑟 来到他们那里看他们，看哪，他们很忧愁。
GEN|40|7|他就问一同关在他主人府内法老的官员，说：“你们今日为什么面带愁容呢？”
GEN|40|8|他们对他说：“我们各自做了一个梦，却没有人能讲解。” 约瑟 对他们说：“解梦不是出于上帝吗？请你们把梦告诉我。”
GEN|40|9|司酒长就把梦告诉 约瑟 ，对他说：“在我的梦中，看哪，有一棵葡萄树在我面前，
GEN|40|10|树上有三根枝子。枝子发了芽，开了花，结出串串成熟的葡萄。
GEN|40|11|法老的杯在我手中，我就拿葡萄挤在法老的杯里，把杯递到他手中。”
GEN|40|12|约瑟 对他说：“梦的解释是这样：三根枝子就是三天；
GEN|40|13|三天之内，法老要让你抬起头来，叫你官复原职。你仍要递杯在法老的手中，像先前作他的司酒长一样。
GEN|40|14|但你得福的时候，请你记得我，向我施慈爱，在法老面前提起我，救我出这监牢。
GEN|40|15|我实在是从 希伯来 人之地被拐来的，我在这里也没有做过什么，好叫他们把我关在牢里。”
GEN|40|16|司膳长见梦解得好，就对 约瑟 说：“在我梦中，看哪，我头上顶着三个装饼的篮子；
GEN|40|17|最上面的篮子里有为法老烤的各样食物，有飞鸟来吃我头上篮子里的食物。”
GEN|40|18|约瑟 说：“梦的解释是这样：三个篮子就是三天；
GEN|40|19|三天之内，法老要让你抬起头来，身首异处，把你挂在木架上，必有飞鸟来吃你身上的肉。”
GEN|40|20|到了第三天，正是法老的生日，他为众臣仆摆设宴席，使司酒长和司膳长从众臣仆中抬起头来，
GEN|40|21|让司酒长官复原职，仍旧递杯在法老手中，
GEN|40|22|却把司膳长挂起来，正如 约瑟 向他们所讲解的。
GEN|40|23|然而，司酒长不记得 约瑟 ，竟忘了他。
GEN|41|1|过了两年，法老做梦，看哪，自己站在 尼罗河 边，
GEN|41|2|看哪，有七头母牛从 尼罗河 里上来，长相俊美，肌肉肥壮，在芦苇中吃草。
GEN|41|3|看哪，随后又有七头母牛从 尼罗河 里上来，长相丑陋，肌肉干瘦，与那七头母牛一同站在河边。
GEN|41|4|这长相丑陋，肌肉干瘦的七头母牛吃了那长相俊美又肥壮的七头母牛。法老就醒了。
GEN|41|5|他又睡着，第二次做梦，看哪，一株麦杆长了七个穗子，又肥大又佳美，
GEN|41|6|看哪，随后又长出七个穗子，又细弱又被东风吹焦了。
GEN|41|7|这细弱的穗子吞了那七个又肥大又饱满的穗子。法老醒了，看哪，是个梦。
GEN|41|8|到了早晨，法老心里不安，就派人把 埃及 所有的术士和智慧人都召来。法老把所做的梦告诉他们，但是没有人能为法老解梦。
GEN|41|9|那时司酒长对法老说：“我今日想起我的罪来。
GEN|41|10|从前法老对臣仆发怒，把我和司膳长关在护卫长府内的监牢里。
GEN|41|11|我们两人在同一晚上各做一梦，每个梦都有各自的解释。
GEN|41|12|同我们在一起有一个 希伯来 的年轻人，是护卫长的仆人。我们告诉他，他就为我们解梦，照着各人的梦讲解。
GEN|41|13|后来事情正如他给我们讲解的实现了，我官复原职，司膳长被挂起来了。”
GEN|41|14|于是法老派人去召 约瑟 ，他们就急忙把他从牢里提出来。他就剃头刮脸，换衣服，进到法老面前。
GEN|41|15|法老对 约瑟 说：“我做了一个梦，没有人能讲解。我听人说，你听了梦就能讲解。”
GEN|41|16|约瑟 回答法老说：“这不在乎我。上帝必应允法老平安。”
GEN|41|17|法老对 约瑟 说：“在我的梦中，看哪，我站在 尼罗河 边，
GEN|41|18|看哪，有七头母牛从 尼罗河 里上来，肌肉肥壮，外形俊美，在芦苇中吃草。
GEN|41|19|看哪，随后又有七头母牛上来，虚弱，外形很丑陋，肌肉又干瘦，在 埃及 全地，我没有见过这样丑陋的牛。
GEN|41|20|这干瘦又丑陋的母牛吃了那先前的七头肥母牛，
GEN|41|21|进了肚子以后却看不出已经进了肚子，那丑陋的长相仍旧和先前一样。我就醒了。
GEN|41|22|我又在梦中观看，看哪，一株麦杆长了七个穗子，又饱满又佳美，
GEN|41|23|看哪，随后又长出七个穗子，枯槁，细弱，又被东风吹焦了。
GEN|41|24|这些细弱的穗子吞了那七个佳美的穗子。我告诉术士，却没有人能为我讲解。”
GEN|41|25|约瑟 对法老说：“法老的梦是同一个。上帝已把要做的事指示法老了。
GEN|41|26|七头好母牛是七年，七个佳美的穗子也是七年，这是同一个梦。
GEN|41|27|那随后上来的七头干瘦又丑陋的母牛是七年；那七个空心，被东风吹焦的穗子也一样，都是七个荒年。
GEN|41|28|这就是我对法老所说，上帝已把要做的事显明给法老了。
GEN|41|29|看哪，必有七个大丰年来到 埃及 全地，
GEN|41|30|随后又有七个荒年，甚至 埃及 地的人都忘了先前的丰收，这地必被饥荒所灭。
GEN|41|31|因为那后来的饥荒非常严重，就不觉得这地先前有丰收。
GEN|41|32|至于法老两次做梦，是因为上帝已经确定这事，上帝必速速成就。
GEN|41|33|现在，请法老选一个聪明又有智慧的人，委派他治理 埃及 地。
GEN|41|34|请法老这样做，委派官员治理这地，在七个丰年的期间，征收 埃及 地出产的五分之一，
GEN|41|35|叫他们聚集未来丰年一切的粮食，积存五谷归在法老的手下作粮食，储藏在各城里。
GEN|41|36|这粮食可以为这地作储备，为了 埃及 地要来的七个荒年，免得这地被饥荒所灭。”
GEN|41|37|这事在法老和他众臣仆眼中都觉得好。
GEN|41|38|法老对臣仆说：“像这样的人，有上帝的灵在他里面，我们岂能找得着呢？”
GEN|41|39|法老对 约瑟 说：“上帝既指示你这一切事，就没有人像你这样聪明又有智慧。
GEN|41|40|你可以治理我的家；我的百姓都必服从你口中的命令。惟独在宝座上，我比你大。”
GEN|41|41|法老又对 约瑟 说：“看，我委派你治理 埃及 全地。”
GEN|41|42|法老就脱下手上带印的戒指，戴在 约瑟 的手上，给他穿上细麻衣，把金链戴在他的颈项上，
GEN|41|43|又给 约瑟 坐他的副座车，在他前面有人呼叫说：“跪下 。”于是，法老委派他治理 埃及 全地。
GEN|41|44|法老对 约瑟 说：“我是法老，若没有你的命令， 埃及 全地的人都不可擅自办事 。”
GEN|41|45|法老给 约瑟 起名叫 撒发那特．巴内亚 ，又将 安城 的祭司 波提．非拉 的女儿 亚西纳 给他为妻。 约瑟 就出去治理 埃及 地。
GEN|41|46|约瑟 在 埃及 王法老面前侍立的时候年三十岁。 约瑟 从法老面前出去，巡行 埃及 全地。
GEN|41|47|七个丰年之内，地的出产极其丰盛 ，
GEN|41|48|约瑟 聚集 埃及 地七年一切的粮食，把粮食积存在各城里，就是把各城周围田地的粮食都积存在该城里。
GEN|41|49|约瑟 积存的五谷很多，如同海边的沙，无法计算，数也数不清。
GEN|41|50|荒年未到以前， 安城 的祭司 波提．非拉 的女儿 亚西纳 为 约瑟 生了两个儿子。
GEN|41|51|约瑟 给长子起名叫 玛拿西 ，因为他说：“上帝使我忘了一切的困苦和我父的全家。”
GEN|41|52|他给次子起名叫 以法莲 ，因为他说：“上帝使我在受苦的地方兴盛。”
GEN|41|53|埃及 地的七个丰年一过，
GEN|41|54|七个荒年就来了，正如 约瑟 所说的。各地都有饥荒，惟独 埃及 全地有粮食。
GEN|41|55|等到 埃及 全地也有了饥荒，众百姓就向法老哀求粮食。法老对所有的 埃及 人说：“你们到 约瑟 那里去，凡他所说的，你们都要做。”
GEN|41|56|当时饥荒遍满了全地， 约瑟 就开了各处的粮仓 ，卖粮食给 埃及 人。 埃及 地的饥荒非常严重。
GEN|41|57|各地的人都去 埃及 ，到 约瑟 那里买粮食，因为全地的饥荒非常严重。
GEN|42|1|雅各 见 埃及 有粮，就对儿子们说：“你们为什么彼此对看呢？”
GEN|42|2|他又说：“看哪，我听见 埃及 有粮，你们可以下到那里，从那里为我们买些粮来，我们就可以存活，不至于死。”
GEN|42|3|于是， 约瑟 的十个哥哥都下去，到 埃及 买粮食。
GEN|42|4|至于 约瑟 的弟弟 便雅悯 ， 雅各 没有派他和哥哥们同去，因为 雅各 说：“恐怕他遭难。”
GEN|42|5|以色列 的儿子们来了，在前来的人当中，为要买粮食，因为 迦南 地也有饥荒。
GEN|42|6|当时在 埃及 地掌权的人是 约瑟 ，卖粮给各地众百姓的就是他。 约瑟 的哥哥们来了，脸伏于地，向他下拜。
GEN|42|7|约瑟 看见他哥哥们，就认出他们，却对他们装作陌生人，向他们说严厉的话，对他们说：“你们从哪里来？”他们说：“我们从 迦南 地来买粮。”
GEN|42|8|约瑟 认得他哥哥们，他们却不认得他。
GEN|42|9|约瑟 想起从前所做的那两个梦，就对他们说：“你们是奸细，你们来是要窥探这地的虚实。”
GEN|42|10|他们对他说：“我主啊，不是的，仆人们是来买粮的。
GEN|42|11|我们都是同一个人的儿子，我们是诚实的人。仆人们并不是奸细。”
GEN|42|12|约瑟 对他们说：“不，你们一定是窥探这地的虚实来的。”
GEN|42|13|他们说：“仆人们本是兄弟十二人，我们都是 迦南 地同一个人的儿子。看哪，最小的今日在我们父亲那里，有一个不在了。”
GEN|42|14|约瑟 对他们说：“我刚才对你们说过了，你们是奸细！
GEN|42|15|我指着法老的性命起誓，若是你们最小的弟弟不到这里来，你们就不可以离开这里；这样你们就可以证实自己了。
GEN|42|16|要派你们当中的一个人去，把你们的弟弟带来。至于你们，都要关在这里，好证实你们的话是不是真的。若不是，我指着法老的性命起誓，你们一定是奸细。”
GEN|42|17|于是 约瑟 把他们一起都关在监里三天。
GEN|42|18|第三天， 约瑟 对他们说：“我是敬畏上帝的，你们这么做就可以活。
GEN|42|19|如果你们是诚实的人，留你们兄弟中的一个关在监牢里，你们带粮食回去，救你们家的饥荒，
GEN|42|20|再把你们最小的弟弟带到我这里来。如此，你们的话就是真的了，你们也不至于死。”他们就照样做了。
GEN|42|21|他们彼此说：“我们在弟弟身上实在犯了罪。他哀求我们的时候，我们看见他的痛苦，却不肯听，所以这场苦难临到我们。”
GEN|42|22|吕便 回答他们说：“我不是对你们说过，不可伤害那孩子吗？只是你们不肯听，看哪，他的血在追讨了。”
GEN|42|23|他们不知道 约瑟 在听，因为在他们之间有传译官。
GEN|42|24|约瑟 转身离开他们，哭了一场，又回来对他们说话，就从他们中间抓了 西缅 ，在他们眼前捆绑他。
GEN|42|25|约瑟 吩咐人把他们的器皿装满粮食，把各人的银子退还在各人的袋里，又给他们路上需用的食物。人就为他们这样做了。
GEN|42|26|他们把粮食驮在驴上，离开那里去了。
GEN|42|27|到了住宿的地方，有一个人打开袋子，要拿饲料喂驴，就看见自己的银子，看哪，仍在袋口上。
GEN|42|28|他对兄弟们说：“我的银子退回来了，看哪，还在我袋子里！”他们战战兢兢，心都快跳出来了，彼此说：“上帝向我们做的是什么呢？”
GEN|42|29|他们来到 迦南 地他们的父亲 雅各 那里，把所遭遇的事都告诉他，说：
GEN|42|30|“那地的主对我们说严厉的话，把我们当作窥探那地的奸细。
GEN|42|31|我们对他说：‘我们是诚实的人，并不是奸细。
GEN|42|32|我们本是兄弟十二人，都是同一个父亲的儿子，有一个不在了，最小的今日和我们父亲在 迦南 地。’
GEN|42|33|那地的主对我们说：‘只有这样我才知道你们是诚实的人：留你们兄弟中的一个在我这里，你们带粮食回去，救你们家的饥荒，
GEN|42|34|再把你们最小的弟弟带到我这里来，我就知道你们不是奸细，是诚实的人。然后，我就把你们的兄弟交还你们，你们也可以在此地做买卖。’”
GEN|42|35|后来他们倒空袋子，看哪，各人的银囊都在袋子里。他们和父亲看见银囊就都害怕。
GEN|42|36|他们的父亲 雅各 对他们说：“你们害我丧失了我的儿子： 约瑟 不在了， 西缅 也不在了，你们还要带走 便雅悯 ！这些事都临到我身上了。”
GEN|42|37|吕便 对他父亲说：“我若不带他回来给你，你可以杀我的两个儿子。只管把他交在我手里，我必带他回来给你。”
GEN|42|38|雅各 说：“我的儿子不可与你们一同下去。他哥哥死了，只剩下他。他若在你们行走的路上遭难，你们就害我白发苍苍、悲悲惨惨下阴间去了。”
GEN|43|1|那地的饥荒非常严重。
GEN|43|2|他们从 埃及 带来的粮食吃完了，父亲对他们说：“你们再去给我们买些粮来。”
GEN|43|3|犹大 对他说：“那人严厉地警告我们说：‘你们的弟弟若不和你们同来，你们就不要来见我的面。’
GEN|43|4|你若派我们的弟弟跟我们同去，我们就下去给你买粮；
GEN|43|5|你若不派他去，我们就不下去，因为那人对我们说：‘你们的弟弟若不和你们同来，你们就不要来见我的面。’”
GEN|43|6|以色列 说：“你们为什么这样害我，告诉那人你们还有弟弟呢？”
GEN|43|7|他们说：“那人详细问到我们和我们的家人，说：‘你们的父亲还在吗？你们还有兄弟吗？’我们就按着他的这些话告诉他，我们怎么知道他会说：‘把你们的弟弟带下来’呢？”
GEN|43|8|犹大 又对他父亲 以色列 说：“请派这年轻人和我同去，我们就动身前去，好叫我们和你，以及我们的孩子都得存活，不至于死。
GEN|43|9|我为他担保，你可以从我手中要人，我若不带他回来交在你面前，我就对你永远担当这罪。
GEN|43|10|我们若没有耽搁，现在第二趟都回来了。”
GEN|43|11|父亲 以色列 对他们说：“如果必须如此，你们要这样做：把本地土产中最好的乳香、蜂蜜、香料、没药、坚果、杏仁各取一点，放在器皿里，带下去送给那人作礼物。
GEN|43|12|手里要带双倍的银子，把退还在你们袋口的银子亲手带回去；或许那是个失误。
GEN|43|13|带着你们的弟弟，动身再去见那人。
GEN|43|14|愿全能的上帝使你们在那人面前蒙怜悯，放你们另一个兄弟和 便雅悯 回来。我若要失丧儿子，就丧了吧！”
GEN|43|15|于是，他们拿着那些礼物，手里也带双倍的银子，并且带着 便雅悯 ，动身下到 埃及 ，站在 约瑟 面前。
GEN|43|16|约瑟 见 便雅悯 和他们同来，就对管家说：“把这些人领到屋里。要宰杀牲畜，预备宴席，因为中午这些人要跟我吃饭。”
GEN|43|17|那人就照 约瑟 所说的去做，领他们进 约瑟 的屋里。
GEN|43|18|这些人因为被领到 约瑟 的屋里，就害怕，说：“领我们到这里来，必是因为当初退还在我们袋里的银子，要设计害我们，抓我们去当奴隶，抢夺我们的驴。”
GEN|43|19|他们就挨近 约瑟 的管家，在屋子门口和他说话，
GEN|43|20|说：“我主啊，求求你，我们当初下来，真的是要买粮食。
GEN|43|21|后来到了住宿的地方，我们打开袋子，看哪，各人的银子还在自己的袋口上，银子的分量一点不少。现在我们亲手把它带回来，
GEN|43|22|我们手里又带了另外的银子来买粮食。我们不知道是谁把银子放在我们袋里的。”
GEN|43|23|他说：“你们平安！不要害怕，是你们的上帝和你们父亲的上帝把财宝放在你们的袋里。你们的银子，我已经收了。”他就把 西缅 带出来，交给他们。
GEN|43|24|那人领这些人进 约瑟 的屋里，给他们水洗脚，又给他们饲料喂驴。
GEN|43|25|他们预备好礼物，等候 约瑟 中午来，因为他们听说他们要在那里吃饭。
GEN|43|26|约瑟 来到家里，他们就把手中的礼物拿进屋里给他，俯伏在地，向他下拜。
GEN|43|27|约瑟 问他们安，又说：“你们的父亲，就是你们所说的那位老人家平安吗？他还在吗？”
GEN|43|28|他们说：“你仆人，我们的父亲平安，他还在。”于是他们低头下拜。
GEN|43|29|约瑟 举目看见他同母的弟弟 便雅悯 ，就说：“你们向我所说那最小的弟弟就是这位吗？”又说：“我儿啊，愿上帝赐恩给你！”
GEN|43|30|约瑟 爱弟之情激动，就急忙找个地方去哭。他进入自己的房间，哭了一场。
GEN|43|31|他洗了脸出来，勉强忍住，就说：“开饭吧！”
GEN|43|32|他们为 约瑟 单独摆了一席，为那些人又摆了一席，也为和 约瑟 同吃饭的 埃及 人另摆了一席，因为 埃及 人不和 希伯来 人一同吃饭；那是 埃及 人所厌恶的。
GEN|43|33|兄弟们被安排在 约瑟 面前坐席，都按着长幼的次序，这些人彼此感到诧异。
GEN|43|34|约瑟 把他面前的食物分给他们，但 便雅悯 所得的比别人多五倍。他们就喝酒，和 约瑟 一同畅饮。
GEN|44|1|约瑟 吩咐管家说：“按照他们的驴子所能驮的，把这些人的袋子装满粮食，再把各人的银子放在各人的袋口上，
GEN|44|2|我的杯，就是那个银杯，要和买粮的银子一同放在最年轻的那个人的袋口上。”管家就照 约瑟 所说的话去做了。
GEN|44|3|天一亮，这些人和他们的驴子就被送走了。
GEN|44|4|他们出城走了不远， 约瑟 对管家说：“起来，去追那些人，追上了就对他们说：‘你们为什么以恶报善呢？
GEN|44|5|这不是我主人用来饮酒，确实用它来占卜的吗？你们这么做是不对的！’”
GEN|44|6|管家追上他们，把这些话对他们说了。
GEN|44|7|他们对他说：“我主为什么说这样的话呢？你仆人们绝不会做这样的事。
GEN|44|8|看哪，我们从前在袋口上发现的银子，尚且从 迦南 地带来还你，我们又怎么会从你主人家里偷窃金银呢？
GEN|44|9|你仆人中无论在谁那里找到杯子，就叫他死，我们也要作我主的奴隶。”
GEN|44|10|管家说：“现在就照你们的话做吧！在谁那里找到杯子，谁就作我的奴隶，其余的人都没有罪。”
GEN|44|11|于是他们各人急忙把袋子卸在地上，各人打开自己的袋子。
GEN|44|12|管家就搜查，从年长的开始到年幼的为止，那杯竟在 便雅悯 的袋子里找到了。
GEN|44|13|他们就撕裂衣服，各人把驮子抬在驴上，回城去了。
GEN|44|14|犹大 和他兄弟们来到 约瑟 的屋里， 约瑟 还在那里，他们就在他面前俯伏于地。
GEN|44|15|约瑟 对他们说：“你们做的是什么事呢？你们岂不知像我这样的人必懂得占卜吗？”
GEN|44|16|犹大 说：“我们对我主能说什么呢？还有什么话可说呢？我们还能为自己表白吗？上帝已经查出你仆人的罪孽了。看哪，我们与那在他手中找到杯子的人都是我主的奴隶。”
GEN|44|17|约瑟 说：“我绝不能做这样的事！谁的手中找到杯子，谁就作我的奴隶。至于你们，可以平平安安上到你们父亲那里去。”
GEN|44|18|犹大 挨近他，说：“我主啊，求求你，让仆人说一句话给我主听，不要向仆人发烈怒，因为你如同法老一样。
GEN|44|19|我主曾问仆人们说：‘你们有父亲、兄弟没有？’
GEN|44|20|我们对我主说：‘我们有父亲，他已经年老，还有他老年所生的一个小儿子。他哥哥死了，他的母亲只剩下他一个孩子，父亲也疼爱他。’
GEN|44|21|你对仆人说：‘把他带下到我这里来，让我亲眼看看他。’
GEN|44|22|我们对我主说：‘这年轻人不能离开他父亲，若是离开，父亲就会死。’
GEN|44|23|你对仆人说：‘你们最小的弟弟若不和你们一同下来，你们就不要来见我的面。’
GEN|44|24|我们上到你仆人，我们父亲那里，就把我主的话告诉了他。
GEN|44|25|后来，我们的父亲说：‘你们再去给我买些粮来。’
GEN|44|26|我们说：‘我们不能下去。最小的弟弟若和我们同去，我们就可以下去。因为，最小的弟弟若不和我们同去，我们必不能见那人的面。’
GEN|44|27|你仆人，我父亲对我们说：‘你们知道我的妻子给我生了两个儿子。
GEN|44|28|一个离开我走了，我说他必是被野兽撕碎了，直到如今我再没有见过他；
GEN|44|29|现在你们又要把这个从我面前带走。倘若他遭难，那么你们就害我白发苍苍、悲悲惨惨下阴间去了。’
GEN|44|30|如今我回到你仆人，我父亲那里，若没有这年轻人和我们同去，我父亲的命是与这年轻人的命相连的，
GEN|44|31|当我们的父亲看见没有了这年轻人，他就会死。这样，我们就害你仆人，我们的父亲白发苍苍、悲悲惨惨下阴间去了。
GEN|44|32|仆人曾向我父亲为这年轻人担保，说：‘我若不带他回来交给父亲，我就在父亲面前永远担当这罪。’
GEN|44|33|现在，求你把仆人留下，代替这年轻人作我主的奴隶，让这年轻人和他哥哥们一同上去。
GEN|44|34|若这年轻人不和我一起，我怎能上到我父亲那里呢？恐怕我要看到灾祸临到我父亲了。”
GEN|45|1|约瑟 在所有侍立在他旁边的人面前情不自禁，就喊叫说：“每一个人都离开我，出去吧！” 约瑟 和兄弟相认的时候没有一人站在他那里。
GEN|45|2|他放声大哭， 埃及 人听见了，法老家中的人也听见了。
GEN|45|3|约瑟 对他兄弟们说：“我就是 约瑟 。我的父亲还在吗？”他兄弟们不敢回答他，因为他们在他面前都很惊惶。
GEN|45|4|约瑟 又对他兄弟们说：“靠近我一点。”他们就近前来。他说：“我是被你们卖到 埃及 的兄弟 约瑟 。
GEN|45|5|现在，不要因为把我卖到这里而忧伤，对自己生气，因为上帝差我在你们以先来，为要保全性命。
GEN|45|6|现在这地的饥荒已经二年了，还有五年不能耕种，没有收成。
GEN|45|7|上帝差我在你们以先来，为要给你们在世上存留余种，大施拯救，保全你们的性命。
GEN|45|8|这样看来，差我到这里来的不是你们，而是上帝。他又使我如同法老之父，作他全家之主，和 埃及 全地掌权的人。
GEN|45|9|你们要赶紧上到我父亲那里，对他说：‘你儿子 约瑟 这样说：上帝已立我作全 埃及 之主，请你下到我这里来，不要耽搁。
GEN|45|10|你和你的儿子孙子，羊群牛群，以及一切所有的，都可以住在 歌珊 地，与我相近。
GEN|45|11|我要在那里奉养你，因为还有五年的饥荒，免得你和你的家属，以及一切所有的，都陷入穷困中。’
GEN|45|12|看哪，你们的眼睛和我弟弟 便雅悯 的眼睛都看见，是我亲口对你们说话。
GEN|45|13|你们要把我在 埃及 一切的尊荣和你们所有看见的事情都告诉我父亲，也要赶紧请我父亲下到这里来。”
GEN|45|14|于是 约瑟 伏在他弟弟 便雅悯 的颈项上哭， 便雅悯 也在他的颈项上哭。
GEN|45|15|他又亲众兄弟，伏着他们哭。过后，他的兄弟就和他说话。
GEN|45|16|这消息传到法老的宫里，说：“ 约瑟 的兄弟们来了。”法老和他的臣仆眼中都看为好。
GEN|45|17|法老对 约瑟 说：“你要吩咐你的兄弟们说：‘你们要这样做：把驮子抬在牲口上，动身到 迦南 地去，
GEN|45|18|请你们的父亲和你们的家属都到我这里来，我要把 埃及 地的美物赐给你们，你们也要吃这地肥美的出产。’
GEN|45|19|你要吩咐他们：‘要这样做：从 埃及 地带着车辆去，把你们的孩子和妻子，以及你们的父亲都接来。
GEN|45|20|你们的眼不要顾惜你们的家具，因为 埃及 全地的美物都是你们的。’”
GEN|45|21|以色列 的儿子们就照样做了。 约瑟 遵照法老的吩咐，给他们车辆和路上需用的食物。
GEN|45|22|他又给所有哥哥每人一套衣服， 却给 便雅悯 三百银子，五套衣服。
GEN|45|23|他也送给父亲十匹公驴，驮着 埃及 的美物，以及十匹母驴，驮着给他父亲在路上需用的谷物、饼和粮食。
GEN|45|24|于是 约瑟 送他的兄弟们回去，对他们说：“你们不要在路上争吵。”
GEN|45|25|他们从 埃及 上去，来到 迦南 地他们的父亲 雅各 那里，
GEN|45|26|告诉他说：“ 约瑟 还活着，并且作了 埃及 全地掌权的人。” 雅各 心里冰凉，因为不信他们。
GEN|45|27|他们就把 约瑟 对他们所说一切的话都告诉了他。他看见 约瑟 派来接他的车辆，他们父亲 雅各 的灵就苏醒了。
GEN|45|28|以色列 说：“够了！我的儿子 约瑟 还活着，我要趁我未死之前去见他。”
GEN|46|1|以色列 带着一切所有的，起程到 别是巴 去，献祭给他父亲 以撒 的上帝。
GEN|46|2|夜间，上帝在异象中对 以色列 说：“ 雅各 ！ 雅各 ！”他说：“我在这里。”
GEN|46|3|上帝说：“我是上帝，你父亲的上帝。不要害怕下 埃及 去，因为我必使你在那里成为大国。
GEN|46|4|我要和你同下 埃及 去，也必定带你上来； 约瑟 要亲手合上你的眼睛。”
GEN|46|5|雅各 就从 别是巴 起行。 以色列 的儿子让他们的父亲 雅各 和他们的孩子、妻子都坐在法老为 雅各 派来的车上。
GEN|46|6|他们也带着 迦南 地所得的牲畜和财物来到 埃及 。 雅各 和他所有的子孙都一同来了。
GEN|46|7|他把他的儿子、孙子、女儿、孙女，他所有的子孙一同带到 埃及 。
GEN|46|8|这些是来到 埃及 的 以色列 人， 雅各 和他子孙的名字： 雅各 的长子是 吕便 。
GEN|46|9|吕便 的儿子是 哈诺 、 法路 、 希斯伦 、 迦米 。
GEN|46|10|西缅 的儿子是 耶母利 、 雅悯 、 阿辖 、 雅斤 、 琐辖 ，还有 迦南 女子生的儿子 扫罗 。
GEN|46|11|利未 的儿子是 革顺 、 哥辖 、 米拉利 。
GEN|46|12|犹大 的儿子是 珥 、 俄南 、 示拉 、 法勒斯 、 谢拉 ； 珥 与 俄南 死在 迦南 地。 法勒斯 的儿子是 希斯仑 、 哈母勒 。
GEN|46|13|以萨迦 的儿子是 陀拉 、 普瓦 、 约伯 、 伸仑 。
GEN|46|14|西布伦 的儿子是 西烈 、 以伦 、 雅利 。
GEN|46|15|这是 利亚 在 巴旦．亚兰 为 雅各 所生的儿孙，还有女儿 底拿 ，儿孙共三十三人。
GEN|46|16|迦得 的儿子是 洗非芸 、 哈基 、 书尼 、 以斯本 、 以利 、 亚罗底 、 亚列利 。
GEN|46|17|亚设 的儿子是 音拿 、 亦施瓦 、 亦施韦 、 比利亚 ，还有他们的妹妹 西拉 。 比利亚 的儿子是 希别 、 玛结 。
GEN|46|18|这是 拉班 给他女儿 利亚 的婢女 悉帕 的儿孙，她为 雅各 所生的共有十六人。
GEN|46|19|雅各 之妻 拉结 的儿子是 约瑟 和 便雅悯 。
GEN|46|20|约瑟 在 埃及 地生了 玛拿西 和 以法莲 ，是 安城 的祭司 波提非拉 的女儿 亚西纳 为 约瑟 生的。
GEN|46|21|便雅悯 的儿子是 比拉 、 比结 、 亚实别 、 基拉 、 乃幔 、 以希 、 罗实 、 母平 、 户平 、 亚勒 。
GEN|46|22|这是 拉结 为 雅各 所生的儿孙，共有十四人。
GEN|46|23|但 的儿子是 户伸 。
GEN|46|24|拿弗他利 的儿子是 雅薛 、 沽尼 、 耶色 、 示冷 。
GEN|46|25|这是 拉班 给他女儿 拉结 的婢女 辟拉 的儿孙，她为 雅各 所生的共有七人。
GEN|46|26|那与 雅各 同到 埃及 的，除了他媳妇之外，凡从他生的共有六十六人。
GEN|46|27|还有 约瑟 在 埃及 所生的两个儿子。到 埃及 的 雅各 全家共有七十人。
GEN|46|28|雅各 派 犹大 先到 约瑟 那里，请他先指示到 歌珊 去的路；于是他们来到了 歌珊 地。
GEN|46|29|约瑟 备好座车，上 歌珊 去迎接他的父亲 以色列 。他见到父亲，就伏在父亲的颈项上，在父亲的颈项上哭了许久。
GEN|46|30|以色列 对 约瑟 说：“我见了你的面，知道你还活着，现在我可以死了。”
GEN|46|31|约瑟 对他兄弟和他父亲的全家说：“我要上去告诉法老，对他说：‘我在 迦南 地的兄弟和我父亲的全家，都到我这里来了。
GEN|46|32|他们是牧羊人，是牧放牲畜的人；他们把羊群牛群和一切所有的都带来了。’
GEN|46|33|等到法老召见你们，说：‘你们是做什么的？’
GEN|46|34|你们就说：‘你的仆人，从幼年直到现在，都是牧放牲畜的人，我们和我们的祖宗都是这样。’如此，你们就可以住在 歌珊 地，因为凡牧羊的都被 埃及 人厌恶。”
GEN|47|1|约瑟 进去告诉法老说：“我的父亲和我的兄弟带着羊群牛群，以及他们一切所有的，从 迦南 地来了。看哪，他们正在 歌珊 地。”
GEN|47|2|约瑟 从他所有兄弟中挑选五个人，引他们到法老面前。
GEN|47|3|法老对 约瑟 的兄弟说：“你们是做什么的？”他们对法老说：“你仆人是牧羊的，我们和我们的祖宗都是这样。”
GEN|47|4|他们又对法老说：“ 迦南 地的饥荒非常严重，仆人的羊群没有牧草，所以我们来到这地寄居。现在求你准许仆人住在 歌珊 地。”
GEN|47|5|法老对 约瑟 说：“你的父亲和你的兄弟到你这里来了，
GEN|47|6|埃及 地都在你面前，只管让你父亲和你兄弟住在最好的地，他们可以住在 歌珊 地。你若知道他们中间有能干的人，就派他们看管我的牲畜。”
GEN|47|7|约瑟 带他父亲 雅各 来，站在法老面前， 雅各 就为法老祝福。
GEN|47|8|法老对 雅各 说：“你平生的年日是多少呢？”
GEN|47|9|雅各 对法老说：“我在世寄居的年日是一百三十年，我一生的岁月又短又苦，比不上我祖先在世寄居的年日。”
GEN|47|10|雅各 又为法老祝福，就从法老面前退出去了。
GEN|47|11|约瑟 安顿他的父亲和兄弟，遵照法老的命令，把 埃及 境内最好的地，就是 兰塞 地，给他们作为产业。
GEN|47|12|约瑟 用粮食供给他父亲和兄弟们，以及他父亲全家的人，照扶养亲属的人口供给。
GEN|47|13|饥荒非常严重，全地都绝了粮， 埃及 地和 迦南 地都因饥荒耗损了。
GEN|47|14|约瑟 收集了 埃及 地和 迦南 地所有的银子，就是众人买粮的银子， 约瑟 就把那些银子都带到法老的宫里。
GEN|47|15|埃及 地和 迦南 地的银子都花光了， 埃及 众人到 约瑟 那里，说：“我们的银子都用完了，求你给我们粮食吧！我们为什么要死在你面前呢？”
GEN|47|16|约瑟 说：“银子若是用完了，可以把你们的牲畜卖给我，我就以你们的牲畜换粮食给你们。”
GEN|47|17|于是他们把牲畜带到 约瑟 那里， 约瑟 就拿粮食换了他们的马、羊、牛、驴；那一年他因换他们一切的牲畜，用粮食养活他们。
GEN|47|18|那一年过去，第二年他们又来到 约瑟 那里，对他说：“不瞒我主，我们的银子都花光了，牲畜也都归于我主了。我们在我主面前，除了自己的身体和土地以外，一无所剩。
GEN|47|19|你为什么要眼看着我们人死地荒呢？求你用粮食买我们和我们的地，我们和我们的地就要为法老效力。求你给我们种子，使我们可以存活，不致死亡，土地也不致荒芜。”
GEN|47|20|于是， 约瑟 为法老买了 埃及 所有的土地， 埃及 人因饥荒所迫，都卖了自己的田地；那些地都归给法老了。
GEN|47|21|至于百姓，从 埃及 边界的一端到另一端， 约瑟 使他们作奴隶。
GEN|47|22|只有祭司的土地， 约瑟 没有买，因为祭司从法老领取薪俸，靠法老的薪俸过活，所以没有卖自己的土地。
GEN|47|23|约瑟 对百姓说：“看哪，我今日为法老买了你们和你们的土地。看，这些种子是给你们的，你们可以耕种土地。
GEN|47|24|将来收割的时候，你们要把五分之一纳给法老，另外四分可以给你们作田地的种子，作你们和你们全家大小的食物。”
GEN|47|25|他们说：“你救了我们的性命，愿我们在我主眼前蒙恩，我们情愿作法老的奴隶。”
GEN|47|26|于是 约瑟 为 埃及 的土地立下定例，直到今日，就是收成的五分之一要归法老。惟独祭司的土地例外，不归于法老。
GEN|47|27|以色列 人住在 埃及 境内的 歌珊 地。他们在那里得了产业，并且生养众多。
GEN|47|28|雅各 住在 埃及 地十七年。 雅各 一生的年日是一百四十七年。
GEN|47|29|以色列 的死期快到了，就叫了他儿子 约瑟 来，对他说：“我若在你眼前蒙恩，把你的手放在我大腿底下，以慈爱和诚实向我承诺，必不将我葬在 埃及 。
GEN|47|30|我与我祖先同睡的时候，你要将我带出 埃及 ，把我葬在他们所葬的地方。” 约瑟 说：“我必遵照你的吩咐去做。”
GEN|47|31|雅各 说：“你向我起誓吧！” 约瑟 就向他起了誓。于是 以色列 在床头 敬拜。
GEN|48|1|这些事以后，有人告诉 约瑟 说：“看哪，你的父亲病了。”他就带着两个儿子 玛拿西 和 以法莲 同去。
GEN|48|2|有人告诉 雅各 说：“看哪，你的儿子 约瑟 到你这里来了。” 以色列 就勉强在床上坐起来。
GEN|48|3|雅各 对 约瑟 说：“全能的上帝曾在 迦南 地的 路斯 向我显现，赐福给我，
GEN|48|4|对我说：‘看哪，我必使你生养众多，成为许多民族，又要将这地赐给你的后裔，永远为业。’
GEN|48|5|我未到 埃及 你那里之前，你在 埃及 地所生的 以法莲 和 玛拿西 这两个儿子，现在他们是我的，正如 吕便 和 西缅 是我的一样。
GEN|48|6|你在他们以后所生的后裔就是你的，这些后裔可以在自己兄弟的名下得产业。
GEN|48|7|至于我，我从 巴旦 回来的时候， 拉结 在我身旁死了，就是在往 迦南 地的路上，离 以法他 还有一段路程。我就把她葬在往 以法他 的路旁； 以法他 就是 伯利恒 。”
GEN|48|8|以色列 看见 约瑟 的儿子，就说：“这些是谁？”
GEN|48|9|约瑟 对他父亲说：“这是上帝在这里赐给我的儿子。” 以色列 说：“领他们到我跟前，我要为他们祝福。”
GEN|48|10|以色列 年纪老迈，眼睛昏花，不能看见。 约瑟 领他们到他跟前，他就和他们亲吻，抱着他们。
GEN|48|11|以色列 对 约瑟 说：“我没有想到能够见你的面。看哪，上帝还让我看见你的儿子。”
GEN|48|12|约瑟 把他们从 以色列 两膝中间领出来，自己脸伏于地下拜。
GEN|48|13|然后， 约瑟 牵着他们两个，带到父亲跟前，右手牵 以法莲 到 以色列 的左边，左手牵 玛拿西 到 以色列 的右边。
GEN|48|14|以色列 却伸出右手来，按在次子 以法莲 的头上，又交叉伸出左手来，按在长子 玛拿西 的头上。
GEN|48|15|他就为 约瑟 祝福说： “愿我祖父 亚伯拉罕 和我父亲 以撒 所事奉的上帝， 就是一生牧养我直到今日的上帝，
GEN|48|16|救赎我脱离一切患难的那位使者，赐福给这两个孩子。 愿我的名，我祖父 亚伯拉罕 和我父亲 以撒 的名藉着他们得以流传。 又愿他们在全地上多多繁衍。”
GEN|48|17|约瑟 见父亲把右手按在 以法莲 的头上，他看为不好，就提起他父亲的手，要从 以法莲 的头上移到 玛拿西 的头上。
GEN|48|18|约瑟 对父亲说：“我父，不是这样。这个才是长子，请你把右手按在他头上。”
GEN|48|19|他父亲却不肯，说：“我知道，我儿，我知道。他也要成为一族，也要强大。可是他的弟弟将来比他还要强大；他弟弟的后裔要成为许多国家。”
GEN|48|20|以色列 就在当日为他们祝福，说：“ 以色列 人要指着你们祝福，说：‘愿上帝使你如 以法莲 、 玛拿西 一样。’”于是他立 以法莲 在 玛拿西 之上。
GEN|48|21|以色列 又对 约瑟 说：“看哪，我快要死了，但上帝必与你们同在，领你们回到你们祖先之地。
GEN|48|22|从前我用刀用弓从 亚摩利 人手下夺取的那一份，我要把它赐给你，使你比你的兄弟多得一份 。”
GEN|49|1|雅各 叫了他的儿子来，说：“你们都来聚集，让我把你们日后要遇到的事告诉你们。
GEN|49|2|雅各 的儿子们，你们要聚集，要聆听， 听你们父亲 以色列 的话。
GEN|49|3|吕便 啊，你是我的长子，我的力量， 我壮年头生之子， 极有尊荣，权力超群。
GEN|49|4|你却放纵如水，必不得居首位； 因为你上了你父亲的床， 你 上了我的榻，污辱了它！
GEN|49|5|西缅 和 利未 是兄弟； 他们的刀剑是残暴的兵器。
GEN|49|6|愿我的心不与他们同谋， 愿我的灵 不与他们合伙； 因为他们在烈怒中杀人， 任意割断牛腿的筋。
GEN|49|7|他们火爆的烈怒可诅， 他们凶残的愤恨可咒！ 我要把他们分散在 雅各 中， 使他们散居在 以色列 。
GEN|49|8|犹大 啊，你的兄弟必赞美你， 你的手必掐住仇敌的颈项， 你父亲的儿子要向你下拜。
GEN|49|9|犹大 是只小狮子； 我儿啊，你捕获了猎物就上去。 他蹲伏，他躺卧，如公狮， 又如母狮，谁敢惹他呢？
GEN|49|10|权杖必不离 犹大 ， 统治者的杖必不离他两脚之间， 直等细罗 来到， 万民都要归顺他。
GEN|49|11|犹大 把小驴拴在葡萄树上， 把驴驹拴在佳美的葡萄树上。 他在葡萄酒中洗衣服， 在葡萄汁 中洗长袍。
GEN|49|12|他的眼睛比 酒红润， 他的牙齿比奶洁白。
GEN|49|13|西布伦 必住在海边， 必成为停船的港口； 他的疆界必延到 西顿 。
GEN|49|14|以萨迦 是匹强壮的驴， 卧在羊圈之中。
GEN|49|15|他看见居所安舒， 土地肥美， 就屈肩负重， 成为服劳役的仆人。
GEN|49|16|但 必为他的百姓伸冤 ， 作为 以色列 支派之一。
GEN|49|17|但 必作道旁的蛇， 路边的毒蛇， 咬伤马蹄， 使骑马的人向后坠落。
GEN|49|18|耶和华啊，我等候你的救恩。
GEN|49|19|迦得 必被袭击者袭击 ， 他却要袭击他们的脚跟。
GEN|49|20|亚设 必出丰盛的粮食， 要供应君王的佳肴。
GEN|49|21|拿弗他利 是被释放的母鹿， 他要生出可爱的小鹿 。
GEN|49|22|约瑟 是多结果子的树枝， 是泉旁多结果的枝子； 他的枝条伸出墙外。
GEN|49|23|弓箭手恶意攻击他， 敌对他，向他射箭。
GEN|49|24|但他的弓仍旧坚硬， 他的手臂灵活敏捷， 这是因 雅各 的大能者的手， 从那里，他是 以色列 的牧者， 以色列 的磐石 。
GEN|49|25|你父亲的上帝必帮助你； 全能者必赐福给你： 天上的福， 深渊下面蕴藏的福， 以及生育哺养的福。
GEN|49|26|你父亲的福 胜过我祖先的福， 直到永世山岭的极限。 这些福必降在 约瑟 的头上， 临到那与兄弟有分别之人的头顶上。
GEN|49|27|便雅悯 是只抓撕掠物的狼， 早晨要吃他的猎物， 晚上要分他的掳物。”
GEN|49|28|这一切是 以色列 的十二个支派。这是他们的父亲对他们所说的话，他按照各人的福分为他们祝福。
GEN|49|29|他又吩咐他们说：“我快要归到我祖先 那里。你们要将我葬在 赫 人 以弗仑 田间的洞里，与我的祖先在一处，
GEN|49|30|就是在 迦南 地 幔利 对面的 麦比拉 田间的洞里，那田是 亚伯拉罕 向 赫 人 以弗仑 买来作坟地的产业。
GEN|49|31|亚伯拉罕 和他的妻子 撒拉 葬在那里； 以撒 和他的妻子 利百加 也葬在那里。我也在那里葬了 利亚 。
GEN|49|32|那块田和田间的洞是向 赫 人买的。”
GEN|49|33|雅各 嘱咐众子完毕后，就把脚收在床上断了气，归到他祖先 那里去了。
GEN|50|1|约瑟 伏在他父亲的脸上，在他脸上哭，又亲他。
GEN|50|2|约瑟 吩咐伺候他的医生们用香料涂他父亲，医生就用香料涂了 以色列 。
GEN|50|3|四十天满了，就是涂香料所规定的日子满了。 埃及 人为他哀哭了七十天。
GEN|50|4|过了哀悼的日子， 约瑟 对法老家中的人说：“我若在你们眼前蒙恩，请你们对法老说：
GEN|50|5|‘我父亲曾叫我起誓说：看哪，我快要死了，你要将我葬在 迦南 地，在我为自己所掘的坟墓里。’现在求你准我上去葬我父亲，然后我必回来。”
GEN|50|6|法老说：“你可以上去，照你父亲叫你起的誓，将他安葬。”
GEN|50|7|于是 约瑟 上去葬他父亲。与他一同上去的有法老的众臣仆和法老家中的长老，以及 埃及 地所有的长老，
GEN|50|8|还有 约瑟 的全家和他的兄弟们，以及他父亲的家属；只留下他们的孩子和羊群牛群在 歌珊 地。
GEN|50|9|又有车辆和驾驶兵和他一同上去，队伍非常庞大。
GEN|50|10|他们到了 约旦河 东 亚达 的禾场，就在那里大大地号啕痛哭。 约瑟 为他父亲哀哭了七天。
GEN|50|11|迦南 的居民看见 亚达 禾场上的哀哭，就说：“这是 埃及 人一场极大的哀哭。”因此那地方名叫 亚伯．麦西 ，是在 约旦河 东。
GEN|50|12|雅各 的儿子们遵照父亲的吩咐去办了，
GEN|50|13|他们把他送到 迦南 地，葬在 幔利 对面的 麦比拉 田间的洞里；那田是 亚伯拉罕 向 赫 人 以弗仑 买来作坟地的产业。
GEN|50|14|约瑟 葬了他父亲以后，就和他的兄弟，以及所有同他上去葬他父亲的人，都回 埃及 去了。
GEN|50|15|约瑟 的哥哥们见父亲死了，就说：“也许 约瑟 仍然怀恨我们，会照我们从前待他一切的恶，重重报复我们。”
GEN|50|16|他们就传口信给 约瑟 说：“你父亲未死之前曾吩咐说：
GEN|50|17|‘你们要对 约瑟 这样说：从前你哥哥们恶待你，你要饶恕他们的过犯和罪恶。’现在求你饶恕你父亲的上帝之仆人们的过犯。”他们对 约瑟 说了这话， 约瑟 就哭了。
GEN|50|18|他的哥哥们又来俯伏在他面前，说：“看哪，我们是你的奴隶。”
GEN|50|19|约瑟 对他们说：“不要怕，我岂能代替上帝呢？
GEN|50|20|从前你们的意思是要害我，但上帝的意思原是好的，要使许多百姓得以存活，成就今日的光景。
GEN|50|21|现在你们不要害怕，我必养活你们和你们的孩子。”于是 约瑟 安慰他们，讲了使他们安心的话。
GEN|50|22|约瑟 和他父亲的家属都住在 埃及 。 约瑟 活了一百一十年。
GEN|50|23|约瑟 看到 以法莲 第三代的子孙。 玛拿西 的孙子， 玛吉 的儿子，出生时都放在 约瑟 的膝上。
GEN|50|24|约瑟 对他的兄弟说：“我快要死了，但上帝必定看顾你们，领你们从这地上去，到他起誓应许给 亚伯拉罕 、 以撒 、 雅各 之地。”
GEN|50|25|约瑟 叫 以色列 的子孙起誓：“上帝必定眷顾你们，你们要把我的骸骨从这里带上去。”
GEN|50|26|约瑟 死了，那时他一百一十岁。人用香料涂了他，把他收殓在棺材里，停放在 埃及 。
