JOHN|1|1|In the beginning was the Word, and the Word was with God, and the Word was God.
JOHN|1|2|He was in the beginning with God.
JOHN|1|3|All things were made through him, and without him was not any thing made that was made.
JOHN|1|4|In him was life, and the life was the light of men.
JOHN|1|5|The light shines in the darkness, and the darkness has not overcome it.
JOHN|1|6|There was a man sent from God, whose name was John.
JOHN|1|7|He came as a witness, to bear witness about the light, that all might believe through him.
JOHN|1|8|He was not the light, but came to bear witness about the light.
JOHN|1|9|The true light, which enlightens everyone, was coming into the world.
JOHN|1|10|He was in the world, and the world was made through him, yet the world did not know him.
JOHN|1|11|He came to his own, and his own people did not receive him.
JOHN|1|12|But to all who did receive him, who believed in his name, he gave the right to become children of God.
JOHN|1|13|who were born, not of blood nor of the will of the flesh nor of the will of man, but of God.
JOHN|1|14|And the Word became flesh and dwelt among us, and we have seen his glory, glory as of the only Son from the Father, full of grace and truth.
JOHN|1|15|(John bore witness about him, and cried out, "This was he of whom I said, 'He who comes after me ranks before me, because he was before me.'")
JOHN|1|16|And from his fullness we have all received, grace upon grace.
JOHN|1|17|For the law was given through Moses; grace and truth came through Jesus Christ.
JOHN|1|18|No one has ever seen God; the only God, who is at the Father's side, he has made him known.
JOHN|1|19|And this is the testimony of John, when the Jews sent priests and Levites from Jerusalem to ask him, "Who are you?"
JOHN|1|20|He confessed, and did not deny, but confessed, "I am not the Christ."
JOHN|1|21|And they asked him, "What then? Are you Elijah?" He said, "I am not." "Are you the Prophet?" And he answered, "No."
JOHN|1|22|So they said to him, "Who are you? We need to give an answer to those who sent us. What do you say about yourself?"
JOHN|1|23|He said, "I am the voice of one crying out in the wilderness, 'Make straight the way of the Lord,' as the prophet Isaiah said."
JOHN|1|24|(Now they had been sent from the Pharisees.)
JOHN|1|25|They asked him, "Then why are you baptizing, if you are neither the Christ, nor Elijah, nor the Prophet?"
JOHN|1|26|John answered them, "I baptize with water, but among you stands one you do not know,
JOHN|1|27|even he who comes after me, the strap of whose sandal I am not worthy to untie."
JOHN|1|28|These things took place in Bethany across the Jordan, where John was baptizing.
JOHN|1|29|The next day he saw Jesus coming toward him, and said, "Behold, the Lamb of God, who takes away the sin of the world!
JOHN|1|30|This is he of whom I said, 'After me comes a man who ranks before me, because he was before me.'
JOHN|1|31|I myself did not know him, but for this purpose I came baptizing with water, that he might be revealed to Israel."
JOHN|1|32|And John bore witness: "I saw the Spirit descend from heaven like a dove, and it remained on him.
JOHN|1|33|I myself did not know him, but he who sent me to baptize with water said to me, 'He on whom you see the Spirit descend and remain, this is he who baptizes with the Holy Spirit.'
JOHN|1|34|And I have seen and have borne witness that this is the Son of God."
JOHN|1|35|The next day again John was standing with two of his disciples,
JOHN|1|36|and he looked at Jesus as he walked by and said, "Behold, the Lamb of God!"
JOHN|1|37|The two disciples heard him say this, and they followed Jesus.
JOHN|1|38|Jesus turned and saw them following and said to them, "What are you seeking?" And they said to him, "Rabbi" (which means Teacher), "where are you staying?"
JOHN|1|39|He said to them, "Come and you will see." So they came and saw where he was staying, and they stayed with him that day, for it was about the tenth hour.
JOHN|1|40|One of the two who heard John speak and followed Jesus was Andrew, Simon Peter's brother.
JOHN|1|41|He first found his own brother Simon and said to him, "We have found the Messiah" (which means Christ).
JOHN|1|42|He brought him to Jesus. Jesus looked at him and said, "So you are Simon the son of John? You shall be called Cephas" (which means Peter).
JOHN|1|43|The next day Jesus decided to go to Galilee. He found Philip and said to him, "Follow me."
JOHN|1|44|Now Philip was from Bethsaida, the city of Andrew and Peter.
JOHN|1|45|Philip found Nathanael and said to him, "We have found him of whom Moses in the Law and also the prophets wrote, Jesus of Nazareth, the son of Joseph."
JOHN|1|46|Nathanael said to him, "Can anything good come out of Nazareth?" Philip said to him, "Come and see."
JOHN|1|47|Jesus saw Nathanael coming toward him and said of him, "Behold, an Israelite indeed, in whom there is no deceit!"
JOHN|1|48|Nathanael said to him, "How do you know me?" Jesus answered him, "Before Philip called you, when you were under the fig tree, I saw you."
JOHN|1|49|Nathanael answered him, "Rabbi, you are the Son of God! You are the King of Israel!"
JOHN|1|50|Jesus answered him, "Because I said to you, 'I saw you under the fig tree,' do you believe? You will see greater things than these."
JOHN|1|51|And he said to him, "Truly, truly, I say to you, you will see heaven opened, and the angels of God ascending and descending on the Son of Man."
JOHN|2|1|On the third day there was a wedding at Cana in Galilee, and the mother of Jesus was there.
JOHN|2|2|Jesus also was invited to the wedding with his disciples.
JOHN|2|3|When the wine ran out, the mother of Jesus said to him, "They have no wine."
JOHN|2|4|And Jesus said to her, "Woman, what does this have to do with me? My hour has not yet come."
JOHN|2|5|His mother said to the servants, "Do whatever he tells you."
JOHN|2|6|Now there were six stone water jars there for the Jewish rites of purification, each holding twenty or thirty gallons.
JOHN|2|7|Jesus said to the servants, "Fill the jars with water." And they filled them up to the brim.
JOHN|2|8|And he said to them, "Now draw some out and take it to the master of the feast." So they took it.
JOHN|2|9|When the master of the feast tasted the water now become wine, and did not know where it came from (though the servants who had drawn the water knew), the master of the feast called the bridegroom
JOHN|2|10|and said to him, "Everyone serves the good wine first, and when people have drunk freely, then the poor wine. But you have kept the good wine until now."
JOHN|2|11|This, the first of his signs, Jesus did at Cana in Galilee, and manifested his glory. And his disciples believed in him.
JOHN|2|12|After this he went down to Capernaum, with his mother and his brothers and his disciples, and they stayed there for a few days.
JOHN|2|13|The Passover of the Jews was at hand, and Jesus went up to Jerusalem.
JOHN|2|14|In the temple he found those who were selling oxen and sheep and pigeons, and the money-changers sitting there.
JOHN|2|15|And making a whip of cords, he drove them all out of the temple, with the sheep and oxen. And he poured out the coins of the money-changers and overturned their tables.
JOHN|2|16|And he told those who sold the pigeons, "Take these things away; do not make my Father's house a house of trade."
JOHN|2|17|His disciples remembered that it was written, "Zeal for your house will consume me."
JOHN|2|18|So the Jews said to him, "What sign do you show us for doing these things?"
JOHN|2|19|Jesus answered them, "Destroy this temple, and in three days I will raise it up."
JOHN|2|20|The Jews then said, "It has taken forty-six years to build this temple, and will you raise it up in three days?"
JOHN|2|21|But he was speaking about the temple of his body.
JOHN|2|22|When therefore he was raised from the dead, his disciples remembered that he had said this, and they believed the Scripture and the word that Jesus had spoken.
JOHN|2|23|Now when he was in Jerusalem at the Passover Feast, many believed in his name when they saw the signs that he was doing.
JOHN|2|24|But Jesus on his part did not entrust himself to them, because he knew all people
JOHN|2|25|and needed no one to bear witness about man, for he himself knew what was in man.
JOHN|3|1|Now there was a man of the Pharisees named Nicodemus, a ruler of the Jews.
JOHN|3|2|This man came to Jesus by night and said to him, "Rabbi, we know that you are a teacher come from God, for no one can do these signs that you do unless God is with him."
JOHN|3|3|Jesus answered him, "Truly, truly, I say to you, unless one is born again he cannot see the kingdom of God."
JOHN|3|4|Nicodemus said to him, "How can a man be born when he is old? Can he enter a second time into his mother's womb and be born?"
JOHN|3|5|Jesus answered, "Truly, truly, I say to you, unless one is born of water and the Spirit, he cannot enter the kingdom of God.
JOHN|3|6|That which is born of the flesh is flesh, and that which is born of the Spirit is spirit.
JOHN|3|7|Do not marvel that I said to you, 'You must be born again.'
JOHN|3|8|The wind blows where it wishes, and you hear its sound, but you do not know where it comes from or where it goes. So it is with everyone who is born of the Spirit."
JOHN|3|9|Nicodemus said to him, "How can these things be?"
JOHN|3|10|Jesus answered him, "Are you the teacher of Israel and yet you do not understand these things?
JOHN|3|11|Truly, truly, I say to you, we speak of what we know, and bear witness to what we have seen, but you do not receive our testimony.
JOHN|3|12|If I have told you earthly things and you do not believe, how can you believe if I tell you heavenly things?
JOHN|3|13|No one has ascended into heaven except him who descended from heaven, the Son of Man.
JOHN|3|14|And as Moses lifted up the serpent in the wilderness, so must the Son of Man be lifted up,
JOHN|3|15|that whoever believes in him may have eternal life."
JOHN|3|16|For God so loved the world, that he gave his only Son, that whoever believes in him should not perish but have eternal life.
JOHN|3|17|For God did not send his Son into the world to condemn the world, but in order that the world might be saved through him.
JOHN|3|18|Whoever believes in him is not condemned, but whoever does not believe is condemned already, because he has not believed in the name of the only Son of God.
JOHN|3|19|And this is the judgment: the light has come into the world, and people loved the darkness rather than the light because their deeds were evil.
JOHN|3|20|For everyone who does wicked things hates the light and does not come to the light, lest his deeds should be exposed.
JOHN|3|21|But whoever does what is true comes to the light, so that it may be clearly seen that his deeds have been carried out in God.
JOHN|3|22|After this Jesus and his disciples went into the Judean countryside, and he remained there with them and was baptizing.
JOHN|3|23|John also was baptizing at Aenon near Salim, because water was plentiful there, and people were coming and being baptized
JOHN|3|24|(for John had not yet been put in prison).
JOHN|3|25|Now a discussion arose between some of John's disciples and a Jew over purification.
JOHN|3|26|And they came to John and said to him, "Rabbi, he who was with you across the Jordan, to whom you bore witness- look, he is baptizing, and all are going to him."
JOHN|3|27|John answered, "A person cannot receive even one thing unless it is given him from heaven.
JOHN|3|28|You yourselves bear me witness, that I said, 'I am not the Christ, but I have been sent before him.'
JOHN|3|29|The one who has the bride is the bridegroom. The friend of the bridegroom, who stands and hears him, rejoices greatly at the bridegroom's voice. Therefore this joy of mine is now complete.
JOHN|3|30|He must increase, but I must decrease."
JOHN|3|31|He who comes from above is above all. He who is of the earth belongs to the earth and speaks in an earthly way. He who comes from heaven is above all.
JOHN|3|32|He bears witness to what he has seen and heard, yet no one receives his testimony.
JOHN|3|33|Whoever receives his testimony sets his seal to this, that God is true.
JOHN|3|34|For he whom God has sent utters the words of God, for he gives the Spirit without measure.
JOHN|3|35|The Father loves the Son and has given all things into his hand.
JOHN|3|36|Whoever believes in the Son has eternal life; whoever does not obey the Son shall not see life, but the wrath of God remains on him.
JOHN|4|1|Now when Jesus learned that the Pharisees had heard that Jesus was making and baptizing more disciples than John
JOHN|4|2|(although Jesus himself did not baptize, but only his disciples),
JOHN|4|3|he left Judea and departed again for Galilee.
JOHN|4|4|And he had to pass through Samaria.
JOHN|4|5|So he came to a town of Samaria called Sychar, near the field that Jacob had given to his son Joseph.
JOHN|4|6|Jacob's well was there; so Jesus, wearied as he was from his journey, was sitting beside the well. It was about the sixth hour.
JOHN|4|7|There came a woman of Samaria to draw water. Jesus said to her, "Give me a drink."
JOHN|4|8|(For his disciples had gone away into the city to buy food.)
JOHN|4|9|The Samaritan woman said to him, "How is it that you, a Jew, ask for a drink from me, a woman of Samaria?" (For Jews have no dealings with Samaritans.)
JOHN|4|10|Jesus answered her, "If you knew the gift of God, and who it is that is saying to you, 'Give me a drink,' you would have asked him, and he would have given you living water."
JOHN|4|11|The woman said to him, "Sir, you have nothing to draw water with, and the well is deep. Where do you get that living water?
JOHN|4|12|Are you greater than our father Jacob? He gave us the well and drank from it himself, as did his sons and his livestock."
JOHN|4|13|Jesus said to her, "Everyone who drinks of this water will be thirsty again,
JOHN|4|14|but whoever drinks of the water that I will give him will never be thirsty forever. The water that I will give him will become in him a spring of water welling up to eternal life."
JOHN|4|15|The woman said to him, "Sir, give me this water, so that I will not be thirsty or have to come here to draw water."
JOHN|4|16|Jesus said to her, "Go, call your husband, and come here."
JOHN|4|17|The woman answered him, "I have no husband." Jesus said to her, "You are right in saying, 'I have no husband';
JOHN|4|18|for you have had five husbands, and the one you now have is not your husband. What you have said is true."
JOHN|4|19|The woman said to him, "Sir, I perceive that you are a prophet.
JOHN|4|20|Our fathers worshiped on this mountain, but you say that in Jerusalem is the place where people ought to worship."
JOHN|4|21|Jesus said to her, "Woman, believe me, the hour is coming when neither on this mountain nor in Jerusalem will you worship the Father.
JOHN|4|22|You worship what you do not know; we worship what we know, for salvation is from the Jews.
JOHN|4|23|But the hour is coming, and is now here, when the true worshipers will worship the Father in spirit and truth, for the Father is seeking such people to worship him.
JOHN|4|24|God is spirit, and those who worship him must worship in spirit and truth."
JOHN|4|25|The woman said to him, "I know that Messiah is coming (he who is called Christ). When he comes, he will tell us all things."
JOHN|4|26|Jesus said to her, "I who speak to you am he."
JOHN|4|27|Just then his disciples came back. They marveled that he was talking with a woman, but no one said, "What do you seek?" or, "Why are you talking with her?"
JOHN|4|28|So the woman left her water jar and went away into town and said to the people,
JOHN|4|29|"Come, see a man who told me all that I ever did. Can this be the Christ?"
JOHN|4|30|They went out of the town and were coming to him.
JOHN|4|31|Meanwhile the disciples were urging him, saying, "Rabbi, eat."
JOHN|4|32|But he said to them, "I have food to eat that you do not know about."
JOHN|4|33|So the disciples said to one another, "Has anyone brought him something to eat?"
JOHN|4|34|Jesus said to them, "My food is to do the will of him who sent me and to accomplish his work.
JOHN|4|35|Do you not say, 'There are yet four months, then comes the harvest'? Look, I tell you, lift up your eyes, and see that the fields are white for harvest.
JOHN|4|36|Already the one who reaps is receiving wages and gathering fruit for eternal life, so that sower and reaper may rejoice together.
JOHN|4|37|For here the saying holds true, 'One sows and another reaps.'
JOHN|4|38|I sent you to reap that for which you did not labor. Others have labored, and you have entered into their labor."
JOHN|4|39|Many Samaritans from that town believed in him because of the woman's testimony, "He told me all that I ever did."
JOHN|4|40|So when the Samaritans came to him, they asked him to stay with them, and he stayed there two days.
JOHN|4|41|And many more believed because of his word.
JOHN|4|42|They said to the woman, "It is no longer because of what you said that we believe, for we have heard for ourselves, and we know that this is indeed the Savior of the world."
JOHN|4|43|After the two days he departed for Galilee.
JOHN|4|44|(For Jesus himself had testified that a prophet has no honor in his own hometown.)
JOHN|4|45|So when he came to Galilee, the Galileans welcomed him, having seen all that he had done in Jerusalem at the feast. For they too had gone to the feast.
JOHN|4|46|So he came again to Cana in Galilee, where he had made the water wine. And at Capernaum there was an official whose son was ill.
JOHN|4|47|When this man heard that Jesus had come from Judea to Galilee, he went to him and asked him to come down and heal his son, for he was at the point of death.
JOHN|4|48|So Jesus said to him, "Unless you see signs and wonders you will not believe."
JOHN|4|49|The official said to him, "Sir, come down before my child dies."
JOHN|4|50|Jesus said to him, "Go; your son will live." The man believed the word that Jesus spoke to him and went on his way.
JOHN|4|51|As he was going down, his servants met him and told him that his son was recovering.
JOHN|4|52|So he asked them the hour when he began to get better, and they said to him, "Yesterday at the seventh hour the fever left him."
JOHN|4|53|The father knew that was the hour when Jesus had said to him, "Your son will live." And he himself believed, and all his household.
JOHN|4|54|This was now the second sign that Jesus did when he had come from Judea to Galilee.
JOHN|5|1|After this there was a feast of the Jews, and Jesus went up to Jerusalem.
JOHN|5|2|Now there is in Jerusalem by the Sheep Gate a pool, in Aramaic called Bethesda, which has five roofed colonnades.
JOHN|5|3|In these lay a multitude of invalids- blind, lame, and paralyzed.
JOHN|5|4|***
JOHN|5|5|One man was there who had been an invalid for thirty-eight years.
JOHN|5|6|When Jesus saw him lying there and knew that he had already been there a long time, he said to him, "Do you want to be healed?"
JOHN|5|7|The sick man answered him, "Sir, I have no one to put me into the pool when the water is stirred up, and while I am going another steps down before me."
JOHN|5|8|Jesus said to him, "Get up, take up your bed, and walk."
JOHN|5|9|And at once the man was healed, and he took up his bed and walked. Now that day was the Sabbath.
JOHN|5|10|So the Jews said to the man who had been healed, "It is the Sabbath, and it is not lawful for you to take up your bed."
JOHN|5|11|But he answered them, "The man who healed me, that man said to me, 'Take up your bed, and walk.'"
JOHN|5|12|They asked him, "Who is the man who said to you, 'Take up your bed and walk'?"
JOHN|5|13|Now the man who had been healed did not know who it was, for Jesus had withdrawn, as there was a crowd in the place.
JOHN|5|14|Afterward Jesus found him in the temple and said to him, "See, you are well! Sin no more, that nothing worse may happen to you."
JOHN|5|15|The man went away and told the Jews that it was Jesus who had healed him.
JOHN|5|16|And this was why the Jews were persecuting Jesus, because he was doing these things on the Sabbath.
JOHN|5|17|But Jesus answered them, "My Father is working until now, and I am working."
JOHN|5|18|This was why the Jews were seeking all the more to kill him, because not only was he breaking the Sabbath, but he was even calling God his own Father, making himself equal with God.
JOHN|5|19|So Jesus said to them, "Truly, truly, I say to you, the Son can do nothing of his own accord, but only what he sees the Father doing. For whatever the Father does, that the Son does likewise.
JOHN|5|20|For the Father loves the Son and shows him all that he himself is doing. And greater works than these will he show him, so that you may marvel.
JOHN|5|21|For as the Father raises the dead and gives them life, so also the Son gives life to whom he will.
JOHN|5|22|The Father judges no one, but has given all judgment to the Son,
JOHN|5|23|that all may honor the Son, just as they honor the Father. Whoever does not honor the Son does not honor the Father who sent him.
JOHN|5|24|Truly, truly, I say to you, whoever hears my word and believes him who sent me has eternal life. He does not come into judgment, but has passed from death to life.
JOHN|5|25|"Truly, truly, I say to you, an hour is coming, and is now here, when the dead will hear the voice of the Son of God, and those who hear will live.
JOHN|5|26|For as the Father has life in himself, so he has granted the Son also to have life in himself.
JOHN|5|27|And he has given him authority to execute judgment, because he is the Son of Man.
JOHN|5|28|Do not marvel at this, for an hour is coming when all who are in the tombs will hear his voice
JOHN|5|29|and come out, those who have done good to the resurrection of life, and those who have done evil to the resurrection of judgment.
JOHN|5|30|"I can do nothing on my own. As I hear, I judge, and my judgment is just, because I seek not my own will but the will of him who sent me.
JOHN|5|31|If I alone bear witness about myself, my testimony is not deemed true.
JOHN|5|32|There is another who bears witness about me, and I know that the testimony that he bears about me is true.
JOHN|5|33|You sent to John, and he has borne witness to the truth.
JOHN|5|34|Not that the testimony that I receive is from man, but I say these things so that you may be saved.
JOHN|5|35|He was a burning and shining lamp, and you were willing to rejoice for a while in his light.
JOHN|5|36|But the testimony that I have is greater than that of John. For the works that the Father has given me to accomplish, the very works that I am doing, bear witness about me that the Father has sent me.
JOHN|5|37|And the Father who sent me has himself borne witness about me. His voice you have never heard, his form you have never seen,
JOHN|5|38|and you do not have his word abiding in you, for you do not believe the one whom he has sent.
JOHN|5|39|You search the Scriptures because you think that in them you have eternal life; and it is they that bear witness about me,
JOHN|5|40|yet you refuse to come to me that you may have life.
JOHN|5|41|I do not receive glory from people.
JOHN|5|42|But I know that you do not have the love of God within you.
JOHN|5|43|I have come in my Father's name, and you do not receive me. If another comes in his own name, you will receive him.
JOHN|5|44|How can you believe, when you receive glory from one another and do not seek the glory that comes from the only God?
JOHN|5|45|Do not think that I will accuse you to the Father. There is one who accuses you: Moses, on whom you have set your hope.
JOHN|5|46|If you believed Moses, you would believe me; for he wrote of me.
JOHN|5|47|But if you do not believe his writings, how will you believe my words?"
JOHN|6|1|After this Jesus went away to the other side of the Sea of Galilee, which is the Sea of Tiberias.
JOHN|6|2|And a large crowd was following him, because they saw the signs that he was doing on the sick.
JOHN|6|3|Jesus went up on the mountain, and there he sat down with his disciples.
JOHN|6|4|Now the Passover, the feast of the Jews, was at hand.
JOHN|6|5|Lifting up his eyes, then, and seeing that a large crowd was coming toward him, Jesus said to Philip, "Where are we to buy bread, so that these people may eat?"
JOHN|6|6|He said this to test him, for he himself knew what he would do.
JOHN|6|7|Philip answered him, "Two hundred denarii would not buy enough bread for each of them to get a little."
JOHN|6|8|One of his disciples, Andrew, Simon Peter's brother, said to him,
JOHN|6|9|"There is a boy here who has five barley loaves and two fish, but what are they for so many?"
JOHN|6|10|Jesus said, "Have the people sit down." Now there was much grass in the place. So the men sat down, about five thousand in number.
JOHN|6|11|Jesus then took the loaves, and when he had given thanks, he distributed them to those who were seated. So also the fish, as much as they wanted.
JOHN|6|12|And when they had eaten their fill, he told his disciples, "Gather up the leftover fragments, that nothing may be lost."
JOHN|6|13|So they gathered them up and filled twelve baskets with fragments from the five barley loaves, left by those who had eaten.
JOHN|6|14|When the people saw the sign that he had done, they said, "This is indeed the Prophet who is to come into the world!"
JOHN|6|15|Perceiving then that they were about to come and take him by force to make him king, Jesus withdrew again to the mountain by himself.
JOHN|6|16|When evening came, his disciples went down to the sea,
JOHN|6|17|got into a boat, and started across the sea to Capernaum. It was now dark, and Jesus had not yet come to them.
JOHN|6|18|The sea became rough because a strong wind was blowing.
JOHN|6|19|When they had rowed about three or four miles, they saw Jesus walking on the sea and coming near the boat, and they were frightened.
JOHN|6|20|But he said to them, "It is I; do not be afraid."
JOHN|6|21|Then they were glad to take him into the boat, and immediately the boat was at the land to which they were going.
JOHN|6|22|On the next day the crowd that remained on the other side of the sea saw that there had been only one boat there, and that Jesus had not entered the boat with his disciples, but that his disciples had gone away alone.
JOHN|6|23|Other boats from Tiberias came near the place where they had eaten the bread after the Lord had given thanks.
JOHN|6|24|So when the crowd saw that Jesus was not there, nor his disciples, they themselves got into the boats and went to Capernaum, seeking Jesus.
JOHN|6|25|When they found him on the other side of the sea, they said to him, "Rabbi, when did you come here?"
JOHN|6|26|Jesus answered them, "Truly, truly, I say to you, you are seeking me, not because you saw signs, but because you ate your fill of the loaves.
JOHN|6|27|Do not labor for the food that perishes, but for the food that endures to eternal life, which the Son of Man will give to you. For on him God the Father has set his seal."
JOHN|6|28|Then they said to him, "What must we do, to be doing the works of God?"
JOHN|6|29|Jesus answered them, "This is the work of God, that you believe in him whom he has sent."
JOHN|6|30|So they said to him, "Then what sign do you do, that we may see and believe you? What work do you perform?
JOHN|6|31|Our fathers ate the manna in the wilderness; as it is written, 'He gave them bread from heaven to eat.'"
JOHN|6|32|Jesus then said to them, "Truly, truly, I say to you, it was not Moses who gave you the bread from heaven, but my Father gives you the true bread from heaven.
JOHN|6|33|For the bread of God is he who comes down from heaven and gives life to the world."
JOHN|6|34|They said to him, "Sir, give us this bread always."
JOHN|6|35|Jesus said to them, "I am the bread of life; whoever comes to me shall not hunger, and whoever believes in me shall never thirst.
JOHN|6|36|But I said to you that you have seen me and yet do not believe.
JOHN|6|37|All that the Father gives me will come to me, and whoever comes to me I will never cast out.
JOHN|6|38|For I have come down from heaven, not to do my own will but the will of him who sent me.
JOHN|6|39|And this is the will of him who sent me, that I should lose nothing of all that he has given me, but raise it up on the last day.
JOHN|6|40|For this is the will of my Father, that everyone who looks on the Son and believes in him should have eternal life, and I will raise him up on the last day."
JOHN|6|41|So the Jews grumbled about him, because he said, "I am the bread that came down from heaven."
JOHN|6|42|They said, "Is not this Jesus, the son of Joseph, whose father and mother we know? How does he now say, 'I have come down from heaven'?"
JOHN|6|43|Jesus answered them, "Do not grumble among yourselves.
JOHN|6|44|No one can come to me unless the Father who sent me draws him. And I will raise him up on the last day.
JOHN|6|45|It is written in the Prophets, 'And they will all be taught by God.' Everyone who has heard and learned from the Father comes to me-
JOHN|6|46|not that anyone has seen the Father except him who is from God; he has seen the Father.
JOHN|6|47|Truly, truly, I say to you, whoever believes has eternal life.
JOHN|6|48|I am the bread of life.
JOHN|6|49|Your fathers ate the manna in the wilderness, and they died.
JOHN|6|50|This is the bread that comes down from heaven, so that one may eat of it and not die.
JOHN|6|51|I am the living bread that came down from heaven. If anyone eats of this bread, he will live forever. And the bread that I will give for the life of the world is my flesh."
JOHN|6|52|The Jews then disputed among themselves, saying, "How can this man give us his flesh to eat?"
JOHN|6|53|So Jesus said to them, "Truly, truly, I say to you, unless you eat the flesh of the Son of Man and drink his blood, you have no life in you.
JOHN|6|54|Whoever feeds on my flesh and drinks my blood has eternal life, and I will raise him up on the last day.
JOHN|6|55|For my flesh is true food, and my blood is true drink.
JOHN|6|56|Whoever feeds on my flesh and drinks my blood abides in me, and I in him.
JOHN|6|57|As the living Father sent me, and I live because of the Father, so whoever feeds on me, he also will live because of me.
JOHN|6|58|This is the bread that came down from heaven, not as the fathers ate and died. Whoever feeds on this bread will live forever."
JOHN|6|59|Jesus said these things in the synagogue, as he taught at Capernaum.
JOHN|6|60|When many of his disciples heard it, they said, "This is a hard saying; who can listen to it?"
JOHN|6|61|But Jesus, knowing in himself that his disciples were grumbling about this, said to them, "Do you take offense at this?
JOHN|6|62|Then what if you were to see the Son of Man ascending to where he was before?
JOHN|6|63|It is the Spirit who gives life; the flesh is of no avail. The words that I have spoken to you are spirit and life.
JOHN|6|64|But there are some of you who do not believe." (For Jesus knew from the beginning who those were who did not believe, and who it was who would betray him.)
JOHN|6|65|And he said, "This is why I told you that no one can come to me unless it is granted him by the Father."
JOHN|6|66|After this many of his disciples turned back and no longer walked with him.
JOHN|6|67|So Jesus said to the Twelve, "Do you want to go away as well?"
JOHN|6|68|Simon Peter answered him, "Lord, to whom shall we go? You have the words of eternal life,
JOHN|6|69|and we have believed, and have come to know, that you are the Holy One of God."
JOHN|6|70|Jesus answered them, "Did I not choose you, the Twelve? And yet one of you is a devil."
JOHN|6|71|He spoke of Judas the son of Simon Iscariot, for he, one of the Twelve, was going to betray him.
JOHN|7|1|After this Jesus went about in Galilee. He would not go about in Judea, because the Jews were seeking to kill him.
JOHN|7|2|Now the Jews' Feast of Booths was at hand.
JOHN|7|3|So his brothers said to him, "Leave here and go to Judea, that your disciples also may see the works you are doing.
JOHN|7|4|For no one works in secret if he seeks to be known openly. If you do these things, show yourself to the world."
JOHN|7|5|For not even his brothers believed in him.
JOHN|7|6|Jesus said to them, "My time has not yet come, but your time is always here.
JOHN|7|7|The world cannot hate you, but it hates me because I testify about it that its works are evil.
JOHN|7|8|You go up to the feast. I am not going up to this feast, for my time has not yet fully come."
JOHN|7|9|After saying this, he remained in Galilee.
JOHN|7|10|But after his brothers had gone up to the feast, then he also went up, not publicly but in private.
JOHN|7|11|The Jews were looking for him at the feast, and saying, "Where is he?"
JOHN|7|12|And there was much muttering about him among the people. While some said, "He is a good man," others said, "No, he is leading the people astray."
JOHN|7|13|Yet for fear of the Jews no one spoke openly of him.
JOHN|7|14|About the middle of the feast Jesus went up into the temple and began teaching.
JOHN|7|15|The Jews therefore marveled, saying, "How is it that this man has learning, when he has never studied?"
JOHN|7|16|So Jesus answered them, "My teaching is not mine, but his who sent me.
JOHN|7|17|If anyone's will is to do God's will, he will know whether the teaching is from God or whether I am speaking on my own authority.
JOHN|7|18|The one who speaks on his own authority seeks his own glory, but the one who seeks the glory of him who sent him is true, and in him there is no falsehood.
JOHN|7|19|Has not Moses given you the law? Yet none of you keeps the law. Why do you seek to kill me?"
JOHN|7|20|The crowd answered, "You have a demon! Who is seeking to kill you?"
JOHN|7|21|Jesus answered them, "I did one deed, and you all marvel at it.
JOHN|7|22|Moses gave you circumcision (not that it is from Moses, but from the fathers), and you circumcise a man on the Sabbath.
JOHN|7|23|If on the Sabbath a man receives circumcision, so that the law of Moses may not be broken, are you angry with me because on the Sabbath I made a man's whole body well?
JOHN|7|24|Do not judge by appearances, but judge with right judgment."
JOHN|7|25|Some of the people of Jerusalem therefore said, "Is not this the man whom they seek to kill?
JOHN|7|26|And here he is, speaking openly, and they say nothing to him! Can it be that the authorities really know that this is the Christ?
JOHN|7|27|But we know where this man comes from, and when the Christ appears, no one will know where he comes from."
JOHN|7|28|So Jesus proclaimed, as he taught in the temple, "You know me, and you know where I come from? But I have not come of my own accord. He who sent me is true, and him you do not know.
JOHN|7|29|I know him, for I come from him, and he sent me."
JOHN|7|30|So they were seeking to arrest him, but no one laid a hand on him, because his hour had not yet come.
JOHN|7|31|Yet many of the people believed in him. They said, "When the Christ appears, will he do more signs than this man has done?"
JOHN|7|32|The Pharisees heard the crowd muttering these things about him, and the chief priests and Pharisees sent officers to arrest him.
JOHN|7|33|Jesus then said, "I will be with you a little longer, and then I am going to him who sent me.
JOHN|7|34|You will seek me and you will not find me. Where I am you cannot come."
JOHN|7|35|The Jews said to one another, "Where does this man intend to go that we will not find him? Does he intend to go to the Dispersion among the Greeks and teach the Greeks?
JOHN|7|36|What does he mean by saying, 'You will seek me and you will not find me,' and, 'Where I am you cannot come'?"
JOHN|7|37|On the last day of the feast, the great day, Jesus stood up and cried out, "If anyone thirsts, let him come to me and drink.
JOHN|7|38|Whoever believes in me, as the Scripture has said, 'Out of his heart will flow rivers of living water.'"
JOHN|7|39|Now this he said about the Spirit, whom those who believed in him were to receive, for as yet the Spirit had not been given, because Jesus was not yet glorified.
JOHN|7|40|When they heard these words, some of the people said, "This really is the Prophet."
JOHN|7|41|Others said, "This is the Christ." But some said, "Is the Christ to come from Galilee?
JOHN|7|42|Has not the Scripture said that the Christ comes from the offspring of David, and comes from Bethlehem, the village where David was?"
JOHN|7|43|So there was a division among the people over him.
JOHN|7|44|Some of them wanted to arrest him, but no one laid hands on him.
JOHN|7|45|The officers then came to the chief priests and Pharisees, who said to them, "Why did you not bring him?"
JOHN|7|46|The officers answered, "No one ever spoke like this man!"
JOHN|7|47|The Pharisees answered them, "Have you also been deceived?
JOHN|7|48|Have any of the authorities or the Pharisees believed in him?
JOHN|7|49|But this crowd that does not know the law is accursed."
JOHN|7|50|Nicodemus, who had gone to him before, and who was one of them, said to them,
JOHN|7|51|"Does our law judge a man without first giving him a hearing and learning what he does?"
JOHN|7|52|They replied, "Are you from Galilee too? Search and see that no prophet arises from Galilee." [THE EARLIEST MANUSCRIPTS DO NOT INCLUDE JOHN 7:53-8:11]
JOHN|7|53|[[They went each to his own house,
JOHN|8|1|but Jesus went to the Mount of Olives.
JOHN|8|2|Early in the morning he came again to the temple. All the people came to him, and he sat down and taught them.
JOHN|8|3|The scribes and the Pharisees brought a woman who had been caught in adultery, and placing her in the midst
JOHN|8|4|they said to him, "Teacher, this woman has been caught in the act of adultery.
JOHN|8|5|Now in the Law Moses commanded us to stone such women. So what do you say?"
JOHN|8|6|This they said to test him, that they might have some charge to bring against him. Jesus bent down and wrote with his finger on the ground.
JOHN|8|7|And as they continued to ask him, he stood up and said to them, "Let him who is without sin among you be the first to throw a stone at her."
JOHN|8|8|And once more he bent down and wrote on the ground.
JOHN|8|9|But when they heard it, they went away one by one, beginning with the older ones, and Jesus was left alone with the woman standing before him.
JOHN|8|10|Jesus stood up and said to her, "Woman, where are they? Has no one condemned you?"
JOHN|8|11|She said, "No one, Lord." And Jesus said, "Neither do I condemn you; go, and from now on sin no more."]]
JOHN|8|12|Again Jesus spoke to them, saying, "I am the light of the world. Whoever follows me will not walk in darkness, but will have the light of life."
JOHN|8|13|So the Pharisees said to him, "You are bearing witness about yourself; your testimony is not true."
JOHN|8|14|Jesus answered, "Even if I do bear witness about myself, my testimony is true, for I know where I came from and where I am going, but you do not know where I come from or where I am going.
JOHN|8|15|You judge according to the flesh; I judge no one.
JOHN|8|16|Yet even if I do judge, my judgment is true, for it is not I alone who judge, but I and the Father who sent me.
JOHN|8|17|In your Law it is written that the testimony of two men is true.
JOHN|8|18|I am the one who bears witness about myself, and the Father who sent me bears witness about me."
JOHN|8|19|They said to him therefore, "Where is your Father?" Jesus answered, "You know neither me nor my Father. If you knew me, you would know my Father also."
JOHN|8|20|These words he spoke in the treasury, as he taught in the temple; but no one arrested him, because his hour had not yet come.
JOHN|8|21|So he said to them again, "I am going away, and you will seek me, and you will die in your sin. Where I am going, you cannot come."
JOHN|8|22|So the Jews said, "Will he kill himself, since he says, 'Where I am going, you cannot come'?"
JOHN|8|23|He said to them, "You are from below; I am from above. You are of this world; I am not of this world.
JOHN|8|24|I told you that you would die in your sins, for unless you believe that I am he you will die in your sins."
JOHN|8|25|So they said to him, "Who are you?" Jesus said to them, "Just what I have been telling you from the beginning.
JOHN|8|26|I have much to say about you and much to judge, but he who sent me is true, and I declare to the world what I have heard from him."
JOHN|8|27|They did not understand that he had been speaking to them about the Father.
JOHN|8|28|So Jesus said to them, "When you have lifted up the Son of Man, then you will know that I am he, and that I do nothing on my own authority, but speak just as the Father taught me.
JOHN|8|29|And he who sent me is with me. He has not left me alone, for I always do the things that are pleasing to him."
JOHN|8|30|As he was saying these things, many believed in him.
JOHN|8|31|So Jesus said to the Jews who had believed in him, "If you abide in my word, you are truly my disciples,
JOHN|8|32|and you will know the truth, and the truth will set you free."
JOHN|8|33|They answered him, "We are offspring of Abraham and have never been enslaved to anyone. How is it that you say, 'You will become free'?"
JOHN|8|34|Jesus answered them, "Truly, truly, I say to you, everyone who commits sin is a slave to sin.
JOHN|8|35|The slave does not remain in the house forever; the son remains forever.
JOHN|8|36|So if the Son sets you free, you will be free indeed.
JOHN|8|37|I know that you are offspring of Abraham; yet you seek to kill me because my word finds no place in you.
JOHN|8|38|I speak of what I have seen with my Father, and you do what you have heard from your father."
JOHN|8|39|They answered him, "Abraham is our father." Jesus said to them, "If you were Abraham's children, you would be doing what Abraham did,
JOHN|8|40|but now you seek to kill me, a man who has told you the truth that I heard from God. This is not what Abraham did.
JOHN|8|41|You are doing what your father did." They said to him, "We were not born of sexual immorality. We have one Father- even God."
JOHN|8|42|Jesus said to them, "If God were your Father, you would love me, for I came from God and I am here. I came not of my own accord, but he sent me.
JOHN|8|43|Why do you not understand what I say? It is because you cannot bear to hear my word.
JOHN|8|44|You are of your father the devil, and your will is to do your father's desires. He was a murderer from the beginning, and has nothing to do with the truth, because there is no truth in him. When he lies, he speaks out of his own character, for he is a liar and the father of lies.
JOHN|8|45|But because I tell the truth, you do not believe me.
JOHN|8|46|Which one of you convicts me of sin? If I tell the truth, why do you not believe me?
JOHN|8|47|Whoever is of God hears the words of God. The reason why you do not hear them is that you are not of God."
JOHN|8|48|The Jews answered him, "Are we not right in saying that you are a Samaritan and have a demon?"
JOHN|8|49|Jesus answered, "I do not have a demon, but I honor my Father, and you dishonor me.
JOHN|8|50|Yet I do not seek my own glory; there is One who seeks it, and he is the judge.
JOHN|8|51|Truly, truly, I say to you, if anyone keeps my word, he will never see death."
JOHN|8|52|The Jews said to him, "Now we know that you have a demon! Abraham died, as did the prophets, yet you say, 'If anyone keeps my word, he will never taste death.'
JOHN|8|53|Are you greater than our father Abraham, who died? And the prophets died! Who do you make yourself out to be?"
JOHN|8|54|Jesus answered, "If I glorify myself, my glory is nothing. It is my Father who glorifies me, of whom you say, 'He is our God.'
JOHN|8|55|But you have not known him. I know him. If I were to say that I do not know him, I would be a liar like you, but I do know him and I keep his word.
JOHN|8|56|Your father Abraham rejoiced that he would see my day. He saw it and was glad."
JOHN|8|57|So the Jews said to him, "You are not yet fifty years old, and have you seen Abraham?"
JOHN|8|58|Jesus said to them, "Truly, truly, I say to you, before Abraham was, I am."
JOHN|8|59|So they picked up stones to throw at him, but Jesus hid himself and went out of the temple.
JOHN|9|1|As he passed by, he saw a man blind from birth.
JOHN|9|2|And his disciples asked him, "Rabbi, who sinned, this man or his parents, that he was born blind?"
JOHN|9|3|Jesus answered, "It was not that this man sinned, or his parents, but that the works of God might be displayed in him.
JOHN|9|4|We must work the works of him who sent me while it is day; night is coming, when no one can work.
JOHN|9|5|As long as I am in the world, I am the light of the world."
JOHN|9|6|Having said these things, he spat on the ground and made mud with the saliva. Then he anointed the man's eyes with the mud
JOHN|9|7|and said to him, "Go, wash in the pool of Siloam" (which means Sent). So he went and washed and came back seeing.
JOHN|9|8|The neighbors and those who had seen him before as a beggar were saying, "Is this not the man who used to sit and beg?"
JOHN|9|9|Some said, "It is he." Others said, "No, but he is like him." He kept saying, "I am the man."
JOHN|9|10|So they said to him, "Then how were your eyes opened?"
JOHN|9|11|He answered, "The man called Jesus made mud and anointed my eyes and said to me, 'Go to Siloam and wash.' So I went and washed and received my sight."
JOHN|9|12|They said to him, "Where is he?" He said, "I do not know."
JOHN|9|13|They brought to the Pharisees the man who had formerly been blind.
JOHN|9|14|Now it was a Sabbath day when Jesus made the mud and opened his eyes.
JOHN|9|15|So the Pharisees again asked him how he had received his sight. And he said to them, "He put mud on my eyes, and I washed, and I see."
JOHN|9|16|Some of the Pharisees said, "This man is not from God, for he does not keep the Sabbath." But others said, "How can a man who is a sinner do such signs?" And there was a division among them.
JOHN|9|17|So they said again to the blind man, "What do you say about him, since he has opened your eyes?" He said, "He is a prophet."
JOHN|9|18|The Jews did not believe that he had been blind and had received his sight, until they called the parents of the man who had received his sight
JOHN|9|19|and asked them, "Is this your son, who you say was born blind? How then does he now see?"
JOHN|9|20|His parents answered, "We know that this is our son and that he was born blind.
JOHN|9|21|But how he now sees we do not know, nor do we know who opened his eyes. Ask him; he is of age. He will speak for himself."
JOHN|9|22|(His parents said these things because they feared the Jews, for the Jews had already agreed that if anyone should confess Jesus to be Christ, he was to be put out of the synagogue.)
JOHN|9|23|Therefore his parents said, "He is of age; ask him."
JOHN|9|24|So for the second time they called the man who had been blind and said to him, "Give glory to God. We know that this man is a sinner."
JOHN|9|25|He answered, "Whether he is a sinner I do not know. One thing I do know, that though I was blind, now I see."
JOHN|9|26|They said to him, "What did he do to you? How did he open your eyes?"
JOHN|9|27|He answered them, "I have told you already, and you would not listen. Why do you want to hear it again? Do you also want to become his disciples?"
JOHN|9|28|And they reviled him, saying, "You are his disciple, but we are disciples of Moses.
JOHN|9|29|We know that God has spoken to Moses, but as for this man, we do not know where he comes from."
JOHN|9|30|The man answered, "Why, this is an amazing thing! You do not know where he comes from, and yet he opened my eyes.
JOHN|9|31|We know that God does not listen to sinners, but if anyone is a worshiper of God and does his will, God listens to him.
JOHN|9|32|Never since the world began has it been heard that anyone opened the eyes of a man born blind.
JOHN|9|33|If this man were not from God, he could do nothing."
JOHN|9|34|They answered him, "You were born in utter sin, and would you teach us?" And they cast him out.
JOHN|9|35|Jesus heard that they had cast him out, and having found him he said, "Do you believe in the Son of Man?"
JOHN|9|36|He answered, "And who is he, sir, that I may believe in him?"
JOHN|9|37|Jesus said to him, "You have seen him, and it is he who is speaking to you."
JOHN|9|38|He said, "Lord, I believe," and he worshiped him.
JOHN|9|39|Jesus said, "For judgment I came into this world, that those who do not see may see, and those who see may become blind."
JOHN|9|40|Some of the Pharisees near him heard these things, and said to him, "Are we also blind?"
JOHN|9|41|Jesus said to them, "If you were blind, you would have no guilt; but now that you say, 'We see,' your guilt remains.
JOHN|10|1|"Truly, truly, I say to you, he who does not enter the sheepfold by the door but climbs in by another way, that man is a thief and a robber.
JOHN|10|2|But he who enters by the door is the shepherd of the sheep.
JOHN|10|3|To him the gatekeeper opens. The sheep hear his voice, and he calls his own sheep by name and leads them out.
JOHN|10|4|When he has brought out all his own, he goes before them, and the sheep follow him, for they know his voice.
JOHN|10|5|A stranger they will not follow, but they will flee from him, for they do not know the voice of strangers."
JOHN|10|6|This figure of speech Jesus used with them, but they did not understand what he was saying to them.
JOHN|10|7|So Jesus again said to them, "Truly, truly, I say to you, I am the door of the sheep.
JOHN|10|8|All who came before me are thieves and robbers, but the sheep did not listen to them.
JOHN|10|9|I am the door. If anyone enters by me, he will be saved and will go in and out and find pasture.
JOHN|10|10|The thief comes only to steal and kill and destroy. I came that they may have life and have it abundantly.
JOHN|10|11|I am the good shepherd. The good shepherd lays down his life for the sheep.
JOHN|10|12|He who is a hired hand and not a shepherd, who does not own the sheep, sees the wolf coming and leaves the sheep and flees, and the wolf snatches them and scatters them.
JOHN|10|13|He flees because he is a hired hand and cares nothing for the sheep.
JOHN|10|14|I am the good shepherd. I know my own and my own know me,
JOHN|10|15|just as the Father knows me and I know the Father; and I lay down my life for the sheep.
JOHN|10|16|And I have other sheep that are not of this fold. I must bring them also, and they will listen to my voice. So there will be one flock, one shepherd.
JOHN|10|17|For this reason the Father loves me, because I lay down my life that I may take it up again.
JOHN|10|18|No one takes it from me, but I lay it down of my own accord. I have authority to lay it down, and I have authority to take it up again. This charge I have received from my Father."
JOHN|10|19|There was again a division among the Jews because of these words.
JOHN|10|20|Many of them said, "He has a demon, and is insane; why listen to him?"
JOHN|10|21|Others said, "These are not the words of one who is oppressed by a demon. Can a demon open the eyes of the blind?"
JOHN|10|22|At that time the Feast of Dedication took place at Jerusalem. It was winter,
JOHN|10|23|and Jesus was walking in the temple, in the colonnade of Solomon.
JOHN|10|24|So the Jews gathered around him and said to him, "How long will you keep us in suspense? If you are the Christ, tell us plainly."
JOHN|10|25|Jesus answered them, "I told you, and you do not believe. The works that I do in my Father's name bear witness about me,
JOHN|10|26|but you do not believe because you are not part of my flock.
JOHN|10|27|My sheep hear my voice, and I know them, and they follow me.
JOHN|10|28|I give them eternal life, and they will never perish, and no one will snatch them out of my hand.
JOHN|10|29|My Father, who has given them to me, is greater than all, and no one is able to snatch them out of the Father's hand.
JOHN|10|30|I and the Father are one."
JOHN|10|31|The Jews picked up stones again to stone him.
JOHN|10|32|Jesus answered them, "I have shown you many good works from the Father; for which of them are you going to stone me?"
JOHN|10|33|The Jews answered him, "It is not for a good work that we are going to stone you but for blasphemy, because you, being a man, make yourself God."
JOHN|10|34|Jesus answered them, "Is it not written in your Law, 'I said, you are gods'?
JOHN|10|35|If he called them gods to whom the word of God came- and Scripture cannot be broken-
JOHN|10|36|do you say of him whom the Father consecrated and sent into the world, 'You are blaspheming,' because I said, 'I am the Son of God'?
JOHN|10|37|If I am not doing the works of my Father, then do not believe me;
JOHN|10|38|but if I do them, even though you do not believe me, believe the works, that you may know and understand that the Father is in me and I am in the Father."
JOHN|10|39|Again they sought to arrest him, but he escaped from their hands.
JOHN|10|40|He went away again across the Jordan to the place where John had been baptizing at first, and there he remained.
JOHN|10|41|And many came to him. And they said, "John did no sign, but everything that John said about this man was true."
JOHN|10|42|And many believed in him there.
JOHN|11|1|Now a certain man was ill, Lazarus of Bethany, the village of Mary and her sister Martha.
JOHN|11|2|It was Mary who anointed the Lord with ointment and wiped his feet with her hair, whose brother Lazarus was ill.
JOHN|11|3|So the sisters sent to him, saying, "Lord, he whom you love is ill."
JOHN|11|4|But when Jesus heard it he said, "This illness does not lead to death. It is for the glory of God, so that the Son of God may be glorified through it."
JOHN|11|5|Now Jesus loved Martha and her sister and Lazarus.
JOHN|11|6|So, when he heard that Lazarus was ill, he stayed two days longer in the place where he was.
JOHN|11|7|Then after this he said to the disciples, "Let us go to Judea again."
JOHN|11|8|The disciples said to him, "Rabbi, the Jews were just now seeking to stone you, and are you going there again?"
JOHN|11|9|Jesus answered, "Are there not twelve hours in the day? If anyone walks in the day, he does not stumble, because he sees the light of this world.
JOHN|11|10|But if anyone walks in the night, he stumbles, because the light is not in him."
JOHN|11|11|After saying these things, he said to them, "Our friend Lazarus has fallen asleep, but I go to awaken him."
JOHN|11|12|The disciples said to him, "Lord, if he has fallen asleep, he will recover."
JOHN|11|13|Now Jesus had spoken of his death, but they thought that he meant taking rest in sleep.
JOHN|11|14|Then Jesus told them plainly, "Lazarus has died,
JOHN|11|15|and for your sake I am glad that I was not there, so that you may believe. But let us go to him."
JOHN|11|16|So Thomas, called the Twin, said to his fellow disciples, "Let us also go, that we may die with him."
JOHN|11|17|Now when Jesus came, he found that Lazarus had already been in the tomb four days.
JOHN|11|18|Bethany was near Jerusalem, about two miles off,
JOHN|11|19|and many of the Jews had come to Martha and Mary to console them concerning their brother.
JOHN|11|20|So when Martha heard that Jesus was coming, she went and met him, but Mary remained seated in the house.
JOHN|11|21|Martha said to Jesus, "Lord, if you had been here, my brother would not have died.
JOHN|11|22|But even now I know that whatever you ask from God, God will give you."
JOHN|11|23|Jesus said to her, "Your brother will rise again."
JOHN|11|24|Martha said to him, "I know that he will rise again in the resurrection on the last day."
JOHN|11|25|Jesus said to her, "I am the resurrection and the life. Whoever believes in me, though he die, yet shall he live,
JOHN|11|26|and everyone who lives and believes in me shall never die. Do you believe this?"
JOHN|11|27|She said to him, "Yes, Lord; I believe that you are the Christ, the Son of God, who is coming into the world."
JOHN|11|28|When she had said this, she went and called her sister Mary, saying in private, "The Teacher is here and is calling for you."
JOHN|11|29|And when she heard it, she rose quickly and went to him.
JOHN|11|30|Now Jesus had not yet come into the village, but was still in the place where Martha had met him.
JOHN|11|31|When the Jews who were with her in the house, consoling her, saw Mary rise quickly and go out, they followed her, supposing that she was going to the tomb to weep there.
JOHN|11|32|Now when Mary came to where Jesus was and saw him, she fell at his feet, saying to him, "Lord, if you had been here, my brother would not have died."
JOHN|11|33|When Jesus saw her weeping, and the Jews who had come with her also weeping, he was deeply moved in his spirit and greatly troubled.
JOHN|11|34|And he said, "Where have you laid him?" They said to him, "Lord, come and see."
JOHN|11|35|Jesus wept.
JOHN|11|36|So the Jews said, "See how he loved him!"
JOHN|11|37|But some of them said, "Could not he who opened the eyes of the blind man also have kept this man from dying?"
JOHN|11|38|Then Jesus, deeply moved again, came to the tomb. It was a cave, and a stone lay against it.
JOHN|11|39|Jesus said, "Take away the stone." Martha, the sister of the dead man, said to him, "Lord, by this time there will be an odor, for he has been dead four days."
JOHN|11|40|Jesus said to her, "Did I not tell you that if you believed you would see the glory of God?"
JOHN|11|41|So they took away the stone. And Jesus lifted up his eyes and said, "Father, I thank you that you have heard me.
JOHN|11|42|I knew that you always hear me, but I said this on account of the people standing around, that they may believe that you sent me."
JOHN|11|43|When he had said these things, he cried out with a loud voice, "Lazarus, come out."
JOHN|11|44|The man who had died came out, his hands and feet bound with linen strips, and his face wrapped with a cloth. Jesus said to them, "Unbind him, and let him go."
JOHN|11|45|Many of the Jews therefore, who had come with Mary and had seen what he did, believed in him,
JOHN|11|46|but some of them went to the Pharisees and told them what Jesus had done.
JOHN|11|47|So the chief priests and the Pharisees gathered the Council and said, "What are we to do? For this man performs many signs.
JOHN|11|48|If we let him go on like this, everyone will believe in him, and the Romans will come and take away both our place and our nation."
JOHN|11|49|But one of them, Caiaphas, who was high priest that year, said to them, "You know nothing at all.
JOHN|11|50|Nor do you understand that it is better for you that one man should die for the people, not that the whole nation should perish."
JOHN|11|51|He did not say this of his own accord, but being high priest that year he prophesied that Jesus would die for the nation,
JOHN|11|52|and not for the nation only, but also to gather into one the children of God who are scattered abroad.
JOHN|11|53|So from that day on they made plans to put him to death.
JOHN|11|54|Jesus therefore no longer walked openly among the Jews, but went from there to the region near the wilderness, to a town called Ephraim, and there he stayed with the disciples.
JOHN|11|55|Now the Passover of the Jews was at hand, and many went up from the country to Jerusalem before the Passover to purify themselves.
JOHN|11|56|They were looking for Jesus and saying to one another as they stood in the temple, "What do you think? That he will not come to the feast at all?"
JOHN|11|57|Now the chief priests and the Pharisees had given orders that if anyone knew where he was, he should let them know, so that they might arrest him.
JOHN|12|1|Six days before the Passover, Jesus therefore came to Bethany, where Lazarus was, whom Jesus had raised from the dead.
JOHN|12|2|So they gave a dinner for him there. Martha served, and Lazarus was one of those reclining with him at the table.
JOHN|12|3|Mary therefore took a pound of expensive ointment made from pure nard, and anointed the feet of Jesus and wiped his feet with her hair. The house was filled with the fragrance of the perfume.
JOHN|12|4|But Judas Iscariot, one of his disciples (he who was about to betray him), said,
JOHN|12|5|"Why was this ointment not sold for three hundred denarii and given to the poor?"
JOHN|12|6|He said this, not because he cared about the poor, but because he was a thief, and having charge of the moneybag he used to help himself to what was put into it.
JOHN|12|7|Jesus said, "Leave her alone, so that she may keep it for the day of my burial.
JOHN|12|8|The poor you always have with you, but you do not always have me."
JOHN|12|9|When the large crowd of the Jews learned that Jesus was there, they came, not only on account of him but also to see Lazarus, whom he had raised from the dead.
JOHN|12|10|So the chief priests made plans to put Lazarus to death as well,
JOHN|12|11|because on account of him many of the Jews were going away and believing in Jesus.
JOHN|12|12|The next day the large crowd that had come to the feast heard that Jesus was coming to Jerusalem.
JOHN|12|13|So they took branches of palm trees and went out to meet him, crying out, "Hosanna! Blessed is he who comes in the name of the Lord, even the King of Israel!"
JOHN|12|14|And Jesus found a young donkey and sat on it, just as it is written,
JOHN|12|15|"Fear not, daughter of Zion; behold, your king is coming, sitting on a donkey's colt!"
JOHN|12|16|His disciples did not understand these things at first, but when Jesus was glorified, then they remembered that these things had been written about him and had been done to him.
JOHN|12|17|The crowd that had been with him when he called Lazarus out of the tomb and raised him from the dead continued to bear witness.
JOHN|12|18|The reason why the crowd went to meet him was that they heard he had done this sign.
JOHN|12|19|So the Pharisees said to one another, "You see that you are gaining nothing. Look, the world has gone after him."
JOHN|12|20|Now among those who went up to worship at the feast were some Greeks.
JOHN|12|21|So these came to Philip, who was from Bethsaida in Galilee, and asked him, "Sir, we wish to see Jesus."
JOHN|12|22|Philip went and told Andrew; Andrew and Philip went and told Jesus.
JOHN|12|23|And Jesus answered them, "The hour has come for the Son of Man to be glorified.
JOHN|12|24|Truly, truly, I say to you, unless a grain of wheat falls into the earth and dies, it remains alone; but if it dies, it bears much fruit.
JOHN|12|25|Whoever loves his life loses it, and whoever hates his life in this world will keep it for eternal life.
JOHN|12|26|If anyone serves me, he must follow me; and where I am, there will my servant be also. If anyone serves me, the Father will honor him.
JOHN|12|27|"Now is my soul troubled. And what shall I say? 'Father, save me from this hour'? But for this purpose I have come to this hour.
JOHN|12|28|Father, glorify your name." Then a voice came from heaven: "I have glorified it, and I will glorify it again."
JOHN|12|29|The crowd that stood there and heard it said that it had thundered. Others said, "An angel has spoken to him."
JOHN|12|30|Jesus answered, "This voice has come for your sake, not mine.
JOHN|12|31|Now is the judgment of this world; now will the ruler of this world be cast out.
JOHN|12|32|And I, when I am lifted up from the earth, will draw all people to myself."
JOHN|12|33|He said this to show by what kind of death he was going to die.
JOHN|12|34|So the crowd answered him, "We have heard from the Law that the Christ remains forever. How can you say that the Son of Man must be lifted up? Who is this Son of Man?"
JOHN|12|35|So Jesus said to them, "The light is among you for a little while longer. Walk while you have the light, lest darkness overtake you. The one who walks in the darkness does not know where he is going.
JOHN|12|36|While you have the light, believe in the light, that you may become sons of light." When Jesus had said these things, he departed and hid himself from them.
JOHN|12|37|Though he had done so many signs before them, they still did not believe in him,
JOHN|12|38|so that the word spoken by the prophet Isaiah might be fulfilled: "Lord, who has believed what he heard from us, and to whom has the arm of the Lord been revealed?"
JOHN|12|39|Therefore they could not believe. For again Isaiah said,
JOHN|12|40|"He has blinded their eyes and hardened their heart, lest they see with their eyes, and understand with their heart, and turn, and I would heal them."
JOHN|12|41|Isaiah said these things because he saw his glory and spoke of him.
JOHN|12|42|Nevertheless, many even of the authorities believed in him, but for fear of the Pharisees they did not confess it, so that they would not be put out of the synagogue;
JOHN|12|43|for they loved the glory that comes from man more than the glory that comes from God.
JOHN|12|44|And Jesus cried out and said, "Whoever believes in me, believes not in me but in him who sent me.
JOHN|12|45|And whoever sees me sees him who sent me.
JOHN|12|46|I have come into the world as light, so that whoever believes in me may not remain in darkness.
JOHN|12|47|If anyone hears my words and does not keep them, I do not judge him; for I did not come to judge the world but to save the world.
JOHN|12|48|The one who rejects me and does not receive my words has a judge; the word that I have spoken will judge him on the last day.
JOHN|12|49|For I have not spoken on my own authority, but the Father who sent me has himself given me a commandment- what to say and what to speak.
JOHN|12|50|And I know that his commandment is eternal life. What I say, therefore, I say as the Father has told me."
JOHN|13|1|Now before the Feast of the Passover, when Jesus knew that his hour had come to depart out of this world to the Father, having loved his own who were in the world, he loved them to the end.
JOHN|13|2|During supper, when the devil had already put it into the heart of Judas Iscariot, Simon's son, to betray him,
JOHN|13|3|Jesus, knowing that the Father had given all things into his hands, and that he had come from God and was going back to God,
JOHN|13|4|rose from supper. He laid aside his outer garments, and taking a towel, tied it around his waist.
JOHN|13|5|Then he poured water into a basin and began to wash the disciples' feet and to wipe them with the towel that was wrapped around him.
JOHN|13|6|He came to Simon Peter, who said to him, "Lord, do you wash my feet?"
JOHN|13|7|Jesus answered him, "What I am doing you do not understand now, but afterward you will understand."
JOHN|13|8|Peter said to him, "You shall never wash my feet." Jesus answered him, "If I do not wash you, you have no share with me."
JOHN|13|9|Simon Peter said to him, "Lord, not my feet only but also my hands and my head!"
JOHN|13|10|Jesus said to him, "The one who has bathed does not need to wash, except for his feet, but is completely clean. And you are clean, but not every one of you."
JOHN|13|11|For he knew who was to betray him; that was why he said, "Not all of you are clean."
JOHN|13|12|When he had washed their feet and put on his outer garments and resumed his place, he said to them, "Do you understand what I have done to you?
JOHN|13|13|You call me Teacher and Lord, and you are right, for so I am.
JOHN|13|14|If I then, your Lord and Teacher, have washed your feet, you also ought to wash one another's feet.
JOHN|13|15|For I have given you an example, that you also should do just as I have done to you.
JOHN|13|16|Truly, truly, I say to you, a servant is not greater than his master, nor is a messenger greater than the one who sent him.
JOHN|13|17|If you know these things, blessed are you if you do them.
JOHN|13|18|I am not speaking of all of you; I know whom I have chosen. But the Scripture will be fulfilled, 'He who ate my bread has lifted his heel against me.'
JOHN|13|19|I am telling you this now, before it takes place, that when it does take place you may believe that I am he.
JOHN|13|20|Truly, truly, I say to you, whoever receives the one I send receives me, and whoever receives me receives the one who sent me."
JOHN|13|21|After saying these things, Jesus was troubled in his spirit, and testified, "Truly, truly, I say to you, one of you will betray me."
JOHN|13|22|The disciples looked at one another, uncertain of whom he spoke.
JOHN|13|23|One of his disciples, whom Jesus loved, was reclining at table close to Jesus,
JOHN|13|24|so Simon Peter motioned to him to ask Jesus of whom he was speaking.
JOHN|13|25|So that disciple, leaning back against Jesus, said to him, "Lord, who is it?"
JOHN|13|26|Jesus answered, "It is he to whom I will give this morsel of bread when I have dipped it." So when he had dipped the morsel, he gave it to Judas, the son of Simon Iscariot.
JOHN|13|27|Then after he had taken the morsel, Satan entered into him. Jesus said to him, "What you are going to do, do quickly."
JOHN|13|28|Now no one at the table knew why he said this to him.
JOHN|13|29|Some thought that, because Judas had the moneybag, Jesus was telling him, "Buy what we need for the feast," or that he should give something to the poor.
JOHN|13|30|So, after receiving the morsel of bread, he immediately went out. And it was night.
JOHN|13|31|When he had gone out, Jesus said, "Now is the Son of Man glorified, and God is glorified in him.
JOHN|13|32|If God is glorified in him, God will also glorify him in himself, and glorify him at once.
JOHN|13|33|Little children, yet a little while I am with you. You will seek me, and just as I said to the Jews, so now I also say to you, 'Where I am going you cannot come.'
JOHN|13|34|A new commandment I give to you, that you love one another: just as I have loved you, you also are to love one another.
JOHN|13|35|By this all people will know that you are my disciples, if you have love for one another."
JOHN|13|36|Simon Peter said to him, "Lord, where are you going?" Jesus answered him, "Where I am going you cannot follow me now, but you will follow afterward."
JOHN|13|37|Peter said to him, "Lord, why can I not follow you now? I will lay down my life for you."
JOHN|13|38|Jesus answered, "Will you lay down your life for me? Truly, truly, I say to you, the rooster will not crow till you have denied me three times.
JOHN|14|1|"Let not your hearts be troubled. Believe in God; believe also in me.
JOHN|14|2|In my Father's house are many rooms. If it were not so, would I have told you that I go to prepare a place for you?
JOHN|14|3|And if I go and prepare a place for you, I will come again and will take you to myself, that where I am you may be also.
JOHN|14|4|And you know the way to where I am going."
JOHN|14|5|Thomas said to him, "Lord, we do not know where you are going. How can we know the way?"
JOHN|14|6|Jesus said to him, "I am the way, and the truth, and the life. No one comes to the Father except through me.
JOHN|14|7|If you had known me, you would have known my Father also. From now on you do know him and have seen him."
JOHN|14|8|Philip said to him, "Lord, show us the Father, and it is enough for us."
JOHN|14|9|Jesus said to him, "Have I been with you so long, and you still do not know me, Philip? Whoever has seen me has seen the Father. How can you say, 'Show us the Father'?
JOHN|14|10|Do you not believe that I am in the Father and the Father is in me? The words that I say to you I do not speak on my own authority, but the Father who dwells in me does his works.
JOHN|14|11|Believe me that I am in the Father and the Father is in me, or else believe on account of the works themselves.
JOHN|14|12|"Truly, truly, I say to you, whoever believes in me will also do the works that I do; and greater works than these will he do, because I am going to the Father.
JOHN|14|13|Whatever you ask in my name, this I will do, that the Father may be glorified in the Son.
JOHN|14|14|If you ask me anything in my name, I will do it.
JOHN|14|15|"If you love me, you will keep my commandments.
JOHN|14|16|And I will ask the Father, and he will give you another Helper, to be with you forever,
JOHN|14|17|even the Spirit of truth, whom the world cannot receive, because it neither sees him nor knows him. You know him, for he dwells with you and will be in you.
JOHN|14|18|"I will not leave you as orphans; I will come to you.
JOHN|14|19|Yet a little while and the world will see me no more, but you will see me. Because I live, you also will live.
JOHN|14|20|In that day you will know that I am in my Father, and you in me, and I in you.
JOHN|14|21|Whoever has my commandments and keeps them, he it is who loves me. And he who loves me will be loved by my Father, and I will love him and manifest myself to him."
JOHN|14|22|Judas (not Iscariot) said to him, "Lord, how is it that you will manifest yourself to us, and not to the world?"
JOHN|14|23|Jesus answered him, "If anyone loves me, he will keep my word, and my Father will love him, and we will come to him and make our home with him.
JOHN|14|24|Whoever does not love me does not keep my words. And the word that you hear is not mine but the Father's who sent me.
JOHN|14|25|"These things I have spoken to you while I am still with you.
JOHN|14|26|But the Helper, the Holy Spirit, whom the Father will send in my name, he will teach you all things and bring to your remembrance all that I have said to you.
JOHN|14|27|Peace I leave with you; my peace I give to you. Not as the world gives do I give to you. Let not your hearts be troubled, neither let them be afraid.
JOHN|14|28|You heard me say to you, 'I am going away, and I will come to you.' If you loved me, you would have rejoiced, because I am going to the Father, for the Father is greater than I.
JOHN|14|29|And now I have told you before it takes place, so that when it does take place you may believe.
JOHN|14|30|I will no longer talk much with you, for the ruler of this world is coming. He has no claim on me,
JOHN|14|31|but I do as the Father has commanded me, so that the world may know that I love the Father. Rise, let us go from here.
JOHN|15|1|"I am the true vine, and my Father is the vinedresser.
JOHN|15|2|Every branch of mine that does not bear fruit he takes away, and every branch that does bear fruit he prunes, that it may bear more fruit.
JOHN|15|3|Already you are clean because of the word that I have spoken to you.
JOHN|15|4|Abide in me, and I in you. As the branch cannot bear fruit by itself, unless it abides in the vine, neither can you, unless you abide in me.
JOHN|15|5|I am the vine; you are the branches. Whoever abides in me and I in him, he it is that bears much fruit, for apart from me you can do nothing.
JOHN|15|6|If anyone does not abide in me he is thrown away like a branch and withers; and the branches are gathered, thrown into the fire, and burned.
JOHN|15|7|If you abide in me, and my words abide in you, ask whatever you wish, and it will be done for you.
JOHN|15|8|By this my Father is glorified, that you bear much fruit and so prove to be my disciples.
JOHN|15|9|As the Father has loved me, so have I loved you. Abide in my love.
JOHN|15|10|If you keep my commandments, you will abide in my love, just as I have kept my Father's commandments and abide in his love.
JOHN|15|11|These things I have spoken to you, that my joy may be in you, and that your joy may be full.
JOHN|15|12|"This is my commandment, that you love one another as I have loved you.
JOHN|15|13|Greater love has no one than this, that someone lays down his life for his friends.
JOHN|15|14|You are my friends if you do what I command you.
JOHN|15|15|No longer do I call you servants, for the servant does not know what his master is doing; but I have called you friends, for all that I have heard from my Father I have made known to you.
JOHN|15|16|You did not choose me, but I chose you and appointed you that you should go and bear fruit and that your fruit should abide, so that whatever you ask the Father in my name, he may give it to you.
JOHN|15|17|These things I command you, so that you will love one another.
JOHN|15|18|"If the world hates you, know that it has hated me before it hated you.
JOHN|15|19|If you were of the world, the world would love you as its own; but because you are not of the world, but I chose you out of the world, therefore the world hates you.
JOHN|15|20|Remember the word that I said to you: 'A servant is not greater than his master.' If they persecuted me, they will also persecute you. If they kept my word, they will also keep yours.
JOHN|15|21|But all these things they will do to you on account of my name, because they do not know him who sent me.
JOHN|15|22|If I had not come and spoken to them, they would not have been guilty of sin, but now they have no excuse for their sin.
JOHN|15|23|Whoever hates me hates my Father also.
JOHN|15|24|If I had not done among them the works that no one else did, they would not be guilty of sin, but now they have seen and hated both me and my Father.
JOHN|15|25|But the word that is written in their Law must be fulfilled: 'They hated me without a cause.'
JOHN|15|26|"But when the Helper comes, whom I will send to you from the Father, the Spirit of truth, who proceeds from the Father, he will bear witness about me.
JOHN|15|27|And you also will bear witness, because you have been with me from the beginning.
JOHN|16|1|"I have said all these things to you to keep you from falling away.
JOHN|16|2|They will put you out of the synagogues. Indeed, the hour is coming when whoever kills you will think he is offering service to God.
JOHN|16|3|And they will do these things because they have not known the Father, nor me.
JOHN|16|4|But I have said these things to you, that when their hour comes you may remember that I told them to you. "I did not say these things to you from the beginning, because I was with you.
JOHN|16|5|But now I am going to him who sent me, and none of you asks me, 'Where are you going?'
JOHN|16|6|But because I have said these things to you, sorrow has filled your heart.
JOHN|16|7|Nevertheless, I tell you the truth: it is to your advantage that I go away, for if I do not go away, the Helper will not come to you. But if I go, I will send him to you.
JOHN|16|8|And when he comes, he will convict the world concerning sin and righteousness and judgment:
JOHN|16|9|concerning sin, because they do not believe in me;
JOHN|16|10|concerning righteousness, because I go to the Father, and you will see me no longer;
JOHN|16|11|concerning judgment, because the ruler of this world is judged.
JOHN|16|12|"I still have many things to say to you, but you cannot bear them now.
JOHN|16|13|When the Spirit of truth comes, he will guide you into all the truth, for he will not speak on his own authority, but whatever he hears he will speak, and he will declare to you the things that are to come.
JOHN|16|14|He will glorify me, for he will take what is mine and declare it to you.
JOHN|16|15|All that the Father has is mine; therefore I said that he will take what is mine and declare it to you.
JOHN|16|16|"A little while, and you will see me no longer; and again a little while, and you will see me."
JOHN|16|17|So some of his disciples said to one another, "What is this that he says to us, 'A little while, and you will not see me, and again a little while, and you will see me'; and, 'because I am going to the Father'?"
JOHN|16|18|So they were saying, "What does he mean by 'a little while'? We do not know what he is talking about."
JOHN|16|19|Jesus knew that they wanted to ask him, so he said to them, "Is this what you are asking yourselves, what I meant by saying, 'A little while and you will not see me, and again a little while and you will see me'?
JOHN|16|20|Truly, truly, I say to you, you will weep and lament, but the world will rejoice. You will be sorrowful, but your sorrow will turn into joy.
JOHN|16|21|When a woman is giving birth, she has sorrow because her hour has come, but when she has delivered the baby, she no longer remembers the anguish, for joy that a human being has been born into the world.
JOHN|16|22|So also you have sorrow now, but I will see you again and your hearts will rejoice, and no one will take your joy from you.
JOHN|16|23|In that day you will ask nothing of me. Truly, truly, I say to you, whatever you ask of the Father in my name, he will give it to you.
JOHN|16|24|Until now you have asked nothing in my name. Ask, and you will receive, that your joy may be full.
JOHN|16|25|"I have said these things to you in figures of speech. The hour is coming when I will no longer speak to you in figures of speech but will tell you plainly about the Father.
JOHN|16|26|In that day you will ask in my name, and I do not say to you that I will ask the Father on your behalf;
JOHN|16|27|for the Father himself loves you, because you have loved me and have believed that I came from God.
JOHN|16|28|I came from the Father and have come into the world, and now I am leaving the world and going to the Father."
JOHN|16|29|His disciples said, "Ah, now you are speaking plainly and not using figurative speech!
JOHN|16|30|Now we know that you know all things and do not need anyone to question you; this is why we believe that you came from God."
JOHN|16|31|Jesus answered them, "Do you now believe?
JOHN|16|32|Behold, the hour is coming, indeed it has come, when you will be scattered, each to his own home, and will leave me alone. Yet I am not alone, for the Father is with me.
JOHN|16|33|I have said these things to you, that in me you may have peace. In the world you will have tribulation. But take heart; I have overcome the world."
JOHN|17|1|When Jesus had spoken these words, he lifted up his eyes to heaven, and said, "Father, the hour has come; glorify your Son that the Son may glorify you,
JOHN|17|2|since you have given him authority over all flesh, to give eternal life to all whom you have given him.
JOHN|17|3|And this is eternal life, that they know you the only true God, and Jesus Christ whom you have sent.
JOHN|17|4|I glorified you on earth, having accomplished the work that you gave me to do.
JOHN|17|5|And now, Father, glorify me in your own presence with the glory that I had with you before the world existed.
JOHN|17|6|"I have manifested your name to the people whom you gave me out of the world. Yours they were, and you gave them to me, and they have kept your word.
JOHN|17|7|Now they know that everything that you have given me is from you.
JOHN|17|8|For I have given them the words that you gave me, and they have received them and have come to know in truth that I came from you; and they have believed that you sent me.
JOHN|17|9|I am praying for them. I am not praying for the world but for those whom you have given me, for they are yours.
JOHN|17|10|All mine are yours, and yours are mine, and I am glorified in them.
JOHN|17|11|And I am no longer in the world, but they are in the world, and I am coming to you. Holy Father, keep them in your name, which you have given me, that they may be one, even as we are one.
JOHN|17|12|While I was with them, I kept them in your name, which you have given me. I have guarded them, and not one of them has been lost except the son of destruction, that the Scripture might be fulfilled.
JOHN|17|13|But now I am coming to you, and these things I speak in the world, that they may have my joy fulfilled in themselves.
JOHN|17|14|I have given them your word, and the world has hated them because they are not of the world, just as I am not of the world.
JOHN|17|15|I do not ask that you take them out of the world, but that you keep them from the evil one.
JOHN|17|16|They are not of the world, just as I am not of the world.
JOHN|17|17|Sanctify them in the truth; your word is truth.
JOHN|17|18|As you sent me into the world, so I have sent them into the world.
JOHN|17|19|And for their sake I consecrate myself, that they also may be sanctified in truth.
JOHN|17|20|"I do not ask for these only, but also for those who will believe in me through their word,
JOHN|17|21|that they may all be one, just as you, Father, are in me, and I in you, that they also may be in us, so that the world may believe that you have sent me.
JOHN|17|22|The glory that you have given me I have given to them, that they may be one even as we are one,
JOHN|17|23|I in them and you in me, that they may become perfectly one, so that the world may know that you sent me and loved them even as you loved me.
JOHN|17|24|Father, I desire that they also, whom you have given me, may be with me where I am, to see my glory that you have given me because you loved me before the foundation of the world.
JOHN|17|25|O righteous Father, even though the world does not know you, I know you, and these know that you have sent me.
JOHN|17|26|I made known to them your name, and I will continue to make it known, that the love with which you have loved me may be in them, and I in them."
JOHN|18|1|When Jesus had spoken these words, he went out with his disciples across the Kidron Valley, where there was a garden, which he and his disciples entered.
JOHN|18|2|Now Judas, who betrayed him, also knew the place, for Jesus often met there with his disciples.
JOHN|18|3|So Judas, having procured a band of soldiers and some officers from the chief priests and the Pharisees, went there with lanterns and torches and weapons.
JOHN|18|4|Then Jesus, knowing all that would happen to him, came forward and said to them, "Whom do you seek?"
JOHN|18|5|They answered him, "Jesus of Nazareth." Jesus said to them, "I am he." Judas, who betrayed him, was standing with them.
JOHN|18|6|When Jesus said to them, "I am he," they drew back and fell to the ground.
JOHN|18|7|So he asked them again, "Whom do you seek?" And they said, "Jesus of Nazareth."
JOHN|18|8|Jesus answered, "I told you that I am he. So, if you seek me, let these men go."
JOHN|18|9|This was to fulfill the word that he had spoken: "Of those whom you gave me I have lost not one."
JOHN|18|10|Then Simon Peter, having a sword, drew it and struck the high priest's servant and cut off his right ear. (The servant's name was Malchus.)
JOHN|18|11|So Jesus said to Peter, "Put your sword into its sheath; shall I not drink the cup that the Father has given me?"
JOHN|18|12|So the band of soldiers and their captain and the officers of the Jews arrested Jesus and bound him.
JOHN|18|13|First they led him to Annas, for he was the father-in-law of Caiaphas, who was high priest that year.
JOHN|18|14|It was Caiaphas who had advised the Jews that it would be expedient that one man should die for the people.
JOHN|18|15|Simon Peter followed Jesus, and so did another disciple. Since that disciple was known to the high priest, he entered with Jesus into the court of the high priest,
JOHN|18|16|but Peter stood outside at the door. So the other disciple, who was known to the high priest, went out and spoke to the servant girl who kept watch at the door, and brought Peter in.
JOHN|18|17|The servant girl at the door said to Peter, "You also are not one of this man's disciples, are you?" He said, "I am not."
JOHN|18|18|Now the servants and officers had made a charcoal fire, because it was cold, and they were standing and warming themselves. Peter also was with them, standing and warming himself.
JOHN|18|19|The high priest then questioned Jesus about his disciples and his teaching.
JOHN|18|20|Jesus answered him, "I have spoken openly to the world. I have always taught in synagogues and in the temple, where all Jews come together. I have said nothing in secret.
JOHN|18|21|Why do you ask me? Ask those who have heard me what I said to them; they know what I said."
JOHN|18|22|When he had said these things, one of the officers standing by struck Jesus with his hand, saying, "Is that how you answer the high priest?"
JOHN|18|23|Jesus answered him, "If what I said is wrong, bear witness about the wrong; but if what I said is right, why do you strike me?"
JOHN|18|24|Annas then sent him bound to Caiaphas the high priest.
JOHN|18|25|Now Simon Peter was standing and warming himself. So they said to him, "You also are not one of his disciples, are you?" He denied it and said, "I am not."
JOHN|18|26|One of the servants of the high priest, a relative of the man whose ear Peter had cut off, asked, "Did I not see you in the garden with him?"
JOHN|18|27|Peter again denied it, and at once a rooster crowed.
JOHN|18|28|Then they led Jesus from the house of Caiaphas to the governor's headquarters. It was early morning. They themselves did not enter the governor's headquarters, so that they would not be defiled, but could eat the Passover.
JOHN|18|29|So Pilate went outside to them and said, "What accusation do you bring against this man?"
JOHN|18|30|They answered him, "If this man were not doing evil, we would not have delivered him over to you."
JOHN|18|31|Pilate said to them, "Take him yourselves and judge him by your own law." The Jews said to him, "It is not lawful for us to put anyone to death."
JOHN|18|32|This was to fulfill the word that Jesus had spoken to show by what kind of death he was going to die.
JOHN|18|33|So Pilate entered his headquarters again and called Jesus and said to him, "Are you the King of the Jews?"
JOHN|18|34|Jesus answered, "Do you say this of your own accord, or did others say it to you about me?"
JOHN|18|35|Pilate answered, "Am I a Jew? Your own nation and the chief priests have delivered you over to me. What have you done?"
JOHN|18|36|Jesus answered, "My kingdom is not of this world. If my kingdom were of this world, my servants would have been fighting, that I might not be delivered over to the Jews. But my kingdom is not from the world."
JOHN|18|37|Then Pilate said to him, "So you are a king?" Jesus answered, "You say that I am a king. For this purpose I was born and for this purpose I have come into the world- to bear witness to the truth. Everyone who is of the truth listens to my voice."
JOHN|18|38|Pilate said to him, "What is truth?" After he had said this, he went back outside to the Jews and told them, "I find no guilt in him.
JOHN|18|39|But you have a custom that I should release one man for you at the Passover. So do you want me to release to you the King of the Jews?"
JOHN|18|40|They cried out again, "Not this man, but Barabbas!" Now Barabbas was a robber.
JOHN|19|1|Then Pilate took Jesus and flogged him.
JOHN|19|2|And the soldiers twisted together a crown of thorns and put it on his head and arrayed him in a purple robe.
JOHN|19|3|They came up to him, saying, "Hail, King of the Jews!" and struck him with their hands.
JOHN|19|4|Pilate went out again and said to them, "See, I am bringing him out to you that you may know that I find no guilt in him."
JOHN|19|5|So Jesus came out, wearing the crown of thorns and the purple robe. Pilate said to them, "Behold the man!"
JOHN|19|6|When the chief priests and the officers saw him, they cried out, "Crucify him, crucify him!" Pilate said to them, "Take him yourselves and crucify him, for I find no guilt in him."
JOHN|19|7|The Jews answered him, "We have a law, and according to that law he ought to die because he has made himself the Son of God."
JOHN|19|8|When Pilate heard this statement, he was even more afraid.
JOHN|19|9|He entered his headquarters again and said to Jesus, "Where are you from?" But Jesus gave him no answer.
JOHN|19|10|So Pilate said to him, "You will not speak to me? Do you not know that I have authority to release you and authority to crucify you?"
JOHN|19|11|Jesus answered him, "You would have no authority over me at all unless it had been given you from above. Therefore he who delivered me over to you has the greater sin."
JOHN|19|12|From then on Pilate sought to release him, but the Jews cried out, "If you release this man, you are not Caesar's friend. Everyone who makes himself a king opposes Caesar."
JOHN|19|13|So when Pilate heard these words, he brought Jesus out and sat down on the judgment seat at a place called The Stone Pavement, and in Aramaic Gabbatha.
JOHN|19|14|Now it was the day of Preparation of the Passover. It was about the sixth hour. He said to the Jews, "Behold your King!"
JOHN|19|15|They cried out, "Away with him, away with him, crucify him!" Pilate said to them, "Shall I crucify your King?" The chief priests answered, "We have no king but Caesar."
JOHN|19|16|So he delivered him over to them to be crucified. So they took Jesus,
JOHN|19|17|and he went out, bearing his own cross, to the place called the place of a skull, which in Aramaic is called Golgotha.
JOHN|19|18|There they crucified him, and with him two others, one on either side, and Jesus between them.
JOHN|19|19|Pilate also wrote an inscription and put it on the cross. It read, "Jesus of Nazareth, the King of the Jews."
JOHN|19|20|Many of the Jews read this inscription, for the place where Jesus was crucified was near the city, and it was written in Aramaic, in Latin, and in Greek.
JOHN|19|21|So the chief priests of the Jews said to Pilate, "Do not write, 'The King of the Jews,' but rather, 'This man said, I am King of the Jews.'"
JOHN|19|22|Pilate answered, "What I have written I have written."
JOHN|19|23|When the soldiers had crucified Jesus, they took his garments and divided them into four parts, one part for each soldier; also his tunic. But the tunic was seamless, woven in one piece from top to bottom,
JOHN|19|24|so they said to one another, "Let us not tear it, but cast lots for it to see whose it shall be." This was to fulfill the Scripture which says, "They divided my garments among them, and for my clothing they cast lots." So the soldiers did these things,
JOHN|19|25|but standing by the cross of Jesus were his mother and his mother's sister, Mary the wife of Clopas, and Mary Magdalene.
JOHN|19|26|When Jesus saw his mother and the disciple whom he loved standing nearby, he said to his mother, "Woman, behold, your son!"
JOHN|19|27|Then he said to the disciple, "Behold, your mother!" And from that hour the disciple took her to his own home.
JOHN|19|28|After this, Jesus, knowing that all was now finished, said (to fulfill the Scripture), "I thirst."
JOHN|19|29|A jar full of sour wine stood there, so they put a sponge full of the sour wine on a hyssop branch and held it to his mouth.
JOHN|19|30|When Jesus had received the sour wine, he said, "It is finished," and he bowed his head and gave up his spirit.
JOHN|19|31|Since it was the day of Preparation, and so that the bodies would not remain on the cross on the Sabbath (for that Sabbath was a high day), the Jews asked Pilate that their legs might be broken and that they might be taken away.
JOHN|19|32|So the soldiers came and broke the legs of the first, and of the other who had been crucified with him.
JOHN|19|33|But when they came to Jesus and saw that he was already dead, they did not break his legs.
JOHN|19|34|But one of the soldiers pierced his side with a spear, and at once there came out blood and water.
JOHN|19|35|He who saw it has borne witness- his testimony is true, and he knows that he is telling the truth- that you also may believe.
JOHN|19|36|For these things took place that the Scripture might be fulfilled: "Not one of his bones will be broken."
JOHN|19|37|And again another Scripture says, "They will look on him whom they have pierced."
JOHN|19|38|After these things Joseph of Arimathea, who was a disciple of Jesus, but secretly for fear of the Jews, asked Pilate that he might take away the body of Jesus, and Pilate gave him permission. So he came and took away his body.
JOHN|19|39|Nicodemus also, who earlier had come to Jesus by night, came bringing a mixture of myrrh and aloes, about seventy-five pounds in weight.
JOHN|19|40|So they took the body of Jesus and bound it in linen cloths with the spices, as is the burial custom of the Jews.
JOHN|19|41|Now in the place where he was crucified there was a garden, and in the garden a new tomb in which no one had yet been laid.
JOHN|19|42|So because of the Jewish day of Preparation, since the tomb was close at hand, they laid Jesus there.
JOHN|20|1|Now on the first day of the week Mary Magdalene came to the tomb early, while it was still dark, and saw that the stone had been taken away from the tomb.
JOHN|20|2|So she ran and went to Simon Peter and the other disciple, the one whom Jesus loved, and said to them, "They have taken the Lord out of the tomb, and we do not know where they have laid him."
JOHN|20|3|So Peter went out with the other disciple, and they were going toward the tomb.
JOHN|20|4|Both of them were running together, but the other disciple outran Peter and reached the tomb first.
JOHN|20|5|And stooping to look in, he saw the linen cloths lying there, but he did not go in.
JOHN|20|6|Then Simon Peter came, following him, and went into the tomb. He saw the linen cloths lying there,
JOHN|20|7|and the face cloth, which had been on Jesus' head, not lying with the linen cloths but folded up in a place by itself.
JOHN|20|8|Then the other disciple, who had reached the tomb first, also went in, and he saw and believed;
JOHN|20|9|for as yet they did not understand the Scripture, that he must rise from the dead.
JOHN|20|10|Then the disciples went back to their homes.
JOHN|20|11|But Mary stood weeping outside the tomb, and as she wept she stooped to look into the tomb.
JOHN|20|12|And she saw two angels in white, sitting where the body of Jesus had lain, one at the head and one at the feet.
JOHN|20|13|They said to her, "Woman, why are you weeping?" She said to them, "They have taken away my Lord, and I do not know where they have laid him."
JOHN|20|14|Having said this, she turned around and saw Jesus standing, but she did not know that it was Jesus.
JOHN|20|15|Jesus said to her, "Woman, why are you weeping? Whom are you seeking?" Supposing him to be the gardener, she said to him, "Sir, if you have carried him away, tell me where you have laid him, and I will take him away."
JOHN|20|16|Jesus said to her, "Mary." She turned and said to him in Aramaic, "Rabboni!" (which means Teacher).
JOHN|20|17|Jesus said to her, "Do not cling to me, for I have not yet ascended to the Father; but go to my brothers and say to them, 'I am ascending to my Father and your Father, to my God and your God.'"
JOHN|20|18|Mary Magdalene went and announced to the disciples, "I have seen the Lord"- and that he had said these things to her.
JOHN|20|19|On the evening of that day, the first day of the week, the doors being locked where the disciples were for fear of the Jews, Jesus came and stood among them and said to them, "Peace be with you."
JOHN|20|20|When he had said this, he showed them his hands and his side. Then the disciples were glad when they saw the Lord.
JOHN|20|21|Jesus said to them again, "Peace be with you. As the Father has sent me, even so I am sending you."
JOHN|20|22|And when he had said this, he breathed on them and said to them, "Receive the Holy Spirit.
JOHN|20|23|If you forgive the sins of anyone, they are forgiven; if you withhold forgiveness from anyone, it is withheld."
JOHN|20|24|Now Thomas, one of the Twelve, called the Twin, was not with them when Jesus came.
JOHN|20|25|So the other disciples told him, "We have seen the Lord." But he said to them, "Unless I see in his hands the mark of the nails, and place my finger into the mark of the nails, and place my hand into his side, I will never believe."
JOHN|20|26|Eight days later, his disciples were inside again, and Thomas was with them. Although the doors were locked, Jesus came and stood among them and said, "Peace be with you."
JOHN|20|27|Then he said to Thomas, "Put your finger here, and see my hands; and put out your hand, and place it in my side. Do not disbelieve, but believe."
JOHN|20|28|Thomas answered him, "My Lord and my God!"
JOHN|20|29|Jesus said to him, "Have you believed because you have seen me? Blessed are those who have not seen and yet have believed."
JOHN|20|30|Now Jesus did many other signs in the presence of the disciples, which are not written in this book;
JOHN|20|31|but these are written so that you may believe that Jesus is the Christ, the Son of God, and that by believing you may have life in his name.
JOHN|21|1|After this Jesus revealed himself again to the disciples by the Sea of Tiberias, and he revealed himself in this way.
JOHN|21|2|Simon Peter, Thomas (called the Twin), Nathanael of Cana in Galilee, the sons of Zebedee, and two others of his disciples were together.
JOHN|21|3|Simon Peter said to them, "I am going fishing." They said to him, "We will go with you." They went out and got into the boat, but that night they caught nothing.
JOHN|21|4|Just as day was breaking, Jesus stood on the shore; yet the disciples did not know that it was Jesus.
JOHN|21|5|Jesus said to them, "Children, do you have any fish?" They answered him, "No."
JOHN|21|6|He said to them, "Cast the net on the right side of the boat, and you will find some." So they cast it, and now they were not able to haul it in, because of the quantity of fish.
JOHN|21|7|That disciple whom Jesus loved therefore said to Peter, "It is the Lord!" When Simon Peter heard that it was the Lord, he put on his outer garment, for he was stripped for work, and threw himself into the sea.
JOHN|21|8|The other disciples came in the boat, dragging the net full of fish, for they were not far from the land, but about a hundred yards off.
JOHN|21|9|When they got out on land, they saw a charcoal fire in place, with fish laid out on it, and bread.
JOHN|21|10|Jesus said to them, "Bring some of the fish that you have just caught."
JOHN|21|11|So Simon Peter went aboard and hauled the net ashore, full of large fish, 153 of them. And although there were so many, the net was not torn.
JOHN|21|12|Jesus said to them, "Come and have breakfast." Now none of the disciples dared ask him, "Who are you?" They knew it was the Lord.
JOHN|21|13|Jesus came and took the bread and gave it to them, and so with the fish.
JOHN|21|14|This was now the third time that Jesus was revealed to the disciples after he was raised from the dead.
JOHN|21|15|When they had finished breakfast, Jesus said to Simon Peter, "Simon, son of John, do you love me more than these?" He said to him, "Yes, Lord; you know that I love you." He said to him, "Feed my lambs."
JOHN|21|16|He said to him a second time, "Simon, son of John, do you love me?" He said to him, "Yes, Lord; you know that I love you." He said to him, "Tend my sheep."
JOHN|21|17|He said to him the third time, "Simon, son of John, do you love me?" Peter was grieved because he said to him the third time, "Do you love me?" and he said to him, "Lord, you know everything; you know that I love you." Jesus said to him, "Feed my sheep.
JOHN|21|18|Truly, truly, I say to you, when you were young, you used to dress yourself and walk wherever you wanted, but when you are old, you will stretch out your hands, and another will dress you and carry you where you do not want to go."
JOHN|21|19|(This he said to show by what kind of death he was to glorify God.) And after saying this he said to him, "Follow me."
JOHN|21|20|Peter turned and saw the disciple whom Jesus loved following them, the one who had been reclining at table close to him and had said, "Lord, who is it that is going to betray you?"
JOHN|21|21|When Peter saw him, he said to Jesus, "Lord, what about this man?"
JOHN|21|22|Jesus said to him, "If it is my will that he remain until I come, what is that to you? You follow me!"
JOHN|21|23|So the saying spread abroad among the brothers that this disciple was not to die; yet Jesus did not say to him that he was not to die, but, "If it is my will that he remain until I come, what is that to you?"
JOHN|21|24|This is the disciple who is bearing witness about these things, and who has written these things, and we know that his testimony is true.
JOHN|21|25|Now there are also many other things that Jesus did. Were every one of them to be written, I suppose that the world itself could not contain the books that would be written.
