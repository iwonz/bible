1THESS|1|1|Paulus et Silvanus et Timo theus ecclesiae Thessalonicen sium in Deo Patre et Domino Iesu Christo: gratia vobis et pax.
1THESS|1|2|Gratias agimus Deo semper pro omnibus vobis, memoriam facientes in orationibus nostris, sine intermissione;
1THESS|1|3|memores operis fidei vestrae et laboris caritatis et sustinentiae spei Domini nostri Iesu Christi ante Deum et Patrem nostrum;
1THESS|1|4|scientes, fratres, dilecti a Deo, electionem vestram,
1THESS|1|5|quia evangelium nostrum non fuit ad vos in sermone tantum sed et in virtute et in Spiritu Sancto et in plenitudine multa, sicut scitis quales fuerimus vobis propter vos.
1THESS|1|6|Et vos imitatores nostri facti estis et Domini, excipientes verbum in tribulatione multa cum gaudio Spiritus Sancti,
1THESS|1|7|ita ut facti sitis forma omnibus credentibus in Macedonia et in Achaia.
1THESS|1|8|A vobis enim diffamatus est sermo Domini non solum in Macedonia et in Achaia, sed in omni loco fides vestra, quae est ad Deum, profecta est, ita ut non sit nobis necesse quidquam loqui;
1THESS|1|9|ipsi enim de nobis annuntiant qualem introitum habuerimus ad vos, et quomodo conversi estis ad Deum a simulacris, servire Deo vivo et vero
1THESS|1|10|et exspectare Filium eius de caelis, quem suscitavit ex mortuis, Iesum, qui eripit nos ab ira ventura.
1THESS|2|1|Nam ipsi scitis, fratres, introi tum nostrum ad vos, quia non inanis fuit;
1THESS|2|2|sed ante passi et contumeliis affecti, sicut scitis, in Philippis, fiduciam habuimus in Deo nostro loqui ad vos evangelium Dei in multa sollicitudine.
1THESS|2|3|Exhortatio enim nostra non ex errore neque ex immunditia neque in dolo,
1THESS|2|4|sed sicut probati sumus a Deo, ut crederetur nobis evangelium, ita loquimur non quasi hominibus placentes, sed Deo, qui probat corda nostra.
1THESS|2|5|Neque enim aliquando fuimus in sermone adulationis, sicut scitis, neque sub praetextu avaritiae, Deus testis,
1THESS|2|6|nec quaerentes ab hominibus gloriam, neque a vobis neque ab aliis;
1THESS|2|7|cum possemus oneri esse ut Christi apostoli, sed facti sumus parvuli in medio vestrum, tamquam si nutrix foveat filios suos;
1THESS|2|8|ita desiderantes vos, cupide volebamus tradere vobis non solum evangelium Dei sed etiam animas nostras, quoniam carissimi nobis facti estis.
1THESS|2|9|Memores enim estis, fratres, laboris nostri et fatigationis; nocte et die operantes, ne quem vestrum gravaremus, praedicavimus in vobis evangelium Dei.
1THESS|2|10|Vos testes estis et Deus, quam sancte et iuste et sine querela vobis, qui credidistis, fuimus;
1THESS|2|11|sicut scitis qualiter unumquemque vestrum, tamquam pater filios suos,
1THESS|2|12|deprecantes vos et consolantes testificati sumus, ut ambularetis digne Deo, qui vocat vos in suum regnum et gloriam.
1THESS|2|13|Ideo et nos gratias agimus Deo sine intermissione, quoniam cum accepissetis a nobis verbum auditus Dei, accepistis non ut verbum hominum sed, sicut est vere, verbum Dei, quod et operatur in vobis, qui creditis.
1THESS|2|14|Vos enim imitatores facti estis, fratres, ecclesiarum Dei, quae sunt in Iudaea in Christo Iesu; quia eadem passi estis et vos a contribulibus vestris, sicut et ipsi a Iudaeis,
1THESS|2|15|qui et Dominum occiderunt Iesum et prophetas et nos persecuti sunt et Deo non placent et omnibus hominibus adversantur,
1THESS|2|16|prohibentes nos gentibus loqui, ut salvae fiant, ut impleant peccata sua semper. Pervenit autem ira Dei super illos usque in finem.
1THESS|2|17|Nos autem, fratres, desolati a vobis ad tempus horae, facie non corde, abundantius festinavimus faciem vestram videre cum multo desiderio.
1THESS|2|18|Propter quod voluimus venire ad vos, ego quidem Paulus et semel et iterum; et impedivit nos Satanas.
1THESS|2|19|Quae est enim nostra spes aut gaudium aut corona gloriae - nonne et vos ante Dominum nostrum Iesum in adventu eius?
1THESS|2|20|Vos enim estis gloria nostra et gaudium.
1THESS|3|1|Propter quod non sustinentes amplius, placuit nobis, ut relin queremur Athenis soli,
1THESS|3|2|et misimus Timotheum, fratrem nostrum et cooperatorem Dei in evangelio Christi, ad confirmandos vos et exhortandos pro fide vestra,
1THESS|3|3|ut nemo turbetur in tribulationibus istis. Ipsi enim scitis quod in hoc positi sumus;
1THESS|3|4|nam et cum apud vos essemus, praedicebamus vobis passuros nos tribulationes, sicut et factum est et scitis.
1THESS|3|5|Propterea et ego amplius non sustinens, misi ad cognoscendam fidem vestram, ne forte tentaverit vos is qui tentat, et inanis fiat labor noster.
1THESS|3|6|Nunc autem, veniente Timotheo ad nos a vobis et annuntiante nobis fidem et caritatem vestram, et quia memoriam nostri habetis bonam semper, desiderantes nos videre, sicut nos quoque vos;
1THESS|3|7|ideo consolati sumus, fratres, propter vos in omni necessitate et tribulatione nostra per vestram fidem;
1THESS|3|8|quoniam nunc vivimus, si vos statis in Domino.
1THESS|3|9|Quam enim gratiarum actionem possumus Deo retribuere pro vobis in omni gaudio, quo gaudemus propter vos ante Deum nostrum,
1THESS|3|10|nocte et die abundantius orantes, ut videamus faciem vestram et compleamus ea, quae desunt fidei vestrae?
1THESS|3|11|Ipse autem Deus et Pater noster et Dominus noster Iesus dirigat viam nostram ad vos;
1THESS|3|12|vos autem Dominus abundare et superabundare faciat caritate in invicem et in omnes, quemadmodum et nos in vos;
1THESS|3|13|ad confirmanda corda vestra sine querela in sanctitate ante Deum et Patrem nostrum, in adventu Domini nostri Iesu cum omnibus sanctis eius. Amen.
1THESS|4|1|De cetero ergo, fratres, rogamus vos et obsecramus in Domino Iesu, ut - quemadmodum accepistis a nobis quomodo vos oporteat ambulare et placere Deo, sicut et ambulatis - ut abundetis magis.
1THESS|4|2|Scitis enim, quae praecepta dederimus vobis per Dominum Iesum.
1THESS|4|3|Haec est enim voluntas Dei, sanctificatio vestra,
1THESS|4|4|ut abstineatis a fornicatione; ut sciat unusquisque vestrum suum vas possidere in sanctificatione et honore,
1THESS|4|5|non in passione desiderii, sicut et gentes, quae ignorant Deum;
1THESS|4|6|ut ne quis supergrediatur neque circumveniat in negotio fratrem suum, quoniam vindex est Dominus de his omnibus, sicut et praediximus vobis et testificati sumus.
1THESS|4|7|Non enim vocavit nos Deus in immunditiam sed in sanctificationem.
1THESS|4|8|Itaque, qui spernit, non hominem spernit sed Deum, qui etiam dat Spiritum suum Sanctum in vos.
1THESS|4|9|De caritate autem fraternitatis non necesse habetis, ut vobis scribam; ipsi enim vos a Deo edocti estis, ut diligatis invicem;
1THESS|4|10|etenim facitis illud in omnes fratres in universa Macedonia. Rogamus autem vos, fratres, ut abundetis magis;
1THESS|4|11|et operam detis, ut quieti sitis et ut vestrum negotium agatis et operemini manibus vestris, sicut praecipimus vobis;
1THESS|4|12|ut honeste ambuletis ad eos, qui foris sunt, et nullius aliquid desideretis.
1THESS|4|13|Nolumus autem vos ignorare, fratres, de dormientibus, ut non contristemini sicut et ceteri, qui spem non habent.
1THESS|4|14|Si enim credimus quod Iesus mortuus est et resurrexit, ita et Deus eos, qui dormierunt, per Iesum adducet cum eo.
1THESS|4|15|Hoc enim vobis dicimus in verbo Domini, quia nos, qui vivimus, qui relinquimur in adventum Domini, non praeveniemus eos, qui dormierunt;
1THESS|4|16|quoniam ipse Dominus in iussu, in voce archangeli et in tuba Dei descendet de caelo, et mortui, qui in Christo sunt, resurgent primi;
1THESS|4|17|deinde nos, qui vivimus, qui relinquimur, simul rapiemur cum illis in nubibus obviam Domino in aera, et sic semper cum Domino erimus.
1THESS|4|18|Itaque consolamini invicem in verbis istis.
1THESS|5|1|De temporibus autem et mo mentis, fratres, non indigetis, ut scribatur vobis;
1THESS|5|2|ipsi enim diligenter scitis quia dies Domini, sicut fur in nocte, ita veniet.
1THESS|5|3|Cum enim dixerint: " Pax et securitas ", tunc repentinus eis superveniet interitus, sicut dolor in utero habenti, et non effugient.
1THESS|5|4|Vos autem, fratres, non estis in tenebris, ut vos dies ille tamquam fur comprehendat;
1THESS|5|5|omnes enim vos filii lucis estis et filii diei. Non sumus noctis neque tenebrarum;
1THESS|5|6|igitur non dormiamus sicut ceteri, sed vigilemus et sobrii simus.
1THESS|5|7|Qui enim dormiunt, nocte dormiunt; et, qui ebrii sunt, nocte inebriantur.
1THESS|5|8|Nos autem, qui diei sumus, sobrii simus, induti loricam fidei et caritatis et galeam spem salutis;
1THESS|5|9|quoniam non posuit nos Deus in iram sed in acquisitionem salutis per Dominum nostrum Iesum Christum,
1THESS|5|10|qui mortuus est pro nobis, ut sive vigilemus sive dormiamus, simul cum illo vivamus.
1THESS|5|11|Propter quod consolamini invicem et aedificate alterutrum, sicut et facitis.
1THESS|5|12|Rogamus autem vos, fratres, ut noveritis eos, qui laborant inter vos et praesunt vobis in Domino et monent vos,
1THESS|5|13|ut habeatis illos superabundanter in caritate propter opus illorum. Pacem habete inter vos.
1THESS|5|14|Hortamur autem vos, fratres: corripite inquietos, consolamini pusillanimes, suscipite infirmos, longanimes estote ad omnes.
1THESS|5|15|Videte, ne quis malum pro malo alicui reddat, sed semper, quod bonum est, sectamini et in invicem et in omnes.
1THESS|5|16|Semper gaudete,
1THESS|5|17|sine intermissione orate,
1THESS|5|18|in omnibus gratias agite; haec enim voluntas Dei est in Christo Iesu erga vos.
1THESS|5|19|Spiritum nolite exstinguere,
1THESS|5|20|prophetias nolite spernere;
1THESS|5|21|omnia autem probate, quod bonum est tenete,
1THESS|5|22|ab omni specie mala abstinete vos.
1THESS|5|23|Ipse autem Deus pacis sanctificet vos per omnia, et integer spiritus vester et anima et corpus sine querela in adventu Domini nostri Iesu Christi servetur.
1THESS|5|24|Fidelis est, qui vocat vos, qui etiam faciet.
1THESS|5|25|Fratres, orate etiam pro nobis.
1THESS|5|26|Salutate fratres omnes in osculo sancto.
1THESS|5|27|Adiuro vos per Dominum, ut legatur epistula omnibus fratribus.
1THESS|5|28|Gratia Domini nostri Iesu Christi vobiscum.
