HAB|1|1|Oraculum, quod vidit Habacuc propheta.
HAB|1|2|Usquequo, Domine, clamabo,et non exaudis?Vociferabor ad te: " Violentia! ",et non salvas?
HAB|1|3|Quare ostendisti mihi iniquitatemet malitiam vides?Et vastitas et violentia est coram me,et facta est contentio, et iurgium exoritur.
HAB|1|4|Propter hoc languet lex,et non pervenit usque ad finem iudicium.Quia impius praevalet adversus iustum,propterea egreditur iudicium perversum.
HAB|1|5|" Aspicite in gentibus et videte,admiramini et obstupescite,quia opus facio in diebus vestris,quod nemo credet, cum narrabitur.
HAB|1|6|Quia ecce ego suscitabo Chaldaeos,gentem amaram et velocem,ambulantem super latitudinem terrae,ut possideat tabernacula non sua.
HAB|1|7|Horribilis et terribilis est,ex semetipsa iudicium eiuset maiestas eius egredietur.
HAB|1|8|Leviores pardis equi eiuset saeviores lupis deserti;et accurrunt equites eius:equites namque eius de longe venient,volabunt quasi aquilafestinans ad comedendum.
HAB|1|9|Omnes, ut violentiam faciant, venient,omnes facies eorum ventus urens;et congregabunt quasi arenam captivos.
HAB|1|10|Et ipsa reges subsannabit,tyrannis illudet;ipsa super omnem munitionem ridebitet comportabit aggerem et capiet eam.
HAB|1|11|Tunc ultra progrediens quasi ventus pertransibitet constituet fortitudinem suam deum suum ".
HAB|1|12|Numquid non tu a principio, Domine,Deus meus, sanctus meus,qui non morieris?Domine, ad iudicium posuisti eam; petra mea, ad corripiendum fundasti eam.
HAB|1|13|Mundi sunt oculi tui, ne videas malum;et respicere ad iniquitatem non poteris.Quare respicis super inique agentes et taces, devorante impio iustiorem se?
HAB|1|14|Fecisti homines quasi pisces maris,quasi reptile non habens principem super se.
HAB|1|15|Omnes in hamo sublevat,trahit eos in sagena suaet congregat in rete suo;super hoc laetatur et exsultat.
HAB|1|16|Propterea immolat sagenae suaeet sacrificat reti suo,quia in ipsis incrassata est portio eius,et cibus eius pinguis.
HAB|1|17|Propter hoc ergo evaginabit gladium suum semper,ut interficiat gentes sine misericordia?
HAB|2|1|Super custodiam meam staboet consistam super speculamet contemplabor, ut videam quid dicat mihiet quid respondeat ad querelam meam.
HAB|2|2|Et respondit mihi Dominus et dixit: Scribe visumet explana eum super tabulas,ut percurrat, qui legerit eum.
HAB|2|3|Quia adhuc visus ad tempus constitutum,sed anhelat in finem et non mentietur;si moram fecerit, exspecta illum,quia veniens veniet et non tardabit.
HAB|2|4|Ecce languidus, in quo non est anima recta;iustus autem in fide sua vivet ".
HAB|2|5|Et profecto divitiae decipiunt virum superbum,et non perveniet ad finem;qui dilatat quasi infernus fauces suaset ipse quasi mors et non adimpletur:et congregat ad se omnes genteset coacervat ad se omnes populos.
HAB|2|6|Numquid non omnes isti super eum parabolam sumentet loquelam aenigmatum dicentes: Vae ei, qui multiplicat non sua - usquequo? Cet aggravat pignora super se! ".
HAB|2|7|Numquid non repente consurgent, qui mordeant te,et evigilabunt agitantes te,et eris in rapinam eis?
HAB|2|8|Quia tu spoliasti gentes multas,spoliabunt te omnes, qui reliqui fuerint de populis;propter sanguinem hominum et oppressionem terrae,civitatum et omnium habitantium in eis.
HAB|2|9|Vae, qui congregat lucrum iniustum in malum domui suae,ut ponat in excelso nidum suumet salvet se de manu mali!
HAB|2|10|Consilium cepisti in confusionem domui tuaeconcidendi populos multoset peccasti in animam tuam.
HAB|2|11|Quia lapis de pariete clamabit,et trabes de contignatione respondebit ei.
HAB|2|12|Vae, qui aedificat civitatem in sanguinibuset condit urbem in iniquitate!
HAB|2|13|Numquid non haec a Domino sunt exercituum,ut laborent populi pro igne,et gentes in vacuum fatigentur?
HAB|2|14|Quia replebitur terra cognitione gloriae Domini,sicut aquae operiunt mare.
HAB|2|15|Vae, qui potum dat amico suomittens venenum suum et inebrians eum,ut aspiciat nuditatem eius!
HAB|2|16|Repleris ignominia pro gloria;bibe tu quoque et denudare!Transibit ad te calix dexterae Domini,et veniet ignominia super gloriam tuam.
HAB|2|17|Quia vastitas Libani operiet te,et miseria animalium deterrebit tepropter sanguinem hominum et oppressionem terrae,civitatum et omnium habitantium in eis.
HAB|2|18|Quid prodest sculptile,quia sculpsit illud fictor suus;conflatile et oraculum mendax,quia speravit in figmento fictor eius, ut faceret simulacra muta?
HAB|2|19|Vae, qui dicit ligno: " Expergiscere! ", " Surge! " lapidi tacenti!Numquid ipse docere poterit?Ecce iste coopertus est auro et argento,et omnis spiritus non est in visceribus eius.
HAB|2|20|Dominus autem in templo sancto suo; sileat a facie eius omnis terra.
HAB|3|1|Oratio Habacuc prophetae.Secundum melodiam lamentationum.
HAB|3|2|Domine, audivi auditionem tuamet timui, Domine, opus tuum.In medio annorum vivifica illud,in medio annorum notum facies.Cum iratus fueris, misericordiae recordaberis.
HAB|3|3|Deus a Theman veniet,et Sanctus de monte Pharan. - Selah.Operit caelos gloria eius,et laudis eius plena est terra.
HAB|3|4|Splendor eius ut lux erit,radii ex manibus eius:ibi abscondita est fortitudo eius.
HAB|3|5|Ante faciem eius ibit mors,et egredietur pestis post pedes eius.
HAB|3|6|Stetit et concussit terram,aspexit et dissolvit gentes.Et contriti sunt montes saeculi,incurvati sunt colles antiquiab itineribus aeternitatis eius.
HAB|3|7|In afflictione vidi tentoria Chusan;turbantur pelles terrae Madian.
HAB|3|8|Numquid in fluminibus iratus es, Domine,aut in fluminibus furor tuusvel in mari indignatio tua?Quia ascendes super equos tuos,quadrigas tuas victrices.
HAB|3|9|Suscitans suscitabis arcum tuum,sagittis replevisti pharetram tuam. - Selah.In fluvios scindes terram,
HAB|3|10|viderunt te et doluerunt montes.Effuderunt aquas nubes,dedit abyssus vocem suam,in altum levavit manus suas.
HAB|3|11|Sol et luna steterunt in habitaculo suo,prae luce sagittarum tuarum discedunt,prae splendore fulgurantis hastae tuae.
HAB|3|12|In fremitu calcabis terram,in furore conteres gentes.
HAB|3|13|Egressus es in salutem populi tui,in salutem cum christo tuo.Percussisti caput de domo impii,denudasti fundamentum usque ad petram. - Selah.
HAB|3|14|Confodisti iaculis tuis caput bellatorum eius,venientium ut turbo ad dispergendum me;exsultatio eorum, sicut eius, qui devorat pauperem in abscondito.
HAB|3|15|Viam fecisti in mari equis tuis,in luto aquarum multarum.
HAB|3|16|Audivi, et conturbatus est venter meus,ad vocem contremuerunt labia mea. Ingreditur putredo in ossibus meis, et subter me vacillant gressus mei.Conquiescam in die tribulationis,ut ascendat super populum, qui invadit nos.
HAB|3|17|Ficus enim non florebit,et non erit fructus in vineis;mentietur opus olivae,et arva non afferent cibum;abscissum est de ovili pecus,et non est armentum in praesepibus.
HAB|3|18|Ego autem in Domino gaudeboet exsultabo in Deo salvatore meo.
HAB|3|19|Dominus Deus fortitudo meaet ponet pedes meos quasi cervorum et super excelsa mea deducet me.Magistro chori. Ad sonitum chordarum.
