PHLM|1|1|Павел, узник Иисуса Христа, и Тимофей брат, Филимону возлюбленному и сотруднику нашему,
PHLM|1|2|и Апфии, (сестре) возлюбленной, и Архиппу, сподвижнику нашему, и домашней твоей церкви:
PHLM|1|3|благодать вам и мир от Бога Отца нашего и Господа Иисуса Христа.
PHLM|1|4|Благодарю Бога моего, всегда вспоминая о тебе в молитвах моих,
PHLM|1|5|слыша о твоей любви и вере, которую имеешь к Господу Иисусу и ко всем святым,
PHLM|1|6|дабы общение веры твоей оказалось деятельным в познании всякого у вас добра во Христе Иисусе.
PHLM|1|7|Ибо мы имеем великую радость и утешение в любви твоей, потому что тобою, брат, успокоены сердца святых.
PHLM|1|8|Посему, имея великое во Христе дерзновение приказывать тебе, что должно,
PHLM|1|9|по любви лучше прошу, не иной кто, как я, Павел старец, а теперь и узник Иисуса Христа;
PHLM|1|10|прошу тебя о сыне моем Онисиме, которого родил я в узах моих:
PHLM|1|11|он был некогда негоден для тебя, а теперь годен тебе и мне; я возвращаю его;
PHLM|1|12|ты же прими его, как мое сердце.
PHLM|1|13|Я хотел при себе удержать его, дабы он вместо тебя послужил мне в узах [за] благовествование;
PHLM|1|14|но без твоего согласия ничего не хотел сделать, чтобы доброе дело твое было не вынужденно, а добровольно.
PHLM|1|15|Ибо, может быть, он для того на время отлучился, чтобы тебе принять его навсегда,
PHLM|1|16|не как уже раба, но выше раба, брата возлюбленного, особенно мне, а тем больше тебе, и по плоти и в Господе.
PHLM|1|17|Итак, если ты имеешь общение со мною, то прими его, как меня.
PHLM|1|18|Если же он чем обидел тебя, или должен, считай это на мне.
PHLM|1|19|Я, Павел, написал моею рукою: я заплачу; не говорю тебе о том, что ты и самим собою мне должен.
PHLM|1|20|Так, брат, дай мне воспользоваться от тебя в Господе; успокой мое сердце в Господе.
PHLM|1|21|Надеясь на послушание твое, я написал к тебе, зная, что ты сделаешь и более, нежели говорю.
PHLM|1|22|А вместе приготовь для меня и помещение; ибо надеюсь, что по молитвам вашим я буду дарован вам.
PHLM|1|23|Приветствует тебя Епафрас, узник вместе со мною ради Христа Иисуса,
PHLM|1|24|Марк, Аристарх, Димас, Лука, сотрудники мои.
PHLM|1|25|Благодать Господа нашего Иисуса Христа со духом вашим. Аминь.
