TITUS|1|1|Paul, a servant of God, and an apostle of Jesus Christ, according to the faith of God's elect, and the acknowledging of the truth which is after godliness;
TITUS|1|2|In hope of eternal life, which God, that cannot lie, promised before the world began;
TITUS|1|3|But hath in due times manifested his word through preaching, which is committed unto me according to the commandment of God our Saviour;
TITUS|1|4|To Titus, mine own son after the common faith: Grace, mercy, and peace, from God the Father and the Lord Jesus Christ our Saviour.
TITUS|1|5|For this cause left I thee in Crete, that thou shouldest set in order the things that are wanting, and ordain elders in every city, as I had appointed thee:
TITUS|1|6|If any be blameless, the husband of one wife, having faithful children not accused of riot or unruly.
TITUS|1|7|For a bishop must be blameless, as the steward of God; not selfwilled, not soon angry, not given to wine, no striker, not given to filthy lucre;
TITUS|1|8|But a lover of hospitality, a lover of good men, sober, just, holy, temperate;
TITUS|1|9|Holding fast the faithful word as he hath been taught, that he may be able by sound doctrine both to exhort and to convince the gainsayers.
TITUS|1|10|For there are many unruly and vain talkers and deceivers, specially they of the circumcision:
TITUS|1|11|Whose mouths must be stopped, who subvert whole houses, teaching things which they ought not, for filthy lucre's sake.
TITUS|1|12|One of themselves, even a prophet of their own, said, The Cretians are alway liars, evil beasts, slow bellies.
TITUS|1|13|This witness is true. Wherefore rebuke them sharply, that they may be sound in the faith;
TITUS|1|14|Not giving heed to Jewish fables, and commandments of men, that turn from the truth.
TITUS|1|15|Unto the pure all things are pure: but unto them that are defiled and unbelieving is nothing pure; but even their mind and conscience is defiled.
TITUS|1|16|They profess that they know God; but in works they deny him, being abominable, and disobedient, and unto every good work reprobate.
TITUS|2|1|But speak thou the things which become sound doctrine:
TITUS|2|2|That the aged men be sober, grave, temperate, sound in faith, in charity, in patience.
TITUS|2|3|The aged women likewise, that they be in behaviour as becometh holiness, not false accusers, not given to much wine, teachers of good things;
TITUS|2|4|That they may teach the young women to be sober, to love their husbands, to love their children,
TITUS|2|5|To be discreet, chaste, keepers at home, good, obedient to their own husbands, that the word of God be not blasphemed.
TITUS|2|6|Young men likewise exhort to be sober minded.
TITUS|2|7|In all things shewing thyself a pattern of good works: in doctrine shewing uncorruptness, gravity, sincerity,
TITUS|2|8|Sound speech, that cannot be condemned; that he that is of the contrary part may be ashamed, having no evil thing to say of you.
TITUS|2|9|Exhort servants to be obedient unto their own masters, and to please them well in all things; not answering again;
TITUS|2|10|Not purloining, but shewing all good fidelity; that they may adorn the doctrine of God our Saviour in all things.
TITUS|2|11|For the grace of God that bringeth salvation hath appeared to all men,
TITUS|2|12|Teaching us that, denying ungodliness and worldly lusts, we should live soberly, righteously, and godly, in this present world;
TITUS|2|13|Looking for that blessed hope, and the glorious appearing of the great God and our Saviour Jesus Christ;
TITUS|2|14|Who gave himself for us, that he might redeem us from all iniquity, and purify unto himself a peculiar people, zealous of good works.
TITUS|2|15|These things speak, and exhort, and rebuke with all authority. Let no man despise thee.
TITUS|3|1|Put them in mind to be subject to principalities and powers, to obey magistrates, to be ready to every good work,
TITUS|3|2|To speak evil of no man, to be no brawlers, but gentle, shewing all meekness unto all men.
TITUS|3|3|For we ourselves also were sometimes foolish, disobedient, deceived, serving divers lusts and pleasures, living in malice and envy, hateful, and hating one another.
TITUS|3|4|But after that the kindness and love of God our Saviour toward man appeared,
TITUS|3|5|Not by works of righteousness which we have done, but according to his mercy he saved us, by the washing of regeneration, and renewing of the Holy Ghost;
TITUS|3|6|Which he shed on us abundantly through Jesus Christ our Saviour;
TITUS|3|7|That being justified by his grace, we should be made heirs according to the hope of eternal life.
TITUS|3|8|This is a faithful saying, and these things I will that thou affirm constantly, that they which have believed in God might be careful to maintain good works. These things are good and profitable unto men.
TITUS|3|9|But avoid foolish questions, and genealogies, and contentions, and strivings about the law; for they are unprofitable and vain.
TITUS|3|10|A man that is an heretick after the first and second admonition reject;
TITUS|3|11|Knowing that he that is such is subverted, and sinneth, being condemned of himself.
TITUS|3|12|When I shall send Artemas unto thee, or Tychicus, be diligent to come unto me to Nicopolis: for I have determined there to winter.
TITUS|3|13|Bring Zenas the lawyer and Apollos on their journey diligently, that nothing be wanting unto them.
TITUS|3|14|And let our's also learn to maintain good works for necessary uses, that they be not unfruitful.
TITUS|3|15|All that are with me salute thee. Greet them that love us in the faith. Grace be with you all. Amen.
