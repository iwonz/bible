HEB|1|1|古時候，上帝藉著眾先知多次多方向列祖說話，
HEB|1|2|末世，藉著他兒子向我們說話，又立他為承受萬有的，也藉著他創造宇宙。
HEB|1|3|他是上帝榮耀的光輝，是上帝本體的真像，常用他大能的命令托住萬有。他洗淨了人的罪，就坐在高天至大者的右邊。
HEB|1|4|他所承受的名比天使的名更尊貴，所以他遠比天使崇高。
HEB|1|5|上帝曾對哪一個天使說過： 「你是我的兒子； 我今日生了你」？ 又說過： 「我要作他的父； 他要作我的子」呢？
HEB|1|6|再者，上帝引領他長子 進入世界的時候，說： 「上帝的使者都要拜他。」
HEB|1|7|關於使者，他說： 「上帝以風為使者， 以火焰為僕役。」
HEB|1|8|關於子，他卻說： 「上帝啊，你的寶座是永永遠遠的； 你國度的權杖是正直的權杖。
HEB|1|9|你喜愛公義，恨惡罪惡； 所以上帝，就是你的上帝，用喜樂油膏你， 勝過膏你的同伴。」
HEB|1|10|他又說： 「主啊，你起初立了地的根基， 天也是你手所造的。
HEB|1|11|天地都會消滅，你卻長存； 天地都會像衣服漸漸舊了；
HEB|1|12|你要將天地捲起來，像捲一件外衣， 天地像衣服都會改變。 你卻永不改變； 你的年數沒有窮盡。」
HEB|1|13|上帝曾對哪一個天使說： 「你坐在我的右邊， 等我使你的仇敵作你的腳凳」？
HEB|1|14|眾天使不都是事奉的靈，奉差遣為那將要承受救恩的人服務的嗎？
HEB|2|1|所以，我們必須越發注意所聽見的道，免得我們隨流失去。
HEB|2|2|既然那藉著天使所傳的話是確定的，凡違背不聽從的，都受了該受的報應；
HEB|2|3|我們若忽略這麼大的救恩，怎能逃避呢？這拯救起先是主親自講的，後來是聽見的人給我們證實了。
HEB|2|4|上帝又按自己的旨意，更用神蹟奇事、百般的異能，和聖靈所給的恩賜，與他們一同作見證。
HEB|2|5|我們所說將來的世界，上帝沒有交給天使管轄。
HEB|2|6|但有人在某處證明說： 「人算甚麼，你竟顧念他； 世人算甚麼，你竟眷顧他。
HEB|2|7|你使他暫時比天使微小 ， 賜他榮耀尊貴為冠冕， 你派他管理你手所造的，
HEB|2|8|使萬物都服在他的腳下。」 既然使萬物都服他 ，就沒有剩下一樣不服他的了。只是如今我們還不見萬物都服他；
HEB|2|9|惟獨見那成為暫時比天使微小的耶穌，因為受了死的痛苦，得了尊貴榮耀為冠冕，好使他因著上帝的恩，為人人經歷了死亡。
HEB|2|10|原來那為萬物所屬、為萬物所本的，為要領許多兒子進入榮耀，使救他們的元帥因受苦難而得以完全，本是合宜的。
HEB|2|11|因那使人成聖的，和那些得以成聖的，都是出於一。為這緣故，他稱他們為弟兄也不以為恥，
HEB|2|12|說： 「我要將你的名傳給我的弟兄， 在會眾中我要頌揚你。」
HEB|2|13|他又說： 「我要依賴他。」 他又說： 「看哪！我與上帝所給我的兒女都在這裏。」
HEB|2|14|既然兒女同有血肉之軀，他也照樣親自成了血肉之軀，為能藉著死敗壞那掌管死權的，就是魔鬼，
HEB|2|15|並要釋放那些一生因怕死而作奴隸的人。
HEB|2|16|誠然，他並沒有幫助天使，而是幫助了 亞伯拉罕 的後裔。
HEB|2|17|所以，他凡事應當與他的弟兄相同，為要在上帝的事上成為慈悲忠信的大祭司，為百姓的罪獻上贖罪祭。
HEB|2|18|既然他自己被試探而受苦，他能幫助被試探的人。
HEB|3|1|同蒙天召的聖潔弟兄啊，要思想我們所宣認為使者、為大祭司的耶穌；
HEB|3|2|他向指派他的盡忠，如同 摩西 向上帝的全 家盡忠一樣。
HEB|3|3|他比 摩西 配得更多的榮耀，好像建造房屋的人比房屋更尊榮；
HEB|3|4|因為房屋都必有人建造，但建造萬物的是上帝。
HEB|3|5|摩西 作為僕人，向上帝的全家盡忠，為將來要談論的事作證；
HEB|3|6|但是基督作為兒子，治理上帝的家。我們若堅持因盼望而有的膽量和誇耀，我們就是他的家了。
HEB|3|7|所以，正如聖靈所說： 「今日，你們若聽他的話，
HEB|3|8|就不可硬著心，像在背叛之時， 就如在曠野受試探之日。
HEB|3|9|在那裏，你們的祖宗試探我， 並且觀看我的作為，
HEB|3|10|有四十年之久。 所以，我厭煩那世代， 說：他們的心常常迷糊， 竟不知道我的道路！
HEB|3|11|我在怒中起誓： 他們斷不可進入我的安息！」
HEB|3|12|弟兄們，你們要謹慎，免得你們中間有人存著邪惡不信的心，離棄了永生的上帝。
HEB|3|13|總要趁著還有今日，天天彼此相勸，免得你們中間有人被罪迷惑，心腸剛硬了。
HEB|3|14|只要我們將起初確實的信心堅持到底，就在基督裏有份了。
HEB|3|15|經上說： 「今日，你們若聽他的話， 就不可硬著心，像在背叛之時。」
HEB|3|16|聽見他而又背叛他的是誰呢？豈不是跟著 摩西 從 埃及 出來的眾人嗎？
HEB|3|17|上帝向誰發怒四十年之久呢？豈不是那些犯罪而陳屍在曠野的人嗎？
HEB|3|18|他向誰起誓，不容他們進入他的安息呢？豈不是向那些不信從的人嗎？
HEB|3|19|這樣看來，他們不能進入安息是因為不信的緣故了。
HEB|4|1|所以，既然進入他安息的應許依舊存在，我們就該存畏懼的心，免得我們 中間有人似乎沒有得到安息。
HEB|4|2|因為的確有福音傳給我們像傳給他們一樣；只是所聽見的道對他們無益，因為他們沒有以信心與所聽見的道配合。
HEB|4|3|但我們已經信的人進入安息，正如上帝所說： 「我在怒中起誓： 他們斷不可進入我的安息！」 其實造物之工，從創世以來已經完成了。
HEB|4|4|論到第七日，有一處說：「到第七日，上帝就歇了他一切工作。」
HEB|4|5|又有一處說：「他們斷不可進入我的安息！」
HEB|4|6|既有這安息保留著讓一些人進入，那些先前聽見福音的人，因不信從而不得進去，
HEB|4|7|所以上帝多年後藉著 大衛 的書，又定了一天—「今日」，如以上所引的說： 「今日，你們若聽他的話， 就不可硬著心。」
HEB|4|8|若是 約書亞 已使他們享了安息，後來上帝就不會再提別的日子了。
HEB|4|9|這樣看來，另有一安息日的安息為上帝的子民保留著。
HEB|4|10|因為那些進入安息的，也是歇了自己的工作，正如上帝歇了他的工作一樣。
HEB|4|11|所以，我們務必竭力進入那安息，免得有人學了不順從而跌倒了。
HEB|4|12|上帝的道是活潑的，是有功效的，比一切兩刃的劍更鋒利，甚至魂與靈、骨節與骨髓，都能刺入、剖開，連心中的思念和主意都能辨明。
HEB|4|13|被造的，沒有一樣在他面前不是顯露的；萬物在他眼前都是赤露敞開的，我們必須向他交賬。
HEB|4|14|既然我們有一位偉大、進入高天的大祭司，就是耶穌—上帝的兒子，我們應當持定所宣認的道。
HEB|4|15|因為我們的大祭司並非不能體恤我們的軟弱；他也在各方面受過試探，與我們一樣，只是他沒有犯罪。
HEB|4|16|所以，我們只管坦然無懼地來到施恩的寶座前，為要得憐憫，蒙恩惠，作及時的幫助。
HEB|5|1|凡從人間挑選的大祭司都是奉派替人辦理屬上帝的事，要為罪獻上禮物和祭物 。
HEB|5|2|他能體諒無知和迷失的人，因為他自己也是被軟弱所困，
HEB|5|3|因此他理當為百姓和自己的罪獻祭。
HEB|5|4|沒有人可擅自取得大祭司的尊榮，惟有蒙上帝所選召的才可以，像 亞倫 一樣。
HEB|5|5|同樣，基督也沒有自取作大祭司的榮耀，而是在乎向他說話的那一位，他說： 「你是我的兒子， 我今日生了你。」
HEB|5|6|就如又有一處說： 「你是照著 麥基洗德 的體系 永遠為祭司。」
HEB|5|7|基督在他肉身的日子，曾大聲哀哭，流淚禱告，懇求那能救他免死的上帝，就因他的虔誠蒙了應允。
HEB|5|8|他雖然為兒子，還是因所受的苦難學了順從。
HEB|5|9|既然他得以完全，就為凡順從他的人成了永遠得救的根源，
HEB|5|10|並蒙上帝照著 麥基洗德 的體系宣稱他為大祭司。
HEB|5|11|論到這事，我們有好些話要說，可是很難解釋，因為你們聽不進去。
HEB|5|12|按時間說，你們早該作教師了，誰知還需要有人再將上帝聖言基礎的要道教導你們；你們成了那需要吃奶、不能吃乾糧的人。
HEB|5|13|凡只能吃奶的，就不熟練仁義的道理，因為他是嬰孩。
HEB|5|14|惟獨長大成人的才能吃乾糧，他們的心竅因練習而靈活，能分辨善惡了。
HEB|6|1|所以，我們應當離開基督道理的基礎，竭力進到成熟的地步；不必再立根基，就如懊悔致死的行為、信靠上帝、
HEB|6|2|各樣洗禮、按手禮、死人復活，以及永遠的審判等的教導。
HEB|6|3|上帝若准許，我們就這樣做。
HEB|6|4|論到那些已經蒙了光照、嘗過天恩的滋味、又於聖靈有份、並嘗過上帝的話的美味，和來世權能的人，若再離棄真道，就不可能使他們重新懊悔了；因為他們親自把上帝的兒子重釘十字架，公然羞辱他。
HEB|6|5|
HEB|6|6|
HEB|6|7|就如一塊田地吸收過屢次下的雨水，生長蔬菜，合乎耕種的人用，就從上帝得福。
HEB|6|8|這塊田地若長荊棘和蒺藜，必被廢棄，近於詛咒，結局就是焚燒。
HEB|6|9|親愛的，雖然這樣說，我們仍深信你們有更好的情況，更接近救恩。
HEB|6|10|因為上帝並非不公義，竟忘記你們的工作和你們為他的名所顯的愛心，就是你們過去和現在伺候聖徒的愛心。
HEB|6|11|我們盼望你們各人都顯出同樣的熱忱，一直到底，好達成所確信的指望。
HEB|6|12|這樣你們才不會懶惰，卻成為效法那些藉著信和忍耐承受應許的人。
HEB|6|13|當初上帝應許 亞伯拉罕 的時候，因為沒有比自己更大的可以指著起誓，就指著自己起誓，
HEB|6|14|說：「我必多多賜福給你；我必使你大大增多。」
HEB|6|15|這樣， 亞伯拉罕 因恆心等待而得了所應許的。
HEB|6|16|人都是指著比自己大的起誓，並且以起誓作保證，了結各樣的爭論。
HEB|6|17|照樣，上帝願意為那承受應許的人更有力地顯明他的旨意不可更改，他以起誓作保證。
HEB|6|18|藉這兩件不可更改的事—在這些事上，上帝絕不會說謊—我們這些逃往避難所的人能得到強有力的鼓勵，去抓住那擺在我們前頭的指望。
HEB|6|19|我們有這指望，如同靈魂的錨，又堅固又牢靠，進入幔子後面的至聖所。
HEB|6|20|為我們作先鋒的耶穌，既照著 麥基洗德 的體系成了永遠的大祭司，已經進入了。
HEB|7|1|這 麥基洗德 就是 撒冷 王，是至高上帝的祭司。他在 亞伯拉罕 打敗諸王回來的時候迎接他，並給他祝福。
HEB|7|2|亞伯拉罕 也將自己所得來的一切，取十分之一給他。他頭一個名字翻譯出來是「公義的王」，他又名「 撒冷 王」，是和平王的意思。
HEB|7|3|他無父、無母、無族譜、無生之始、無命之終，是與上帝的兒子相似，他永遠作祭司。
HEB|7|4|你們想一想，這個人多麼偉大啊！連先祖 亞伯拉罕 都拿戰利品的十分之一給他。
HEB|7|5|那得祭司職分的 利未 子孫，奉命照例向百姓取十分之一，這百姓是自己的弟兄，雖是從 亞伯拉罕 親身生的，還是照例取十分之一。
HEB|7|6|惟獨 麥基洗德 那不與他們同族譜的，從 亞伯拉罕 收取了十分之一，並且給蒙應許的 亞伯拉罕 祝福。
HEB|7|7|向來位分大的給位分小的祝福，這是無可爭議的。
HEB|7|8|在這事上，一方面，收取十分之一的都是必死的人；另一方面，收取十分之一的卻是那位被證實是活著的。
HEB|7|9|我們可以說，那接受十分之一的 利未 也是藉著 亞伯拉罕 納了十分之一，
HEB|7|10|因為 麥基洗德 迎接 亞伯拉罕 的時候， 利未 還在他先祖的身體裏面。
HEB|7|11|那麼，如果百姓藉著 利未 人的祭司職任能達到完全—因為百姓是在這職分下領受律法的—為甚麼還需要按照 麥基洗德 的體系另外興起一位祭司，而不按照 亞倫 的體系呢？
HEB|7|12|既然祭司的職分已更改，律法也需要更改。
HEB|7|13|因為這些話所指的人本屬別的支派，那支派裏從來沒有一人在祭壇前事奉的。
HEB|7|14|很明顯地，我們的主是從 猶大 出來的；但關於這支派， 摩西 並沒有提到祭司。
HEB|7|15|倘若有另一位像 麥基洗德 的祭司興起來，我的話就更顯而易見了。
HEB|7|16|他成為祭司，並不是照屬肉身的條例，而是照無窮 生命的大能。
HEB|7|17|因為有給他作見證的說： 「你是照著 麥基洗德 的體系 永遠為祭司。」
HEB|7|18|一方面，先前的誡命因軟弱無能而廢掉了，
HEB|7|19|（律法本來就不能成就甚麼）；另一方面，一個更好的指望被引進來，靠這指望，我們就可以親近上帝。
HEB|7|20|再者，耶穌成為祭司，並不是沒有上帝的誓言；其他的祭司被指派時並沒有這種誓言，
HEB|7|21|只有耶穌是起誓立的，因為那位立他的對他說： 「主起了誓， 絕不改變。 你是永遠為祭司。」
HEB|7|22|既是起誓立的，耶穌也作了更美之約的中保。
HEB|7|23|一方面，那些成為祭司的數目本來多，是因為受死亡限制不能長久留住。
HEB|7|24|另一方面，這位既是永遠留住的，他具有不可更換的祭司職任。
HEB|7|25|所以，凡靠著他進到上帝面前的人，他都能拯救到底，因為他長遠活著為他們祈求。
HEB|7|26|這樣一位聖潔、無邪惡、無玷污、遠離罪人、高過諸天的大祭司，對我們是最合適的；
HEB|7|27|他不像那些大祭司，每日必須先為自己的罪，後為百姓的罪獻祭，因為他只一次將自己獻上就把這事成全了。
HEB|7|28|律法所立的大祭司本是有弱點的人，但在律法以後，上帝以起誓的話立了兒子為大祭司，成為完全，直到永遠。
HEB|8|1|我們所講的事，其中第一要緊的就是：我們有這樣一位大祭司，他已經坐在天上至大者寶座的右邊，
HEB|8|2|在聖所，就是在真帳幕裏作僕役；這帳幕是主所支搭的，不是人所支搭的。
HEB|8|3|凡大祭司都是為獻禮物和祭物設立的，所以這位大祭司也必須有所獻上。
HEB|8|4|他若在地上，就不用作祭司，因為已經有照律法獻禮物的祭司了。
HEB|8|5|他們所供奉的本是天上之事的樣式和影像，正如 摩西 將要造帳幕的時候，上帝警戒他，說：「要謹慎，一切都要照著在山上指示你的樣式去做。」
HEB|8|6|如今耶穌已經得了更優越的事奉，正如他作更美之約的中保；這約原是憑更美之應許立的。
HEB|8|7|第一個約若沒有瑕疵，就無須尋求第二個約了。
HEB|8|8|所以上帝指責他們說： 「主說，看哪，日子將到， 我要與 以色列 家 和 猶大 家另立新的約；
HEB|8|9|不像我拉著他們祖宗的手 領他們出 埃及 地的時候， 與他們所立的約； 因為他們不恆心守我的約， 所以我也不理他們；這是主說的。
HEB|8|10|主又說： 那些日子以後， 我與 以色列 家所立的約是這樣： 我要將我的律法放在他們的心思裏， 寫在他們的心上； 我要作他們的上帝， 他們要作我的子民。
HEB|8|11|他們各人不用教導自己的鄉親和自己的弟兄，說：你要認識主； 因為從最小的到最大的， 他們都要認識我。
HEB|8|12|我要寬恕他們的不義， 絕不再記得他們的罪惡。」
HEB|8|13|既然上帝提到「新的約」，那麼第一個約就成為舊的了；而那漸舊漸衰的必然很快消逝了。
HEB|9|1|原來連第一個約都有敬拜的禮儀和屬世界的聖幕。
HEB|9|2|因為那預備好了的帳幕，第一層叫聖所，裏面有燈臺、供桌和供餅。
HEB|9|3|第二層幔子後又有一層帳幕，叫至聖所，
HEB|9|4|有金香壇和四周包金的約櫃，櫃裏有盛嗎哪的金罐、 亞倫 那根發過芽的杖和兩塊約版；
HEB|9|5|櫃上面有榮耀的基路伯罩著施恩座。有關這一切我現在不能一一細說。
HEB|9|6|這些物件既如此預備齊了，眾祭司就不斷地進第一層帳幕行拜上帝的禮。
HEB|9|7|至於第二層帳幕，惟有大祭司一年一次獨自進去，沒有一次不帶著血，為自己獻上，也為百姓無意所犯的過錯獻上。
HEB|9|8|聖靈藉此指明，第一層帳幕仍存在的時候，進入至聖所的路還沒有顯示。
HEB|9|9|那第一層帳幕是現今時代的一個預表，表示所獻的禮物和祭物都不能使敬拜的人在良心上得以完全。
HEB|9|10|這些事只不過是有關飲食和各種潔淨的規矩，是屬肉體的條例，它的功效是直到新次序的時期來到為止。
HEB|9|11|但現在基督已經來到，作了已實現的美事的大祭司，經過那更大更全備的帳幕，不是人手所造，也不是屬於這世界的；
HEB|9|12|他不用山羊和牛犢的血，而是用自己的血，只一次進入至聖所就獲得了永遠的贖罪。
HEB|9|13|若山羊和公牛的血，以及母牛犢的灰，灑在不潔的人身上，尚且使人成聖，身體潔淨，
HEB|9|14|何況基督的血，他藉著永遠的靈把自己無瑕疵地獻給上帝，更能洗淨我們 的良心，除去致死的行為，好事奉那位永生的上帝。
HEB|9|15|為此，基督作了新約的中保；因為他的死，贖了人在第一個約之時所犯的罪過，使蒙召的人能得著所應許永遠的產業。
HEB|9|16|凡有遺囑，必須證實立遺囑的人已經死了。
HEB|9|17|因為人死了，遺囑才有效力；立遺囑的人尚在，遺囑就不能生效。
HEB|9|18|所以，第一個約也是用血立的。
HEB|9|19|因為 摩西 當日照著律法將各樣誡命傳給眾百姓，就拿朱紅色絨和牛膝草，把牛犢、山羊 的血和水灑在書上，又灑在眾百姓身上，
HEB|9|20|說：「這血就是上帝與你們立約的憑據。」
HEB|9|21|他又照樣把血灑在帳幕和敬拜用的各樣器皿上。
HEB|9|22|按著律法，幾乎每樣東西都是用血潔淨的；沒有流血，就沒有赦罪。
HEB|9|23|這樣，照著天上樣式做的物件必須用這些禮儀去潔淨，但那天上的一切，自然當用更美的祭物去潔淨。
HEB|9|24|因為基督並沒有進了人手所造的聖所—這不過是真聖所的影像—而是進到天上，如今為我們出現在上帝面前。
HEB|9|25|他也無須多次將自己獻上，像大祭司每年帶著牛羊的血進入至聖所。
HEB|9|26|如果這樣，他從創世以來就必須多次受苦了。但如今，他在今世的末期顯現，僅一次把自己獻為祭，好除掉罪。
HEB|9|27|按著命定，人人都有一死，死後且有審判。
HEB|9|28|同樣，基督既然一次獻上，擔當了許多人的罪，將來要第二次顯現，與罪無關，而是為了拯救熱切等候他的人。
HEB|10|1|既然律法只不過是未來美好事物的影子，不是本體的真像，就不能藉著每年常獻一樣的祭物，使那些進前來的人完全。
HEB|10|2|若不然，獻祭的事豈不早已停止了嗎？因為敬拜的人僅只一次潔淨，良心就不再覺得有罪了。
HEB|10|3|但是這些祭物使人每年都想起罪來，
HEB|10|4|因為公牛和山羊的血不能除罪。
HEB|10|5|所以，基督到世上來的時候，就說： 「祭物和禮物不是你所要的， 但你曾給我預備了身體。
HEB|10|6|燔祭和贖罪祭 是你不喜歡的。
HEB|10|7|那時我說： 看哪！我來了，我的事在經卷上已經記載了； 上帝啊！我來為要照你的旨意行。」
HEB|10|8|以上說：「祭物和禮物，以及燔祭和贖罪祭，不是你所要的，也不是你喜歡的。」這都是按著律法獻的。
HEB|10|9|他接著說：「看哪！我來了，為要照你的旨意行。」可見他除去在先的，為要立定在後的。
HEB|10|10|我們憑著這旨意，藉著耶穌基督，僅只一次獻上他的身體就得以成聖。
HEB|10|11|所有的祭司天天站著事奉上帝，屢次獻上一樣的祭物，這祭物永不能除罪。
HEB|10|12|但基督獻了一次永遠有效的贖罪祭，就坐在上帝的右邊，
HEB|10|13|從此等候他的仇敵成為他的腳凳。
HEB|10|14|因為他僅只一次獻祭，就使那些得以成聖的人永遠完全。
HEB|10|15|聖靈也對我們作證，因為他說過：
HEB|10|16|「主說：那些日子以後， 我與他們所立的約是這樣的： 我要將我的律法放在他們的心上， 又要寫在他們的心思裏。」
HEB|10|17|並說： 「他們的罪惡和他們的過犯， 我絕不再記得。」
HEB|10|18|這些罪過既已蒙赦免，就不用再為罪獻祭了。
HEB|10|19|所以，弟兄們，既然我們靠著耶穌的血得以坦然進入至聖所，
HEB|10|20|是藉著他給我們開了一條又新又活的路，從幔子經過，這幔子就是他的身體。
HEB|10|21|既然我們有一位偉大祭司治理上帝的家，
HEB|10|22|那麼，我們該用誠心和充足的信心，同已蒙潔淨、無虧的良心，和清水洗淨了的身體來親近上帝。
HEB|10|23|我們要堅守所宣認的指望，毫不動搖，因為應許我們的那位是信實的。
HEB|10|24|我們要彼此相顧，激發愛心，勉勵行善；
HEB|10|25|不可停止聚會，好像那些停止慣了的人，倒要彼此勸勉，既然知道那日子臨近，就更當如此。
HEB|10|26|如果我們領受真理的知識以後仍故意犯罪，就不再有贖罪的祭物，
HEB|10|27|惟有戰戰兢兢等候審判和那將吞滅眾敵人的烈火了。
HEB|10|28|任何人干犯 摩西 的律法，憑兩個或三個證人，尚且必須處死，不得寬赦，
HEB|10|29|更何況踐踏上帝兒子的人，他們將那使他成聖之約的血當作不潔淨，又褻慢施恩的聖靈的人，你們想，他不該受更嚴厲的懲罰嗎？
HEB|10|30|因為我們知道誰說： 「伸冤在我， 我必報應。」 又說： 「主要審判他的百姓。」
HEB|10|31|落在永生上帝的手裏真是可怕呀！
HEB|10|32|你們要追念往日；你們蒙了光照以後，忍受了許多痛苦的掙扎：
HEB|10|33|一面在眾人面前公然被毀謗，遭患難；一面陪伴那些受這樣苦難的人。
HEB|10|34|你們同情那些遭監禁的人，也欣然忍受你們的家業被人搶去，因為你們知道自己有更美好更長存的家業。
HEB|10|35|所以，不可丟棄你們無懼的心，存這樣的心必得大賞賜。
HEB|10|36|你們必須忍耐，使你們行完了上帝的旨意，可以獲得所應許的。
HEB|10|37|因為 「還有一點點時候， 那要來的就來，必不遲延。
HEB|10|38|只是我的義人必因信得生； 他若退縮，我心就不喜歡他。」
HEB|10|39|我們卻不是退縮以致沉淪的那等人，而是有信心以致得生命的人。
HEB|11|1|信就是對所盼望之事有把握，對未見之事有確據。
HEB|11|2|古人因著這信獲得了讚許。
HEB|11|3|因著信，我們知道這宇宙是藉上帝的話造成的。這樣，看得見的是從看不見的造出來的。
HEB|11|4|因著信， 亞伯 獻祭給上帝比 該隱 所獻的更美，因此獲得了讚許為義人，上帝親自悅納了他的禮物。他雖然死了，卻因這信仍舊在說話。
HEB|11|5|因著信， 以諾 被接去，得以不見死，人也找不著他，因為上帝已經把他接去了；只是他被接去以前，已討得上帝的喜悅而蒙讚許。
HEB|11|6|沒有信，就不能討上帝的喜悅，因為到上帝面前來的人必須信有上帝，並且信他會賞賜尋求他的人。
HEB|11|7|因著信， 挪亞 既蒙上帝指示他未見的事，動了敬畏的心，造了方舟，使他全家得救。藉此他定了那世代的罪，自己也承受了那從信而來的義。
HEB|11|8|因著信， 亞伯拉罕 蒙召的時候就遵命出去，往將來要承受為基業的地方去；他出去的時候還不知往哪裏去。
HEB|11|9|因著信，他就在所應許之地作客，好像在異鄉，居住在帳棚裏，與蒙同一個應許的 以撒 和 雅各 一樣。
HEB|11|10|因為他等候著那座有根基的城，就是上帝所設計和建造的。
HEB|11|11|因著信， 撒拉 自己已過了生育的年齡還能懷孕，因為她認為應許她的那位是可信的 ；
HEB|11|12|所以，從一個彷彿已死的人竟生出子孫，如同天上的星那樣眾多，海邊的沙那樣無數。
HEB|11|13|這些人都是存著信心死的，並沒有得著所應許的，卻從遠處觀望，且歡喜迎接。他們承認自己在地上是客旅，是寄居的。
HEB|11|14|說這樣話的人是表明自己要尋找一個家鄉。
HEB|11|15|他們若想念所離開的家鄉，還有回去的機會。
HEB|11|16|其實他們所羨慕的是一個更美的，就是在天上的家鄉。所以，上帝並不因他們稱他為上帝 而覺得羞恥，因為他已經為他們預備了一座城。
HEB|11|17|因著信， 亞伯拉罕 被考驗的時候把 以撒 獻上，這就是那領受了應許的人甘心把自己獨生的兒子獻上。
HEB|11|18|論到這兒子，上帝曾說：「從 以撒 生的才要稱為你的後裔。」
HEB|11|19|他認為上帝甚至能使人從死人中復活，意味著他得回了他的兒子。
HEB|11|20|因著信， 以撒 指著將來的事給 雅各 、 以掃 祝福。
HEB|11|21|因著信， 雅各 臨死的時候給 約瑟 的兩個兒子個別祝福，扶著枴杖敬拜上帝。
HEB|11|22|因著信， 約瑟 臨終的時候提到 以色列 人將來要出 埃及 ，並為自己的骸骨留下遺言。
HEB|11|23|因著信， 摩西 生下來，他的父母見他是個俊美的孩子，把他藏了三個月，並不怕王的命令。
HEB|11|24|因著信， 摩西 長大了不肯稱為法老女兒之子。
HEB|11|25|他寧可和上帝的百姓一同受苦，也不願在罪中享受片刻的歡樂。
HEB|11|26|他把為彌賽亞受凌辱看得比 埃及 的財物更寶貴，因為他想望所要得的賞賜。
HEB|11|27|因著信，他離開 埃及 ，不怕王的憤怒，因為他恆心忍耐，如同看見那不能看見的上帝。
HEB|11|28|因著信，他設立逾越節，在門上灑血，免得那毀滅者加害 以色列 人的長子。
HEB|11|29|因著信，他們過 紅海 如行乾地； 埃及 人試著要過去就被淹沒了。
HEB|11|30|因著信， 以色列 人圍繞 耶利哥城 七日，城牆就倒塌了。
HEB|11|31|因著信，妓女 喇合 曾友善地接待探子，就沒有跟那些不順從的人一同滅亡。
HEB|11|32|我還要說甚麼呢？若要一一細說 基甸 、 巴拉 、 參孫 、 耶弗他 、 大衛 、 撒母耳 和眾先知的事，時間就不夠了。
HEB|11|33|他們藉著信，制伏了敵國，行了公義，得了應許，堵住了獅子的口，
HEB|11|34|滅了烈火的威力，在鋒利的刀劍下逃生，從軟弱變為剛強，爭戰中顯出勇猛，打退外邦的全軍。
HEB|11|35|有些婦人得回從死人中復活的親人。又有人忍受嚴刑，拒絕被釋放，為要得著更美好的復活。
HEB|11|36|又有人忍受戲弄、鞭打、捆鎖、監禁、各等的磨煉；
HEB|11|37|他們被石頭打死，被鋸鋸死， 被刀殺，披著綿羊山羊的皮各處奔跑，受貧窮、患難、虐待。
HEB|11|38|這世界配不上他們，他們在曠野、山嶺、山洞、地穴，飄流無定。
HEB|11|39|這些人都是因信獲得了讚許，卻仍未得著所應許的，
HEB|11|40|因為上帝給我們預備了更美好的事，若沒有我們，他們就不能達到完全。
HEB|12|1|所以，既然我們有這許多見證人如同雲彩圍繞著我們，就該卸下各樣重擔和緊緊纏累的罪，以堅忍的心奔那擺在我們前頭的路程，
HEB|12|2|仰望我們信心的創始成終者耶穌，他因那擺在前面的喜樂，輕看羞辱，忍受了十字架的苦難，如今已坐在上帝寶座的右邊。
HEB|12|3|你們要仔細想想這位忍受了罪人如此頂撞的耶穌，你們就不致心灰意懶了。
HEB|12|4|你們與罪惡爭鬥，還沒有抵抗到流血的地步。
HEB|12|5|你們又忘了上帝勸你們如同勸兒女的那些話，說： 「我兒啊，不可輕看主的管教， 被他責備的時候不可灰心；
HEB|12|6|因為主所愛的，他必管教， 又鞭打他所接納的每一個孩子。」
HEB|12|7|為了受管教，你們要忍受。上帝待你們如同待兒女。哪有兒女不被父親管教的呢？
HEB|12|8|管教原是眾兒女共同所領受的；你們若不受管教，就是私生子，不是兒女了。
HEB|12|9|再者，我們曾有肉身之父管教我們，我們尚且敬重他，何況靈性之父，我們豈不更當順服他而得生命嗎？
HEB|12|10|肉身之父都是短時間隨己意管教我們，惟有靈性之父管教我們是要我們得益處，使我們在他的聖潔上有份。
HEB|12|11|凡管教的事，當時不覺得快樂，反覺得痛苦；後來卻為那經過鍛鍊的人結出平安的果子，就是義的果子。
HEB|12|12|所以，你們要把下垂的手舉起來，發酸的腿挺直；
HEB|12|13|要為自己的腳把道路修直了，使瘸了的腿不再脫臼，反而得到痊癒。
HEB|12|14|你們要追求與眾人和睦，並要追求聖潔；人非聖潔不能見主。
HEB|12|15|要謹慎，免得有人失去了上帝的恩典；免得有毒根生出來擾亂你們，因而使許多人沾染污穢，
HEB|12|16|免得有人淫亂，或不敬虔如 以掃 ，他因一點點食物把自己長子的名分賣了。
HEB|12|17|後來你們知道，他想要承受父親的祝福，竟被拒絕，雖然流著淚苦求，卻得不著門路使他父親回心轉意。
HEB|12|18|你們不是來到那可觸摸的山，那裏有火焰、密雲、黑暗、暴風、
HEB|12|19|角聲，和說話的聲音；當時那些聽見這聲音的，都求不要再向他們說話，
HEB|12|20|因為他們擔當不起所命令他們的話，說：「靠近這山的，即使是走獸，也要用石頭打死。」
HEB|12|21|所見的景象極其可怕，以致 摩西 說：「我恐懼戰兢。」
HEB|12|22|但是你們是來到 錫安山 ，永生上帝的城，就是天上的 耶路撒冷 ，那裏有千千萬萬的天使，
HEB|12|23|有名字記錄在天上眾長子的盛會，有審判眾人的上帝和成為完全的義人的靈魂，
HEB|12|24|並新約的中保耶穌，以及所灑的血；這血所說的信息比 亞伯 的血所說的更美。
HEB|12|25|你們總要謹慎，不可拒絕那向你們說話的，因為那些拒絕了在地上警戒他們的，尚且不能逃罪，何況我們違背那從天上警戒我們的呢？
HEB|12|26|當時他的聲音震動了地，但如今他應許說：「再一次我不單要震動地，還要震動天。」
HEB|12|27|這「再一次」的話是指明被震動的要像受造之物一樣被挪去，使那不被震動的能常存。
HEB|12|28|所以，既然我們得了不能被震動的國度，就要感恩，照著上帝所喜悅的，用虔誠、敬畏的心事奉上帝，
HEB|12|29|因為我們的上帝是吞滅的火。
HEB|13|1|你們務要常存弟兄相愛的心。
HEB|13|2|不可忘記用愛心接待旅客，因為曾經有人這樣做，在無意中接待了天使。
HEB|13|3|要記念受監禁的人，好像與他們同受監禁；要記念受虐待的人，好像你們也親身受虐待一樣。
HEB|13|4|婚姻，人人都當尊重，共眠的床也不可污穢，因為淫亂和通姦的人，上帝必審判。
HEB|13|5|不可貪愛錢財，要以自己所有的為滿足，因為上帝曾說：「我絕不撇下你，也絕不丟棄你。」
HEB|13|6|所以，我們可以勇敢地說： 「主是我的幫助， 我必不懼怕。 人能把我怎麼樣呢？」
HEB|13|7|從前引導你們、傳上帝的道給你們的人，你們要記念他們，效法他們的信心，回顧他們為人的結局。
HEB|13|8|耶穌基督昨日、今日，一直到永遠，是一樣的。
HEB|13|9|你們不要被種種怪異的教訓勾引了去，因為人的心靠恩典得堅固才是好的，並不是靠飲食。那在飲食上用心的，從來沒有得到益處。
HEB|13|10|我們有一祭壇，上面的祭物是那些在會幕中供職的人無權可吃的。
HEB|13|11|因為牲畜的血被大祭司帶入至聖所作贖罪祭，牲畜的體卻在營外燒掉。
HEB|13|12|所以，耶穌也在城門外受苦，為要用自己的血使百姓成聖。
HEB|13|13|這樣，我們也當走出營外，到他那裏去，忍受他所受的凌辱。
HEB|13|14|在這裏，我們本沒有永存的城，而是在尋求那將要來的城。
HEB|13|15|我們應當藉著耶穌，常常以頌讚為祭獻給上帝，這是那宣認他名的人嘴唇所結的果子。
HEB|13|16|只是不可忘記行善和分享，因為這樣的祭物是上帝所喜悅的。
HEB|13|17|你們要服從那些引導你們的，並且要順服，因為他們為你們的靈魂時刻警醒，像在上帝面前交賬的人，讓他們在交賬的時候有喜樂，而不是嘆息，嘆息就對你們無益了。
HEB|13|18|請你們為我們禱告；因為我們自覺良心無虧，願意凡事按正道而行。
HEB|13|19|我更求你們為我禱告，使我快些回到你們那裏去。
HEB|13|20|但願賜平安 的上帝，就是那憑永約之血，把群羊的大牧人—我們主耶穌從死人中領出來的上帝，
HEB|13|21|在各樣善事上裝備你們，使你們遵行他的旨意；又藉著耶穌基督在我們 裏面行他所喜悅的事。願榮耀歸給他，直到永永遠遠 。阿們！
HEB|13|22|弟兄們，我簡略地寫信給你們，希望你們聽我勸勉的話。
HEB|13|23|你們該知道，我們的弟兄 提摩太 已經重獲自由了；他若很快就來，我必同他去見你們。
HEB|13|24|請你們向帶領你們的諸位和眾聖徒問安。從 意大利 來的人也向你們問安。
HEB|13|25|願恩惠與你們眾人同在。
