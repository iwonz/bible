NEH|1|1|The words of Nehemiah son of Hacaliah: In the month of Kislev in the twentieth year, while I was in the citadel of Susa,
NEH|1|2|Hanani, one of my brothers, came from Judah with some other men, and I questioned them about the Jewish remnant that survived the exile, and also about Jerusalem.
NEH|1|3|They said to me, "Those who survived the exile and are back in the province are in great trouble and disgrace. The wall of Jerusalem is broken down, and its gates have been burned with fire."
NEH|1|4|When I heard these things, I sat down and wept. For some days I mourned and fasted and prayed before the God of heaven.
NEH|1|5|Then I said: "O LORD, God of heaven, the great and awesome God, who keeps his covenant of love with those who love him and obey his commands,
NEH|1|6|let your ear be attentive and your eyes open to hear the prayer your servant is praying before you day and night for your servants, the people of Israel. I confess the sins we Israelites, including myself and my father's house, have committed against you.
NEH|1|7|We have acted very wickedly toward you. We have not obeyed the commands, decrees and laws you gave your servant Moses.
NEH|1|8|"Remember the instruction you gave your servant Moses, saying, 'If you are unfaithful, I will scatter you among the nations,
NEH|1|9|but if you return to me and obey my commands, then even if your exiled people are at the farthest horizon, I will gather them from there and bring them to the place I have chosen as a dwelling for my Name.'
NEH|1|10|"They are your servants and your people, whom you redeemed by your great strength and your mighty hand.
NEH|1|11|O Lord, let your ear be attentive to the prayer of this your servant and to the prayer of your servants who delight in revering your name. Give your servant success today by granting him favor in the presence of this man." I was cupbearer to the king.
NEH|2|1|In the month of Nisan in the twentieth year of King Artaxerxes, when wine was brought for him, I took the wine and gave it to the king. I had not been sad in his presence before;
NEH|2|2|so the king asked me, "Why does your face look so sad when you are not ill? This can be nothing but sadness of heart." I was very much afraid,
NEH|2|3|but I said to the king, "May the king live forever! Why should my face not look sad when the city where my fathers are buried lies in ruins, and its gates have been destroyed by fire?"
NEH|2|4|The king said to me, "What is it you want?" Then I prayed to the God of heaven,
NEH|2|5|and I answered the king, "If it pleases the king and if your servant has found favor in his sight, let him send me to the city in Judah where my fathers are buried so that I can rebuild it."
NEH|2|6|Then the king, with the queen sitting beside him, asked me, "How long will your journey take, and when will you get back?" It pleased the king to send me; so I set a time.
NEH|2|7|I also said to him, "If it pleases the king, may I have letters to the governors of Trans-Euphrates, so that they will provide me safe-conduct until I arrive in Judah?
NEH|2|8|And may I have a letter to Asaph, keeper of the king's forest, so he will give me timber to make beams for the gates of the citadel by the temple and for the city wall and for the residence I will occupy?" And because the gracious hand of my God was upon me, the king granted my requests.
NEH|2|9|So I went to the governors of Trans-Euphrates and gave them the king's letters. The king had also sent army officers and cavalry with me.
NEH|2|10|When Sanballat the Horonite and Tobiah the Ammonite official heard about this, they were very much disturbed that someone had come to promote the welfare of the Israelites.
NEH|2|11|I went to Jerusalem, and after staying there three days
NEH|2|12|I set out during the night with a few men. I had not told anyone what my God had put in my heart to do for Jerusalem. There were no mounts with me except the one I was riding on.
NEH|2|13|By night I went out through the Valley Gate toward the Jackal Well and the Dung Gate, examining the walls of Jerusalem, which had been broken down, and its gates, which had been destroyed by fire.
NEH|2|14|Then I moved on toward the Fountain Gate and the King's Pool, but there was not enough room for my mount to get through;
NEH|2|15|so I went up the valley by night, examining the wall. Finally, I turned back and reentered through the Valley Gate.
NEH|2|16|The officials did not know where I had gone or what I was doing, because as yet I had said nothing to the Jews or the priests or nobles or officials or any others who would be doing the work.
NEH|2|17|Then I said to them, "You see the trouble we are in: Jerusalem lies in ruins, and its gates have been burned with fire. Come, let us rebuild the wall of Jerusalem, and we will no longer be in disgrace."
NEH|2|18|I also told them about the gracious hand of my God upon me and what the king had said to me. They replied, "Let us start rebuilding." So they began this good work.
NEH|2|19|But when Sanballat the Horonite, Tobiah the Ammonite official and Geshem the Arab heard about it, they mocked and ridiculed us. "What is this you are doing?" they asked. "Are you rebelling against the king?"
NEH|2|20|I answered them by saying, "The God of heaven will give us success. We his servants will start rebuilding, but as for you, you have no share in Jerusalem or any claim or historic right to it."
NEH|3|1|Eliashib the high priest and his fellow priests went to work and rebuilt the Sheep Gate. They dedicated it and set its doors in place, building as far as the Tower of the Hundred, which they dedicated, and as far as the Tower of Hananel.
NEH|3|2|The men of Jericho built the adjoining section, and Zaccur son of Imri built next to them.
NEH|3|3|The Fish Gate was rebuilt by the sons of Hassenaah. They laid its beams and put its doors and bolts and bars in place.
NEH|3|4|Meremoth son of Uriah, the son of Hakkoz, repaired the next section. Next to him Meshullam son of Berekiah, the son of Meshezabel, made repairs, and next to him Zadok son of Baana also made repairs.
NEH|3|5|The next section was repaired by the men of Tekoa, but their nobles would not put their shoulders to the work under their supervisors.
NEH|3|6|The Jeshanah Gate was repaired by Joiada son of Paseah and Meshullam son of Besodeiah. They laid its beams and put its doors and bolts and bars in place.
NEH|3|7|Next to them, repairs were made by men from Gibeon and Mizpah-Melatiah of Gibeon and Jadon of Meronoth-places under the authority of the governor of Trans-Euphrates.
NEH|3|8|Uzziel son of Harhaiah, one of the goldsmiths, repaired the next section; and Hananiah, one of the perfume-makers, made repairs next to that. They restored Jerusalem as far as the Broad Wall.
NEH|3|9|Rephaiah son of Hur, ruler of a half-district of Jerusalem, repaired the next section.
NEH|3|10|Adjoining this, Jedaiah son of Harumaph made repairs opposite his house, and Hattush son of Hashabneiah made repairs next to him.
NEH|3|11|Malkijah son of Harim and Hasshub son of Pahath-Moab repaired another section and the Tower of the Ovens.
NEH|3|12|Shallum son of Hallohesh, ruler of a half-district of Jerusalem, repaired the next section with the help of his daughters.
NEH|3|13|The Valley Gate was repaired by Hanun and the residents of Zanoah. They rebuilt it and put its doors and bolts and bars in place. They also repaired five hundred yards of the wall as far as the Dung Gate.
NEH|3|14|The Dung Gate was repaired by Malkijah son of Recab, ruler of the district of Beth Hakkerem. He rebuilt it and put its doors and bolts and bars in place.
NEH|3|15|The Fountain Gate was repaired by Shallun son of Col-Hozeh, ruler of the district of Mizpah. He rebuilt it, roofing it over and putting its doors and bolts and bars in place. He also repaired the wall of the Pool of Siloam, by the King's Garden, as far as the steps going down from the City of David.
NEH|3|16|Beyond him, Nehemiah son of Azbuk, ruler of a half-district of Beth Zur, made repairs up to a point opposite the tombs of David, as far as the artificial pool and the House of the Heroes.
NEH|3|17|Next to him, the repairs were made by the Levites under Rehum son of Bani. Beside him, Hashabiah, ruler of half the district of Keilah, carried out repairs for his district.
NEH|3|18|Next to him, the repairs were made by their countrymen under Binnui son of Henadad, ruler of the other half-district of Keilah.
NEH|3|19|Next to him, Ezer son of Jeshua, ruler of Mizpah, repaired another section, from a point facing the ascent to the armory as far as the angle.
NEH|3|20|Next to him, Baruch son of Zabbai zealously repaired another section, from the angle to the entrance of the house of Eliashib the high priest.
NEH|3|21|Next to him, Meremoth son of Uriah, the son of Hakkoz, repaired another section, from the entrance of Eliashib's house to the end of it.
NEH|3|22|The repairs next to him were made by the priests from the surrounding region.
NEH|3|23|Beyond them, Benjamin and Hasshub made repairs in front of their house; and next to them, Azariah son of Maaseiah, the son of Ananiah, made repairs beside his house.
NEH|3|24|Next to him, Binnui son of Henadad repaired another section, from Azariah's house to the angle and the corner,
NEH|3|25|and Palal son of Uzai worked opposite the angle and the tower projecting from the upper palace near the court of the guard. Next to him, Pedaiah son of Parosh
NEH|3|26|and the temple servants living on the hill of Ophel made repairs up to a point opposite the Water Gate toward the east and the projecting tower.
NEH|3|27|Next to them, the men of Tekoa repaired another section, from the great projecting tower to the wall of Ophel.
NEH|3|28|Above the Horse Gate, the priests made repairs, each in front of his own house.
NEH|3|29|Next to them, Zadok son of Immer made repairs opposite his house. Next to him, Shemaiah son of Shecaniah, the guard at the East Gate, made repairs.
NEH|3|30|Next to him, Hananiah son of Shelemiah, and Hanun, the sixth son of Zalaph, repaired another section. Next to them, Meshullam son of Berekiah made repairs opposite his living quarters.
NEH|3|31|Next to him, Malkijah, one of the goldsmiths, made repairs as far as the house of the temple servants and the merchants, opposite the Inspection Gate, and as far as the room above the corner;
NEH|3|32|and between the room above the corner and the Sheep Gate the goldsmiths and merchants made repairs.
NEH|4|1|When Sanballat heard that we were rebuilding the wall, he became angry and was greatly incensed. He ridiculed the Jews,
NEH|4|2|and in the presence of his associates and the army of Samaria, he said, "What are those feeble Jews doing? Will they restore their wall? Will they offer sacrifices? Will they finish in a day? Can they bring the stones back to life from those heaps of rubble-burned as they are?"
NEH|4|3|Tobiah the Ammonite, who was at his side, said, "What they are building-if even a fox climbed up on it, he would break down their wall of stones!"
NEH|4|4|Hear us, O our God, for we are despised. Turn their insults back on their own heads. Give them over as plunder in a land of captivity.
NEH|4|5|Do not cover up their guilt or blot out their sins from your sight, for they have thrown insults in the face of the builders.
NEH|4|6|So we rebuilt the wall till all of it reached half its height, for the people worked with all their heart.
NEH|4|7|But when Sanballat, Tobiah, the Arabs, the Ammonites and the men of Ashdod heard that the repairs to Jerusalem's walls had gone ahead and that the gaps were being closed, they were very angry.
NEH|4|8|They all plotted together to come and fight against Jerusalem and stir up trouble against it.
NEH|4|9|But we prayed to our God and posted a guard day and night to meet this threat.
NEH|4|10|Meanwhile, the people in Judah said, "The strength of the laborers is giving out, and there is so much rubble that we cannot rebuild the wall."
NEH|4|11|Also our enemies said, "Before they know it or see us, we will be right there among them and will kill them and put an end to the work."
NEH|4|12|Then the Jews who lived near them came and told us ten times over, "Wherever you turn, they will attack us."
NEH|4|13|Therefore I stationed some of the people behind the lowest points of the wall at the exposed places, posting them by families, with their swords, spears and bows.
NEH|4|14|After I looked things over, I stood up and said to the nobles, the officials and the rest of the people, "Don't be afraid of them. Remember the Lord, who is great and awesome, and fight for your brothers, your sons and your daughters, your wives and your homes."
NEH|4|15|When our enemies heard that we were aware of their plot and that God had frustrated it, we all returned to the wall, each to his own work.
NEH|4|16|From that day on, half of my men did the work, while the other half were equipped with spears, shields, bows and armor. The officers posted themselves behind all the people of Judah
NEH|4|17|who were building the wall. Those who carried materials did their work with one hand and held a weapon in the other,
NEH|4|18|and each of the builders wore his sword at his side as he worked. But the man who sounded the trumpet stayed with me.
NEH|4|19|Then I said to the nobles, the officials and the rest of the people, "The work is extensive and spread out, and we are widely separated from each other along the wall.
NEH|4|20|Wherever you hear the sound of the trumpet, join us there. Our God will fight for us!"
NEH|4|21|So we continued the work with half the men holding spears, from the first light of dawn till the stars came out.
NEH|4|22|At that time I also said to the people, "Have every man and his helper stay inside Jerusalem at night, so they can serve us as guards by night and workmen by day."
NEH|4|23|Neither I nor my brothers nor my men nor the guards with me took off our clothes; each had his weapon, even when he went for water.
NEH|5|1|Now the men and their wives raised a great outcry against their Jewish brothers.
NEH|5|2|Some were saying, "We and our sons and daughters are numerous; in order for us to eat and stay alive, we must get grain."
NEH|5|3|Others were saying, "We are mortgaging our fields, our vineyards and our homes to get grain during the famine."
NEH|5|4|Still others were saying, "We have had to borrow money to pay the king's tax on our fields and vineyards.
NEH|5|5|Although we are of the same flesh and blood as our countrymen and though our sons are as good as theirs, yet we have to subject our sons and daughters to slavery. Some of our daughters have already been enslaved, but we are powerless, because our fields and our vineyards belong to others."
NEH|5|6|When I heard their outcry and these charges, I was very angry.
NEH|5|7|I pondered them in my mind and then accused the nobles and officials. I told them, "You are exacting usury from your own countrymen!" So I called together a large meeting to deal with them
NEH|5|8|and said: "As far as possible, we have bought back our Jewish brothers who were sold to the Gentiles. Now you are selling your brothers, only for them to be sold back to us!" They kept quiet, because they could find nothing to say.
NEH|5|9|So I continued, "What you are doing is not right. Shouldn't you walk in the fear of our God to avoid the reproach of our Gentile enemies?
NEH|5|10|I and my brothers and my men are also lending the people money and grain. But let the exacting of usury stop!
NEH|5|11|Give back to them immediately their fields, vineyards, olive groves and houses, and also the usury you are charging them-the hundredth part of the money, grain, new wine and oil."
NEH|5|12|"We will give it back," they said. "And we will not demand anything more from them. We will do as you say." Then I summoned the priests and made the nobles and officials take an oath to do what they had promised.
NEH|5|13|I also shook out the folds of my robe and said, "In this way may God shake out of his house and possessions every man who does not keep this promise. So may such a man be shaken out and emptied!" At this the whole assembly said, "Amen," and praised the LORD. And the people did as they had promised.
NEH|5|14|Moreover, from the twentieth year of King Artaxerxes, when I was appointed to be their governor in the land of Judah, until his thirty-second year-twelve years-neither I nor my brothers ate the food allotted to the governor.
NEH|5|15|But the earlier governors-those preceding me-placed a heavy burden on the people and took forty shekels of silver from them in addition to food and wine. Their assistants also lorded it over the people. But out of reverence for God I did not act like that.
NEH|5|16|Instead, I devoted myself to the work on this wall. All my men were assembled there for the work; we did not acquire any land.
NEH|5|17|Furthermore, a hundred and fifty Jews and officials ate at my table, as well as those who came to us from the surrounding nations.
NEH|5|18|Each day one ox, six choice sheep and some poultry were prepared for me, and every ten days an abundant supply of wine of all kinds. In spite of all this, I never demanded the food allotted to the governor, because the demands were heavy on these people.
NEH|5|19|Remember me with favor, O my God, for all I have done for these people.
NEH|6|1|When word came to Sanballat, Tobiah, Geshem the Arab and the rest of our enemies that I had rebuilt the wall and not a gap was left in it-though up to that time I had not set the doors in the gates-
NEH|6|2|Sanballat and Geshem sent me this message: "Come, let us meet together in one of the villages on the plain of Ono." But they were scheming to harm me;
NEH|6|3|so I sent messengers to them with this reply: "I am carrying on a great project and cannot go down. Why should the work stop while I leave it and go down to you?"
NEH|6|4|Four times they sent me the same message, and each time I gave them the same answer.
NEH|6|5|Then, the fifth time, Sanballat sent his aide to me with the same message, and in his hand was an unsealed letter
NEH|6|6|in which was written: "It is reported among the nations-and Geshem says it is true-that you and the Jews are plotting to revolt, and therefore you are building the wall. Moreover, according to these reports you are about to become their king
NEH|6|7|and have even appointed prophets to make this proclamation about you in Jerusalem: 'There is a king in Judah!' Now this report will get back to the king; so come, let us confer together."
NEH|6|8|I sent him this reply: "Nothing like what you are saying is happening; you are just making it up out of your head."
NEH|6|9|They were all trying to frighten us, thinking, "Their hands will get too weak for the work, and it will not be completed." But I prayed, "Now strengthen my hands."
NEH|6|10|One day I went to the house of Shemaiah son of Delaiah, the son of Mehetabel, who was shut in at his home. He said, "Let us meet in the house of God, inside the temple, and let us close the temple doors, because men are coming to kill you-by night they are coming to kill you."
NEH|6|11|But I said, "Should a man like me run away? Or should one like me go into the temple to save his life? I will not go!"
NEH|6|12|I realized that God had not sent him, but that he had prophesied against me because Tobiah and Sanballat had hired him.
NEH|6|13|He had been hired to intimidate me so that I would commit a sin by doing this, and then they would give me a bad name to discredit me.
NEH|6|14|Remember Tobiah and Sanballat, O my God, because of what they have done; remember also the prophetess Noadiah and the rest of the prophets who have been trying to intimidate me.
NEH|6|15|So the wall was completed on the twenty-fifth of Elul, in fifty-two days.
NEH|6|16|When all our enemies heard about this, all the surrounding nations were afraid and lost their self-confidence, because they realized that this work had been done with the help of our God.
NEH|6|17|Also, in those days the nobles of Judah were sending many letters to Tobiah, and replies from Tobiah kept coming to them.
NEH|6|18|For many in Judah were under oath to him, since he was son-in-law to Shecaniah son of Arah, and his son Jehohanan had married the daughter of Meshullam son of Berekiah.
NEH|6|19|Moreover, they kept reporting to me his good deeds and then telling him what I said. And Tobiah sent letters to intimidate me.
NEH|7|1|After the wall had been rebuilt and I had set the doors in place, the gatekeepers and the singers and the Levites were appointed.
NEH|7|2|I put in charge of Jerusalem my brother Hanani, along with Hananiah the commander of the citadel, because he was a man of integrity and feared God more than most men do.
NEH|7|3|I said to them, "The gates of Jerusalem are not to be opened until the sun is hot. While the gatekeepers are still on duty, have them shut the doors and bar them. Also appoint residents of Jerusalem as guards, some at their posts and some near their own houses."
NEH|7|4|Now the city was large and spacious, but there were few people in it, and the houses had not yet been rebuilt.
NEH|7|5|So my God put it into my heart to assemble the nobles, the officials and the common people for registration by families. I found the genealogical record of those who had been the first to return. This is what I found written there:
NEH|7|6|These are the people of the province who came up from the captivity of the exiles whom Nebuchadnezzar king of Babylon had taken captive (they returned to Jerusalem and Judah, each to his own town,
NEH|7|7|in company with Zerubbabel, Jeshua, Nehemiah, Azariah, Raamiah, Nahamani, Mordecai, Bilshan, Mispereth, Bigvai, Nehum and Baanah): The list of the men of Israel:
NEH|7|8|the descendants of Parosh 2,172
NEH|7|9|of Shephatiah 372
NEH|7|10|of Arah 652
NEH|7|11|of Pahath-Moab (through the line of Jeshua and Joab) 2,818
NEH|7|12|of Elam 1,254
NEH|7|13|of Zattu 845
NEH|7|14|of Zaccai 760
NEH|7|15|of Binnui 648
NEH|7|16|of Bebai 628
NEH|7|17|of Azgad 2,322
NEH|7|18|of Adonikam 667
NEH|7|19|of Bigvai 2,067
NEH|7|20|of Adin 655
NEH|7|21|of Ater (through Hezekiah) 98
NEH|7|22|of Hashum 328
NEH|7|23|of Bezai 324
NEH|7|24|of Hariph 112
NEH|7|25|of Gibeon 95
NEH|7|26|the men of Bethlehem and Netophah 188
NEH|7|27|of Anathoth 128
NEH|7|28|of Beth Azmaveth 42
NEH|7|29|of Kiriath Jearim, Kephirah and Beeroth 743
NEH|7|30|of Ramah and Geba 621
NEH|7|31|of Micmash 122
NEH|7|32|of Bethel and Ai 123
NEH|7|33|of the other Nebo 52
NEH|7|34|of the other Elam 1,254
NEH|7|35|of Harim 320
NEH|7|36|of Jericho 345
NEH|7|37|of Lod, Hadid and Ono 721
NEH|7|38|of Senaah 3,930
NEH|7|39|The priests: the descendants of Jedaiah (through the family of Jeshua) 973
NEH|7|40|of Immer 1,052
NEH|7|41|of Pashhur 1,247
NEH|7|42|of Harim 1,017
NEH|7|43|The Levites: the descendants of Jeshua (through Kadmiel through the line of Hodaviah) 74
NEH|7|44|The singers: the descendants of Asaph 148
NEH|7|45|The gatekeepers: the descendants of Shallum, Ater, Talmon, Akkub, Hatita and Shobai 138
NEH|7|46|The temple servants: the descendants of Ziha, Hasupha, Tabbaoth,
NEH|7|47|Keros, Sia, Padon,
NEH|7|48|Lebana, Hagaba, Shalmai,
NEH|7|49|Hanan, Giddel, Gahar,
NEH|7|50|Reaiah, Rezin, Nekoda,
NEH|7|51|Gazzam, Uzza, Paseah,
NEH|7|52|Besai, Meunim, Nephussim,
NEH|7|53|Bakbuk, Hakupha, Harhur,
NEH|7|54|Bazluth, Mehida, Harsha,
NEH|7|55|Barkos, Sisera, Temah,
NEH|7|56|Neziah and Hatipha
NEH|7|57|The descendants of the servants of Solomon: the descendants of Sotai, Sophereth, Perida,
NEH|7|58|Jaala, Darkon, Giddel,
NEH|7|59|Shephatiah, Hattil, Pokereth-Hazzebaim and Amon
NEH|7|60|The temple servants and the descendants of the servants of Solomon 392
NEH|7|61|The following came up from the towns of Tel Melah, Tel Harsha, Kerub, Addon and Immer, but they could not show that their families were descended from Israel:
NEH|7|62|the descendants of Delaiah, Tobiah and Nekoda 642
NEH|7|63|And from among the priests: the descendants of Hobaiah, Hakkoz and Barzillai (a man who had married a daughter of Barzillai the Gileadite and was called by that name).
NEH|7|64|These searched for their family records, but they could not find them and so were excluded from the priesthood as unclean.
NEH|7|65|The governor, therefore, ordered them not to eat any of the most sacred food until there should be a priest ministering with the Urim and Thummim.
NEH|7|66|The whole company numbered 42,360,
NEH|7|67|besides their 7,337 menservants and maidservants; and they also had 245 men and women singers.
NEH|7|68|There were 736 horses, 245 mules,
NEH|7|69|435 camels and 6,720 donkeys.
NEH|7|70|Some of the heads of the families contributed to the work. The governor gave to the treasury 1,000 drachmas of gold, 50 bowls and 530 garments for priests.
NEH|7|71|Some of the heads of the families gave to the treasury for the work 20,000 drachmas of gold and 2,200 minas of silver.
NEH|7|72|The total given by the rest of the people was 20,000 drachmas of gold, 2,000 minas of silver and 67 garments for priests.
NEH|7|73|The priests, the Levites, the gatekeepers, the singers and the temple servants, along with certain of the people and the rest of the Israelites, settled in their own towns. When the seventh month came and the Israelites had settled in their towns,
NEH|8|1|all the people assembled as one man in the square before the Water Gate. They told Ezra the scribe to bring out the Book of the Law of Moses, which the LORD had commanded for Israel.
NEH|8|2|So on the first day of the seventh month Ezra the priest brought the Law before the assembly, which was made up of men and women and all who were able to understand.
NEH|8|3|He read it aloud from daybreak till noon as he faced the square before the Water Gate in the presence of the men, women and others who could understand. And all the people listened attentively to the Book of the Law.
NEH|8|4|Ezra the scribe stood on a high wooden platform built for the occasion. Beside him on his right stood Mattithiah, Shema, Anaiah, Uriah, Hilkiah and Maaseiah; and on his left were Pedaiah, Mishael, Malkijah, Hashum, Hashbaddanah, Zechariah and Meshullam.
NEH|8|5|Ezra opened the book. All the people could see him because he was standing above them; and as he opened it, the people all stood up.
NEH|8|6|Ezra praised the LORD, the great God; and all the people lifted their hands and responded, "Amen! Amen!" Then they bowed down and worshiped the LORD with their faces to the ground.
NEH|8|7|The Levites-Jeshua, Bani, Sherebiah, Jamin, Akkub, Shabbethai, Hodiah, Maaseiah, Kelita, Azariah, Jozabad, Hanan and Pelaiah-instructed the people in the Law while the people were standing there.
NEH|8|8|They read from the Book of the Law of God, making it clear and giving the meaning so that the people could understand what was being read.
NEH|8|9|Then Nehemiah the governor, Ezra the priest and scribe, and the Levites who were instructing the people said to them all, "This day is sacred to the LORD your God. Do not mourn or weep." For all the people had been weeping as they listened to the words of the Law.
NEH|8|10|Nehemiah said, "Go and enjoy choice food and sweet drinks, and send some to those who have nothing prepared. This day is sacred to our Lord. Do not grieve, for the joy of the LORD is your strength."
NEH|8|11|The Levites calmed all the people, saying, "Be still, for this is a sacred day. Do not grieve."
NEH|8|12|Then all the people went away to eat and drink, to send portions of food and to celebrate with great joy, because they now understood the words that had been made known to them.
NEH|8|13|On the second day of the month, the heads of all the families, along with the priests and the Levites, gathered around Ezra the scribe to give attention to the words of the Law.
NEH|8|14|They found written in the Law, which the LORD had commanded through Moses, that the Israelites were to live in booths during the feast of the seventh month
NEH|8|15|and that they should proclaim this word and spread it throughout their towns and in Jerusalem: "Go out into the hill country and bring back branches from olive and wild olive trees, and from myrtles, palms and shade trees, to make booths"-as it is written.
NEH|8|16|So the people went out and brought back branches and built themselves booths on their own roofs, in their courtyards, in the courts of the house of God and in the square by the Water Gate and the one by the Gate of Ephraim.
NEH|8|17|The whole company that had returned from exile built booths and lived in them. From the days of Joshua son of Nun until that day, the Israelites had not celebrated it like this. And their joy was very great.
NEH|8|18|Day after day, from the first day to the last, Ezra read from the Book of the Law of God. They celebrated the feast for seven days, and on the eighth day, in accordance with the regulation, there was an assembly.
NEH|9|1|On the twenty-fourth day of the same month, the Israelites gathered together, fasting and wearing sackcloth and having dust on their heads.
NEH|9|2|Those of Israelite descent had separated themselves from all foreigners. They stood in their places and confessed their sins and the wickedness of their fathers.
NEH|9|3|They stood where they were and read from the Book of the Law of the LORD their God for a quarter of the day, and spent another quarter in confession and in worshiping the LORD their God.
NEH|9|4|Standing on the stairs were the Levites-Jeshua, Bani, Kadmiel, Shebaniah, Bunni, Sherebiah, Bani and Kenani-who called with loud voices to the LORD their God.
NEH|9|5|And the Levites-Jeshua, Kadmiel, Bani, Hashabneiah, Sherebiah, Hodiah, Shebaniah and Pethahiah-said: "Stand up and praise the LORD your God, who is from everlasting to everlasting. Blessed be your glorious name, and may it be exalted above all blessing and praise.
NEH|9|6|You alone are the LORD. You made the heavens, even the highest heavens, and all their starry host, the earth and all that is on it, the seas and all that is in them. You give life to everything, and the multitudes of heaven worship you.
NEH|9|7|"You are the LORD God, who chose Abram and brought him out of Ur of the Chaldeans and named him Abraham.
NEH|9|8|You found his heart faithful to you, and you made a covenant with him to give to his descendants the land of the Canaanites, Hittites, Amorites, Perizzites, Jebusites and Girgashites. You have kept your promise because you are righteous.
NEH|9|9|"You saw the suffering of our forefathers in Egypt; you heard their cry at the Red Sea.
NEH|9|10|You sent miraculous signs and wonders against Pharaoh, against all his officials and all the people of his land, for you knew how arrogantly the Egyptians treated them. You made a name for yourself, which remains to this day.
NEH|9|11|You divided the sea before them, so that they passed through it on dry ground, but you hurled their pursuers into the depths, like a stone into mighty waters.
NEH|9|12|By day you led them with a pillar of cloud, and by night with a pillar of fire to give them light on the way they were to take.
NEH|9|13|"You came down on Mount Sinai; you spoke to them from heaven. You gave them regulations and laws that are just and right, and decrees and commands that are good.
NEH|9|14|You made known to them your holy Sabbath and gave them commands, decrees and laws through your servant Moses.
NEH|9|15|In their hunger you gave them bread from heaven and in their thirst you brought them water from the rock; you told them to go in and take possession of the land you had sworn with uplifted hand to give them.
NEH|9|16|"But they, our forefathers, became arrogant and stiff-necked, and did not obey your commands.
NEH|9|17|They refused to listen and failed to remember the miracles you performed among them. They became stiff-necked and in their rebellion appointed a leader in order to return to their slavery. But you are a forgiving God, gracious and compassionate, slow to anger and abounding in love. Therefore you did not desert them,
NEH|9|18|even when they cast for themselves an image of a calf and said, 'This is your god, who brought you up out of Egypt,' or when they committed awful blasphemies.
NEH|9|19|"Because of your great compassion you did not abandon them in the desert. By day the pillar of cloud did not cease to guide them on their path, nor the pillar of fire by night to shine on the way they were to take.
NEH|9|20|You gave your good Spirit to instruct them. You did not withhold your manna from their mouths, and you gave them water for their thirst.
NEH|9|21|For forty years you sustained them in the desert; they lacked nothing, their clothes did not wear out nor did their feet become swollen.
NEH|9|22|"You gave them kingdoms and nations, allotting to them even the remotest frontiers. They took over the country of Sihon king of Heshbon and the country of Og king of Bashan.
NEH|9|23|You made their sons as numerous as the stars in the sky, and you brought them into the land that you told their fathers to enter and possess.
NEH|9|24|Their sons went in and took possession of the land. You subdued before them the Canaanites, who lived in the land; you handed the Canaanites over to them, along with their kings and the peoples of the land, to deal with them as they pleased.
NEH|9|25|They captured fortified cities and fertile land; they took possession of houses filled with all kinds of good things, wells already dug, vineyards, olive groves and fruit trees in abundance. They ate to the full and were well-nourished; they reveled in your great goodness.
NEH|9|26|"But they were disobedient and rebelled against you; they put your law behind their backs. They killed your prophets, who had admonished them in order to turn them back to you; they committed awful blasphemies.
NEH|9|27|So you handed them over to their enemies, who oppressed them. But when they were oppressed they cried out to you. From heaven you heard them, and in your great compassion you gave them deliverers, who rescued them from the hand of their enemies.
NEH|9|28|"But as soon as they were at rest, they again did what was evil in your sight. Then you abandoned them to the hand of their enemies so that they ruled over them. And when they cried out to you again, you heard from heaven, and in your compassion you delivered them time after time.
NEH|9|29|"You warned them to return to your law, but they became arrogant and disobeyed your commands. They sinned against your ordinances, by which a man will live if he obeys them. Stubbornly they turned their backs on you, became stiff-necked and refused to listen.
NEH|9|30|For many years you were patient with them. By your Spirit you admonished them through your prophets. Yet they paid no attention, so you handed them over to the neighboring peoples.
NEH|9|31|But in your great mercy you did not put an end to them or abandon them, for you are a gracious and merciful God.
NEH|9|32|"Now therefore, O our God, the great, mighty and awesome God, who keeps his covenant of love, do not let all this hardship seem trifling in your eyes-the hardship that has come upon us, upon our kings and leaders, upon our priests and prophets, upon our fathers and all your people, from the days of the kings of Assyria until today.
NEH|9|33|In all that has happened to us, you have been just; you have acted faithfully, while we did wrong.
NEH|9|34|Our kings, our leaders, our priests and our fathers did not follow your law; they did not pay attention to your commands or the warnings you gave them.
NEH|9|35|Even while they were in their kingdom, enjoying your great goodness to them in the spacious and fertile land you gave them, they did not serve you or turn from their evil ways.
NEH|9|36|"But see, we are slaves today, slaves in the land you gave our forefathers so they could eat its fruit and the other good things it produces.
NEH|9|37|Because of our sins, its abundant harvest goes to the kings you have placed over us. They rule over our bodies and our cattle as they please. We are in great distress.
NEH|9|38|"In view of all this, we are making a binding agreement, putting it in writing, and our leaders, our Levites and our priests are affixing their seals to it."
NEH|10|1|Those who sealed it were: Nehemiah the governor, the son of Hacaliah. Zedekiah,
NEH|10|2|Seraiah, Azariah, Jeremiah,
NEH|10|3|Pashhur, Amariah, Malkijah,
NEH|10|4|Hattush, Shebaniah, Malluch,
NEH|10|5|Harim, Meremoth, Obadiah,
NEH|10|6|Daniel, Ginnethon, Baruch,
NEH|10|7|Meshullam, Abijah, Mijamin,
NEH|10|8|Maaziah, Bilgai and Shemaiah. These were the priests.
NEH|10|9|The Levites: Jeshua son of Azaniah, Binnui of the sons of Henadad, Kadmiel,
NEH|10|10|and their associates: Shebaniah, Hodiah, Kelita, Pelaiah, Hanan,
NEH|10|11|Mica, Rehob, Hashabiah,
NEH|10|12|Zaccur, Sherebiah, Shebaniah,
NEH|10|13|Hodiah, Bani and Beninu.
NEH|10|14|The leaders of the people: Parosh, Pahath-Moab, Elam, Zattu, Bani,
NEH|10|15|Bunni, Azgad, Bebai,
NEH|10|16|Adonijah, Bigvai, Adin,
NEH|10|17|Ater, Hezekiah, Azzur,
NEH|10|18|Hodiah, Hashum, Bezai,
NEH|10|19|Hariph, Anathoth, Nebai,
NEH|10|20|Magpiash, Meshullam, Hezir,
NEH|10|21|Meshezabel, Zadok, Jaddua,
NEH|10|22|Pelatiah, Hanan, Anaiah,
NEH|10|23|Hoshea, Hananiah, Hasshub,
NEH|10|24|Hallohesh, Pilha, Shobek,
NEH|10|25|Rehum, Hashabnah, Maaseiah,
NEH|10|26|Ahiah, Hanan, Anan,
NEH|10|27|Malluch, Harim and Baanah.
NEH|10|28|"The rest of the people-priests, Levites, gatekeepers, singers, temple servants and all who separated themselves from the neighboring peoples for the sake of the Law of God, together with their wives and all their sons and daughters who are able to understand-
NEH|10|29|all these now join their brothers the nobles, and bind themselves with a curse and an oath to follow the Law of God given through Moses the servant of God and to obey carefully all the commands, regulations and decrees of the LORD our Lord.
NEH|10|30|"We promise not to give our daughters in marriage to the peoples around us or take their daughters for our sons.
NEH|10|31|"When the neighboring peoples bring merchandise or grain to sell on the Sabbath, we will not buy from them on the Sabbath or on any holy day. Every seventh year we will forgo working the land and will cancel all debts.
NEH|10|32|"We assume the responsibility for carrying out the commands to give a third of a shekel each year for the service of the house of our God:
NEH|10|33|for the bread set out on the table; for the regular grain offerings and burnt offerings; for the offerings on the Sabbaths, New Moon festivals and appointed feasts; for the holy offerings; for sin offerings to make atonement for Israel; and for all the duties of the house of our God.
NEH|10|34|"We-the priests, the Levites and the people-have cast lots to determine when each of our families is to bring to the house of our God at set times each year a contribution of wood to burn on the altar of the LORD our God, as it is written in the Law.
NEH|10|35|"We also assume responsibility for bringing to the house of the LORD each year the firstfruits of our crops and of every fruit tree.
NEH|10|36|"As it is also written in the Law, we will bring the firstborn of our sons and of our cattle, of our herds and of our flocks to the house of our God, to the priests ministering there.
NEH|10|37|"Moreover, we will bring to the storerooms of the house of our God, to the priests, the first of our ground meal, of our grain offerings, of the fruit of all our trees and of our new wine and oil. And we will bring a tithe of our crops to the Levites, for it is the Levites who collect the tithes in all the towns where we work.
NEH|10|38|A priest descended from Aaron is to accompany the Levites when they receive the tithes, and the Levites are to bring a tenth of the tithes up to the house of our God, to the storerooms of the treasury.
NEH|10|39|The people of Israel, including the Levites, are to bring their contributions of grain, new wine and oil to the storerooms where the articles for the sanctuary are kept and where the ministering priests, the gatekeepers and the singers stay. "We will not neglect the house of our God."
NEH|11|1|Now the leaders of the people settled in Jerusalem, and the rest of the people cast lots to bring one out of every ten to live in Jerusalem, the holy city, while the remaining nine were to stay in their own towns.
NEH|11|2|The people commended all the men who volunteered to live in Jerusalem.
NEH|11|3|These are the provincial leaders who settled in Jerusalem (now some Israelites, priests, Levites, temple servants and descendants of Solomon's servants lived in the towns of Judah, each on his own property in the various towns,
NEH|11|4|while other people from both Judah and Benjamin lived in Jerusalem): From the descendants of Judah: Athaiah son of Uzziah, the son of Zechariah, the son of Amariah, the son of Shephatiah, the son of Mahalalel, a descendant of Perez;
NEH|11|5|and Maaseiah son of Baruch, the son of Col-Hozeh, the son of Hazaiah, the son of Adaiah, the son of Joiarib, the son of Zechariah, a descendant of Shelah.
NEH|11|6|The descendants of Perez who lived in Jerusalem totaled 468 able men.
NEH|11|7|From the descendants of Benjamin: Sallu son of Meshullam, the son of Joed, the son of Pedaiah, the son of Kolaiah, the son of Maaseiah, the son of Ithiel, the son of Jeshaiah,
NEH|11|8|and his followers, Gabbai and Sallai-928 men.
NEH|11|9|Joel son of Zicri was their chief officer, and Judah son of Hassenuah was over the Second District of the city.
NEH|11|10|From the priests: Jedaiah; the son of Joiarib; Jakin;
NEH|11|11|Seraiah son of Hilkiah, the son of Meshullam, the son of Zadok, the son of Meraioth, the son of Ahitub, supervisor in the house of God,
NEH|11|12|and their associates, who carried on work for the temple-822 men; Adaiah son of Jeroham, the son of Pelaliah, the son of Amzi, the son of Zechariah, the son of Pashhur, the son of Malkijah,
NEH|11|13|and his associates, who were heads of families-242 men; Amashsai son of Azarel, the son of Ahzai, the son of Meshillemoth, the son of Immer,
NEH|11|14|and his associates, who were able men-128. Their chief officer was Zabdiel son of Haggedolim.
NEH|11|15|From the Levites: Shemaiah son of Hasshub, the son of Azrikam, the son of Hashabiah, the son of Bunni;
NEH|11|16|Shabbethai and Jozabad, two of the heads of the Levites, who had charge of the outside work of the house of God;
NEH|11|17|Mattaniah son of Mica, the son of Zabdi, the son of Asaph, the director who led in thanksgiving and prayer; Bakbukiah, second among his associates; and Abda son of Shammua, the son of Galal, the son of Jeduthun.
NEH|11|18|The Levites in the holy city totaled 284.
NEH|11|19|The gatekeepers: Akkub, Talmon and their associates, who kept watch at the gates-172 men.
NEH|11|20|The rest of the Israelites, with the priests and Levites, were in all the towns of Judah, each on his ancestral property.
NEH|11|21|The temple servants lived on the hill of Ophel, and Ziha and Gishpa were in charge of them.
NEH|11|22|The chief officer of the Levites in Jerusalem was Uzzi son of Bani, the son of Hashabiah, the son of Mattaniah, the son of Mica. Uzzi was one of Asaph's descendants, who were the singers responsible for the service of the house of God.
NEH|11|23|The singers were under the king's orders, which regulated their daily activity.
NEH|11|24|Pethahiah son of Meshezabel, one of the descendants of Zerah son of Judah, was the king's agent in all affairs relating to the people.
NEH|11|25|As for the villages with their fields, some of the people of Judah lived in Kiriath Arba and its surrounding settlements, in Dibon and its settlements, in Jekabzeel and its villages,
NEH|11|26|in Jeshua, in Moladah, in Beth Pelet,
NEH|11|27|in Hazar Shual, in Beersheba and its settlements,
NEH|11|28|in Ziklag, in Meconah and its settlements,
NEH|11|29|in En Rimmon, in Zorah, in Jarmuth,
NEH|11|30|Zanoah, Adullam and their villages, in Lachish and its fields, and in Azekah and its settlements. So they were living all the way from Beersheba to the Valley of Hinnom.
NEH|11|31|The descendants of the Benjamites from Geba lived in Micmash, Aija, Bethel and its settlements,
NEH|11|32|in Anathoth, Nob and Ananiah,
NEH|11|33|in Hazor, Ramah and Gittaim,
NEH|11|34|in Hadid, Zeboim and Neballat,
NEH|11|35|in Lod and Ono, and in the Valley of the Craftsmen.
NEH|11|36|Some of the divisions of the Levites of Judah settled in Benjamin.
NEH|12|1|These were the priests and Levites who returned with Zerubbabel son of Shealtiel and with Jeshua: Seraiah, Jeremiah, Ezra,
NEH|12|2|Amariah, Malluch, Hattush,
NEH|12|3|Shecaniah, Rehum, Meremoth,
NEH|12|4|Iddo, Ginnethon, Abijah,
NEH|12|5|Mijamin, Moadiah, Bilgah,
NEH|12|6|Shemaiah, Joiarib, Jedaiah,
NEH|12|7|Sallu, Amok, Hilkiah and Jedaiah. These were the leaders of the priests and their associates in the days of Jeshua.
NEH|12|8|The Levites were Jeshua, Binnui, Kadmiel, Sherebiah, Judah, and also Mattaniah, who, together with his associates, was in charge of the songs of thanksgiving.
NEH|12|9|Bakbukiah and Unni, their associates, stood opposite them in the services.
NEH|12|10|Jeshua was the father of Joiakim, Joiakim the father of Eliashib, Eliashib the father of Joiada,
NEH|12|11|Joiada the father of Jonathan, and Jonathan the father of Jaddua.
NEH|12|12|In the days of Joiakim, these were the heads of the priestly families: of Seraiah's family, Meraiah; of Jeremiah's, Hananiah;
NEH|12|13|of Ezra's, Meshullam; of Amariah's, Jehohanan;
NEH|12|14|of Malluch's, Jonathan; of Shecaniah's, Joseph;
NEH|12|15|of Harim's, Adna; of Meremoth's, Helkai;
NEH|12|16|of Iddo's, Zechariah; of Ginnethon's, Meshullam;
NEH|12|17|of Abijah's, Zicri; of Miniamin's and of Moadiah's, Piltai;
NEH|12|18|of Bilgah's, Shammua; of Shemaiah's, Jehonathan;
NEH|12|19|of Joiarib's, Mattenai; of Jedaiah's, Uzzi;
NEH|12|20|of Sallu's, Kallai; of Amok's, Eber;
NEH|12|21|of Hilkiah's, Hashabiah; of Jedaiah's, Nethanel.
NEH|12|22|The family heads of the Levites in the days of Eliashib, Joiada, Johanan and Jaddua, as well as those of the priests, were recorded in the reign of Darius the Persian.
NEH|12|23|The family heads among the descendants of Levi up to the time of Johanan son of Eliashib were recorded in the book of the annals.
NEH|12|24|And the leaders of the Levites were Hashabiah, Sherebiah, Jeshua son of Kadmiel, and their associates, who stood opposite them to give praise and thanksgiving, one section responding to the other, as prescribed by David the man of God.
NEH|12|25|Mattaniah, Bakbukiah, Obadiah, Meshullam, Talmon and Akkub were gatekeepers who guarded the storerooms at the gates.
NEH|12|26|They served in the days of Joiakim son of Jeshua, the son of Jozadak, and in the days of Nehemiah the governor and of Ezra the priest and scribe.
NEH|12|27|At the dedication of the wall of Jerusalem, the Levites were sought out from where they lived and were brought to Jerusalem to celebrate joyfully the dedication with songs of thanksgiving and with the music of cymbals, harps and lyres.
NEH|12|28|The singers also were brought together from the region around Jerusalem-from the villages of the Netophathites,
NEH|12|29|from Beth Gilgal, and from the area of Geba and Azmaveth, for the singers had built villages for themselves around Jerusalem.
NEH|12|30|When the priests and Levites had purified themselves ceremonially, they purified the people, the gates and the wall.
NEH|12|31|I had the leaders of Judah go up on top of the wall. I also assigned two large choirs to give thanks. One was to proceed on top of the wall to the right, toward the Dung Gate.
NEH|12|32|Hoshaiah and half the leaders of Judah followed them,
NEH|12|33|along with Azariah, Ezra, Meshullam,
NEH|12|34|Judah, Benjamin, Shemaiah, Jeremiah,
NEH|12|35|as well as some priests with trumpets, and also Zechariah son of Jonathan, the son of Shemaiah, the son of Mattaniah, the son of Micaiah, the son of Zaccur, the son of Asaph,
NEH|12|36|and his associates-Shemaiah, Azarel, Milalai, Gilalai, Maai, Nethanel, Judah and Hanani-with musical instruments prescribed by David the man of God. Ezra the scribe led the procession.
NEH|12|37|At the Fountain Gate they continued directly up the steps of the City of David on the ascent to the wall and passed above the house of David to the Water Gate on the east.
NEH|12|38|The second choir proceeded in the opposite direction. I followed them on top of the wall, together with half the people-past the Tower of the Ovens to the Broad Wall,
NEH|12|39|over the Gate of Ephraim, the Jeshanah Gate, the Fish Gate, the Tower of Hananel and the Tower of the Hundred, as far as the Sheep Gate. At the Gate of the Guard they stopped.
NEH|12|40|The two choirs that gave thanks then took their places in the house of God; so did I, together with half the officials,
NEH|12|41|as well as the priests-Eliakim, Maaseiah, Miniamin, Micaiah, Elioenai, Zechariah and Hananiah with their trumpets-
NEH|12|42|and also Maaseiah, Shemaiah, Eleazar, Uzzi, Jehohanan, Malkijah, Elam and Ezer. The choirs sang under the direction of Jezrahiah.
NEH|12|43|And on that day they offered great sacrifices, rejoicing because God had given them great joy. The women and children also rejoiced. The sound of rejoicing in Jerusalem could be heard far away.
NEH|12|44|At that time men were appointed to be in charge of the storerooms for the contributions, firstfruits and tithes. From the fields around the towns they were to bring into the storerooms the portions required by the Law for the priests and the Levites, for Judah was pleased with the ministering priests and Levites.
NEH|12|45|They performed the service of their God and the service of purification, as did also the singers and gatekeepers, according to the commands of David and his son Solomon.
NEH|12|46|For long ago, in the days of David and Asaph, there had been directors for the singers and for the songs of praise and thanksgiving to God.
NEH|12|47|So in the days of Zerubbabel and of Nehemiah, all Israel contributed the daily portions for the singers and gatekeepers. They also set aside the portion for the other Levites, and the Levites set aside the portion for the descendants of Aaron.
NEH|13|1|On that day the Book of Moses was read aloud in the hearing of the people and there it was found written that no Ammonite or Moabite should ever be admitted into the assembly of God,
NEH|13|2|because they had not met the Israelites with food and water but had hired Balaam to call a curse down on them. (Our God, however, turned the curse into a blessing.)
NEH|13|3|When the people heard this law, they excluded from Israel all who were of foreign descent.
NEH|13|4|Before this, Eliashib the priest had been put in charge of the storerooms of the house of our God. He was closely associated with Tobiah,
NEH|13|5|and he had provided him with a large room formerly used to store the grain offerings and incense and temple articles, and also the tithes of grain, new wine and oil prescribed for the Levites, singers and gatekeepers, as well as the contributions for the priests.
NEH|13|6|But while all this was going on, I was not in Jerusalem, for in the thirty-second year of Artaxerxes king of Babylon I had returned to the king. Some time later I asked his permission
NEH|13|7|and came back to Jerusalem. Here I learned about the evil thing Eliashib had done in providing Tobiah a room in the courts of the house of God.
NEH|13|8|I was greatly displeased and threw all Tobiah's household goods out of the room.
NEH|13|9|I gave orders to purify the rooms, and then I put back into them the equipment of the house of God, with the grain offerings and the incense.
NEH|13|10|I also learned that the portions assigned to the Levites had not been given to them, and that all the Levites and singers responsible for the service had gone back to their own fields.
NEH|13|11|So I rebuked the officials and asked them, "Why is the house of God neglected?" Then I called them together and stationed them at their posts.
NEH|13|12|All Judah brought the tithes of grain, new wine and oil into the storerooms.
NEH|13|13|I put Shelemiah the priest, Zadok the scribe, and a Levite named Pedaiah in charge of the storerooms and made Hanan son of Zaccur, the son of Mattaniah, their assistant, because these men were considered trustworthy. They were made responsible for distributing the supplies to their brothers.
NEH|13|14|Remember me for this, O my God, and do not blot out what I have so faithfully done for the house of my God and its services.
NEH|13|15|In those days I saw men in Judah treading winepresses on the Sabbath and bringing in grain and loading it on donkeys, together with wine, grapes, figs and all other kinds of loads. And they were bringing all this into Jerusalem on the Sabbath. Therefore I warned them against selling food on that day.
NEH|13|16|Men from Tyre who lived in Jerusalem were bringing in fish and all kinds of merchandise and selling them in Jerusalem on the Sabbath to the people of Judah.
NEH|13|17|I rebuked the nobles of Judah and said to them, "What is this wicked thing you are doing-desecrating the Sabbath day?
NEH|13|18|Didn't your forefathers do the same things, so that our God brought all this calamity upon us and upon this city? Now you are stirring up more wrath against Israel by desecrating the Sabbath."
NEH|13|19|When evening shadows fell on the gates of Jerusalem before the Sabbath, I ordered the doors to be shut and not opened until the Sabbath was over. I stationed some of my own men at the gates so that no load could be brought in on the Sabbath day.
NEH|13|20|Once or twice the merchants and sellers of all kinds of goods spent the night outside Jerusalem.
NEH|13|21|But I warned them and said, "Why do you spend the night by the wall? If you do this again, I will lay hands on you." From that time on they no longer came on the Sabbath.
NEH|13|22|Then I commanded the Levites to purify themselves and go and guard the gates in order to keep the Sabbath day holy. Remember me for this also, O my God, and show mercy to me according to your great love.
NEH|13|23|Moreover, in those days I saw men of Judah who had married women from Ashdod, Ammon and Moab.
NEH|13|24|Half of their children spoke the language of Ashdod or the language of one of the other peoples, and did not know how to speak the language of Judah.
NEH|13|25|I rebuked them and called curses down on them. I beat some of the men and pulled out their hair. I made them take an oath in God's name and said: "You are not to give your daughters in marriage to their sons, nor are you to take their daughters in marriage for your sons or for yourselves.
NEH|13|26|Was it not because of marriages like these that Solomon king of Israel sinned? Among the many nations there was no king like him. He was loved by his God, and God made him king over all Israel, but even he was led into sin by foreign women.
NEH|13|27|Must we hear now that you too are doing all this terrible wickedness and are being unfaithful to our God by marrying foreign women?"
NEH|13|28|One of the sons of Joiada son of Eliashib the high priest was son-in-law to Sanballat the Horonite. And I drove him away from me.
NEH|13|29|Remember them, O my God, because they defiled the priestly office and the covenant of the priesthood and of the Levites.
NEH|13|30|So I purified the priests and the Levites of everything foreign, and assigned them duties, each to his own task.
NEH|13|31|I also made provision for contributions of wood at designated times, and for the firstfruits. Remember me with favor, O my God.
