EXOD|1|1|Вот имена сынов Израилевых, которые вошли в Египет с Иаковом, вошли каждый с домом своим:
EXOD|1|2|Рувим, Симеон, Левий и Иуда,
EXOD|1|3|Иссахар, Завулон и Вениамин,
EXOD|1|4|Дан и Неффалим, Гад и Асир.
EXOD|1|5|Всех же душ, происшедших от чресл Иакова, было семьдесят, а Иосиф был [уже] в Египте.
EXOD|1|6|И умер Иосиф и все братья его и весь род их;
EXOD|1|7|а сыны Израилевы расплодились и размножились, и возросли и усилились чрезвычайно, и наполнилась ими земля та.
EXOD|1|8|И восстал в Египте новый царь, который не знал Иосифа,
EXOD|1|9|и сказал народу своему: вот, народ сынов Израилевых многочислен и сильнее нас;
EXOD|1|10|перехитрим же его, чтобы он не размножался; иначе, когда случится война, соединится и он с нашими неприятелями, и вооружится против нас, и выйдет из земли [нашей].
EXOD|1|11|И поставили над ним начальников работ, чтобы изнуряли его тяжкими работами. И он построил фараону Пифом и Раамсес, города для запасов.
EXOD|1|12|Но чем более изнуряли его, тем более он умножался и тем более возрастал, так что опасались сынов Израилевых.
EXOD|1|13|И потому Египтяне с жестокостью принуждали сынов Израилевых к работам
EXOD|1|14|и делали жизнь их горькою от тяжкой работы над глиною и кирпичами и от всякой работы полевой, от всякой работы, к которой принуждали их с жестокостью.
EXOD|1|15|Царь Египетский повелел повивальным бабкам Евреянок, из коих одной имя Шифра, а другой Фуа,
EXOD|1|16|и сказал: когда вы будете повивать у Евреянок, то наблюдайте при родах: если будет сын, то умерщвляйте его, а если дочь, то пусть живет.
EXOD|1|17|Но повивальные бабки боялись Бога и не делали так, как говорил им царь Египетский, и оставляли детей в живых.
EXOD|1|18|Царь Египетский призвал повивальных бабок и сказал им: для чего вы делаете такое дело, что оставляете детей в живых?
EXOD|1|19|Повивальные бабки сказали фараону: Еврейские женщины не так, как Египетские; они здоровы, ибо прежде нежели придет к ним повивальная бабка, они уже рождают.
EXOD|1|20|За сие Бог делал добро повивальным бабкам, а народ умножался и весьма усиливался.
EXOD|1|21|И так как повивальные бабки боялись Бога, то Он устроял домы их.
EXOD|1|22|Тогда фараон всему народу своему повелел, говоря: всякого новорожденного [у Евреев] сына бросайте в реку, а всякую дочь оставляйте в живых.
EXOD|2|1|Некто из племени Левиина пошел и взял себе жену из того же племени.
EXOD|2|2|Жена зачала и родила сына и, видя, что он очень красив, скрывала его три месяца;
EXOD|2|3|но не могши долее скрывать его, взяла корзинку из тростника и осмолила ее асфальтом и смолою и, положив в нее младенца, поставила в тростнике у берега реки,
EXOD|2|4|а сестра его стала вдали наблюдать, что с ним будет.
EXOD|2|5|И вышла дочь фараонова на реку мыться, а прислужницы ее ходили по берегу реки. Она увидела корзинку среди тростника и послала рабыню свою взять ее.
EXOD|2|6|Открыла и увидела младенца; и вот, дитя плачет; и сжалилась над ним и сказала: это из Еврейских детей.
EXOD|2|7|И сказала сестра его дочери фараоновой: не сходить ли мне и не позвать ли к тебе кормилицу из Евреянок, чтоб она вскормила тебе младенца?
EXOD|2|8|Дочь фараонова сказала ей: сходи. Девица пошла и призвала мать младенца.
EXOD|2|9|Дочь фараонова сказала ей: возьми младенца сего и вскорми его мне; я дам тебе плату. Женщина взяла младенца и кормила его.
EXOD|2|10|И вырос младенец, и она привела его к дочери фараоновой, и он был у нее вместо сына, и нарекла имя ему: Моисей, потому что, говорила она, я из воды вынула его.
EXOD|2|11|Спустя много времени, когда Моисей вырос, случилось, что он вышел к братьям своим [сынам Израилевым] и увидел тяжкие работы их; и увидел, что Египтянин бьет одного Еврея из братьев его.
EXOD|2|12|Посмотрев туда и сюда и видя, что нет никого, он убил Египтянина и скрыл его в песке.
EXOD|2|13|И вышел он на другой день, и вот, два Еврея ссорятся; и сказал он обижающему: зачем ты бьешь ближнего твоего?
EXOD|2|14|А тот сказал: кто поставил тебя начальником и судьею над нами? не думаешь ли убить меня, как убил Египтянина? Моисей испугался и сказал: верно, узнали об этом деле.
EXOD|2|15|И услышал фараон об этом деле и хотел убить Моисея; но Моисей убежал от фараона и остановился в земле Мадиамской, и сел у колодезя.
EXOD|2|16|У священника Мадиамского [было] семь дочерей. Они пришли, начерпали [воды] и наполнили корыта, чтобы напоить овец отца своего.
EXOD|2|17|И пришли пастухи и отогнали их. Тогда встал Моисей и защитил их, и напоил овец их.
EXOD|2|18|И пришли они к Рагуилу, отцу своему, и он сказал: что вы так скоро пришли сегодня?
EXOD|2|19|Они сказали: какой–то Египтянин защитил нас от пастухов, и даже начерпал нам воды и напоил овец.
EXOD|2|20|Он сказал дочерям своим: где же он? зачем вы его оставили? позовите его, и пусть он ест хлеб.
EXOD|2|21|Моисею понравилось жить у сего человека; и он выдал за Моисея дочь свою Сепфору.
EXOD|2|22|Она родила сына, и [Моисей] нарек ему имя: Гирсам, потому что, говорил он, я стал пришельцем в чужой земле.
EXOD|2|23|Спустя долгое время, умер царь Египетский. И стенали сыны Израилевы от работы и вопияли, и вопль их от работы восшел к Богу.
EXOD|2|24|И услышал Бог стенание их, и вспомнил Бог завет Свой с Авраамом, Исааком и Иаковом.
EXOD|2|25|И увидел Бог сынов Израилевых, и призрел их Бог.
EXOD|3|1|Моисей пас овец у Иофора, тестя своего, священника Мадиамского. Однажды провел он стадо далеко в пустыню и пришел к горе Божией, Хориву.
EXOD|3|2|И явился ему Ангел Господень в пламени огня из среды тернового куста. И увидел он, что терновый куст горит огнем, но куст не сгорает.
EXOD|3|3|Моисей сказал: пойду и посмотрю на сие великое явление, отчего куст не сгорает.
EXOD|3|4|Господь увидел, что он идет смотреть, и воззвал к нему Бог из среды куста, и сказал: Моисей! Моисей! Он сказал: вот я!
EXOD|3|5|И сказал Бог: не подходи сюда; сними обувь твою с ног твоих, ибо место, на котором ты стоишь, есть земля святая.
EXOD|3|6|И сказал: Я Бог отца твоего, Бог Авраама, Бог Исаака и Бог Иакова. Моисей закрыл лице свое, потому что боялся воззреть на Бога.
EXOD|3|7|И сказал Господь: Я увидел страдание народа Моего в Египте и услышал вопль его от приставников его; Я знаю скорби его
EXOD|3|8|и иду избавить его от руки Египтян и вывести его из земли сей в землю хорошую и пространную, где течет молоко и мед, в землю Хананеев, Хеттеев, Аморреев, Ферезеев, Евеев и Иевусеев.
EXOD|3|9|И вот, уже вопль сынов Израилевых дошел до Меня, и Я вижу угнетение, каким угнетают их Египтяне.
EXOD|3|10|Итак пойди: Я пошлю тебя к фараону; и выведи из Египта народ Мой, сынов Израилевых.
EXOD|3|11|Моисей сказал Богу: кто я, чтобы мне идти к фараону и вывести из Египта сынов Израилевых?
EXOD|3|12|И сказал [Бог]: Я буду с тобою, и вот тебе знамение, что Я послал тебя: когда ты выведешь народ из Египта, вы совершите служение Богу на этой горе.
EXOD|3|13|И сказал Моисей Богу: вот, я приду к сынам Израилевым и скажу им: Бог отцов ваших послал меня к вам. А они скажут мне: как Ему имя? Что сказать мне им?
EXOD|3|14|Бог сказал Моисею: Я есмь Сущий. И сказал: так скажи сынам Израилевым: Сущий [Иегова] послал меня к вам.
EXOD|3|15|И сказал еще Бог Моисею: так скажи сынам Израилевым: Господь, Бог отцов ваших, Бог Авраама, Бог Исаака и Бог Иакова послал меня к вам. Вот имя Мое на веки, и памятование о Мне из рода в род.
EXOD|3|16|Пойди, собери старейшин Израилевых и скажи им: Господь, Бог отцов ваших, явился мне, Бог Авраама, Исаака и Иакова, и сказал: Я посетил вас и [увидел], что делается с вами в Египте.
EXOD|3|17|И сказал: Я выведу вас от угнетения Египетского в землю Хананеев, Хеттеев, Аморреев, Ферезеев, Евеев и Иевусеев, в землю, где течет молоко и мед.
EXOD|3|18|И они послушают голоса твоего, и пойдешь ты и старейшины Израилевы к царю Египетскому, и скажете ему: Господь, Бог Евреев, призвал нас; итак отпусти нас в пустыню, на три дня пути, чтобы принести жертву Господу, Богу нашему.
EXOD|3|19|Но Я знаю, что царь Египетский не позволит вам идти, если [не принудить его] рукою крепкою;
EXOD|3|20|и простру руку Мою и поражу Египет всеми чудесами Моими, которые сделаю среди его; и после того он отпустит вас.
EXOD|3|21|И дам народу сему милость в глазах Египтян; и когда пойдете, то пойдете не с пустыми руками:
EXOD|3|22|каждая женщина выпросит у соседки своей и у живущей в доме ее вещей серебряных и вещей золотых, и одежд, и вы нарядите ими и сыновей ваших и дочерей ваших, и оберете Египтян.
EXOD|4|1|И отвечал Моисей и сказал: а если они не поверят мне и не послушают голоса моего и скажут: не явился тебе Господь?
EXOD|4|2|И сказал ему Господь: что это в руке у тебя? Он отвечал: жезл.
EXOD|4|3|[Господь] сказал: брось его на землю. Он бросил его на землю, и жезл превратился в змея, и Моисей побежал от него.
EXOD|4|4|И сказал Господь Моисею: простри руку твою и возьми его за хвост. Он простер руку свою, и взял его; и он стал жезлом в руке его.
EXOD|4|5|Это для того, чтобы поверили, что явился тебе Господь, Бог отцов их, Бог Авраама, Бог Исаака и Бог Иакова.
EXOD|4|6|Еще сказал ему Господь: положи руку твою к себе в пазуху. И он положил руку свою к себе в пазуху, вынул ее, и вот, рука его побелела от проказы, как снег.
EXOD|4|7|[Еще] сказал: положи опять руку твою к себе в пазуху. И он положил руку свою к себе в пазуху; и вынул ее из пазухи своей, и вот, она опять стала такою же, как тело его.
EXOD|4|8|Если они не поверят тебе и не послушают голоса первого знамения, то поверят голосу знамения другого;
EXOD|4|9|если же не поверят и двум сим знамениям и не послушают голоса твоего, то возьми воды [из] реки и вылей на сушу; и вода, взятая из реки, сделается кровью на суше.
EXOD|4|10|И сказал Моисей Господу: о, Господи! человек я не речистый, [и] [таков был] и вчера и третьего дня, и когда Ты начал говорить с рабом Твоим: я тяжело говорю и косноязычен.
EXOD|4|11|Господь сказал: кто дал уста человеку? кто делает немым, или глухим, или зрячим, или слепым? не Я ли Господь?
EXOD|4|12|итак пойди, и Я буду при устах твоих и научу тебя, что тебе говорить.
EXOD|4|13|[Моисей] сказал: Господи! пошли другого, кого можешь послать.
EXOD|4|14|И возгорелся гнев Господень на Моисея, и Он сказал: разве нет у тебя Аарона брата, Левитянина? Я знаю, что он может говорить, и вот, он выйдет навстречу тебе, и, увидев тебя, возрадуется в сердце своем;
EXOD|4|15|ты будешь ему говорить и влагать слова в уста его, а Я буду при устах твоих и при устах его и буду учить вас, что вам делать;
EXOD|4|16|и будет говорить он вместо тебя к народу; итак он будет твоими устами, а ты будешь ему вместо Бога;
EXOD|4|17|и жезл сей возьми в руку твою: им ты будешь творить знамения.
EXOD|4|18|И пошел Моисей, и возвратился к Иофору, тестю своему, и сказал ему: пойду я, и возвращусь к братьям моим, которые в Египте, и посмотрю, живы ли еще они? И сказал Иофор Моисею: иди с миром.
EXOD|4|19|И сказал Господь Моисею в [земле] Мадиамской: пойди, возвратись в Египет, ибо умерли все, искавшие души твоей.
EXOD|4|20|И взял Моисей жену свою и сыновей своих, посадил их на осла и отправился в землю Египетскую. И жезл Божий Моисей взял в руку свою.
EXOD|4|21|И сказал Господь Моисею: когда пойдешь и возвратишься в Египет, смотри, все чудеса, которые Я поручил тебе, сделай пред лицем фараона, а Я ожесточу сердце его, и он не отпустит народа.
EXOD|4|22|И скажи фараону: так говорит Господь: Израиль [есть] сын Мой, первенец Мой;
EXOD|4|23|Я говорю тебе: отпусти сына Моего, чтобы он совершил Мне служение; а если не отпустишь его, то вот, Я убью сына твоего, первенца твоего.
EXOD|4|24|Дорогою на ночлеге случилось, что встретил его Господь и хотел умертвить его.
EXOD|4|25|Тогда Сепфора, взяв каменный нож, обрезала крайнюю плоть сына своего и, бросив к ногам его, сказала: ты жених крови у меня.
EXOD|4|26|И отошел от него [Господь]. Тогда сказала она: жених крови – по обрезанию.
EXOD|4|27|И Господь сказал Аарону: пойди навстречу Моисею в пустыню. И он пошел, и встретился с ним при горе Божией, и поцеловал его.
EXOD|4|28|И пересказал Моисей Аарону все слова Господа, Который его послал, и все знамения, которые Он заповедал.
EXOD|4|29|И пошел Моисей с Аароном, и собрали они всех старейшин сынов Израилевых,
EXOD|4|30|и пересказал Аарон все слова, которые говорил Господь Моисею; и сделал [Моисей] знамения пред глазами народа,
EXOD|4|31|и поверил народ; и услышали, что Господь посетил сынов Израилевых и увидел страдание их, и преклонились они и поклонились.
EXOD|5|1|После сего Моисей и Аарон пришли к фараону и сказали: так говорит Господь, Бог Израилев: отпусти народ Мой, чтоб он совершил Мне праздник в пустыне.
EXOD|5|2|Но фараон сказал: кто такой Господь, чтоб я послушался голоса Его [и] отпустил Израиля? я не знаю Господа и Израиля не отпущу.
EXOD|5|3|Они сказали: Бог Евреев призвал нас; отпусти нас в пустыню на три дня пути принести жертву Господу, Богу нашему, чтобы Он не поразил нас язвою, или мечом.
EXOD|5|4|И сказал им царь Египетский: для чего вы, Моисей и Аарон, отвлекаете народ от дел его? ступайте на свою работу.
EXOD|5|5|И сказал фараон: вот, народ в земле сей многочислен, и вы отвлекаете его от работ его.
EXOD|5|6|И в тот же день фараон дал повеление приставникам над народом и надзирателям, говоря:
EXOD|5|7|не давайте впредь народу соломы для делания кирпича, как вчера и третьего дня, пусть они сами ходят и собирают себе солому,
EXOD|5|8|а кирпичей наложите на них то же урочное число, какое они делали вчера и третьего дня, и не убавляйте; они праздны, потому и кричат: пойдем, принесем жертву Богу нашему;
EXOD|5|9|дать им больше работы, чтоб они работали и не занимались пустыми речами.
EXOD|5|10|И вышли приставники народа и надзиратели его и сказали народу: так говорит фараон: не даю вам соломы;
EXOD|5|11|сами пойдите, берите себе солому, где найдете, а от работы вашей ничего не убавляется.
EXOD|5|12|И рассеялся народ по всей земле Египетской собирать жниво вместо соломы.
EXOD|5|13|Приставники же понуждали, говоря: выполняйте работу свою каждый день, как и тогда, когда была [у вас] солома.
EXOD|5|14|А надзирателей из сынов Израилевых, которых поставили над ними приставники фараоновы, били, говоря: почему вы вчера и сегодня не изготовляете урочного числа кирпичей, как было до сих пор?
EXOD|5|15|И пришли надзиратели сынов Израилевых и возопили к фараону, говоря: для чего ты так поступаешь с рабами твоими?
EXOD|5|16|соломы не дают рабам твоим, а кирпичи, говорят нам, делайте. И вот, рабов твоих бьют; грех народу твоему.
EXOD|5|17|Но он сказал: праздны вы, праздны, поэтому и говорите: пойдем, принесем жертву Господу.
EXOD|5|18|Пойдите же, работайте; соломы не дадут вам, а положенное число кирпичей давайте.
EXOD|5|19|И увидели надзиратели сынов Израилевых беду свою в словах: не убавляйте числа кирпичей, какое [положено] на каждый день.
EXOD|5|20|И когда они вышли от фараона, то встретились с Моисеем и Аароном, которые стояли, ожидая их,
EXOD|5|21|и сказали им: да видит и судит вам Господь за то, что вы сделали нас ненавистными в глазах фараона и рабов его и дали им меч в руки, чтобы убить нас.
EXOD|5|22|И обратился Моисей к Господу и сказал: Господи! для чего Ты подвергнул такому бедствию народ сей, для чего послал меня?
EXOD|5|23|ибо с того времени, как я пришел к фараону и стал говорить именем Твоим, он начал хуже поступать с народом сим; избавить же, – Ты не избавил народа Твоего.
EXOD|6|1|И сказал Господь Моисею: теперь увидишь ты, что Я сделаю с фараоном; по действию руки крепкой он отпустит их; по действию руки крепкой даже выгонит их из земли своей.
EXOD|6|2|И говорил Бог Моисею и сказал ему: Я Господь.
EXOD|6|3|Являлся Я Аврааму, Исааку и Иакову с [именем] "Бог Всемогущий", а с именем [Моим] "Господь" не открылся им;
EXOD|6|4|и Я поставил завет Мой с ними, чтобы дать им землю Ханаанскую, землю странствования их, в которой они странствовали.
EXOD|6|5|И Я услышал стенание сынов Израилевых о том, что Египтяне держат их в рабстве, и вспомнил завет Мой.
EXOD|6|6|Итак скажи сынам Израилевым: Я Господь, и выведу вас из–под ига Египтян, и избавлю вас от рабства их, и спасу вас мышцею простертою и судами великими;
EXOD|6|7|и приму вас Себе в народ и буду вам Богом, и вы узнаете, что Я Господь, Бог ваш, изведший вас из–под ига Египетского;
EXOD|6|8|и введу вас в ту землю, о которой Я, подняв руку Мою, [клялся] дать ее Аврааму, Исааку и Иакову, и дам вам ее в наследие. Я Господь.
EXOD|6|9|Моисей пересказал это сынам Израилевым; но они не послушали Моисея по малодушию и тяжести работ.
EXOD|6|10|И сказал Господь Моисею, говоря:
EXOD|6|11|войди, скажи фараону, царю Египетскому, чтобы он отпустил сынов Израилевых из земли своей.
EXOD|6|12|И сказал Моисей пред Господом, говоря: вот, сыны Израилевы не слушают меня; как же послушает меня фараон? а я не словесен.
EXOD|6|13|И говорил Господь Моисею и Аарону, и давал им повеления к сынам Израилевым и к фараону, царю Египетскому, чтобы вывести сынов Израилевых из земли Египетской.
EXOD|6|14|Вот начальники поколений их: сыны Рувима, первенца Израилева: Ханох и Фаллу, Хецрон и Харми: это семейства Рувимовы.
EXOD|6|15|Сыны Симеона: Иемуил и Иамин, и Огад, и Иахин, и Цохар, и Саул, сын Хананеянки: это семейства Симеона.
EXOD|6|16|Вот имена сынов Левия по родам их: Гирсон и Кааф и Мерари. А лет жизни Левия было сто тридцать семь.
EXOD|6|17|Сыны Гирсона: Ливни и Шимеи с семействами их.
EXOD|6|18|Сыны Каафовы: Амрам и Ицгар, и Хеврон, и Узиил. А лет жизни Каафа было сто тридцать три года.
EXOD|6|19|Сыны Мерари: Махли и Муши. Это семейства Левия по родам их.
EXOD|6|20|Амрам взял Иохаведу, тетку свою, себе в жену, и она родила ему Аарона и Моисея. А лет жизни Амрама было сто тридцать семь.
EXOD|6|21|Сыны Ицгаровы: Корей и Нефег и Зихри.
EXOD|6|22|Сыны Узииловы: Мисаил и Елцафан и Сифри.
EXOD|6|23|Аарон взял себе в жену Елисавету, дочь Аминадава, сестру Наассона, и она родила ему Надава и Авиуда, Елеазара и Ифамара.
EXOD|6|24|Сыны Корея: Асир, Елкана и Авиасаф: это семейства Кореевы.
EXOD|6|25|Елеазар, сын Аарона, взял себе в жену [одну] из дочерей Футииловых, и она родила ему Финееса. Вот начальники поколений левитских по семействам их.
EXOD|6|26|Аарон и Моисей, это – те, которым сказал Господь: выведите сынов Израилевых из земли Египетской по ополчениям их.
EXOD|6|27|Они–то говорили фараону, царю Египетскому, чтобы вывести сынов Израилевых из Египта; это – Моисей и Аарон.
EXOD|6|28|Итак в то время, когда Господь говорил Моисею в земле Египетской,
EXOD|6|29|Господь сказал Моисею, говоря: Я Господь! скажи фараону, царю Египетскому, все, что Я говорю тебе.
EXOD|6|30|Моисей же сказал пред Господом: вот, я несловесен: как же послушает меня фараон?
EXOD|7|1|Но Господь сказал Моисею: смотри, Я поставил тебя Богом фараону, а Аарон, брат твой, будет твоим пророком:
EXOD|7|2|ты будешь говорить все, что Я повелю тебе, а Аарон, брат твой, будет говорить фараону, чтобы он отпустил сынов Израилевых из земли своей;
EXOD|7|3|но Я ожесточу сердце фараоново, и явлю множество знамений Моих и чудес Моих в земле Египетской;
EXOD|7|4|фараон не послушает вас, и Я наложу руку Мою на Египет и выведу воинство Мое, народ Мой, сынов Израилевых, из земли Египетской – судами великими;
EXOD|7|5|тогда узнают Египтяне, что Я Господь, когда простру руку Мою на Египет и выведу сынов Израилевых из среды их.
EXOD|7|6|И сделали Моисей и Аарон, как повелел им Господь, так они и сделали.
EXOD|7|7|Моисей [был] восьмидесяти, а Аарон восьмидесяти трех лет, когда стали говорить они к фараону.
EXOD|7|8|И сказал Господь Моисею и Аарону, говоря:
EXOD|7|9|если фараон скажет вам: сделайте чудо, то ты скажи Аарону: возьми жезл твой и брось пред фараоном – он сделается змеем.
EXOD|7|10|Моисей и Аарон пришли к фараону, и сделали так, как повелел Господь. И бросил Аарон жезл свой пред фараоном и пред рабами его, и он сделался змеем.
EXOD|7|11|И призвал фараон мудрецов и чародеев; и эти волхвы Египетские сделали то же своими чарами:
EXOD|7|12|каждый из них бросил свой жезл, и они сделались змеями, но жезл Ааронов поглотил их жезлы.
EXOD|7|13|Сердце фараоново ожесточилось, и он не послушал их, как и говорил Господь.
EXOD|7|14|И сказал Господь Моисею: упорно сердце фараоново: он не хочет отпустить народ.
EXOD|7|15|Пойди к фараону завтра: вот, он выйдет к воде, ты стань на пути его, на берегу реки, и жезл, который превращался в змея, возьми в руку твою
EXOD|7|16|и скажи ему: Господь, Бог Евреев, послал меня сказать тебе: отпусти народ Мой, чтобы он совершил Мне служение в пустыне; но вот, ты доселе не послушался.
EXOD|7|17|Так говорит Господь: из сего узнаешь, что Я Господь: вот этим жезлом, который в руке моей, я ударю по воде, которая в реке, и она превратится в кровь,
EXOD|7|18|и рыба в реке умрет, и река воссмердит, и Египтянам омерзительно будет пить воду из реки.
EXOD|7|19|И сказал Господь Моисею: скажи Аарону: возьми жезл твой, и простри руку твою на воды Египтян: на реки их, на потоки их, на озера их и на всякое вместилище вод их, – и превратятся в кровь, и будет кровь по всей земле Египетской и в деревянных и в каменных сосудах.
EXOD|7|20|И сделали Моисей и Аарон, как повелел Господь. И поднял [Аарон] жезл и ударил по воде речной пред глазами фараона и пред глазами рабов его, и вся вода в реке превратилась в кровь,
EXOD|7|21|и рыба в реке вымерла, и река воссмердела, и Египтяне не могли пить воды из реки; и была кровь по всей земле Египетской.
EXOD|7|22|И волхвы Египетские чарами своими сделали то же. И ожесточилось сердце фараона, и не послушал их, как и говорил Господь.
EXOD|7|23|И оборотился фараон, и пошел в дом свой; и сердце его не тронулось и сим.
EXOD|7|24|И стали копать все Египтяне около реки [чтобы найти] воду для питья, потому что не могли пить воды из реки.
EXOD|7|25|И исполнилось семь дней после того, как Господь поразил реку.
EXOD|7|26|И сказал Господь Моисею: пойди к фараону и скажи ему: так говорит Господь: отпусти народ Мой, чтобы он совершил Мне служение;
EXOD|7|27|если же ты не согласишься отпустить, то вот, Я поражаю всю область твою жабами;
EXOD|7|28|и воскишит река жабами, и они выйдут и войдут в дом твой, и в спальню твою, и на постель твою, и в домы рабов твоих и народа твоего, и в печи твои, и в квашни твои,
EXOD|7|29|и на тебя, и на народ твой, и на всех рабов твоих взойдут жабы.
EXOD|8|1|И сказал Господь Моисею: скажи Аарону: простри руку твою с жезлом твоим на реки, на потоки и на озера и выведи жаб на землю Египетскую.
EXOD|8|2|Аарон простер руку свою на воды Египетские; и вышли жабы и покрыли землю Египетскую.
EXOD|8|3|То же сделали и волхвы чарами своими и вывели жаб на землю Египетскую.
EXOD|8|4|И призвал фараон Моисея и Аарона и сказал: помолитесь Господу, чтоб Он удалил жаб от меня и от народа моего, и я отпущу народ [Израильский] принести жертву Господу.
EXOD|8|5|Моисей сказал фараону: назначь мне сам, когда помолиться за тебя, за рабов твоих и за народ твой, чтобы жабы исчезли у тебя, в домах твоих, и остались только в реке.
EXOD|8|6|Он сказал: завтра. [Моисей] отвечал: [будет] по слову твоему, дабы ты узнал, что нет никого, как Господь Бог наш;
EXOD|8|7|и удалятся жабы от тебя, от домов твоих, и от рабов твоих и от твоего народа; только в реке они останутся.
EXOD|8|8|Моисей и Аарон вышли от фараона, и Моисей воззвал к Господу о жабах, которых Он навел на фараона.
EXOD|8|9|И сделал Господь по слову Моисея: жабы вымерли в домах, на дворах и на полях;
EXOD|8|10|и собрали их в груды, и воссмердела земля.
EXOD|8|11|И увидел фараон, что сделалось облегчение, и ожесточил сердце свое, и не послушал их, как и говорил Господь.
EXOD|8|12|И сказал Господь Моисею: скажи Аарону: простри жезл твой и ударь в персть земную, и сделается [персмь] мошками по всей земле Египетской.
EXOD|8|13|Так они и сделали: Аарон простер руку свою с жезлом своим и ударил в персть земную, и явились мошки на людях и на скоте. Вся персть земная сделалась мошками по всей земле Египетской.
EXOD|8|14|Старались также и волхвы чарами своими произвести мошек, но не могли. И были мошки на людях и на скоте.
EXOD|8|15|И сказали волхвы фараону: это перст Божий. Но сердце фараоново ожесточилось, и он не послушал их, как и говорил Господь.
EXOD|8|16|И сказал Господь Моисею: завтра встань рано и явись пред лице фараона. Вот, он пойдет к воде, и ты скажи ему: так говорит Господь: отпусти народ Мой, чтобы он совершил Мне служение.
EXOD|8|17|а если не отпустишь народа Моего, то вот, Я пошлю на тебя и на рабов твоих, и на народ твой, и в домы твои песьих мух, и наполнятся домы Египтян песьими мухами и самая земля, на которой они [живут];
EXOD|8|18|и отделю в тот день землю Гесем, на которой пребывает народ Мой, и там не будет песьих мух, дабы ты знал, что Я Господь среди земли;
EXOD|8|19|Я сделаю разделение между народом Моим и между народом твоим. Завтра будет сие знамение.
EXOD|8|20|Так и сделал Господь: налетело множество песьих мух в дом фараонов, и в домы рабов его, и на всю землю Египетскую: погибала земля от песьих мух.
EXOD|8|21|И призвал фараон Моисея и Аарона и сказал: пойдите, принесите жертву Богу вашему в сей земле.
EXOD|8|22|Но Моисей сказал: нельзя сего сделать, ибо отвратительно для Египтян жертвоприношение наше Господу, Богу нашему: если мы отвратительную для Египтян жертву станем приносить в глазах их, то не побьют ли они нас камнями?
EXOD|8|23|мы пойдем в пустыню, на три дня пути, и принесем жертву Господу, Богу нашему, как скажет нам.
EXOD|8|24|И сказал фараон: я отпущу вас принести жертву Господу Богу вашему в пустыне, только не уходите далеко; помолитесь обо мне.
EXOD|8|25|Моисей сказал: вот, я выхожу от тебя и помолюсь Господу, и удалятся песьи мухи от фараона, и от рабов его, и от народа его завтра, только фараон пусть перестанет обманывать, не отпуская народа принести жертву Господу.
EXOD|8|26|И вышел Моисей от фараона и помолился Господу.
EXOD|8|27|И сделал Господь по слову Моисея и удалил песьих мух от фараона, от рабов его и от народа его: не осталось ни одной.
EXOD|8|28|Но фараон ожесточил сердце свое и на этот раз и не отпустил народа.
EXOD|9|1|И сказал Господь Моисею: пойди к фараону и скажи ему: так говорит Господь, Бог Евреев: отпусти народ Мой, чтобы он совершил Мне служение;
EXOD|9|2|ибо если ты не захочешь отпустить и еще будешь удерживать его,
EXOD|9|3|то вот, рука Господня будет на скоте твоем, который в поле, на конях, на ослах, на верблюдах, на волах и овцах: будет моровая язва весьма тяжкая;
EXOD|9|4|и разделит Господь между скотом Израильским и скотом Египетским, и из всего [скота] сынов Израилевых не умрет ничего.
EXOD|9|5|И назначил Господь время, сказав: завтра сделает это Господь в земле сей.
EXOD|9|6|И сделал это Господь на другой день, и вымер весь скот Египетский; из скота же сынов Израилевых не умерло ничего.
EXOD|9|7|Фараон послал [узнать], и вот, из скота Израилевых не умерло ничего. Но сердце фараоново ожесточилось, и он не отпустил народа.
EXOD|9|8|И сказал Господь Моисею и Аарону: возьмите по полной горсти пепла из печи, и пусть бросит его Моисей к небу в глазах фараона;
EXOD|9|9|и поднимется пыль по всей земле Египетской, и будет на людях и на скоте воспаление с нарывами, во всей земле Египетской.
EXOD|9|10|Они взяли пепла из печи и предстали пред лице фараона. Моисей бросил его к небу, и сделалось воспаление с нарывами на людях и на скоте.
EXOD|9|11|И не могли волхвы устоять пред Моисеем по причине воспаления, потому что воспаление было на волхвах и на всех Египтянах.
EXOD|9|12|Но Господь ожесточил сердце фараона, и он не послушал их, как и говорил Господь Моисею.
EXOD|9|13|И сказал Господь Моисею: завтра встань рано и явись пред лице фараона, и скажи ему: так говорит Господь, Бог Евреев: отпусти народ Мой, чтобы он совершил Мне служение;
EXOD|9|14|ибо в этот раз Я пошлю все язвы Мои в сердце твое, и на рабов твоих, и на народ твой, дабы ты узнал, что нет подобного Мне на всей земле;
EXOD|9|15|так как Я простер руку Мою, то поразил бы тебя и народ твой язвою, и ты истреблен был бы с земли:
EXOD|9|16|но для того Я сохранил тебя, чтобы показать на тебе силу Мою, и чтобы возвещено было имя Мое по всей земле;
EXOD|9|17|ты еще противостоишь народу Моему, чтобы не отпускать его, –
EXOD|9|18|вот, Я пошлю завтра, в это самое время, град весьма сильный, которому подобного не было в Египте со дня основания его доныне;
EXOD|9|19|итак пошли собрать стада твои и все, что есть у тебя в поле: на всех людей и скот, которые останутся в поле и не соберутся в домы, падет град, и они умрут.
EXOD|9|20|Те из рабов фараоновых, которые убоялись слова Господня, поспешно собрали рабов своих и стада свои в домы;
EXOD|9|21|а кто не обратил сердца своего к слову Господню, тот оставил рабов своих и стада свои в поле.
EXOD|9|22|И сказал Господь Моисею: простри руку твою к небу, и падет град на всю землю Египетскую, на людей, на скот и на всю траву полевую в земле Египетской.
EXOD|9|23|И простер Моисей жезл свой к небу, и Господь произвел гром и град, и огонь разливался по земле; и послал Господь град на землю Египетскую;
EXOD|9|24|и был град и огонь между градом, [град] весьма сильный, какого не было во всей земле Египетской со времени населения ее.
EXOD|9|25|И побил град по всей земле Египетской все, что было в поле, от человека до скота, и всю траву полевую побил град, и все деревья в поле поломал;
EXOD|9|26|только в земле Гесем, где жили сыны Израилевы, не было града.
EXOD|9|27|И послал фараон, и призвал Моисея и Аарона, и сказал им: на этот раз я согрешил; Господь праведен, а я и народ мой виновны;
EXOD|9|28|помолитесь Господу: пусть перестанут громы Божии и град; и отпущу вас и не буду более удерживать.
EXOD|9|29|Моисей сказал ему: как скоро я выйду из города, простру руки мои к Господу; громы перестанут, и града более не будет, дабы ты узнал, что Господня земля;
EXOD|9|30|но я знаю, что ты и рабы твои еще не убоитесь Господа Бога.
EXOD|9|31|Лен и ячмень были побиты, потому что ячмень выколосился, а лен осеменился;
EXOD|9|32|а пшеница и полба не побиты, потому что они были поздние.
EXOD|9|33|И вышел Моисей от фараона из города и простер руки свои к Господу, и прекратились гром и град, и дождь перестал литься на землю.
EXOD|9|34|И увидел фараон, что перестал дождь и град и гром, и продолжал грешить, и отягчил сердце свое сам и рабы его.
EXOD|9|35|И ожесточилось сердце фараона, и он не отпустил сынов Израилевых, как и говорил Господь чрез Моисея.
EXOD|10|1|И сказал Господь Моисею: войди к фараону, ибо Я отягчил сердце его и сердце рабов его, чтобы явить между ними сии знамения Мои,
EXOD|10|2|и чтобы ты рассказывал сыну твоему и сыну сына твоего о том, что Я сделал в Египте, и о знамениях Моих, которые Я показал в нем, и чтобы вы знали, что Я Господь.
EXOD|10|3|Моисей и Аарон пришли к фараону и сказали ему: так говорит Господь, Бог Евреев: долго ли ты не смиришься предо Мною? отпусти народ Мой, чтобы он совершил Мне служение;
EXOD|10|4|а если ты не отпустишь народа Моего, то вот, завтра Я наведу саранчу на твою область:
EXOD|10|5|она покроет лице земли так, что нельзя будет видеть земли, и поест у вас оставшееся, уцелевшее от града; объест также все дерева, растущие у вас в поле,
EXOD|10|6|и наполнит домы твои, домы всех рабов твоих и домы всех Египтян, чего не видели отцы твои, ни отцы отцов твоих со дня, как живут на земле, даже до сего дня. [Моисей] обратился и вышел от фараона.
EXOD|10|7|Тогда рабы фараоновы сказали ему: долго ли он будет мучить нас? отпусти сих людей, пусть они совершат служение Господу, Богу своему; неужели ты еще не видишь, что Египет гибнет?
EXOD|10|8|И возвратили Моисея и Аарона к фараону, и [фараон] сказал им: пойдите, совершите служение Господу, Богу вашему; кто же и кто пойдет?
EXOD|10|9|И сказал Моисей: пойдем с малолетними нашими и стариками нашими, с сыновьями нашими и дочерями нашими, и с овцами нашими и с волами нашими пойдем, ибо у нас праздник Господу.
EXOD|10|10|[Фараон] сказал им: пусть будет так, Господь с вами! я готов отпустить вас: но зачем с детьми? видите, у вас худое намерение!
EXOD|10|11|нет: пойдите [одни] мужчины и совершите служение Господу, так как вы сего просили. И выгнали их от фараона.
EXOD|10|12|Тогда Господь сказал Моисею: простри руку твою на землю Египетскую, и пусть нападет саранча на землю Египетскую и поест всю траву земную [и] все, что уцелело от града.
EXOD|10|13|И простер Моисей жезл свой на землю Египетскую, и Господь навел на сию землю восточный ветер, [продолжавшийся] весь тот день и всю ночь. Настало утро, и восточный ветер нанес саранчу.
EXOD|10|14|И напала саранча на всю землю Египетскую и легла по всей стране Египетской в великом множестве: прежде не бывало такой саранчи, и после сего не будет такой;
EXOD|10|15|она покрыла лице всей земли, так что земли не было видно, и поела всю траву земную и все плоды древесные, уцелевшие от града, и не осталось никакой зелени ни на деревах, ни на траве полевой во всей земле Египетской.
EXOD|10|16|Фараон поспешно призвал Моисея и Аарона и сказал: согрешил я пред Господом, Богом вашим, и пред вами;
EXOD|10|17|теперь простите грех мой еще раз и помолитесь Господу Богу вашему, чтобы Он только отвратил от меня сию смерть.
EXOD|10|18|[Моисей] вышел от фараона и помолился Господу.
EXOD|10|19|И воздвигнул Господь с противной стороны западный весьма сильный ветер, и он понес саранчу и бросил ее в Чермное море: не осталось ни одной саранчи во всей стране Египетской.
EXOD|10|20|Но Господь ожесточил сердце фараона, и он не отпустил сынов Израилевых.
EXOD|10|21|И сказал Господь Моисею: простри руку твою к небу, и будет тьма на земле Египетской, осязаемая тьма.
EXOD|10|22|Моисей простер руку свою к небу, и была густая тьма по всей земле Египетской три дня;
EXOD|10|23|не видели друг друга, и никто не вставал с места своего три дня; у всех же сынов Израилевых был свет в жилищах их.
EXOD|10|24|Фараон призвал Моисея и сказал: пойдите, совершите служение Господу, пусть только останется мелкий и крупный скот ваш, а дети ваши пусть идут с вами.
EXOD|10|25|Но Моисей сказал: дай также в руки наши жертвы и всесожжения, чтобы принести Господу Богу нашему;
EXOD|10|26|пусть пойдут и стада наши с нами, не останется ни копыта; ибо из них мы возьмем на жертву Господу, Богу нашему; но доколе не придем туда, мы не знаем, что принести в жертву Господу.
EXOD|10|27|И ожесточил Господь сердце фараона, и он не захотел отпустить их.
EXOD|10|28|И сказал ему фараон: пойди от меня; берегись, не являйся более пред лице мое; в тот день, когда ты увидишь лице мое, умрешь.
EXOD|10|29|И сказал Моисей: как сказал ты, так и будет; я не увижу более лица твоего.
EXOD|11|1|И сказал Господь Моисею: еще одну казнь Я наведу на фараона и на Египтян; после того он отпустит вас отсюда; когда же он будет отпускать, с поспешностью будет гнать вас отсюда;
EXOD|11|2|внуши народу, чтобы каждый у ближнего своего и каждая женщина у ближней своей выпросили вещей серебряных и вещей золотых.
EXOD|11|3|И дал Господь милость народу [Своему] в глазах Египтян, да и Моисей был весьма велик в земле Египетской, в глазах рабов фараоновых и в глазах народа.
EXOD|11|4|И сказал Моисей: так говорит Господь: в полночь Я пройду посреди Египта,
EXOD|11|5|и умрет всякий первенец в земле Египетской от первенца фараона, который сидит на престоле своем, до первенца рабыни, которая при жерновах, и все первородное из скота;
EXOD|11|6|и будет вопль великий по всей земле Египетской, какого не бывало и какого не будет более;
EXOD|11|7|у всех же сынов Израилевых ни на человека, ни на скот не пошевелит пес языком своим, дабы вы знали, какое различие делает Господь между Египтянами и между Израильтянами.
EXOD|11|8|И придут все рабы твои сии ко мне и поклонятся мне, говоря: выйди ты и весь народ, которым ты предводительствуешь. После сего я и выйду. И вышел [Моисей] от фараона с гневом.
EXOD|11|9|И сказал Господь Моисею: не послушал вас фараон, чтобы умножились чудеса Мои в земле Египетской.
EXOD|11|10|Моисей и Аарон сделали все сии чудеса пред фараоном; но Господь ожесточил сердце фараона, и он не отпустил сынов Израилевых из земли своей.
EXOD|12|1|И сказал Господь Моисею и Аарону в земле Египетской, говоря:
EXOD|12|2|месяц сей [да будет] у вас началом месяцев, первым [да] [будет] он у вас между месяцами года.
EXOD|12|3|Скажите всему обществу Израилевых: в десятый [день] сего месяца пусть возьмут себе каждый одного агнца по семействам, по агнцу на семейство;
EXOD|12|4|а если семейство так мало, что не [съест] агнца, то пусть возьмет с соседом своим, ближайшим к дому своему, по числу душ: по той мере, сколько каждый съест, расчислитесь на агнца.
EXOD|12|5|Агнец у вас должен быть без порока, мужеского пола, однолетний; возьмите его от овец, или от коз,
EXOD|12|6|и пусть он хранится у вас до четырнадцатого дня сего месяца: тогда пусть заколет его все собрание общества Израильского вечером,
EXOD|12|7|и пусть возьмут от крови [его] и помажут на обоих косяках и на перекладине дверей в домах, где будут есть его;
EXOD|12|8|пусть съедят мясо его в сию самую ночь, испеченное на огне; с пресным хлебом и с горькими [травами] пусть съедят его;
EXOD|12|9|не ешьте от него недопеченного, или сваренного в воде, но ешьте испеченное на огне, голову с ногами и внутренностями;
EXOD|12|10|не оставляйте от него до утра; но оставшееся от него до утра сожгите на огне.
EXOD|12|11|Ешьте же его так: пусть будут чресла ваши препоясаны, обувь ваша на ногах ваших и посохи ваши в руках ваших, и ешьте его с поспешностью: это – Пасха Господня.
EXOD|12|12|А Я в сию самую ночь пройду по земле Египетской и поражу всякого первенца в земле Египетской, от человека до скота, и над всеми богами Египетскими произведу суд. Я Господь.
EXOD|12|13|И будет у вас кровь знамением на домах, где вы находитесь, и увижу кровь и пройду мимо вас, и не будет между вами язвы губительной, когда буду поражать землю Египетскую.
EXOD|12|14|И да будет вам день сей памятен, и празднуйте в оный праздник Господу во [все] роды ваши; [как] установление вечное празднуйте его.
EXOD|12|15|Семь дней ешьте пресный хлеб; с самого первого дня уничтожьте квасное в домах ваших, ибо кто будет есть квасное с первого дня до седьмого дня, душа та истреблена будет из среды Израиля.
EXOD|12|16|И в первый день да будет у вас священное собрание, и в седьмой день священное собрание: никакой работы не должно делать в них; только что есть каждому, одно то можно делать вам.
EXOD|12|17|Наблюдайте опресноки, ибо в сей самый день Я вывел ополчения ваши из земли Египетской, и наблюдайте день сей в роды ваши, как установление вечное.
EXOD|12|18|С четырнадцатого дня первого месяца, с вечера ешьте пресный хлеб до вечера двадцать первого дня того же месяца;
EXOD|12|19|семь дней не должно быть закваски в домах ваших, ибо кто будет есть квасное, душа та истреблена будет из общества Израилевых – пришлец ли то, или природный житель земли той.
EXOD|12|20|Ничего квасного не ешьте; во всяком местопребывании вашем ешьте пресный хлеб.
EXOD|12|21|И созвал Моисей всех старейшин Израилевых и сказал им: выберите и возьмите себе агнцев по семействам вашим и заколите пасху;
EXOD|12|22|и возьмите пучок иссопа, и обмочите в кровь, которая в сосуде, и помажьте перекладину и оба косяка дверей кровью, которая в сосуде; а вы никто не выходите за двери дома своего до утра.
EXOD|12|23|И пойдет Господь поражать Египет, и увидит кровь на перекладине и на обоих косяках, и пройдет Господь мимо дверей, и не попустит губителю войти в домы ваши для поражения.
EXOD|12|24|Храните сие, как закон для себя и для сынов своих на веки.
EXOD|12|25|Когда войдете в землю, которую Господь даст вам, как Он говорил, соблюдайте сие служение.
EXOD|12|26|И когда скажут вам дети ваши: что это за служение?
EXOD|12|27|скажите: это пасхальная жертва Господу, Который прошел мимо домов сынов Израилевых в Египте, когда поражал Египтян, и домы наши избавил. И преклонился народ и поклонился.
EXOD|12|28|И пошли сыны Израилевы и сделали: как повелел Господь Моисею и Аарону, так и сделали.
EXOD|12|29|В полночь Господь поразил всех первенцев в земле Египетской, от первенца фараона, сидевшего на престоле своем, до первенца узника, находившегося в темнице, и все первородное из скота.
EXOD|12|30|И встал фараон ночью сам и все рабы его и весь Египет; и сделался великий вопль в [земле] Египетской, ибо не было дома, где не было бы мертвеца.
EXOD|12|31|И призвал [фараон] Моисея и Аарона ночью и сказал: встаньте, выйдите из среды народа моего, как вы, так и сыны Израилевы, и пойдите, совершите служение Господу, как говорили вы;
EXOD|12|32|и мелкий и крупный скот ваш возьмите, как вы говорили; и пойдите и благословите меня.
EXOD|12|33|И понуждали Египтяне народ, чтобы скорее выслать его из земли той; ибо говорили они: мы все помрем.
EXOD|12|34|И понес народ тесто свое, прежде нежели оно вскисло; квашни их, завязанные в одеждах их, были на плечах их.
EXOD|12|35|И сделали сыны Израилевы по слову Моисея и просили у Египтян вещей серебряных и вещей золотых и одежд.
EXOD|12|36|Господь же дал милость народу [Своему] в глазах Египтян: и они давали ему, и обобрал он Египтян.
EXOD|12|37|И отправились сыны Израилевы из Раамсеса в Сокхоф до шестисот тысяч пеших мужчин, кроме детей;
EXOD|12|38|и множество разноплеменных людей вышли с ними, и мелкий и крупный скот, стадо весьма большое.
EXOD|12|39|И испекли они из теста, которое вынесли из Египта, пресные лепешки, ибо оно еще не вскисло, потому что они выгнаны были из Египта и не могли медлить, и даже пищи не приготовили себе на дорогу.
EXOD|12|40|Времени же, в которое сыны Израилевы обитали в Египте, было четыреста тридцать лет.
EXOD|12|41|По прошествии четырехсот тридцати лет, в этот самый день вышло все ополчение Господне из земли Египетской ночью.
EXOD|12|42|Это – ночь бдения Господу за изведение их из земли Египетской; эта самая ночь – бдение Господу у всех сынов Израилевых в роды их.
EXOD|12|43|И сказал Господь Моисею и Аарону: вот устав Пасхи: никакой иноплеменник не должен есть ее;
EXOD|12|44|а всякий раб, купленный за серебро, когда обрежешь его, может есть ее;
EXOD|12|45|поселенец и наемник не должен есть ее.
EXOD|12|46|В одном доме должно есть ее, не выносите мяса вон из дома и костей ее не сокрушайте.
EXOD|12|47|Все общество Израиля должно совершать ее.
EXOD|12|48|Если же поселится у тебя пришлец и захочет совершить Пасху Господу, то обрежь у него всех мужеского пола, и тогда пусть он приступит к совершению ее и будет как природный житель земли; а никакой необрезанный не должен есть ее;
EXOD|12|49|один закон да будет и для природного жителя и для пришельца, поселившегося между вами.
EXOD|12|50|И сделали все сыны Израилевы: как повелел Господь Моисею и Аарону, так и сделали.
EXOD|12|51|В этот самый день Господь вывел сынов Израилевых из земли Египетской по ополчениям их.
EXOD|13|1|И сказал Господь Моисею, говоря:
EXOD|13|2|освяти Мне каждого первенца, разверзающего всякие ложесна между сынами Израилевыми, от человека до скота: Мои они.
EXOD|13|3|И сказал Моисей народу: помните сей день, в который вышли вы из Египта, из дома рабства, ибо рукою крепкою вывел вас Господь оттоле, и не ешьте квасного:
EXOD|13|4|сегодня выходите вы, в месяце Авиве.
EXOD|13|5|И когда введет тебя Господь в землю Хананеев и Хеттеев, и Аморреев, и Евеев, и Иевусеев, о которой клялся Он отцам твоим, что даст тебе землю, где течет молоко и мед, то совершай сие служение в сем месяце;
EXOD|13|6|семь дней ешь пресный хлеб, и в седьмой день – праздник Господу;
EXOD|13|7|пресный хлеб должно есть семь дней, и не должно находиться у тебя квасного хлеба, и не должно находиться у тебя квасного во всех пределах твоих.
EXOD|13|8|И объяви в день тот сыну твоему, говоря: это ради того, что Господь сделал со мною, когда я вышел из Египта.
EXOD|13|9|И да будет тебе это знаком на руке твоей и памятником пред глазами твоими, дабы закон Господень был в устах твоих, ибо рукою крепкою вывел тебя Господь из Египта.
EXOD|13|10|Исполняй же устав сей в назначенное время, из года в год.
EXOD|13|11|И когда введет тебя Господь в землю Ханаанскую, как Он клялся тебе и отцам твоим, и даст ее тебе, –
EXOD|13|12|отделяй Господу все, разверзающее ложесна; и все первородное из скота, какой у тебя будет, мужеского пола, – Господу,
EXOD|13|13|а всякого из ослов, разверзающего, заменяй агнцем; а если не заменишь, выкупи его; и каждого первенца человеческого из сынов твоих выкупай.
EXOD|13|14|И когда после спросит тебя сын твой, говоря: что это? то скажи ему: рукою крепкою вывел нас Господь из Египта, из дома рабства;
EXOD|13|15|ибо когда фараон упорствовал отпустить нас, Господь умертвил всех первенцев в земле Египетской, от первенца человеческого до первенца из скота, – посему я приношу в жертву Господу все, разверзающее ложесна, мужеского пола, а всякого первенца [из] сынов моих выкупаю;
EXOD|13|16|и да будет это знаком на руке твоей и вместо повязки над глазами твоими, ибо рукою крепкою Господь вывел нас из Египта.
EXOD|13|17|Когда же фараон отпустил народ, Бог не повел [его] по дороге земли Филистимской, потому что она близка; ибо сказал Бог: чтобы не раскаялся народ, увидев войну, и не возвратился в Египет.
EXOD|13|18|И обвел Бог народ дорогою пустынною к Чермному морю. И вышли сыны Израилевы вооруженные из земли Египетской.
EXOD|13|19|И взял Моисей с собою кости Иосифа, ибо [Иосиф] клятвою заклял сынов Израилевых, сказав: посетит вас Бог, и вы с собою вынесите кости мои отсюда.
EXOD|13|20|И двинулись [сыны Израилевы] из Сокхофа и расположились станом в Ефаме, в конце пустыни.
EXOD|13|21|Господь же шел пред ними днем в столпе облачном, показывая им путь, а ночью в столпе огненном, светя им, дабы идти им и днем и ночью.
EXOD|13|22|Не отлучался столп облачный днем и столп огненный ночью от лица народа.
EXOD|14|1|И сказал Господь Моисею, говоря:
EXOD|14|2|скажи сынам Израилевым, чтобы они обратились и расположились станом пред Пи–Гахирофом, между Мигдолом и между морем, пред Ваал–Цефоном; напротив его поставьте стан у моря.
EXOD|14|3|И скажет фараон о сынах Израилевых: они заблудились в земле сей, заперла их пустыня.
EXOD|14|4|А Я ожесточу сердце фараона, и он погонится за ними, и покажу славу Мою на фараоне и на всем войске его; и познают Египтяне, что Я Господь. И сделали так.
EXOD|14|5|И возвещено было царю Египетскому, что народ бежал; и обратилось сердце фараона и рабов его против народа сего, и они сказали: что это мы сделали? зачем отпустили Израильтян, чтобы они не работали нам?
EXOD|14|6|[Фараон] запряг колесницу свою и народ свой взял с собою;
EXOD|14|7|и взял шестьсот колесниц отборных и все колесницы Египетские, и начальников над всеми ими.
EXOD|14|8|И ожесточил Господь сердце фараона, царя Египетского, и он погнался за сынами Израилевыми; сыны же Израилевы шли под рукою высокою.
EXOD|14|9|И погнались за ними Египтяне, и все кони с колесницами фараона, и всадники, и все войско его, и настигли их расположившихся у моря, при Пи–Гахирофе пред Ваал–Цефоном.
EXOD|14|10|Фараон приблизился, и сыны Израилевы оглянулись, и вот, Египтяне идут за ними: и весьма устрашились и возопили сыны Израилевы к Господу,
EXOD|14|11|и сказали Моисею: разве нет гробов в Египте, что ты привел нас умирать в пустыне? что это ты сделал с нами, выведя нас из Египта?
EXOD|14|12|Не это ли самое говорили мы тебе в Египте, сказав: оставь нас, пусть мы работаем Египтянам? Ибо лучше быть нам в рабстве у Египтян, нежели умереть в пустыне.
EXOD|14|13|Но Моисей сказал народу: не бойтесь, стойте – и увидите спасение Господне, которое Он соделает вам ныне, ибо Египтян, которых видите вы ныне, более не увидите во веки;
EXOD|14|14|Господь будет поборать за вас, а вы будьте спокойны.
EXOD|14|15|И сказал Господь Моисею: что ты вопиешь ко Мне? скажи сынам Израилевым, чтоб они шли,
EXOD|14|16|а ты подними жезл твой и простри руку твою на море, и раздели его, и пройдут сыны Израилевы среди моря по суше;
EXOD|14|17|Я же ожесточу сердце Египтян, и они пойдут вслед за ними; и покажу славу Мою на фараоне и на всем войске его, на колесницах его и на всадниках его;
EXOD|14|18|и узнают Египтяне, что Я Господь, когда покажу славу Мою на фараоне, на колесницах его и на всадниках его.
EXOD|14|19|И двинулся Ангел Божий, шедший пред станом Израилевых, и пошел позади их; двинулся и столп облачный от лица их и стал позади их;
EXOD|14|20|и вошел в средину между станом Египетским и между станом Израилевых, и был облаком и мраком [для одних] и освещал ночь [для других], и не сблизились одни с другими во всю ночь.
EXOD|14|21|И простер Моисей руку свою на море, и гнал Господь море сильным восточным ветром всю ночь и сделал море сушею, и расступились воды.
EXOD|14|22|И пошли сыны Израилевы среди моря по суше: воды же были им стеною по правую и по левую сторону.
EXOD|14|23|Погнались Египтяне, и вошли за ними в средину моря все кони фараона, колесницы его и всадники его.
EXOD|14|24|И в утреннюю стражу воззрел Господь на стан Египтян из столпа огненного и облачного и привел в замешательство стан Египтян;
EXOD|14|25|и отнял колеса у колесниц их, так что они влекли их с трудом. И сказали Египтяне: побежим от Израильтян, потому что Господь поборает за них против Египтян.
EXOD|14|26|И сказал Господь Моисею: простри руку твою на море, и да обратятся воды на Египтян, на колесницы их и на всадников их.
EXOD|14|27|И простер Моисей руку свою на море, и к утру вода возвратилась в свое место; а Египтяне бежали на встречу [воде]. Так потопил Господь Египтян среди моря.
EXOD|14|28|И вода возвратилась и покрыла колесницы и всадников всего войска фараонова, вошедших за ними в море; не осталось ни одного из них.
EXOD|14|29|А сыны Израилевы прошли по суше среди моря: воды [были] им стеною по правую и по левую сторону.
EXOD|14|30|И избавил Господь в день тот Израильтян из рук Египтян, и увидели Израилевы Египтян мертвыми на берегу моря.
EXOD|14|31|И увидели Израильтяне руку великую, которую явил Господь над Египтянами, и убоялся народ Господа и поверил Господу и Моисею, рабу Его. Тогда Моисей и сыны Израилевы воспели Господу песнь сию и говорили:
EXOD|15|1|Пою Господу, ибо Он высоко превознесся; коня и всадника его ввергнул в море.
EXOD|15|2|Господь крепость моя и слава моя, Он был мне спасением. Он Бог мой, и прославлю Его; Бог отца моего, и превознесу Его.
EXOD|15|3|Господь муж брани, Иегова имя Ему.
EXOD|15|4|Колесницы фараона и войско его ввергнул Он в море, и избранные военачальники его потонули в Чермном море.
EXOD|15|5|Пучины покрыли их: они пошли в глубину, как камень.
EXOD|15|6|Десница Твоя, Господи, прославилась силою; десница Твоя, Господи, сразила врага.
EXOD|15|7|Величием славы Твоей Ты низложил восставших против Тебя. Ты послал гнев Твой, и он попалил их, как солому.
EXOD|15|8|От дуновения Твоего расступились воды, влага стала, как стена, огустели пучины в сердце моря.
EXOD|15|9|Враг сказал: погонюсь, настигну, разделю добычу; насытится ими душа моя, обнажу меч мой, истребит их рука моя.
EXOD|15|10|Ты дунул духом Твоим, и покрыло их море: они погрузились, как свинец, в великих водах.
EXOD|15|11|Кто, как Ты, Господи, между богами? Кто, как Ты, величествен святостью, досточтим хвалами, Творец чудес?
EXOD|15|12|Ты простер десницу Твою: поглотила их земля.
EXOD|15|13|Ты ведешь милостью Твоею народ сей, который Ты избавил, – сопровождаешь силою Твоею в жилище святыни Твоей.
EXOD|15|14|Услышали народы и трепещут: ужас объял жителей Филистимских;
EXOD|15|15|тогда смутились князья Едомовы, трепет объял вождей Моавитских, уныли все жители Ханаана.
EXOD|15|16|Да нападет на них страх и ужас; от величия мышцы Твоей да онемеют они, как камень, доколе проходит народ Твой, Господи, доколе проходит сей народ, который Ты приобрел.
EXOD|15|17|Введи его и насади его на горе достояния Твоего, на месте, которое Ты соделал жилищем Себе, Господи, во святилище, [которое] создали руки Твои, Владыка!
EXOD|15|18|Господь будет царствовать во веки и в вечность.
EXOD|15|19|Когда вошли кони фараона с колесницами его и с всадниками его в море, то Господь обратил на них воды морские, а сыны Израилевы прошли по суше среди моря.
EXOD|15|20|И взяла Мариам пророчица, сестра Ааронова, в руку свою тимпан, и вышли за нею все женщины с тимпанами и ликованием.
EXOD|15|21|И воспела Мариам пред ними: пойте Господу, ибо высоко превознесся Он, коня и всадника его ввергнул в море.
EXOD|15|22|И повел Моисей Израильтян от Чермного моря, и они вступили в пустыню Сур; и шли они три дня по пустыне и не находили воды.
EXOD|15|23|Пришли в Мерру – и не могли пить воды в Мерре, ибо она была горька, почему и наречено тому [месту] имя: Мерра.
EXOD|15|24|И возроптал народ на Моисея, говоря: что нам пить?
EXOD|15|25|[Моисей] возопил к Господу, и Господь показал ему дерево, и он бросил его в воду, и вода сделалась сладкою. Там [Бог] дал [народу] устав и закон и там испытывал его.
EXOD|15|26|И сказал: если ты будешь слушаться гласа Господа, Бога твоего, и делать угодное пред очами Его, и внимать заповедям Его, и соблюдать все уставы Его, то не наведу на тебя ни одной из болезней, которые навел Я на Египет, ибо Я Господь, целитель твой.
EXOD|15|27|И пришли в Елим; там [было] двенадцать источников воды и семьдесят финиковых дерев, и расположились там станом при водах.
EXOD|16|1|И двинулись из Елима, и пришло все общество сынов Израилевых в пустыню Син, что между Елимом и между Синаем, в пятнадцатый день второго месяца по выходе их из земли Египетской.
EXOD|16|2|И возроптало все общество сынов Израилевых на Моисея и Аарона в пустыне,
EXOD|16|3|и сказали им сыны Израилевы: о, если бы мы умерли от руки Господней в земле Египетской, когда мы сидели у котлов с мясом, когда мы ели хлеб досыта! ибо вывели вы нас в эту пустыню, чтобы все собрание это уморить голодом.
EXOD|16|4|И сказал Господь Моисею: вот, Я одождю вам хлеб с неба, и пусть народ выходит и собирает ежедневно, сколько нужно на день, чтобы Мне испытать его, будет ли он поступать по закону Моему, или нет;
EXOD|16|5|а в шестой день пусть заготовляют, что принесут, и будет вдвое против того, по скольку собирают в прочие дни.
EXOD|16|6|И сказали Моисей и Аарон всему [обществу] сынов Израилевых: вечером узнаете вы, что Господь вывел вас из земли Египетской,
EXOD|16|7|и утром увидите славу Господню, ибо услышал Он ропот ваш на Господа: а мы что такое, что ропщете на нас?
EXOD|16|8|И сказал Моисей: [узнаете], когда Господь вечером даст вам мяса в пищу, а утром хлеба досыта, ибо Господь услышал ропот ваш, который вы подняли против Него: а мы что? не на нас ропот ваш, но на Господа.
EXOD|16|9|И сказал Моисей Аарону: скажи всему обществу сынов Израилевых: предстаньте пред лице Господа, ибо Он услышал ропот ваш.
EXOD|16|10|И когда говорил Аарон ко всему обществу сынов Израилевых, то они оглянулись к пустыне, и вот, слава Господня явилась в облаке.
EXOD|16|11|И сказал Господь Моисею, говоря:
EXOD|16|12|Я услышал ропот сынов Израилевых; скажи им: вечером будете есть мясо, а поутру насытитесь хлебом – и узнаете, что Я Господь, Бог ваш.
EXOD|16|13|Вечером налетели перепелы и покрыли стан, а поутру лежала роса около стана;
EXOD|16|14|роса поднялась, и вот, на поверхности пустыни [нечто] мелкое, круповидное, мелкое, как иней на земле.
EXOD|16|15|И увидели сыны Израилевы и говорили друг другу: что это? Ибо не знали, что это. И Моисей сказал им: это хлеб, который Господь дал вам в пищу;
EXOD|16|16|вот что повелел Господь: собирайте его каждый по стольку, сколько ему съесть; по гомору на человека, по числу душ, сколько у кого в шатре, собирайте.
EXOD|16|17|И сделали так сыны Израилевы и собрали, кто много, кто мало;
EXOD|16|18|и меряли гомором, и у того, кто собрал много, не было лишнего, и у того, кто мало, не было недостатка: каждый собрал, сколько ему съесть.
EXOD|16|19|И сказал им Моисей: никто не оставляй сего до утра.
EXOD|16|20|Но не послушали они Моисея, и оставили от сего некоторые до утра, – и завелись черви, и оно воссмердело. И разгневался на них Моисей.
EXOD|16|21|И собирали его рано поутру, каждый сколько ему съесть; когда же обогревало солнце, оно таяло.
EXOD|16|22|В шестой же день собрали хлеба вдвое, по два гомора на каждого. И пришли все начальники общества и донесли Моисею.
EXOD|16|23|И [он] сказал им: вот что сказал Господь: завтра покой, святая суббота Господня; что надобно печь, пеките, и что надобно варить, варите [сегодня], а что останется, отложите и сберегите до утра.
EXOD|16|24|И отложили то до утра, как повелел Моисей, и оно не воссмердело, и червей не было в нем.
EXOD|16|25|И сказал Моисей: ешьте его сегодня, ибо сегодня суббота Господня; сегодня не найдете его на поле;
EXOD|16|26|шесть дней собирайте его, а в седьмой день – суббота: не будет его в [этот день].
EXOD|16|27|[Но некоторые] из народа вышли в седьмой день собирать – и не нашли.
EXOD|16|28|И сказал Господь Моисею: долго ли будете вы уклоняться от соблюдения заповедей Моих и законов Моих?
EXOD|16|29|смотрите, Господь дал вам субботу, посему Он и дает в шестой день хлеба на два дня: оставайтесь каждый у себя, никто не выходи от места своего в седьмой день.
EXOD|16|30|И покоился народ в седьмой день.
EXOD|16|31|И нарек дом Израилев [хлебу] тому имя: манна; она была, как кориандровое семя, белая, вкусом же как лепешка с медом.
EXOD|16|32|И сказал Моисей: вот что повелел Господь: наполните [манною] гомор для хранения в роды ваши, дабы видели хлеб, которым Я питал вас в пустыне, когда вывел вас из земли Египетской.
EXOD|16|33|И сказал Моисей Аарону: возьми один сосуд, и положи в него полный гомор манны, и поставь его пред Господом, для хранения в роды ваши.
EXOD|16|34|И поставил его Аарон пред ковчегом свидетельства для хранения, как повелел Господь Моисею.
EXOD|16|35|Сыны Израилевы ели манну сорок лет, доколе не пришли в землю обитаемую; манну ели они, доколе не пришли к пределам земли Ханаанской.
EXOD|16|36|А гомор есть десятая часть ефы.
EXOD|17|1|И двинулось все общество сынов Израилевых из пустыни Син в путь свой, по повелению Господню, и расположилось станом в Рефидиме, и не было воды пить народу.
EXOD|17|2|И укорял народ Моисея, и говорили: дайте нам воды пить. И сказал им Моисей: что вы укоряете меня? что искушаете Господа?
EXOD|17|3|И жаждал там народ воды, и роптал народ на Моисея, говоря: зачем ты вывел нас из Египта, уморить жаждою нас и детей наших и стада наши?
EXOD|17|4|Моисей возопил к Господу и сказал: что мне делать с народом сим? еще немного, и побьют меня камнями.
EXOD|17|5|И сказал Господь Моисею: пройди перед народом, и возьми с собою [некоторых] из старейшин Израильских, и жезл твой, которым ты ударил по воде, возьми в руку твою, и пойди;
EXOD|17|6|вот, Я стану пред тобою там на скале в Хориве, и ты ударишь в скалу, и пойдет из нее вода, и будет пить народ. И сделал так Моисей в глазах старейшин Израильских.
EXOD|17|7|И нарек месту тому имя: Масса и Мерива, по причине укорения сынов Израилевых и потому, что они искушали Господа, говоря: есть ли Господь среди нас, или нет?
EXOD|17|8|И пришли Амаликитяне и воевали с Израильтянами в Рефидиме.
EXOD|17|9|Моисей сказал Иисусу: выбери нам мужей, и пойди, сразись с Амаликитянами; завтра я стану на вершине холма, и жезл Божий будет в руке моей.
EXOD|17|10|И сделал Иисус, как сказал ему Моисей, и [пошел] сразиться с Амаликитянами; а Моисей и Аарон и Ор взошли на вершину холма.
EXOD|17|11|И когда Моисей поднимал руки свои, одолевал Израиль, а когда опускал руки свои, одолевал Амалик;
EXOD|17|12|но руки Моисеевы отяжелели, и тогда взяли камень и подложили под него, и он сел на нем, Аарон же и Ор поддерживали руки его, один с одной, а другой с другой [стороны]. И были руки его подняты до захождения солнца.
EXOD|17|13|И низложил Иисус Амалика и народ его острием меча.
EXOD|17|14|И сказал Господь Моисею: напиши сие для памяти в книгу и внуши Иисусу, что Я совершенно изглажу память Амаликитян из поднебесной.
EXOD|17|15|И устроил Моисей жертвенник и нарек ему имя: Иегова Нисси.
EXOD|17|16|Ибо, сказал он, рука на престоле Господа: брань у Господа против Амалика из рода в род.
EXOD|18|1|И услышал Иофор, священник Мадиамский, тесть Моисеев, о всем, что сделал Бог для Моисея и для Израиля, народа Своего, когда вывел Господь Израиля из Египта,
EXOD|18|2|и взял Иофор, тесть Моисеев, Сепфору, жену Моисееву, пред тем возвращенную,
EXOD|18|3|и двух сынов ее, из которых одному имя Гирсам, потому что говорил [Моисей]: я пришлец в земле чужой;
EXOD|18|4|а другому имя Елиезер, потому что [говорил он] Бог отца моего был мне помощником и избавил меня от меча фараонова.
EXOD|18|5|И пришел Иофор, тесть Моисея, с сыновьями его и женою его к Моисею в пустыню, где он расположился станом у горы Божией,
EXOD|18|6|и дал знать Моисею: я, тесть твой Иофор, иду к тебе, и жена твоя, и два сына ее с нею.
EXOD|18|7|Моисей вышел навстречу тестю своему, и поклонился, и целовал его, и после взаимного приветствия они вошли в шатер.
EXOD|18|8|И рассказал Моисей тестю своему о всем, что сделал Господь с фараоном и с Египтянами за Израиля, и о всех трудностях, какие встретили их на пути, и как избавил их Господь.
EXOD|18|9|Иофор радовался о всех благодеяниях, которые Господь явил Израилю, когда избавил его из руки Египтян.
EXOD|18|10|и сказал Иофор: благословен Господь, Который избавил вас из руки Египтян и из руки фараоновой, Который избавил народ сей из–под власти Египтян;
EXOD|18|11|ныне узнал я, что Господь велик паче всех богов, в том самом, чем они превозносились над [Израильтянами].
EXOD|18|12|И принес Иофор, тесть Моисеев, всесожжение и жертвы Богу; и пришел Аарон и все старейшины Израилевы есть хлеба с тестем Моисеевым пред Богом.
EXOD|18|13|На другой день сел Моисей судить народ, и стоял народ пред Моисеем с утра до вечера.
EXOD|18|14|И видел тесть Моисеев, все, что он делает с народом, и сказал: что это такое делаешь ты с народом? для чего ты сидишь один, а весь народ стоит пред тобою с утра до вечера?
EXOD|18|15|И сказал Моисей тестю своему: народ приходит ко мне просить суда у Бога;
EXOD|18|16|когда случается у них какое дело, они приходят ко мне, и я сужу между тем и другим и объявляю уставы Божии и законы Его.
EXOD|18|17|Но тесть Моисеев сказал ему: не хорошо это ты делаешь:
EXOD|18|18|ты измучишь и себя и народ сей, который с тобою, ибо слишком тяжело для тебя это дело: ты один не можешь исправлять его;
EXOD|18|19|итак послушай слов моих; я дам тебе совет, и будет Бог с тобою: будь ты для народа посредником пред Богом и представляй Богу дела [его];
EXOD|18|20|научай их уставам и законам [Божиим], указывай им путь [Его], по которому они должны идти, и дела, которые они должны делать;
EXOD|18|21|ты же усмотри из всего народа людей способных, боящихся Бога, людей правдивых, ненавидящих корысть, и поставь [их] над ним тысяченачальниками, стоначальниками, пятидесятиначальниками и десятиначальниками;
EXOD|18|22|пусть они судят народ во всякое время и о всяком важном деле доносят тебе, а все малые дела судят сами: и будет тебе легче, и они понесут с тобою [бремя];
EXOD|18|23|если ты сделаешь это, и Бог повелит тебе, то ты можешь устоять, и весь народ сей будет отходить в свое место с миром.
EXOD|18|24|И послушал Моисей слов тестя своего и сделал все, что он говорил;
EXOD|18|25|и выбрал Моисей из всего Израиля способных людей и поставил их начальниками народа, тысяченачальниками, стоначальниками, пятидесятиначальниками и десятиначальниками.
EXOD|18|26|и судили они народ во всякое время; о делах важных доносили Моисею, а все малые дела судили сами.
EXOD|18|27|И отпустил Моисей тестя своего, и он пошел в землю свою.
EXOD|19|1|В третий месяц по исходе сынов Израиля из земли Египетской, в самый день новолуния, пришли они в пустыню Синайскую.
EXOD|19|2|И двинулись они из Рефидима, и пришли в пустыню Синайскую, и расположились там станом в пустыне; и расположился там Израиль станом против горы.
EXOD|19|3|Моисей взошел к Богу [на гору], и воззвал к нему Господь с горы, говоря: так скажи дому Иаковлеву и возвести сынам Израилевым:
EXOD|19|4|вы видели, что Я сделал Египтянам, и как Я носил вас [как бы] на орлиных крыльях, и принес вас к Себе;
EXOD|19|5|итак, если вы будете слушаться гласа Моего и соблюдать завет Мой, то будете Моим уделом из всех народов, ибо Моя вся земля,
EXOD|19|6|а вы будете у Меня царством священников и народом святым; вот слова, которые ты скажешь сынам Израилевым.
EXOD|19|7|И пришел Моисей и созвал старейшин народа и предложил им все сии слова, которые заповедал ему Господь.
EXOD|19|8|И весь народ отвечал единогласно, говоря: все, что сказал Господь, исполним. И донес Моисей слова народа Господу.
EXOD|19|9|И сказал Господь Моисею: вот, Я приду к тебе в густом облаке, дабы слышал народ, как Я буду говорить с тобою, и поверил тебе навсегда. И Моисей объявил слова народа Господу.
EXOD|19|10|И сказал Господь Моисею: пойди к народу, и освяти его сегодня и завтра; пусть вымоют одежды свои,
EXOD|19|11|чтоб быть готовыми к третьему дню: ибо в третий день сойдет Господь пред глазами всего народа на гору Синай;
EXOD|19|12|и проведи для народа черту со всех сторон и скажи: берегитесь восходить на гору и прикасаться к подошве ее; всякий, кто прикоснется к горе, предан будет смерти;
EXOD|19|13|рука да не прикоснется к нему, а пусть побьют его камнями, или застрелят стрелою; скот ли то, или человек, да не останется в живых; во время протяжного трубного звука могут они взойти на гору.
EXOD|19|14|И сошел Моисей с горы к народу и освятил народ, и они вымыли одежду свою.
EXOD|19|15|И сказал народу: будьте готовы к третьему дню; не прикасайтесь к женам.
EXOD|19|16|На третий день, при наступлении утра, были громы и молнии, и густое облако над горою, и трубный звук весьма сильный; и вострепетал весь народ, бывший в стане.
EXOD|19|17|И вывел Моисей народ из стана в сретение Богу, и стали у подошвы горы.
EXOD|19|18|Гора же Синай вся дымилась от того, что Господь сошел на нее в огне; и восходил от нее дым, как дым из печи, и вся гора сильно колебалась;
EXOD|19|19|и звук трубный становился сильнее и сильнее. Моисей говорил, и Бог отвечал ему голосом.
EXOD|19|20|И сошел Господь на гору Синай, на вершину горы, и призвал Господь Моисея на вершину горы, и взошел Моисей.
EXOD|19|21|И сказал Господь Моисею: сойди и подтверди народу, чтобы он не порывался к Господу видеть [Его], и чтобы не пали многие из него;
EXOD|19|22|священники же, приближающиеся к Господу, должны освятить себя, чтобы не поразил их Господь.
EXOD|19|23|И сказал Моисей Господу: не может народ взойти на гору Синай, потому что Ты предостерег нас, сказав: проведи черту вокруг горы и освяти ее.
EXOD|19|24|И Господь сказал ему: пойди, сойди, потом взойди ты и с тобою Аарон; а священники и народ да не порываются восходить к Господу, чтобы не поразил их.
EXOD|19|25|И сошел Моисей к народу и пересказал ему.
EXOD|20|1|И изрек Бог все слова сии, говоря:
EXOD|20|2|Я Господь, Бог твой, Который вывел тебя из земли Египетской, из дома рабства;
EXOD|20|3|да не будет у тебя других богов пред лицем Моим.
EXOD|20|4|Не делай себе кумира и никакого изображения того, что на небе вверху, и что на земле внизу, и что в воде ниже земли;
EXOD|20|5|не поклоняйся им и не служи им, ибо Я Господь, Бог твой, Бог ревнитель, наказывающий детей за вину отцов до третьего и четвертого [рода], ненавидящих Меня,
EXOD|20|6|и творящий милость до тысячи родов любящим Меня и соблюдающим заповеди Мои.
EXOD|20|7|Не произноси имени Господа, Бога твоего, напрасно, ибо Господь не оставит без наказания того, кто произносит имя Его напрасно.
EXOD|20|8|Помни день субботний, чтобы святить его;
EXOD|20|9|шесть дней работай и делай всякие дела твои,
EXOD|20|10|а день седьмой – суббота Господу, Богу твоему: не делай в оный никакого дела ни ты, ни сын твой, ни дочь твоя, ни раб твой, ни рабыня твоя, ни скот твой, ни пришлец, который в жилищах твоих;
EXOD|20|11|ибо в шесть дней создал Господь небо и землю, море и все, что в них, а в день седьмой почил; посему благословил Господь день субботний и освятил его.
EXOD|20|12|Почитай отца твоего и мать твою, чтобы продлились дни твои на земле, которую Господь, Бог твой, дает тебе.
EXOD|20|13|Не убивай.
EXOD|20|14|Не прелюбодействуй.
EXOD|20|15|Не кради.
EXOD|20|16|Не произноси ложного свидетельства на ближнего твоего.
EXOD|20|17|Не желай дома ближнего твоего; не желай жены ближнего твоего, ни раба его, ни рабыни его, ни вола его, ни осла его, ничего, что у ближнего твоего.
EXOD|20|18|Весь народ видел громы и пламя, и звук трубный, и гору дымящуюся; и увидев [то], народ отступил и стал вдали.
EXOD|20|19|И сказали Моисею: говори ты с нами, и мы будем слушать, но чтобы не говорил с нами Бог, дабы нам не умереть.
EXOD|20|20|И сказал Моисей народу: не бойтесь; Бог пришел, чтобы испытать вас и чтобы страх Его был пред лицем вашим, дабы вы не грешили.
EXOD|20|21|И стоял народ вдали, а Моисей вступил во мрак, где Бог.
EXOD|20|22|И сказал Господь Моисею: так скажи сынам Израилевым: вы видели, как Я с неба говорил вам;
EXOD|20|23|не делайте предо Мною богов серебряных, или богов золотых, не делайте себе:
EXOD|20|24|сделай Мне жертвенник из земли и приноси на нем всесожжения твои и мирные жертвы твои, овец твоих и волов твоих; на всяком месте, где Я положу память имени Моего, Я приду к тебе и благословлю тебя;
EXOD|20|25|если же будешь делать Мне жертвенник из камней, то не сооружай его из тесаных, ибо, как скоро наложишь на них тесло твое, то осквернишь их;
EXOD|20|26|и не всходи по ступеням к жертвеннику Моему, дабы не открылась при нем нагота твоя.
EXOD|21|1|И вот законы, которые ты объявишь им:
EXOD|21|2|если купишь раба Еврея, пусть он работает шесть лет, а в седьмой пусть выйдет на волю даром;
EXOD|21|3|если он пришел один, пусть один и выйдет; а если он женатый, пусть выйдет с ним и жена его;
EXOD|21|4|если же господин его дал ему жену и она родила ему сынов, или дочерей, то жена и дети ее пусть останутся у господина ее, а он выйдет один;
EXOD|21|5|но если раб скажет: люблю господина моего, жену мою и детей моих, не пойду на волю, –
EXOD|21|6|то пусть господин его приведет его пред богов и поставит его к двери, или к косяку, и проколет ему господин его ухо шилом, и он останется рабом его вечно.
EXOD|21|7|Если кто продаст дочь свою в рабыни, то она не может выйти, как выходят рабы;
EXOD|21|8|если она не угодна господину своему и он не обручит ее, пусть позволит выкупить ее; а чужому народу продать ее не властен, когда сам пренебрег ее;
EXOD|21|9|если он обручит ее сыну своему, пусть поступит с нею по праву дочерей;
EXOD|21|10|если же другую возьмет за него, то она не должна лишаться пищи, одежды и супружеского сожития;
EXOD|21|11|а если он сих трех [вещей] не сделает для нее, пусть она отойдет даром, без выкупа.
EXOD|21|12|Кто ударит человека так, что он умрет, да будет предан смерти;
EXOD|21|13|но если кто не злоумышлял, а Бог попустил ему попасть под руки его, то Я назначу у тебя место, куда убежать [убийце];
EXOD|21|14|а если кто с намерением умертвит ближнего коварно, то [и] от жертвенника Моего бери его на смерть.
EXOD|21|15|Кто ударит отца своего, или свою мать, того должно предать смерти.
EXOD|21|16|Кто украдет человека и продаст его, или найдется он в руках у него, то должно предать его смерти.
EXOD|21|17|Кто злословит отца своего, или свою мать, того должно предать смерти.
EXOD|21|18|Когда ссорятся, и один человек ударит другого камнем, или кулаком, и тот не умрет, но сляжет в постель,
EXOD|21|19|то, если он встанет и будет выходить из дома с помощью палки, ударивший не будет повинен [смерти]; только пусть заплатит за остановку в его работе и даст на лечение его.
EXOD|21|20|А если кто ударит раба своего, или служанку свою палкою, и они умрут под рукою его, то он должен быть наказан;
EXOD|21|21|но если они день или два дня переживут, то не должно наказывать его, ибо это его серебро.
EXOD|21|22|Когда дерутся люди, и ударят беременную женщину, и она выкинет, но не будет [другого] вреда, то взять с [виновного] пеню, какую наложит на него муж той женщины, и он должен заплатить оную при посредниках;
EXOD|21|23|а если будет вред, то отдай душу за душу,
EXOD|21|24|глаз за глаз, зуб за зуб, руку за руку, ногу за ногу,
EXOD|21|25|обожжение за обожжение, рану за рану, ушиб за ушиб.
EXOD|21|26|Если кто раба своего ударит в глаз, или служанку свою в глаз, и повредит его, пусть отпустит их на волю за глаз;
EXOD|21|27|и если выбьет зуб рабу своему, или рабе своей, пусть отпустит их на волю за зуб.
EXOD|21|28|Если вол забодает мужчину или женщину до смерти, то вола побить камнями и мяса его не есть; а хозяин вола не виноват;
EXOD|21|29|но если вол бодлив был и вчера и третьего дня, и хозяин его, быв извещен о сем, не стерег его, а он убил мужчину или женщину, то вола побить камнями, и хозяина его предать смерти;
EXOD|21|30|если на него наложен будет выкуп, пусть даст выкуп за душу свою, какой наложен будет на него.
EXOD|21|31|Сына ли забодает, дочь ли забодает, – по сему же закону поступать с ним.
EXOD|21|32|Если вол забодает раба или рабу, то господину их заплатить тридцать сиклей серебра, а вола побить камнями.
EXOD|21|33|Если кто раскроет яму, или если выкопает яму и не покроет ее, и упадет в нее вол или осел,
EXOD|21|34|то хозяин ямы должен заплатить, отдать серебро хозяину их, а труп будет его.
EXOD|21|35|Если чей–нибудь вол забодает до смерти вола у соседа его, пусть продадут живого вола и разделят пополам цену его; также и убитого пусть разделят пополам;
EXOD|21|36|а если известно было, что вол бодлив был и вчера и третьего дня, но хозяин его не стерег его, то должен он заплатить вола за вола, а убитый будет его.
EXOD|21|37|Если кто украдет вола или овцу и заколет или продаст, то пять волов заплатит за вола и четыре овцы за овцу.
EXOD|22|1|Если [кто] застанет вора подкапывающего и ударит его, так что он умрет, то кровь не [вменится] ему;
EXOD|22|2|но если взошло над ним солнце, то [вменится] ему кровь. [Укравший] должен заплатить; а если нечем, то пусть продадут его [для уплаты] за украденное им;
EXOD|22|3|если украденное найдется у него в руках живым, вол ли то, или осел, или овца, пусть заплатит вдвое.
EXOD|22|4|Если кто потравит поле, или виноградник, пустив скот свой травить чужое поле, пусть вознаградит лучшим из поля своего и лучшим из виноградника своего.
EXOD|22|5|Если появится огонь и охватит терн и выжжет копны, или жатву, или поле, то должен заплатить, кто произвел сей пожар.
EXOD|22|6|Если кто отдаст ближнему на сохранение серебро или вещи, и они украдены будут из дома его, то, если найдется вор, пусть он заплатит вдвое;
EXOD|22|7|а если не найдется вор, пусть хозяин дома придет пред судей [и поклянется], что не простер руки своей на собственность ближнего своего.
EXOD|22|8|О всякой вещи спорной, о воле, об осле, об овце, об одежде, о всякой вещи потерянной, о которой кто–нибудь скажет, что она его, дело обоих должно быть доведено до судей: кого обвинят судьи, тот заплатит ближнему своему вдвое.
EXOD|22|9|Если кто отдаст ближнему своему осла, или вола, или овцу, или какой другой скот на сбережение, а он умрет, или будет поврежден, или уведен, так что никто сего не увидит, –
EXOD|22|10|клятва пред Господом да будет между обоими в том, что [взявший] не простер руки своей на собственность ближнего своего; и хозяин должен принять, а [тот] не будет платить;
EXOD|22|11|а если украден будет у него, то должен заплатить хозяину его;
EXOD|22|12|если же будет [зверем] растерзан, то пусть в доказательство представит растерзанное: за растерзанное он не платит.
EXOD|22|13|Если кто займет у ближнего своего скот, и он будет поврежден, или умрет, а хозяина его не было при нем, то должен заплатить;
EXOD|22|14|если же хозяин его был при нем, то не должен платить; если он взят был в наймы за деньги, то пусть и пойдет за ту цену.
EXOD|22|15|Если обольстит кто девицу необрученную и переспит с нею, пусть даст ей вено [и возьмет ее] себе в жену;
EXOD|22|16|а если отец не согласится выдать ее за него, пусть заплатит [столько] серебра, сколько [полагается] на вено девицам.
EXOD|22|17|Ворожеи не оставляй в живых.
EXOD|22|18|Всякий скотоложник да будет предан смерти.
EXOD|22|19|Приносящий жертву богам, кроме одного Господа, да будет истреблен.
EXOD|22|20|Пришельца не притесняй и не угнетай его, ибо вы сами были пришельцами в земле Египетской.
EXOD|22|21|Ни вдовы, ни сироты не притесняйте;
EXOD|22|22|если же ты притеснишь их, то, когда они возопиют ко Мне, Я услышу вопль их,
EXOD|22|23|и воспламенится гнев Мой, и убью вас мечом, и будут жены ваши вдовами и дети ваши сиротами.
EXOD|22|24|Если дашь деньги взаймы бедному из народа Моего, то не притесняй его и не налагай на него роста.
EXOD|22|25|Если возьмешь в залог одежду ближнего твоего, до захождения солнца возврати ее,
EXOD|22|26|ибо она есть единственный покров у него, она – одеяние тела его: в чем будет он спать? итак, когда он возопиет ко Мне, Я услышу, ибо Я милосерд.
EXOD|22|27|Судей не злословь и начальника в народе твоем не поноси.
EXOD|22|28|Не медли [приносить Мне] начатки от гумна твоего и от точила твоего; отдавай Мне первенца из сынов твоих;
EXOD|22|29|то же делай с волом твоим и с овцою твоею. семь дней пусть они будут при матери своей, а в восьмой день отдавай их Мне.
EXOD|22|30|И будете у Меня людьми святыми; и мяса, растерзанного зверем в поле, не ешьте, псам бросайте его.
EXOD|23|1|Не внимай пустому слуху, не давай руки твоей нечестивому, чтоб быть свидетелем неправды.
EXOD|23|2|Не следуй за большинством на зло, и не решай тяжбы, отступая по большинству от правды;
EXOD|23|3|и бедному не потворствуй в тяжбе его.
EXOD|23|4|Если найдешь вола врага твоего, или осла его заблудившегося, приведи его к нему;
EXOD|23|5|если увидишь осла врага твоего упавшим под ношею своею, то не оставляй его; развьючь вместе с ним.
EXOD|23|6|Не суди превратно тяжбы бедного твоего.
EXOD|23|7|Удаляйся от неправды и не умерщвляй невинного и правого, ибо Я не оправдаю беззаконника.
EXOD|23|8|Даров не принимай, ибо дары слепыми делают зрячих и превращают дело правых.
EXOD|23|9|Пришельца не обижай: вы знаете душу пришельца, потому что сами были пришельцами в земле Египетской.
EXOD|23|10|Шесть лет засевай землю твою и собирай произведения ее,
EXOD|23|11|а в седьмой оставляй ее в покое, чтобы питались убогие из твоего народа, а остатками после них питались звери полевые; так же поступай с виноградником твоим и с маслиною твоею.
EXOD|23|12|Шесть дней делай дела твои, а в седьмой день покойся, чтобы отдохнул вол твой и осел твой и успокоился сын рабы твоей и пришлец.
EXOD|23|13|Соблюдайте все, что Я сказал вам, и имени других богов не упоминайте; да не слышится оно из уст твоих.
EXOD|23|14|Три раза в году празднуй Мне:
EXOD|23|15|наблюдай праздник опресноков: семь дней ешь пресный хлеб, как Я повелел тебе, в назначенное время месяца Авива, ибо в оном ты вышел из Египта; и пусть не являются пред лице Мое с пустыми [руками];
EXOD|23|16|[наблюдай] и праздник жатвы первых плодов труда твоего, какие ты сеял на поле, и праздник собирания плодов в конце года, когда уберешь с поля работу твою.
EXOD|23|17|Три раза в году должен являться весь мужеский пол твой пред лице Владыки, Господа.
EXOD|23|18|не изливай крови жертвы Моей на квасное, и тук от праздничной жертвы Моей не должен оставаться до утра.
EXOD|23|19|Начатки плодов земли твоей приноси в дом Господа, Бога твоего. Не вари козленка в молоке матери его.
EXOD|23|20|Вот, Я посылаю пред тобою Ангела хранить тебя на пути и ввести тебя в то место, которое Я приготовил.
EXOD|23|21|блюди себя пред лицем Его и слушай гласа Его; не упорствуй против Него, потому что Он не простит греха вашего, ибо имя Мое в Нем.
EXOD|23|22|Если ты будешь слушать гласа Его и исполнять все, что скажу, то врагом буду врагов твоих и противником противников твоих.
EXOD|23|23|Когда пойдет пред тобою Ангел Мой и поведет тебя к Аморреям, Хеттеям, Ферезеям, Хананеям, Евеям и Иевусеям, и истреблю их:
EXOD|23|24|то не поклоняйся богам их, и не служи им, и не подражай делам их, но сокруши их и разрушь столбы их:
EXOD|23|25|служите Господу, Богу вашему, и Он благословит хлеб твой и воду твою; и отвращу от вас болезни.
EXOD|23|26|Не будет преждевременно рождающих и бесплодных в земле твоей; число дней твоих сделаю полным.
EXOD|23|27|Ужас Мой пошлю пред тобою, и в смущение приведу всякий народ, к которому ты придешь, и буду обращать к тебе тыл всех врагов твоих;
EXOD|23|28|пошлю пред тобою шершней, и они погонят от лица твоего Евеев, Хананеев и Хеттеев;
EXOD|23|29|не выгоню их от лица твоего в один год, чтобы земля не сделалась пуста и не умножились против тебя звери полевые:
EXOD|23|30|мало–помалу буду прогонять их от тебя, доколе ты не размножишься и не возьмешь во владение земли сей.
EXOD|23|31|Проведу пределы твои от моря Чермного до моря Филистимского и от пустыни до реки; ибо предам в руки ваши жителей сей земли, и прогонишь их от лица твоего;
EXOD|23|32|не заключай союза ни с ними, ни с богами их;
EXOD|23|33|не должны они жить в земле твоей, чтобы они не ввели тебя в грех против Меня; ибо если ты будешь служить богам их, то это будет тебе сетью.
EXOD|24|1|И Моисею сказал Он: взойди к Господу ты и Аарон, Надав и Авиуд и семьдесят из старейшин Израилевых, и поклонитесь издали;
EXOD|24|2|Моисей один пусть приблизится к Господу, а они пусть не приближаются, и народ пусть не восходит с ним.
EXOD|24|3|И пришел Моисей и пересказал народу все слова Господни и все законы. И отвечал весь народ в один голос, и сказали: все, что сказал Господь, сделаем.
EXOD|24|4|И написал Моисей все слова Господни и, встав рано поутру, поставил под горою жертвенник и двенадцать камней, по [числу] двенадцати колен Израилевых;
EXOD|24|5|и послал юношей из сынов Израилевых, и принесли они всесожжения, и заклали тельцов в мирную жертву Господу.
EXOD|24|6|Моисей, взяв половину крови, влил в чаши, а [другою] половиною окропил жертвенник;
EXOD|24|7|и взял книгу завета и прочитал вслух народу, и сказали они: все, что сказал Господь, сделаем и будем послушны.
EXOD|24|8|И взял Моисей крови и окропил народ, говоря: вот кровь завета, который Господь заключил с вами о всех словах сих.
EXOD|24|9|Потом взошел Моисей и Аарон, Надав и Авиуд и семьдесят из старейшин Израилевых,
EXOD|24|10|и видели Бога Израилева; и под ногами Его нечто подобное работе из чистого сапфира и, как самое небо, ясное.
EXOD|24|11|И Он не простер руки Своей на избранных из сынов Израилевых: они видели Бога, и ели и пили.
EXOD|24|12|И сказал Господь Моисею: взойди ко Мне на гору и будь там; и дам тебе скрижали каменные, и закон и заповеди, которые Я написал для научения их.
EXOD|24|13|И встал Моисей с Иисусом, служителем своим, и пошел Моисей на гору Божию,
EXOD|24|14|а старейшинам сказал: оставайтесь здесь, доколе мы не возвратимся к вам; вот Аарон и Ор с вами; кто будет иметь дело, пусть приходит к ним.
EXOD|24|15|И взошел Моисей на гору, и покрыло облако гору,
EXOD|24|16|и слава Господня осенила гору Синай; и покрывало ее облако шесть дней, а в седьмой день [Господь] воззвал к Моисею из среды облака.
EXOD|24|17|Вид же славы Господней на вершине горы был пред глазами сынов Израилевых, как огонь поядающий.
EXOD|24|18|Моисей вступил в средину облака и взошел на гору; и был Моисей на горе сорок дней и сорок ночей.
EXOD|25|1|И сказал Господь Моисею, говоря:
EXOD|25|2|скажи сынам Израилевым, чтобы они сделали Мне приношения; от всякого человека, у которого будет усердие, принимайте приношения Мне.
EXOD|25|3|Вот приношения, которые вы должны принимать от них: золото и серебро и медь,
EXOD|25|4|и [шерсть] голубую, пурпуровую и червленую, и виссон, и козью,
EXOD|25|5|и кожи бараньи красные, и кожи синие, и дерева ситтим,
EXOD|25|6|елей для светильника, ароматы для елея помазания и для благовонного курения,
EXOD|25|7|камень оникс и камни вставные для ефода и для наперсника.
EXOD|25|8|И устроят они Мне святилище, и буду обитать посреди их;
EXOD|25|9|все, как Я показываю тебе, и образец скинии и образец всех сосудов ее; так и сделайте.
EXOD|25|10|Сделайте ковчег из дерева ситтим: длина ему два локтя с половиною, и ширина ему полтора локтя, и высота ему полтора локтя;
EXOD|25|11|и обложи его чистым золотом, изнутри и снаружи покрой его; и сделай наверху вокруг его золотой венец.
EXOD|25|12|и вылей для него четыре кольца золотых и утверди на четырех нижних углах его: два кольца на одной стороне его, два кольца на другой стороне его.
EXOD|25|13|Сделай из дерева ситтим шесты и обложи их золотом;
EXOD|25|14|и вложи шесты в кольца, по сторонам ковчега, чтобы посредством их носить ковчег;
EXOD|25|15|в кольцах ковчега должны быть шесты и не должны отниматься от него.
EXOD|25|16|И положи в ковчег откровение, которое Я дам тебе.
EXOD|25|17|Сделай также крышку из чистого золота: длина ее два локтя с половиною, а ширина ее полтора локтя;
EXOD|25|18|и сделай из золота двух херувимов: чеканной работы сделай их на обоих концах крышки;
EXOD|25|19|сделай одного херувима с одного края, а другого херувима с другого края; [выдавшимися] из крышки сделайте херувимов на обоих краях ее;
EXOD|25|20|и будут херувимы с распростертыми вверх крыльями, покрывая крыльями своими крышку, а лицами своими [будут] друг к другу: к крышке будут лица херувимов.
EXOD|25|21|И положи крышку на ковчег сверху, в ковчег же положи откровение, которое Я дам тебе;
EXOD|25|22|там Я буду открываться тебе и говорить с тобою над крышкою, посреди двух херувимов, которые над ковчегом откровения, о всем, что ни буду заповедывать чрез тебя сынам Израилевым.
EXOD|25|23|И сделай стол из дерева ситтим, длиною в два локтя, шириною в локоть, и вышиною в полтора локтя,
EXOD|25|24|и обложи его золотом чистым, и сделай вокруг него золотой венец.
EXOD|25|25|и сделай вокруг него стенки в ладонь и у стенок его сделай золотой венец вокруг;
EXOD|25|26|и сделай для него четыре кольца золотых и утверди кольца на четырех углах у четырех ножек его;
EXOD|25|27|при стенках должны быть кольца, чтобы влагать шесты, для ношения на них стола;
EXOD|25|28|а шесты сделай из дерева ситтим и обложи их золотом, и будут носить на них сей стол;
EXOD|25|29|сделай также для него блюдо, кадильницы, чаши и кружки, чтобы возливать ими: из золота чистого сделай их;
EXOD|25|30|и полагай на стол хлебы предложения пред лицем Моим постоянно.
EXOD|25|31|И сделай светильник из золота чистого; чеканный должен быть сей светильник; стебель его, ветви его, чашечки его, яблоки его и цветы его должны выходить из него;
EXOD|25|32|шесть ветвей должны выходить из боков его: три ветви светильника из одного бока его и три ветви светильника из другого бока его;
EXOD|25|33|три чашечки наподобие миндального цветка, с яблоком и цветами, должны быть на одной ветви, и три чашечки наподобие миндального цветка на другой ветви, с яблоком и цветами: так на [всех] шести ветвях, выходящих из светильника;
EXOD|25|34|а на [стебле] светильника должны быть четыре чашечки наподобие миндального цветка с яблоками и цветами;
EXOD|25|35|у шести ветвей, выходящих из [стебля] светильника, яблоко под двумя ветвями его, и яблоко под другими двумя ветвями, и яблоко под [третьими] двумя ветвями его.
EXOD|25|36|яблоки и ветви их из него должны выходить: он весь [должен] [быть] чеканный, цельный, из чистого золота.
EXOD|25|37|И сделай к нему семь лампад и поставь на него лампады его, чтобы светили на переднюю сторону его;
EXOD|25|38|и щипцы к нему и лотки к нему из чистого золота;
EXOD|25|39|из таланта золота чистого пусть сделают его со всеми сими принадлежностями.
EXOD|25|40|Смотри, сделай их по тому образцу, какой показан тебе на горе.
EXOD|26|1|Скинию же сделай из десяти покрывал крученого виссона и из голубой, пурпуровой и червленой [шерсти], и херувимов сделай на них искусною работою;
EXOD|26|2|длина каждого покрывала двадцать восемь локтей, а ширина каждого покрывала четыре локтя: мера одна всем покрывалам.
EXOD|26|3|Пять покрывал пусть будут соединены одно с другим, и [другие] пять покрывал соединены одно с другим.
EXOD|26|4|Сделай петли голубого [цвета] на краю первого покрывала, в конце соединяющего обе половины; так сделай и на краю последнего покрывала, соединяющего обе половины;
EXOD|26|5|пятьдесят петлей сделай у одного покрывала и пятьдесят петлей сделай на краю покрывала, которое соединяется с другим; петли [должны] соответствовать одна другой;
EXOD|26|6|и сделай пятьдесят крючков золотых и крючками соедини покрывала одно с другим, и будет скиния одно [целое].
EXOD|26|7|И сделай покрывала на козьей [шерсти], чтобы покрывать скинию; одиннадцать покрывал сделай таких;
EXOD|26|8|длина одного покрывала тридцать локтей, а ширина четыре локтя; [это] одно покрывало: одиннадцати покрывалам одна мера.
EXOD|26|9|И соедини пять покрывал особо и шесть покрывал особо; шестое покрывало сделай двойное с передней стороны скинии.
EXOD|26|10|Сделай пятьдесят петлей на краю крайнего покрывала, для соединения его [с другим], и пятьдесят петлей на краю другого покрывала, для соединения с ним;
EXOD|26|11|сделай пятьдесят крючков медных, и вложи крючки в петли, и соедини покров, чтобы он составлял одно.
EXOD|26|12|А излишек, остающийся от покрывал скиний, – половина излишнего покрывала пусть будет свешена на задней стороне скинии;
EXOD|26|13|а излишек от длины покрывал скинии, на локоть с одной и на локоть с другой стороны, пусть будет свешен по бокам скинии с той и с другой стороны, для покрытия ее.
EXOD|26|14|И сделай покрышку для покрова из кож бараньих красных и еще покров верхний из кож синих.
EXOD|26|15|И сделай брусья для скинии из дерева ситтим, чтобы они стояли:
EXOD|26|16|длиною в десять локтей брус, и полтора локтя каждому брусу ширина;
EXOD|26|17|у каждого бруса по два шипа: один против другого: так сделай у всех брусьев скинии.
EXOD|26|18|Так сделай брусья для скинии: двадцать брусьев для полуденной стороны к югу,
EXOD|26|19|и под двадцать брусьев сделай сорок серебряных подножий: два подножия под один брус для двух шипов его, и два подножия под другой брус для двух шипов его;
EXOD|26|20|и двадцать брусьев для другой стороны скинии к северу,
EXOD|26|21|и для них сорок подножий серебряных: два подножия под один брус, и два подножия под другой брус.
EXOD|26|22|для задней же стороны скинии к западу сделай шесть брусьев
EXOD|26|23|и два бруса сделай для углов скинии на заднюю сторону;
EXOD|26|24|они должны быть соединены внизу и соединены вверху к одному кольцу: так должно быть с ними обоими; для обоих углов пусть они будут;
EXOD|26|25|и так будет восемь брусьев, и для них серебряных подножий шестнадцать: два подножия под один брус, и два подножия под другой брус.
EXOD|26|26|И сделай шесты из дерева ситтим, пять для брусьев одной стороны скинии,
EXOD|26|27|и пять шестов для брусьев другой стороны скинии, и пять шестов для брусьев задней стороны сзади скинии, к западу;
EXOD|26|28|а внутренний шест будет проходить по средине брусьев от одного конца до другого;
EXOD|26|29|брусья же обложи золотом, и кольца, для вкладывания шестов, сделай из золота, и шесты обложи золотом.
EXOD|26|30|И поставь скинию по образцу, который показан тебе на горе.
EXOD|26|31|И сделай завесу из голубой, пурпуровой и червленой шерсти и крученого виссона; искусною работою должны быть сделаны на ней херувимы;
EXOD|26|32|и повесь ее на четырех столбах из ситтим, обложенных золотом, с золотыми крючками, на четырех подножиях серебряных;
EXOD|26|33|и повесь завесу на крючках и внеси туда за завесу ковчег откровения; и будет завеса отделять вам святилище от Святаго–святых.
EXOD|26|34|И положи крышку на ковчег откровения во Святом–святых.
EXOD|26|35|И поставь стол вне завесы и светильник против стола на стороне скинии к югу; стол же поставь на северной стороне.
EXOD|26|36|И сделай завесу для входа в скинию из голубой и пурпуровой и червленой [шерсти] и из крученого виссона узорчатой работы;
EXOD|26|37|и сделай для завесы пять столбов из ситтим и обложи их золотом; крючки к ним золотые; и вылей для них пять подножий медных.
EXOD|27|1|И сделай жертвенник из дерева ситтим длиною пяти локтей и шириною пяти локтей, так чтобы он был четыреугольный, и вышиною трех локтей.
EXOD|27|2|И сделай роги на четырех углах его, так чтобы роги выходили из него; и обложи его медью.
EXOD|27|3|Сделай к нему горшки для высыпания в них пепла, и лопатки, и чаши, и вилки, и угольницы; все принадлежности сделай из меди.
EXOD|27|4|Сделай к нему решетку, род сетки, из меди, и сделай на сетке, на четырех углах ее, четыре кольца медных;
EXOD|27|5|и положи ее по окраине жертвенника внизу, так чтобы сетка была до половины жертвенника.
EXOD|27|6|И сделай шесты для жертвенника, шесты из дерева ситтим, и обложи их медью;
EXOD|27|7|и вкладывай шесты его в кольца, так чтобы шесты были по обоим бокам жертвенника, когда нести его.
EXOD|27|8|Сделай его пустой внутри, досчатый: как показано тебе на горе, так пусть сделают.
EXOD|27|9|Сделай двор скинии: с полуденной стороны к югу завесы для двора должны быть из крученого виссона, длиною во сто локтей по одной стороне;
EXOD|27|10|столбов для них двадцать, и подножий для них двадцать медных; крючки у столбов и связи на них из серебра.
EXOD|27|11|Также и вдоль по северной стороне – завесы ста локтей длиною; столбов для них двадцать, и подножий для них двадцать медных; крючки у столбов и связи на них из серебра.
EXOD|27|12|В ширину же двора с западной стороны – завесы пятидесяти локтей; столбов для них десять, и подножий к ним десять.
EXOD|27|13|И в ширину двора с передней стороны к востоку – [завесы] пятидесяти локтей.
EXOD|27|14|К одной стороне – завесы в пятнадцать локтей; столбов для них три, и подножий для них три;
EXOD|27|15|и к другой стороне – завесы в пятнадцать [локтей]; столбов для них три, и подножий для них три.
EXOD|27|16|А для ворот двора завеса в двадцать локтей из голубой и пурпуровой и червленой шерсти и из крученого виссона узорчатой работы; столбов для нее четыре, и подножий к ним четыре.
EXOD|27|17|Все столбы вокруг двора должны быть соединены связями из серебра; крючки у них из серебра, а подножия к ним из меди.
EXOD|27|18|Длина двора сто локтей, а ширина по всему протяжению пятьдесят, высота пять локтей; [завесы] из крученого виссона, а подножия [у] [столбов] из меди.
EXOD|27|19|Все принадлежности скинии для всякого употребления в ней, и все колья ее, и все колья двора – из меди.
EXOD|27|20|И вели сынам Израилевым, чтобы они приносили тебе елей чистый, выбитый из маслин, для освещения, чтобы горел светильник во всякое время;
EXOD|27|21|в скинии собрания вне завесы, которая пред [ковчегом] откровения, будет зажигать его Аарон и сыновья его, от вечера до утра, пред лицем Господним. [Это] устав вечный для поколений их от сынов Израилевых.
EXOD|28|1|И возьми к себе Аарона, брата твоего, и сынов его с ним, от среды сынов Израилевых, чтоб он был священником Мне, Аарона и Надава, Авиуда, Елеазара и Ифамара, сынов Аароновых.
EXOD|28|2|И сделай священные одежды Аарону, брату твоему, для славы и благолепия.
EXOD|28|3|И скажи всем мудрым сердцем, которых Я исполнил духа премудрости, чтобы они сделали Аарону одежды для посвящения его, чтобы он был священником Мне.
EXOD|28|4|Вот одежды, которые должны они сделать: наперсник, ефод, верхняя риза, хитон стяжной, кидар и пояс. Пусть сделают священные одежды Аарону, брату твоему, и сынам его, чтобы он был священником Мне.
EXOD|28|5|Пусть они возьмут золота, голубой и пурпуровой и червленой шерсти и виссона,
EXOD|28|6|и сделают ефод из золота, из голубой, пурпуровой и червленой [шерсти], и из крученого виссона, искусною работою.
EXOD|28|7|У него должны быть на обоих концах его два связывающие нарамника, чтобы он был связан.
EXOD|28|8|И пояс ефода, который поверх его, должен быть одинаковой с ним работы, из золота, из голубой, пурпуровой и червленой [шерсти] и из крученого виссона.
EXOD|28|9|И возьми два камня оникса и вырежь на них имена сынов Израилевых:
EXOD|28|10|шесть имен их на одном камне и шесть имен остальных на другом камне, по [порядку] рождения их;
EXOD|28|11|чрез резчика на камне, который вырезывает печати, вырежь на двух камнях имена сынов Израилевых; и вставь их в золотые гнезда
EXOD|28|12|и положи два камня сии на нарамники ефода: [это] камни на память сынам Израилевым; и будет Аарон носить имена их пред Господом на обоих раменах своих для памяти.
EXOD|28|13|И сделай гнезда из золота;
EXOD|28|14|и две цепочки из чистого золота, витыми сделай их работою плетеною, и прикрепи витые цепочки к гнездам.
EXOD|28|15|Сделай наперсник судный искусною работою; сделай его такою же работою, как ефод: из золота, из голубой, пурпуровой и червленой [шерсти] и из крученого виссона сделай его;
EXOD|28|16|он должен быть четыреугольный, двойной, в пядень длиною и в пядень шириною;
EXOD|28|17|и вставь в него оправленные камни в четыре ряда; рядом: рубин, топаз, изумруд, – это один ряд;
EXOD|28|18|второй ряд: карбункул, сапфир и алмаз;
EXOD|28|19|третий ряд: яхонт, агат и аметист;
EXOD|28|20|четвертый ряд: хризолит, оникс и яспис; в золотых гнездах должны быть вставлены они.
EXOD|28|21|Сих камней должно быть двенадцать, по [числу сынов Израилевых], по именам их; на каждом, как на печати, должно быть вырезано по одному имени из числа двенадцати колен.
EXOD|28|22|К наперснику сделай цепочки витые плетеною работою из чистого золота;
EXOD|28|23|и сделай к наперснику два кольца из золота и прикрепи два кольца к двум концам наперсника;
EXOD|28|24|и вдень две плетеные цепочки из золота в оба кольца по концам наперсника,
EXOD|28|25|а два конца двух цепочек прикрепи к двум гнездам и прикрепи к нарамникам ефода с лицевой стороны его;
EXOD|28|26|еще сделай два кольца золотых и прикрепи их к двум [другим] концам наперсника, на той стороне, которая лежит к ефоду внутрь;
EXOD|28|27|также сделай два кольца золотых и прикрепи их к двум нарамникам ефода снизу, с лицевой стороны его, у соединения его, над поясом ефода;
EXOD|28|28|и прикрепят наперсник кольцами его к кольцам ефода шнуром из голубой шерсти, чтобы он был над поясом ефода, и чтоб не спадал наперсник с ефода.
EXOD|28|29|И будет носить Аарон имена сынов Израилевых на наперснике судном у сердца своего, когда будет входить во святилище, для постоянной памяти пред Господом.
EXOD|28|30|На наперсник судный возложи урим и туммим, и они будут у сердца Ааронова, когда будет он входить [во святилище] пред лице Господне; и будет Аарон всегда носить суд сынов Израилевых у сердца своего пред лицем Господним.
EXOD|28|31|И сделай верхнюю ризу к ефоду всю голубого [цвета];
EXOD|28|32|среди ее должно быть отверстие для головы; у отверстия ее вокруг должна быть обшивка тканая, подобно как у отверстия брони, чтобы не дралось;
EXOD|28|33|по подолу ее сделай яблоки из [нитей] голубого, яхонтового, пурпурового и червленого [цвета], вокруг по подолу ее; позвонки золотые между ними кругом:
EXOD|28|34|золотой позвонок и яблоко, золотой позвонок и яблоко, по подолу верхней ризы кругом;
EXOD|28|35|она будет на Аароне в служении, дабы слышен был от него звук, когда он будет входить во святилище пред лице Господне и когда будет выходить, чтобы ему не умереть.
EXOD|28|36|И сделай полированную дощечку из чистого золота, и вырежь на ней, как вырезывают на печати: "Святыня Господня",
EXOD|28|37|и прикрепи ее шнуром голубого цвета к кидару, так чтобы она была на передней стороне кидара;
EXOD|28|38|и будет она на челе Аароновом, и понесет на себе Аарон недостатки приношений, посвящаемых от сынов Израилевых, и всех даров, ими приносимых; и будет она непрестанно на челе его, для благоволения Господня к ним.
EXOD|28|39|И сделай хитон из виссона и кидар из виссона и сделай пояс узорчатой работы;
EXOD|28|40|сделай и сынам Аароновым хитоны, сделай им поясы, и головные повязки сделай им для славы и благолепия,
EXOD|28|41|и облеки в них Аарона, брата твоего, и сынов его с ним, и помажь их, и наполни руки их, и посвяти их, и они будут священниками Мне.
EXOD|28|42|И сделай им нижнее платье льняное, для прикрытия телесной наготы от чресл до голеней,
EXOD|28|43|и да будут они на Аароне и на сынах его, когда будут они входить в скинию собрания, или приступать к жертвеннику для служения во святилище, чтобы им не навести [на себя] греха и не умереть. [Это] устав вечный для него и для потомков его по нем.
EXOD|29|1|Вот что должен ты совершить над ними, чтобы посвятить их во священники Мне: возьми одного тельца из волов, и двух овнов без порока,
EXOD|29|2|и хлебов пресных, и опресноков, смешанных с елеем, и лепешек пресных, помазанных елеем: из муки пшеничной сделай их,
EXOD|29|3|и положи их в одну корзину, и принеси их в корзине, и вместе тельца и двух овнов.
EXOD|29|4|Аарона же и сынов его приведи ко входу в скинию собрания и омой их водою.
EXOD|29|5|И возьми одежды, и облеки Аарона в хитон и в верхнюю ризу, в ефод и в наперсник, и опояшь его по ефоду;
EXOD|29|6|и возложи ему на голову кидар и укрепи диадиму святыни на кидаре;
EXOD|29|7|и возьми елей помазания, и возлей ему на голову, и помажь его.
EXOD|29|8|И приведи также сынов его и облеки их в хитоны;
EXOD|29|9|и опояшь их поясом, Аарона и сынов его, и возложи на них повязки и будет им принадлежать священство по уставу на веки; и наполни руки Аарона и сынов его.
EXOD|29|10|И приведи тельца пред скинию собрания, и возложат Аарон и сыны его руки свои на голову тельца,
EXOD|29|11|и заколи тельца пред лицем Господним при входе в скинию собрания;
EXOD|29|12|возьми крови тельца и возложи перстом твоим на роги жертвенника, а всю кровь вылей у основания жертвенника;
EXOD|29|13|возьми весь тук, покрывающий внутренности, и сальник с печени, и обе почки и тук, который на них, и воскури на жертвеннике;
EXOD|29|14|а мясо тельца и кожу его и нечистоты его сожги на огне вне стана: это – [жертва] за грех.
EXOD|29|15|И возьми одного овна, и возложат Аарон и сыны его руки свои на голову овна;
EXOD|29|16|и заколи овна, и возьми крови его, и покропи на жертвенник со всех сторон;
EXOD|29|17|рассеки овна на части, вымой внутренности его и голени его, и положи [их] на рассеченные части его и на голову его;
EXOD|29|18|и сожги всего овна на жертвеннике. Это всесожжение Господу, благоухание приятное, жертва Господу.
EXOD|29|19|Возьми и другого овна, и возложат Аарон и сыны его руки свои на голову овна;
EXOD|29|20|и заколи овна, и возьми крови его, и возложи на край правого уха Ааронова и на край правого уха сынов его, и на большой палец правой руки их, и на большой палец правой ноги их; и покропи кровью на жертвенник со всех сторон;
EXOD|29|21|и возьми крови, которая на жертвеннике, и елея помазания, и покропи на Аарона и на одежды его, и на сынов его, и на одежды сынов его с ним, – и будут освящены, он и одежды его, и сыны его и одежды их с ним.
EXOD|29|22|И возьми от овна тук и курдюк, и тук, покрывающий внутренности, и сальник с печени, и обе почки и тук, который на них, правое плечо,
EXOD|29|23|и один круглый хлеб, одну лепешку на елее и один опреснок из корзины, которая пред Господом,
EXOD|29|24|и положи все на руки Аарону и на руки сынам его, и принеси это, потрясая пред лицем Господним;
EXOD|29|25|и возьми это с рук их и сожги на жертвеннике со всесожжением, в благоухание пред Господом: это жертва Господу.
EXOD|29|26|И возьми грудь от овна вручения, который для Аарона, и принеси ее, потрясая пред лицем Господним, – и это будет твоя доля;
EXOD|29|27|и освяти грудь приношения, которая потрясаема была и плечо возношения, которое было возносимо, от овна вручения, который для Аарона и для сынов его, –
EXOD|29|28|и будет [это] Аарону и сынам его в участок вечный от сынов Израилевых, ибо это – возношение; возношение должно быть от сынов Израилевых при мирных жертвах, возношение их Господу.
EXOD|29|29|А священные одежды, которые для Аарона, перейдут после него к сынам его, чтобы в них помазывать их и вручать им [священство];
EXOD|29|30|семь дней должен облачаться в них священник из сынов его, заступающий его место, который будет входить в скинию собрания для служения во святилище.
EXOD|29|31|Овна же вручения возьми и свари мясо его на месте святом;
EXOD|29|32|и пусть съедят Аарон и сыны его мясо овна сего из корзины, у дверей скинии собрания,
EXOD|29|33|ибо чрез это совершено очищение для вручения им священства и для посвящения их; посторонний не должен есть [сего], ибо это святыня;
EXOD|29|34|если останется от мяса вручения и от хлеба до утра, то сожги остаток на огне: не должно есть его, ибо это святыня.
EXOD|29|35|И поступи с Аароном и с сынами его во всем так, как Я повелел тебе; в семь дней наполняй руки их.
EXOD|29|36|И тельца за грех приноси каждый день для очищения, и жертву за грех совершай на жертвеннике для очищения его, и помажь его для освящения его;
EXOD|29|37|семь дней очищай жертвенник, и освяти его, и будет жертвенник святыня великая: все, прикасающееся к жертвеннику, освятится.
EXOD|29|38|Вот что будешь ты приносить на жертвеннике: двух агнцев однолетних каждый день постоянно.
EXOD|29|39|одного агнца приноси поутру, а другого агнца приноси вечером,
EXOD|29|40|и десятую [часть ефы] пшеничной муки, смешанной с четвертью гина битого елея, а для возлияния четверть гина вина, для одного агнца;
EXOD|29|41|другого агнца приноси вечером: с мучным даром, подобным утреннему, и с таким же возлиянием приноси его в благоухание приятное, в жертву Господу.
EXOD|29|42|Это – всесожжение постоянное в роды ваши пред дверями скинии собрания пред Господом, где буду открываться вам, чтобы говорить с тобою;
EXOD|29|43|там буду открываться сынам Израилевым, и освятится [место сие] славою Моею.
EXOD|29|44|И освящу скинию собрания и жертвенник; и Аарона и сынов его освящу, чтобы они священнодействовали Мне;
EXOD|29|45|и буду обитать среди сынов Израилевых, и буду им Богом,
EXOD|29|46|и узнают, что Я Господь, Бог их, Который вывел их из земли Египетской, чтобы Мне обитать среди них. Я Господь, Бог их.
EXOD|30|1|И сделай жертвенник для приношения курений, из дерева ситтим сделай его:
EXOD|30|2|длина ему локоть, и ширина ему локоть; он должен быть четыреугольный; а вышина ему два локтя; из него [должны выходить] роги его;
EXOD|30|3|обложи его чистым золотом, верх его и бока его кругом, и роги его; и сделай к нему золотой венец вокруг;
EXOD|30|4|под венцом его на двух углах его сделай два кольца из золота; сделай их с двух сторон его; и будут они влагалищем для шестов, чтобы носить его на них;
EXOD|30|5|шесты сделай из дерева ситтим и обложи их золотом.
EXOD|30|6|И поставь его пред завесою, которая пред ковчегом откровения, против крышки, которая на [ковчеге] откровения, где Я буду открываться тебе.
EXOD|30|7|На нем Аарон будет курить благовонным курением; каждое утро, когда он приготовляет лампады, будет курить им;
EXOD|30|8|и когда Аарон зажигает лампады вечером, он будет курить им: [это] – всегдашнее курение пред Господом в роды ваши.
EXOD|30|9|Не приносите на нем никакого иного курения, ни всесожжения, ни приношения хлебного, и возлияния не возливайте на него.
EXOD|30|10|И будет совершать Аарон очищение над рогами его однажды в год; кровью очистительной [жертвы] за грех он будет очищать его однажды в год в роды ваши. Это святыня великая у Господа.
EXOD|30|11|И сказал Господь Моисею, говоря:
EXOD|30|12|когда будешь делать исчисление сынов Израилевых при пересмотре их, то пусть каждый даст выкуп за душу свою Господу при исчислении их, и не будет между ними язвы губительной при исчислении их;
EXOD|30|13|всякий, поступающий в исчисление, должен давать половину сикля, сикля священного; в сикле двадцать гер: полсикля приношение Господу;
EXOD|30|14|всякий, поступающий в исчисление от двадцати лет и выше, должен давать приношение Господу;
EXOD|30|15|богатый не больше и бедный не меньше полсикля должны давать в приношение Господу, для выкупа душ ваших;
EXOD|30|16|и возьми серебро выкупа от сынов Израилевых и употребляй его на служение скинии собрания; и будет это для сынов Израилевых в память пред Господом, для искупления душ ваших.
EXOD|30|17|И сказал Господь Моисею, говоря:
EXOD|30|18|сделай умывальник медный для омовения и подножие его медное, и поставь его между скиниею собрания и между жертвенником, и налей в него воды;
EXOD|30|19|и пусть Аарон и сыны его омывают из него руки свои и ноги свои;
EXOD|30|20|когда они должны входить в скинию собрания, пусть они омываются водою, чтобы им не умереть; или когда должны приступать к жертвеннику для служения, для жертвоприношения Господу,
EXOD|30|21|пусть они омывают руки свои и ноги свои водою, чтобы им не умереть; и будет им это уставом вечным, ему и потомкам его в роды их.
EXOD|30|22|И сказал Господь Моисею, говоря:
EXOD|30|23|возьми себе самых лучших благовонных веществ: смирны самоточной пятьсот [сиклей], корицы благовонной половину против того, двести пятьдесят, тростника благовонного двести пятьдесят,
EXOD|30|24|касии пятьсот [сиклей], по сиклю священному, и масла оливкового гин;
EXOD|30|25|и сделай из сего миро для священного помазания, масть составную, искусством составляющего масти: это будет миро для священного помазания;
EXOD|30|26|и помажь им скинию собрания и ковчег откровения,
EXOD|30|27|и стол и все принадлежности его, и светильник и все принадлежности его, и жертвенник курения,
EXOD|30|28|и жертвенник всесожжения и все принадлежности его, и умывальник и подножие его;
EXOD|30|29|и освяти их, и будет святыня великая: все, прикасающееся к ним, освятится;
EXOD|30|30|помажь и Аарона и сынов его и посвяти их, чтобы они были священниками Мне.
EXOD|30|31|А сынам Израилевым скажи: это будет у Меня миро священного помазания в роды ваши;
EXOD|30|32|тела прочих людей не должно помазывать им, и по составу его не делайте подобного ему; оно – святыня: святынею должно быть для вас;
EXOD|30|33|кто составит подобное ему или кто помажет им постороннего, тот истребится из народа своего.
EXOD|30|34|И сказал Господь Моисею: возьми себе благовонных веществ: стакти, ониха, халвана душистого и чистого ливана, всего половину,
EXOD|30|35|и сделай из них искусством составляющего масти курительный состав, стертый, чистый, святый,
EXOD|30|36|и истолки его мелко, и полагай его пред [ковчегом] откровения в скинии собрания, где Я буду открываться тебе: это будет святыня великая для вас;
EXOD|30|37|курения, сделанного по сему составу, не делайте себе: святынею да будет оно у тебя для Господа;
EXOD|30|38|кто сделает подобное, чтобы курить им, истребится из народа своего.
EXOD|31|1|И сказал Господь Моисею, говоря:
EXOD|31|2|смотри, Я назначаю именно Веселеила, сына Уриева, сына Орова, из колена Иудина;
EXOD|31|3|и Я исполнил его Духом Божиим, мудростью, разумением, ведением и всяким искусством,
EXOD|31|4|работать из золота, серебра и меди,
EXOD|31|5|резать камни для вставливания и резать дерево для всякого дела;
EXOD|31|6|и вот, Я даю ему помощником Аголиава, сына Ахисамахова, из колена Данова, и в сердце всякого мудрого вложу мудрость, дабы они сделали все, что Я повелел тебе:
EXOD|31|7|скинию собрания и ковчег откровения и крышку на него, и все принадлежности скинии,
EXOD|31|8|и стол и принадлежности его, и светильник из чистого золота и все принадлежности его, и жертвенник курения,
EXOD|31|9|и жертвенник всесожжения и все принадлежности его, и умывальник и подножие его,
EXOD|31|10|и одежды служебные и одежды священные Аарону священнику, и одежды сынам его, для священнослужения,
EXOD|31|11|и елей помазания и курение благовонное для святилища: все так, как Я повелел тебе, они сделают.
EXOD|31|12|И сказал Господь Моисею, говоря:
EXOD|31|13|скажи сынам Израилевым так: субботы Мои соблюдайте, ибо это – знамение между Мною и вами в роды ваши, дабы вы знали, что Я Господь, освящающий вас;
EXOD|31|14|и соблюдайте субботу, ибо она свята для вас: кто осквернит ее, тот да будет предан смерти; кто станет в оную делать дело, та душа должна быть истреблена из среды народа своего;
EXOD|31|15|шесть дней пусть делают дела, а в седьмой – суббота покоя, посвященная Господу: всякий, кто делает дело в день субботний, да будет предан смерти;
EXOD|31|16|и пусть хранят сыны Израилевы субботу, празднуя субботу в роды свои, как завет вечный;
EXOD|31|17|это – знамение между Мною и сынами Израилевыми на веки, потому что в шесть дней сотворил Господь небо и землю, а в день седьмой почил и покоился.
EXOD|31|18|И когда [Бог] перестал говорить с Моисеем на горе Синае, дал ему две скрижали откровения, скрижали каменные, на которых написано было перстом Божиим.
EXOD|32|1|Когда народ увидел, что Моисей долго не сходит с горы, то собрался к Аарону и сказал ему: встань и сделай нам бога, который бы шел перед нами, ибо с этим человеком, с Моисеем, который вывел нас из земли Египетской, не знаем, что сделалось.
EXOD|32|2|И сказал им Аарон: выньте золотые серьги, которые в ушах ваших жен, ваших сыновей и ваших дочерей, и принесите ко мне.
EXOD|32|3|И весь народ вынул золотые серьги из ушей своих и принесли к Аарону.
EXOD|32|4|Он взял их из рук их, и сделал из них литого тельца, и обделал его резцом. И сказали они: вот бог твой, Израиль, который вывел тебя из земли Египетской!
EXOD|32|5|Увидев [сие], Аарон поставил пред ним жертвенник, и провозгласил Аарон, говоря: завтра праздник Господу.
EXOD|32|6|На другой день они встали рано и принесли всесожжения и привели жертвы мирные: и сел народ есть и пить, а после встал играть.
EXOD|32|7|И сказал Господь Моисею: поспеши сойти; ибо развратился народ твой, который ты вывел из земли Египетской;
EXOD|32|8|скоро уклонились они от пути, который Я заповедал им: сделали себе литого тельца и поклонились ему, и принесли ему жертвы и сказали: вот бог твой, Израиль, который вывел тебя из земли Египетской!
EXOD|32|9|И сказал Господь Моисею: Я вижу народ сей, и вот, народ он – жестоковыйный;
EXOD|32|10|итак оставь Меня, да воспламенится гнев Мой на них, и истреблю их, и произведу многочисленный народ от тебя.
EXOD|32|11|Но Моисей стал умолять Господа, Бога Своего, и сказал: да не воспламеняется, Господи, гнев Твой на народ Твой, который Ты вывел из земли Египетской силою великою и рукою крепкою,
EXOD|32|12|чтобы Египтяне не говорили: на погибель Он вывел их, чтобы убить их в горах и истребить их с лица земли; отврати пламенный гнев Твой и отмени погубление народа Твоего;
EXOD|32|13|вспомни Авраама, Исаака и Израиля, рабов Твоих, которым клялся Ты Собою, говоря: умножая умножу семя ваше, как звезды небесные, и всю землю сию, о которой Я сказал, дам семени вашему, и будут владеть вечно.
EXOD|32|14|И отменил Господь зло, о котором сказал, что наведет его на народ Свой.
EXOD|32|15|И обратился и сошел Моисей с горы; в руке его [были] две скрижали откровения, на которых написано было с обеих сторон: и на той и на другой стороне написано было;
EXOD|32|16|скрижали были дело Божие, и письмена, начертанные на скрижалях, были письмена Божии.
EXOD|32|17|И услышал Иисус голос народа шумящего и сказал Моисею: военный крик в стане.
EXOD|32|18|Но [Моисей] сказал: это не крик побеждающих и не вопль поражаемых; я слышу голос поющих.
EXOD|32|19|Когда же он приблизился к стану и увидел тельца и пляски, тогда он воспламенился гневом и бросил из рук своих скрижали и разбил их под горою;
EXOD|32|20|и взял тельца, которого они сделали, и сжег его в огне, и стер в прах, и рассыпал по воде, и дал ее пить сынам Израилевым.
EXOD|32|21|И сказал Моисей Аарону: что сделал тебе народ сей, что ты ввел его в грех великий?
EXOD|32|22|Но Аарон сказал: да не возгорается гнев господина моего; ты знаешь этот народ, что он буйный.
EXOD|32|23|Они сказали мне: сделай нам бога, который шел бы перед нами; ибо с Моисеем, с этим человеком, который вывел нас из земли Египетской, не знаем, что сделалось.
EXOD|32|24|И я сказал им: у кого есть золото, снимите с себя. и отдали мне; я бросил его в огонь, и вышел этот телец.
EXOD|32|25|Моисей увидел, что это народ необузданный, ибо Аарон допустил его до необузданности, к посрамлению пред врагами его.
EXOD|32|26|И стал Моисей в воротах стана и сказал: кто Господень, – ко мне! И собрались к нему все сыны Левиины.
EXOD|32|27|И он сказал им: так говорит Господь Бог Израилев: возложите каждый свой меч на бедро свое, пройдите по стану от ворот до ворот и обратно, и убивайте каждый брата своего, каждый друга своего, каждый ближнего своего.
EXOD|32|28|И сделали сыны Левиины по слову Моисея: и пало в тот день из народа около трех тысяч человек.
EXOD|32|29|Ибо Моисей сказал: сегодня посвятите руки ваши Господу, каждый в сыне своем и брате своем, да ниспошлет Он вам сегодня благословение.
EXOD|32|30|На другой день сказал Моисей народу: вы сделали великий грех; итак я взойду к Господу, не заглажу ли греха вашего.
EXOD|32|31|И возвратился Моисей к Господу и сказал: о, народ сей сделал великий грех: сделал себе золотого бога;
EXOD|32|32|прости им грех их, а если нет, то изгладь и меня из книги Твоей, в которую Ты вписал.
EXOD|32|33|Господь сказал Моисею: того, кто согрешил предо Мною, изглажу из книги Моей;
EXOD|32|34|итак, иди, веди народ сей, куда Я сказал тебе; вот Ангел Мой пойдет пред тобою, и в день посещения Моего Я посещу их за грех их.
EXOD|32|35|И поразил Господь народ за сделанного тельца, которого сделал Аарон.
EXOD|33|1|И сказал Господь Моисею: пойди, иди отсюда ты и народ, который ты вывел из земли Египетской, в землю, о которой Я клялся Аврааму, Исааку и Иакову, говоря: потомству твоему дам ее;
EXOD|33|2|и пошлю пред тобою Ангела, и прогоню Хананеев, Аморреев, Хеттеев, Ферезеев, Евеев и Иевусеев,
EXOD|33|3|[и введет он вас] в землю, где течет молоко и мед; ибо Сам не пойду среди вас, чтобы не погубить Мне вас на пути, потому что вы народ жестоковыйный.
EXOD|33|4|Народ, услышав грозное слово сие, возрыдал, и никто не возложил на себя украшений своих.
EXOD|33|5|Ибо Господь сказал Моисею: скажи сынам Израилевым: вы народ жестоковыйный; если Я пойду среди вас, то в одну минуту истреблю вас; итак снимите с себя украшения свои; Я посмотрю, что Мне делать с вами.
EXOD|33|6|Сыны Израилевы сняли с себя украшения свои у горы Хорива.
EXOD|33|7|Моисей же взял и поставил себе шатер вне стана, вдали от стана, и назвал его скиниею собрания; и каждый, ищущий Господа, приходил в скинию собрания, находившуюся вне стана.
EXOD|33|8|И когда Моисей выходил к скинии, весь народ вставал, и становился каждый у входа в свой шатер и смотрел вслед Моисею, доколе он не входил в скинию.
EXOD|33|9|Когда же Моисей входил в скинию, тогда спускался столп облачный и становился у входа в скинию, и [Господь] говорил с Моисеем.
EXOD|33|10|И видел весь народ столп облачный, стоявший у входа в скинию; и вставал весь народ, и поклонялся каждый у входа в шатер свой.
EXOD|33|11|И говорил Господь с Моисеем лицем к лицу, как бы говорил кто с другом своим; и он возвращался в стан; а служитель его Иисус, сын Навин, юноша, не отлучался от скинии.
EXOD|33|12|Моисей сказал Господу: вот, Ты говоришь мне: веди народ сей, а не открыл мне, кого пошлешь со мною, хотя Ты сказал: "Я знаю тебя по имени, и ты приобрел благоволение в очах Моих";
EXOD|33|13|итак, если я приобрел благоволение в очах Твоих, то молю: открой мне путь Твой, дабы я познал Тебя, чтобы приобрести благоволение в очах Твоих; и помысли, что сии люди Твой народ.
EXOD|33|14|[Господь] сказал: Сам Я пойду, и введу тебя в покой.
EXOD|33|15|[Моисей] сказал Ему: если не пойдешь Ты Сам [с нами], то и не выводи нас отсюда,
EXOD|33|16|ибо по чему узнать, что я и народ Твой обрели благоволение в очах Твоих? не по тому ли, когда Ты пойдешь с нами? тогда я и народ Твой будем славнее всякого народа на земле.
EXOD|33|17|И сказал Господь Моисею: и то, о чем ты говорил, Я сделаю, потому что ты приобрел благоволение в очах Моих, и Я знаю тебя по имени.
EXOD|33|18|[Моисей] сказал: покажи мне славу Твою.
EXOD|33|19|И сказал [Господь]: Я проведу пред тобою всю славу Мою и провозглашу имя Иеговы пред тобою, и кого помиловать – помилую, кого пожалеть – пожалею.
EXOD|33|20|И потом сказал Он: лица Моего не можно тебе увидеть, потому что человек не может увидеть Меня и остаться в живых.
EXOD|33|21|И сказал Господь: вот место у Меня, стань на этой скале;
EXOD|33|22|когда же будет проходить слава Моя, Я поставлю тебя в расселине скалы и покрою тебя рукою Моею, доколе не пройду;
EXOD|33|23|и когда сниму руку Мою, ты увидишь Меня сзади, а лице Мое не будет видимо.
EXOD|34|1|И сказал Господь Моисею: вытеши себе две скрижали каменные, подобные прежним, и Я напишу на сих скрижалях слова, какие были на прежних скрижалях, которые ты разбил;
EXOD|34|2|и будь готов к утру, и взойди утром на гору Синай, и предстань предо Мною там на вершине горы;
EXOD|34|3|но никто не должен восходить с тобою, и никто не должен показываться на всей горе; даже скот, мелкий и крупный, не должен пастись близ горы сей.
EXOD|34|4|И вытесал Моисей две скрижали каменные, подобные прежним, и, встав рано поутру, взошел на гору Синай, как повелел ему Господь; и взял в руки свои две скрижали каменные.
EXOD|34|5|И сошел Господь в облаке, и остановился там близ него, и провозгласил имя Иеговы.
EXOD|34|6|И прошел Господь пред лицем его и возгласил: Господь, Господь, Бог человеколюбивый и милосердый, долготерпеливый и многомилостивый и истинный,
EXOD|34|7|сохраняющий милость в тысячи [родов], прощающий вину и преступление и грех, но не оставляющий без наказания, наказывающий вину отцов в детях и в детях детей до третьего и четвертого рода.
EXOD|34|8|Моисей тотчас пал на землю и поклонился [Богу]
EXOD|34|9|и сказал: если я приобрел благоволение в очах Твоих, Владыка, то да пойдет Владыка посреди нас; ибо народ сей жестоковыен; прости беззакония наши и грехи наши и сделай нас наследием Твоим.
EXOD|34|10|И сказал [Господь]: вот, Я заключаю завет: пред всем народом твоим соделаю чудеса, каких не было по всей земле и ни у каких народов; и увидит весь народ, среди которого ты находишься, дело Господа; ибо страшно будет то, что Я сделаю для тебя;
EXOD|34|11|сохрани то, что повелеваю тебе ныне: вот, Я изгоняю от лица твоего Аморреев, Хананеев, Хеттеев, Ферезеев, Евеев, и Иевусеев;
EXOD|34|12|смотри, не вступай в союз с жителями той земли, в которую ты войдешь, дабы они не сделались сетью среди вас.
EXOD|34|13|Жертвенники их разрушьте, столбы их сокрушите, вырубите [священные] рощи их.
EXOD|34|14|ибо ты не должен поклоняться богу иному, кроме Господа; потому что имя Его – ревнитель; Он Бог ревнитель.
EXOD|34|15|Не вступай в союз с жителями той земли, чтобы, когда они будут блудодействовать вслед богов своих и приносить жертвы богам своим, не пригласили и тебя, и ты не вкусил бы жертвы их;
EXOD|34|16|и не бери из дочерей их жен сынам своим, дабы дочери их, блудодействуя вслед богов своих, не ввели и сынов твоих в блужение вслед богов своих.
EXOD|34|17|Не делай себе богов литых.
EXOD|34|18|Праздник опресноков соблюдай: семь дней ешь пресный хлеб, как Я повелел тебе, в назначенное время месяца Авива, ибо в месяце Авиве вышел ты из Египта.
EXOD|34|19|Все, разверзающее ложесна – Мне, как и весь скот твой мужеского пола, разверзающий ложесна, из волов и овец;
EXOD|34|20|первородное из ослов заменяй агнцем, а если не заменишь, то выкупи его; всех первенцев из сынов твоих выкупай; пусть не являются пред лице Мое с пустыми руками.
EXOD|34|21|Шесть дней работай, а в седьмой день покойся; покойся и во время посева и жатвы.
EXOD|34|22|И праздник седмиц совершай, праздник начатков жатвы пшеницы и праздник собирания [плодов] в конце года;
EXOD|34|23|три раза в году должен являться весь мужеский пол твой пред лице Владыки, Господа Бога Израилева,
EXOD|34|24|ибо Я прогоню народы от лица твоего и распространю пределы твои, и никто не пожелает земли твоей, если ты будешь являться пред лице Господа Бога твоего три раза в году.
EXOD|34|25|Не изливай крови жертвы Моей на квасное, и жертва праздника Пасхи не должна переночевать до утра.
EXOD|34|26|Самые первые плоды земли твоей принеси в дом Господа Бога твоего. Не вари козленка в молоке матери его.
EXOD|34|27|И сказал Господь Моисею: напиши себе слова сии, ибо в сих словах Я заключаю завет с тобою и с Израилем.
EXOD|34|28|И пробыл там [Моисей] у Господа сорок дней и сорок ночей, хлеба не ел и воды не пил; и написал на скрижалях слова завета, десятословие.
EXOD|34|29|Когда сходил Моисей с горы Синая, и две скрижали откровения были в руке у Моисея при сошествии его с горы, то Моисей не знал, что лице его стало сиять лучами от того, что [Бог] говорил с ним.
EXOD|34|30|И увидел Моисея Аарон и все сыны Израилевы, и вот, лице его сияет, и боялись подойти к нему.
EXOD|34|31|И призвал их Моисей, и пришли к нему Аарон и все начальники общества, и разговаривал Моисей с ними.
EXOD|34|32|После сего приблизились все сыны Израилевы, и он заповедал им все, что говорил ему Господь на горе Синае.
EXOD|34|33|И когда Моисей перестал разговаривать с ними, то положил на лице свое покрывало.
EXOD|34|34|Когда же входил Моисей пред лице Господа, чтобы говорить с Ним, тогда снимал покрывало, доколе не выходил; а выйдя пересказывал сынам Израилевым все, что заповедано было.
EXOD|34|35|И видели сыны Израилевы, что сияет лице Моисеево, и Моисей опять полагал покрывало на лице свое, доколе не входил говорить с Ним.
EXOD|35|1|И собрал Моисей все общество сынов Израилевых и сказал им: вот что заповедал Господь делать:
EXOD|35|2|шесть дней делайте дела, а день седьмой должен быть у вас святым, суббота покоя Господу: всякий, кто будет делать в нее дело, предан будет смерти;
EXOD|35|3|не зажигайте огня во всех жилищах ваших в день субботы.
EXOD|35|4|И сказал Моисей всему обществу сынов Израилевых: вот что заповедал Господь:
EXOD|35|5|сделайте от себя приношения Господу: каждый по усердию пусть принесет приношение Господу, золото, серебро, медь,
EXOD|35|6|[шерсть] голубого, пурпурового и червленого [цвета], и виссон, и козью шерсть,
EXOD|35|7|кожи бараньи красные, и кожи синие, и дерево ситтим,
EXOD|35|8|и елей для светильника, и ароматы для елея помазания и для благовонных курений,
EXOD|35|9|камень оникс и камни вставные для ефода и наперсника.
EXOD|35|10|И всякий из вас мудрый сердцем пусть придет и сделает все, что повелел Господь:
EXOD|35|11|скинию и покров ее и [верхнюю] покрышку ее, крючки и брусья ее, шесты ее, столбы ее и подножия ее,
EXOD|35|12|ковчег и шесты его, крышку и завесу для преграды,
EXOD|35|13|стол и шесты его и все принадлежности его, и хлебы предложения,
EXOD|35|14|и светильник для освещения с принадлежностями его, и лампады его и елей для освещения,
EXOD|35|15|и жертвенник для курений и шесты его, и елей помазания, и благовонные курения, и завесу ко входу скинии,
EXOD|35|16|жертвенник всесожжения и решетку медную для него, и шесты его и все принадлежности его, умывальник и подножие его,
EXOD|35|17|завесы двора, столбы его и подножия их, и завесу у входа во двор,
EXOD|35|18|колья скинии, и колья двора и веревки их,
EXOD|35|19|одежды служебные для служения во святилище, и священные одежды Аарону священнику и одежды сынам его для священнодействия.
EXOD|35|20|И пошло все общество сынов Израилевых от Моисея.
EXOD|35|21|И приходили все, которых влекло к тому сердце, и все, которых располагал дух, и приносили приношения Господу для устроения скинии собрания и для всех потребностей ее и для священных одежд;
EXOD|35|22|и приходили мужья с женами, и все по расположению сердца приносили кольца, серьги, перстни и привески, всякие золотые вещи, каждый, кто только хотел приносить золото Господу;
EXOD|35|23|и каждый, у кого была [шерсть] голубого, пурпурового и червленого [цвета], виссон и козья шерсть, кожи бараньи красные и кожи синие, приносил их;
EXOD|35|24|и каждый, кто жертвовал серебро или медь, приносил сие в дар Господу; и каждый, у кого было дерево ситтим, приносил сие на всякую потребность [для скинии];
EXOD|35|25|и все женщины, мудрые сердцем, пряли своими руками и приносили пряжу голубого, пурпурового и червленого [цвета] и виссон;
EXOD|35|26|и все женщины, которых влекло сердце, умевшие прясть, пряли козью шерсть;
EXOD|35|27|князья же приносили камень оникс и камни вставные для ефода и наперсника,
EXOD|35|28|также и благовония, и елей для светильника и для [составления] елея помазания и для благовонных курений;
EXOD|35|29|и все мужья и жены из сынов Израилевых, которых влекло сердце принести на всякое дело, какое Господь чрез Моисея повелел сделать, приносили добровольный дар Господу.
EXOD|35|30|И сказал Моисей сынам Израилевым: смотрите, Господь назначил именно Веселеила, сына Урии, сына Ора, из колена Иудина,
EXOD|35|31|и исполнил его Духом Божиим, мудростью, разумением, ведением и всяким искусством,
EXOD|35|32|составлять искусные ткани, работать из золота, серебра и меди,
EXOD|35|33|и резать камни для вставливания, и резать дерево, и делать всякую художественную работу;
EXOD|35|34|и способность учить [других] вложил в сердце его, его и Аголиава, сына Ахисамахова, из колена Данова;
EXOD|35|35|он исполнил сердце их мудростью, чтобы делать всякую работу резчика и искусного ткача, и вышивателя по голубой, пурпуровой, червленой и виссонной ткани, и ткачей, делающих всякую работу и составляющих искусные ткани.
EXOD|36|1|И стал работать Веселеил и Аголиав и все мудрые сердцем, которым Господь дал мудрость и разумение, чтоб уметь сделать всякую работу, потребную для святилища, как повелел Господь.
EXOD|36|2|И призвал Моисей Веселеила и Аголиава и всех мудрых сердцем, которым Господь дал мудрость, и всех, коих влекло сердце приступить к работе и работать.
EXOD|36|3|И взяли они от Моисея все приношения, которые принесли сыны Израилевы, на потребности святилища, чтобы работать. Между тем еще продолжали приносить к нему добровольные дары каждое утро.
EXOD|36|4|Тогда пришли все мудрые сердцем, производившие всякие работы святилища, каждый от своей работы, какою кто занимался,
EXOD|36|5|и сказали Моисею, говоря: народ много приносит, более нежели потребно для работ, какие повелел Господь сделать.
EXOD|36|6|И приказал Моисей, и объявлено было в стане, чтобы ни мужчина, ни женщина не делали уже ничего для приношения во святилище; и перестал народ приносить.
EXOD|36|7|Запаса было достаточно на всякие работы, какие надлежало делать, и даже осталось.
EXOD|36|8|И сделали все мудрые сердцем, занимавшиеся работою скинии: десять покрывал из крученого виссона и из голубой, пурпуровой и червленой [шерсти]; и херувимов сделали на них искусною работою;
EXOD|36|9|длина каждого покрывала двадцать восемь локтей, и ширина каждого покрывала четыре локтя: всем покрывалам одна мера.
EXOD|36|10|И соединил он пять покрывал одно с другим, и [другие] пять покрывал соединил одно с другим.
EXOD|36|11|И сделал петли голубого [цвета] на краю одного покрывала, где оно соединяется с другим; так же сделал он и на краю последнего покрывала, для соединения его с другим;
EXOD|36|12|пятьдесят петлей сделал он у одного покрывала, и пятьдесят петлей сделал в конце покрывала, где оно соединяется с другим; петли сии соответствовали одна другой;
EXOD|36|13|и сделал пятьдесят крючков золотых, и крючками соединил одно покрывало с другим, и стала скиния одно [целое].
EXOD|36|14|Потом сделал покрывала из козьей шерсти для покрытия скинии: одиннадцать покрывал сделал таких;
EXOD|36|15|длиною покрывало тридцать локтей, и шириною покрывало четыре локтя: одиннадцати покрывалам мера одна.
EXOD|36|16|И соединил он пять покрывал особо и шесть покрывал особо.
EXOD|36|17|И сделал пятьдесят петлей на краю покрывала крайнего, где оно соединяется с другим, и пятьдесят петлей сделал на краю покрывала, соединяющегося с другим;
EXOD|36|18|и сделал пятьдесят медных крючков для соединения покрова, чтоб составилось одно [целое].
EXOD|36|19|И сделал для скинии покров из красных бараньих кож и покрышку сверху из кож синих.
EXOD|36|20|И сделал брусья для скинии из дерева ситтим прямостоящие:
EXOD|36|21|десять локтей длина бруса, и полтора локтя ширина каждого бруса;
EXOD|36|22|у каждого бруса по два шипа, один против другого: так сделал он все брусья скинии.
EXOD|36|23|И сделал для скинии двадцать таких брусьев для полуденной стороны,
EXOD|36|24|и сорок серебряных подножий сделал под двадцать брусьев: два подножия под один брус для двух шипов его, и два подножия под другой брус для двух шипов его;
EXOD|36|25|и для другой стороны скинии, к северу, сделал двадцать брусьев
EXOD|36|26|и сорок серебряных подножий: два подножия под один брус, и два подножия под другой брус;
EXOD|36|27|а для задней стороны скинии, к западу, сделал шесть брусьев,
EXOD|36|28|и два бруса сделал для угла в скинии на заднюю сторону;
EXOD|36|29|и были они соединены внизу и соединены вверху к одному кольцу: так сделал он с ними обоими на обоих углах;
EXOD|36|30|и было восемь брусьев и серебряных подножий шестнадцать, по два подножия под каждый брус.
EXOD|36|31|И сделал шесты из дерева ситтим, пять для брусьев одной стороны скинии,
EXOD|36|32|и пять шестов для брусьев другой стороны скинии, и пять шестов для брусьев задней стороны скинии;
EXOD|36|33|и сделал внутренний шест, который проходил бы по средине брусьев от одного конца до другого;
EXOD|36|34|брусья обложил золотом, и кольца, в которые вкладываются шесты, сделал из золота, и шесты обложил золотом.
EXOD|36|35|И сделал завесу из голубой, пурпуровой и червленой [шерсти] и из крученого виссона, и искусною работою сделал на ней херувимов;
EXOD|36|36|и сделал для нее четыре столба из ситтим и обложил их золотом, с золотыми крючками, и вылил для них четыре серебряных подножия.
EXOD|36|37|И сделал завесу ко входу скинии из голубой, пурпуровой и червленой [шерсти] и из крученого виссона, узорчатой работы,
EXOD|36|38|и пять столбов для нее с крючками; и обложил верхи их и связи их золотом, и [вылил] пять медных подножий.
EXOD|37|1|И сделал Веселеил ковчег из дерева ситтим; длина его два локтя с половиною, ширина его полтора локтя и высота его полтора локтя;
EXOD|37|2|и обложил его чистым золотом внутри и снаружи и сделал вокруг него золотой венец;
EXOD|37|3|и вылил для него четыре кольца золотых, на четырех нижних углах его: два кольца на одной стороне его и два кольца на другой стороне его.
EXOD|37|4|И сделал шесты из дерева ситтим и обложил их золотом;
EXOD|37|5|и вложил шесты в кольца, по сторонам ковчега, чтобы носить ковчег.
EXOD|37|6|И сделал крышку из чистого золота: длина ее два локтя с половиною, а ширина полтора локтя.
EXOD|37|7|И сделал двух херувимов из золота: чеканной работы сделал их на обоих концах крышки,
EXOD|37|8|одного херувима с одного конца, а другого херувима с другого конца: выдавшимися из крышки сделал херувимов с обоих концов ее;
EXOD|37|9|и были херувимы с распростертыми вверх крыльями и покрывали крыльями своими крышку, а лицами своими были [обращены] друг к другу; к крышке [были] лица херувимов.
EXOD|37|10|И сделал стол из дерева ситтим длиною в два локтя, шириною в локоть и вышиною в полтора локтя,
EXOD|37|11|и обложил его золотом чистым, и сделал вокруг него золотой венец;
EXOD|37|12|и сделал вокруг него стенки в ладонь и сделал золотой венец у стенок его;
EXOD|37|13|и вылил для него четыре кольца золотых и утвердил кольца на четырех углах, у четырех ножек его;
EXOD|37|14|при стенках были кольца, чтобы влагать шесты для ношения стола;
EXOD|37|15|и сделал шесты из дерева ситтим и обложил их золотом для ношения стола.
EXOD|37|16|Потом сделал сосуды, принадлежавшие к столу: блюда, кадильницы, кружки и чаши, чтобы возливать ими, из чистого золота.
EXOD|37|17|И сделал светильник из золота чистого, чеканный сделал светильник; стебель его, ветви его, чашечки его, яблоки его и цветы его [выходили] из него;
EXOD|37|18|шесть ветвей выходило из боков его: три ветви светильника из одного бока его и три ветви светильника из другого бока его;
EXOD|37|19|три чашечки были наподобие миндального цветка, яблоко и цветы на одной ветви, и три чашечки наподобие миндального цветка, яблоко и цветы на другой ветви: так на [всех] шести ветвях, выходящих из светильника;
EXOD|37|20|а на [стебле] светильника было четыре чашечки наподобие миндального цветка с яблоками и цветами;
EXOD|37|21|у шести ветвей, выходящих из него, яблоко под первыми двумя ветвями, и яблоко под [вторыми] двумя ветвями, и яблоко под [третьими] двумя ветвями;
EXOD|37|22|яблоки и ветви их выходили из него; весь он [был] чеканный, цельный, из чистого золота.
EXOD|37|23|И сделал к нему семь лампад, и щипцы к нему и лотки к нему, из чистого золота;
EXOD|37|24|из таланта чистого золота сделал его со всеми принадлежностями его.
EXOD|37|25|И сделал жертвенник курения из дерева ситтим: длина его локоть и ширина его локоть, четыреугольный, вышина его два локтя; из него выходили роги его;
EXOD|37|26|и обложил его чистым золотом, верх его и стороны его кругом, и роги его, и сделал к нему золотой венец вокруг;
EXOD|37|27|под венцом его на двух углах его сделал два кольца золотых; с двух сторон его сделал их, чтобы вкладывать в них шесты для ношения его;
EXOD|37|28|шесты сделал из дерева ситтим и обложил их золотом.
EXOD|37|29|И сделал миро для священного помазания и курение благовонное, чистое, искусством составляющего масти.
EXOD|38|1|И сделал жертвенник всесожжения из дерева ситтим длиною в пять локтей и шириною в пять локтей, четыреугольный, вышиною в три локтя;
EXOD|38|2|и сделал роги на четырех углах его, так что из него выходили роги, и обложил его медью.
EXOD|38|3|И сделал все принадлежности жертвенника: горшки, лопатки, чаши, вилки и угольницы; все принадлежности его сделал из меди.
EXOD|38|4|И сделал для жертвенника решетку, род сетки, из меди, по окраине его внизу до половины его;
EXOD|38|5|и сделал четыре кольца на четырех углах медной решетки для вкладывания шестов.
EXOD|38|6|И сделал шесты из дерева ситтим, и обложил их медью,
EXOD|38|7|и вложил шесты в кольца на боках жертвенника, чтобы носить его посредством их; пустой внутри из досок сделал его.
EXOD|38|8|И сделал умывальник из меди и подножие его из меди с изящными изображениями, украшающими вход скинии собрания.
EXOD|38|9|И сделал двор: с полуденной стороны, к югу, завесы из крученого виссона, длиною во сто локтей;
EXOD|38|10|столбов для них двадцать и подножий к ним двадцать медных; крючки у столбов и связи их из серебра.
EXOD|38|11|И по северной стороне – [завесы] во сто локтей; столбов для них двадцать и подножий к ним двадцать медных; крючки у столбов и связи их из серебра.
EXOD|38|12|И с западной стороны – завесы в пятьдесят локтей, столбов для них десять и подножий к ним десять; крючки у столбов и связи их из серебра.
EXOD|38|13|И с передней стороны к востоку – [завесы] в пятьдесят локтей.
EXOD|38|14|Для одной стороны [ворот двора] – завесы в пятнадцать локтей, столбов для них три и подножий к ним три;
EXOD|38|15|и для другой стороны – завесы в пятнадцать локтей, столбов для них три и подножий к ним три.
EXOD|38|16|Все завесы во все стороны двора из крученого виссона,
EXOD|38|17|а подножия у столбов из меди, крючки у столбов и связи их из серебра; верхи же у них обложены серебром, и все столбы двора соединены связями серебряными.
EXOD|38|18|Завеса же для ворот двора узорчатой работы из голубой, пурпуровой и червленой [шерсти] и из крученого виссона, длиною в двадцать локтей, вышиною в пять локтей, по всему протяжению, подобно завесам двора;
EXOD|38|19|и столбов для нее четыре, и подножий к ним четыре медных; крючки у них серебряные, а верхи их обложены серебром, и связи их серебряные.
EXOD|38|20|Все колья вокруг скинии и двора медные.
EXOD|38|21|Вот исчисление того, что употреблено для скинии откровения, сделанное по повелению Моисея, посредством левитов под надзором Ифамара, сына Ааронова, священника.
EXOD|38|22|Делал же все, что повелел Господь Моисею, Веселеил, сын Урии, сына Ора, из колена Иудина,
EXOD|38|23|и с ним Аголиав, сын Ахисамахов, из колена Данова, резчик и искусный ткач и вышиватель по голубой, пурпуровой, червленой и виссоновой [ткани].
EXOD|38|24|Всего золота, употребленного в дело на все принадлежности святилища, золота, принесенного в дар, было двадцать девять талантов и семьсот тридцать сиклей, сиклей священных;
EXOD|38|25|серебра же от исчисленных [лиц] общества сто талантов и тысяча семьсот семьдесят пять сиклей, сиклей священных;
EXOD|38|26|с шестисот трех тысяч пятисот пятидесяти человек, с каждого поступившего в исчисление, от двадцати лет и выше, по полсиклю с человека, считая на сикль священный.
EXOD|38|27|Сто талантов серебра употреблено на вылитие подножий святилища и подножий у завесы; сто подножий из ста талантов, по таланту на подножие;
EXOD|38|28|а из тысячи семисот семидесяти пяти [сиклей] сделал он крючки у столбов и покрыл верхи их и сделал связи для них.
EXOD|38|29|Меди же, принесенной в дар, было семьдесят талантов и две тысячи четыреста сиклей;
EXOD|38|30|из нее сделал он подножия [для столбов] у входа в скинию свидетельства, и жертвенник медный, и решетку медную для него, и все сосуды жертвенника,
EXOD|38|31|и подножия [для столбов] всего двора, и подножия [для] [столбов] ворот двора, и все колья скинии и все колья вокруг двора.
EXOD|39|1|Из голубой же, пурпуровой и червленой [шерсти] сделали они служебные одежды, для служения во святилище; также сделали священные одежды Аарону, как повелел Господь Моисею.
EXOD|39|2|И сделал ефод из золота, из голубой, пурпуровой и червленой [шерсти] и из крученого виссона;
EXOD|39|3|и разбили они золото в листы и вытянули нити, чтобы воткать их между голубыми, пурпуровыми, червлеными и виссонными [нитями], искусною работою.
EXOD|39|4|И сделали у него нарамники связывающие; на обоих концах своих он был связан.
EXOD|39|5|И пояс ефода, который поверх его, одинаковой с ним работы, [сделан] [был] из золота, из голубой, пурпуровой и червленой [шерсти] и крученого виссона, как повелел Господь Моисею.
EXOD|39|6|И обделали камни ониксовые, вставив их в золотые гнезда и вырезав на них имена сынов Израилевых, как вырезывают на печати;
EXOD|39|7|и положил он их на нарамники ефода, в память сынов Израилевых, как повелел Господь Моисею.
EXOD|39|8|И сделал наперсник искусною работою, такою же работою, как ефод, из золота, из голубой, пурпуровой и червленой [шерсти] и из крученого виссона;
EXOD|39|9|он был четыреугольный; двойной сделали они наперсник в пядень длиною и в пядень шириною, двойной он был;
EXOD|39|10|и вставили в него в четыре ряда камни. Рядом: рубин, топаз, изумруд, – это первый ряд;
EXOD|39|11|во втором ряду: карбункул, сапфир и алмаз;
EXOD|39|12|в третьем ряду: яхонт, агат и аметист;
EXOD|39|13|в четвертом ряду: хризолит, оникс и яспис; и вставлены они в золотых гнездах.
EXOD|39|14|Камней было по числу имен сынов Израилевых: двенадцать было их, по числу имен их, и на каждом из них вырезано было, [как] на печати, по одному имени, для двенадцати колен.
EXOD|39|15|К наперснику сделали толстые цепочки витою работою из чистого золота;
EXOD|39|16|и сделали два золотых гнезда и два золотых кольца и прикрепили два кольца к двум концам наперсника;
EXOD|39|17|и вдели обе плетеные цепочки из золота в два кольца по концам наперсника,
EXOD|39|18|а два конца двух цепочек прикрепили к двум гнездам и прикрепили их к нарамникам ефода с лицевой стороны его;
EXOD|39|19|еще сделали два кольца золотых и прикрепили к двум [другим] концам наперсника, на той стороне, которая находится к ефоду внутрь;
EXOD|39|20|и еще сделали два кольца золотых и прикрепили их к двум нарамникам ефода снизу, с лицевой стороны его, у соединения его над поясом ефода;
EXOD|39|21|и прикрепили наперсник кольцами его к кольцам ефода посредством шнура из голубой [шерсти], чтобы он был над поясом ефода, и чтобы не отставал наперсник от ефода, как повелел Господь Моисею.
EXOD|39|22|И сделал верхнюю ризу к ефоду, тканую, всю из голубой [шерсти],
EXOD|39|23|и среди верхней ризы отверстие, как отверстие у брони, и вокруг него обшивку, чтобы не дралось;
EXOD|39|24|по подолу верхней ризы сделали они яблоки из голубой, пурпуровой и червленой [шерсти];
EXOD|39|25|и сделали позвонки из чистого золота и повесили позвонки между яблоками по подолу верхней ризы кругом;
EXOD|39|26|позвонок и яблоко, позвонок и яблоко, по подолу верхней ризы кругом для служения, как повелел Господь Моисею.
EXOD|39|27|И сделали для Аарона и для сыновей его хитоны из виссона, тканые,
EXOD|39|28|и кидар из виссона, и головные повязки из виссона, и нижнее льняное платье из крученого виссона,
EXOD|39|29|и пояс из крученого виссона и из голубой, пурпуровой и червленой [шерсти], узорчатой работы, как повелел Господь Моисею.
EXOD|39|30|И сделали полированную дощечку, диадиму святыни, из чистого золота, и начертали на ней письмена, как вырезывают на печати: Святыня Господня;
EXOD|39|31|и прикрепили к ней шнур из голубой [шерсти], чтобы привязать ее к кидару сверху, как повелел Господь Моисею.
EXOD|39|32|Так кончена была вся работа для скинии собрания; и сделали сыны Израилевы все: как повелел Господь Моисею, так и сделали.
EXOD|39|33|И принесли к Моисею скинию, покров и все принадлежности ее, крючки ее, брусья ее, шесты ее, столбы ее и подножия ее,
EXOD|39|34|покров из кож бараньих красных и покров из кож синих и завесу закрывающую,
EXOD|39|35|ковчег откровения и шесты его, и крышку,
EXOD|39|36|стол со всеми принадлежностями его и хлебы предложения,
EXOD|39|37|светильник из чистого золота, лампады его, лампады расставленные на нем и все принадлежности его, и елей для освещения,
EXOD|39|38|золотой жертвенник и елей помазания, и благовония для курения, и завесу ко входу в скинию,
EXOD|39|39|жертвенник медный и медную решетку к нему, шесты его и все принадлежности его, умывальник и подножие его,
EXOD|39|40|завесы двора, столбы и подножия, завесу к воротам двора, веревки и колья и все вещи, принадлежащие к служению в скинии собрания,
EXOD|39|41|одежды служебные для служения во святилище, священные одежды Аарону священнику и одежды сыновьям его для священнодействия.
EXOD|39|42|Как повелел Господь Моисею, так и сделали сыны Израилевы все сии работы.
EXOD|39|43|И увидел Моисей всю работу, и вот они сделали ее: как повелел Господь, так и сделали. И благословил их Моисей.
EXOD|40|1|И сказал Господь Моисею, говоря:
EXOD|40|2|в первый месяц, в первый день месяца поставь скинию собрания,
EXOD|40|3|и поставь в ней ковчег откровения, и закрой ковчег завесою;
EXOD|40|4|и внеси стол и расставь на нем все вещи его, и внеси светильник и поставь на нем лампады его;
EXOD|40|5|и поставь золотой жертвенник для курения пред ковчегом откровения и повесь завесу у входа в скинию.
EXOD|40|6|и поставь жертвенник всесожжения пред входом в скинию собрания;
EXOD|40|7|и поставь умывальник между скиниею собрания и между жертвенником и влей в него воды;
EXOD|40|8|и поставь двор кругом и повесь завесу в воротах двора.
EXOD|40|9|И возьми елея помазания, и помажь скинию и все, что в ней, и освяти ее и все принадлежности ее, и будет свята;
EXOD|40|10|помажь жертвенник всесожжения и все принадлежности его, и освяти жертвенник, и будет жертвенник святыня великая;
EXOD|40|11|и помажь умывальник и подножие его и освяти его.
EXOD|40|12|И приведи Аарона и сынов его ко входу в скинию собрания и омой их водою,
EXOD|40|13|и облеки Аарона в священные одежды, и помажь его, и освяти его, чтобы он был священником Мне.
EXOD|40|14|И сынов его приведи, и одень их в хитоны,
EXOD|40|15|и помажь их, как помазал ты отца их, чтобы они были священниками Мне, и помазание их посвятит их в вечное священство в роды их.
EXOD|40|16|И сделал Моисей все, как повелел ему Господь, так и сделал.
EXOD|40|17|В первый месяц второго года, в первый [день] месяца поставлена скиния.
EXOD|40|18|И поставил Моисей скинию, положил подножия ее, поставил брусья ее, положил шесты и поставил столбы ее,
EXOD|40|19|распростер покров над скиниею, и положил покрышку поверх сего покрова, как повелел Господь Моисею.
EXOD|40|20|И взял и положил откровение в ковчег, и вложил шесты в [кольца] ковчега, и положил крышку на ковчег сверху;
EXOD|40|21|и внес ковчег в скинию, и повесил завесу, и закрыл ковчег откровения, как повелел Господь Моисею.
EXOD|40|22|И поставил стол в скинии собрания, на северной стороне скинии, вне завесы,
EXOD|40|23|и разложил на нем ряд хлебов пред Господом, как повелел Господь Моисею.
EXOD|40|24|И поставил светильник в скинии собрания против стола, на южной стороне скинии,
EXOD|40|25|и поставил лампады пред Господом, как повелел Господь Моисею.
EXOD|40|26|И поставил золотой жертвенник в скинии собрания пред завесою
EXOD|40|27|и воскурил на нем благовонное курение, как повелел Господь Моисею.
EXOD|40|28|И повесил завесу при входе в скинию;
EXOD|40|29|и жертвенник всесожжения поставил у входа в скинию собрания и принес на нем всесожжения и приношение хлебное, как повелел Господь Моисею.
EXOD|40|30|И поставил умывальник между скиниею собрания и жертвенником и налил в него воды для омовения,
EXOD|40|31|и омывали из него Моисей и Аарон и сыны его руки свои и ноги свои:
EXOD|40|32|когда они входили в скинию собрания и подходили к жертвеннику, тогда омывались, как повелел Господь Моисею.
EXOD|40|33|И поставил двор вокруг скинии и жертвенника и повесил завесу в воротах двора. И так окончил Моисей дело.
EXOD|40|34|И покрыло облако скинию собрания, и слава Господня наполнила скинию;
EXOD|40|35|и не мог Моисей войти в скинию собрания, потому что осеняло ее облако, и слава Господня наполняла скинию.
EXOD|40|36|Когда поднималось облако от скинии, тогда отправлялись в путь сыны Израилевы во все путешествие свое;
EXOD|40|37|если же не поднималось облако, то и они не отправлялись в путь, доколе оно не поднималось,
EXOD|40|38|ибо облако Господне стояло над скиниею днем, и огонь был ночью в ней пред глазами всего дома Израилева во все путешествие их.
