JOHN|1|1|in principio erat Verbum et Verbum erat apud Deum et Deus erat Verbum
JOHN|1|2|hoc erat in principio apud Deum
JOHN|1|3|omnia per ipsum facta sunt et sine ipso factum est nihil quod factum est
JOHN|1|4|in ipso vita erat et vita erat lux hominum
JOHN|1|5|et lux in tenebris lucet et tenebrae eam non conprehenderunt
JOHN|1|6|fuit homo missus a Deo cui nomen erat Iohannes
JOHN|1|7|hic venit in testimonium ut testimonium perhiberet de lumine ut omnes crederent per illum
JOHN|1|8|non erat ille lux sed ut testimonium perhiberet de lumine
JOHN|1|9|erat lux vera quae inluminat omnem hominem venientem in mundum
JOHN|1|10|in mundo erat et mundus per ipsum factus est et mundus eum non cognovit
JOHN|1|11|in propria venit et sui eum non receperunt
JOHN|1|12|quotquot autem receperunt eum dedit eis potestatem filios Dei fieri his qui credunt in nomine eius
JOHN|1|13|qui non ex sanguinibus neque ex voluntate carnis neque ex voluntate viri sed ex Deo nati sunt
JOHN|1|14|et Verbum caro factum est et habitavit in nobis et vidimus gloriam eius gloriam quasi unigeniti a Patre plenum gratiae et veritatis
JOHN|1|15|Iohannes testimonium perhibet de ipso et clamat dicens hic erat quem dixi vobis qui post me venturus est ante me factus est quia prior me erat
JOHN|1|16|et de plenitudine eius nos omnes accepimus et gratiam pro gratia
JOHN|1|17|quia lex per Mosen data est gratia et veritas per Iesum Christum facta est
JOHN|1|18|Deum nemo vidit umquam unigenitus Filius qui est in sinu Patris ipse enarravit
JOHN|1|19|et hoc est testimonium Iohannis quando miserunt Iudaei ab Hierosolymis sacerdotes et Levitas ad eum ut interrogarent eum tu quis es
JOHN|1|20|et confessus est et non negavit et confessus est quia non sum ego Christus
JOHN|1|21|et interrogaverunt eum quid ergo Helias es tu et dicit non sum propheta es tu et respondit non
JOHN|1|22|dixerunt ergo ei quis es ut responsum demus his qui miserunt nos quid dicis de te ipso
JOHN|1|23|ait ego vox clamantis in deserto dirigite viam Domini sicut dixit Esaias propheta
JOHN|1|24|et qui missi fuerant erant ex Pharisaeis
JOHN|1|25|et interrogaverunt eum et dixerunt ei quid ergo baptizas si tu non es Christus neque Helias neque propheta
JOHN|1|26|respondit eis Iohannes dicens ego baptizo in aqua medius autem vestrum stetit quem vos non scitis
JOHN|1|27|ipse est qui post me venturus est qui ante me factus est cuius ego non sum dignus ut solvam eius corrigiam calciamenti
JOHN|1|28|haec in Bethania facta sunt trans Iordanen ubi erat Iohannes baptizans
JOHN|1|29|altera die videt Iohannes Iesum venientem ad se et ait ecce agnus Dei qui tollit peccatum mundi
JOHN|1|30|hic est de quo dixi post me venit vir qui ante me factus est quia prior me erat
JOHN|1|31|et ego nesciebam eum sed ut manifestaretur Israhel propterea veni ego in aqua baptizans
JOHN|1|32|et testimonium perhibuit Iohannes dicens quia vidi Spiritum descendentem quasi columbam de caelo et mansit super eum
JOHN|1|33|et ego nesciebam eum sed qui misit me baptizare in aqua ille mihi dixit super quem videris Spiritum descendentem et manentem super eum hic est qui baptizat in Spiritu Sancto
JOHN|1|34|et ego vidi et testimonium perhibui quia hic est Filius Dei
JOHN|1|35|altera die iterum stabat Iohannes et ex discipulis eius duo
JOHN|1|36|et respiciens Iesum ambulantem dicit ecce agnus Dei
JOHN|1|37|et audierunt eum duo discipuli loquentem et secuti sunt Iesum
JOHN|1|38|conversus autem Iesus et videns eos sequentes dicit eis quid quaeritis qui dixerunt ei rabbi quod dicitur interpretatum magister ubi habitas
JOHN|1|39|dicit eis venite et videte venerunt et viderunt ubi maneret et apud eum manserunt die illo hora autem erat quasi decima
JOHN|1|40|erat autem Andreas frater Simonis Petri unus ex duobus qui audierant ab Iohanne et secuti fuerant eum
JOHN|1|41|invenit hic primum fratrem suum Simonem et dicit ei invenimus Messiam quod est interpretatum Christus
JOHN|1|42|et adduxit eum ad Iesum intuitus autem eum Iesus dixit tu es Simon filius Iohanna tu vocaberis Cephas quod interpretatur Petrus
JOHN|1|43|in crastinum voluit exire in Galilaeam et invenit Philippum et dicit ei Iesus sequere me
JOHN|1|44|erat autem Philippus a Bethsaida civitate Andreae et Petri
JOHN|1|45|invenit Philippus Nathanahel et dicit ei quem scripsit Moses in lege et prophetae invenimus Iesum filium Ioseph a Nazareth
JOHN|1|46|et dixit ei Nathanahel a Nazareth potest aliquid boni esse dicit ei Philippus veni et vide
JOHN|1|47|vidit Iesus Nathanahel venientem ad se et dicit de eo ecce vere Israhelita in quo dolus non est
JOHN|1|48|dicit ei Nathanahel unde me nosti respondit Iesus et dixit ei priusquam te Philippus vocaret cum esses sub ficu vidi te
JOHN|1|49|respondit ei Nathanahel et ait rabbi tu es Filius Dei tu es rex Israhel
JOHN|1|50|respondit Iesus et dixit ei quia dixi tibi vidi te sub ficu credis maius his videbis
JOHN|1|51|et dicit ei amen amen dico vobis videbitis caelum apertum et angelos Dei ascendentes et descendentes supra Filium hominis
JOHN|2|1|et die tertio nuptiae factae sunt in Cana Galilaeae et erat mater Iesu ibi
JOHN|2|2|vocatus est autem ibi et Iesus et discipuli eius ad nuptias
JOHN|2|3|et deficiente vino dicit mater Iesu ad eum vinum non habent
JOHN|2|4|et dicit ei Iesus quid mihi et tibi est mulier nondum venit hora mea
JOHN|2|5|dicit mater eius ministris quodcumque dixerit vobis facite
JOHN|2|6|erant autem ibi lapideae hydriae sex positae secundum purificationem Iudaeorum capientes singulae metretas binas vel ternas
JOHN|2|7|dicit eis Iesus implete hydrias aqua et impleverunt eas usque ad summum
JOHN|2|8|et dicit eis Iesus haurite nunc et ferte architriclino et tulerunt
JOHN|2|9|ut autem gustavit architriclinus aquam vinum factam et non sciebat unde esset ministri autem sciebant qui haurierant aquam vocat sponsum architriclinus
JOHN|2|10|et dicit ei omnis homo primum bonum vinum ponit et cum inebriati fuerint tunc id quod deterius est tu servasti bonum vinum usque adhuc
JOHN|2|11|hoc fecit initium signorum Iesus in Cana Galilaeae et manifestavit gloriam suam et crediderunt in eum discipuli eius
JOHN|2|12|post hoc descendit Capharnaum ipse et mater eius et fratres eius et discipuli eius et ibi manserunt non multis diebus
JOHN|2|13|et prope erat pascha Iudaeorum et ascendit Hierosolyma Iesus
JOHN|2|14|et invenit in templo vendentes boves et oves et columbas et nummularios sedentes
JOHN|2|15|et cum fecisset quasi flagellum de funiculis omnes eiecit de templo oves quoque et boves et nummulariorum effudit aes et mensas subvertit
JOHN|2|16|et his qui columbas vendebant dixit auferte ista hinc nolite facere domum Patris mei domum negotiationis
JOHN|2|17|recordati vero sunt discipuli eius quia scriptum est zelus domus tuae comedit me
JOHN|2|18|responderunt ergo Iudaei et dixerunt ei quod signum ostendis nobis quia haec facis
JOHN|2|19|respondit Iesus et dixit eis solvite templum hoc et in tribus diebus excitabo illud
JOHN|2|20|dixerunt ergo Iudaei quadraginta et sex annis aedificatum est templum hoc et tu tribus diebus excitabis illud
JOHN|2|21|ille autem dicebat de templo corporis sui
JOHN|2|22|cum ergo resurrexisset a mortuis recordati sunt discipuli eius quia hoc dicebat et crediderunt scripturae et sermoni quem dixit Iesus
JOHN|2|23|cum autem esset Hierosolymis in pascha in die festo multi crediderunt in nomine eius videntes signa eius quae faciebat
JOHN|2|24|ipse autem Iesus non credebat semet ipsum eis eo quod ipse nosset omnes
JOHN|2|25|et quia opus ei non erat ut quis testimonium perhiberet de homine ipse enim sciebat quid esset in homine
JOHN|3|1|erat autem homo ex Pharisaeis Nicodemus nomine princeps Iudaeorum
JOHN|3|2|hic venit ad eum nocte et dixit ei rabbi scimus quia a Deo venisti magister nemo enim potest haec signa facere quae tu facis nisi fuerit Deus cum eo
JOHN|3|3|respondit Iesus et dixit ei amen amen dico tibi nisi quis natus fuerit denuo non potest videre regnum Dei
JOHN|3|4|dicit ad eum Nicodemus quomodo potest homo nasci cum senex sit numquid potest in ventrem matris suae iterato introire et nasci
JOHN|3|5|respondit Iesus amen amen dico tibi nisi quis renatus fuerit ex aqua et Spiritu non potest introire in regnum Dei
JOHN|3|6|quod natum est ex carne caro est et quod natum est ex Spiritu spiritus est
JOHN|3|7|non mireris quia dixi tibi oportet vos nasci denuo
JOHN|3|8|Spiritus ubi vult spirat et vocem eius audis sed non scis unde veniat et quo vadat sic est omnis qui natus est ex Spiritu
JOHN|3|9|respondit Nicodemus et dixit ei quomodo possunt haec fieri
JOHN|3|10|respondit Iesus et dixit ei tu es magister Israhel et haec ignoras
JOHN|3|11|amen amen dico tibi quia quod scimus loquimur et quod vidimus testamur et testimonium nostrum non accipitis
JOHN|3|12|si terrena dixi vobis et non creditis quomodo si dixero vobis caelestia credetis
JOHN|3|13|et nemo ascendit in caelum nisi qui descendit de caelo Filius hominis qui est in caelo
JOHN|3|14|et sicut Moses exaltavit serpentem in deserto ita exaltari oportet Filium hominis
JOHN|3|15|ut omnis qui credit in ipso non pereat sed habeat vitam aeternam
JOHN|3|16|sic enim dilexit Deus mundum ut Filium suum unigenitum daret ut omnis qui credit in eum non pereat sed habeat vitam aeternam
JOHN|3|17|non enim misit Deus Filium suum in mundum ut iudicet mundum sed ut salvetur mundus per ipsum
JOHN|3|18|qui credit in eum non iudicatur qui autem non credit iam iudicatus est quia non credidit in nomine unigeniti Filii Dei
JOHN|3|19|hoc est autem iudicium quia lux venit in mundum et dilexerunt homines magis tenebras quam lucem erant enim eorum mala opera
JOHN|3|20|omnis enim qui mala agit odit lucem et non venit ad lucem ut non arguantur opera eius
JOHN|3|21|qui autem facit veritatem venit ad lucem ut manifestentur eius opera quia in Deo sunt facta
JOHN|3|22|post haec venit Iesus et discipuli eius in iudaeam terram et illic demorabatur cum eis et baptizabat
JOHN|3|23|erat autem et Iohannes baptizans in Aenon iuxta Salim quia aquae multae erant illic et adveniebant et baptizabantur
JOHN|3|24|nondum enim missus fuerat in carcerem Iohannes
JOHN|3|25|facta est ergo quaestio ex discipulis Iohannis cum Iudaeis de purificatione
JOHN|3|26|et venerunt ad Iohannem et dixerunt ei rabbi qui erat tecum trans Iordanen cui tu testimonium perhibuisti ecce hic baptizat et omnes veniunt ad eum
JOHN|3|27|respondit Iohannes et dixit non potest homo accipere quicquam nisi fuerit ei datum de caelo
JOHN|3|28|ipsi vos mihi testimonium perhibetis quod dixerim ego non sum Christus sed quia missus sum ante illum
JOHN|3|29|qui habet sponsam sponsus est amicus autem sponsi qui stat et audit eum gaudio gaudet propter vocem sponsi hoc ergo gaudium meum impletum est
JOHN|3|30|illum oportet crescere me autem minui
JOHN|3|31|qui desursum venit supra omnes est qui est de terra de terra est et de terra loquitur qui de caelo venit supra omnes est
JOHN|3|32|et quod vidit et audivit hoc testatur et testimonium eius nemo accipit
JOHN|3|33|qui accipit eius testimonium signavit quia Deus verax est
JOHN|3|34|quem enim misit Deus verba Dei loquitur non enim ad mensuram dat Deus Spiritum
JOHN|3|35|Pater diligit Filium et omnia dedit in manu eius
JOHN|3|36|qui credit in Filium habet vitam aeternam qui autem incredulus est Filio non videbit vitam sed ira Dei manet super eum
JOHN|4|1|ut ergo cognovit Iesus quia audierunt Pharisaei quia Iesus plures discipulos facit et baptizat quam Iohannes
JOHN|4|2|quamquam Iesus non baptizaret sed discipuli eius
JOHN|4|3|reliquit Iudaeam et abiit iterum in Galilaeam
JOHN|4|4|oportebat autem eum transire per Samariam
JOHN|4|5|venit ergo in civitatem Samariae quae dicitur Sychar iuxta praedium quod dedit Iacob Ioseph filio suo
JOHN|4|6|erat autem ibi fons Iacob Iesus ergo fatigatus ex itinere sedebat sic super fontem hora erat quasi sexta
JOHN|4|7|venit mulier de Samaria haurire aquam dicit ei Iesus da mihi bibere
JOHN|4|8|discipuli enim eius abierant in civitatem ut cibos emerent
JOHN|4|9|dicit ergo ei mulier illa samaritana quomodo tu Iudaeus cum sis bibere a me poscis quae sum mulier samaritana non enim coutuntur Iudaei Samaritanis
JOHN|4|10|respondit Iesus et dixit ei si scires donum Dei et quis est qui dicit tibi da mihi bibere tu forsitan petisses ab eo et dedisset tibi aquam vivam
JOHN|4|11|dicit ei mulier Domine neque in quo haurias habes et puteus altus est unde ergo habes aquam vivam
JOHN|4|12|numquid tu maior es patre nostro Iacob qui dedit nobis puteum et ipse ex eo bibit et filii eius et pecora eius
JOHN|4|13|respondit Iesus et dixit ei omnis qui bibit ex aqua hac sitiet iterum qui autem biberit ex aqua quam ego dabo ei non sitiet in aeternum
JOHN|4|14|sed aqua quam dabo ei fiet in eo fons aquae salientis in vitam aeternam
JOHN|4|15|dicit ad eum mulier Domine da mihi hanc aquam ut non sitiam neque veniam huc haurire
JOHN|4|16|dicit ei Iesus vade voca virum tuum et veni huc
JOHN|4|17|respondit mulier et dixit non habeo virum dicit ei Iesus bene dixisti quia non habeo virum
JOHN|4|18|quinque enim viros habuisti et nunc quem habes non est tuus vir hoc vere dixisti
JOHN|4|19|dicit ei mulier Domine video quia propheta es tu
JOHN|4|20|patres nostri in monte hoc adoraverunt et vos dicitis quia Hierosolymis est locus ubi adorare oportet
JOHN|4|21|dicit ei Iesus mulier crede mihi quia veniet hora quando neque in monte hoc neque in Hierosolymis adorabitis Patrem
JOHN|4|22|vos adoratis quod nescitis nos adoramus quod scimus quia salus ex Iudaeis est
JOHN|4|23|sed venit hora et nunc est quando veri adoratores adorabunt Patrem in spiritu et veritate nam et Pater tales quaerit qui adorent eum
JOHN|4|24|spiritus est Deus et eos qui adorant eum in spiritu et veritate oportet adorare
JOHN|4|25|dicit ei mulier scio quia Messias venit qui dicitur Christus cum ergo venerit ille nobis adnuntiabit omnia
JOHN|4|26|dicit ei Iesus ego sum qui loquor tecum
JOHN|4|27|et continuo venerunt discipuli eius et mirabantur quia cum muliere loquebatur nemo tamen dixit quid quaeris aut quid loqueris cum ea
JOHN|4|28|reliquit ergo hydriam suam mulier et abiit in civitatem et dicit illis hominibus
JOHN|4|29|venite videte hominem qui dixit mihi omnia quaecumque feci numquid ipse est Christus
JOHN|4|30|exierunt de civitate et veniebant ad eum
JOHN|4|31|interea rogabant eum discipuli dicentes rabbi manduca
JOHN|4|32|ille autem dixit eis ego cibum habeo manducare quem vos nescitis
JOHN|4|33|dicebant ergo discipuli ad invicem numquid aliquis adtulit ei manducare
JOHN|4|34|dicit eis Iesus meus cibus est ut faciam voluntatem eius qui misit me ut perficiam opus eius
JOHN|4|35|nonne vos dicitis quod adhuc quattuor menses sunt et messis venit ecce dico vobis levate oculos vestros et videte regiones quia albae sunt iam ad messem
JOHN|4|36|et qui metit mercedem accipit et congregat fructum in vitam aeternam ut et qui seminat simul gaudeat et qui metit
JOHN|4|37|in hoc enim est verbum verum quia alius est qui seminat et alius est qui metit
JOHN|4|38|ego misi vos metere quod vos non laborastis alii laboraverunt et vos in laborem eorum introistis
JOHN|4|39|ex civitate autem illa multi crediderunt in eum Samaritanorum propter verbum mulieris testimonium perhibentis quia dixit mihi omnia quaecumque feci
JOHN|4|40|cum venissent ergo ad illum Samaritani rogaverunt eum ut ibi maneret et mansit ibi duos dies
JOHN|4|41|et multo plures crediderunt propter sermonem eius
JOHN|4|42|et mulieri dicebant quia iam non propter tuam loquellam credimus ipsi enim audivimus et scimus quia hic est vere salvator mundi
JOHN|4|43|post duos autem dies exiit inde et abiit in Galilaeam
JOHN|4|44|ipse enim Iesus testimonium perhibuit quia propheta in sua patria honorem non habet
JOHN|4|45|cum ergo venisset in Galilaeam exceperunt eum Galilaei cum omnia vidissent quae fecerat Hierosolymis in die festo et ipsi enim venerant in diem festum
JOHN|4|46|venit ergo iterum in Cana Galilaeae ubi fecit aquam vinum et erat quidam regulus cuius filius infirmabatur Capharnaum
JOHN|4|47|hic cum audisset quia Iesus adveniret a Iudaea in Galilaeam abiit ad eum et rogabat eum ut descenderet et sanaret filium eius incipiebat enim mori
JOHN|4|48|dixit ergo Iesus ad eum nisi signa et prodigia videritis non creditis
JOHN|4|49|dicit ad eum regulus Domine descende priusquam moriatur filius meus
JOHN|4|50|dicit ei Iesus vade filius tuus vivit credidit homo sermoni quem dixit ei Iesus et ibat
JOHN|4|51|iam autem eo descendente servi occurrerunt ei et nuntiaverunt dicentes quia filius eius viveret
JOHN|4|52|interrogabat ergo horam ab eis in qua melius habuerit et dixerunt ei quia heri hora septima reliquit eum febris
JOHN|4|53|cognovit ergo pater quia illa hora erat in qua dixit ei Iesus filius tuus vivit et credidit ipse et domus eius tota
JOHN|4|54|hoc iterum secundum signum fecit Iesus cum venisset a Iudaea in Galilaeam
JOHN|5|1|post haec erat dies festus Iudaeorum et ascendit Iesus Hierosolymis
JOHN|5|2|est autem Hierosolymis super Probatica piscina quae cognominatur hebraice Bethsaida quinque porticus habens
JOHN|5|3|in his iacebat multitudo magna languentium caecorum claudorum aridorum expectantium aquae motum
JOHN|5|4|
JOHN|5|5|erat autem quidam homo ibi triginta et octo annos habens in infirmitate sua
JOHN|5|6|hunc cum vidisset Iesus iacentem et cognovisset quia multum iam tempus habet dicit ei vis sanus fieri
JOHN|5|7|respondit ei languidus Domine hominem non habeo ut cum turbata fuerit aqua mittat me in piscinam dum venio enim ego alius ante me descendit
JOHN|5|8|dicit ei Iesus surge tolle grabattum tuum et ambula
JOHN|5|9|et statim sanus factus est homo et sustulit grabattum suum et ambulabat erat autem sabbatum in illo die
JOHN|5|10|dicebant Iudaei illi qui sanatus fuerat sabbatum est non licet tibi tollere grabattum tuum
JOHN|5|11|respondit eis qui me fecit sanum ille mihi dixit tolle grabattum tuum et ambula
JOHN|5|12|interrogaverunt ergo eum quis est ille homo qui dixit tibi tolle grabattum tuum et ambula
JOHN|5|13|is autem qui sanus fuerat effectus nesciebat quis esset Iesus enim declinavit turba constituta in loco
JOHN|5|14|postea invenit eum Iesus in templo et dixit illi ecce sanus factus es iam noli peccare ne deterius tibi aliquid contingat
JOHN|5|15|abiit ille homo et nuntiavit Iudaeis quia Iesus esset qui fecit eum sanum
JOHN|5|16|propterea persequebantur Iudaei Iesum quia haec faciebat in sabbato
JOHN|5|17|Iesus autem respondit eis Pater meus usque modo operatur et ego operor
JOHN|5|18|propterea ergo magis quaerebant eum Iudaei interficere quia non solum solvebat sabbatum sed et Patrem suum dicebat Deum aequalem se faciens Deo respondit itaque Iesus et dixit eis
JOHN|5|19|amen amen dico vobis non potest Filius a se facere quicquam nisi quod viderit Patrem facientem quaecumque enim ille fecerit haec et Filius similiter facit
JOHN|5|20|Pater enim diligit Filium et omnia demonstrat ei quae ipse facit et maiora his demonstrabit ei opera ut vos miremini
JOHN|5|21|sicut enim Pater suscitat mortuos et vivificat sic et Filius quos vult vivificat
JOHN|5|22|neque enim Pater iudicat quemquam sed iudicium omne dedit Filio
JOHN|5|23|ut omnes honorificent Filium sicut honorificant Patrem qui non honorificat Filium non honorificat Patrem qui misit illum
JOHN|5|24|amen amen dico vobis quia qui verbum meum audit et credit ei qui misit me habet vitam aeternam et in iudicium non venit sed transit a morte in vitam
JOHN|5|25|amen amen dico vobis quia venit hora et nunc est quando mortui audient vocem Filii Dei et qui audierint vivent
JOHN|5|26|sicut enim Pater habet vitam in semet ipso sic dedit et Filio vitam habere in semet ipso
JOHN|5|27|et potestatem dedit ei et iudicium facere quia Filius hominis est
JOHN|5|28|nolite mirari hoc quia venit hora in qua omnes qui in monumentis sunt audient vocem eius
JOHN|5|29|et procedent qui bona fecerunt in resurrectionem vitae qui vero mala egerunt in resurrectionem iudicii
JOHN|5|30|non possum ego a me ipso facere quicquam sicut audio iudico et iudicium meum iustum est quia non quaero voluntatem meam sed voluntatem eius qui misit me
JOHN|5|31|si ego testimonium perhibeo de me testimonium meum non est verum
JOHN|5|32|alius est qui testimonium perhibet de me et scio quia verum est testimonium quod perhibet de me
JOHN|5|33|vos misistis ad Iohannem et testimonium perhibuit veritati
JOHN|5|34|ego autem non ab homine testimonium accipio sed haec dico ut vos salvi sitis
JOHN|5|35|ille erat lucerna ardens et lucens vos autem voluistis exultare ad horam in luce eius
JOHN|5|36|ego autem habeo testimonium maius Iohanne opera enim quae dedit mihi Pater ut perficiam ea ipsa opera quae ego facio testimonium perhibent de me quia Pater me misit
JOHN|5|37|et qui misit me Pater ipse testimonium perhibuit de me neque vocem eius umquam audistis neque speciem eius vidistis
JOHN|5|38|et verbum eius non habetis in vobis manens quia quem misit ille huic vos non creditis
JOHN|5|39|scrutamini scripturas quia vos putatis in ipsis vitam aeternam habere et illae sunt quae testimonium perhibent de me
JOHN|5|40|et non vultis venire ad me ut vitam habeatis
JOHN|5|41|claritatem ab hominibus non accipio
JOHN|5|42|sed cognovi vos quia dilectionem Dei non habetis in vobis
JOHN|5|43|ego veni in nomine Patris mei et non accipitis me si alius venerit in nomine suo illum accipietis
JOHN|5|44|quomodo potestis vos credere qui gloriam ab invicem accipitis et gloriam quae a solo est Deo non quaeritis
JOHN|5|45|nolite putare quia ego accusaturus sim vos apud Patrem est qui accuset vos Moses in quo vos speratis
JOHN|5|46|si enim crederetis Mosi crederetis forsitan et mihi de me enim ille scripsit
JOHN|5|47|si autem illius litteris non creditis quomodo meis verbis credetis
JOHN|6|1|post haec abiit Iesus trans mare Galilaeae quod est Tiberiadis
JOHN|6|2|et sequebatur eum multitudo magna quia videbant signa quae faciebat super his qui infirmabantur
JOHN|6|3|subiit ergo in montem Iesus et ibi sedebat cum discipulis suis
JOHN|6|4|erat autem proximum pascha dies festus Iudaeorum
JOHN|6|5|cum sublevasset ergo oculos Iesus et vidisset quia multitudo maxima venit ad eum dicit ad Philippum unde ememus panes ut manducent hii
JOHN|6|6|hoc autem dicebat temptans eum ipse enim sciebat quid esset facturus
JOHN|6|7|respondit ei Philippus ducentorum denariorum panes non sufficiunt eis ut unusquisque modicum quid accipiat
JOHN|6|8|dicit ei unus ex discipulis eius Andreas frater Simonis Petri
JOHN|6|9|est puer unus hic qui habet quinque panes hordiacios et duos pisces sed haec quid sunt inter tantos
JOHN|6|10|dixit ergo Iesus facite homines discumbere erat autem faenum multum in loco discubuerunt ergo viri numero quasi quinque milia
JOHN|6|11|accepit ergo panes Iesus et cum gratias egisset distribuit discumbentibus similiter et ex piscibus quantum volebant
JOHN|6|12|ut autem impleti sunt dixit discipulis suis colligite quae superaverunt fragmenta ne pereant
JOHN|6|13|collegerunt ergo et impleverunt duodecim cofinos fragmentorum ex quinque panibus hordiaciis quae superfuerunt his qui manducaverunt
JOHN|6|14|illi ergo homines cum vidissent quod fecerat signum dicebant quia hic est vere propheta qui venturus est in mundum
JOHN|6|15|Iesus ergo cum cognovisset quia venturi essent ut raperent eum et facerent eum regem fugit iterum in montem ipse solus
JOHN|6|16|ut autem sero factum est descenderunt discipuli eius ad mare
JOHN|6|17|et cum ascendissent navem venerunt trans mare in Capharnaum et tenebrae iam factae erant et non venerat ad eos Iesus
JOHN|6|18|mare autem vento magno flante exsurgebat
JOHN|6|19|cum remigassent ergo quasi stadia viginti quinque aut triginta vident Iesum ambulantem super mare et proximum navi fieri et timuerunt
JOHN|6|20|ille autem dicit eis ego sum nolite timere
JOHN|6|21|voluerunt ergo accipere eum in navi et statim fuit navis ad terram quam ibant
JOHN|6|22|altera die turba quae stabat trans mare vidit quia navicula alia non erat ibi nisi una et quia non introisset cum discipulis suis Iesus in navem sed soli discipuli eius abissent
JOHN|6|23|aliae vero supervenerunt naves a Tiberiade iuxta locum ubi manducaverant panem gratias agente Domino
JOHN|6|24|cum ergo vidisset turba quia Iesus non esset ibi neque discipuli eius ascenderunt naviculas et venerunt Capharnaum quaerentes Iesum
JOHN|6|25|et cum invenissent eum trans mare dixerunt ei rabbi quando huc venisti
JOHN|6|26|respondit eis Iesus et dixit amen amen dico vobis quaeritis me non quia vidistis signa sed quia manducastis ex panibus et saturati estis
JOHN|6|27|operamini non cibum qui perit sed qui permanet in vitam aeternam quem Filius hominis vobis dabit hunc enim Pater signavit Deus
JOHN|6|28|dixerunt ergo ad eum quid faciemus ut operemur opera Dei
JOHN|6|29|respondit Iesus et dixit eis hoc est opus Dei ut credatis in eum quem misit ille
JOHN|6|30|dixerunt ergo ei quod ergo tu facis signum ut videamus et credamus tibi quid operaris
JOHN|6|31|patres nostri manna manducaverunt in deserto sicut scriptum est panem de caelo dedit eis manducare
JOHN|6|32|dixit ergo eis Iesus amen amen dico vobis non Moses dedit vobis panem de caelo sed Pater meus dat vobis panem de caelo verum
JOHN|6|33|panis enim Dei est qui descendit de caelo et dat vitam mundo
JOHN|6|34|dixerunt ergo ad eum Domine semper da nobis panem hunc
JOHN|6|35|dixit autem eis Iesus ego sum panis vitae qui veniet ad me non esuriet et qui credit in me non sitiet umquam
JOHN|6|36|sed dixi vobis quia et vidistis me et non creditis
JOHN|6|37|omne quod dat mihi Pater ad me veniet et eum qui venit ad me non eiciam foras
JOHN|6|38|quia descendi de caelo non ut faciam voluntatem meam sed voluntatem eius qui misit me
JOHN|6|39|haec est autem voluntas eius qui misit me Patris ut omne quod dedit mihi non perdam ex eo sed resuscitem illum novissimo die
JOHN|6|40|haec est enim voluntas Patris mei qui misit me ut omnis qui videt Filium et credit in eum habeat vitam aeternam et resuscitabo ego eum in novissimo die
JOHN|6|41|murmurabant ergo Iudaei de illo quia dixisset ego sum panis qui de caelo descendi
JOHN|6|42|et dicebant nonne hic est Iesus filius Ioseph cuius nos novimus patrem et matrem quomodo ergo dicit hic quia de caelo descendi
JOHN|6|43|respondit ergo Iesus et dixit eis nolite murmurare in invicem
JOHN|6|44|nemo potest venire ad me nisi Pater qui misit me traxerit eum et ego resuscitabo eum novissimo die
JOHN|6|45|est scriptum in prophetis et erunt omnes docibiles Dei omnis qui audivit a Patre et didicit venit ad me
JOHN|6|46|non quia Patrem vidit quisquam nisi is qui est a Deo hic vidit Patrem
JOHN|6|47|amen amen dico vobis qui credit in me habet vitam aeternam
JOHN|6|48|ego sum panis vitae
JOHN|6|49|patres vestri manducaverunt in deserto manna et mortui sunt
JOHN|6|50|hic est panis de caelo descendens ut si quis ex ipso manducaverit non moriatur
JOHN|6|51|ego sum panis vivus qui de caelo descendi
JOHN|6|52|si quis manducaverit ex hoc pane vivet in aeternum et panis quem ego dabo caro mea est pro mundi vita
JOHN|6|53|litigabant ergo Iudaei ad invicem dicentes quomodo potest hic nobis carnem suam dare ad manducandum
JOHN|6|54|dixit ergo eis Iesus amen amen dico vobis nisi manducaveritis carnem Filii hominis et biberitis eius sanguinem non habetis vitam in vobis
JOHN|6|55|qui manducat meam carnem et bibit meum sanguinem habet vitam aeternam et ego resuscitabo eum in novissimo die
JOHN|6|56|caro enim mea vere est cibus et sanguis meus vere est potus
JOHN|6|57|qui manducat meam carnem et bibit meum sanguinem in me manet et ego in illo
JOHN|6|58|sicut misit me vivens Pater et ego vivo propter Patrem et qui manducat me et ipse vivet propter me
JOHN|6|59|hic est panis qui de caelo descendit non sicut manducaverunt patres vestri manna et mortui sunt qui manducat hunc panem vivet in aeternum
JOHN|6|60|haec dixit in synagoga docens in Capharnaum
JOHN|6|61|multi ergo audientes ex discipulis eius dixerunt durus est hic sermo quis potest eum audire
JOHN|6|62|sciens autem Iesus apud semet ipsum quia murmurarent de hoc discipuli eius dixit eis hoc vos scandalizat
JOHN|6|63|si ergo videritis Filium hominis ascendentem ubi erat prius
JOHN|6|64|spiritus est qui vivificat caro non prodest quicquam verba quae ego locutus sum vobis spiritus et vita sunt
JOHN|6|65|sed sunt quidam ex vobis qui non credunt sciebat enim ab initio Iesus qui essent credentes et quis traditurus esset eum
JOHN|6|66|et dicebat propterea dixi vobis quia nemo potest venire ad me nisi fuerit ei datum a Patre meo
JOHN|6|67|ex hoc multi discipulorum eius abierunt retro et iam non cum illo ambulabant
JOHN|6|68|dixit ergo Iesus ad duodecim numquid et vos vultis abire
JOHN|6|69|respondit ergo ei Simon Petrus Domine ad quem ibimus verba vitae aeternae habes
JOHN|6|70|et nos credidimus et cognovimus quia tu es Christus Filius Dei
JOHN|6|71|respondit eis Iesus nonne ego vos duodecim elegi et ex vobis unus diabolus est
JOHN|6|72|dicebat autem Iudam Simonis Scariotis hic enim erat traditurus eum cum esset unus ex duodecim
JOHN|7|1|post haec ambulabat Iesus in Galilaeam non enim volebat in Iudaeam ambulare quia quaerebant eum Iudaei interficere
JOHN|7|2|erat autem in proximo dies festus Iudaeorum scenopegia
JOHN|7|3|dixerunt autem ad eum fratres eius transi hinc et vade in Iudaeam ut et discipuli tui videant opera tua quae facis
JOHN|7|4|nemo quippe in occulto quid facit et quaerit ipse in palam esse si haec facis manifesta te ipsum mundo
JOHN|7|5|neque enim fratres eius credebant in eum
JOHN|7|6|dicit ergo eis Iesus tempus meum nondum advenit tempus autem vestrum semper est paratum
JOHN|7|7|non potest mundus odisse vos me autem odit quia ego testimonium perhibeo de illo quia opera eius mala sunt
JOHN|7|8|vos ascendite ad diem festum hunc ego non ascendo ad diem festum istum quia meum tempus nondum impletum est
JOHN|7|9|haec cum dixisset ipse mansit in Galilaea
JOHN|7|10|ut autem ascenderunt fratres eius tunc et ipse ascendit ad diem festum non manifeste sed quasi in occulto
JOHN|7|11|Iudaei ergo quaerebant eum in die festo et dicebant ubi est ille
JOHN|7|12|et murmur multus de eo erat in turba; quidam enim dicebant quia bonus est alii autem dicebant non sed seducit turbas
JOHN|7|13|nemo tamen palam loquebatur de illo propter metum Iudaeorum
JOHN|7|14|iam autem die festo mediante ascendit Iesus in templum et docebat
JOHN|7|15|et mirabantur Iudaei dicentes quomodo hic litteras scit cum non didicerit
JOHN|7|16|respondit eis Iesus et dixit mea doctrina non est mea sed eius qui misit me
JOHN|7|17|si quis voluerit voluntatem eius facere cognoscet de doctrina utrum ex Deo sit an ego a me ipso loquar
JOHN|7|18|qui a semet ipso loquitur gloriam propriam quaerit qui autem quaerit gloriam eius qui misit illum hic verax est et iniustitia in illo non est
JOHN|7|19|nonne Moses dedit vobis legem et nemo ex vobis facit legem
JOHN|7|20|quid me quaeritis interficere respondit turba et dixit daemonium habes quis te quaerit interficere
JOHN|7|21|respondit Iesus et dixit eis unum opus feci et omnes miramini
JOHN|7|22|propterea Moses dedit vobis circumcisionem non quia ex Mose est sed ex patribus et in sabbato circumciditis hominem
JOHN|7|23|si circumcisionem accipit homo in sabbato ut non solvatur lex Mosi mihi indignamini quia totum hominem sanum feci in sabbato
JOHN|7|24|nolite iudicare secundum faciem sed iustum iudicium iudicate
JOHN|7|25|dicebant ergo quidam ex Hierosolymis nonne hic est quem quaerunt interficere
JOHN|7|26|et ecce palam loquitur et nihil ei dicunt numquid vere cognoverunt principes quia hic est Christus
JOHN|7|27|sed hunc scimus unde sit Christus autem cum venerit nemo scit unde sit
JOHN|7|28|clamabat ergo docens in templo Iesus et dicens et me scitis et unde sim scitis et a me ipso non veni sed est verus qui misit me quem vos non scitis
JOHN|7|29|ego scio eum quia ab ipso sum et ipse me misit
JOHN|7|30|quaerebant ergo eum adprehendere et nemo misit in illum manus quia nondum venerat hora eius
JOHN|7|31|de turba autem multi crediderunt in eum et dicebant Christus cum venerit numquid plura signa faciet quam quae hic facit
JOHN|7|32|audierunt Pharisaei turbam murmurantem de illo haec et miserunt principes et Pharisaei ministros ut adprehenderent eum
JOHN|7|33|dixit ergo Iesus adhuc modicum tempus vobiscum sum et vado ad eum qui misit me
JOHN|7|34|quaeretis me et non invenietis et ubi sum ego vos non potestis venire
JOHN|7|35|dixerunt ergo Iudaei ad se ipsos quo hic iturus est quia non inveniemus eum numquid in dispersionem gentium iturus est et docturus gentes
JOHN|7|36|quis est hic sermo quem dixit quaeretis me et non invenietis et ubi sum ego non potestis venire
JOHN|7|37|in novissimo autem die magno festivitatis stabat Iesus et clamabat dicens si quis sitit veniat ad me et bibat
JOHN|7|38|qui credit in me sicut dixit scriptura flumina de ventre eius fluent aquae vivae
JOHN|7|39|hoc autem dixit de Spiritu quem accepturi erant credentes in eum non enim erat Spiritus quia Iesus nondum fuerat glorificatus
JOHN|7|40|ex illa ergo turba cum audissent hos sermones eius dicebant hic est vere propheta
JOHN|7|41|alii dicebant hic est Christus quidam autem dicebant numquid a Galilaea Christus venit
JOHN|7|42|nonne scriptura dicit quia ex semine David et Bethleem castello ubi erat David venit Christus
JOHN|7|43|dissensio itaque facta est in turba propter eum
JOHN|7|44|quidam autem ex ipsis volebant adprehendere eum sed nemo misit super illum manus
JOHN|7|45|venerunt ergo ministri ad pontifices et Pharisaeos et dixerunt eis illi quare non adduxistis eum
JOHN|7|46|responderunt ministri numquam sic locutus est homo sicut hic homo
JOHN|7|47|responderunt ergo eis Pharisaei numquid et vos seducti estis
JOHN|7|48|numquid aliquis ex principibus credidit in eum aut ex Pharisaeis
JOHN|7|49|sed turba haec quae non novit legem maledicti sunt
JOHN|7|50|dicit Nicodemus ad eos ille qui venit ad eum nocte qui unus erat ex ipsis
JOHN|7|51|numquid lex nostra iudicat hominem nisi audierit ab ipso prius et cognoverit quid faciat
JOHN|7|52|responderunt et dixerunt ei numquid et tu Galilaeus es scrutare et vide quia propheta a Galilaea non surgit
JOHN|7|53|et reversi sunt unusquisque in domum suam
JOHN|8|1|Iesus autem perrexit in montem Oliveti
JOHN|8|2|et diluculo iterum venit in templum et omnis populus venit ad eum et sedens docebat eos
JOHN|8|3|adducunt autem scribae et Pharisaei mulierem in adulterio deprehensam et statuerunt eam in medio
JOHN|8|4|et dixerunt ei magister haec mulier modo deprehensa est in adulterio
JOHN|8|5|in lege autem Moses mandavit nobis huiusmodi lapidare tu ergo quid dicis
JOHN|8|6|haec autem dicebant temptantes eum ut possent accusare eum Iesus autem inclinans se deorsum digito scribebat in terra
JOHN|8|7|cum autem perseverarent interrogantes eum erexit se et dixit eis qui sine peccato est vestrum primus in illam lapidem mittat
JOHN|8|8|et iterum se inclinans scribebat in terra
JOHN|8|9|audientes autem unus post unum exiebant incipientes a senioribus et remansit solus et mulier in medio stans
JOHN|8|10|erigens autem se Iesus dixit ei mulier ubi sunt nemo te condemnavit
JOHN|8|11|quae dixit nemo Domine dixit autem Iesus nec ego te condemnabo vade et amplius iam noli peccare
JOHN|8|12|iterum ergo locutus est eis Iesus dicens ego sum lux mundi qui sequitur me non ambulabit in tenebris sed habebit lucem vitae
JOHN|8|13|dixerunt ergo ei Pharisaei tu de te ipso testimonium perhibes testimonium tuum non est verum
JOHN|8|14|respondit Iesus et dixit eis et si ego testimonium perhibeo de me ipso verum est testimonium meum quia scio unde veni et quo vado vos autem nescitis unde venio aut quo vado
JOHN|8|15|vos secundum carnem iudicatis ego non iudico quemquam
JOHN|8|16|et si iudico ego iudicium meum verum est quia solus non sum sed ego et qui me misit Pater
JOHN|8|17|et in lege vestra scriptum est quia duorum hominum testimonium verum est
JOHN|8|18|ego sum qui testimonium perhibeo de me ipso et testimonium perhibet de me qui misit me Pater
JOHN|8|19|dicebant ergo ei ubi est Pater tuus respondit Iesus neque me scitis neque Patrem meum si me sciretis forsitan et Patrem meum sciretis
JOHN|8|20|haec verba locutus est in gazofilacio docens in templo et nemo adprehendit eum quia necdum venerat hora eius
JOHN|8|21|dixit ergo iterum eis Iesus ego vado et quaeretis me et in peccato vestro moriemini quo ego vado vos non potestis venire
JOHN|8|22|dicebant ergo Iudaei numquid interficiet semet ipsum quia dicit quo ego vado vos non potestis venire
JOHN|8|23|et dicebat eis vos de deorsum estis ego de supernis sum vos de mundo hoc estis ego non sum de hoc mundo
JOHN|8|24|dixi ergo vobis quia moriemini in peccatis vestris si enim non credideritis quia ego sum moriemini in peccato vestro
JOHN|8|25|dicebant ergo ei tu quis es dixit eis Iesus principium quia et loquor vobis
JOHN|8|26|multa habeo de vobis loqui et iudicare sed qui misit me verax est et ego quae audivi ab eo haec loquor in mundo
JOHN|8|27|et non cognoverunt quia Patrem eis dicebat
JOHN|8|28|dixit ergo eis Iesus cum exaltaveritis Filium hominis tunc cognoscetis quia ego sum et a me ipso facio nihil sed sicut docuit me Pater haec loquor
JOHN|8|29|et qui me misit mecum est non reliquit me solum quia ego quae placita sunt ei facio semper
JOHN|8|30|haec illo loquente multi crediderunt in eum
JOHN|8|31|dicebat ergo Iesus ad eos qui crediderunt ei Iudaeos si vos manseritis in sermone meo vere discipuli mei eritis
JOHN|8|32|et cognoscetis veritatem et veritas liberabit vos
JOHN|8|33|responderunt ei semen Abrahae sumus et nemini servivimus umquam quomodo tu dicis liberi eritis
JOHN|8|34|respondit eis Iesus amen amen dico vobis quia omnis qui facit peccatum servus est peccati
JOHN|8|35|servus autem non manet in domo in aeternum filius manet in aeternum
JOHN|8|36|si ergo Filius vos liberaverit vere liberi eritis
JOHN|8|37|scio quia filii Abrahae estis sed quaeritis me interficere quia sermo meus non capit in vobis
JOHN|8|38|ego quod vidi apud Patrem loquor et vos quae vidistis apud patrem vestrum facitis
JOHN|8|39|responderunt et dixerunt ei pater noster Abraham est dicit eis Iesus si filii Abrahae estis opera Abrahae facite
JOHN|8|40|nunc autem quaeritis me interficere hominem qui veritatem vobis locutus sum quam audivi a Deo hoc Abraham non fecit
JOHN|8|41|vos facitis opera patris vestri dixerunt itaque ei nos ex fornicatione non sumus nati unum patrem habemus Deum
JOHN|8|42|dixit ergo eis Iesus si Deus pater vester esset diligeretis utique me ego enim ex Deo processi et veni neque enim a me ipso veni sed ille me misit
JOHN|8|43|quare loquellam meam non cognoscitis quia non potestis audire sermonem meum
JOHN|8|44|vos ex patre diabolo estis et desideria patris vestri vultis facere ille homicida erat ab initio et in veritate non stetit quia non est veritas in eo cum loquitur mendacium ex propriis loquitur quia mendax est et pater eius
JOHN|8|45|ego autem quia veritatem dico non creditis mihi
JOHN|8|46|quis ex vobis arguit me de peccato si veritatem dico quare vos non creditis mihi
JOHN|8|47|qui est ex Deo verba Dei audit propterea vos non auditis quia ex Deo non estis
JOHN|8|48|responderunt igitur Iudaei et dixerunt ei nonne bene dicimus nos quia Samaritanus es tu et daemonium habes
JOHN|8|49|respondit Iesus ego daemonium non habeo sed honorifico Patrem meum et vos inhonoratis me
JOHN|8|50|ego autem non quaero gloriam meam est qui quaerit et iudicat
JOHN|8|51|amen amen dico vobis si quis sermonem meum servaverit mortem non videbit in aeternum
JOHN|8|52|dixerunt ergo Iudaei nunc cognovimus quia daemonium habes Abraham mortuus est et prophetae et tu dicis si quis sermonem meum servaverit non gustabit mortem in aeternum
JOHN|8|53|numquid tu maior es patre nostro Abraham qui mortuus est et prophetae mortui sunt quem te ipsum facis
JOHN|8|54|respondit Iesus si ego glorifico me ipsum gloria mea nihil est est Pater meus qui glorificat me quem vos dicitis quia Deus noster est
JOHN|8|55|et non cognovistis eum ego autem novi eum et si dixero quia non scio eum ero similis vobis mendax sed scio eum et sermonem eius servo
JOHN|8|56|Abraham pater vester exultavit ut videret diem meum et vidit et gavisus est
JOHN|8|57|dixerunt ergo Iudaei ad eum quinquaginta annos nondum habes et Abraham vidisti
JOHN|8|58|dixit eis Iesus amen amen dico vobis antequam Abraham fieret ego sum
JOHN|8|59|tulerunt ergo lapides ut iacerent in eum Iesus autem abscondit se et exivit de templo
JOHN|9|1|et praeteriens vidit hominem caecum a nativitate
JOHN|9|2|et interrogaverunt eum discipuli sui rabbi quis peccavit hic aut parentes eius ut caecus nasceretur
JOHN|9|3|respondit Iesus neque hic peccavit neque parentes eius sed ut manifestetur opera Dei in illo
JOHN|9|4|me oportet operari opera eius qui misit me donec dies est venit nox quando nemo potest operari
JOHN|9|5|quamdiu in mundo sum lux sum mundi
JOHN|9|6|haec cum dixisset expuit in terram et fecit lutum ex sputo et linuit lutum super oculos eius
JOHN|9|7|et dixit ei vade lava in natatoria Siloae quod interpretatur Missus abiit ergo et lavit et venit videns
JOHN|9|8|itaque vicini et qui videbant eum prius quia mendicus erat dicebant nonne hic est qui sedebat et mendicabat alii dicebant quia hic est
JOHN|9|9|alii autem nequaquam sed similis est eius ille dicebat quia ego sum
JOHN|9|10|dicebant ergo ei quomodo aperti sunt oculi tibi
JOHN|9|11|respondit ille homo qui dicitur Iesus lutum fecit et unxit oculos meos et dixit mihi vade ad natatoriam Siloae et lava et abii et lavi et vidi
JOHN|9|12|dixerunt ei ubi est ille ait nescio
JOHN|9|13|adducunt eum ad Pharisaeos qui caecus fuerat
JOHN|9|14|erat autem sabbatum quando lutum fecit Iesus et aperuit oculos eius
JOHN|9|15|iterum ergo interrogabant eum Pharisaei quomodo vidisset ille autem dixit eis lutum posuit mihi super oculos et lavi et video
JOHN|9|16|dicebant ergo ex Pharisaeis quidam non est hic homo a Deo quia sabbatum non custodit alii dicebant quomodo potest homo peccator haec signa facere et scisma erat in eis
JOHN|9|17|dicunt ergo caeco iterum tu quid dicis de eo qui aperuit oculos tuos ille autem dixit quia propheta est
JOHN|9|18|non crediderunt ergo Iudaei de illo quia caecus fuisset et vidisset donec vocaverunt parentes eius qui viderat
JOHN|9|19|et interrogaverunt eos dicentes hic est filius vester quem vos dicitis quia caecus natus est quomodo ergo nunc videt
JOHN|9|20|responderunt eis parentes eius et dixerunt scimus quia hic est filius noster et quia caecus natus est
JOHN|9|21|quomodo autem nunc videat nescimus aut quis eius aperuit oculos nos nescimus ipsum interrogate aetatem habet ipse de se loquatur
JOHN|9|22|haec dixerunt parentes eius quia timebant Iudaeos iam enim conspiraverant Iudaei ut si quis eum confiteretur Christum extra synagogam fieret
JOHN|9|23|propterea parentes eius dixerunt quia aetatem habet ipsum interrogate
JOHN|9|24|vocaverunt ergo rursum hominem qui fuerat caecus et dixerunt ei da gloriam Deo nos scimus quia hic homo peccator est
JOHN|9|25|dixit ergo ille si peccator est nescio unum scio quia caecus cum essem modo video
JOHN|9|26|dixerunt ergo illi quid fecit tibi quomodo aperuit tibi oculos
JOHN|9|27|respondit eis dixi vobis iam et audistis quid iterum vultis audire numquid et vos vultis discipuli eius fieri
JOHN|9|28|maledixerunt ei et dixerunt tu discipulus illius es nos autem Mosi discipuli sumus
JOHN|9|29|nos scimus quia Mosi locutus est Deus hunc autem nescimus unde sit
JOHN|9|30|respondit ille homo et dixit eis in hoc enim mirabile est quia vos nescitis unde sit et aperuit meos oculos
JOHN|9|31|scimus autem quia peccatores Deus non audit sed si quis Dei cultor est et voluntatem eius facit hunc exaudit
JOHN|9|32|a saeculo non est auditum quia aperuit quis oculos caeci nati
JOHN|9|33|nisi esset hic a Deo non poterat facere quicquam
JOHN|9|34|responderunt et dixerunt ei in peccatis natus es totus et tu doces nos et eiecerunt eum foras
JOHN|9|35|audivit Iesus quia eiecerunt eum foras et cum invenisset eum dixit ei tu credis in Filium Dei
JOHN|9|36|respondit ille et dixit quis est Domine ut credam in eum
JOHN|9|37|et dixit ei Iesus et vidisti eum et qui loquitur tecum ipse est
JOHN|9|38|at ille ait credo Domine et procidens adoravit eum
JOHN|9|39|dixit ei Iesus in iudicium ego in hunc mundum veni ut qui non vident videant et qui vident caeci fiant
JOHN|9|40|et audierunt ex Pharisaeis qui cum ipso erant et dixerunt ei numquid et nos caeci sumus
JOHN|9|41|dixit eis Iesus si caeci essetis non haberetis peccatum nunc vero dicitis quia videmus peccatum vestrum manet
JOHN|10|1|amen amen dico vobis qui non intrat per ostium in ovile ovium sed ascendit aliunde ille fur est et latro
JOHN|10|2|qui autem intrat per ostium pastor est ovium
JOHN|10|3|huic ostiarius aperit et oves vocem eius audiunt et proprias oves vocat nominatim et educit eas
JOHN|10|4|et cum proprias oves emiserit ante eas vadit et oves illum sequuntur quia sciunt vocem eius
JOHN|10|5|alienum autem non sequuntur sed fugient ab eo quia non noverunt vocem alienorum
JOHN|10|6|hoc proverbium dixit eis Iesus illi autem non cognoverunt quid loqueretur eis
JOHN|10|7|dixit ergo eis iterum Iesus amen amen dico vobis quia ego sum ostium ovium
JOHN|10|8|omnes quotquot venerunt fures sunt et latrones sed non audierunt eos oves
JOHN|10|9|ego sum ostium per me si quis introierit salvabitur et ingredietur et egredietur et pascua inveniet
JOHN|10|10|fur non venit nisi ut furetur et mactet et perdat ego veni ut vitam habeant et abundantius habeant
JOHN|10|11|ego sum pastor bonus bonus pastor animam suam dat pro ovibus
JOHN|10|12|mercennarius et qui non est pastor cuius non sunt oves propriae videt lupum venientem et dimittit oves et fugit et lupus rapit et dispergit oves
JOHN|10|13|mercennarius autem fugit quia mercennarius est et non pertinet ad eum de ovibus
JOHN|10|14|ego sum pastor bonus et cognosco meas et cognoscunt me meae
JOHN|10|15|sicut novit me Pater et ego agnosco Patrem et animam meam pono pro ovibus
JOHN|10|16|et alias oves habeo quae non sunt ex hoc ovili et illas oportet me adducere et vocem meam audient et fiet unum ovile unus pastor
JOHN|10|17|propterea me Pater diligit quia ego pono animam meam ut iterum sumam eam
JOHN|10|18|nemo tollit eam a me sed ego pono eam a me ipso potestatem habeo ponendi eam et potestatem habeo iterum sumendi eam hoc mandatum accepi a Patre meo
JOHN|10|19|dissensio iterum facta est inter Iudaeos propter sermones hos
JOHN|10|20|dicebant autem multi ex ipsis daemonium habet et insanit quid eum auditis
JOHN|10|21|alii dicebant haec verba non sunt daemonium habentis numquid daemonium potest caecorum oculos aperire
JOHN|10|22|facta sunt autem encenia in Hierosolymis et hiemps erat
JOHN|10|23|et ambulabat Iesus in templo in porticu Salomonis
JOHN|10|24|circumdederunt ergo eum Iudaei et dicebant ei quousque animam nostram tollis si tu es Christus dic nobis palam
JOHN|10|25|respondit eis Iesus loquor vobis et non creditis opera quae ego facio in nomine Patris mei haec testimonium perhibent de me
JOHN|10|26|sed vos non creditis quia non estis ex ovibus meis
JOHN|10|27|oves meae vocem meam audiunt et ego cognosco eas et sequuntur me
JOHN|10|28|et ego vitam aeternam do eis et non peribunt in aeternum et non rapiet eas quisquam de manu mea
JOHN|10|29|Pater meus quod dedit mihi maius omnibus est et nemo potest rapere de manu Patris mei
JOHN|10|30|ego et Pater unum sumus
JOHN|10|31|sustulerunt lapides Iudaei ut lapidarent eum
JOHN|10|32|respondit eis Iesus multa opera bona ostendi vobis ex Patre meo propter quod eorum opus me lapidatis
JOHN|10|33|responderunt ei Iudaei de bono opere non lapidamus te sed de blasphemia et quia tu homo cum sis facis te ipsum Deum
JOHN|10|34|respondit eis Iesus nonne scriptum est in lege vestra quia ego dixi dii estis
JOHN|10|35|si illos dixit deos ad quos sermo Dei factus est et non potest solvi scriptura
JOHN|10|36|quem Pater sanctificavit et misit in mundum vos dicitis quia blasphemas quia dixi Filius Dei sum
JOHN|10|37|si non facio opera Patris mei nolite credere mihi
JOHN|10|38|si autem facio et si mihi non vultis credere operibus credite ut cognoscatis et credatis quia in me est Pater et ego in Patre
JOHN|10|39|quaerebant ergo eum prendere et exivit de manibus eorum
JOHN|10|40|et abiit iterum trans Iordanen in eum locum ubi erat Iohannes baptizans primum et mansit illic
JOHN|10|41|et multi venerunt ad eum et dicebant quia Iohannes quidem signum fecit nullum
JOHN|10|42|omnia autem quaecumque dixit Iohannes de hoc vera erant et multi crediderunt in eum
JOHN|11|1|erat autem quidam languens Lazarus a Bethania de castello Mariae et Marthae sororis eius
JOHN|11|2|Maria autem erat quae unxit Dominum unguento et extersit pedes eius capillis suis cuius frater Lazarus infirmabatur
JOHN|11|3|miserunt ergo sorores ad eum dicentes Domine ecce quem amas infirmatur
JOHN|11|4|audiens autem Iesus dixit eis infirmitas haec non est ad mortem sed pro gloria Dei ut glorificetur Filius Dei per eam
JOHN|11|5|diligebat autem Iesus Martham et sororem eius Mariam et Lazarum
JOHN|11|6|ut ergo audivit quia infirmabatur tunc quidem mansit in eodem loco duobus diebus
JOHN|11|7|deinde post haec dicit discipulis suis eamus in Iudaeam iterum
JOHN|11|8|dicunt ei discipuli rabbi nunc quaerebant te Iudaei lapidare et iterum vadis illuc
JOHN|11|9|respondit Iesus nonne duodecim horae sunt diei si quis ambulaverit in die non offendit quia lucem huius mundi videt
JOHN|11|10|si autem ambulaverit nocte offendit quia lux non est in eo
JOHN|11|11|haec ait et post hoc dicit eis Lazarus amicus noster dormit sed vado ut a somno exsuscitem eum
JOHN|11|12|dixerunt ergo discipuli eius Domine si dormit salvus erit
JOHN|11|13|dixerat autem Iesus de morte eius illi autem putaverunt quia de dormitione somni diceret
JOHN|11|14|tunc ergo dixit eis Iesus manifeste Lazarus mortuus est
JOHN|11|15|et gaudeo propter vos ut credatis quoniam non eram ibi sed eamus ad eum
JOHN|11|16|dixit ergo Thomas qui dicitur Didymus ad condiscipulos eamus et nos ut moriamur cum eo
JOHN|11|17|venit itaque Iesus et invenit eum quattuor dies iam in monumento habentem
JOHN|11|18|erat autem Bethania iuxta Hierosolyma quasi stadiis quindecim
JOHN|11|19|multi autem ex Iudaeis venerant ad Martham et Mariam ut consolarentur eas de fratre suo
JOHN|11|20|Martha ergo ut audivit quia Iesus venit occurrit illi Maria autem domi sedebat
JOHN|11|21|dixit ergo Martha ad Iesum Domine si fuisses hic frater meus non fuisset mortuus
JOHN|11|22|sed et nunc scio quia quaecumque poposceris a Deo dabit tibi Deus
JOHN|11|23|dicit illi Iesus resurget frater tuus
JOHN|11|24|dicit ei Martha scio quia resurget in resurrectione in novissima die
JOHN|11|25|dixit ei Iesus ego sum resurrectio et vita qui credit in me et si mortuus fuerit vivet
JOHN|11|26|et omnis qui vivit et credit in me non morietur in aeternum credis hoc
JOHN|11|27|ait illi utique Domine ego credidi quia tu es Christus Filius Dei qui in mundum venisti
JOHN|11|28|et cum haec dixisset abiit et vocavit Mariam sororem suam silentio dicens magister adest et vocat te
JOHN|11|29|illa ut audivit surgit cito et venit ad eum
JOHN|11|30|nondum enim venerat Iesus in castellum sed erat adhuc in illo loco ubi occurrerat ei Martha
JOHN|11|31|Iudaei igitur qui erant cum ea in domo et consolabantur eam cum vidissent Mariam quia cito surrexit et exiit secuti sunt eam dicentes quia vadit ad monumentum ut ploret ibi
JOHN|11|32|Maria ergo cum venisset ubi erat Iesus videns eum cecidit ad pedes eius et dixit ei Domine si fuisses hic non esset mortuus frater meus
JOHN|11|33|Iesus ergo ut vidit eam plorantem et Iudaeos qui venerant cum ea plorantes fremuit spiritu et turbavit se ipsum
JOHN|11|34|et dixit ubi posuistis eum dicunt ei Domine veni et vide
JOHN|11|35|et lacrimatus est Iesus
JOHN|11|36|dixerunt ergo Iudaei ecce quomodo amabat eum
JOHN|11|37|quidam autem dixerunt ex ipsis non poterat hic qui aperuit oculos caeci facere ut et hic non moreretur
JOHN|11|38|Iesus ergo rursum fremens in semet ipso venit ad monumentum erat autem spelunca et lapis superpositus erat ei
JOHN|11|39|ait Iesus tollite lapidem dicit ei Martha soror eius qui mortuus fuerat Domine iam fetet quadriduanus enim est
JOHN|11|40|dicit ei Iesus nonne dixi tibi quoniam si credideris videbis gloriam Dei
JOHN|11|41|tulerunt ergo lapidem Iesus autem elevatis sursum oculis dixit Pater gratias ago tibi quoniam audisti me
JOHN|11|42|ego autem sciebam quia semper me audis sed propter populum qui circumstat dixi ut credant quia tu me misisti
JOHN|11|43|haec cum dixisset voce magna clamavit Lazare veni foras
JOHN|11|44|et statim prodiit qui fuerat mortuus ligatus pedes et manus institis et facies illius sudario erat ligata dicit Iesus eis solvite eum et sinite abire
JOHN|11|45|multi ergo ex Iudaeis qui venerant ad Mariam et viderant quae fecit crediderunt in eum
JOHN|11|46|quidam autem ex ipsis abierunt ad Pharisaeos et dixerunt eis quae fecit Iesus
JOHN|11|47|collegerunt ergo pontifices et Pharisaei concilium et dicebant quid facimus quia hic homo multa signa facit
JOHN|11|48|si dimittimus eum sic omnes credent in eum et venient Romani et tollent nostrum et locum et gentem
JOHN|11|49|unus autem ex ipsis Caiaphas cum esset pontifex anni illius dixit eis vos nescitis quicquam
JOHN|11|50|nec cogitatis quia expedit nobis ut unus moriatur homo pro populo et non tota gens pereat
JOHN|11|51|hoc autem a semet ipso non dixit sed cum esset pontifex anni illius prophetavit quia Iesus moriturus erat pro gente
JOHN|11|52|et non tantum pro gente sed et ut filios Dei qui erant dispersi congregaret in unum
JOHN|11|53|ab illo ergo die cogitaverunt ut interficerent eum
JOHN|11|54|Iesus ergo iam non in palam ambulabat apud Iudaeos sed abiit in regionem iuxta desertum in civitatem quae dicitur Efrem et ibi morabatur cum discipulis
JOHN|11|55|proximum autem erat pascha Iudaeorum et ascenderunt multi Hierosolyma de regione ante pascha ut sanctificarent se ipsos
JOHN|11|56|quaerebant ergo Iesum et conloquebantur ad invicem in templo stantes quid putatis quia non veniat ad diem festum
JOHN|11|57|dederant autem pontifices et Pharisaei mandatum ut si quis cognoverit ubi sit indicet ut adprehendant eum
JOHN|12|1|Iesus ergo ante sex dies paschae venit Bethaniam ubi fuerat Lazarus mortuus quem suscitavit Iesus
JOHN|12|2|fecerunt autem ei cenam ibi et Martha ministrabat Lazarus vero unus erat ex discumbentibus cum eo
JOHN|12|3|Maria ergo accepit libram unguenti nardi pistici pretiosi unxit pedes Iesu et extersit capillis suis pedes eius et domus impleta est ex odore unguenti
JOHN|12|4|dicit ergo unus ex discipulis eius Iudas Scariotis qui erat eum traditurus
JOHN|12|5|quare hoc unguentum non veniit trecentis denariis et datum est egenis
JOHN|12|6|dixit autem hoc non quia de egenis pertinebat ad eum sed quia fur erat et loculos habens ea quae mittebantur portabat
JOHN|12|7|dixit ergo Iesus sine illam ut in die sepulturae meae servet illud
JOHN|12|8|pauperes enim semper habetis vobiscum me autem non semper habetis
JOHN|12|9|cognovit ergo turba multa ex Iudaeis quia illic est et venerunt non propter Iesum tantum sed ut Lazarum viderent quem suscitavit a mortuis
JOHN|12|10|cogitaverunt autem principes sacerdotum ut et Lazarum interficerent
JOHN|12|11|quia multi propter illum abibant ex Iudaeis et credebant in Iesum
JOHN|12|12|in crastinum autem turba multa quae venerat ad diem festum cum audissent quia venit Iesus Hierosolyma
JOHN|12|13|acceperunt ramos palmarum et processerunt obviam ei et clamabant osanna benedictus qui venit in nomine Domini rex Israhel
JOHN|12|14|et invenit Iesus asellum et sedit super eum sicut scriptum est
JOHN|12|15|noli timere filia Sion ecce rex tuus venit sedens super pullum asinae
JOHN|12|16|haec non cognoverunt discipuli eius primum sed quando glorificatus est Iesus tunc recordati sunt quia haec erant scripta de eo et haec fecerunt ei
JOHN|12|17|testimonium ergo perhibebat turba quae erat cum eo quando Lazarum vocavit de monumento et suscitavit eum a mortuis
JOHN|12|18|propterea et obviam venit ei turba quia audierunt eum fecisse hoc signum
JOHN|12|19|Pharisaei ergo dixerunt ad semet ipsos videtis quia nihil proficimus ecce mundus totus post eum abiit
JOHN|12|20|erant autem gentiles quidam ex his qui ascenderant ut adorarent in die festo
JOHN|12|21|hii ergo accesserunt ad Philippum qui erat a Bethsaida Galilaeae et rogabant eum dicentes domine volumus Iesum videre
JOHN|12|22|venit Philippus et dicit Andreae Andreas rursum et Philippus dixerunt Iesu
JOHN|12|23|Iesus autem respondit eis dicens venit hora ut clarificetur Filius hominis
JOHN|12|24|amen amen dico vobis nisi granum frumenti cadens in terram mortuum fuerit
JOHN|12|25|ipsum solum manet si autem mortuum fuerit multum fructum adfert qui amat animam suam perdet eam et qui odit animam suam in hoc mundo in vitam aeternam custodit eam
JOHN|12|26|si quis mihi ministrat me sequatur et ubi sum ego illic et minister meus erit si quis mihi ministraverit honorificabit eum Pater meus
JOHN|12|27|nunc anima mea turbata est et quid dicam Pater salvifica me ex hora hac sed propterea veni in horam hanc
JOHN|12|28|Pater clarifica tuum nomen venit ergo vox de caelo et clarificavi et iterum clarificabo
JOHN|12|29|turba ergo quae stabat et audierat dicebant tonitruum factum esse alii dicebant angelus ei locutus est
JOHN|12|30|respondit Iesus et dixit non propter me vox haec venit sed propter vos
JOHN|12|31|nunc iudicium est mundi nunc princeps huius mundi eicietur foras
JOHN|12|32|et ego si exaltatus fuero a terra omnia traham ad me ipsum
JOHN|12|33|hoc autem dicebat significans qua morte esset moriturus
JOHN|12|34|respondit ei turba nos audivimus ex lege quia Christus manet in aeternum et quomodo tu dicis oportet exaltari Filium hominis quis est iste Filius hominis
JOHN|12|35|dixit ergo eis Iesus adhuc modicum lumen in vobis est ambulate dum lucem habetis ut non tenebrae vos conprehendant et qui ambulat in tenebris nescit quo vadat
JOHN|12|36|dum lucem habetis credite in lucem ut filii lucis sitis haec locutus est Iesus et abiit et abscondit se ab eis
JOHN|12|37|cum autem tanta signa fecisset coram eis non credebant in eum
JOHN|12|38|ut sermo Esaiae prophetae impleretur quem dixit Domine quis credidit auditui nostro et brachium Domini cui revelatum est
JOHN|12|39|propterea non poterant credere quia iterum dixit Esaias
JOHN|12|40|excaecavit oculos eorum et induravit eorum cor ut non videant oculis et intellegant corde et convertantur et sanem eos
JOHN|12|41|haec dixit Esaias quando vidit gloriam eius et locutus est de eo
JOHN|12|42|verumtamen et ex principibus multi crediderunt in eum sed propter Pharisaeos non confitebantur ut de synagoga non eicerentur
JOHN|12|43|dilexerunt enim gloriam hominum magis quam gloriam Dei
JOHN|12|44|Iesus autem clamavit et dixit qui credit in me non credit in me sed in eum qui misit me
JOHN|12|45|et qui videt me videt eum qui misit me
JOHN|12|46|ego lux in mundum veni ut omnis qui credit in me in tenebris non maneat
JOHN|12|47|et si quis audierit verba mea et non custodierit ego non iudico eum non enim veni ut iudicem mundum sed ut salvificem mundum
JOHN|12|48|qui spernit me et non accipit verba mea habet qui iudicet eum sermo quem locutus sum ille iudicabit eum in novissimo die
JOHN|12|49|quia ego ex me ipso non sum locutus sed qui misit me Pater ipse mihi mandatum dedit quid dicam et quid loquar
JOHN|12|50|et scio quia mandatum eius vita aeterna est quae ergo ego loquor sicut dixit mihi Pater sic loquor
JOHN|13|1|ante diem autem festum paschae sciens Iesus quia venit eius hora ut transeat ex hoc mundo ad Patrem cum dilexisset suos qui erant in mundo in finem dilexit eos
JOHN|13|2|et cena facta cum diabolus iam misisset in corde ut traderet eum Iudas Simonis Scariotis
JOHN|13|3|sciens quia omnia dedit ei Pater in manus et quia a Deo exivit et ad Deum vadit
JOHN|13|4|surgit a cena et ponit vestimenta sua et cum accepisset linteum praecinxit se
JOHN|13|5|deinde mittit aquam in pelvem et coepit lavare pedes discipulorum et extergere linteo quo erat praecinctus
JOHN|13|6|venit ergo ad Simonem Petrum et dicit ei Petrus Domine tu mihi lavas pedes
JOHN|13|7|respondit Iesus et dicit ei quod ego facio tu nescis modo scies autem postea
JOHN|13|8|dicit ei Petrus non lavabis mihi pedes in aeternum respondit Iesus ei si non lavero te non habes partem mecum
JOHN|13|9|dicit ei Simon Petrus Domine non tantum pedes meos sed et manus et caput
JOHN|13|10|dicit ei Iesus qui lotus est non indiget ut lavet sed est mundus totus et vos mundi estis sed non omnes
JOHN|13|11|sciebat enim quisnam esset qui traderet eum propterea dixit non estis mundi omnes
JOHN|13|12|postquam ergo lavit pedes eorum et accepit vestimenta sua cum recubuisset iterum dixit eis scitis quid fecerim vobis
JOHN|13|13|vos vocatis me magister et Domine et bene dicitis sum etenim
JOHN|13|14|si ergo ego lavi vestros pedes Dominus et magister et vos debetis alter alterius lavare pedes
JOHN|13|15|exemplum enim dedi vobis ut quemadmodum ego feci vobis ita et vos faciatis
JOHN|13|16|amen amen dico vobis non est servus maior domino suo neque apostolus maior eo qui misit illum
JOHN|13|17|si haec scitis beati eritis si feceritis ea
JOHN|13|18|non de omnibus vobis dico ego scio quos elegerim sed ut impleatur scriptura qui manducat mecum panem levavit contra me calcaneum suum
JOHN|13|19|amodo dico vobis priusquam fiat ut credatis cum factum fuerit quia ego sum
JOHN|13|20|amen amen dico vobis qui accipit si quem misero me accipit qui autem me accipit accipit eum qui me misit
JOHN|13|21|cum haec dixisset Iesus turbatus est spiritu et protestatus est et dixit amen amen dico vobis quia unus ex vobis tradet me
JOHN|13|22|aspiciebant ergo ad invicem discipuli haesitantes de quo diceret
JOHN|13|23|erat ergo recumbens unus ex discipulis eius in sinu Iesu quem diligebat Iesus
JOHN|13|24|innuit ergo huic Simon Petrus et dicit ei quis est de quo dicit
JOHN|13|25|itaque cum recubuisset ille supra pectus Iesu dicit ei Domine quis est
JOHN|13|26|respondit Iesus ille est cui ego intinctum panem porrexero et cum intinxisset panem dedit Iudae Simonis Scariotis
JOHN|13|27|et post buccellam tunc introivit in illum Satanas dicit ei Iesus quod facis fac citius
JOHN|13|28|hoc autem nemo scivit discumbentium ad quid dixerit ei
JOHN|13|29|quidam enim putabant quia loculos habebat Iudas quia dicit ei Iesus eme ea quae opus sunt nobis ad diem festum aut egenis ut aliquid daret
JOHN|13|30|cum ergo accepisset ille buccellam exivit continuo erat autem nox
JOHN|13|31|cum ergo exisset dicit Iesus nunc clarificatus est Filius hominis et Deus clarificatus est in eo
JOHN|13|32|si Deus clarificatus est in eo et Deus clarificabit eum in semet ipso et continuo clarificabit eum
JOHN|13|33|filioli adhuc modicum vobiscum sum quaeretis me et sicut dixi Iudaeis quo ego vado vos non potestis venire et vobis dico modo
JOHN|13|34|mandatum novum do vobis ut diligatis invicem sicut dilexi vos ut et vos diligatis invicem
JOHN|13|35|in hoc cognoscent omnes quia mei discipuli estis si dilectionem habueritis ad invicem
JOHN|13|36|dicit ei Simon Petrus Domine quo vadis respondit Iesus quo ego vado non potes me modo sequi sequeris autem postea
JOHN|13|37|dicit ei Petrus quare non possum sequi te modo animam meam pro te ponam
JOHN|13|38|respondit Iesus animam tuam pro me ponis amen amen dico tibi non cantabit gallus donec me ter neges
JOHN|14|1|non turbetur cor vestrum creditis in Deum et in me credite
JOHN|14|2|in domo Patris mei mansiones multae sunt si quo minus dixissem vobis quia vado parare vobis locum
JOHN|14|3|et si abiero et praeparavero vobis locum iterum venio et accipiam vos ad me ipsum ut ubi sum ego et vos sitis
JOHN|14|4|et quo ego vado scitis et viam scitis
JOHN|14|5|dicit ei Thomas Domine nescimus quo vadis et quomodo possumus viam scire
JOHN|14|6|dicit ei Iesus ego sum via et veritas et vita nemo venit ad Patrem nisi per me
JOHN|14|7|si cognovissetis me et Patrem meum utique cognovissetis et amodo cognoscitis eum et vidistis eum
JOHN|14|8|dicit ei Philippus Domine ostende nobis Patrem et sufficit nobis
JOHN|14|9|dicit ei Iesus tanto tempore vobiscum sum et non cognovistis me Philippe qui vidit me vidit et Patrem quomodo tu dicis ostende nobis Patrem
JOHN|14|10|non credis quia ego in Patre et Pater in me est verba quae ego loquor vobis a me ipso non loquor Pater autem in me manens ipse facit opera
JOHN|14|11|non creditis quia ego in Patre et Pater in me est
JOHN|14|12|alioquin propter opera ipsa credite amen amen dico vobis qui credit in me opera quae ego facio et ipse faciet et maiora horum faciet quia ego ad Patrem vado
JOHN|14|13|et quodcumque petieritis in nomine meo hoc faciam ut glorificetur Pater in Filio
JOHN|14|14|si quid petieritis me in nomine meo hoc faciam
JOHN|14|15|si diligitis me mandata mea servate
JOHN|14|16|et ego rogabo Patrem et alium paracletum dabit vobis ut maneat vobiscum in aeternum
JOHN|14|17|Spiritum veritatis quem mundus non potest accipere quia non videt eum nec scit eum vos autem cognoscitis eum quia apud vos manebit et in vobis erit
JOHN|14|18|non relinquam vos orfanos veniam ad vos
JOHN|14|19|adhuc modicum et mundus me iam non videt vos autem videtis me quia ego vivo et vos vivetis
JOHN|14|20|in illo die vos cognoscetis quia ego sum in Patre meo et vos in me et ego in vobis
JOHN|14|21|qui habet mandata mea et servat ea ille est qui diligit me qui autem diligit me diligetur a Patre meo et ego diligam eum et manifestabo ei me ipsum
JOHN|14|22|dicit ei Iudas non ille Scariotis Domine quid factum est quia nobis manifestaturus es te ipsum et non mundo
JOHN|14|23|respondit Iesus et dixit ei si quis diligit me sermonem meum servabit et Pater meus diliget eum et ad eum veniemus et mansiones apud eum faciemus
JOHN|14|24|qui non diligit me sermones meos non servat et sermonem quem audistis non est meus sed eius qui misit me Patris
JOHN|14|25|haec locutus sum vobis apud vos manens
JOHN|14|26|paracletus autem Spiritus Sanctus quem mittet Pater in nomine meo ille vos docebit omnia et suggeret vobis omnia quaecumque dixero vobis
JOHN|14|27|pacem relinquo vobis pacem meam do vobis non quomodo mundus dat ego do vobis non turbetur cor vestrum neque formidet
JOHN|14|28|audistis quia ego dixi vobis vado et venio ad vos si diligeretis me gauderetis utique quia vado ad Patrem quia Pater maior me est
JOHN|14|29|et nunc dixi vobis priusquam fiat ut cum factum fuerit credatis
JOHN|14|30|iam non multa loquar vobiscum venit enim princeps mundi huius et in me non habet quicquam
JOHN|14|31|sed ut cognoscat mundus quia diligo Patrem et sicut mandatum dedit mihi Pater sic facio surgite eamus hinc
JOHN|15|1|ego sum vitis vera et Pater meus agricola est
JOHN|15|2|omnem palmitem in me non ferentem fructum tollet eum et omnem qui fert fructum purgabit eum ut fructum plus adferat
JOHN|15|3|iam vos mundi estis propter sermonem quem locutus sum vobis
JOHN|15|4|manete in me et ego in vobis sicut palmes non potest ferre fructum a semet ipso nisi manserit in vite sic nec vos nisi in me manseritis
JOHN|15|5|ego sum vitis vos palmites qui manet in me et ego in eo hic fert fructum multum quia sine me nihil potestis facere
JOHN|15|6|si quis in me non manserit mittetur foras sicut palmes et aruit et colligent eos et in ignem mittunt et ardent
JOHN|15|7|si manseritis in me et verba mea in vobis manserint quodcumque volueritis petetis et fiet vobis
JOHN|15|8|in hoc clarificatus est Pater meus ut fructum plurimum adferatis et efficiamini mei discipuli
JOHN|15|9|sicut dilexit me Pater et ego dilexi vos manete in dilectione mea
JOHN|15|10|si praecepta mea servaveritis manebitis in dilectione mea sicut et ego Patris mei praecepta servavi et maneo in eius dilectione
JOHN|15|11|haec locutus sum vobis ut gaudium meum in vobis sit et gaudium vestrum impleatur
JOHN|15|12|hoc est praeceptum meum ut diligatis invicem sicut dilexi vos
JOHN|15|13|maiorem hac dilectionem nemo habet ut animam suam quis ponat pro amicis suis
JOHN|15|14|vos amici mei estis si feceritis quae ego praecipio vobis
JOHN|15|15|iam non dico vos servos quia servus nescit quid facit dominus eius vos autem dixi amicos quia omnia quaecumque audivi a Patre meo nota feci vobis
JOHN|15|16|non vos me elegistis sed ego elegi vos et posui vos ut eatis et fructum adferatis et fructus vester maneat ut quodcumque petieritis Patrem in nomine meo det vobis
JOHN|15|17|haec mando vobis ut diligatis invicem
JOHN|15|18|si mundus vos odit scitote quia me priorem vobis odio habuit
JOHN|15|19|si de mundo fuissetis mundus quod suum erat diligeret quia vero de mundo non estis sed ego elegi vos de mundo propterea odit vos mundus
JOHN|15|20|mementote sermonis mei quem ego dixi vobis non est servus maior domino suo si me persecuti sunt et vos persequentur si sermonem meum servaverunt et vestrum servabunt
JOHN|15|21|sed haec omnia facient vobis propter nomen meum quia nesciunt eum qui misit me
JOHN|15|22|si non venissem et locutus fuissem eis peccatum non haberent nunc autem excusationem non habent de peccato suo
JOHN|15|23|qui me odit et Patrem meum odit
JOHN|15|24|si opera non fecissem in eis quae nemo alius fecit peccatum non haberent nunc autem et viderunt et oderunt et me et Patrem meum
JOHN|15|25|sed ut impleatur sermo qui in lege eorum scriptus est quia odio me habuerunt gratis
JOHN|15|26|cum autem venerit paracletus quem ego mittam vobis a Patre Spiritum veritatis qui a Patre procedit ille testimonium perhibebit de me
JOHN|15|27|et vos testimonium perhibetis quia ab initio mecum estis
JOHN|16|1|haec locutus sum vobis ut non scandalizemini
JOHN|16|2|absque synagogis facient vos sed venit hora ut omnis qui interficit vos arbitretur obsequium se praestare Deo
JOHN|16|3|et haec facient quia non noverunt Patrem neque me
JOHN|16|4|sed haec locutus sum vobis ut cum venerit hora eorum reminiscamini quia ego dixi vobis
JOHN|16|5|haec autem vobis ab initio non dixi quia vobiscum eram at nunc vado ad eum qui me misit et nemo ex vobis interrogat me quo vadis
JOHN|16|6|sed quia haec locutus sum vobis tristitia implevit cor vestrum
JOHN|16|7|sed ego veritatem dico vobis expedit vobis ut ego vadam si enim non abiero paracletus non veniet ad vos si autem abiero mittam eum ad vos
JOHN|16|8|et cum venerit ille arguet mundum de peccato et de iustitia et de iudicio
JOHN|16|9|de peccato quidem quia non credunt in me
JOHN|16|10|de iustitia vero quia ad Patrem vado et iam non videbitis me
JOHN|16|11|de iudicio autem quia princeps mundi huius iudicatus est
JOHN|16|12|adhuc multa habeo vobis dicere sed non potestis portare modo
JOHN|16|13|cum autem venerit ille Spiritus veritatis docebit vos in omnem veritatem non enim loquetur a semet ipso sed quaecumque audiet loquetur et quae ventura sunt adnuntiabit vobis
JOHN|16|14|ille me clarificabit quia de meo accipiet et adnuntiabit vobis
JOHN|16|15|omnia quaecumque habet Pater mea sunt propterea dixi quia de meo accipit et adnuntiabit vobis
JOHN|16|16|modicum et iam non videbitis me et iterum modicum et videbitis me quia vado ad Patrem
JOHN|16|17|dixerunt ergo ex discipulis eius ad invicem quid est hoc quod dicit nobis modicum et non videbitis me et iterum modicum et videbitis me et quia vado ad Patrem
JOHN|16|18|dicebant ergo quid est hoc quod dicit modicum nescimus quid loquitur
JOHN|16|19|cognovit autem Iesus quia volebant eum interrogare et dixit eis de hoc quaeritis inter vos quia dixi modicum et non videbitis me et iterum modicum et videbitis me
JOHN|16|20|amen amen dico vobis quia plorabitis et flebitis vos mundus autem gaudebit vos autem contristabimini sed tristitia vestra vertetur in gaudium
JOHN|16|21|mulier cum parit tristitiam habet quia venit hora eius cum autem pepererit puerum iam non meminit pressurae propter gaudium quia natus est homo in mundum
JOHN|16|22|et vos igitur nunc quidem tristitiam habetis iterum autem videbo vos et gaudebit cor vestrum et gaudium vestrum nemo tollit a vobis
JOHN|16|23|et in illo die me non rogabitis quicquam amen amen dico vobis si quid petieritis Patrem in nomine meo dabit vobis
JOHN|16|24|usque modo non petistis quicquam in nomine meo petite et accipietis ut gaudium vestrum sit plenum
JOHN|16|25|haec in proverbiis locutus sum vobis venit hora cum iam non in proverbiis loquar vobis sed palam de Patre adnuntiabo vobis
JOHN|16|26|illo die in nomine meo petetis et non dico vobis quia ego rogabo Patrem de vobis
JOHN|16|27|ipse enim Pater amat vos quia vos me amastis et credidistis quia ego a Deo exivi
JOHN|16|28|exivi a Patre et veni in mundum iterum relinquo mundum et vado ad Patrem
JOHN|16|29|dicunt ei discipuli eius ecce nunc palam loqueris et proverbium nullum dicis
JOHN|16|30|nunc scimus quia scis omnia et non opus est tibi ut quis te interroget in hoc credimus quia a Deo existi
JOHN|16|31|respondit eis Iesus modo creditis
JOHN|16|32|ecce venit hora et iam venit ut dispergamini unusquisque in propria et me solum relinquatis et non sum solus quia Pater mecum est
JOHN|16|33|haec locutus sum vobis ut in me pacem habeatis in mundo pressuram habetis sed confidite ego vici mundum
JOHN|17|1|haec locutus est Iesus et sublevatis oculis in caelum dixit Pater venit hora clarifica Filium tuum ut Filius tuus clarificet te
JOHN|17|2|sicut dedisti ei potestatem omnis carnis ut omne quod dedisti ei det eis vitam aeternam
JOHN|17|3|haec est autem vita aeterna ut cognoscant te solum verum Deum et quem misisti Iesum Christum
JOHN|17|4|ego te clarificavi super terram opus consummavi quod dedisti mihi ut faciam
JOHN|17|5|et nunc clarifica me tu Pater apud temet ipsum claritatem quam habui priusquam mundus esset apud te
JOHN|17|6|manifestavi nomen tuum hominibus quos dedisti mihi de mundo tui erant et mihi eos dedisti et sermonem tuum servaverunt
JOHN|17|7|nunc cognoverunt quia omnia quae dedisti mihi abs te sunt
JOHN|17|8|quia verba quae dedisti mihi dedi eis et ipsi acceperunt et cognoverunt vere quia a te exivi et crediderunt quia tu me misisti
JOHN|17|9|ego pro eis rogo non pro mundo rogo sed pro his quos dedisti mihi quia tui sunt
JOHN|17|10|et mea omnia tua sunt et tua mea sunt et clarificatus sum in eis
JOHN|17|11|et iam non sum in mundo et hii in mundo sunt et ego ad te venio Pater sancte serva eos in nomine tuo quos dedisti mihi ut sint unum sicut et nos
JOHN|17|12|cum essem cum eis ego servabam eos in nomine tuo quos dedisti mihi custodivi et nemo ex his perivit nisi filius perditionis ut scriptura impleatur
JOHN|17|13|nunc autem ad te venio et haec loquor in mundo ut habeant gaudium meum impletum in semet ipsis
JOHN|17|14|ego dedi eis sermonem tuum et mundus odio eos habuit quia non sunt de mundo sicut et ego non sum de mundo
JOHN|17|15|non rogo ut tollas eos de mundo sed ut serves eos ex malo
JOHN|17|16|de mundo non sunt sicut et ego non sum de mundo
JOHN|17|17|sanctifica eos in veritate sermo tuus veritas est
JOHN|17|18|sicut me misisti in mundum et ego misi eos in mundum
JOHN|17|19|et pro eis ego sanctifico me ipsum ut sint et ipsi sanctificati in veritate
JOHN|17|20|non pro his autem rogo tantum sed et pro eis qui credituri sunt per verbum eorum in me
JOHN|17|21|ut omnes unum sint sicut tu Pater in me et ego in te ut et ipsi in nobis unum sint ut mundus credat quia tu me misisti
JOHN|17|22|et ego claritatem quam dedisti mihi dedi eis ut sint unum sicut nos unum sumus
JOHN|17|23|ego in eis et tu in me ut sint consummati in unum et cognoscat mundus quia tu me misisti et dilexisti eos sicut me dilexisti
JOHN|17|24|Pater quos dedisti mihi volo ut ubi ego sum et illi sint mecum ut videant claritatem meam quam dedisti mihi quia dilexisti me ante constitutionem mundi
JOHN|17|25|Pater iuste et mundus te non cognovit ego autem te cognovi et hii cognoverunt quia tu me misisti
JOHN|17|26|et notum feci eis nomen tuum et notum faciam ut dilectio qua dilexisti me in ipsis sit et ego in ipsis
JOHN|18|1|haec cum dixisset Iesus egressus est cum discipulis suis trans torrentem Cedron ubi erat hortus in quem introivit ipse et discipuli eius
JOHN|18|2|sciebat autem et Iudas qui tradebat eum ipsum locum quia frequenter Iesus convenerat illuc cum discipulis suis
JOHN|18|3|Iudas ergo cum accepisset cohortem et a pontificibus et Pharisaeis ministros venit illuc cum lanternis et facibus et armis
JOHN|18|4|Iesus itaque sciens omnia quae ventura erant super eum processit et dicit eis quem quaeritis
JOHN|18|5|responderunt ei Iesum Nazarenum dicit eis Iesus ego sum stabat autem et Iudas qui tradebat eum cum ipsis
JOHN|18|6|ut ergo dixit eis ego sum abierunt retrorsum et ceciderunt in terram
JOHN|18|7|iterum ergo eos interrogavit quem quaeritis illi autem dixerunt Iesum Nazarenum
JOHN|18|8|respondit Iesus dixi vobis quia ego sum si ergo me quaeritis sinite hos abire
JOHN|18|9|ut impleretur sermo quem dixit quia quos dedisti mihi non perdidi ex ipsis quemquam
JOHN|18|10|Simon ergo Petrus habens gladium eduxit eum et percussit pontificis servum et abscidit eius auriculam dextram erat autem nomen servo Malchus
JOHN|18|11|dixit ergo Iesus Petro mitte gladium in vaginam calicem quem dedit mihi Pater non bibam illum
JOHN|18|12|cohors ergo et tribunus et ministri Iudaeorum conprehenderunt Iesum et ligaverunt eum
JOHN|18|13|et adduxerunt eum ad Annam primum erat enim socer Caiaphae qui erat pontifex anni illius
JOHN|18|14|erat autem Caiaphas qui consilium dederat Iudaeis quia expedit unum hominem mori pro populo
JOHN|18|15|sequebatur autem Iesum Simon Petrus et alius discipulus discipulus autem ille erat notus pontifici et introivit cum Iesu in atrium pontificis
JOHN|18|16|Petrus autem stabat ad ostium foris exivit ergo discipulus alius qui erat notus pontifici et dixit ostiariae et introduxit Petrum
JOHN|18|17|dicit ergo Petro ancilla ostiaria numquid et tu ex discipulis es hominis istius dicit ille non sum
JOHN|18|18|stabant autem servi et ministri ad prunas quia frigus erat et calefiebant erat autem cum eis et Petrus stans et calefaciens se
JOHN|18|19|pontifex ergo interrogavit Iesum de discipulis suis et de doctrina eius
JOHN|18|20|respondit ei Iesus ego palam locutus sum mundo ego semper docui in synagoga et in templo quo omnes Iudaei conveniunt et in occulto locutus sum nihil
JOHN|18|21|quid me interrogas interroga eos qui audierunt quid locutus sum ipsis ecce hii sciunt quae dixerim ego
JOHN|18|22|haec autem cum dixisset unus adsistens ministrorum dedit alapam Iesu dicens sic respondes pontifici
JOHN|18|23|respondit ei Iesus si male locutus sum testimonium perhibe de malo si autem bene quid me caedis
JOHN|18|24|et misit eum Annas ligatum ad Caiaphan pontificem
JOHN|18|25|erat autem Simon Petrus stans et calefaciens se dixerunt ergo ei numquid et tu ex discipulis eius es negavit ille et dixit non sum
JOHN|18|26|dicit unus ex servis pontificis cognatus eius cuius abscidit Petrus auriculam nonne ego te vidi in horto cum illo
JOHN|18|27|iterum ergo negavit Petrus et statim gallus cantavit
JOHN|18|28|adducunt ergo Iesum a Caiapha in praetorium erat autem mane et ipsi non introierunt in praetorium ut non contaminarentur sed manducarent pascha
JOHN|18|29|exivit ergo Pilatus ad eos foras et dixit quam accusationem adfertis adversus hominem hunc
JOHN|18|30|responderunt et dixerunt ei si non esset hic malefactor non tibi tradidissemus eum
JOHN|18|31|dixit ergo eis Pilatus accipite eum vos et secundum legem vestram iudicate eum dixerunt ergo ei Iudaei nobis non licet interficere quemquam
JOHN|18|32|ut sermo Iesu impleretur quem dixit significans qua esset morte moriturus
JOHN|18|33|introivit ergo iterum in praetorium Pilatus et vocavit Iesum et dixit ei tu es rex Iudaeorum
JOHN|18|34|et respondit Iesus a temet ipso hoc dicis an alii tibi dixerunt de me
JOHN|18|35|respondit Pilatus numquid ego Iudaeus sum gens tua et pontifices tradiderunt te mihi quid fecisti
JOHN|18|36|respondit Iesus regnum meum non est de mundo hoc si ex hoc mundo esset regnum meum ministri mei decertarent ut non traderer Iudaeis nunc autem meum regnum non est hinc
JOHN|18|37|dixit itaque ei Pilatus ergo rex es tu respondit Iesus tu dicis quia rex sum ego ego in hoc natus sum et ad hoc veni in mundum ut testimonium perhibeam veritati omnis qui est ex veritate audit meam vocem
JOHN|18|38|dicit ei Pilatus quid est veritas et cum hoc dixisset iterum exivit ad Iudaeos et dicit eis ego nullam invenio in eo causam
JOHN|18|39|est autem consuetudo vobis ut unum dimittam vobis in pascha vultis ergo dimittam vobis regem Iudaeorum
JOHN|18|40|clamaverunt rursum omnes dicentes non hunc sed Barabban erat autem Barabbas latro
JOHN|19|1|tunc ergo adprehendit Pilatus Iesum et flagellavit
JOHN|19|2|et milites plectentes coronam de spinis inposuerunt capiti eius et veste purpurea circumdederunt eum
JOHN|19|3|et veniebant ad eum et dicebant have rex Iudaeorum et dabant ei alapas
JOHN|19|4|exiit iterum Pilatus foras et dicit eis ecce adduco vobis eum foras
JOHN|19|5|ut cognoscatis quia in eo nullam causam invenio et purpureum vestimentum et dicit eis ecce homo
JOHN|19|6|cum ergo vidissent eum pontifices et ministri clamabant dicentes crucifige crucifige dicit eis Pilatus accipite eum vos et crucifigite ego enim non invenio in eo causam
JOHN|19|7|responderunt ei Iudaei nos legem habemus et secundum legem debet mori quia Filium Dei se fecit
JOHN|19|8|cum ergo audisset Pilatus hunc sermonem magis timuit
JOHN|19|9|et ingressus est praetorium iterum et dicit ad Iesum unde es tu Iesus autem responsum non dedit ei
JOHN|19|10|dicit ergo ei Pilatus mihi non loqueris nescis quia potestatem habeo crucifigere te et potestatem habeo dimittere te
JOHN|19|11|respondit Iesus non haberes potestatem adversum me ullam nisi tibi esset datum desuper propterea qui tradidit me tibi maius peccatum habet
JOHN|19|12|exinde quaerebat Pilatus dimittere eum Iudaei autem clamabant dicentes si hunc dimittis non es amicus Caesaris omnis qui se regem facit contradicit Caesari
JOHN|19|13|Pilatus ergo cum audisset hos sermones adduxit foras Iesum et sedit pro tribunali in locum qui dicitur Lithostrotus hebraice autem Gabbatha
JOHN|19|14|erat autem parasceve paschae hora quasi sexta et dicit Iudaeis ecce rex vester
JOHN|19|15|illi autem clamabant tolle tolle crucifige eum dixit eis Pilatus regem vestrum crucifigam responderunt pontifices non habemus regem nisi Caesarem
JOHN|19|16|tunc ergo tradidit eis illum ut crucifigeretur susceperunt autem Iesum et eduxerunt
JOHN|19|17|et baiulans sibi crucem exivit in eum qui dicitur Calvariae locum hebraice Golgotha
JOHN|19|18|ubi eum crucifixerunt et cum eo alios duos hinc et hinc medium autem Iesum
JOHN|19|19|scripsit autem et titulum Pilatus et posuit super crucem erat autem scriptum Iesus Nazarenus rex Iudaeorum
JOHN|19|20|hunc ergo titulum multi legerunt Iudaeorum quia prope civitatem erat locus ubi crucifixus est Iesus et erat scriptum hebraice graece et latine
JOHN|19|21|dicebant ergo Pilato pontifices Iudaeorum noli scribere rex Iudaeorum sed quia ipse dixit rex sum Iudaeorum
JOHN|19|22|respondit Pilatus quod scripsi scripsi
JOHN|19|23|milites ergo cum crucifixissent eum acceperunt vestimenta eius et fecerunt quattuor partes unicuique militi partem et tunicam erat autem tunica inconsutilis desuper contexta per totum
JOHN|19|24|dixerunt ergo ad invicem non scindamus eam sed sortiamur de illa cuius sit ut scriptura impleatur dicens partiti sunt vestimenta mea sibi et in vestem meam miserunt sortem et milites quidem haec fecerunt
JOHN|19|25|stabant autem iuxta crucem Iesu mater eius et soror matris eius Maria Cleopae et Maria Magdalene
JOHN|19|26|cum vidisset ergo Iesus matrem et discipulum stantem quem diligebat dicit matri suae mulier ecce filius tuus
JOHN|19|27|deinde dicit discipulo ecce mater tua et ex illa hora accepit eam discipulus in sua
JOHN|19|28|postea sciens Iesus quia iam omnia consummata sunt ut consummaretur scriptura dicit sitio
JOHN|19|29|vas ergo positum erat aceto plenum illi autem spongiam plenam aceto hysopo circumponentes obtulerunt ori eius
JOHN|19|30|cum ergo accepisset Iesus acetum dixit consummatum est et inclinato capite tradidit spiritum
JOHN|19|31|Iudaei ergo quoniam parasceve erat ut non remanerent in cruce corpora sabbato erat enim magnus dies ille sabbati rogaverunt Pilatum ut frangerentur eorum crura et tollerentur
JOHN|19|32|venerunt ergo milites et primi quidem fregerunt crura et alterius qui crucifixus est cum eo
JOHN|19|33|ad Iesum autem cum venissent ut viderunt eum iam mortuum non fregerunt eius crura
JOHN|19|34|sed unus militum lancea latus eius aperuit et continuo exivit sanguis et aqua
JOHN|19|35|et qui vidit testimonium perhibuit et verum est eius testimonium et ille scit quia vera dicit ut et vos credatis
JOHN|19|36|facta sunt enim haec ut scriptura impleatur os non comminuetis ex eo
JOHN|19|37|et iterum alia scriptura dicit videbunt in quem transfixerunt
JOHN|19|38|post haec autem rogavit Pilatum Ioseph ab Arimathia eo quod esset discipulus Iesu occultus autem propter metum Iudaeorum ut tolleret corpus Iesu et permisit Pilatus venit ergo et tulit corpus Iesu
JOHN|19|39|venit autem et Nicodemus qui venerat ad Iesum nocte primum ferens mixturam murrae et aloes quasi libras centum
JOHN|19|40|acceperunt ergo corpus Iesu et ligaverunt eum linteis cum aromatibus sicut mos Iudaeis est sepelire
JOHN|19|41|erat autem in loco ubi crucifixus est hortus et in horto monumentum novum in quo nondum quisquam positus erat
JOHN|19|42|ibi ergo propter parasceven Iudaeorum quia iuxta erat monumentum posuerunt Iesum
JOHN|20|1|una autem sabbati Maria Magdalene venit mane cum adhuc tenebrae essent ad monumentum et videt lapidem sublatum a monumento
JOHN|20|2|cucurrit ergo et venit ad Simonem Petrum et ad alium discipulum quem amabat Iesus et dicit eis tulerunt Dominum de monumento et nescimus ubi posuerunt eum
JOHN|20|3|exiit ergo Petrus et ille alius discipulus et venerunt ad monumentum
JOHN|20|4|currebant autem duo simul et ille alius discipulus praecucurrit citius Petro et venit primus ad monumentum
JOHN|20|5|et cum se inclinasset videt posita linteamina non tamen introivit
JOHN|20|6|venit ergo Simon Petrus sequens eum et introivit in monumentum et videt linteamina posita
JOHN|20|7|et sudarium quod fuerat super caput eius non cum linteaminibus positum sed separatim involutum in unum locum
JOHN|20|8|tunc ergo introivit et ille discipulus qui venerat primus ad monumentum et vidit et credidit
JOHN|20|9|nondum enim sciebant scripturam quia oportet eum a mortuis resurgere
JOHN|20|10|abierunt ergo iterum ad semet ipsos discipuli
JOHN|20|11|Maria autem stabat ad monumentum foris plorans dum ergo fleret inclinavit se et prospexit in monumentum
JOHN|20|12|et vidit duos angelos in albis sedentes unum ad caput et unum ad pedes ubi positum fuerat corpus Iesu
JOHN|20|13|dicunt ei illi mulier quid ploras dicit eis quia tulerunt Dominum meum et nescio ubi posuerunt eum
JOHN|20|14|haec cum dixisset conversa est retrorsum et videt Iesum stantem et non sciebat quia Iesus est
JOHN|20|15|dicit ei Iesus mulier quid ploras quem quaeris illa existimans quia hortulanus esset dicit ei domine si tu sustulisti eum dicito mihi ubi posuisti eum et ego eum tollam
JOHN|20|16|dicit ei Iesus Maria conversa illa dicit ei rabboni quod dicitur magister
JOHN|20|17|dicit ei Iesus noli me tangere nondum enim ascendi ad Patrem meum vade autem ad fratres meos et dic eis ascendo ad Patrem meum et Patrem vestrum et Deum meum et Deum vestrum
JOHN|20|18|venit Maria Magdalene adnuntians discipulis quia vidi Dominum et haec dixit mihi
JOHN|20|19|cum esset ergo sero die illo una sabbatorum et fores essent clausae ubi erant discipuli propter metum Iudaeorum venit Iesus et stetit in medio et dicit eis pax vobis
JOHN|20|20|et hoc cum dixisset ostendit eis manus et latus gavisi sunt ergo discipuli viso Domino
JOHN|20|21|dixit ergo eis iterum pax vobis sicut misit me Pater et ego mitto vos
JOHN|20|22|hoc cum dixisset insuflavit et dicit eis accipite Spiritum Sanctum
JOHN|20|23|quorum remiseritis peccata remittuntur eis quorum retinueritis detenta sunt
JOHN|20|24|Thomas autem unus ex duodecim qui dicitur Didymus non erat cum eis quando venit Iesus
JOHN|20|25|dixerunt ergo ei alii discipuli vidimus Dominum ille autem dixit eis nisi videro in manibus eius figuram clavorum et mittam digitum meum in locum clavorum et mittam manum meam in latus eius non credam
JOHN|20|26|et post dies octo iterum erant discipuli eius intus et Thomas cum eis venit Iesus ianuis clausis et stetit in medio et dixit pax vobis
JOHN|20|27|deinde dicit Thomae infer digitum tuum huc et vide manus meas et adfer manum tuam et mitte in latus meum et noli esse incredulus sed fidelis
JOHN|20|28|respondit Thomas et dixit ei Dominus meus et Deus meus
JOHN|20|29|dicit ei Iesus quia vidisti me credidisti beati qui non viderunt et crediderunt
JOHN|20|30|multa quidem et alia signa fecit Iesus in conspectu discipulorum suorum quae non sunt scripta in libro hoc
JOHN|20|31|haec autem scripta sunt ut credatis quia Iesus est Christus Filius Dei et ut credentes vitam habeatis in nomine eius
JOHN|21|1|postea manifestavit se iterum Iesus ad mare Tiberiadis manifestavit autem sic
JOHN|21|2|erant simul Simon Petrus et Thomas qui dicitur Didymus et Nathanahel qui erat a Cana Galilaeae et filii Zebedaei et alii ex discipulis eius duo
JOHN|21|3|dicit eis Simon Petrus vado piscari dicunt ei venimus et nos tecum et exierunt et ascenderunt in navem et illa nocte nihil prendiderunt
JOHN|21|4|mane autem iam facto stetit Iesus in litore non tamen cognoverunt discipuli quia Iesus est
JOHN|21|5|dicit ergo eis Iesus pueri numquid pulmentarium habetis responderunt ei non
JOHN|21|6|dixit eis mittite in dexteram navigii rete et invenietis miserunt ergo et iam non valebant illud trahere a multitudine piscium
JOHN|21|7|dicit ergo discipulus ille quem diligebat Iesus Petro Dominus est Simon Petrus cum audisset quia Dominus est tunicam succinxit se erat enim nudus et misit se in mare
JOHN|21|8|alii autem discipuli navigio venerunt non enim longe erant a terra sed quasi a cubitis ducentis trahentes rete piscium
JOHN|21|9|ut ergo descenderunt in terram viderunt prunas positas et piscem superpositum et panem
JOHN|21|10|dicit eis Iesus adferte de piscibus quos prendidistis nunc
JOHN|21|11|ascendit Simon Petrus et traxit rete in terram plenum magnis piscibus centum quinquaginta tribus et cum tanti essent non est scissum rete
JOHN|21|12|dicit eis Iesus venite prandete et nemo audebat discentium interrogare eum tu quis es scientes quia Dominus esset
JOHN|21|13|et venit Iesus et accepit panem et dat eis et piscem similiter
JOHN|21|14|hoc iam tertio manifestatus est Iesus discipulis cum surrexisset a mortuis
JOHN|21|15|cum ergo prandissent dicit Simoni Petro Iesus Simon Iohannis diligis me plus his dicit ei etiam Domine tu scis quia amo te dicit ei pasce agnos meos
JOHN|21|16|dicit ei iterum Simon Iohannis diligis me ait illi etiam Domine tu scis quia amo te dicit ei pasce agnos meos
JOHN|21|17|dicit ei tertio Simon Iohannis amas me contristatus est Petrus quia dixit ei tertio amas me et dicit ei Domine tu omnia scis tu scis quia amo te dicit ei pasce oves meas
JOHN|21|18|amen amen dico tibi cum esses iunior cingebas te et ambulabas ubi volebas cum autem senueris extendes manus tuas et alius te cinget et ducet quo non vis
JOHN|21|19|hoc autem dixit significans qua morte clarificaturus esset Deum et hoc cum dixisset dicit ei sequere me
JOHN|21|20|conversus Petrus vidit illum discipulum quem diligebat Iesus sequentem qui et recubuit in cena super pectus eius et dixit Domine quis est qui tradit te
JOHN|21|21|hunc ergo cum vidisset Petrus dicit Iesu Domine hic autem quid
JOHN|21|22|dicit ei Iesus si sic eum volo manere donec veniam quid ad te tu me sequere
JOHN|21|23|exivit ergo sermo iste in fratres quia discipulus ille non moritur et non dixit ei Iesus non moritur sed si sic eum volo manere donec venio quid ad te
JOHN|21|24|hic est discipulus qui testimonium perhibet de his et scripsit haec et scimus quia verum est testimonium eius
JOHN|21|25|sunt autem et alia multa quae fecit Iesus quae si scribantur per singula nec ipsum arbitror mundum capere eos qui scribendi sunt libros amen
