NEH|1|1|verba Neemiae filii Echliae et factum est in mense casleu anno vicesimo et ego eram in Susis castro
NEH|1|2|et venit Anani unus de fratribus meis ipse et viri ex Iuda et interrogavi eos de Iudaeis qui remanserant et supererant de captivitate et de Hierusalem
NEH|1|3|et dixerunt mihi qui remanserunt et derelicti sunt de captivitate ibi in provincia in adflictione magna sunt et in obprobrio et murus Hierusalem dissipatus est et portae eius conbustae sunt igni
NEH|1|4|cumque audissem verba huiuscemodi sedi et flevi et luxi diebus et ieiunabam et orabam ante faciem Dei caeli
NEH|1|5|et dixi quaeso Domine Deus caeli fortis magne atque terribilis qui custodis pactum et misericordiam cum his qui te diligunt et custodiunt mandata tua
NEH|1|6|fiat auris tua auscultans et oculi tui aperti ut audias orationem servi tui quam ego oro coram te hodie nocte et die pro filiis Israhel servis tuis et confiteor pro peccatis filiorum Israhel quibus peccaverunt tibi et ego et domus patris mei peccavimus
NEH|1|7|vanitate seducti sumus et non custodivimus mandatum et caerimonias et iudicia quae praecepisti Mosi servo tuo
NEH|1|8|memento verbi quod mandasti Mosi famulo tuo dicens cum transgressi fueritis ego dispergam vos in populos
NEH|1|9|et si revertamini ad me et custodiatis mandata mea et faciatis ea etiam si abducti fueritis ad extrema caeli inde congregabo vos et inducam in locum quem elegi ut habitaret nomen meum ibi
NEH|1|10|et ipsi servi tui et populus tuus quos redemisti in fortitudine tua magna et in manu tua valida
NEH|1|11|obsecro Domine sit auris tua adtendens ad orationem servi tui et ad orationem servorum tuorum qui volunt timere nomen tuum et dirige servum tuum hodie et da ei misericordiam ante virum hunc ego enim eram pincerna regis
NEH|2|1|factum est autem in mense nisan anno vicesimo Artarxersis regis et vinum erat ante eum et levavi vinum et dedi regi et non eram quasi languidus ante faciem eius
NEH|2|2|dixitque mihi rex quare vultus tuus tristis cum te aegrotum non videam non est hoc frustra sed malum nescio quid in corde tuo est et timui valde ac nimis
NEH|2|3|et dixi regi rex in aeternum vive quare non maereat vultus meus quia civitas domus sepulchrorum patris mei deserta est et portae eius conbustae sunt igni
NEH|2|4|et ait mihi rex pro qua re postulas et oravi Deum caeli
NEH|2|5|et dixi ad regem si videtur regi bonum et si placet servus tuus ante faciem tuam ut mittas me in Iudaeam ad civitatem sepulchri patris mei et aedificabo eam
NEH|2|6|dixitque mihi rex et regina quae sedebat iuxta eum usque ad quod tempus erit iter tuum et quando reverteris et placuit ante vultum regis et misit me et constitui ei tempus
NEH|2|7|et dixi regi si regi videtur bonum epistulas det mihi ad duces regionis trans Flumen ut transducant me donec veniam in Iudaeam
NEH|2|8|et epistulam ad Asaph custodem saltus regis ut det mihi ligna et tegere possim portas turris domus et muri civitatis et domum quam ingressus fuero et dedit mihi rex iuxta manum Dei mei bonam mecum
NEH|2|9|et veni ad duces regionis trans Flumen dedique eis epistulas regis miserat autem mecum rex principes militum et equites
NEH|2|10|et audierunt Sanaballat Horonites et Tobias servus ammanites et contristati sunt adflictione magna quod venisset homo qui quaereret prosperitatem filiorum Israhel
NEH|2|11|et veni Hierusalem et eram ibi diebus tribus
NEH|2|12|et surrexi nocte ego et viri pauci mecum et non indicavi cuiquam quid Deus dedisset in corde meo ut facerem in Hierusalem et iumentum non erat mecum nisi animal cui sedebam
NEH|2|13|et egressus sum per portam Vallis nocte et ante fontem Draconis et ad portam Stercoris et considerabam murum Hierusalem dissipatum et portas eius consumptas igni
NEH|2|14|et transivi ad portam Fontis et ad aquaeductum Regis et non erat locus iumento cui sedebam ut transiret
NEH|2|15|et ascendi per torrentem nocte et considerabam murum et reversus veni ad portam Vallis et redii
NEH|2|16|magistratus autem nesciebant quo abissem aut quid ego facerem sed et Iudaeis et sacerdotibus et optimatibus et magistratibus et reliquis qui faciebant opus usque ad id locorum nihil indicaveram
NEH|2|17|et dixi eis vos nostis adflictionem in qua sumus quia Hierusalem deserta est et portae eius consumptae sunt igni venite et aedificemus muros Hierusalem et non simus ultra obprobrium
NEH|2|18|et indicavi eis manum Dei mei quod esset bona mecum et verba regis quae locutus est mihi et aio surgamus et aedificemus et confortatae sunt manus eorum in bono
NEH|2|19|audierunt autem Sanaballat Horonites et Tobias servus ammanites et Gosem Arabs et subsannaverunt nos et despexerunt dixeruntque quae est haec res quam facitis numquid contra regem vos rebellatis
NEH|2|20|et reddidi eis sermonem dixique ad eos Deus caeli ipse nos iuvat et nos servi eius sumus surgamus et aedificemus vobis autem non est pars et iustitia et memoria in Hierusalem
NEH|3|1|et surrexit Eliasib sacerdos magnus et fratres eius sacerdotes et aedificaverunt portam Gregis ipsi sanctificaverunt eam et statuerunt valvas eius et usque ad turrem centum cubitorum sanctificaverunt eam usque ad turrem Ananehel
NEH|3|2|et iuxta eum aedificaverunt viri Hiericho et iuxta eum aedificavit Zecchur filius Amri
NEH|3|3|portam autem Piscium aedificaverunt filii Asanaa ipsi texerunt eam et statuerunt valvas eius et seras et vectes et iuxta eos aedificavit Marimuth filius Uriae filii Accus
NEH|3|4|et iuxta eos aedificavit Mosollam filius Barachiae filii Mesezebel et iuxta eos aedificavit Sadoc filius Baana
NEH|3|5|et iuxta eos aedificaverunt Thecueni optimates autem eorum non subposuerunt colla sua in opere Domini sui
NEH|3|6|et portam Veterem aedificaverunt Ioiada filius Fasea et Mosollam filius Besodia ipsi texerunt eam et statuerunt valvas eius et seras et vectes
NEH|3|7|et iuxta eos aedificavit Meletias Gabaonites et Iadon Meronathites viri de Gabaon et Maspha pro duce qui erat in regione trans Flumen
NEH|3|8|et iuxta eum aedificavit Ezihel filius Araia aurifex et iuxta eum aedificavit Anania filius pigmentarii et dimiserunt Hierusalem usque ad murum plateae latioris
NEH|3|9|et iuxta eum aedificavit Rafaia filius Ahur princeps vici Hierusalem
NEH|3|10|et iuxta eos aedificavit Ieiada filius Aromath contra domum suam et iuxta eum aedificavit Attus filius Asebeniae
NEH|3|11|mediam partem vici aedificavit Melchias filius Erem et Asub filius Phaethmoab et turrem Furnorum
NEH|3|12|iuxta eum aedificavit Sellum filius Alloes princeps mediae partis vici Hierusalem ipse et filiae eius
NEH|3|13|et portam Vallis aedificavit Anun et habitatores Zanoe ipsi aedificaverunt eam et statuerunt valvas eius et seras et vectes et mille cubitos in muro usque ad portam Sterquilinii
NEH|3|14|et portam Sterquilinii aedificavit Melchias filius Rechab princeps vici Bethaccharem ipse aedificavit eam et statuit valvas eius et seras et vectes
NEH|3|15|et portam Fontis aedificavit Sellum filius Choloozai princeps pagi Maspha ipse aedificavit eam et texit et statuit valvas eius et seras et vectes et muros piscinae Siloae in hortum regis et usque ad gradus qui descendunt de civitate David
NEH|3|16|post eum aedificavit Neemias filius Azboc princeps dimidiae partis vici Bethsur usque contra sepulchra David et usque ad piscinam quae grandi opere constructa est et usque ad domum Fortium
NEH|3|17|post eum aedificaverunt Levitae Reum filius Benni post eum aedificavit Asebias princeps dimidiae partis vici Ceilae in vico suo
NEH|3|18|post eum aedificaverunt fratres eorum Behui filius Enadad princeps dimidiae partis Ceila
NEH|3|19|et aedificavit iuxta eum Azer filius Iosue princeps Maspha mensuram secundam contra ascensum firmissimi anguli
NEH|3|20|post eum in monte aedificavit Baruch filius Zacchai mensuram secundam ab angulo usque ad portam domus Eliasib sacerdotis magni
NEH|3|21|post eum aedificavit Meremuth filius Uriae filii Accus mensuram secundam a porta domus Eliasib donec extenderetur domus Eliasib
NEH|3|22|et post eum aedificaverunt sacerdotes viri de campestribus Iordanis
NEH|3|23|post eum aedificavit Beniamin et Asub contra domum suam et post eum aedificavit Azarias filius Maasiae filii Ananiae contra domum suam
NEH|3|24|post eum aedificavit Bennui filius Enadda mensuram secundam a domo Azariae usque ad flexuram et usque ad angulum
NEH|3|25|Falel filius Ozi contra flexuram et turrem quae eminet de domo regis excelsa id est in atrio carceris post eum Phadaia filius Pheros
NEH|3|26|Nathinnei autem habitabant in Ofel usque contra portam Aquarum ad orientem et turrem quae prominebat
NEH|3|27|post eum aedificaverunt Thecueni mensuram secundam e regione a turre magna et eminenti usque ad murum templi
NEH|3|28|sursum autem a porta Equorum aedificaverunt sacerdotes unusquisque contra domum suam
NEH|3|29|post eos aedificavit Seddo filius Emmer contra domum suam et post eum aedificavit Semeia filius Secheniae custos portae orientalis
NEH|3|30|post eum aedificavit Anania filius Selemiae et Anon filius Selo sextus mensuram secundam post eum aedificavit Mosollam filius Barachiae contra gazofilacium suum post eum aedificavit Melchias filius aurificis usque ad domum Nathinneorum et scruta vendentium contra portam Iudicialem et usque ad cenaculum Anguli
NEH|3|31|et inter cenaculum Anguli in porta Gregis aedificaverunt artifices et negotiatores
NEH|4|1|factum est autem cum audisset Sanaballat quod aedificaremus murum iratus est valde et motus nimis subsannavit Iudaeos
NEH|4|2|et dixit coram fratribus suis et frequentia Samaritanorum quid Iudaei inbecilli faciunt num dimittent eos gentes num sacrificabunt et conplebunt in una die numquid aedificare poterunt lapides de acervis pulveris qui conbusti sunt
NEH|4|3|sed et Tobias Ammanites proximus eius ait aedificent si ascenderit vulpis transiliet murum eorum lapideum
NEH|4|4|audi Deus noster quia facti sumus despectio converte obprobrium super caput eorum et da eos in despectionem in terra captivitatis
NEH|4|5|ne operias iniquitatem eorum et peccatum eorum coram facie tua non deleatur quia inriserunt aedificantes
NEH|4|6|itaque aedificavimus murum et coniunximus totum usque ad partem dimidiam et provocatum est cor populi ad operandum
NEH|4|7|factum est autem cum audisset Sanaballat et Tobias et Arabes et Ammanitae et Azotii quod obducta esset cicatrix muri Hierusalem et quod coepissent interrupta concludi irati sunt nimis
NEH|4|8|et congregati omnes pariter ut venirent et pugnarent contra Hierusalem et molirentur insidias
NEH|4|9|et oravimus Deum nostrum et posuimus custodes super murum die et nocte contra eos
NEH|4|10|dixit autem Iudas debilitata est fortitudo portantis et humus nimia est et nos non poterimus aedificare murum
NEH|4|11|et dixerunt hostes nostri nesciant et ignorent donec veniamus in medio eorum et interficiamus eos et cessare faciamus opus
NEH|4|12|factum est autem venientibus Iudaeis qui habitabant iuxta eos et dicentibus nobis per decem vices ex omnibus locis quibus venerant ad nos
NEH|4|13|statui in loco post murum per circuitum populum in ordine cum gladiis suis et lanceis et arcis
NEH|4|14|perspexi atque surrexi et aio ad optimates et ad magistratus et ad reliquam partem vulgi nolite timere a facie eorum Domini magni et terribilis mementote et pugnate pro fratribus vestris filiis vestris et filiabus vestris uxoribus vestris et domibus
NEH|4|15|factum est autem cum audissent inimici nostri nuntiatum esse nobis dissipavit Deus consilium eorum et reversi sumus omnes ad muros unusquisque ad opus suum
NEH|4|16|et factum est a die illa media pars iuvenum eorum faciebant opus et media parata erat ad bellum et lanceae et scuta et arcus et loricae et principes post eos in omni domo Iuda
NEH|4|17|aedificantium in muro et portantium onera et inponentium una manu sua faciebat opus et altera tenebat gladium
NEH|4|18|aedificantium enim unusquisque gladio erat accinctus renes et aedificabant et clangebant bucina iuxta me
NEH|4|19|et dixi ad optimates et ad magistratus et ad reliquam partem vulgi opus grande est et latum et nos separati sumus in muro procul alter ab altero
NEH|4|20|in loco quocumque audieritis clangorem tubae illuc concurrite ad nos Deus noster pugnabit pro nobis
NEH|4|21|et nos ipsi faciamus opus et media pars nostrum teneat lanceas ab ascensu aurorae donec egrediantur astra
NEH|4|22|in tempore quoque illo dixi populo unusquisque cum puero suo maneat in medio Hierusalem et sint vobis vices per noctem et diem ad operandum
NEH|4|23|ego autem et fratres mei et pueri mei et custodes qui erant post me non deponebamus vestimenta nostra unusquisque tantum nudabatur ad baptismum
NEH|5|1|et factus est clamor populi et uxorum eius magnus adversus fratres suos iudaeos
NEH|5|2|et erant qui dicerent filii nostri et filiae nostrae multae sunt nimis accipiamus pro pretio eorum frumentum et comedamus et vivamus
NEH|5|3|et erant qui dicerent agros nostros et vineas et domos nostras opponamus et accipiamus frumentum in fame
NEH|5|4|et alii dicebant mutuo sumamus pecunias in tributa regis demusque agros nostros et vineas
NEH|5|5|et nunc sicut carnes fratrum nostrorum sic carnes nostrae sunt sicut filii eorum ita filii nostri ecce nos subiugamus filios nostros et filias nostras in servitutem et de filiabus nostris sunt famulae nec habemus unde possint redimi et agros nostros et vineas alii possident
NEH|5|6|et iratus sum nimis cum audissem clamorem eorum secundum verba haec
NEH|5|7|cogitavitque cor meum mecum et increpui optimates et magistratus et dixi eis usurasne singuli a fratribus vestris exigatis et congregavi adversus eos contionem magnam
NEH|5|8|et dixi eis nos ut scitis redemimus fratres nostros iudaeos qui venditi fuerant gentibus secundum possibilitatem nostram et vos igitur vendite fratres vestros et emimus eos et siluerunt nec invenerunt quid responderent
NEH|5|9|dixique ad eos non est bona res quam facitis quare non in timore Dei nostri ambulatis ne exprobretur nobis a gentibus inimicis nostris
NEH|5|10|et ego et fratres mei et pueri mei commodavimus plurimis pecuniam et frumentum non repetamus in commune istud aes alienum concedamus quod debetur nobis
NEH|5|11|reddite eis hodie agros suos vineas suas oliveta sua et domos suas quin potius et centesimam pecuniae frumenti vini et olei quam exigere soletis ab eis date pro illis
NEH|5|12|et dixerunt reddimus et ab eis nihil quaerimus sicque faciemus ut loqueris et vocavi sacerdotes et adiuravi eos ut facerent iuxta quod dixeram
NEH|5|13|insuper et sinum meum excussi et dixi sic excutiat Deus omnem virum qui non conpleverit verbum istud de domo sua et de laboribus suis sic excutiatur et vacuus fiat et dixit universa multitudo amen et laudaverunt Deum fecit ergo populus sicut dictum erat
NEH|5|14|a die autem illa qua praeceperat mihi ut essem dux in terra Iuda ab anno vicesimo usque ad annum tricesimum secundum Artarxersis regis per annos duodecim ego et fratres mei annonas quae ducibus debebantur non comedimus
NEH|5|15|duces autem primi qui fuerant ante me gravaverunt populum et acceperunt ab eis in pane vino et pecunia cotidie siclos quadraginta sed et ministri eorum depresserant populum ego autem non feci ita propter timorem Dei
NEH|5|16|quin potius in opere muri aedificavi et agrum non emi et omnes pueri mei congregati ad opus erant
NEH|5|17|Iudaei quoque et magistratus centum quinquaginta viri et qui veniebant ad nos de gentibus quae in circuitu nostro sunt in mensa mea erant
NEH|5|18|parabatur autem mihi per dies singulos bos unus arietes sex electi exceptis volatilibus et inter dies decem vina diversa et alia multa tribuebam insuper et annonas ducatus mei non quaesivi valde enim erat adtenuatus populus
NEH|5|19|memento mei Deus meus in bonum secundum omnia quae feci populo huic
NEH|6|1|factum est autem cum audisset Sanaballat et Tobia et Gosem Arabs et ceteri inimici nostri quod aedificassem ego murum et non esset in ipso residua interruptio usque ad tempus autem illud valvas non posueram in portis
NEH|6|2|miserunt Sanaballat et Gosem ad me dicentes veni et percutiamus foedus pariter in viculis in campo Ono ipsi autem cogitabant ut facerent mihi malum
NEH|6|3|misi ergo ad eos nuntios dicens opus grande ego facio et non possum descendere ne forte neglegatur cum venero et descendero ad vos
NEH|6|4|miserunt autem ad me secundum verbum hoc per quattuor vices et respondi eis iuxta sermonem priorem
NEH|6|5|et misit ad me Sanaballat iuxta verbum prius quinta vice puerum suum et epistulam habebat in manu scriptam hoc modo
NEH|6|6|in gentibus auditum est et Gosem dixit quod tu et Iudaei cogitetis rebellare et propterea aedifices murum et levare te velis super eos regem propter quam causam
NEH|6|7|et prophetas posueris qui praedicent de te in Hierusalem dicentes rex in Iudaea est auditurus est rex verba haec idcirco nunc veni ut ineamus consilium pariter
NEH|6|8|et misi ad eos dicens non est factum secundum verba haec quae tu loqueris de corde enim tuo tu conponis haec
NEH|6|9|omnes autem hii terrebant nos cogitantes quod cessarent manus nostrae ab opere et quiesceremus quam ob causam magis confortavi manus meas
NEH|6|10|et ingressus sum domum Samaiae filii Dalaiae filii Metabehel secreto qui ait tractemus nobiscum in domo Dei in medio templi et claudamus portas aedis quia venturi sunt ut interficiant te et nocte venturi sunt ad occidendum te
NEH|6|11|et dixi num quisquam similis mei fugit et quis ut ego ingredietur templum et vivet non ingrediar
NEH|6|12|et intellexi quod Deus non misisset eum sed quasi vaticinans locutus esset ad me et Tobia et Sanaballat conduxissent eum
NEH|6|13|acceperat enim pretium ut territus facerem et peccarem et haberent malum quod exprobrarent mihi
NEH|6|14|memento Domine mei pro Tobia et Sanaballat iuxta opera eorum talia sed et Noadiae prophetae et ceterorum prophetarum qui terrebant me
NEH|6|15|conpletus est autem murus vicesimo quinto die mensis elul quinquaginta duobus diebus
NEH|6|16|factum est ergo cum audissent omnes inimici nostri ut timerent universae gentes quae erant in circuitu nostro et conciderent intra semet ipsos et scirent quod a Deo factum esset opus hoc
NEH|6|17|sed et in diebus illis multae optimatium Iudaeorum epistulae mittebantur ad Tobiam et a Tobia veniebant ad eos
NEH|6|18|multi enim erant in Iudaea habentes iuramentum eius quia gener erat Secheniae filii Orei et Iohanan filius eius acceperat filiam Mosollam filii Barachiae
NEH|6|19|sed et laudabant eum coram me et verba mea nuntiabant ei et Tobias mittebat epistulas ut terreret me
NEH|7|1|postquam autem aedificatus est murus et posui valvas et recensui ianitores et cantores et Levitas
NEH|7|2|praecepi Aneni fratri meo et Ananiae principi domus de Hierusalem ipse enim quasi vir verax et timens Deum plus ceteris videbatur
NEH|7|3|et dixi eis non aperiantur portae Hierusalem usque ad calorem solis cumque adhuc adsisterent clausae portae sunt et oppilatae et posui custodes de habitatoribus Hierusalem singulos per vices suas et unumquemque contra domum suam
NEH|7|4|civitas autem erat lata nimis et grandis et populus parvus in medio eius et non erant domus aedificatae
NEH|7|5|dedit autem Deus in corde meo et congregavi optimates et magistratus et vulgum ut recenserem eos et inveni librum census eorum qui ascenderant primum et inventum est scriptum in eo
NEH|7|6|isti filii provinciae qui ascenderunt de captivitate migrantium quos transtulerat Nabuchodonosor rex Babylonis et reversi sunt in Hierusalem et in Iudaeam unusquisque in civitatem suam
NEH|7|7|qui venerunt cum Zorobabel Hiesuae Neemias Azarias Raamias Naamni Mardocheus Belsar Mespharath Beggoai Naum Baana numerus virorum populi Israhel
NEH|7|8|filii Pharos duo milia centum septuaginta duo
NEH|7|9|filii Saphatiae trecenti septuaginta duo
NEH|7|10|filii Area sescenti quinquaginta duo
NEH|7|11|filii Phaethmoab filiorum Hiesuae et Ioab duo milia octingenti decem et octo
NEH|7|12|filii Helam mille octingenti quinquaginta quattuor
NEH|7|13|filii Zethua octingenti quadraginta quinque
NEH|7|14|filii Zacchai septingenti sexaginta
NEH|7|15|filii Bennui sescenti quadraginta octo
NEH|7|16|filii Bebai sescenti viginti octo
NEH|7|17|filii Azgad duo milia trecenti viginti duo
NEH|7|18|filii Adonicam sescenti sexaginta septem
NEH|7|19|filii Baggoaim duo milia sexaginta septem
NEH|7|20|filii Adin sescenti quinquaginta quinque
NEH|7|21|filii Ater filii Ezechiae nonaginta octo
NEH|7|22|filii Asem trecenti viginti octo
NEH|7|23|filii Besai trecenti viginti quattuor
NEH|7|24|filii Areph centum duodecim
NEH|7|25|filii Gabaon nonaginta quinque
NEH|7|26|viri Bethleem et Netupha centum octoginta octo
NEH|7|27|viri Anathoth centum viginti octo
NEH|7|28|viri Bethamoth quadraginta duo
NEH|7|29|viri Cariathiarim Cephira et Beroth septingenti quadraginta tres
NEH|7|30|viri Rama et Geba sescenti viginti unus
NEH|7|31|viri Machmas centum viginti duo
NEH|7|32|viri Bethel et Hai centum viginti tres
NEH|7|33|viri Nebo alterius quinquaginta duo
NEH|7|34|viri Helam alterius mille ducenti quinquaginta quattuor
NEH|7|35|filii Arem trecenti viginti
NEH|7|36|filii Hiericho trecenti quadraginta quinque
NEH|7|37|filii Lod Adid et Ono septingenti viginti unus
NEH|7|38|filii Senaa tria milia nongenti triginta
NEH|7|39|sacerdotes filii Idaia in domo Iosua nongenti septuaginta tres
NEH|7|40|filii Emmer mille quinquaginta duo
NEH|7|41|filii Phassur mille ducenti quadraginta septem
NEH|7|42|filii Arem mille decem et septem Levitae
NEH|7|43|filii Iosue et Cadmihel filiorum
NEH|7|44|Oduia septuaginta quattuor cantores
NEH|7|45|filii Asaph centum quadraginta octo
NEH|7|46|ianitores filii Sellum filii Ater filii Telmon filii Accub filii Atita filii Sobai centum triginta octo
NEH|7|47|Nathinnei filii Soa filii Asfa filii Tebaoth
NEH|7|48|filii Ceros filii Siaa filii Fado filii Lebana filii Agaba filii Selmon
NEH|7|49|filii Anan filii Geddel filii Gaer
NEH|7|50|filii Raaia filii Rasim filii Necoda
NEH|7|51|filii Gezem filii Aza filii Fasea
NEH|7|52|filii Besai filii Munim filii Nephusim
NEH|7|53|filii Becbuc filii Acupha filii Arur
NEH|7|54|filii Besloth filii Meida filii Arsa
NEH|7|55|filii Bercos filii Sisara filii Thema
NEH|7|56|filii Nesia filii Atipha
NEH|7|57|filii servorum Salomonis filii Sotai filii Sophereth filii Pherida
NEH|7|58|filii Iahala filii Dercon filii Geddel
NEH|7|59|filii Saphatia filii Athil filii Phocereth qui erat ortus ex Sabaim filio Amon
NEH|7|60|omnes Nathinnei et filii servorum Salomonis trecenti nonaginta duo
NEH|7|61|hii sunt autem qui ascenderunt de Thelmella Thelarsa Cherub Addon et Emmer et non potuerunt indicare domum patrum suorum et semen suum utrum ex Israhel essent
NEH|7|62|filii Dalaia filii Tobia filii Necoda sescenti quadraginta duo
NEH|7|63|et de sacerdotibus filii Abia filii Accos filii Berzellai qui accepit de filiabus Berzellai Galaditis uxorem et vocatus est nomine eorum
NEH|7|64|hii quaesierunt scripturam suam in censu et non invenerunt et eiecti sunt de sacerdotio
NEH|7|65|dixitque Athersatha eis ut non manducarent de sanctis sanctorum donec staret sacerdos doctus et eruditus
NEH|7|66|omnis multitudo quasi unus quadraginta duo milia sescenti sexaginta
NEH|7|67|absque servis et ancillis eorum qui erant septem milia trecenti triginta et septem et inter eos cantores et cantrices ducentae quadraginta quinque
NEH|7|68|
NEH|7|69|cameli quadringenti triginta quinque asini sex milia septingenti viginti
NEH|7|70|nonnulli autem de principibus familiarum dederunt in opus Athersatha dedit in thesaurum auri dragmas mille fialas quinquaginta tunicas sacerdotales quingentas triginta
NEH|7|71|et de principibus familiarum dederunt in thesaurum operis auri dragmas viginti milia et argenti minas duo milia ducentas
NEH|7|72|et quod dedit reliquus populus auri dragmas viginti milia et argenti minas duo milia et tunicas sacerdotales sexaginta septem
NEH|7|73|habitaverunt autem sacerdotes et Levitae et ianitores et cantores et reliquum vulgus et Nathinnei et omnis Israhel in civitatibus suis
NEH|8|1|et venerat mensis septimus filii autem Israhel erant in civitatibus suis congregatusque est omnis populus quasi vir unus ad plateam quae est ante portam Aquarum et dixerunt Ezrae scribae ut adferret librum legis Mosi quam praecepit Dominus Israheli
NEH|8|2|adtulit ergo Ezras sacerdos legem coram multitudine virorum et mulierum cunctisque qui poterant intellegere in die prima mensis septimi
NEH|8|3|et legit in eo aperte in platea quae erat ante portam Aquarum de mane usque ad mediam diem in conspectu virorum et mulierum et sapientium et aures omnis populi erant erectae ad librum
NEH|8|4|stetit autem Ezras scriba super gradum ligneum quem fecerat ad loquendum et steterunt iuxta eum Matthathia et Sema et Ania et Uria et Helcia et Maasia ad dextram eius et ad sinistram Phadaia Misahel et Melchia et Asum et Asephdana Zaccharia et Mosollam
NEH|8|5|et aperuit Ezras librum coram omni populo super universum quippe populum eminebat et cum aperuisset eum stetit omnis populus
NEH|8|6|et benedixit Ezras Domino Deo magno et respondit omnis populus amen amen elevans manus suas et incurvati sunt et adoraverunt Deum proni in terram
NEH|8|7|porro Hiesue et Baani et Serebia Iamin Accub Septhai Odia Maasia Celita Azarias Iozabed Anam Phalaia Levitae silentium faciebant in populo ad audiendam legem populus autem stabat in gradu suo
NEH|8|8|et legerunt in libro legis Dei distincte et adposite ad intellegendum et intellexerunt cum legeretur
NEH|8|9|dixit autem Neemias ipse est Athersatha et Ezras sacerdos scriba et Levitae interpretantes universo populo dies sanctificatus est Domino Deo nostro nolite lugere et nolite flere flebat enim omnis populus cum audiret verba legis
NEH|8|10|et dixit eis ite comedite pinguia et bibite mulsum et mittite partes ei qui non praeparavit sibi quia sanctus dies Domini est et nolite contristari gaudium enim Domini est fortitudo nostra
NEH|8|11|Levitae autem silentium faciebant in omni populo dicentes tacete quia dies sanctus est et nolite dolere
NEH|8|12|abiit itaque omnis populus ut comederet et biberet et mitteret partes et faceret laetitiam magnam quia intellexerant verba quae docuerat eos
NEH|8|13|et in die secundo congregati sunt principes familiarum universi populi sacerdotes et Levitae ad Ezram scribam ut interpretaretur eis verba legis
NEH|8|14|et invenerunt scriptum in lege praecepisse Dominum in manu Mosi ut habitent filii Israhel in tabernaculis in die sollemni mense septimo
NEH|8|15|et ut praedicent et divulgent vocem in universis urbibus suis et in Hierusalem dicentes egredimini in montem et adferte frondes olivae et frondes ligni pulcherrimi frondes myrti et ramos palmarum et frondes ligni nemorosi ut fiant tabernacula sicut scriptum est
NEH|8|16|et egressus est populus et adtulerunt feceruntque sibi tabernacula unusquisque in domate suo et in atriis suis et in atriis domus Dei et in platea portae Aquarum et in platea portae Ephraim
NEH|8|17|fecit ergo universa ecclesia eorum qui redierant de captivitate tabernacula et habitaverunt in tabernaculis non enim fecerant a diebus Iosue filii Nun taliter filii Israhel usque ad diem illum et fuit laetitia magna nimis
NEH|8|18|legit autem in libro legis Dei per dies singulos a die primo usque ad diem novissimum et fecerunt sollemnitatem septem diebus et in die octavo collectum iuxta ritum
NEH|9|1|in die autem vicesimo quarto mensis huius convenerunt filii Israhel in ieiunio et in saccis et humus super eos
NEH|9|2|et separatum est semen filiorum Israhel ab omni filio alienigena et steterunt et confitebantur peccata sua et iniquitates patrum suorum
NEH|9|3|et consurrexerunt ad standum et legerunt in volumine legis Domini Dei sui quater in die et quater confitebantur et adorabant Dominum Deum suum
NEH|9|4|surrexit autem super gradum Levitarum Iosue et Bani Cedmihel Sebnia Bani Sarebias Bani Chanani et inclamaverunt voce magna Dominum Deum suum
NEH|9|5|et dixerunt Levitae Iosue et Cedmihel Bonni Asebia Serebia Odoia Sebna Fataia surgite benedicite Domino Deo vestro ab aeterno usque in aeternum et benedicant nomini gloriae tuae excelso in omni benedictione et laude
NEH|9|6|tu ipse Domine solus tu fecisti caelum caelum caelorum et omnem exercitum eorum terram et universa quae in ea sunt maria et omnia quae in eis sunt et tu vivificas omnia haec et exercitus caeli te adorat
NEH|9|7|tu ipse Domine Deus qui elegisti Abram et eduxisti eum de igne Chaldeorum et posuisti nomen eius Abraham
NEH|9|8|et invenisti cor eius fidele coram te et percussisti cum eo foedus ut dares ei terram Chananei Chetthei Amorrei et Ferezei et Iebusei et Gergesei ut dares semini eius et implesti verba tua quoniam iustus es
NEH|9|9|et vidisti adflictionem patrum nostrorum in Aegypto clamoremque eorum audisti super mare Rubrum
NEH|9|10|et dedisti signa et portenta in Pharao et in universis servis eius et in omni populo terrae illius cognovisti enim quia superbe egerant contra eos et fecisti tibi nomen sicut et in hac die
NEH|9|11|et mare divisisti ante eos et transierunt per medium maris in sicca persecutores autem eorum proiecisti in profundum quasi lapidem in aquas validas
NEH|9|12|et in columna nubis ductor eorum fuisti per diem et in columna ignis per noctem ut appareret eis via per quam ingrediebantur
NEH|9|13|ad montem quoque Sinai descendisti et locutus es cum eis de caelo et dedisti eis iudicia recta et legem veritatis caerimonias et praecepta bona
NEH|9|14|et sabbatum sanctificatum tuum ostendisti eis et mandata et caerimonias et legem praecepisti eis in manu Mosi servi tui
NEH|9|15|panem quoque de caelo dedisti eis in fame eorum et aquam de petra eduxisti eis sitientibus et dixisti eis ut ingrederentur et possiderent terram super quam levasti manum tuam ut traderes eis
NEH|9|16|ipsi vero et patres nostri superbe egerunt et induraverunt cervices suas et non audierunt mandata tua
NEH|9|17|et noluerunt audire et non sunt recordati mirabilium tuorum quae feceras eis et induraverunt cervices suas et dederunt caput ut converterentur ad servitutem suam quasi per contentionem tu autem Deus propitius clemens et misericors longanimis et multae miserationis non dereliquisti eos
NEH|9|18|et quidem cum fecissent sibi vitulum conflatilem et dixissent iste est Deus tuus qui eduxit te de Aegypto feceruntque blasphemias magnas
NEH|9|19|tu autem in misericordiis tuis multis non dimisisti eos in deserto columna nubis non recessit ab eis per diem ut duceret eos in via et columna ignis in nocte ut ostenderet eis iter per quod ingrederentur
NEH|9|20|et spiritum tuum bonum dedisti qui doceret eos et manna tuum non prohibuisti ab ore eorum et aquam dedisti eis in siti
NEH|9|21|quadraginta annis pavisti eos in deserto nihilque eis defuit vestimenta eorum non inveteraverunt et pedes eorum non sunt adtriti
NEH|9|22|et dedisti eis regna et populos et partitus es eis sortes et possederunt terram Seon et terram regis Esebon et terram Og regis Basan
NEH|9|23|et filios eorum multiplicasti sicut stellas caeli et adduxisti eos ad terram de qua dixeras patribus eorum ut ingrederentur et possiderent
NEH|9|24|et venerunt filii et possederunt terram et humiliasti coram eis habitatores terrae Chananeos et dedisti eos in manu eorum et reges eorum et populos terrae ut facerent eis sicut placebat illis
NEH|9|25|ceperunt itaque urbes munitas et humum pinguem et possederunt domos plenas cunctis bonis cisternas ab aliis fabricatas vineas et oliveta et ligna pomifera multa et comederunt et saturati sunt et inpinguati sunt et abundavere deliciis in bonitate tua magna
NEH|9|26|provocaverunt autem te ad iracundiam et recesserunt a te et proiecerunt legem tuam post terga sua et prophetas tuos occiderunt qui contestabantur eos ut reverterentur ad te feceruntque blasphemias grandes
NEH|9|27|et dedisti eos in manu hostium suorum et adflixerunt eos et in tempore tribulationis suae clamaverunt ad te et tu de caelo audisti et secundum miserationes tuas multas dedisti eis salvatores qui salvaverunt eos de manu hostium suorum
NEH|9|28|cumque requievissent reversi sunt ut facerent malum in conspectu tuo et dereliquisti eos in manu inimicorum suorum et possederunt eos conversique sunt et clamaverunt ad te tu autem de caelo audisti et liberasti eos in misericordiis tuis multis temporibus
NEH|9|29|et contestatus es eos ut reverterentur ad legem tuam ipsi vero superbe egerunt et non audierunt mandata tua et in iudiciis tuis peccaverunt quae faciet homo et vivet in eis et dederunt umerum recedentem et cervicem suam induraverunt nec audierunt
NEH|9|30|et protraxisti super eos annos multos et contestatus es eos in spiritu tuo per manum prophetarum tuorum et non audierunt et tradidisti eos in manu populorum terrarum
NEH|9|31|in misericordiis autem tuis plurimis non fecisti eos in consumptione nec dereliquisti eos quoniam Deus miserationum et clemens tu es
NEH|9|32|nunc itaque Deus noster Deus magne fortis et terribilis custodiens pactum et misericordiam ne avertas a facie tua omnem laborem qui invenit nos reges nostros principes nostros et sacerdotes nostros prophetas nostros et patres nostros et omnem populum tuum a diebus regis Assur usque in diem hanc
NEH|9|33|et tu iustus in omnibus quae venerunt super nos quia veritatem fecisti nos autem impie egimus
NEH|9|34|reges nostri principes nostri sacerdotes nostri et patres nostri non fecerunt legem tuam et non adtenderunt mandata tua et testimonia tua quae testificatus es in eis
NEH|9|35|et ipsi in regnis suis bonis et in bonitate tua multa quam dederas eis et in terra latissima et pingui quam tradideras in conspectu eorum non servierunt tibi nec reversi sunt ab studiis suis pessimis
NEH|9|36|ecce nos ipsi hodie servi sumus et terram quam dedisti patribus nostris ut comederent panem eius et quae bona sunt eius et nos ipsi servi sumus in ea
NEH|9|37|et fruges eius multiplicantur regibus quos posuisti super nos propter peccata nostra et in corporibus nostris dominantur et in iumentis nostris secundum voluntatem suam et in tribulatione magna sumus
NEH|9|38|super omnibus ergo his nos ipsi percutimus foedus et scribimus et signant principes nostri Levitae nostri et sacerdotes nostri
NEH|10|1|signatores autem fuerunt Neemias Athersatha filius Achelai et Sedecias
NEH|10|2|Saraias Azarias Hieremias
NEH|10|3|Phessur Amaria Melchia
NEH|10|4|Attus Sebenia Melluc
NEH|10|5|Arem Mermuth Obdias
NEH|10|6|Danihel Genton Baruch
NEH|10|7|Mosollam Abia Miamin
NEH|10|8|Mazia Belga Semaia hii sacerdotes
NEH|10|9|porro Levitae Iosue filius Azaniae Bennui de filiis Enadad Cedmihel
NEH|10|10|et fratres eorum Sechenia Odevia Celita Phalaia Anan
NEH|10|11|Micha Roob Asebia
NEH|10|12|Zacchur Serebia Sabania
NEH|10|13|Odia Bani Baninu
NEH|10|14|capita populi Pheros Phaethmoab Helam Zethu Bani
NEH|10|15|Bonni Azgad Bebai
NEH|10|16|Adonia Beggoai Adin
NEH|10|17|Ater Ezechia Azur
NEH|10|18|Odevia Asum Besai
NEH|10|19|Ares Anathoth Nebai
NEH|10|20|Mecphia Mosollam Azir
NEH|10|21|Mesizabel Sadoc Ieddua
NEH|10|22|Felthia Anan Ania
NEH|10|23|Osee Anania Asub
NEH|10|24|Aloes Phaleam Sobec
NEH|10|25|Reum Asebna Madsia
NEH|10|26|et Haia Hanam Anan
NEH|10|27|Melluc Arem Baana
NEH|10|28|et reliqui de populo sacerdotes Levitae ianitores et cantores Nathinnei et omnes qui se separaverunt de populis terrarum ad legem Dei uxores eorum filii eorum et filiae eorum
NEH|10|29|omnis qui poterat sapere spondentes pro fratribus suis optimates eorum et qui veniebant ad pollicendum et iurandum ut ambularent in lege Dei quam dederat in manu Mosi servi Dei ut facerent et custodirent universa mandata Domini Dei nostri et iudicia eius et caerimonias eius
NEH|10|30|et ut non daremus filias nostras populo terrae et filias eorum non acciperemus filiis nostris
NEH|10|31|populi quoque terrae qui inportant venalia et omnia ad usum per diem sabbati ut vendant non accipiemus ab eis in sabbato et in die sanctificata et dimittemus annum septimum et exactionem universae manus
NEH|10|32|et statuemus super nos praecepta ut demus tertiam partem sicli per annum ad opus domus Dei nostri
NEH|10|33|ad panes propositionis et ad sacrificium sempiternum et in holocaustum sempiternum in sabbatis in kalendis in sollemnitatibus et in sanctificatis et pro peccato ut exoretur pro Israhel et in omnem usum domus Dei nostri
NEH|10|34|sortes ergo misimus super oblatione lignorum inter sacerdotes et Levitas et populos ut inferrentur in domum Dei nostri per domos patrum nostrorum per tempora a temporibus anni usque ad annum ut arderent super altare Domini Dei nostri sicut scriptum est in lege Mosi
NEH|10|35|et ut adferremus primogenita terrae nostrae et primitiva universi fructus omnis ligni ab anno in annum in domo Domini
NEH|10|36|et primitiva filiorum nostrorum et pecorum nostrorum sicut scriptum est in lege et primitiva boum nostrorum et ovium nostrarum ut offerrentur in domo Dei nostri sacerdotibus qui ministrant in domo Dei nostri
NEH|10|37|et primitias ciborum nostrorum et libaminum nostrorum et poma omnis ligni vindemiae quoque et olei adferemus sacerdotibus ad gazofilacium Dei nostri et decimam partem terrae nostrae Levitis ipsi Levitae decimas accipient ex omnibus civitatibus operum nostrorum
NEH|10|38|erit autem sacerdos filius Aaron cum Levitis in decimis Levitarum et Levitae offerent decimam partem decimae suae in domum Dei nostri ad gazofilacium in domo thesauri
NEH|10|39|ad gazofilacium enim deportabunt filii Israhel et filii Levi primitias frumenti vini et olei et ibi erunt vasa sanctificata et sacerdotes et cantores et ianitores et ministri et non dimittemus domum Dei nostri
NEH|11|1|habitaverunt autem principes populi in Hierusalem reliqua vero plebs misit sortem ut tollerent unam partem de decem qui habitaturi essent in Hierusalem in civitate sancta novem vero partes in civitatibus
NEH|11|2|benedixit autem populus omnibus viris qui se sponte obtulerunt ut habitarent in Hierusalem
NEH|11|3|hii sunt itaque principes provinciae qui habitaverunt in Hierusalem et in civitatibus Iuda habitavit unusquisque in possessione sua in urbibus suis Israhel sacerdotes Levitae Nathinnei et filii servorum Salomonis
NEH|11|4|et in Hierusalem habitaverunt de filiis Iuda et de filiis Beniamin de filiis Iuda Athaias filius Aziam filii Zacchariae filii Amariae filii Saphatia filii Malelehel de filiis Phares
NEH|11|5|Imaasia filius Baruch filius Coloza filius Azia filius Adaia filius Ioiarib filius Zacchariae filius Silonites
NEH|11|6|omnes filii Phares qui habitaverunt in Hierusalem quadringenti sexaginta octo viri fortes
NEH|11|7|hii sunt autem filii Beniamin Sellum filius Mosollam filius Ioed filius Phadaia filius Colaia filius Masia filius Ethehel filius Isaia
NEH|11|8|et post eum Gabbai Sellai nongenti viginti octo
NEH|11|9|et Iohel filius Zechri praepositus eorum et Iuda filius Sennua super civitatem secundus
NEH|11|10|et de sacerdotibus Idaia filius Ioarib Iachin
NEH|11|11|Saraia filius Elcia filius Mesollam filius Sadoc filius Meraioth filius Ahitub princeps domus Dei
NEH|11|12|et fratres eorum facientes opera templi octingenti viginti duo et Adaia filius Ieroam filius Felelia filius Amsi filius Zacchariae filius Phessur filius Melchiae
NEH|11|13|et fratres eius principes patrum ducenti quadraginta duo et Amassai filius Azrihel filius Aazi filius Mosollamoth filius Emmer
NEH|11|14|et fratres eorum potentes nimis centum viginti octo et praepositus eorum Zabdihel filius potentium
NEH|11|15|et de Levitis Sebenia filius Asob filius Azaricam filius Asabia filius Boni
NEH|11|16|et Sabathai et Iozabed super opera quae erant forinsecus in domo Dei a principibus Levitarum
NEH|11|17|et Mathania filius Micha filius Zebdaei filius Asaph princeps ad laudandum et confitendum in oratione et Becbecia secundus de fratribus eius et Abda filius Sammua filius Galal filius Idithun
NEH|11|18|omnes Levitae in civitate sancta ducenti octoginta quattuor
NEH|11|19|et ianitores Accob Telmon et fratres eorum qui custodiebant ostia centum septuaginta duo
NEH|11|20|et reliqui ex Israhel sacerdotes et Levitae in universis civitatibus Iuda unusquisque in possessione sua
NEH|11|21|et Nathinnei qui habitabant in Ofel et Siaha et Gaspha de Nathinneis
NEH|11|22|et episcopus Levitarum in Hierusalem Azzi filius Bani filius Asabiae filius Matthaniae filius Michae de filiis Asaph cantores in ministerio domus Dei
NEH|11|23|praeceptum quippe regis super eos erat et ordo in cantoribus per dies singulos
NEH|11|24|et Fataia filius Mesezebel de filiis Zera filii Iuda in manu regis iuxta omne verbum populi
NEH|11|25|et in domibus per omnes regiones eorum de filiis Iuda habitaverunt in Cariatharbe et in filiabus eius et in Dibon et in filiabus eius et in Capsel et in viculis eius
NEH|11|26|et in Iesue et in Molada et in Bethfaleth
NEH|11|27|et in Asersual et in Bersabee et in filiabus eius
NEH|11|28|et in Siceleg et in Mochona et in filiabus eius
NEH|11|29|et in Ainremmon et in Sara et in Irimuth
NEH|11|30|Zanoa Odollam et villis earum Lachis et regionibus eius Azeca et filiabus eius et manserunt in Bersabee usque ad vallem Ennom
NEH|11|31|filii autem Beniamin a Geba Mechmas et Aia et Bethel et filiabus eius
NEH|11|32|Anathoth Nob Anania
NEH|11|33|Asor Rama Getthaim
NEH|11|34|Adid Seboim Neballa Loth
NEH|11|35|et Ono valle Artificum
NEH|11|36|et de Levitis partitiones Iuda et Beniamin
NEH|12|1|hii autem sacerdotes et Levitae qui ascenderunt cum Zorobabel filio Salathihel et Iosue Saraia Hieremias Ezra
NEH|12|2|Amaria Melluch Attus
NEH|12|3|Sechenia Reum Meremuth
NEH|12|4|Addo Genthon Abia
NEH|12|5|Miamin Madia Belga
NEH|12|6|Semaia et Ioarib Idaia Sellum Amoc Elceia
NEH|12|7|Idaia isti principes sacerdotum et fratres eorum in diebus Iosue
NEH|12|8|porro Levitae Iesua Bennui Cedmihel Sarabia Iuda Mathanias super hymnos ipsi et fratres eorum
NEH|12|9|et Becbecia atque et Hanni fratres eorum unusquisque in officio suo
NEH|12|10|Hiesue autem genuit Ioachim et Ioachim genuit Eliasib et Eliasib genuit Ioiada
NEH|12|11|et Ioiada genuit Ionathan et Ionathan genuit Ieddoa
NEH|12|12|in diebus autem Ioachim erant sacerdotes principes familiarum Saraiae Amaria Hieremiae Anania
NEH|12|13|Ezrae Mosollam Amariae Iohanan
NEH|12|14|Milico Ionathan Sebeniae Ioseph
NEH|12|15|Arem Edna Maraioth Elci
NEH|12|16|Addaiae Zaccharia Genthon Mosollam
NEH|12|17|Abiae Zecheri Miamin et Moadiae Felti
NEH|12|18|Belgae Sammua Semaiae Ionathan
NEH|12|19|Ioiarib Matthanai Iadaiae Azzi
NEH|12|20|Sellaiae Celai Amoc Eber
NEH|12|21|Elciae Asebia Idaiae Nathanahel
NEH|12|22|Levitae in diebus Eliasib et Ioiada et Ionan et Ieddoa scripti principes familiarum et sacerdotes in regno Darii Persae
NEH|12|23|filii Levi principes familiarum scripti in libro verborum dierum et usque ad dies Ionathan filii Eliasib
NEH|12|24|et principes Levitarum Asebia Serebia et Iesue filius Cedmihel et fratres eorum per vices suas ut laudarent et confiterentur iuxta praeceptum David viri Dei et observarent aeque per ordinem
NEH|12|25|Matthania et Becbecia Obedia Mosollam Thelmon Accub custodes portarum et vestibulorum ante portas
NEH|12|26|hii in diebus Ioachim filii Iesue filii Iosedech et in diebus Neemiae ducis et Ezrae sacerdotis scribaeque
NEH|12|27|in dedicatione autem muri Hierusalem requisierunt Levitas de omnibus locis suis ut adducerent eos in Hierusalem et facerent dedicationem et laetitiam in actione gratiarum et in cantico in cymbalis psalteriis et citharis
NEH|12|28|congregati sunt ergo filii cantorum et de campestribus circa Hierusalem et de villis Netuphati
NEH|12|29|et de domo Galgal et de regionibus Geba et Azmaveth quoniam villas aedificaverunt sibi cantores in circuitu Hierusalem
NEH|12|30|et mundati sunt sacerdotes et Levitae et mundaverunt populum et portas et murum
NEH|12|31|ascendere autem feci principes Iuda super murum et statui duos choros laudantium magnos et ierunt ad dexteram super murum ad portam Sterquilinii
NEH|12|32|et ivit post eos Osaias et media pars principum Iuda
NEH|12|33|et Azarias Ezras et Mosollam Iuda et Beniamin et Semeia et Hieremia
NEH|12|34|et de filiis sacerdotum in tubis Zaccharias filius Ionathan filius Semeiae filius Mathaniae filius Michaiae filius Zecchur filius Asaph
NEH|12|35|et fratres eius Semeia et Azarel Malalai Galalai Maai Nathanel et Iuda et Anani in vasis cantici David viri Dei et Ezras scriba ante eos in porta Fontis
NEH|12|36|et contra eos ascenderunt in gradibus civitatis David in ascensu muri super domum David et usque ad portam Aquarum ad orientem
NEH|12|37|et chorus secundus gratias referentium ibat ex adverso et ego post eum et media pars populi super murum et super turrem Furnorum et usque ad murum latissimum
NEH|12|38|et super portam Ephraim et super portam Antiquam et super portam Piscium et turrem Ananehel et turrem Ema et usque ad portam Gregis et steterunt in porta Custodiae
NEH|12|39|steteruntque duo chori laudantium in domo Dei et ego et dimidia pars magistratuum mecum
NEH|12|40|et sacerdotes Eliachim Maasia Miniamin Michea Elioenai Zaccharia Anania in tubis
NEH|12|41|et Maasia et Semea et Eleazar et Azi et Iohanan et Melchia et Elam et Ezer et clare cecinerunt cantores et Iezraia praepositus
NEH|12|42|et immolaverunt in die illa victimas magnas et laetati sunt Deus enim laetificaverat eos laetitia magna sed et uxores eorum et liberi gavisi sunt et audita est laetitia Hierusalem procul
NEH|12|43|recensuerunt quoque in die illa viros super gazofilacia thesauri ad libamina et ad primitias et ad decimas ut introferrent per eos principes civitatis in decore gratiarum actionis sacerdotes et Levitas quia laetatus est Iuda in sacerdotibus et Levitis adstantibus
NEH|12|44|et custodierunt observationem Dei sui et observationem expiationis et cantores et ianitores iuxta praeceptum David et Salomonis filii eius
NEH|12|45|quia in diebus David et Asaph ab exordio erant principes constituti cantorum in carmine laudantium et confitentium Deo
NEH|12|46|et omnis Israhel in diebus Zorobabel et in diebus Neemiae dabat partes cantoribus et ianitoribus per dies singulos et sanctificabant Levitas et Levitae sanctificabant filios Aaron
NEH|13|1|in die autem illo lectum est in volumine Mosi audiente populo et inventum est scriptum in eo quod non debeat introire Ammanites et Moabites in ecclesiam Dei usque in aeternum
NEH|13|2|eo quod non occurrerint filiis Israhel cum pane et aqua et conduxerint adversum eum Balaam ad maledicendum ei et convertit Deus noster maledictionem in benedictionem
NEH|13|3|factum est autem cum audissent legem separaverunt omnem alienigenam ab Israhel
NEH|13|4|et super hoc erat Eliasib sacerdos qui fuerat positus in gazofilacio domus Dei nostri et proximus Tobiae
NEH|13|5|fecit ergo sibi gazofilacium grande et ibi erant ante eum reponentes munera et tus et vasa et decimam frumenti et vini et olei partes Levitarum et cantorum et ianitorum et primitias sacerdotales
NEH|13|6|in omnibus autem his non fui in Hierusalem quia in anno tricesimo secundo Artarxersis regis Babylonis veni ad regem et in fine dierum rogavi regem
NEH|13|7|et veni in Hierusalem et intellexi malum quod fecerat Eliasib Tobiae ut faceret ei thesaurum in vestibulis domus Dei
NEH|13|8|et malum mihi visum est valde et proieci vasa domus Tobiae foras de gazofilacio
NEH|13|9|praecepique et mundaverunt gazofilacia et rettuli ibi vasa domus Dei sacrificium et tus
NEH|13|10|et cognovi quoniam partes Levitarum non fuissent datae et fugisset unusquisque in regionem suam de Levitis et de cantoribus et de his qui ministrabant
NEH|13|11|et egi causam adversus magistratus et dixi quare dereliquimus domum Dei et congregavi eos et feci stare in stationibus suis
NEH|13|12|et omnis Iuda adportabat decimam frumenti et vini et olei in horrea
NEH|13|13|et constituimus super horrea Selemiam sacerdotem et Sadoc scribam et Phadaiam de Levitis et iuxta eos Anan filium Zacchur filium Matthaniae quoniam fideles conprobati sunt et ipsis creditae sunt partes fratrum suorum
NEH|13|14|memento mei Deus meus pro hoc et ne deleas miserationes meas quas feci in domo Dei mei et in caerimoniis eius
NEH|13|15|in diebus illis vidi in Iuda calcabant torcularia in sabbato portantes acervos et onerantes super asinos vinum et uvas et ficus et omne onus et inferentes Hierusalem in die sabbati et contestatus sum ut in die qua vendere liceret venderent
NEH|13|16|et Tyrii habitaverunt in ea inferentes pisces et omnia venalia et vendebant in sabbatis filiis Iuda et in Hierusalem
NEH|13|17|et obiurgavi optimates Iuda et dixi eis quae est res haec mala quam vos facitis et profanatis diem sabbati
NEH|13|18|numquid non haec fecerunt patres nostri et adduxit Deus noster super nos omne malum hoc et super civitatem hanc et vos additis iracundiam super Israhel violando sabbatum
NEH|13|19|factum est itaque cum quievissent portae Hierusalem die sabbati dixi et cluserunt ianuas et praecepi ut non aperirent eas usque post sabbatum et de pueris meis constitui super portas ut nullus inferret onus in die sabbati
NEH|13|20|et manserunt negotiatores et vendentes universa venalia foris Hierusalem semel et bis
NEH|13|21|et contestatus sum eos et dixi eis quare manetis ex adverso muri si secundo hoc feceritis manum mittam in vos itaque ex tempore illo non venerunt in sabbato
NEH|13|22|dixi quoque Levitis ut mundarentur et venirent ad custodiendas portas et sanctificandum diem sabbati et pro hoc ergo memento mei Deus meus et parce mihi secundum multitudinem miserationum tuarum
NEH|13|23|sed et in diebus illis vidi Iudaeos ducentes uxores azotias ammanitidas et moabitidas
NEH|13|24|et filii eorum ex media parte loquebantur azotice et nesciebant loqui iudaice et loquebantur iuxta linguam populi et populi
NEH|13|25|et obiurgavi eos et maledixi et cecidi ex ipsis viros et decalvavi eos et adiuravi in Deo ut non darent filias suas filiis eorum et non acciperent de filiabus eorum filiis suis et sibimet ipsis dicens
NEH|13|26|numquid non in huiuscemodi re peccavit Salomon rex Israhel et certe in gentibus multis non erat rex similis ei et dilectus Deo suo erat et posuit eum Deus regem super omnem Israhel et ipsum ergo ad peccatum duxerunt mulieres alienigenae
NEH|13|27|numquid et nos inoboedientes faciemus omne malum grande hoc ut praevaricemur in Deo nostro et ducamus uxores peregrinas
NEH|13|28|de filiis autem Ioiada filii Eliasib sacerdotis magni gener erat Sanaballat Horonitis quem fugavi a me
NEH|13|29|recordare Domine Deus meus adversum eos qui polluunt sacerdotium iusque sacerdotale et leviticum
NEH|13|30|igitur mundavi eos ab omnibus alienigenis et constitui ordines sacerdotum et Levitarum unumquemque in ministerio suo
NEH|13|31|et in oblatione lignorum in temporibus constitutis et in primitiis memento mei Deus meus in bonum
