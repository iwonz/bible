HOS|1|1|verbum Domini quod factum est ad Osee filium Beeri in diebus Oziae Ioatham Ahaz Ezechiae regum Iuda et in diebus Hieroboam filii Ioas regis Israhel
HOS|1|2|principium loquendi Dominum in Osee et dixit Dominus ad Osee vade sume tibi uxorem fornicationum et filios fornicationum quia fornicans fornicabitur terra a Domino
HOS|1|3|et abiit et accepit Gomer filiam Debelaim et concepit et peperit filium
HOS|1|4|et dixit Dominus ad eum voca nomen eius Hiezrahel quoniam adhuc modicum et visitabo sanguinem Hiezrahel super domum Hieu et quiescere faciam regnum domus Israhel
HOS|1|5|et in illa die conteram arcum Israhel in valle Hiezrahel
HOS|1|6|et concepit adhuc et peperit filiam et dixit ei voca nomen eius Absque misericordia quia non addam ultra misereri domui Israhel sed oblivione obliviscar eorum
HOS|1|7|et domui Iuda miserebor et salvabo eos in Domino Deo suo et non salvabo eos in arcu et gladio et in bello et in equis et in equitibus
HOS|1|8|et ablactavit eam quae erat absque misericordia et concepit et peperit filium
HOS|1|9|et dixit voca nomen eius Non populus meus quia vos non populus meus et ego non ero vester
HOS|1|10|et erit numerus filiorum Israhel quasi harena maris quae sine mensura est et non numerabitur et erit in loco ubi dicetur eis non populus meus vos dicetur eis filii Dei viventis
HOS|1|11|et congregabuntur filii Iuda et filii Israhel pariter et ponent sibimet caput unum et ascendent de terra quia magnus dies Hiezrahel
HOS|2|1|dicite fratribus vestris Populus meus et sorori vestrae Misericordiam consecuta
HOS|2|2|iudicate matrem vestram iudicate quoniam ipsa non uxor mea et ego non vir eius auferat fornicationes suas a facie sua et adulteria sua de medio uberum suorum
HOS|2|3|ne forte expoliem eam nudam et statuam eam secundum diem nativitatis suae et ponam eam quasi solitudinem et statuam eam velut terram inviam et interficiam eam siti
HOS|2|4|et filiorum illius non miserebor quoniam filii fornicationum sunt
HOS|2|5|quia fornicata est mater eorum confusa est quae concepit eos quia dixit vadam post amatores meos qui dant panes mihi et aquas meas lanam meam et linum meum oleum meum et potum meum
HOS|2|6|propter hoc ecce ego sepiam viam tuam spinis et sepiam eam maceria et semitas suas non inveniet
HOS|2|7|et sequetur amatores suos et non adprehendet eos et quaeret eos et non inveniet et dicet vadam et revertar ad virum meum priorem quia bene mihi erat tunc magis quam nunc
HOS|2|8|et haec nescivit quia ego dedi ei frumentum et vinum et oleum et argentum multiplicavi ei et aurum quae fecerunt Baal
HOS|2|9|idcirco convertar et sumam frumentum meum in tempore suo et vinum meum in tempore suo et liberabo lanam meam et linum meum quae operiebant ignominiam eius
HOS|2|10|et nunc revelabo stultitiam eius in oculis amatorum eius et vir non eruet eam de manu mea
HOS|2|11|et cessare faciam omne gaudium eius sollemnitatem eius neomeniam eius sabbatum eius et omnia festa tempora eius
HOS|2|12|et corrumpam vineam eius et ficum eius de quibus dixit mercedes hae meae sunt quas dederunt mihi amatores mei et ponam eam in saltu et comedet illam bestia agri
HOS|2|13|et visitabo super eam dies Baalim quibus accendebat incensum et ornabatur inaure sua et monili suo et ibat post amatores suos et mei obliviscebatur dicit Dominus
HOS|2|14|propter hoc ecce ego lactabo eam et ducam eam in solitudinem et loquar ad cor eius
HOS|2|15|et dabo ei vinitores eius ex eodem loco et vallem Achor ad aperiendam spem et canet ibi iuxta dies iuventutis suae et iuxta dies ascensionis suae de terra Aegypti
HOS|2|16|et erit in die illo ait Dominus vocabit me Vir meus et non vocabit me ultra Baali
HOS|2|17|et auferam nomina Baalim de ore eius et non recordabitur ultra nominis eorum
HOS|2|18|et percutiam eis foedus in die illa cum bestia agri et cum volucre caeli et cum reptili terrae et arcum et gladium et bellum conteram de terra et dormire eos faciam fiducialiter
HOS|2|19|et sponsabo te mihi in sempiternum et sponsabo te mihi in iustitia et iudicio et in misericordia et miserationibus
HOS|2|20|et sponsabo te mihi in fide et scies quia ego Dominus
HOS|2|21|et erit in illa die exaudiam dicit Dominus exaudiam caelos et illi exaudient terram
HOS|2|22|et terra exaudiet triticum et vinum et oleum et haec exaudient Hiezrahel
HOS|2|23|et seminabo eam mihi in terram et miserebor eius quae fuit absque misericordia
HOS|2|24|et dicam non populo meo populus meus tu et ipse dicet Dominus meus es tu
HOS|3|1|et dixit Dominus ad me adhuc vade dilige mulierem dilectam amico et adulteram sicut diligit Dominus filios Israhel et ipsi respectant ad deos alienos et diligunt vinacea uvarum
HOS|3|2|et fodi eam mihi quindecim argenteis et choro hordei et dimidio choro hordei
HOS|3|3|et dixi ad eam dies multos expectabis me non fornicaberis et non eris viro sed et ego expectabo te
HOS|3|4|quia dies multos sedebunt filii Israhel sine rege et sine principe et sine sacrificio et sine altari et sine ephod et sine therafin
HOS|3|5|et post haec revertentur filii Israhel et quaerent Dominum Deum suum et David regem suum et pavebunt ad Dominum et ad bonum eius in novissimo dierum
HOS|4|1|audite verbum Domini filii Israhel quia iudicium Domino cum habitatoribus terrae non est enim veritas et non est misericordia et non est scientia Dei in terra
HOS|4|2|maledictum et mendacium et homicidium et furtum et adulterium inundaverunt et sanguis sanguinem tetigit
HOS|4|3|propter hoc lugebit terra et infirmabitur omnis qui habitat in ea in bestia agri et in volucre caeli sed et pisces maris congregabuntur
HOS|4|4|verumtamen unusquisque non iudicet et non arguatur vir populus enim tuus sicut hii qui contradicunt sacerdoti
HOS|4|5|et corrues hodie et corruet etiam propheta tecum nocte tacere feci matrem tuam
HOS|4|6|conticuit populus meus eo quod non habuerit scientiam quia tu scientiam reppulisti repellam te ne sacerdotio fungaris mihi et oblita es legis Dei tui obliviscar filiorum tuorum et ego
HOS|4|7|secundum multitudinem eorum sic peccaverunt mihi gloriam eorum in ignominiam commutabo
HOS|4|8|peccata populi mei comedent et ad iniquitatem eorum sublevabunt animas eorum
HOS|4|9|et erit sicut populus sic sacerdos et visitabo super eum vias eius et cogitationes eius reddam ei
HOS|4|10|et comedent et non saturabuntur fornicati sunt et non cessaverunt quoniam Dominum reliquerunt in non custodiendo
HOS|4|11|fornicatio et vinum et ebrietas aufert cor
HOS|4|12|populus meus in ligno suo interrogavit et baculus eius adnuntiavit ei spiritus enim fornicationum decepit eos et fornicati sunt a Deo suo
HOS|4|13|super capita montium sacrificabant et super colles accendebant thymiama subtus quercum et populum et terebinthum quia bona erat umbra eius ideo fornicabuntur filiae vestrae et sponsae vestrae adulterae erunt
HOS|4|14|non visitabo super filias vestras cum fuerint fornicatae et super sponsas vestras cum adulteraverint quoniam ipsi cum meretricibus versabantur et cum effeminatis sacrificabant et populus non intellegens vapulabit
HOS|4|15|si fornicaris tu Israhel non delinquat saltim Iuda et nolite ingredi in Galgala et ne ascenderitis in Bethaven neque iuraveritis vivit Dominus
HOS|4|16|quoniam sicut vacca lasciviens declinavit Israhel nunc pascet eos Dominus quasi agnum in latitudine
HOS|4|17|particeps idolorum Ephraim dimitte eum
HOS|4|18|separatum est convivium eorum fornicatione fornicati sunt dilexerunt adferre ignominiam protectores eius
HOS|4|19|ligavit spiritus eam in alis suis et confundentur a sacrificiis suis
HOS|5|1|audite hoc sacerdotes et adtendite domus Israhel et domus regis auscultate quia vobis iudicium est quoniam laqueus facti estis speculationi et rete expansum super Thabor
HOS|5|2|et victimas declinastis in profundum et ego eruditor omnium eorum
HOS|5|3|ego scio Ephraim et Israhel non est absconditus a me quia nunc fornicatus est Ephraim contaminatus est Israhel
HOS|5|4|non dabunt cogitationes suas ut revertantur ad Dominum suum quia spiritus fornicationis in medio eorum et Dominum non cognoverunt
HOS|5|5|et respondebit arrogantia Israhel in facie eius et Israhel et Ephraim ruent in iniquitate sua ruet etiam Iudas cum eis
HOS|5|6|in gregibus suis et in armentis suis vadent ad quaerendum Dominum et non invenient ablatus est ab eis
HOS|5|7|in Domino praevaricati sunt quia filios alienos genuerunt nunc devorabit eos mensis cum partibus suis
HOS|5|8|clangite bucina in Gabaa tuba in Rama ululate in Bethaven post tergum tuum Beniamin
HOS|5|9|Ephraim in desolatione erit in die correptionis in tribubus Israhel ostendi fidem
HOS|5|10|facti sunt principes Iuda quasi adsumentes terminum super eos effundam quasi aquam iram meam
HOS|5|11|calumniam patiens Ephraim fractus iudicio quoniam coepit abire post sordem
HOS|5|12|et ego quasi tinea Ephraim et quasi putredo domui Iuda
HOS|5|13|et vidit Ephraim languorem suum et Iudas vinculum suum et abiit Ephraim ad Assur et misit ad regem ultorem et ipse non poterit sanare vos nec solvere poterit a vobis vinculum
HOS|5|14|quoniam ego quasi leaena Ephraim et quasi catulus leonis domui Iuda ego ego capiam et vadam tollam et non est qui eruat
HOS|5|15|vadens revertar ad locum meum donec deficiatis et quaeratis faciem meam
HOS|6|1|in tribulatione sua mane consurgunt ad me venite et revertamur ad Dominum
HOS|6|2|quia ipse cepit et sanabit nos percutiet et curabit nos
HOS|6|3|vivificabit nos post duos dies in die tertia suscitabit nos et vivemus in conspectu eius sciemus sequemurque ut cognoscamus Dominum quasi diluculum praeparatus est egressus eius et veniet quasi imber nobis temporaneus et serotinus terrae
HOS|6|4|quid faciam tibi Ephraim quid faciam tibi Iuda misericordia vestra quasi nubes matutina et quasi ros mane pertransiens
HOS|6|5|propter hoc dolavi in prophetis occidi eos in verbis oris mei et iudicia tua quasi lux egredientur
HOS|6|6|quia misericordiam volui et non sacrificium et scientiam Dei plus quam holocausta
HOS|6|7|ipsi autem sicut Adam transgressi sunt pactum ibi praevaricati sunt in me
HOS|6|8|Galaad civitas operantium idolum subplantata sanguine
HOS|6|9|et quasi fauces virorum latronum particeps sacerdotum in via interficientium pergentes de Sychem quia scelus operati sunt
HOS|6|10|in domo Israhel vidi horrendum ibi fornicationes Ephraim contaminatus est Israhel
HOS|6|11|sed et Iuda pone messem tibi cum convertero captivitatem populi mei
HOS|7|1|cum sanare vellem Israhel revelata est iniquitas Ephraim et malitia Samariae quia operati sunt mendacium et fur ingressus est spolians latrunculus foris
HOS|7|2|et ne forte dicant in cordibus suis omnem malitiam eorum me recordatum nunc circumdederunt eos adinventiones suae coram facie mea factae sunt
HOS|7|3|in malitia sua laetificaverunt regem et in mendaciis suis principes
HOS|7|4|omnes adulterantes quasi clibanus succensus a coquente quievit paululum civitas a commixtione fermenti donec fermentaretur totum
HOS|7|5|dies regis nostri coeperunt principes furere a vino extendit manum suam cum inlusoribus
HOS|7|6|quia adplicuerunt quasi clibanum cor suum cum insidiaretur eis tota nocte dormivit coquens eos mane ipse succensus quasi ignis flammae
HOS|7|7|omnes calefacti sunt quasi clibanus et devoraverunt iudices suos omnes reges eorum ceciderunt non est qui clamet in eis ad me
HOS|7|8|Ephraim in populis ipse commiscebatur Ephraim factus est subcinericius qui non reversatur
HOS|7|9|comederunt alieni robur eius et ipse nescivit sed et cani effusi sunt in eo et ipse ignoravit
HOS|7|10|et humiliabitur superbia Israhel in facie eius nec reversi sunt ad Dominum Deum suum et non quaesierunt eum in omnibus his
HOS|7|11|et factus est Ephraim quasi columba seducta non habens cor Aegyptum invocabant ad Assyrios abierunt
HOS|7|12|et cum profecti fuerint expandam super eos rete meum quasi volucrem caeli detraham eos caedam eos secundum auditionem coetus eorum
HOS|7|13|vae eis quoniam recesserunt a me vastabuntur quia praevaricati sunt in me et ego redemi eos et ipsi locuti sunt contra me mendacia
HOS|7|14|et non clamaverunt ad me in corde suo sed ululabant in cubilibus suis super triticum et vinum ruminabant recesserunt a me
HOS|7|15|et ego erudivi et confortavi brachia eorum et in me cogitaverunt malitiam
HOS|7|16|reversi sunt ut essent absque iugo facti sunt quasi arcus dolosus cadent in gladio principes eorum a furore linguae suae ista subsannatio eorum in terra Aegypti
HOS|8|1|in gutture tuo sit tuba quasi aquila super domum Domini pro eo quod transgressi sunt foedus meum et legem meam praevaricati sunt
HOS|8|2|me invocabunt Deus meus cognovimus te Israhel
HOS|8|3|proiecit Israhel bonum inimicus persequetur eum
HOS|8|4|ipsi regnaverunt et non ex me principes extiterunt et non cognovi argentum suum et aurum suum fecerunt sibi idola ut interirent
HOS|8|5|proiectus est vitulus tuus Samaria iratus est furor meus in eis usquequo non poterunt emundari
HOS|8|6|quia ex Israhel et ipse est artifex fecit illum et non est Deus quoniam in aranearum telas erit vitulus Samariae
HOS|8|7|quia ventum seminabunt et turbinem metent culmus stans non est in eis germen non faciet farinam quod si et fecerit alieni comedent eam
HOS|8|8|devoratus est Israhel nunc factus est in nationibus quasi vas inmundum
HOS|8|9|quia ipsi ascenderunt ad Assur onager solitarius sibi Ephraim munera dederunt amatoribus
HOS|8|10|sed et cum mercede conduxerint nationes nunc congregabo eos et quiescent paulisper ab onere regis et principum
HOS|8|11|quia multiplicavit Ephraim altaria ad peccandum factae sunt ei arae in delictum
HOS|8|12|scribam ei multiplices leges meas quae velut alienae conputatae sunt
HOS|8|13|hostias adfer adfer immolabunt carnes et comedent Dominus non suscipiet eas nunc recordabitur iniquitatis eorum et visitabit peccata eorum ipsi in Aegyptum convertentur
HOS|8|14|et oblitus est Israhel factoris sui et aedificavit delubra et Iudas multiplicavit urbes munitas et mittam ignem in civitates eius et devorabit aedes illius
HOS|9|1|noli laetari Israhel noli exultare sicut populi quia fornicatus es a Deo tuo dilexisti mercedem super omnes areas tritici
HOS|9|2|area et torcular non pascet eos et vinum mentietur eis
HOS|9|3|non habitabunt in terra Domini reversus est Ephraim Aegyptum et in Assyriis pollutum comedit
HOS|9|4|non libabunt Domino vinum et non placebunt ei sacrificia eorum quasi panis lugentium omnes qui comedunt eum contaminabuntur quia panis eorum animae ipsorum non intrabit in domum Domini
HOS|9|5|quid facietis in die sollemni in die festivitatis Domini
HOS|9|6|ecce enim profecti sunt a vastitate Aegyptus congregavit eos Memphis sepeliet eos desiderabile argenti eorum urtica hereditabit lappa in tabernaculis eorum
HOS|9|7|venerunt dies visitationis venerunt dies retributionis scitote Israhel stultum prophetam insanum virum spiritalem propter multitudinem iniquitatis tuae et multitudo amentiae
HOS|9|8|speculator Ephraim cum Deo meo propheta laqueus ruinae super omnes vias eius insania in domo Dei eius
HOS|9|9|profunde peccaverunt sicut in diebus Gabaa recordabitur iniquitatis eorum et visitabit peccata eorum
HOS|9|10|quasi uvas in deserto inveni Israhel quasi prima poma ficulneae in cacumine eius vidi patres eorum ipsi autem intraverunt ad Beelphegor et abalienati sunt in confusione et facti sunt abominabiles sicut ea quae dilexerunt
HOS|9|11|Ephraim quasi avis avolavit gloria eorum a partu et ab utero et a conceptu
HOS|9|12|quod si et enutrierint filios suos absque liberis eos faciam in hominibus sed et vae eis cum recessero ab eis
HOS|9|13|Ephraim ut vidi Tyrus erat fundata in pulchritudine et Ephraim educit ad interfectorem filios suos
HOS|9|14|da eis Domine quid dabis eis da eis vulvam sine liberis et ubera arentia
HOS|9|15|omnes nequitiae eorum in Galgal quia ibi exosos habui eos propter malitiam adinventionum eorum de domo mea eiciam eos non addam ut diligam eos omnes principes eorum recedentes
HOS|9|16|percussus est Ephraim radix eorum exsiccata est fructum nequaquam facient quod si et genuerint interficiam amantissima uteri eorum
HOS|9|17|abiciet eos Deus meus quia non audierunt eum et erunt vagi in nationibus
HOS|10|1|vitis frondosa Israhel fructus adaequatus est ei secundum multitudinem fructus sui multiplicavit altaria iuxta ubertatem terrae suae exuberavit simulacris
HOS|10|2|divisum est cor eorum nunc interibunt ipse confringet simulacra eorum depopulabitur aras eorum
HOS|10|3|quia nunc dicent non est rex nobis non enim timemus Dominum et rex quid faciet nobis
HOS|10|4|loquimini verba visionis inutilis et ferietis foedus et germinabit quasi amaritudo iudicium super sulcos agri
HOS|10|5|vaccas Bethaven coluerunt habitatores Samariae quia luxit super eum populus eius et aeditui eius super eum exultaverunt in gloria eius quia migravit ab eo
HOS|10|6|siquidem et ipse in Assur delatus est munus regi ultori confusio Ephraim capiet et confundetur Israhel in voluntate sua
HOS|10|7|transire fecit Samaria regem suum quasi spumam super faciem aquae
HOS|10|8|et disperdentur excelsa idoli peccatum Israhel lappa et tribulus ascendet super aras eorum et dicent montibus operite nos et collibus cadite super nos
HOS|10|9|ex diebus Gabaa peccavit Israhel ibi steterunt non conprehendet eos in Gabaa proelium super filios iniquitatis
HOS|10|10|iuxta desiderium meum corripiam eos congregabuntur super eos populi cum corripientur propter duas iniquitates suas
HOS|10|11|Ephraim vitula docta diligere trituram et ego transivi super pulchritudinem colli eius ascendam super Ephraim arabit Iudas confringet sibi sulcos Iacob
HOS|10|12|seminate vobis in iustitia metite in ore misericordiae innovate vobis novale tempus autem requirendi Dominum cum venerit qui docebit vos iustitiam
HOS|10|13|arastis impietatem iniquitatem messuistis comedistis frugem mendacii quia confisus es in viis tuis in multitudine fortium tuorum
HOS|10|14|consurget tumultus in populo tuo et omnes munitiones tuae vastabuntur sicut vastatus est Salman a domo eius qui iudicavit Baal in die proelii matre super filios adlisa
HOS|10|15|sic fecit vobis Bethel a facie malitiae nequitiarum vestrarum
HOS|11|1|sicuti mane transit pertransiit rex Israhel quia puer Israhel et dilexi eum et ex Aegypto vocavi filium meum
HOS|11|2|vocaverunt eos sic abierunt a facie eorum Baalim immolabant et simulacris sacrificabant
HOS|11|3|et ego quasi nutricius Ephraim portabam eos in brachiis meis et nescierunt quod curarem eos
HOS|11|4|in funiculis Adam traham eos in vinculis caritatis et ero eis quasi exaltans iugum super maxillas eorum et declinavi ad eum ut vesceretur
HOS|11|5|non revertetur in terram Aegypti et Assur ipse rex eius quoniam noluerunt converti
HOS|11|6|coepit gladius in civitatibus eius et consumet electos eius et comedet capita eorum
HOS|11|7|et populus meus pendebit ad reditum meum iugum autem inponetur ei simul quod non auferetur
HOS|11|8|quomodo dabo te Ephraim protegam te Israhel quomodo dabo te sicut Adama ponam te ut Seboim conversum est in me cor meum pariter conturbata est paenitudo mea
HOS|11|9|non faciam furorem irae meae non convertar ut disperdam Ephraim quoniam Deus ego et non homo in medio tui Sanctus et non ingrediar civitatem
HOS|11|10|post Dominum ambulabunt quasi leo rugiet quia ipse rugiet et formidabunt filii maris
HOS|11|11|et avolabunt quasi avis ex Aegypto et quasi columba de terra Assyriorum et conlocabo eos in domibus suis dicit Dominus
HOS|11|12|circumdedit me in negatione Ephraim et in dolo domus Israhel Iudas autem testis descendit cum Deo et cum sanctis fidelis
HOS|12|1|Ephraim pascit ventum et sequitur aestum tota die mendacium et vastitatem multiplicat et foedus cum Assyriis iniit et oleum in Aegyptum ferebat
HOS|12|2|iudicium ergo Domini cum Iuda et visitatio super Iacob iuxta vias eius et iuxta adinventiones eius reddet ei
HOS|12|3|in utero subplantavit fratrem suum et in fortitudine sua directus est cum angelo
HOS|12|4|et invaluit ad angelum et confortatus est flevit et rogavit eum in Bethel invenit eum et ibi locutus est nobiscum
HOS|12|5|et Dominus Deus exercituum Dominus memoriale eius
HOS|12|6|et tu ad Deum tuum converteris misericordiam et iudicium custodi et spera in Deo tuo semper
HOS|12|7|Chanaan in manu eius statera dolosa calumniam dilexit
HOS|12|8|et dixit Ephraim verumtamen dives effectus sum inveni idolum mihi omnes labores mei non invenient mihi iniquitatem quam peccavi
HOS|12|9|et ego Dominus Deus tuus ex terra Aegypti adhuc sedere te faciam in tabernaculis sicut in diebus festivitatis
HOS|12|10|et locutus sum super prophetas et ego visionem multiplicavi et in manu prophetarum adsimilatus sum
HOS|12|11|si Galaad idolum tamen frustra erant in Galgal bubus immolantes nam et altaria eorum quasi acervi super sulcos agri
HOS|12|12|fugit Iacob in regionem Syriae et servivit Israhel in uxore et in uxore servavit
HOS|12|13|in propheta autem eduxit Dominus Israhel de Aegypto et in propheta servatus est
HOS|12|14|ad iracundiam me provocavit Ephraim in amaritudinibus suis et sanguis eius super eum veniet et obprobrium eius restituet ei Dominus suus
HOS|13|1|loquente Ephraim horror invasit Israhel et deliquit in Baal et mortuus est
HOS|13|2|et nunc addiderunt ad peccandum feceruntque sibi conflatile de argento suo quasi similitudinem idolorum factura artificum totum est his ipsi dicunt immolate homines vitulos adorantes
HOS|13|3|idcirco erunt quasi nubes matutina et sicut ros matutinus praeteriens sicut pulvis turbine raptus ex area et sicut fumus de fumario
HOS|13|4|ego autem Dominus Deus tuus ex terra Aegypti et Deum absque me nescies et salvator non est praeter me
HOS|13|5|ego cognovi te in deserto in terra solitudinis
HOS|13|6|iuxta pascua sua et adimpleti sunt et saturati elevaverunt cor suum et obliti sunt mei
HOS|13|7|et ero eis quasi leaena sicut pardus in via Assyriorum
HOS|13|8|occurram eis quasi ursa raptis catulis et disrumpam interiora iecoris eorum et consumam eos ibi quasi leo bestia agri scindet eos
HOS|13|9|perditio tua Israhel tantummodo in me auxilium tuum
HOS|13|10|ubi est rex tuus maxime nunc salvet te in omnibus urbibus tuis et iudices tui de quibus dixisti da mihi regem et principes
HOS|13|11|dabo tibi regem in furore meo et auferam in indignatione mea
HOS|13|12|conligata est iniquitas Ephraim absconditum peccatum eius
HOS|13|13|dolores parturientis venient ei ipse filius non sapiens nunc enim non stabit in contritione filiorum
HOS|13|14|de manu mortis liberabo eos de morte redimam eos ero mors tua o mors ero morsus tuus inferne consolatio abscondita est ab oculis meis
HOS|13|15|quia ipse inter fratres dividet adducet urentem ventum Dominus de deserto ascendentem et siccabit venas eius et desolabit fontem eius et ipse diripiet thesaurum omnis vasis desiderabilis
HOS|14|1|pereat Samaria quoniam ad amaritudinem concitavit Dominum suum in gladio pereat parvuli eorum elidantur et fetae eius discindantur
HOS|14|2|convertere Israhel ad Dominum Deum tuum quoniam corruisti in iniquitate tua
HOS|14|3|tollite vobiscum verba et convertimini ad Dominum dicite ei omnem aufer iniquitatem et accipe bonum et reddemus vitulos labiorum nostrorum
HOS|14|4|Assur non salvabit nos super equum non ascendemus nec dicemus ultra dii nostri opera manuum nostrarum quia eius qui in te est misereberis pupilli
HOS|14|5|sanabo contritiones eorum diligam eos spontanee quia aversus est furor meus ab eo
HOS|14|6|ero quasi ros Israhel germinabit quasi lilium et erumpet radix eius ut Libani
HOS|14|7|ibunt rami eius et erit quasi oliva gloria eius et odor eius ut Libani
HOS|14|8|convertentur sedentes in umbra eius vivent tritico et germinabunt quasi vinea memoriale eius sicut vinum Libani
HOS|14|9|Ephraim quid mihi ultra idola ego exaudiam et dirigam eum ego ut abietem virentem ex me fructus tuus inventus est
HOS|14|10|quis sapiens et intelleget ista intellegens et sciet haec quia rectae viae Domini et iusti ambulabunt in eis praevaricatores vero corruent in eis
