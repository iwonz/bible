HOS|1|1|Слово Господнє, що було до Осії, Беерового сина, за днів Уззійї, Йотама, Ахаза, Єзекії, Юдиних царів, та за днів Єровоама, Йоашового сина, Ізраїлевого царя.
HOS|1|2|Початок того, що Господь говорив через Осію. І сказав Господь до Осії: Іди, візьми собі жінку блудливу, і вона породить дітей блуду, бо сильно блудодіє цей Край, відступивши від Господа.
HOS|1|3|І він пішов, і взяв Ґомер, дочку Дівлаїма, і вона зачала, і породила йому сина.
HOS|1|4|І сказав Господь до нього: Назви ім'я йому Їзреел, бо ще трохи, і покараю кров Їзреелу на домі Єгу, і вчиню кінець царству Ізраїлевого дому.
HOS|1|5|І станеться того дня, і Я зламаю Ізраїлевого лука в долині Їзреел.
HOS|1|6|І зачала вона ще, і породила дочку. І сказав Він йому: Назви ім'я їй Ло-Рухама, бо більше Я вже не змилуюся над Ізраїлевим домом, бо вже більше не прощу Я їм.
HOS|1|7|А над Юдиним домом Я змилуюся, і допоможу їм через Господа, їхнього Бога, але не допоможу їм ані луком, ані мечем, ані війною, кіньми чи верхівцями.
HOS|1|8|І відлучила вона Ло-Рухаму, і зачала знову, і породила сина.
HOS|1|9|А Він сказав: Назви ім'я йому Ло-Аммі, бо ви не народ Мій, і Я не буду ваш!
HOS|1|10|(2-1) І буде число Ізраїлевих синів, як морський пісок, що його не можна ані зміряти, ані злічити. І станеться, замість того, що говориться їм: Ви не народ Мій, буде їм сказано: Ви сини Бога Живого.
HOS|1|11|(2-2) І будуть зібрані разом сини Юдині та сини Ізраїлеві, і настановлять собі одного голову, і повиходять з землі, бо великий день Їзреелу.
HOS|2|1|(2-3) Скажіть своїм братам: Народ Мій, а своїм сестрам: Помилувана.
HOS|2|2|(2-4) Судіться з вашою матір'ю, судіться, бо вона не жінка Моя, а Я не її чоловік, і нехай вона відкине від себе свій блуд, і з-поміж своїх перс свій перелюб,
HOS|2|3|(2-5) щоб Я не роздягнув її до нага, і не поставив її такою, як у день її народження, і щоб не зробив Я її пустинею, і не обернув її на суху землю, і не забив її спрагою.
HOS|2|4|(2-6) Над синами ж її Я не змилуюся, бо вони сини блуду,
HOS|2|5|(2-7) бо їхня мати блудлива була, та, що ними була вагітна, сором чинила, бо казала вона: Я піду за своїми полюбовниками, що дають мені хліб мій та воду мою, мою вовну та льон мій, оливу мою та напої мої.
HOS|2|6|(2-8) Тому то ось Я вкрию твою дорогу тернями, і обгороджу її огорожею, і стежок своїх не знайде вона.
HOS|2|7|(2-9) І буде вона гнатися за своїми полюбовниками, але не дожене їх, і буде шукати їх, та не знайде. І скаже вона: Піду я, і вернуся до мого першого чоловіка, бо краще було мені тоді, як тепер.
HOS|2|8|(2-10) А вона не знає, що то Я давав їй збіжжя, і виноградний сік, і свіжу оливу, і примножив їй срібло та золото, яке вони звернули на Ваала.
HOS|2|9|(2-11) Тому то заберу назад Своє збіжжя в його часі, а Мій сік виноградний в його умовленому часі, і заберу Свою вовну та Свій льон, що був на покриття її наготи.
HOS|2|10|(2-12) А тепер відкрию її наготу на очах її коханців, і ніхто не врятує її від Моєї руки.
HOS|2|11|(2-13) І зроблю кінець усякій радості її, святу її, новомісяччю її, і суботі її, та всякому святковому часові.
HOS|2|12|(2-14) І спустошу її виноградника та її фіґове дерево, про які вона говорила: Це мені дар за блудодійство, що дали мені мої полюбовники. А Я оберну їх на ліс, і їх пожере польова звірина!
HOS|2|13|(2-15) І навіщу її за дні Ваалів, коли вона кадила. І приоздоблювалася ти своєю носовою сережкою та своїм нашийником, і ходила за своїми полюбовниками, а Мене забувала, говорить Господь.
HOS|2|14|(2-16) Тому то ось Я намовлю її, і попроваджу її до пустині, і буду говорити до серця її.
HOS|2|15|(2-17) І дам їй виноградники звідти та долину Ахор за двері надії, і вона буде там співати, як за днів своєї молодости, як за дня виходу її з єгипетського краю.
HOS|2|16|(2-18) І станеться, того дня говорить Господь ти кликатимеш: Чоловіче мій, і не будеш більше кликати Мене: Мій ваале.
HOS|2|17|(2-19) І усуну імена Ваалів з її уст, і вони не будуть більше згадувані своїм іменем.
HOS|2|18|(2-20) І складу їм заповіта того дня з польовою звіриною, і з птаством небесним, та з плазуючим по землі, і лука й меча та війну знищу з землі, і покладу їх безпечно.
HOS|2|19|(2-21) І заручуся з тобою навіки, і заручуся з тобою справедливістю, і правосуддям, і милістю та любов'ю.
HOS|2|20|(2-22) І заручуся з тобою вірністю, і ти пізнаєш Господа.
HOS|2|21|(2-23) І станеться того дня, Я почую, говорить Господь, почую небо, а воно почує землю,
HOS|2|22|(2-24) а земля задоволить збіжжя, і виноградний сік, і оливу, а вони задовольнять Їзреела.
HOS|2|23|(2-25) І обсію її Собі на землі, і змилуюся над Ло-Рухамою, і скажу до Ло-Амі: Ти народ Мій, а він скаже: Мій Боже!
HOS|3|1|І сказав Господь мені ще: Іди, покохай жінку, кохану приятелем, але перелюбну, подібно, як любить Господь Ізраїлевих синів, а вони звертаються до інших богів, і кохаються у виноградних коржиках.
HOS|3|2|І я купив її собі за п'ятнадцять шеклів срібла й хомер ячменю та летех ячменю.
HOS|3|3|І сказав я до неї: Сиди довгі дні в мене, не будь блудлива, і не будь нічия, також і я буду такий до тебе.
HOS|3|4|Бо Ізраїлеві сини будуть сидіти довгі дні без царя та без князя, і без жертви та без камінного стовпа, і без ефода та без домашніх божків.
HOS|3|5|Потому Ізраїлеві сини навернуться, і будуть шукати Господа, Бога свого, та царя свого Давида, і за останніх днів з тремтінням обернуться до Господа та до Його добра.
HOS|4|1|Послухайте слова Господнього, Ізраїлеві сини, бо Господь має прю із мешканцями земними, бо нема на землі ані правди, ні милости, ані богопізнання.
HOS|4|2|Клянуть та неправду говорять, і вбивають та крадуть, і чинять перелюб, поставали насильниками, а кров доторкається крови.
HOS|4|3|Тому то в жалобу земля упаде, і стане нещасним усякий мешканець на ній з польовою звіриною й з птаством небесним, і також морські риби погинуть.
HOS|4|4|Та тільки ніхто хай не свариться, і хай не плямує ніхто! А народ Мій як суперечник з священиком.
HOS|4|5|І спіткнешся ти вдень, і спіткнеться з тобою й пророк уночі, і знищу Я матір твою!
HOS|4|6|Погине народ Мій за те, що не має знання: тому, що знання ти відкинув, відкину й тебе, щоб не був ти для Мене священиком. А тому, що забув ти Закон свого Бога, забуду синів твоїх й Я!
HOS|4|7|Що більше розмножуються, то більше грішать проти Мене. Їхню славу зміню Я на ганьбу!
HOS|4|8|Вони жертву за прогріх народу Мого їдять, і до провини його свою душу схиляють.
HOS|4|9|І буде священикові, як і народові, і дороги його навіщу Я на нім, і йому відплачу згідно вчинків його.
HOS|4|10|І вони будуть їсти, але не наситяться, чинитимуть блуд, та не розмножаться, бо покинули дбати про Господа.
HOS|4|11|Блуд і вино та сік виноградний володіють їхнім серцем.
HOS|4|12|Народ Мій допитується в свого дерева, і об'являє йому його палиця, бо дух блудодійства заводить до блуду, і вони заблудили від Бога свого.
HOS|4|13|На верховинах гірських вони жертви приносять, і кадять на взгір'ях під дубом, і тополею та теребінтом, бо хороша їхня тінь, тому ваші дочки блудливими стали, а ваші невістки вчиняють перелюб.
HOS|4|14|Та не покараю ще ваших дочок, що вони блудодіють, та ваших невісток, що чинять перелюб, як відходять вони з блудодійками і жертви приносять з розпусницями. А народ без знання загибає!
HOS|4|15|Якщо ти блудливий, Ізраїлю, нехай Юда не буде провинний! І не ходіть до Ґілґалу, і не приходьте до Бет-Авену, і не присягайте: Як живий Господь!
HOS|4|16|Бо Ізраїль зробився упертий, немов та уперта корова. Та тепер Господь пастиме їх, як вівцю на привіллі!
HOS|4|17|Прилучивсь до бовванів Єфрем, покинь ти його!
HOS|4|18|Збір п'яниць звироднілих учинився розпусним, їхні провідники покохали нечистість.
HOS|4|19|Вітер їх похапає на крила свої, і вони посоромляться жертов своїх.
HOS|5|1|Послухайте цього, священики, і почуйте, Ізраїлів доме, а ви, царський доме, візьміть до вух, бо вам буде суд, бо ви для Міцпи були пасткою й сіткою, розтягненою на Фавор.
HOS|5|2|І глибоко вгрузли в розпусті вони, та Я поплямую всіх їх.
HOS|5|3|Я знаю Єфрема, а Ізраїль не схований передо Мною, бо тепер блудодійним, Єфреме, ти став, занечистивсь Ізраїль.
HOS|5|4|Не дають їхні вчинки вернутись до Бога, бо дух блудодійства в середині їхній, і не відають Господа.
HOS|5|5|І гордість Ізраїлева засвідчиться перед обличчям його. А Ізраїль й Єфрем упадуть за провину свою, також Юда із ними впаде.
HOS|5|6|З своєю отарою та з своєю худобою вони Господа підуть шукати, але не знайдуть, Він від них віддалився.
HOS|5|7|Вони зрадили Господа, бо породили сторонніх дітей, тепер їх пожере молодик разом із частками їхнього поля.
HOS|5|8|Засурміте у рога в Ґів'ї, сурмою в Рамі, закричіть у Бет-Авені за тобою, Веніямине!
HOS|5|9|В день картання Єфрем за спустошення стане; поміж племенами Ізраїля Я завідомив про певне.
HOS|5|10|Стали зверхники Юди, мов ті, що межу переносять, на них виллю, як воду, Свій гнів!
HOS|5|11|Єфрем став пригноблений, судом розбитий, бо він намагався ходити за марнотою.
HOS|5|12|І Я буду, як міль, для Єфрема, і мов та гнилизна для дому Юди.
HOS|5|13|І побачив Єфрем свою хворість, а Юда свого чиряка, і Єфрем відійшов до Ашшура і послав до царя до великого. Та він вилікувати вас не зможе, і не вигоїть вам чиряка!
HOS|5|14|Бо Я немов лев для Єфрема, і немов той левчук дому Юди. Я, Я розшматую й піду, і ніхто не врятує!
HOS|5|15|Піду, повернуся до місця Свого, аж поки провини своєї вони не признають, і не стануть шукати Мого лиця. Та в утиску будуть шукати Мене!
HOS|6|1|Ходіть, і вернімось до Господа, бо Він пошматував і нас вилікує, ударив і нас перев'яже!
HOS|6|2|Оживить він нас до двох день, а третього дня нас поставить, і будемо жити ми перед обличчям Його.
HOS|6|3|І пізнаймо, намагаймось пізнати ми Господа! Міцно поставлений прихід Його, мов зірниці, і Він прийде до нас, немов дощ, немов дощ весняний, що напоює землю.
HOS|6|4|Що, Єфреме, зроблю Я тобі, що зроблю тобі, Юдо? Бо ваша любов, немов хмара поранку, і мов та роса, що зникає уранці,
HOS|6|5|тому Я тесав їх пророками, позабивав їх прореченням уст Своїх, і суд Мій, як світло те, вийде.
HOS|6|6|Бо Я милости хочу, а не жертви, і Богопізнання більше від цілопалень.
HOS|6|7|Вони заповіта Мого порушили, мов той Адам, вони там Мене зрадили.
HOS|6|8|Ґілеад, місто злочинців, повне кривавих слідів.
HOS|6|9|І як той розбишака чигає, так ватага священиків на дорозі в Сихем учиняють розбій, бо злочин учиняють вони.
HOS|6|10|У домі Ізраїля бачу жахливе, там блуд у Єфрема, занечистивсь Ізраїль.
HOS|6|11|Також, Юдо, для тебе жнива приготовлені, як Я долю народу Свого поверну!
HOS|7|1|Коли Я лікую Ізраїля, то виявляю гріх Єфремів та зло Самарії, бо роблять вони неправдиве, і злодій приходить, грабує на вулиці банда.
HOS|7|2|І не думають в серці своєму, що Я пам'ятаю про все їхнє зло. Тепер їхні вчинки ось їх оточили і перед обличчям Моїм поставали.
HOS|7|3|Вони злістю своєю втішають царя, а своїми обманами зверхників.
HOS|7|4|Усі вони чинять перелюб, мов піч, яку пекар розпалює, що напалювати перестає, як тісто замісить та вкисне воно.
HOS|7|5|У святковий день нашого царя похворіли князі від жару вина, і він простяг до насмішників руку свою.
HOS|7|6|Бо їхнє нутро, як піч, у них палає їхнє серце: всю ніч спить їхній гнів, а на ранок горить, як палючий огонь.
HOS|7|7|Вони всі гарячі, як піч, і суддів своїх пожирають. Усі царі їхні попадали, між ними нікого нема, хто б кликав до Мене.
HOS|7|8|Змішався Єфрем із народами, Єфрем став млинцем, що печеться неперевернений.
HOS|7|9|Його силу чужі пожирають, та про те він не знає, вже й волосся посивіло в нього, а того він не знає.
HOS|7|10|І гордість Ізраїля свідчить на нього, і до Господа, Бога свого вони не вертаються, і не шукають Його у всім цім.
HOS|7|11|А Єфрем став, як голуб, нерозумний, немудрий: закликають в Єгипет, а йдуть в Асирію.
HOS|7|12|Як підуть вони, розтягну Свою сітку над ними, стягну їх додолу, мов птаство небесне, за злобою їхньою Я їх караю.
HOS|7|13|Горе їм, бо від Мене вони відійшли, погуба на них, бо повстали вони проти Мене! Хоч Я викупив їх, та вони проти Мене говорять неправду.
HOS|7|14|І вони в своїм серці не кличуть до Мене, як виють на ложах своїх, точать сварку за хліб та вино, і відступають від Мене.
HOS|7|15|А Я їх картав, їхні рамена зміцняв, а вони зло на Мене задумують...
HOS|7|16|Вони навертаються, та не до Всевишнього, стали, немов той обманливий лук... Упадуть від меча їхні князі за гордість свого язика, це їхня наруга в єгипетськім краї!
HOS|8|1|Рога до уст своїх, та й засурми: на дім Божий спадає неначе орел, бо переступили вони заповіта Мого, і на Закона Мого повстали.
HOS|8|2|До Мене взивають вони: Мій Боже, познали Тебе ми, Ізраїлю!
HOS|8|3|Покинув Ізраїль добро, ворог його пожене!
HOS|8|4|Вони ставлять царя, але не від Мене, вони князя ставлять, але Я не знаю! Вони з срібла свого та із золота свого божків наробили собі, щоб загинути,
HOS|8|5|відкинув теля твоє Я, Самаріє! Мій гнів запалився на них, аж доки не можуть вони від провини очиститись?
HOS|8|6|Бо й воно від Ізраїля. Зробив його майстер, і воно то не Бог, бо теля самарійське на кавалки обернеться.
HOS|8|7|А що вітер вони засівають, то бурю пожнуть, в них не буде й колосся, а зерно не видасть муки, коли ж видасть, чужі поковтають її.
HOS|8|8|Ізраїль проковтнений, став між народами він як та річ, що до неї немає замилування.
HOS|8|9|Бо вони відійшли до Ашшуру, як дикий осел, що самітний собі, а Єфрем за любов дає дари любовні.
HOS|8|10|І хоч вони здобувають прихильників серед поганів, Я їх позбираю тепер, і незабаром вони перестануть помазувати царя, і князів.
HOS|8|11|Бо жертівників був намножив Єфрем, щоб грішити, на провину йому стали ці жертівники!
HOS|8|12|Я можу йому написати Закон Свій хоч тисячу разів, як чуже пораховане буде!
HOS|8|13|Вони ж жертви кохають, ріжуть м'ясо й їдять, та Господь не вподобує їх. Тепер Він згадає про їхню провину та їхні гріхи покарає, вони до Єгипту повернуться!
HOS|8|14|Ізраїль забув про свого Творця та й будує палати, а Юда намножив твердинні міста, та пошлю Я огонь на його ці міста, і пожере він палати його!
HOS|9|1|Не тішся, Ізраїлю, радістю, як ті народи, бо ти чиниш блуд, відступаючи від свого Бога, дар блудодійний кохаєш на всіх токах збіжжевих.
HOS|9|2|Годувати не буде їх тік та чавило, а сік виноградний зведе їх.
HOS|9|3|Не будуть сидіти в Господньому Краї вони, і Єфрем до Єгипту повернеться, і вони будуть їсти нечисте в Асирії.
HOS|9|4|Господеві вина вони лити не будуть, і жертви не будуть приємні Йому; це буде для них, немов хліб похоронний, усі, що будуть його споживати, занечистяться, бо їхній хліб для насичення їх, не для дому Господнього.
HOS|9|5|Що зробите ви на день урочистий та на день свята Господнього?
HOS|9|6|Бо йдуть ось вони до Асирії, їх збирає Єгипет, Мемфіс їх ховає, коштовність їхнього срібла посяде кропива, будяччя по їхніх наметах.
HOS|9|7|Прийшли дні навіщення, прийшли дні заплати, Ізраїль пізнає оце: Нерозумний пророк цей, шалений муж духа, за численність провин твоїх і велике зненавидження!
HOS|9|8|Єфрем сторож із Богом моїм, пророк пастка птахолова на всіх дорогах його, ненависть у домі Бога його.
HOS|9|9|Глибоко зіпсулись вони, як за днів тих Ґів'ї, Він згадає за їхні провини, Він їхні гріхи покарає!
HOS|9|10|Немов виноград на пустині, знайшов Я Ізраїля, як фіґу поранню на фіґовім дереві, Я бачив був ваших батьків на початку його, та вони до Баал-Пеору прийшли, і себе присвятили для Бошета, і стали гидотою, як полюблене ними.
HOS|9|11|Єфремова слава, як птах, відлетить: не буде народження, ані зачаття, ані вагітности.
HOS|9|12|Бо якщо вони викохають свої діти, то їх повбиваю, так що не буде людини, бо горе їм, як відступлю Я від них.
HOS|9|13|Єфрем, як Я бачу, для вловів йому подали його власних дітей, і Єфрем поведе своїх власних дітей на заріз...
HOS|9|14|Дай їм, Господи, що ж Ти даси? дай їм утробу неплідну та висохлі груди!
HOS|9|15|Усе їхнє зло у Ґілґалі, бо там Я зненавидів їх; за зло їхніх учинків Я вижену їх з Свого дому. Не буду їх більше любити, всі їхні князі ворохобники!
HOS|9|16|Побитий Єфрем, їхній корень посох, він плоду не зродить. А коли вони зродять, то Я повбиваю улюблених їхнього лона.
HOS|9|17|Відкине їх Бог мій, бо вони неслухняні для Нього були, і будуть вони мандрувати між народами.
HOS|10|1|Ізраїль буйний виноград, що родить подібне собі. Та за многістю плоду свого він намножує жертівники, за добрістю Краю свого бовванські стовпи прикрашає.
HOS|10|2|Облудне їхнє серце, тому винні тепер вони будуть, Він їхні жертівники понищить поруйнує стовпи їхні.
HOS|10|3|Бо тепер вони кажуть: Нема в нас царя, бо ми не боялися Господа, а цар що нам зробить?
HOS|10|4|Говорять порожні слова, клянуться фальшиво, коли заповіта складають, і на грядках польових цвіте їхнє правосуддя, немов той полин.
HOS|10|5|За телят Бет-Авену бояться мешканці Самарії, бо в жалобі опинився через нього народ його, а жерці будуть плакати над ним, за славу його, що пішла на вигнання від нього.
HOS|10|6|Запроваджений буде і він в Асирію цареві великому в дар. Прийме сором Єфрем, і посоромлений буде Ізраїль за раду свою.
HOS|10|7|Самарія загине; її цар немов тріска ота на поверхні води!
HOS|10|8|І поруйновані будуть висоти Авена, Ізраїлів гріх, тернина й будяччя зросте на їхніх жертівниках, і до гір вони скажуть: Накрийте ви нас! а до взгір'їв: На нас упадіть!
HOS|10|9|Від днів Ґів'ї грішив ти, Ізраїлю! Там вони полишились були, чи ж їх не досягне в Ґів'ї війна проти синів беззаконних?
HOS|10|10|За жаданням Своїм покараю Я їх, і зберуться народи на них, і покарані будуть вони за подвійні провини свої.
HOS|10|11|А Єфрем це привчена телиця, що звикла вона молотити, Сам ярмо накладу на її товсту шию, запряжу Я Єфрема, Юда буде орати, Яків буде собі скородити.
HOS|10|12|Сійте собі на справедливість, за милістю жніть, оріте собі переліг, бо час навернутись до Господа, ще поки Він прийде і правду лине вам дощем.
HOS|10|13|Ви беззаконня орали, пожали ви кривду, плід брехні споживали, бо надіявся ти на дорогу свою, на многість лицарства свого.
HOS|10|14|І станеться шум по народах твоїх, і всі твердині твої поруйновані будуть, як Шалман зруйнував Бет-Арбел в час війни, була мати з синами убита.
HOS|10|15|Отак вам учинить Бет-Ел за зло вашого зла, конче згине Ізраїлів цар на світанку!
HOS|11|1|Як Ізраїль був хлопцем, Я його покохав, і з Єгипту покликав Я сина Свого.
HOS|11|2|Як часто їх кликав, так вони йшли від Мене, приносили жертви Ваалам, і кадили бовванам.
HOS|11|3|Я ж Єфрема ходити навчав, Я їх брав на рамена Свої, та не знали вони, що Я їх лікував.
HOS|11|4|Я тягнув їх шнурками, що людям лицюють, шнурками любови, і був Я для них немов ті, що здіймають ярмо з-над їхньої шиї, і Я їх годував.
HOS|11|5|До краю єгипетського він не вернеться, та Ашшур він буде для нього царем, бо вони не хотіли вернутись до Мене.
HOS|11|6|А містами його ґрасуватиме меч, і засуви його повиламлює він та й пожере їх за задуми їхні.
HOS|11|7|А народ Мій схильний відпадати від Мене, і хоч кличуть його догори, він не підіймається разом.
HOS|11|8|Як тебе Я, Єфреме, віддам, як видам тебе, о Ізраїлю? Як тебе Я віддам, як Адму, учиню тебе, мов Цевоїм? У Мені перевернулося серце Моє, розпалилася разом і жалість Моя!
HOS|11|9|Не вчиню жару гніву Свого, більше нищити Єфрема не буду, бо Бог Я, а не людина, серед тебе Святий, і не прийду в люті гніву.
HOS|11|10|За Господом підуть вони, а Він заричить, немов лев, і Він заричить, і від заходу прийдуть в тремтінні сини.
HOS|11|11|Вони прийдуть в тремтінні, як птах із Єгипту, і як голуб із краю Ашшура, і Я посаджу їх по їхніх домах, говорить Господь.
HOS|11|12|(12-1) Єфрем оточив Мене лжею, лукавством Ізраїлів дім, а Юда держався ще з Богом і з святими був вірний.
HOS|12|1|(12-2) Єфрем пасе вітра й женеться за вітром із сходу. Неправду й руїну розмножує він кожного дня, умову складають з Ашшуром, олива ж несеться в Єгипет.
HOS|12|2|(12-3) Та в Господа з Юдою пря, і Якова Він навістить за путями його, за ділами його йому зверне.
HOS|12|3|(12-4) Він в утробі тримав за п'яту свого брата, а в силі своїй він боровся із Богом,
HOS|12|4|(12-5) і боровся він з Анголом, та й переміг. Плакав він, і благав він Його, у Бет-Елі знайшов Він його, і там з нами говорить.
HOS|12|5|(12-6) А Господь Бог Саваот, Його Ймення Господь.
HOS|12|6|(12-7) А ти через Бога свого навернешся, стережи милість та суд, і завжди надійся на Бога свого!
HOS|12|7|(12-8) Немов Ханаан, у нього в руці неправдива вага, любить він кривду чинити.
HOS|12|8|(12-9) І каже Єфрем: Справді я збагатився, знайшов я маєток собі! У всіх моїх чинах не знайдуть провини мені, що гріхом би була.
HOS|12|9|(12-10) А Я Господь, Бог твій від краю єгипетського, ще в наметах тебе посаджу, немов за днів свята.
HOS|12|10|(12-11) І Я говорив до пророків, і видіння розмножив, і через пророків Я притчі казав.
HOS|12|11|(12-12) Хіба беззаконня лишив Ґілеад, і марнотою стались лиш там? У Ґілґалі приносили в жертву волів, а їхні жертівники мов ті купи каміння на борознах пільних.
HOS|12|12|(12-13) І втік Яків на поле Арама, а Ізраїль за жінку робив, і за жінку отару стеріг.
HOS|12|13|(12-14) І через пророка Господь із Єгипту Ізраїля вивів, і пророком стережений був він.
HOS|12|14|(12-15) Єфрем Господа гірко розгнівав, і тому його вчинки криваві Він лишить на ньому, і поверне йому його сором.
HOS|13|1|Як Єфрем говорив, то тремтіли, він піднесений був ув Ізраїлі, та через Ваала згрішив і помер.
HOS|13|2|А тепер іще більше грішать, бо зробили собі вони відлива з срібла свого, божків за своєю подобою; робота майстрів усе те, розмовляють із ними вони; ті люди, що жертву приносять, цілують телят.
HOS|13|3|Тому вони стануть, як хмара поранку, і мов та роса, що зникає вранці, немов та полова, що з току виноситься бурею, і наче із комина дим.
HOS|13|4|А Я Господь, Бог твій від краю єгипетського, і Бога, крім Мене, не будеш ти знати, і крім Мене немає Спасителя.
HOS|13|5|Я тебе на пустині пізнав, у пересохлому краї.
HOS|13|6|Мали добрі пасовиська й ситі були, наситилися і загордилось їхнє серце, тому то забули про Мене вони!
HOS|13|7|І став Я для них, немов лев, на дорозі чигаю, немов та пантера.
HOS|13|8|Нападу Я на них, немов та ведмедиця, що дітей загубила, і те розірву, у що серце їхнє замкнене, і їх, як левчук, пожеру там, шматуватиме їх польова звірина.
HOS|13|9|Погубив ти себе, о Ізраїлю, бо ти був проти Мене, спасіння свого.
HOS|13|10|Де цар твій тоді? Нехай він поможе тобі по містах твоїх усіх! А де судді твої, що про них ти сказав: Дай нам царя та князів?
HOS|13|11|Я тобі дав царя в Своїм гніві, і забрав у Своїй ревності.
HOS|13|12|Провина Єфремова зв'язана, схований прогріх його.
HOS|13|13|Болі, немов породіллі, надійдуть на нього. Не мудрий він син, бо інакше не був би так довго у матернім нутрі.
HOS|13|14|З рук шеолу Я викуплю їх, від смерти їх вибавлю. Де, смерте, жало твоє? Де, шеоле, твоя перемога? Жаль сховається перед очима Моїми!
HOS|13|15|Хоч він дає плід між братами, але прийде вітер зо сходу, вітер Господній, що зійде з пустині, і всохне його джерело, і пересохне криничка його, понищить він скарб всіх коштовних речей!
HOS|13|16|(14-1) Завинить Самарія, бо стала уперта до Бога свого, поляжуть вони від меча! Порозбивані будуть їхні діти, вагітні їхні розпороті будуть!
HOS|14|1|(14-2) Вернися, Ізраїлю, до Господа, Бога свого, бо спіткнувся ти через провину свою!
HOS|14|2|(14-3) Візьміть із собою слова, та й зверніться до Господа, до Нього промовте: Прости нам усяку провину, та добре прийми, і ми принесемо у жертву плода своїх уст!
HOS|14|3|(14-4) Ашшур не спасе нас, не будемо їздити ми на коні, і не скажемо вже чинові рук наших: боже наш, бо тільки Тобою помилуваний сирота.
HOS|14|4|(14-5) Ворохобність їхню вилікую, добровільно любитиму їх, бо Мій гнів відвернувся від нього.
HOS|14|5|(14-6) Я буду Ізраїлеві, як роса, розцвіте він, неначе лілея, і пустить коріння своє, мов Ліван.
HOS|14|6|(14-7) Розійдуться його пагінці, і буде його пишнота, мов оливне те дерево, а пахощ його мов Ліван.
HOS|14|7|(14-8) Навернуться ті, що сиділи під тінню його, збіжжя оживлять вони й зацвітуть, немов той виноград, будуть згадки про нього, немов про ліванське вино.
HOS|14|8|(14-9) Єфрем, що йому до бовванів іще? Я вислухав вже та побачив його, Я для нього немов кипарис той зелений: з Мене знайдений буде твій плід.
HOS|14|9|(14-10) Хто мудрий, то це зрозуміє, розумний і пізнає, бо прості Господні дороги, і праведні ходять по них, а грішні спіткнуться на них!
