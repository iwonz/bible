1JOHN|1|1|That which was from the beginning, which we have heard, which we have seen with our eyes, which we have looked at and our hands have touched--this we proclaim concerning the Word of life.
1JOHN|1|2|The life appeared; we have seen it and testify to it, and we proclaim to you the eternal life, which was with the Father and has appeared to us.
1JOHN|1|3|We proclaim to you what we have seen and heard, so that you also may have fellowship with us. And our fellowship is with the Father and with his Son, Jesus Christ.
1JOHN|1|4|We write this to make our joy complete.
1JOHN|1|5|This is the message we have heard from him and declare to you: God is light; in him there is no darkness at all.
1JOHN|1|6|If we claim to have fellowship with him yet walk in the darkness, we lie and do not live by the truth.
1JOHN|1|7|But if we walk in the light, as he is in the light, we have fellowship with one another, and the blood of Jesus, his Son, purifies us from all sin.
1JOHN|1|8|If we claim to be without sin, we deceive ourselves and the truth is not in us.
1JOHN|1|9|If we confess our sins, he is faithful and just and will forgive us our sins and purify us from all unrighteousness.
1JOHN|1|10|If we claim we have not sinned, we make him out to be a liar and his word has no place in our lives.
1JOHN|2|1|My dear children, I write this to you so that you will not sin. But if anybody does sin, we have one who speaks to the Father in our defense--Jesus Christ, the Righteous One.
1JOHN|2|2|He is the atoning sacrifice for our sins, and not only for ours but also for the sins of the whole world.
1JOHN|2|3|We know that we have come to know him if we obey his commands.
1JOHN|2|4|The man who says, "I know him," but does not do what he commands is a liar, and the truth is not in him.
1JOHN|2|5|But if anyone obeys his word, God's love is truly made complete in him. This is how we know we are in him:
1JOHN|2|6|Whoever claims to live in him must walk as Jesus did.
1JOHN|2|7|Dear friends, I am not writing you a new command but an old one, which you have had since the beginning. This old command is the message you have heard.
1JOHN|2|8|Yet I am writing you a new command; its truth is seen in him and you, because the darkness is passing and the true light is already shining.
1JOHN|2|9|Anyone who claims to be in the light but hates his brother is still in the darkness.
1JOHN|2|10|Whoever loves his brother lives in the light, and there is nothing in him to make him stumble.
1JOHN|2|11|But whoever hates his brother is in the darkness and walks around in the darkness; he does not know where he is going, because the darkness has blinded him.
1JOHN|2|12|I write to you, dear children, because your sins have been forgiven on account of his name.
1JOHN|2|13|I write to you, fathers, because you have known him who is from the beginning. I write to you, young men, because you have overcome the evil one. I write to you, dear children, because you have known the Father.
1JOHN|2|14|I write to you, fathers, because you have known him who is from the beginning. I write to you, young men, because you are strong, and the word of God lives in you, and you have overcome the evil one.
1JOHN|2|15|Do not love the world or anything in the world. If anyone loves the world, the love of the Father is not in him.
1JOHN|2|16|For everything in the world--the cravings of sinful man, the lust of his eyes and the boasting of what he has and does--comes not from the Father but from the world.
1JOHN|2|17|The world and its desires pass away, but the man who does the will of God lives forever.
1JOHN|2|18|Dear children, this is the last hour; and as you have heard that the antichrist is coming, even now many antichrists have come. This is how we know it is the last hour.
1JOHN|2|19|They went out from us, but they did not really belong to us. For if they had belonged to us, they would have remained with us; but their going showed that none of them belonged to us.
1JOHN|2|20|But you have an anointing from the Holy One, and all of you know the truth.
1JOHN|2|21|I do not write to you because you do not know the truth, but because you do know it and because no lie comes from the truth.
1JOHN|2|22|Who is the liar? It is the man who denies that Jesus is the Christ. Such a man is the antichrist--he denies the Father and the Son.
1JOHN|2|23|No one who denies the Son has the Father; whoever acknowledges the Son has the Father also.
1JOHN|2|24|See that what you have heard from the beginning remains in you. If it does, you also will remain in the Son and in the Father.
1JOHN|2|25|And this is what he promised us--even eternal life.
1JOHN|2|26|I am writing these things to you about those who are trying to lead you astray.
1JOHN|2|27|As for you, the anointing you received from him remains in you, and you do not need anyone to teach you. But as his anointing teaches you about all things and as that anointing is real, not counterfeit--just as it has taught you, remain in him.
1JOHN|2|28|And now, dear children, continue in him, so that when he appears we may be confident and unashamed before him at his coming.
1JOHN|2|29|If you know that he is righteous, you know that everyone who does what is right has been born of him.
1JOHN|3|1|How great is the love the Father has lavished on us, that we should be called children of God! And that is what we are! The reason the world does not know us is that it did not know him.
1JOHN|3|2|Dear friends, now we are children of God, and what we will be has not yet been made known. But we know that when he appears, we shall be like him, for we shall see him as he is.
1JOHN|3|3|Everyone who has this hope in him purifies himself, just as he is pure.
1JOHN|3|4|Everyone who sins breaks the law; in fact, sin is lawlessness.
1JOHN|3|5|But you know that he appeared so that he might take away our sins. And in him is no sin.
1JOHN|3|6|No one who lives in him keeps on sinning. No one who continues to sin has either seen him or known him.
1JOHN|3|7|Dear children, do not let anyone lead you astray. He who does what is right is righteous, just as he is righteous.
1JOHN|3|8|He who does what is sinful is of the devil, because the devil has been sinning from the beginning. The reason the Son of God appeared was to destroy the devil's work.
1JOHN|3|9|No one who is born of God will continue to sin, because God's seed remains in him; he cannot go on sinning, because he has been born of God.
1JOHN|3|10|This is how we know who the children of God are and who the children of the devil are: Anyone who does not do what is right is not a child of God; nor is anyone who does not love his brother.
1JOHN|3|11|This is the message you heard from the beginning: We should love one another.
1JOHN|3|12|Do not be like Cain, who belonged to the evil one and murdered his brother. And why did he murder him? Because his own actions were evil and his brother's were righteous.
1JOHN|3|13|Do not be surprised, my brothers, if the world hates you.
1JOHN|3|14|We know that we have passed from death to life, because we love our brothers. Anyone who does not love remains in death.
1JOHN|3|15|Anyone who hates his brother is a murderer, and you know that no murderer has eternal life in him.
1JOHN|3|16|This is how we know what love is: Jesus Christ laid down his life for us. And we ought to lay down our lives for our brothers.
1JOHN|3|17|If anyone has material possessions and sees his brother in need but has no pity on him, how can the love of God be in him?
1JOHN|3|18|Dear children, let us not love with words or tongue but with actions and in truth.
1JOHN|3|19|This then is how we know that we belong to the truth, and how we set our hearts at rest in his presence
1JOHN|3|20|whenever our hearts condemn us. For God is greater than our hearts, and he knows everything.
1JOHN|3|21|Dear friends, if our hearts do not condemn us, we have confidence before God
1JOHN|3|22|and receive from him anything we ask, because we obey his commands and do what pleases him.
1JOHN|3|23|And this is his command: to believe in the name of his Son, Jesus Christ, and to love one another as he commanded us.
1JOHN|3|24|Those who obey his commands live in him, and he in them. And this is how we know that he lives in us: We know it by the Spirit he gave us.
1JOHN|4|1|Dear friends, do not believe every spirit, but test the spirits to see whether they are from God, because many false prophets have gone out into the world.
1JOHN|4|2|This is how you can recognize the Spirit of God: Every spirit that acknowledges that Jesus Christ has come in the flesh is from God,
1JOHN|4|3|but every spirit that does not acknowledge Jesus is not from God. This is the spirit of the antichrist, which you have heard is coming and even now is already in the world.
1JOHN|4|4|You, dear children, are from God and have overcome them, because the one who is in you is greater than the one who is in the world.
1JOHN|4|5|They are from the world and therefore speak from the viewpoint of the world, and the world listens to them.
1JOHN|4|6|We are from God, and whoever knows God listens to us; but whoever is not from God does not listen to us. This is how we recognize the Spirit of truth and the spirit of falsehood.
1JOHN|4|7|Dear friends, let us love one another, for love comes from God. Everyone who loves has been born of God and knows God.
1JOHN|4|8|Whoever does not love does not know God, because God is love.
1JOHN|4|9|This is how God showed his love among us: He sent his one and only Son into the world that we might live through him.
1JOHN|4|10|This is love: not that we loved God, but that he loved us and sent his Son as an atoning sacrifice for our sins.
1JOHN|4|11|Dear friends, since God so loved us, we also ought to love one another.
1JOHN|4|12|No one has ever seen God; but if we love one another, God lives in us and his love is made complete in us.
1JOHN|4|13|We know that we live in him and he in us, because he has given us of his Spirit.
1JOHN|4|14|And we have seen and testify that the Father has sent his Son to be the Savior of the world.
1JOHN|4|15|If anyone acknowledges that Jesus is the Son of God, God lives in him and he in God.
1JOHN|4|16|And so we know and rely on the love God has for us. God is love. Whoever lives in love lives in God, and God in him.
1JOHN|4|17|In this way, love is made complete among us so that we will have confidence on the day of judgment, because in this world we are like him.
1JOHN|4|18|There is no fear in love. But perfect love drives out fear, because fear has to do with punishment. The one who fears is not made perfect in love.
1JOHN|4|19|We love because he first loved us.
1JOHN|4|20|If anyone says, "I love God," yet hates his brother, he is a liar. For anyone who does not love his brother, whom he has seen, cannot love God, whom he has not seen.
1JOHN|4|21|And he has given us this command: Whoever loves God must also love his brother.
1JOHN|5|1|Everyone who believes that Jesus is the Christ is born of God, and everyone who loves the father loves his child as well.
1JOHN|5|2|This is how we know that we love the children of God: by loving God and carrying out his commands.
1JOHN|5|3|This is love for God: to obey his commands. And his commands are not burdensome,
1JOHN|5|4|for everyone born of God overcomes the world. This is the victory that has overcome the world, even our faith.
1JOHN|5|5|Who is it that overcomes the world? Only he who believes that Jesus is the Son of God.
1JOHN|5|6|This is the one who came by water and blood--Jesus Christ. He did not come by water only, but by water and blood. And it is the Spirit who testifies, because the Spirit is the truth.
1JOHN|5|7|For there are three that testify:
1JOHN|5|8|the Spirit, the water and the blood; and the three are in agreement.
1JOHN|5|9|We accept man's testimony, but God's testimony is greater because it is the testimony of God, which he has given about his Son.
1JOHN|5|10|Anyone who believes in the Son of God has this testimony in his heart. Anyone who does not believe God has made him out to be a liar, because he has not believed the testimony God has given about his Son.
1JOHN|5|11|And this is the testimony: God has given us eternal life, and this life is in his Son.
1JOHN|5|12|He who has the Son has life; he who does not have the Son of God does not have life.
1JOHN|5|13|I write these things to you who believe in the name of the Son of God so that you may know that you have eternal life.
1JOHN|5|14|This is the confidence we have in approaching God: that if we ask anything according to his will, he hears us.
1JOHN|5|15|And if we know that he hears us--whatever we ask--we know that we have what we asked of him.
1JOHN|5|16|If anyone sees his brother commit a sin that does not lead to death, he should pray and God will give him life. I refer to those whose sin does not lead to death. There is a sin that leads to death. I am not saying that he should pray about that.
1JOHN|5|17|All wrongdoing is sin, and there is sin that does not lead to death.
1JOHN|5|18|We know that anyone born of God does not continue to sin; the one who was born of God keeps him safe, and the evil one cannot harm him.
1JOHN|5|19|We know that we are children of God, and that the whole world is under the control of the evil one.
1JOHN|5|20|We know also that the Son of God has come and has given us understanding, so that we may know him who is true. And we are in him who is true--even in his Son Jesus Christ. He is the true God and eternal life.
1JOHN|5|21|Dear children, keep yourselves from idols.
