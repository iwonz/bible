EPH|1|1|Paul, an apostle of Christ Jesus by the will of God, To the saints in Ephesus, the faithful in Christ Jesus:
EPH|1|2|Grace and peace to you from God our Father and the Lord Jesus Christ.
EPH|1|3|Praise be to the God and Father of our Lord Jesus Christ, who has blessed us in the heavenly realms with every spiritual blessing in Christ.
EPH|1|4|For he chose us in him before the creation of the world to be holy and blameless in his sight. In love
EPH|1|5|he predestined us to be adopted as his sons through Jesus Christ, in accordance with his pleasure and will--
EPH|1|6|to the praise of his glorious grace, which he has freely given us in the One he loves.
EPH|1|7|In him we have redemption through his blood, the forgiveness of sins, in accordance with the riches of God's grace
EPH|1|8|that he lavished on us with all wisdom and understanding.
EPH|1|9|And he made known to us the mystery of his will according to his good pleasure, which he purposed in Christ,
EPH|1|10|to be put into effect when the times will have reached their fulfillment--to bring all things in heaven and on earth together under one head, even Christ.
EPH|1|11|In him we were also chosen, having been predestined according to the plan of him who works out everything in conformity with the purpose of his will,
EPH|1|12|in order that we, who were the first to hope in Christ, might be for the praise of his glory.
EPH|1|13|And you also were included in Christ when you heard the word of truth, the gospel of your salvation. Having believed, you were marked in him with a seal, the promised Holy Spirit,
EPH|1|14|who is a deposit guaranteeing our inheritance until the redemption of those who are God's possession--to the praise of his glory.
EPH|1|15|For this reason, ever since I heard about your faith in the Lord Jesus and your love for all the saints,
EPH|1|16|I have not stopped giving thanks for you, remembering you in my prayers.
EPH|1|17|I keep asking that the God of our Lord Jesus Christ, the glorious Father, may give you the Spirit of wisdom and revelation, so that you may know him better.
EPH|1|18|I pray also that the eyes of your heart may be enlightened in order that you may know the hope to which he has called you, the riches of his glorious inheritance in the saints,
EPH|1|19|and his incomparably great power for us who believe. That power is like the working of his mighty strength,
EPH|1|20|which he exerted in Christ when he raised him from the dead and seated him at his right hand in the heavenly realms,
EPH|1|21|far above all rule and authority, power and dominion, and every title that can be given, not only in the present age but also in the one to come.
EPH|1|22|And God placed all things under his feet and appointed him to be head over everything for the church,
EPH|1|23|which is his body, the fullness of him who fills everything in every way.
EPH|2|1|As for you, you were dead in your transgressions and sins,
EPH|2|2|in which you used to live when you followed the ways of this world and of the ruler of the kingdom of the air, the spirit who is now at work in those who are disobedient.
EPH|2|3|All of us also lived among them at one time, gratifying the cravings of our sinful nature and following its desires and thoughts. Like the rest, we were by nature objects of wrath.
EPH|2|4|But because of his great love for us, God, who is rich in mercy,
EPH|2|5|made us alive with Christ even when we were dead in transgressions--it is by grace you have been saved.
EPH|2|6|And God raised us up with Christ and seated us with him in the heavenly realms in Christ Jesus,
EPH|2|7|in order that in the coming ages he might show the incomparable riches of his grace, expressed in his kindness to us in Christ Jesus.
EPH|2|8|For it is by grace you have been saved, through faith--and this not from yourselves, it is the gift of God--
EPH|2|9|not by works, so that no one can boast.
EPH|2|10|For we are God's workmanship, created in Christ Jesus to do good works, which God prepared in advance for us to do.
EPH|2|11|Therefore, remember that formerly you who are Gentiles by birth and called "uncircumcised" by those who call themselves "the circumcision" (that done in the body by the hands of men)--
EPH|2|12|remember that at that time you were separate from Christ, excluded from citizenship in Israel and foreigners to the covenants of the promise, without hope and without God in the world.
EPH|2|13|But now in Christ Jesus you who once were far away have been brought near through the blood of Christ.
EPH|2|14|For he himself is our peace, who has made the two one and has destroyed the barrier, the dividing wall of hostility,
EPH|2|15|by abolishing in his flesh the law with its commandments and regulations. His purpose was to create in himself one new man out of the two, thus making peace,
EPH|2|16|and in this one body to reconcile both of them to God through the cross, by which he put to death their hostility.
EPH|2|17|He came and preached peace to you who were far away and peace to those who were near.
EPH|2|18|For through him we both have access to the Father by one Spirit.
EPH|2|19|Consequently, you are no longer foreigners and aliens, but fellow citizens with God's people and members of God's household,
EPH|2|20|built on the foundation of the apostles and prophets, with Christ Jesus himself as the chief cornerstone.
EPH|2|21|In him the whole building is joined together and rises to become a holy temple in the Lord.
EPH|2|22|And in him you too are being built together to become a dwelling in which God lives by his Spirit.
EPH|3|1|For this reason I, Paul, the prisoner of Christ Jesus for the sake of you Gentiles--
EPH|3|2|Surely you have heard about the administration of God's grace that was given to me for you,
EPH|3|3|that is, the mystery made known to me by revelation, as I have already written briefly.
EPH|3|4|In reading this, then, you will be able to understand my insight into the mystery of Christ,
EPH|3|5|which was not made known to men in other generations as it has now been revealed by the Spirit to God's holy apostles and prophets.
EPH|3|6|This mystery is that through the gospel the Gentiles are heirs together with Israel, members together of one body, and sharers together in the promise in Christ Jesus.
EPH|3|7|I became a servant of this gospel by the gift of God's grace given me through the working of his power.
EPH|3|8|Although I am less than the least of all God's people, this grace was given me: to preach to the Gentiles the unsearchable riches of Christ,
EPH|3|9|and to make plain to everyone the administration of this mystery, which for ages past was kept hidden in God, who created all things.
EPH|3|10|His intent was that now, through the church, the manifold wisdom of God should be made known to the rulers and authorities in the heavenly realms,
EPH|3|11|according to his eternal purpose which he accomplished in Christ Jesus our Lord.
EPH|3|12|In him and through faith in him we may approach God with freedom and confidence.
EPH|3|13|I ask you, therefore, not to be discouraged because of my sufferings for you, which are your glory.
EPH|3|14|For this reason I kneel before the Father,
EPH|3|15|from whom his whole family in heaven and on earth derives its name.
EPH|3|16|I pray that out of his glorious riches he may strengthen you with power through his Spirit in your inner being,
EPH|3|17|so that Christ may dwell in your hearts through faith. And I pray that you, being rooted and established in love,
EPH|3|18|may have power, together with all the saints, to grasp how wide and long and high and deep is the love of Christ,
EPH|3|19|and to know this love that surpasses knowledge--that you may be filled to the measure of all the fullness of God.
EPH|3|20|Now to him who is able to do immeasurably more than all we ask or imagine, according to his power that is at work within us,
EPH|3|21|to him be glory in the church and in Christ Jesus throughout all generations, for ever and ever! Amen.
EPH|4|1|As a prisoner for the Lord, then, I urge you to live a life worthy of the calling you have received.
EPH|4|2|Be completely humble and gentle; be patient, bearing with one another in love.
EPH|4|3|Make every effort to keep the unity of the Spirit through the bond of peace.
EPH|4|4|There is one body and one Spirit--just as you were called to one hope when you were called--
EPH|4|5|one Lord, one faith, one baptism;
EPH|4|6|one God and Father of all, who is over all and through all and in all.
EPH|4|7|But to each one of us grace has been given as Christ apportioned it.
EPH|4|8|This is why it says: "When he ascended on high, he led captives in his train and gave gifts to men."
EPH|4|9|(What does "he ascended" mean except that he also descended to the lower, earthly regions?
EPH|4|10|He who descended is the very one who ascended higher than all the heavens, in order to fill the whole universe.)
EPH|4|11|It was he who gave some to be apostles, some to be prophets, some to be evangelists, and some to be pastors and teachers,
EPH|4|12|to prepare God's people for works of service, so that the body of Christ may be built up
EPH|4|13|until we all reach unity in the faith and in the knowledge of the Son of God and become mature, attaining to the whole measure of the fullness of Christ.
EPH|4|14|Then we will no longer be infants, tossed back and forth by the waves, and blown here and there by every wind of teaching and by the cunning and craftiness of men in their deceitful scheming.
EPH|4|15|Instead, speaking the truth in love, we will in all things grow up into him who is the Head, that is, Christ.
EPH|4|16|From him the whole body, joined and held together by every supporting ligament, grows and builds itself up in love, as each part does its work.
EPH|4|17|So I tell you this, and insist on it in the Lord, that you must no longer live as the Gentiles do, in the futility of their thinking.
EPH|4|18|They are darkened in their understanding and separated from the life of God because of the ignorance that is in them due to the hardening of their hearts.
EPH|4|19|Having lost all sensitivity, they have given themselves over to sensuality so as to indulge in every kind of impurity, with a continual lust for more.
EPH|4|20|You, however, did not come to know Christ that way.
EPH|4|21|Surely you heard of him and were taught in him in accordance with the truth that is in Jesus.
EPH|4|22|You were taught, with regard to your former way of life, to put off your old self, which is being corrupted by its deceitful desires;
EPH|4|23|to be made new in the attitude of your minds;
EPH|4|24|and to put on the new self, created to be like God in true righteousness and holiness.
EPH|4|25|Therefore each of you must put off falsehood and speak truthfully to his neighbor, for we are all members of one body.
EPH|4|26|"In your anger do not sin": Do not let the sun go down while you are still angry,
EPH|4|27|and do not give the devil a foothold.
EPH|4|28|He who has been stealing must steal no longer, but must work, doing something useful with his own hands, that he may have something to share with those in need.
EPH|4|29|Do not let any unwholesome talk come out of your mouths, but only what is helpful for building others up according to their needs, that it may benefit those who listen.
EPH|4|30|And do not grieve the Holy Spirit of God, with whom you were sealed for the day of redemption.
EPH|4|31|Get rid of all bitterness, rage and anger, brawling and slander, along with every form of malice.
EPH|4|32|Be kind and compassionate to one another, forgiving each other, just as in Christ God forgave you.
EPH|5|1|Be imitators of God, therefore, as dearly loved children
EPH|5|2|and live a life of love, just as Christ loved us and gave himself up for us as a fragrant offering and sacrifice to God.
EPH|5|3|But among you there must not be even a hint of sexual immorality, or of any kind of impurity, or of greed, because these are improper for God's holy people.
EPH|5|4|Nor should there be obscenity, foolish talk or coarse joking, which are out of place, but rather thanksgiving.
EPH|5|5|For of this you can be sure: No immoral, impure or greedy person--such a man is an idolater--has any inheritance in the kingdom of Christ and of God.
EPH|5|6|Let no one deceive you with empty words, for because of such things God's wrath comes on those who are disobedient.
EPH|5|7|Therefore do not be partners with them.
EPH|5|8|For you were once darkness, but now you are light in the Lord. Live as children of light
EPH|5|9|(for the fruit of the light consists in all goodness, righteousness and truth)
EPH|5|10|and find out what pleases the Lord.
EPH|5|11|Have nothing to do with the fruitless deeds of darkness, but rather expose them.
EPH|5|12|For it is shameful even to mention what the disobedient do in secret.
EPH|5|13|But everything exposed by the light becomes visible,
EPH|5|14|for it is light that makes everything visible. This is why it is said: "Wake up, O sleeper, rise from the dead, and Christ will shine on you."
EPH|5|15|Be very careful, then, how you live--not as unwise but as wise,
EPH|5|16|making the most of every opportunity, because the days are evil.
EPH|5|17|Therefore do not be foolish, but understand what the Lord's will is.
EPH|5|18|Do not get drunk on wine, which leads to debauchery. Instead, be filled with the Spirit.
EPH|5|19|Speak to one another with psalms, hymns and spiritual songs. Sing and make music in your heart to the Lord,
EPH|5|20|always giving thanks to God the Father for everything, in the name of our Lord Jesus Christ.
EPH|5|21|Submit to one another out of reverence for Christ.
EPH|5|22|Wives, submit to your husbands as to the Lord.
EPH|5|23|For the husband is the head of the wife as Christ is the head of the church, his body, of which he is the Savior.
EPH|5|24|Now as the church submits to Christ, so also wives should submit to their husbands in everything.
EPH|5|25|Husbands, love your wives, just as Christ loved the church and gave himself up for her
EPH|5|26|to make her holy, cleansing her by the washing with water through the word,
EPH|5|27|and to present her to himself as a radiant church, without stain or wrinkle or any other blemish, but holy and blameless.
EPH|5|28|In this same way, husbands ought to love their wives as their own bodies. He who loves his wife loves himself.
EPH|5|29|After all, no one ever hated his own body, but he feeds and cares for it, just as Christ does the church--
EPH|5|30|for we are members of his body.
EPH|5|31|"For this reason a man will leave his father and mother and be united to his wife, and the two will become one flesh."
EPH|5|32|This is a profound mystery--but I am talking about Christ and the church.
EPH|5|33|However, each one of you also must love his wife as he loves himself, and the wife must respect her husband.
EPH|6|1|Children, obey your parents in the Lord, for this is right.
EPH|6|2|"Honor your father and mother"--which is the first commandment with a promise--
EPH|6|3|"that it may go well with you and that you may enjoy long life on the earth."
EPH|6|4|Fathers, do not exasperate your children; instead, bring them up in the training and instruction of the Lord.
EPH|6|5|Slaves, obey your earthly masters with respect and fear, and with sincerity of heart, just as you would obey Christ.
EPH|6|6|Obey them not only to win their favor when their eye is on you, but like slaves of Christ, doing the will of God from your heart.
EPH|6|7|Serve wholeheartedly, as if you were serving the Lord, not men,
EPH|6|8|because you know that the Lord will reward everyone for whatever good he does, whether he is slave or free.
EPH|6|9|And masters, treat your slaves in the same way. Do not threaten them, since you know that he who is both their Master and yours is in heaven, and there is no favoritism with him.
EPH|6|10|Finally, be strong in the Lord and in his mighty power.
EPH|6|11|Put on the full armor of God so that you can take your stand against the devil's schemes.
EPH|6|12|For our struggle is not against flesh and blood, but against the rulers, against the authorities, against the powers of this dark world and against the spiritual forces of evil in the heavenly realms.
EPH|6|13|Therefore put on the full armor of God, so that when the day of evil comes, you may be able to stand your ground, and after you have done everything, to stand.
EPH|6|14|Stand firm then, with the belt of truth buckled around your waist, with the breastplate of righteousness in place,
EPH|6|15|and with your feet fitted with the readiness that comes from the gospel of peace.
EPH|6|16|In addition to all this, take up the shield of faith, with which you can extinguish all the flaming arrows of the evil one.
EPH|6|17|Take the helmet of salvation and the sword of the Spirit, which is the word of God.
EPH|6|18|And pray in the Spirit on all occasions with all kinds of prayers and requests. With this in mind, be alert and always keep on praying for all the saints.
EPH|6|19|Pray also for me, that whenever I open my mouth, words may be given me so that I will fearlessly make known the mystery of the gospel,
EPH|6|20|for which I am an ambassador in chains. Pray that I may declare it fearlessly, as I should.
EPH|6|21|Tychicus, the dear brother and faithful servant in the Lord, will tell you everything, so that you also may know how I am and what I am doing.
EPH|6|22|I am sending him to you for this very purpose, that you may know how we are, and that he may encourage you.
EPH|6|23|Peace to the brothers, and love with faith from God the Father and the Lord Jesus Christ.
EPH|6|24|Grace to all who love our Lord Jesus Christ with an undying love.
