PHLM|1|1|Paul, a prisoner of Christ Jesus, and Timothy our brother,
PHLM|1|2|To Philemon our dear friend and fellow worker, to Apphia our sister, to Archippus our fellow soldier and to the church that meets in your home:
PHLM|1|3|Grace to you and peace from God our Father and the Lord Jesus Christ.
PHLM|1|4|I always thank my God as I remember you in my prayers,
PHLM|1|5|because I hear about your faith in the Lord Jesus and your love for all the saints.
PHLM|1|6|I pray that you may be active in sharing your faith, so that you will have a full understanding of every good thing we have in Christ.
PHLM|1|7|Your love has given me great joy and encouragement, because you, brother, have refreshed the hearts of the saints.
PHLM|1|8|Therefore, although in Christ I could be bold and order you to do what you ought to do,
PHLM|1|9|yet I appeal to you on the basis of love. I then, as Paul--an old man and now also a prisoner of Christ Jesus--
PHLM|1|10|I appeal to you for my son Onesimus, who became my son while I was in chains.
PHLM|1|11|Formerly he was useless to you, but now he has become useful both to you and to me.
PHLM|1|12|I am sending him--who is my very heart--back to you.
PHLM|1|13|I would have liked to keep him with me so that he could take your place in helping me while I am in chains for the gospel.
PHLM|1|14|But I did not want to do anything without your consent, so that any favor you do will be spontaneous and not forced.
PHLM|1|15|Perhaps the reason he was separated from you for a little while was that you might have him back for good--
PHLM|1|16|no longer as a slave, but better than a slave, as a dear brother. He is very dear to me but even dearer to you, both as a man and as a brother in the Lord.
PHLM|1|17|So if you consider me a partner, welcome him as you would welcome me.
PHLM|1|18|If he has done you any wrong or owes you anything, charge it to me.
PHLM|1|19|I, Paul, am writing this with my own hand. I will pay it back--not to mention that you owe me your very self.
PHLM|1|20|I do wish, brother, that I may have some benefit from you in the Lord; refresh my heart in Christ.
PHLM|1|21|Confident of your obedience, I write to you, knowing that you will do even more than I ask.
PHLM|1|22|And one thing more: Prepare a guest room for me, because I hope to be restored to you in answer to your prayers.
PHLM|1|23|Epaphras, my fellow prisoner in Christ Jesus, sends you greetings.
PHLM|1|24|And so do Mark, Aristarchus, Demas and Luke, my fellow workers.
PHLM|1|25|The grace of the Lord Jesus Christ be with your spirit.
