REV|1|1|Об'явлення Ісуса Христа, яке дав Йому Бог, щоб показати Своїм рабам, що незабаром статися має. І Він показав, і послав Своїм Анголом рабові Своєму Іванові,
REV|1|2|який свідчив про Слово Боже, і про свідчення Ісуса Христа, і про все, що він бачив.
REV|1|3|Блаженний, хто читає, і ті, хто слухає слова пророцтва та додержує написане в ньому, час бо близький!
REV|1|4|Іван до семи Церков, що в Азії: благодать вам і мир від Того, Хто є, Хто був і Хто має прийти; і від семи духів, що перед престолом Його,
REV|1|5|та від Ісуса Христа, а Він Свідок вірний, Первенець з мертвих і Владика земних царів. Йому, що нас полюбив і кров'ю Своєю обмив нас від наших гріхів,
REV|1|6|що вчинив нас царями, священиками Богові й Отцеві Своєму, Тому слава та сила на вічні віки! Амінь.
REV|1|7|Ото Він із хмарами йде, і побачить Його кожне око, і ті, що Його прокололи були, і всі племена землі будуть плакати за Ним. Так, амінь!
REV|1|8|Я Альфа й Омега, говорить Господь, Бог, Той, Хто є, і Хто був, і Хто має прийти, Вседержитель!
REV|1|9|Я, Іван, ваш брат і спільник у біді, і в царстві, і в терпінні в Ісусі, був на острові, що зветься Патмос, за Слово Боже і за свідчення Ісуса Христа.
REV|1|10|Я був у дусі Господнього дня, і почув за собою голос гучний, немов сурми,
REV|1|11|який говорив: Що бачиш, напиши те до книги, і пошли до сімох Церков: до Ефесу, і до Смірни, і до Пергаму, і до Тіятирів, і до Сард, і до Філядельфії, і до Лаодикії.
REV|1|12|І я оглянувся, щоб побачити голос, що говорив зо мною. І, оглянувшись, я побачив сім свічників золотих;
REV|1|13|а посеред семи свічників Подібного до Людського Сина, одягненого в довгу одежу і підперезаного по грудях золотим поясом.
REV|1|14|А Його голова та волосся білі, немов біла вовна, як сніг; а очі Його немов полум'я огняне.
REV|1|15|А ноги Його подібні до міді, розпалені, наче в печі; а голос Його немов шум великої води.
REV|1|16|І сім зір Він держав у правиці Своїй, а з уст Його меч обосічний виходив, а обличчя Його, немов сонце, що світить у силі своїй.
REV|1|17|І коли я побачив Його, то до ніг Йому впав, немов мертвий. І поклав Він на мене правицю Свою та й промовив мені: Не лякайся! Я Перший і Останній,
REV|1|18|і Живий. І був Я мертвий, а ось Я Живий на вічні віки. І маю ключі Я від смерти й від аду.
REV|1|19|Отже, напиши, що ти бачив, і що є, і що має бути по цьому!
REV|1|20|Таємниця семи зір, що бачив ти їх на правиці Моїй, і семи свічників золотих: сім зір, то Анголи семи Церков, а сім свічників, що ти бачив, то сім Церков.
REV|2|1|До Ангола Церкви в Ефесі напиши: Оце каже Той, Хто тримає сім зір у правиці Своїй, Хто ходить серед семи свічників золотих:
REV|2|2|Я знаю діла твої, і працю твою, і твою терпеливість, і що не можеш терпіти лихих, і випробував тих, хто себе називає апостолами, але ними не є, і знайшов, що фальшиві вони.
REV|2|3|І ти маєш терпіння, і працював для Ймення Мого, але не знемігся.
REV|2|4|Але маю на тебе, що ти покинув свою першу любов.
REV|2|5|Отож, пам'ятай, звідки ти впав, і покайся, і вчинки давніші роби. Коли ж ні, то до тебе прийду незабаром, і зрушу твого свічника з його місця, якщо не покаєшся.
REV|2|6|Але маєш оце, що ненавидиш учинки Николаїтів, яких і Я ненавиджу.
REV|2|7|Хто має вухо, хай чує, що Дух промовляє Церквам: переможцеві дам їсти від дерева життя, яке в раю Божім.
REV|2|8|А до Ангола Церкви в Смірні напиши: Оце каже Перший й Останній, що був мертвий й ожив:
REV|2|9|Я знаю діла твої, і біду, і убозтво, але ти багатий, і зневагу тих, що говорять про себе, ніби юдеї вони, та ними не є, але вони зборище сатани.
REV|2|10|Не бійся того, що маєш страждати! Ось диявол вкидатиме декого з вас до в'язниць, щоб вас випробувати. І будете мати біду десять день. Будь вірний до смерти, і Я тобі дам вінця життя!
REV|2|11|Хто має вухо, хай чує, що Дух промовляє Церквам: переможець не буде пошкоджений від другої смерти.
REV|2|12|А до Ангола Церкви в Пергамі напиши: Оце каже Той, що має меча обосічного:
REV|2|13|Я знаю діла твої, і що де ти живеш, там престол сатани. І тримаєш ти Ймення Моє, і ти не відкинувся від віри Моєї навіть за днів, коли в вас, де живе сатана, був убитий Антипа, свідок Мій вірний.
REV|2|14|Але трохи Я маю на тебе, бо маєш там тих, хто тримається науки Валаама, що навчав був Балака покласти спотикання перед синами Ізраїля, щоб їли ідольські жертви й розпусту чинили.
REV|2|15|Так маєш і ти таких, що тримаються науки Николаїтської так само.
REV|2|16|Тож покайся! Коли ж ні, то до тебе прийду незабаром, і воюватиму з ними мечем Своїх уст.
REV|2|17|Хто має вухо, хай чує, що Дух промовляє Церквам: переможцеві дам їсти приховану манну, і дам йому білого каменя, а на камені написане ймення нове, якого не знає ніхто, тільки той, хто приймає його.
REV|2|18|І до Ангола Церкви в Тіятирах напиши: Оце каже Син Божий, що має очі Свої, як полум'я огняне, а ноги Його подібні до міді:
REV|2|19|Я знаю діла твої, і любов, і віру, і службу, і твою терпеливість, і останні вчинки твої, що більші за перші.
REV|2|20|Але маю на тебе, що жінці Єзавелі, яка каже, ніби вона пророкиня, ти попускаєш навчати та зводити рабів Моїх, чинити розпусту та їсти ідольські жертви.
REV|2|21|І Я дав був їй часу, щоб покаялася, та вона не схотіла покаятися в розпусті своїй.
REV|2|22|Ось Я кину її на ложе, а тих, що чинять із нею розпусту, у велику біду, коли тільки в учинках своїх не покаються,
REV|2|23|а діти її поб'ю смертю. І пізнають усі Церкви, що Я Той, Хто нирки й серця вивіряє, і Я кожному з вас дам за вчинками вашими.
REV|2|24|А вам, та іншим, що в Тіятирах, що не мають науки цієї, і як кажуть не розуміють так званих глибин сатани, кажу: не накладу на вас іншого тягару,
REV|2|25|тільки те, що ви маєте, тримайте, аж поки прийду.
REV|2|26|А переможцеві, і тому, хто аж до кінця додержує Мої вчинки, Я дам йому владу над поганами,
REV|2|27|і буде пасти їх залізним жезлом; вони, немов глиняний посуд, покрушаться, як і Я одержав владу від Свого Отця,
REV|2|28|і дам Я йому зорю досвітню.
REV|2|29|Хто має вухо, хай чує, що Дух промовляє Церквам!
REV|3|1|А до Ангола Церкви в Сардах напиши: Оце каже Той, Хто має сім Божих духів і сім зір: Я знаю діла твої, що маєш ім'я, ніби живий, а ти мертвий.
REV|3|2|Будь чуйний та решту зміцняй, що мають померти. Бо Я не знайшов твоїх діл закінченими перед Богом Моїм.
REV|3|3|Отож, пам'ятай, як ти взяв і почув, і бережи, і покайся. А коли ти не чуйний, то на тебе прийду, немов злодій, і ти знати не будеш, якої години на тебе прийду.
REV|3|4|Та ти маєш і в Сардах кілька імен, що одежі своєї вони не споганили, і в білій зо Мною ходитимуть, бо гідні вони.
REV|3|5|Переможець зодягнеться в білу одежу, а ймення його Я не змию із книги життя, і ймення його визнаю перед Отцем Своїм і перед Його Анголами.
REV|3|6|Хто має вухо, хай чує, що Дух промовляє Церквам!
REV|3|7|І до Ангола Церкви в Філядельфії напиши: Оце каже Святий, Правдивий, що має ключа Давидового, що Він відчиняє, і ніхто не зачинить, що Він зачиняє, і ніхто не відчинить.
REV|3|8|Я знаю діла твої. Ось Я перед тобою дверей не зачинив, і їх зачинити не може ніхто. Хоч малу маєш силу, але слово Моє ти зберіг, і від Ймення Мого не відкинувся.
REV|3|9|Ось Я зроблю, що декого з зборища сатани, із тих, що себе називають юдеями, та ними не є, але кажуть неправду, ось Я зроблю, що вони прийдуть та вклоняться перед ногами твоїми, і пізнають, що Я полюбив тебе.
REV|3|10|А що ти зберіг слово терпіння Мого, то й Я тебе збережу від години випробовування, що має прийти на ввесь всесвіт, щоб випробувати мешканців землі.
REV|3|11|Я прийду незабаром. Тримай, що ти маєш, щоб твого вінця ніхто не забрав.
REV|3|12|Переможця зроблю Я стовпом у храмі Бога Мого, і він вже не вийде назовні, і на нім напишу Ім'я Бога Мого й ім'я міста Бога Мого, Єрусалиму Нового, що з неба сходить від Бога Мого, та нове Ім'я Своє.
REV|3|13|Хто має вухо, хай чує, що Дух промовляє Церквам!
REV|3|14|І до Ангола Церкви в Лаодикії напиши: Оце каже Амінь, Свідок вірний і правдивий, початок Божого творива:
REV|3|15|Я знаю діла твої, що ти не холодний, ані гарячий. Якби то холодний чи гарячий ти був!
REV|3|16|А що ти літеплий, і ні гарячий, ані холодний, то виплюну тебе з Своїх уст...
REV|3|17|Бо ти кажеш: Я багатий, і збагатів, і не потребую нічого. А не знаєш, що ти нужденний, і мізерний, і вбогий, і сліпий, і голий!
REV|3|18|Раджу тобі купити в Мене золота, в огні перечищеного, щоб збагатитись, і білу одежу, щоб зодягтися, і щоб ганьба наготи твоєї не видна була, а мастю на очі намасти свої очі, щоб бачити.
REV|3|19|Кого Я люблю, тому докоряю й караю того. Будь же ревний і покайся!
REV|3|20|Ось Я стою під дверима та стукаю: коли хто почує Мій голос і двері відчинить, Я до нього ввійду, і буду вечеряти з ним, а він зо Мною.
REV|3|21|Переможцеві сісти Я дам на Моєму престолі зо Мною, як і Я переміг був, і з Отцем Своїм сів на престолі Його.
REV|3|22|Хто має вухо, хай чує, що Дух промовляє Церквам!
REV|4|1|По цьому я поглянув, і ось двері на небі відчинені, і перший голос, що я чув його, як сурму, що зо мною говорив, сказав: Іди сюди, і Я тобі покажу, що статися має по цьому!
REV|4|2|І зараз у дусі я був. І ось престол стояв на небі, а на престолі Сидячий.
REV|4|3|А Сидячий подібний був з вигляду до каменя яспіса й сардиса, а веселка навколо престолу видом подібна була до смарагду.
REV|4|4|А навколо престолу двадцять чотири престоли, а на престолах я бачив двадцятьох чотирьох старців, що сиділи, у шати білі одягнені, а на головах своїх мали вінці золоті.
REV|4|5|А від престолу виходили блискавки, і голоси, і громи. А перед престолом горіли сім свічників огняних, а вони сім духів Божих.
REV|4|6|І перед престолом як море скляне, до кришталю подібне. А серед престолу й навколо престолу четверо тварин, повні очей спереду й ззаду.
REV|4|7|І перша тварина подібна до лева, а друга тварина подібна до теляти, а третя тварина мала лице, як людина, а четверта тварина подібна до орла, що летить.
REV|4|8|І ті чотири тварині, кожна з них мала навколо по шість крил, а всередині повна очей. І спокою не мають вони день і ніч, промовляючи: Свят, свят, свят Господь, Бог Вседержитель, що Він був, і що є, і що має прийти!
REV|4|9|І коли ті тварини складають славу, і честь, і подяку Тому, Хто сидить на престолі й живе віки вічні,
REV|4|10|тоді падають двадцять чотири старці перед Тим, Хто сидить на престолі, і вклоняються Тому, Хто живе віки вічні, і складають вінці свої перед престолом та кажуть:
REV|4|11|Достойний Ти, Господи й Боже наш, прийняти славу, і честь, і силу, бо все Ти створив, і з волі Твоєї існує та створене все!
REV|5|1|І я бачив в правиці Того, Хто сидить на престолі, книгу, написану всередині й назовні, і запечатану сімома печатками.
REV|5|2|І бачив я потужного Ангола, який гучним голосом кликав: Хто гідний розгорнути книгу, і зламати печатки її?
REV|5|3|І не міг ніхто ні на небі, ні на землі, ані під землею розгорнути книги, ані навіть зазирнути в неї.
REV|5|4|І плакав я гірко, що не знайшовся ані один гідний розгорнути й прочитати книгу, ані навіть зазирнути в неї.
REV|5|5|А один із старців промовив до мене: Не плач! Ось Лев, що з племени Юдиного, корень Давидів, переміг так, що може розгорнути книгу, і зламати сім печаток її.
REV|5|6|І я глянув, і ось серед престолу й чотирьох тварин і серед старців стоїть Агнець, як заколений, що має сім рогів і сім очей, а це сім Божих духів, посланих на всю землю.
REV|5|7|І Він підійшов, і взяв книгу з правиці Того, Хто сидить на престолі.
REV|5|8|А коли Він узяв книгу, то чотири тварині й двадцять чотири старці попадали перед Агнцем, а кожен мав гусла й золоті чаші, повні пахощів, а вони молитви святих.
REV|5|9|І нову пісню співають вони, промовляючи: Ти достойний узяти цю книгу, і розкрити печатки її, бо Ти був заколений, і кров'ю Своєю Ти викупив людей Богові з усякого племени, і язика, і народу, і люду.
REV|5|10|І Ти їх зробив для нашого Бога царями, і священиками, і вони на землі царюватимуть!
REV|5|11|І я бачив, і чув голос багатьох Анголів навколо престолу, і тварин, і старців, і число їх було десятки тисяч раз по десять тисяч і тисячі тисяч.
REV|5|12|І казали вони гучним голосом: Достойний Агнець, що заколений, прийняти силу, і багатство, і мудрість, і міць, і честь, і славу, і благословення!
REV|5|13|І кожне створіння, що воно на небі, і на землі, і під землею, і на морі, і все, що в них, чув я, говорило: Тому, Хто сидить на престолі, і Агнцеві благословення, і честь, і слава, і сила на вічні віки!
REV|5|14|А чотири тварині казали: Амінь! І двадцять чотири старці попадали та поклонились Тому, Хто живе повік віку!
REV|6|1|І я бачив, що Агнець розкрив одну з семи печаток, і почув я одну з чотирьох тих тварин, яка говорила, як голосом грому: Підійди!
REV|6|2|І я глянув, і ось кінь білий, а той, хто на ньому сидів, мав лука. І вінця йому дано, і він вийшов, немов переможець, і щоб перемогти.
REV|6|3|І коли другу печатку розкрив, я другу тварину почув, що казала: Підійди!
REV|6|4|І вийшов кінь другий, червоний. А тому, хто на ньому сидів, було дано взяти мир із землі та щоб убивали один одного. І меч великий був даний йому.
REV|6|5|І коли третю печатку розкрив, я третю тварину почув, що казала: Підійди! І я глянув, і ось кінь вороний. А той, хто на ньому сидів, мав вагу в своїй руці.
REV|6|6|І я ніби голос почув посеред чотирьох тих тварин, що казав: Ківш пшениці за динарія, і три ковші ячменю за динарія, а оливи й вина не марнуй!
REV|6|7|А коли Він четверту печатку розкрив, я четверту тварину почув, що казала: Підійди!
REV|6|8|І я глянув, і ось кінь чалий. А той, хто на ньому сидів, на ім'я йому Смерть, за ним же слідом ішов Ад. І дана їм влада була на четвертій частині землі забивати мечем, і голодом, і мором, і земними звірми.
REV|6|9|І коли п'яту печатку розкрив, я побачив під жертівником душі побитих за Боже Слово, і за свідчення, яке вони мали.
REV|6|10|І кликнули вони гучним голосом, кажучи: Аж доки, Владико святий та правдивий, не будеш судити, і не мститимеш тим, хто живе на землі, за кров нашу?
REV|6|11|І кожному з них дано білу одежу, і сказано їм іще трохи спочити, аж поки доповнять число їхні співслуги, і брати їхні, що будуть побиті, як і вони.
REV|6|12|І коли шосту печатку розкрив, я поглянув, і ось сталось велике трясіння землі, і сонце зчорніло, як міх волосяний, і ввесь місяць зробився, як кров...
REV|6|13|І на землю попадали зорі небесні, як фіґове дерево ронить свої недозрілі плоди, коли потрясе сильний вітер...
REV|6|14|І небо сховалось, згорнувшись, немов той сувій пергамену, і кожна гора, і кожен острів порушилися з своїх місць...
REV|6|15|І земні царі, і вельможі та тисячники, і багаті та сильні, і кожен раб та кожен вільний, поховались у печери та в скелі гірські,
REV|6|16|та й кажуть до гір та до скель: Поспадайте на нас, і позакривайте ви нас від лиця Того, Хто сидить на престолі, і від гніву Агнця!...
REV|6|17|Бо прийшов це великий день гніву Його, і хто встояти може?
REV|7|1|А по цьому я бачив чотирьох Анголів, що стояли на чотирьох кутах землі та тримали чотири земні вітри, щоб вітер не віяв на землю, ані на море, ані на жодне дерево.
REV|7|2|І бачив я іншого Ангола, що від схід сонця виходив, і мав печатку Бога Живого. І він гучним голосом крикнув до чотирьох Анголів, що їм дано пошкодити землі та морю,
REV|7|3|говорячи: Не шкодьте ані землі, ані морю, ані дереву, аж поки ми покладемо печатки рабам Бога нашого на їхніх чолах!
REV|7|4|І почув я число попечатаних: сто сорок чотири тисячі попечатаних від усіх племен Ізраїлевих синів:
REV|7|5|з племени Юдиного дванадцять тисяч попечатаних, з племени Рувимового дванадцять тисяч, з племени Ґадового дванадцять тисяч,
REV|7|6|з племени Асирового дванадцять тисяч, з племени Нефталимового дванадцять тисяч, з племени Манасіїного дванадцять тисяч,
REV|7|7|з племени Симеонового дванадцять тисяч, з племени Левіїного дванадцять тисяч, з племени Іссахарового дванадцять тисяч,
REV|7|8|з племени Завулонового дванадцять тисяч, з племени Йосипового дванадцять тисяч, з племени Веніяминового дванадцять тисяч попечатаних.
REV|7|9|Потому я глянув, і ось натовп великий, що його зрахувати не може ніхто, з усякого люду, і племен, і народів, і язиків, стояв перед престолом і перед Агнцем, зодягнені в білу одежу, а в їхніх руках було пальмове віття.
REV|7|10|І взивали вони гучним голосом, кажучи: Спасіння нашому Богові, що сидить на престолі, і Агнцеві!
REV|7|11|А всі Анголи стояли навколо престолу та старців і чотирьох тих тварин. І вони на обличчя попадали перед престолом, і вклонилися Богові,
REV|7|12|кажучи: Амінь! Благословення, і слава, і мудрість, і хвала, і честь, і сила, і міць нашому Богу на вічні віки! Амінь!
REV|7|13|І відповів один із старців, і до мене сказав: Оці, що зодягнені в білу одежу, хто вони й звідкіля поприходили?
REV|7|14|І сказав я йому: Мій пане, ти знаєш! Він же мені відказав: Це ті, що прийшли від великого горя, і випрали одіж свою, та вибілили її в крові Агнця...
REV|7|15|Тому то вони перед Божим престолом, і в храмі Його день і ніч Йому служать. А Той, Хто сидить на престолі, розтягне намета над ними.
REV|7|16|Вони голоду й спраги терпіти не будуть уже, і не буде палити їх сонце, ані спека яка.
REV|7|17|Бо Агнець, що серед престолу, буде їх пасти, і водитиме їх до джерел вод життя. І Бог кожну сльозу з очей їхніх зітре!
REV|8|1|І коли сьому печатку розкрив, німа тиша настала на небі десь на півгодини.
REV|8|2|І я бачив сімох Анголів, що стояли перед Богом. І дано було їм сім сурем.
REV|8|3|І прийшов другий Ангол, та й став перед жертівником із золотою кадильницею. І було йому дано багато кадила, щоб до молитов усіх святих додав на золотого жертівника, що перед престолом.
REV|8|4|І знявся дим кадильний з молитвами святих від руки Ангола перед Бога.
REV|8|5|А Ангол кадильницю взяв, і наповнив її огнем із жертівника, та й кинув на землю. І зчинилися громи, і гуркотнява, і блискавиці та трясіння землі...
REV|8|6|І сім Анголів, що мали сім сурем, приготувалися, щоб сурмити.
REV|8|7|І засурмив перший Ангол, і вчинилися град та огонь, перемішані з кров'ю, і впали на землю. І спалилась третина землі, і згоріла третина дерев, і всіляка зелена трава погоріла...
REV|8|8|І засурмив другий Ангол, і немов би велика гора, розпалена огнем, була вкинена в море. І третина моря зробилася кров'ю,
REV|8|9|і померла третина морського створіння, що мають життя, і загинула третина кораблів...
REV|8|10|І засурмив третій Ангол, і велика зоря спала з неба, палаючи, як смолоскип. І спала вона на третину річок та на водні джерела.
REV|8|11|А ймення зорі тій Полин. І стала третина води, як полин, і багато з людей повмирали з води, бо згіркла вона...
REV|8|12|І засурмив Ангол четвертий, і вдарено третину сонця, і третину місяця, і третину зір, щоб затьмилася їхня третина, щоб третина дня не світила, так само ж і ніч...
REV|8|13|І бачив, і чув я одного орла, що летів серед неба і кликав гучним голосом: Горе, горе, горе тим, хто живе на землі, від голосів сурмових позосталих трьох Анголів, що мають сурмити!...
REV|9|1|І засурмив п'ятий Ангол, і я бачив зорю, що спала із неба додолу. І їй даний був ключ від криниці безодньої.
REV|9|2|І вона відімкнула криницю безодню, і дим повалив із криниці, мов дим із великої печі. І затьмилося сонце й повітря від криничного диму...
REV|9|3|А з диму на землю вийшла сарана, і дано їй міць, як мають міць скорпіони земні.
REV|9|4|І наказано їй, щоб вона не шкодила земній траві, ані жадному зіллю, ані жадному дереву, але тільки тим людям, які на чолах не мають печатки Божої.
REV|9|5|І було дано їй, щоб їх не вбивати, але мучити п'ять місяців; а мука від неї, як мука від скорпіона, коли вкусить людину.
REV|9|6|І в ті дні люди смерти шукатимуть, та не знайдуть її! Померти вони захотять, та втече від них смерть!...
REV|9|7|А вигляд сарани був подібний до коней, на війну приготованих; а на головах у неї немов би вінки, подібні на золото, а обличчя її немов людські обличчя.
REV|9|8|І мала волосся як волосся жіноче, а її зуби були немов лев'ячі.
REV|9|9|І мала вона панцери, немов панцери залізні; а шум її крил немов шум колесниць, коли коней багато біжить на війну.
REV|9|10|І мала хвости, подібні до скорпіонових, та жала, а в неї в хвостах її влада п'ять місяців шкодити людям.
REV|9|11|І мала вона над собою царя, ангола безодні; йому по-єврейському ім'я Аваддон, а по-грецькому звався він Аполліон!
REV|9|12|Одне горе минуло! Ось за ним ще два горя надходять!
REV|9|13|І засурмив шостий Ангол, і я почув один голос із чотирьох рогів золотого жертівника, який перед Богом,
REV|9|14|що казав шостому Анголові, який мав сурму: Розв'яжи чотирьох Анголів, що пов'язані при великій річці Ефраті.
REV|9|15|І були порозв'язувані чотири Анголи, приготовані на годину, і на день, і на місяць, і на рік, щоб убили третину людей.
REV|9|16|А число кінного війська двадцять тисяч раз по десять тисяч; і я чув їхнє число.
REV|9|17|І так бачив я коней в видінні, а на них верхівців, що панцери мали огняні, і гіяцинтові, і сірчані. А голови в коней немов голови лев'ячі, а з їхнього рота виходив огонь, і дим, і сірка.
REV|9|18|І побита була третина людей від цих трьох поразок, від огню, і від диму, і від сірки, що виходили з їхніх ротів.
REV|9|19|Сила бо коней була в їхнім роті та в їхніх хвостах. А хвости їхні подібні до вужів, що мають голови, і ними вони шкоду чинять.
REV|9|20|А решта людей, що не вбита була цими поразками, не покаялася за діла своїх рук, щоб не кланятись демонам, ані ідолам золотим, і срібним, і мідяним, і кам'яним, і дерев'яним, що не можуть вони ані бачити, ані чути, ані ходити.
REV|9|21|І вони не покаялися в своїх убивствах, ані в чарах своїх, ні в розпусті своїй, ні в крадіжках своїх...
REV|10|1|І бачив я іншого потужного Ангола, що сходив із неба. Був одягнений в хмару, і над його головою веселка була, а обличчя його як стовпи огняні,
REV|10|2|і мав у руці своїй книжку розгорнену. І він поставив свою праву ногу на море, а ліву на землю,
REV|10|3|і закричав гучним голосом, як лев той ричить. І як він закричав, то заговорили сім громів голосами своїми.
REV|10|4|А як заговорили сім громів голосами своїми, я хотів був писати. Та я почув голос із неба, що до мене казав: Запечатай оте, що сім громів казали, і того не пиши!
REV|10|5|А Ангол, що я бачив його, як стояв він на морі й землі, зняв до неба правицю свою
REV|10|6|та й поклявся Живучим по вічні віки, Який створив небо та те, що на ньому, і землю та те, що на ній, і море й що в нім, що вже часу не буде,
REV|10|7|а дня голосу сьомого Ангола, коли він засурмить, довершиться Божа таємниця, як Він благовістив був Своїм рабам пророкам.
REV|10|8|І голос, що я чув його з неба, став знов говорити зо мною й казати: Піди, та візьми розгорнену книжку з руки Ангола, що стоїть на морі й землі.
REV|10|9|І пішов я до Ангола та й промовив йому, щоб дав мені книжку. А він мені каже: Візьми, і з'їж її! І гіркість учинить вона для твого живота, та в устах твоїх буде солодка, як мед.
REV|10|10|І я взяв з руки Ангола книжку та й з'їв її. І була вона в устах моїх, немов мед той, солодка. Та коли її з'їв, вона гіркість зробила в моїм животі...
REV|10|11|І сказали мені: Ти мусиш знову пророкувати про народи, і поган, і язики, і про багато царів.
REV|11|1|І дано тростину мені, подібну до палиці, і сказано: Устань, і зміряй храма Божого й жертівника, і тих, хто вклоняється в ньому.
REV|11|2|А двір, що за храмом, лиши та не міряй його, бо він даний поганам, і сорок два місяці будуть топтати вони святе місто.
REV|11|3|І звелю Я двом свідкам Своїм, і будуть вони пророкувати тисячу двісті й шістдесят день, зодягнені в волосяницю.
REV|11|4|Вони дві оливі та два свічники, що стоять перед Богом землі.
REV|11|5|І коли б хто схотів учинити їм кривду, то вийде огонь з їхніх уст, і поїсть ворогів їхніх. А коли хто захоче вчинити їм кривду, той отак мусить бути забитий.
REV|11|6|Вони мають владу небо замкнути, щоб за днів їхніх пророцтва не йшов дощ. І мають владу вони над водою, у кров обертати її, і вдарити землю всілякою карою, скільки разів вони схочуть.
REV|11|7|А коли вони скінчать свідоцтво своє, то звірина, що з безодні виходить, із ними війну поведе, і вона їх переможе та їх повбиває.
REV|11|8|І їхні трупи полишить на майдані великого міста, що зветься духовно Содом і Єгипет, де й Господь наш був розп'ятий.
REV|11|9|І багато з народів, і з племен, і з язиків, і з поган будуть дивитися півчверта дні на їхні трупи, не дозволять покласти в гроби їхніх трупів.
REV|11|10|А мешканці землі будуть тішитися та радіти над ними, і дарунки пошлють один одному, бо мучили ці два пророки мешканців землі.
REV|11|11|А по півчверта днях дух життя ввійшов у них від Бога, і вони повставали на ноги свої. І напав жах великий на тих, хто дивився на них!
REV|11|12|І почули вони гучний голос із неба, що їм говорив: Зійдіть сюди! І на небо зійшли вони в хмарі, і вороги їхні дивились на них.
REV|11|13|І тієї години зчинився страшний землетрус, і десята частина міста того завалилась... І в цім трусі загинуло сім тисяч людських імен, а решта обгорнена жахом була, і вони віддали славу Богу Небесному!...
REV|11|14|Друге горе минуло! Ото незабаром настане за ним третє горе!
REV|11|15|І засурмив сьомий Ангол, і на небі зчинились гучні голоси, що казали: Перейшло панування над світом до Господа нашого та до Христа Його, і Він зацарює на вічні віки!
REV|11|16|І двадцять чотири старці, що на престолах своїх перед Богом сидять, попадали на обличчя свої, та й уклонилися Богові,
REV|11|17|кажучи: Дяку складаємо Тобі, Господи, Боже Вседержителю, що Ти є й що Ти був, що прийняв Свою силу велику та й зацарював!
REV|11|18|А погани розлютилися, та гнів Твій прийшов, і час настав мертвих судити, і дати заплату рабам Твоїм, пророкам і святим, і тим, хто Ймення Твого боїться малим і великим, і знищити тих, хто нищить землю.
REV|11|19|І розкрився храм Божий на небі, і ковчег заповіту Його в Його храмі з'явився. І зчинилися блискавки, і гуркіт, і громи, і землетрус, і великий град...
REV|12|1|І з'явилась на небі велика ознака: Жінка, зодягнена в сонце, а під ногами її місяць, а на її голові вінок із дванадцяти зір.
REV|12|2|І вона мала в утробі, і кричала від болю, та муки терпіла від породу.
REV|12|3|І з'явилася інша ознака на небі, ось змій червоноогняний, великий, що мав сім голів та десять рогів, а на його головах сім вінців.
REV|12|4|Його хвіст змів третину зір із Неба та й кинув додолу. І змій стояв перед жінкою, що мала вродити, щоб з'їсти дитину її, коли вродить...
REV|12|5|І дитину вродила вона чоловічої статі, що всі народи має пасти залізним жезлом. І дитина її була взята до Бога, і до престолу Його.
REV|12|6|А жінка втекла на пустиню, де вона мала місце, від Бога для неї вготоване, щоб там годували її тисячу двісті шістдесят день.
REV|12|7|І сталась на небі війна: Михаїл та його Анголи вчинили зо змієм війну. І змій воював та його анголи,
REV|12|8|та не втрималися, і вже не знайшлося їм місця на небі.
REV|12|9|І скинений був змій великий, вуж стародавній, що зветься диявол і сатана, що зводить усесвіт, і скинений був він додолу, а з ним і його анголи були скинені.
REV|12|10|І я почув гучний голос на небі, який говорив: Тепер настало спасіння, і сила, і царство нашого Бога, і влада Христа Його, бо скинений той, хто братів наших скаржив, хто перед нашим Богом оскаржував їх день і ніч!
REV|12|11|І вони його перемогли кров'ю Агнця та словом свого засвідчення, і не полюбили життя свого навіть до смерти!
REV|12|12|Через це звеселися ти, небо, та ті, хто на нім пробуває! Горе землі та морю, до вас бо диявол зійшов, маючи лютість велику, знаючи, що короткий час має!
REV|12|13|А коли змій побачив, що додолу він скинений, то став переслідувати жінку, що вродила хлоп'я.
REV|12|14|І жінці дані були дві крилі великого орла, щоб від змія летіла в пустиню до місця свого, де будуть її годувати час, і часи, і півчасу.
REV|12|15|І пустив змій за жінкою з уст своїх воду, як річку, щоб річка схопила її.
REV|12|16|Та жінці земля помогла, і розкрила земля свої уста, та й випила річку, яку змій був пустив із своїх уст...
REV|12|17|І змій розлютувався на жінку, і пішов воювати з останком насіння її, що вони бережуть Божі заповіді та мають свідоцтво Ісусове.
REV|13|1|(12-18) І я став на морському піску. (13-1) І я бачив звірину, що виходила з моря, яка мала десять рогів та сім голів, а на рогах її було десять вінців, а на її головах богозневажні імена.
REV|13|2|А звірина, що я її бачив, подібна до рися була, а ноги її як ведмежі, а паща її немов лев'яча паща. І змій дав їй свою силу, і престола свого, і владу велику.
REV|13|3|А одна з її голів була ніби забита на смерть, але рана смертельна її вздоровилась. І вся земля дивувалась, слідкуючи за звіриною!
REV|13|4|І вклонилися змієві, що дав владу звірині. І вклонились звірині, говорячи: Хто до звірини подібний, і хто воювати з нею може?
REV|13|5|І їй дано уста, що говорили зухвале та богозневажне. І їй дано владу діяти сорок два місяці.
REV|13|6|І відкрила вона свої уста на зневагу проти Бога, щоб богозневажати Ім'я Його й оселю Його, та тих, хто на небі живе.
REV|13|7|І їй дано провадити війну зо святими, та їх перемогти. І їй дана влада над кожним племенем, і народом, і язиком, і людом.
REV|13|8|І їй вклоняться всі, хто живе на землі, що їхні імена не написані в книгах життя Агнця, заколеного від закладин світу.
REV|13|9|Коли має хто вухо, нехай слухає:
REV|13|10|Коли хто до полону веде, сам піде в полон. Коли хто мечем убиває, такий мусить сам бути вбитий мечем! Отут терпеливість та віра святих!
REV|13|11|І бачив я іншу звірину, що виходила з землі. І вона мала два роги, подібні ягнячим, та говорила, як змій.
REV|13|12|І вона виконувала всю владу першої звірини перед нею, і робила, щоб земля та ті, хто живе на ній, вклонилися першій звірині, що в неї вздоровлена була її рана смертельна.
REV|13|13|І чинить вона великі ознаки, так що й огонь зводить з неба додолу перед людьми.
REV|13|14|І зводить вона мешканців землі через ознаки, що їх дано їй чинити перед звіриною, намовляючи мешканців землі зробити образа звірини, що має рану від меча, та живе.
REV|13|15|І дано їй вкласти духа образові звірини, щоб заговорив образ звірини, і зробити, щоб усі, хто не поклониться образові звірини, побиті були.
REV|13|16|І зробить вона, щоб усім малим і великим, багатим і вбогим, вільним і рабам було дано знамено на їхню правицю або на їхні чола,
REV|13|17|щоб ніхто не міг ані купити, ані продати, якщо він не має знамена ймення звірини, або числа ймення його...
REV|13|18|Тут мудрість! Хто має розум, нехай порахує число звірини, бо воно число людське. А число її шістсот шістдесят шість.
REV|14|1|І я глянув, і ось Агнець стоїть на Сіонській горі, а з Ним сто сорок чотири тисячі, що мають Ім'я Його й Ім'я Отця Його, написане на своїх чолах.
REV|14|2|І почув я голос із неба, немов шум великої води, і немов гук міцного грому. І почув я голос гуслярів, що грали на гуслах своїх,
REV|14|3|і співали, як пісню нову перед престолом і перед чотирьома тваринами й старцями. І ніхто не міг навчитися пісні, окрім цих ста сорока чотирьох тисяч, викуплених від землі.
REV|14|4|Це ті, хто не осквернився з жінками, бо чисті вони. Вони йдуть за Агнцем, куди Він іде. Вони викуплені від людей, первістки Богові й Агнцеві,
REV|14|5|не знайшлося бо підступу в їхніх устах, бо вони непорочні!
REV|14|6|І побачив я іншого Ангола, що летів серед неба, і мав благовістити вічну Євангелію мешканцям землі, і кожному людові, і племені, і язику, і народові.
REV|14|7|І він говорив гучним голосом: Побійтеся Бога та славу віддайте Йому, бо настала година суду Його, і вклоніться Тому, Хто створив небо, і землю, і море, і водні джерела!
REV|14|8|А інший, другий Ангол летів слідом і казав: Упав, упав Вавилон, город великий, бо лютим вином розпусти своєї він напоїв усі народи!
REV|14|9|А інший, третій Ангол летів услід за ним, гучним голосом кажучи: Коли хто вклоняється звірині та образу її, і приймає знамено на чолі своїм чи на руці своїй,
REV|14|10|то той питиме з вина Божого гніву, вина незмішаного в чаші гніву Його, і буде мучений в огні й сірці перед Анголами святими та перед Агнцем.
REV|14|11|А дим їхніх мук підійматиметься вічні віки. І не мають спокою день і ніч усі ті, хто вклоняється звірині та образу її, і приймає знамено ймення його.
REV|14|12|Тут терпеливість святих, що додержують заповіді Божі та Ісусову віру!
REV|14|13|І почув я голос із неба, що до мене казав: Напиши: Блаженні ті мертві, хто з цього часу вмирає в Господі! Так, каже Дух, вони від праць своїх заспокояться, бо їхні діла йдуть за ними слідом.
REV|14|14|І я глянув, і ото біла хмара, а на хмарі сидить подібний до Людського Сина. Він мав на своїй голові золотого вінця, а в руці його гострий серп.
REV|14|15|І інший Ангол вийшов із храму, і гучним голосом кликнув до того, хто на хмарі сидів: Пошли серпа свого й жни, бо настала година пожати, дозріло бо жниво землі!
REV|14|16|І той, хто на хмарі сидів, скинув додолу серпа свого, і земля була вижата.
REV|14|17|І інший Ангол вийшов із храму, що на небі, і він мав гострого серпа.
REV|14|18|І інший Ангол, що мав владу над огнем, вийшов від жертівника. І він гучним голосом кликнув до того, що мав гострого серпа, говорячи: Пошли свого гострого серпа, і позбирай грона земної виноградини, бо грона її вже доспіли.
REV|14|19|І Ангол кинув додолу серпа свого, і зібрав виноград на землі, і вкинув в велике чавило Божого гніву.
REV|14|20|І потовчене було чавило за містом, і потекла кров із чавила аж до кінських вуздечок, на тисячу шістсот стадій...
REV|15|1|І бачив я інше знамено на небі, велике та дивне, сім Анголів, що сім кар вони мали, бо ними кінчався гнів Божий.
REV|15|2|І я бачив щось, ніби як море скляне, з огнем перемішане. А ті, що перемогли звірину та образа його, і знамено його, і число його ймення, стояли на морі склянім, та мали гусла Божі.
REV|15|3|І співали вони пісню Мойсея, раба Божого, і пісню Агнця, говорячи: Великі та дивні діла Твої, о Господи, Боже Вседержителю! Справедливі й правдиві дороги Твої, о Царю святих!
REV|15|4|Хто Тебе, Господи, не побоїться, та Ймення Твого не прославить? Бо один Ти святий, бо народи всі прийдуть та вклоняться перед Тобою, бо з'явилися суди Твої!
REV|15|5|А по цьому я глянув, і ось відчинився храм скинії свідчення в небі,
REV|15|6|і сім Анголів вийшли з храму, і сім кар вони мали. Вони були вдягнені в шати льняні, чисті й ясні, і підперезані довкола грудей золотими поясами.
REV|15|7|І одна з чотирьох тих тварин дала сімом Анголам сім чаш золотих, наповнених гніву Бога, що живе повік віку.
REV|15|8|І храм переповнився димом від Божої слави, і від сили Його. Та до храму ніхто не спромігся ввійти, аж поки не скінчилися ті сім кар сімох Анголів.
REV|16|1|І я почув гучний голос із храму, що казав до семи Анголів: Ідіть, і вилийте на землю сім чаш гніву Божого!
REV|16|2|І пішов перший Ангол, і вилив на землю чашу свою. І шкідливі та люті болячки обсіли людей, хто мав знамено звірини й вклонявсь її образу.
REV|16|3|А другий Ангол вилив свою чашу до моря. І сталася кров, немов у мерця, і кожна істота жива вмерла в морі.
REV|16|4|Третій же Ангол вилив чашу свою на річки та на водні джерела, і сталася кров.
REV|16|5|І почув я Ангола вод, який говорив: Ти праведний, що Ти є й що Ти був, і святий, що Ти це присудив!
REV|16|6|Бо вони пролили кров святих та пророків, і Ти дав їм напитися крови. Вони варті того!
REV|16|7|І я чув, як жертівник говорив: Так, Господи, Боже Вседержителю! Правдиві й справедливі суди Твої!
REV|16|8|А Ангол четвертий вилив свою чашу на сонце. І дано йому палити людей огнем.
REV|16|9|І спека велика палила людей, і зневажали вони Ім'я Бога, що має владу над карами тими, і вони не покаялися, щоб славу віддати Йому.
REV|16|10|А п'ятий Ангол вилив чашу свою на престола звірини. І затьмилося царство її, і люди від болю кусали свої язики,
REV|16|11|і Бога Небесного вони зневажали від болю свого й від своїх болячок, та в учинках своїх не покаялись!
REV|16|12|Шостий же Ангол вилив чашу свою на річку велику Ефрат, і вода її висохла, щоб приготовити дорогу царям, які від схід сонця.
REV|16|13|І я бачив, що виходили з уст змія, і з уст звірини, і з уст неправдивого пророка три духи нечисті, як жаби,
REV|16|14|це духи демонські, що чинять ознаки. Вони виходять до царів усього всесвіту, щоб зібрати їх на війну того великого дня Вседержителя Бога.
REV|16|15|Ось іду, немов злодій! Блаженний, хто чуйний, і одежу свою береже, щоб нагим не ходити, і щоб не бачили ганьби його!
REV|16|16|І зібрав їх на місце, яке по-єврейському зветься Армагеддон.
REV|16|17|Сьомий же Ангол вилив чашу свою на повітря. І голос гучний залунав від небесного храму з престолу, говорячи: Сталося!
REV|16|18|І сталися блискавки й гуркіт та громи, і сталось велике трясіння землі, якого не було, відколи людина живе на землі... Великий такий землетрус, такий міцний!
REV|16|19|І місто велике розпалося на три частині, і попадали людські міста... І великий Вавилон був згаданий перед Богом, щоб дати йому чашу вина Його лютого гніву...
REV|16|20|І зник кожен острів, і не знайдено гір!...
REV|16|21|І великий град, як важкі тягарі, падав із неба на людей. І люди зневажали Бога за покарання градом, бо кара Його була дуже велика!...
REV|17|1|І прийшов один із семи Анголів, що мають сім чаш, і говорив зо мною, кажучи: Підійди, я покажу тобі засудження великої розпусниці, що сидить над багатьма водами.
REV|17|2|З нею розпусту чинили земні царі, і вином розпусти її впивались мешканці землі.
REV|17|3|І в дусі повів він мене на пустиню. І побачив я жінку, що сиділа на червоній звірині, переповненій іменами богозневажними, яка мала сім голів і десять рогів.
REV|17|4|А жінка була одягнена в порфіру й кармазин, і приоздоблена золотом і дорогоцінним камінням та перлами. У руці своїй мала вона золоту чашу, повну гидоти та нечести розпусти її.
REV|17|5|А на чолі її було написане ім'я, таємниця: Великий Вавилон, мати розпусти й гидоти землі.
REV|17|6|І бачив я жінку, п'яну від крови святих і від крови мучеників Ісусових, і, бачивши її, дивувався я дивом великим.
REV|17|7|А Ангол промовив до мене: Чого ти дивуєшся? Я скажу тобі таємницю жінки й звірини, яка носить її, яка має сім голів і десять рогів.
REV|17|8|Звірина, яку бачив я, була і нема, і має вийти з безодні і піде вона на погибіль. А мешканці землі, що їхні імена не записані в книгу життя від закладин світу, дивуватися будуть, як побачать, що звірина була і нема, і з'явиться.
REV|17|9|Тут розум, що має він мудрість. Сім голів це сім гір, що на них сидить жінка. І сім царів,
REV|17|10|п'ять їх упало, один є, другий іще не прийшов, а як прийде, то мусить він трохи пробути.
REV|17|11|І звірина, що була і нема, і вона сама восьма й з сімох, і йде на погибіль.
REV|17|12|А десять тих рогів, що бачив ти їх, то десять царів, що ще не прийняли царства, але приймуть владу царську із звіриною на одну годину.
REV|17|13|Вони мають одну думку, а силу та владу свою віддадуть звірині.
REV|17|14|Вони воюватимуть проти Агнця та Агнець переможе їх, бо Він Господь над панами та Цар над царями. А ті, хто з Ним, покликані, і вибрані, і вірні.
REV|17|15|І говорить до мене: Води, що бачив ти їх, де сидить та розпусниця, то народи та люди, і племена та язики.
REV|17|16|А десять рогів, що ти бачив їх, та звірина, вони зненавидять розпусницю, спустошать її й обнажать, і з'їдять її тіло, і огнем її спалять.
REV|17|17|Бо Бог дав їм до серця, щоб волю чинили Його, маючи одну думку, і щоб царство своє віддали звірині, аж поки не виповняться слова Божі.
REV|17|18|А жінка, яку ти бачив, то місто велике, що панує над царями земними.
REV|18|1|Після цього побачив я іншого Ангола, що сходив із неба, і що владу велику він мав. І земля освітилась від слави його.
REV|18|2|І він гучним голосом кликнув, говорячи: Упав, упав великий Вавилон! Став він оселею демонів, і сховищем усякому духові нечистому, і сховищем усіх птахів нечистих та ненавидних,
REV|18|3|бо лютим вином розпусти своєї він напоїв всі народи! І земні царі з ним розпусту чинили, а земні купці збагатіли від сили розкоші його!
REV|18|4|І почув я інший голос із неба, який говорив: Вийдіть із нього, люди мої, щоб не сталися ви спільниками гріхів його, і щоб не потрапили в карання його.
REV|18|5|Гріхи бо його досягли аж до неба, і Бог ізгадав про неправди його.
REV|18|6|Відплатіть ви йому, як і він вам платив, і вдвоє подвойте йому за вчинки його! Удвоє налийте до чаші, що нею він вам наливав!
REV|18|7|Скільки він славив себе та розкошував, стільки муки та смутку завдайте йому! Бо в серці своєму говорить: Сиджу, як цариця, і я не вдова, і бачити смутку не буду!
REV|18|8|Через це одного дня прийдуть кари його, смерть, і плач, і голод, і спалений буде огнем, бо міцний Господь, Бог, що судить його!
REV|18|9|І будуть плакати та голосити за ним царі земні, що з ним розпусту чинили та розкошували, коли побачать дим пожежі його.
REV|18|10|Вони через страх його мук стоятимуть здалека та говоритимуть: Горе, горе, о місто велике, Вавилоне, місто могутнє, бо суд твій прийшов однієї години!
REV|18|11|І земні купці будуть плакати та голосити за ним, бо ніхто не купує вже їхнього вантажу,
REV|18|12|вантажу золота, і срібла, і каміння дорогоцінного, і перел, і віссону, і порфіри, і шовку, і кармазину, і всякого дерева запашного, і всякого посуду з слонової кости, і всякого посуду з дорогоцінного дерева, і мідяного, і залізного, і мармурового,
REV|18|13|і кориці, і шафрану, і пахощів, і мирри, і ливану, і вина, і оливи, і тонкої муки, і пшениці, і товару, і вівців, і коней, і возів, і рабів, і душ людських.
REV|18|14|І плоди пожадливости душі твоєї відійшли від тебе, і все сите та світле пропало для тебе, і вже їх ти не знайдеш!
REV|18|15|Купці цими речами, що вони збагатилися з нього, від страху мук його стануть здалека, і будуть плакати та голосити,
REV|18|16|і казати: Горе, горе, місто велике, зодягнене в віссон і порфіру та в кармазин, і прикрашене золотом і дорогоцінним камінням та перлами,
REV|18|17|бо за одну годину згинуло таке велике багатство... І кожен стерник, і кожен, хто пливає на кораблях, і моряки, і всі, хто працює на морі, стали здалека,
REV|18|18|і, бачивши дим від пожежі його, кричали й казали: Котре до великого міста подібне?
REV|18|19|І вони посипали порохом голови свої, і закричали, плачучи та голосячи, і кажучи: Горе, горе, місто велике, що в ньому з його дорогоцінностей збагатилися всі, хто має кораблі на морі, бо за одну годину воно спорожніло!
REV|18|20|Радій з цього, небо, і святі апостоли та пророки, бо Бог виконав суд ваш над ним!
REV|18|21|І один сильний Ангол узяв великого каменя, як жорно, і кинув до моря, говорячи: З таким розгоном буде кинений Вавилон, місто велике, і вже він не знайдеться!
REV|18|22|І голос гуслярів, і співаків, і сопільників, і сурмачів уже не буде чутий в тобі! І вже не знайдеться в тобі жадного мистця й ніякого мистецтва, і шум жорен уже не буде чутий в тобі!
REV|18|23|І світло свічника вже не буде світити в тобі, і голос молодого й молодої вже не буде чутий в тобі. Бо купці твої були земні вельможі, бо твоїм ворожбитством були зведені всі народи!
REV|18|24|Бо в нім знайдена кров пророків, і святих, і побитих усіх на землі...
REV|19|1|По цьому почув я наче гучний голос великого натовпу в небі, який говорив: Алілуя! Спасіння, і слава, і сила Господеві нашому,
REV|19|2|правдиві бо та справедливі суди Його, бо Він засудив ту велику розпусницю, що землю зіпсула своєю розпустою, і помстив за кров Своїх рабів з її рук!
REV|19|3|І вдруге сказали вони: Алілуя! І з неї дим виступає на вічні віки!
REV|19|4|І попадали двадцять чотири старці й чотири тварині, і поклонилися Богові, що сидить на престолі, говорячи: Амінь, алілуя!
REV|19|5|А від престолу вийшов голос, що кликав: Хваліть Бога нашого, усі раби Його, і всі, хто боїться Його, і малі, і великі!
REV|19|6|І почув я ніби голос великого натовпу, і наче шум великої води, і мов голос громів гучних, що вигукували: Алілуя, бо запанував Господь, наш Бог Вседержитель!
REV|19|7|Радіймо та тішмося, і даймо славу Йому, бо весілля Агнця настало, і жона Його себе приготувала!
REV|19|8|І їй дано було зодягнутися в чистий та світлий вісон, бо віссон то праведність святих.
REV|19|9|І сказав він мені: Напиши: Блаженні покликані на весільну вечерю Агнця! І сказав він мені: Це правдиві Божі слова!
REV|19|10|І я впав до його ніг, щоб вклонитись йому. І він каже мені: Таж ні! Я співслуга твій та братів твоїх, хто має засвідчення Ісусове, Богові вклонися! Бо засвідчення Ісусове, то дух пророцтва.
REV|19|11|І побачив я небо відкрите. І ось білий кінь, а Той, Хто на ньому сидів, зветься Вірний і Правдивий, і Він справедливо судить і воює.
REV|19|12|Очі Його немов полум'я огняне, а на голові Його багато вінців. Він ім'я мав написане, якого не знає ніхто, тільки Він Сам.
REV|19|13|І зодягнений був Він у шату, покрашену кров'ю. А Йому на ім'я: Слово Боже.
REV|19|14|А війська небесні, зодягнені в білий та чистий віссон, їхали вслід за Ним на білих конях.
REV|19|15|А з Його уст виходив гострий меч, щоб ним бити народи. І Він пастиме їх залізним жезлом, і Він буде топтати чавило вина лютого гніву Бога Вседержителя!
REV|19|16|І Він має на шаті й на стегнах Своїх написане ймення: Цар над царями, і Господь над панами.
REV|19|17|І бачив я одного Ангола, що на сонці стояв. І він гучним голосом кликнув, кажучи до всіх птахів, що серед неба літали: Ходіть, і зберіться на велику Божу вечерю,
REV|19|18|щоб ви їли тіла царів, і тіла тисячників, і тіла сильних, і тіла коней і тих, хто сидить на них, і тіла всіх вільних і рабів, і малих, і великих...
REV|19|19|І я побачив звірину, і земних царів, і війська їхні, зібрані, щоб учинити війну з Тим, Хто сидить на коні, та з військом Його.
REV|19|20|І схоплена була звірина, а з нею неправдивий пророк, що ознаки чинив перед нею, що ними звів тих, хто знамено звірини прийняв і поклонився був образові її. Обоє вони були вкинені живими до огняного озера, що сіркою горіло...
REV|19|21|А решта побита була мечем Того, Хто сидів на коні, що виходив із уст Його. І все птаство наїлося їхніми трупами...
REV|20|1|І бачив я Ангола, що сходив із неба, що мав ключа від безодні, і кайдани великі в руці своїй.
REV|20|2|І схопив він змія, вужа стародавнього, що диявол він і сатана, і зв'язав його на тисячу років,
REV|20|3|та й кинув його до безодні, і замкнув його, і печатку над ним поклав, щоб народи не зводив уже, аж поки не скінчиться тисяча років. А по цьому він розв'язаний буде на короткий час.
REV|20|4|І бачив я престоли та тих, хто сидів на них, і суд їм був даний, і душі стятих за свідчення про Ісуса й за Слово Боже, які не вклонились звірині, ані образові її, і не прийняли знамена на чола свої та на руку свою. І вони ожили, і царювали з Христом тисячу років.
REV|20|5|А інші померлі не ожили, аж поки не скінчиться тисяча років. Це перше воскресіння.
REV|20|6|Блаженний і святий, хто має частку в першому воскресінні! Над ними друга смерть не матиме влади, але вони будуть священиками Бога й Христа, і царюватимуть з Ним тисячу років.
REV|20|7|Коли ж скінчиться тисяча років, сатана буде випущений із в'язниці своєї.
REV|20|8|І вийде він зводити народи, що вони на чотирьох краях землі, Ґоґа й Маґоґа, щоб зібрати їх до бою, а число їхнє як морський пісок.
REV|20|9|І вийшли вони на ширину землі, і оточили табір святих та улюблене місто. І зійшов огонь з неба, і пожер їх.
REV|20|10|А диявол, що зводив їх, був укинений в озеро огняне та сірчане, де звірина й пророк неправдивий. І мучені будуть вони день і ніч на вічні віки.
REV|20|11|І я бачив престола великого білого, і Того, Хто на ньому сидів, що від лиця Його втекла земля й небо, і місця для них не знайшлося.
REV|20|12|І бачив я мертвих малих і великих, що стояли перед Богом. І розгорнулися книги, і розгорнулась інша книга, то книга життя. І суджено мертвих, як написано в книгах, за вчинками їхніми.
REV|20|13|І дало море мертвих, що в ньому, і смерть і ад дали мертвих, що в них, і суджено їх згідно з їхніми вчинками.
REV|20|14|Смерть же та ад були вкинені в озеро огняне. Це друга смерть, озеро огняне.
REV|20|15|А хто не знайшовся написаний в книзі життя, той укинений буде в озеро огняне...
REV|21|1|І бачив я небо нове й нову землю, перше бо небо та перша земля проминули, і моря вже не було.
REV|21|2|І я, Іван, бачив місто святе, Новий Єрусалим, що сходив із неба від Бога, що був приготований, як невіста, прикрашена для чоловіка свого.
REV|21|3|І почув я гучний голос із престолу, який кликав: Оце оселя Бога з людьми, і Він житиме з ними! Вони будуть народом Його, і Сам Бог буде з ними,
REV|21|4|і Бог кожну сльозу з очей їхніх зітре, і не буде вже смерти. Ані смутку, ані крику, ані болю вже не буде, бо перше минулося!
REV|21|5|І сказав Той, Хто сидить на престолі: Ось нове все творю! І говорить: Напиши, що слова ці правдиві та вірні!
REV|21|6|І сказав Він мені: Сталося! Я Альфа й Омега, Початок і Кінець. Хто прагне, тому дармо Я дам від джерела живої води.
REV|21|7|Переможець наслідить усе, і Я буду Богом для нього, а він Мені буде за сина!
REV|21|8|А лякливим, і невірним, і мерзким, і душогубам, і розпусникам, і чарівникам, і ідолянам, і всім неправдомовцям, їхня частина в озері, що горить огнем та сіркою, а це друга смерть!
REV|21|9|І прийшов до мене один із семи Анголів, що мають сім чаш, наповнених сімома останніми карами, та й промовив до мене, говорячи: Ходи, покажу я тобі невісту, жону Агнця.
REV|21|10|І заніс мене духом на гору велику й високу, і місто велике мені показав, святий Єрусалим, що сходив із неба від Бога.
REV|21|11|Славу Божу він має. А світлість його подібна до каменя дорогоцінного, як каменя ясписа, що блищить, як кришталь.
REV|21|12|Мур воно мало великий і високий, мало дванадцять брам, а на брамах дванадцять Анголів та ймення написані, а вони імення дванадцятьох племен синів Ізраїля.
REV|21|13|Від сходу три брамі, і від півночі три брамі, і від півдня три брамі, і від заходу три брамі.
REV|21|14|І міський мур мав дванадцять підвалин, а на них дванадцять імен дванадцяти апостолів Агнця.
REV|21|15|А той, хто зо мною говорив, мав міру, золоту тростину, щоб зміряти місто, і брами його і його мур.
REV|21|16|А місто чотирикутнє, а довжина його така, як і ширина. І він зміряв місто тростиною на дванадцять тисяч стадій; довжина, і ширина, і вишина його рівні.
REV|21|17|І зміряв він мура його на сто сорок чотири лікті міри людської, яка й міра Ангола.
REV|21|18|Його мур був збудований з яспису, а місто було щире золото, подібне до чистого скла.
REV|21|19|Підвалини муру міського прикрашені були всяким дорогоцінним камінням. Перша підвалина яспис, друга сапфір, третя халкидон, четверта смарагд,
REV|21|20|п'ята сардонікс, шоста сардій, сьома хризоліт, восьма берил, дев'ята топаз, десята хрисопрас, одинадцята якинт, дванадцята аметист.
REV|21|21|А дванадцять брам то дванадцять перлин, і кожна брама зокрема була з однієї перлини. А вулиці міста щире золото, прозорі, як скло.
REV|21|22|А храму не бачив я в ньому, бо Господь, Бог Вседержитель то йому храм і Агнець.
REV|21|23|І місто не має потреби ні в сонці, ні в місяці, щоб у ньому світили, слава бо Божа його освітила, а світильник для нього Агнець.
REV|21|24|І народи ходитимуть у світлі його, а земські царі принесуть свою славу до нього.
REV|21|25|А брами його зачинятись не будуть удень, бо там ночі не буде.
REV|21|26|І принесуть до нього славу й честь народів.
REV|21|27|І не ввійде до нього ніщо нечисте, ані той, хто чинить гидоту й неправду, але тільки ті, хто записаний у книзі життя Агнця.
REV|22|1|І показав він мені чисту ріку живої води, ясну, мов кришталь, що випливала з престолу Бога й Агнця.
REV|22|2|Посеред його вулиці, і по цей бік і по той бік ріки дерево життя, що родить дванадцять раз плоди, кожного місяця приносячи плід свій. А листя дерев на вздоровлення народів.
REV|22|3|І жадного прокляття більше не буде. І буде в ньому Престол Бога та Агнця, а раби Його будуть служити Йому,
REV|22|4|і побачать лице Його, а Ймення Його на їхніх чолах.
REV|22|5|А ночі вже більше не буде, і не буде потреби в світлі світильника, ані в світлі сонця, бо освітлює їх Господь, Бог, а вони царюватимуть вічні віки.
REV|22|6|І сказав він до мене: Це вірні й правдиві слова, а Господь, Бог духів пророчих, послав Свого Ангола, щоб він показав своїм рабам, що незабаром статися мусить.
REV|22|7|Ото, незабаром приходжу. Блаженний, хто зберігає пророчі слова цієї книги!
REV|22|8|І я, Іван, чув і бачив оце. А коли я почув та побачив, я впав до ніг Ангола, що мені це показував, щоб вклонитись йому.
REV|22|9|І сказав він до мене: Таж ні! Бо я співслуга твій і братів твоїх пророків, і тих, хто зберігає слова цієї книги. Богові вклонися!
REV|22|10|І сказав він до мене: Не запечатуй слів пророцтва цієї книги. Час бо близький!
REV|22|11|Неправедний нехай чинить неправду ще, і поганий нехай ще опоганюється. А праведний нехай ще чинить правду, а святий нехай ще освячується!
REV|22|12|Ото, незабаром приходжу, і зо Мною заплата Моя, щоб кожному віддати згідно з ділами його.
REV|22|13|Я Альфа й Омега, Перший і Останній, Початок і Кінець.
REV|22|14|Блаженні, хто випере шати свої, щоб мати право на дерево життя, і ввійти брамами в місто!
REV|22|15|А поза ним будуть пси, і чарівники, і розпусники, і душогуби, і ідоляни, і кожен, хто любить та чинить неправду.
REV|22|16|Я, Ісус, послав Свого Ангола, щоб засвідчити вам це у Церквах. Я корінь і рід Давидів, зоря ясна і досвітня!
REV|22|17|А Дух і невіста говорять: Прийди! А хто чує, хай каже: Прийди! І хто прагне, хай прийде, і хто хоче, хай воду життя бере дармо!
REV|22|18|Свідкую я кожному, хто чує слова пророцтва цієї книги: Коли хто до цього додасть що, то накладе на нього Бог кари, що написані в книзі оцій.
REV|22|19|А коли хто що відійме від слів книги пророцтва цього, то відійме Бог частку його від дерева життя, і від міста святого, що написане в книзі оцій.
REV|22|20|Той, Хто свідкує, говорить оце: Так, незабаром прийду! Амінь. Прийди, Господи Ісусе!
REV|22|21|Благодать Господа нашого Ісуса Христа зо всіма вами! Амінь.
