JAS|1|1|Iacobus Dei et Domini nostri Iesu Christi servus duodecim tribubus quae sunt in dispersione salutem
JAS|1|2|omne gaudium existimate fratres mei cum in temptationibus variis incideritis
JAS|1|3|scientes quod probatio fidei vestrae patientiam operatur
JAS|1|4|patientia autem opus perfectum habeat ut sitis perfecti et integri in nullo deficientes
JAS|1|5|si quis autem vestrum indiget sapientiam postulet a Deo qui dat omnibus affluenter et non inproperat et dabitur ei
JAS|1|6|postulet autem in fide nihil haesitans qui enim haesitat similis est fluctui maris qui a vento movetur et circumfertur
JAS|1|7|non ergo aestimet homo ille quod accipiat aliquid a Domino
JAS|1|8|vir duplex animo inconstans in omnibus viis suis
JAS|1|9|glorietur autem frater humilis in exaltatione sua
JAS|1|10|dives autem in humilitate sua quoniam sicut flos faeni transibit
JAS|1|11|exortus est enim sol cum ardore et arefecit faenum et flos eius decidit et decor vultus eius deperiit ita et dives in itineribus suis marcescet
JAS|1|12|beatus vir qui suffert temptationem quia cum probatus fuerit accipiet coronam vitae quam repromisit Deus diligentibus se
JAS|1|13|nemo cum temptatur dicat quoniam a Deo temptor Deus enim intemptator malorum est ipse autem neminem temptat
JAS|1|14|unusquisque vero temptatur a concupiscentia sua abstractus et inlectus
JAS|1|15|dein concupiscentia cum conceperit parit peccatum peccatum vero cum consummatum fuerit generat mortem
JAS|1|16|nolite itaque errare fratres mei dilectissimi
JAS|1|17|omne datum optimum et omne donum perfectum desursum est descendens a Patre luminum apud quem non est transmutatio nec vicissitudinis obumbratio
JAS|1|18|voluntarie genuit nos verbo veritatis ut simus initium aliquod creaturae eius
JAS|1|19|scitis fratres mei dilecti sit autem omnis homo velox ad audiendum tardus autem ad loquendum et tardus ad iram
JAS|1|20|ira enim viri iustitiam Dei non operatur
JAS|1|21|propter quod abicientes omnem inmunditiam et abundantiam malitiae in mansuetudine suscipite insitum verbum quod potest salvare animas vestras
JAS|1|22|estote autem factores verbi et non auditores tantum fallentes vosmet ipsos
JAS|1|23|quia si quis auditor est verbi et non factor hic conparabitur viro consideranti vultum nativitatis suae in speculo
JAS|1|24|consideravit enim se et abiit et statim oblitus est qualis fuerit
JAS|1|25|qui autem perspexerit in lege perfecta libertatis et permanserit non auditor obliviosus factus sed factor operis hic beatus in facto suo erit
JAS|1|26|si quis autem putat se religiosum esse non refrenans linguam suam sed seducens cor suum huius vana est religio
JAS|1|27|religio munda et inmaculata apud Deum et Patrem haec est visitare pupillos et viduas in tribulatione eorum inmaculatum se custodire ab hoc saeculo
JAS|2|1|fratres mei nolite in personarum acceptione habere fidem Domini nostri Iesu Christi gloriae
JAS|2|2|etenim si introierit in conventu vestro vir aureum anulum habens in veste candida introierit autem et pauper in sordido habitu
JAS|2|3|et intendatis in eum qui indutus est veste praeclara et dixeritis tu sede hic bene pauperi autem dicatis tu sta illic aut sede sub scabillo pedum meorum
JAS|2|4|nonne iudicatis apud vosmet ipsos et facti estis iudices cogitationum iniquarum
JAS|2|5|audite fratres mei dilectissimi nonne Deus elegit pauperes in hoc mundo divites in fide et heredes regni quod repromisit Deus diligentibus se
JAS|2|6|vos autem exhonorastis pauperem nonne divites per potentiam opprimunt vos et ipsi trahunt vos ad iudicia
JAS|2|7|nonne ipsi blasphemant bonum nomen quod invocatum est super vos
JAS|2|8|si tamen legem perficitis regalem secundum scripturas diliges proximum tuum sicut te ipsum bene facitis
JAS|2|9|si autem personas accipitis peccatum operamini redarguti a lege quasi transgressores
JAS|2|10|quicumque autem totam legem servaverit offendat autem in uno factus est omnium reus
JAS|2|11|qui enim dixit non moechaberis dixit et non occides quod si non moechaberis occides autem factus es transgressor legis
JAS|2|12|sic loquimini et sic facite sicut per legem libertatis incipientes iudicari
JAS|2|13|iudicium enim sine misericordia illi qui non fecit misericordiam superexultat autem misericordia iudicio
JAS|2|14|quid proderit fratres mei si fidem quis dicat se habere opera autem non habeat numquid poterit fides salvare eum
JAS|2|15|si autem frater aut soror nudi sunt et indigent victu cotidiano
JAS|2|16|dicat autem aliquis de vobis illis ite in pace calefacimini et saturamini non dederitis autem eis quae necessaria sunt corporis quid proderit
JAS|2|17|sic et fides si non habeat opera mortua est in semet ipsam
JAS|2|18|sed dicet quis tu fidem habes et ego opera habeo ostende mihi fidem tuam sine operibus et ego ostendam tibi ex operibus fidem meam
JAS|2|19|tu credis quoniam unus est Deus bene facis et daemones credunt et contremescunt
JAS|2|20|vis autem scire o homo inanis quoniam fides sine operibus otiosa est
JAS|2|21|Abraham pater noster nonne ex operibus iustificatus est offerens Isaac filium suum super altare
JAS|2|22|vides quoniam fides cooperabatur operibus illius et ex operibus fides consummata est
JAS|2|23|et suppleta est scriptura dicens credidit Abraham Deo et reputatum est illi ad iustitiam et amicus Dei appellatus est
JAS|2|24|videtis quoniam ex operibus iustificatur homo et non ex fide tantum
JAS|2|25|similiter autem et Raab meretrix nonne ex operibus iustificata est suscipiens nuntios et alia via eiciens
JAS|2|26|sicut enim corpus sine spiritu emortuum est ita et fides sine operibus mortua est
JAS|3|1|nolite plures magistri fieri fratres mei scientes quoniam maius iudicium sumitis
JAS|3|2|in multis enim offendimus omnes si quis in verbo non offendit hic perfectus est vir potens etiam freno circumducere totum corpus
JAS|3|3|si autem equorum frenos in ora mittimus ad consentiendum nobis et omne corpus illorum circumferimus
JAS|3|4|ecce et naves cum magnae sint et a ventis validis minentur circumferuntur a modico gubernaculo ubi impetus dirigentis voluerit
JAS|3|5|ita et lingua modicum quidem membrum est et magna exultat ecce quantus ignis quam magnam silvam incendit
JAS|3|6|et lingua ignis est universitas iniquitatis lingua constituitur in membris nostris quae maculat totum corpus et inflammat rotam nativitatis nostrae inflammata a gehenna
JAS|3|7|omnis enim natura bestiarum et volucrum et serpentium etiam ceterorum domantur et domita sunt a natura humana
JAS|3|8|linguam autem nullus hominum domare potest inquietum malum plena veneno mortifero
JAS|3|9|in ipsa benedicimus Dominum et Patrem et in ipsa maledicimus homines qui ad similitudinem Dei facti sunt
JAS|3|10|ex ipso ore procedit benedictio et maledictio non oportet fratres mei haec ita fieri
JAS|3|11|numquid fons de eodem foramine emanat dulcem et amaram aquam
JAS|3|12|numquid potest fratres mei ficus olivas facere aut vitis ficus sic neque salsa dulcem potest facere aquam
JAS|3|13|quis sapiens et disciplinatus inter vos ostendat ex bona conversatione operationem suam in mansuetudine sapientiae
JAS|3|14|quod si zelum amarum habetis et contentiones in cordibus vestris nolite gloriari et mendaces esse adversus veritatem
JAS|3|15|non est ista sapientia desursum descendens sed terrena animalis diabolica
JAS|3|16|ubi enim zelus et contentio ibi inconstantia et omne opus pravum
JAS|3|17|quae autem desursum est sapientia primum quidem pudica est deinde pacifica modesta suadibilis plena misericordia et fructibus bonis non iudicans sine simulatione
JAS|3|18|fructus autem iustitiae in pace seminatur facientibus pacem
JAS|4|1|unde bella et lites in vobis nonne hinc ex concupiscentiis vestris quae militant in membris vestris
JAS|4|2|concupiscitis et non habetis occiditis et zelatis et non potestis adipisci litigatis et belligeratis non habetis propter quod non postulatis
JAS|4|3|petitis et non accipitis eo quod male petatis ut in concupiscentiis vestris insumatis
JAS|4|4|adulteri nescitis quia amicitia huius mundi inimica est Dei quicumque ergo voluerit amicus esse saeculi huius inimicus Dei constituitur
JAS|4|5|aut putatis quia inaniter scriptura dicat ad invidiam concupiscit Spiritus qui inhabitat in nobis
JAS|4|6|maiorem autem dat gratiam propter quod dicit Deus superbis resistit humilibus autem dat gratiam
JAS|4|7|subditi igitur estote Deo resistite autem diabolo et fugiet a vobis
JAS|4|8|adpropiate Domino et adpropinquabit vobis emundate manus peccatores et purificate corda duplices animo
JAS|4|9|miseri estote et lugete et plorate risus vester in luctum convertatur et gaudium in maerorem
JAS|4|10|humiliamini in conspectu Domini et exaltabit vos
JAS|4|11|nolite detrahere de alterutrum fratres qui detrahit fratri aut qui iudicat fratrem suum detrahit legi et iudicat legem si autem iudicas legem non es factor legis sed iudex
JAS|4|12|unus est legislator et iudex qui potest perdere et liberare tu autem quis es qui iudicas proximum
JAS|4|13|ecce nunc qui dicitis hodie aut crastino ibimus in illam civitatem et faciemus quidem ibi annum et mercabimur et lucrum faciemus
JAS|4|14|qui ignoratis quid erit in crastinum quae enim est vita vestra vapor est ad modicum parens deinceps exterminatur
JAS|4|15|pro eo ut dicatis si Dominus voluerit et vixerimus faciemus hoc aut illud
JAS|4|16|nunc autem exultatis in superbiis vestris omnis exultatio talis maligna est
JAS|4|17|scienti igitur bonum facere et non facienti peccatum est illi
JAS|5|1|age nunc divites plorate ululantes in miseriis quae advenient vobis
JAS|5|2|divitiae vestrae putrefactae sunt et vestimenta vestra a tineis comesta sunt
JAS|5|3|aurum et argentum vestrum eruginavit et erugo eorum in testimonium vobis erit et manducabit carnes vestras sicut ignis thesaurizastis in novissimis diebus
JAS|5|4|ecce merces operariorum qui messuerunt regiones vestras qui fraudatus est a vobis clamat et clamor ipsorum in aures Domini Sabaoth introiit
JAS|5|5|epulati estis super terram et in luxuriis enutristis corda vestra in die occisionis
JAS|5|6|addixistis occidistis iustum non resistit vobis
JAS|5|7|patientes igitur estote fratres usque ad adventum Domini ecce agricola expectat pretiosum fructum terrae patienter ferens donec accipiat temporivum et serotinum
JAS|5|8|patientes estote et vos confirmate corda vestra quoniam adventus Domini adpropinquavit
JAS|5|9|nolite ingemescere fratres in alterutrum ut non iudicemini ecce iudex ante ianuam adsistit
JAS|5|10|exemplum accipite fratres laboris et patientiae prophetas qui locuti sunt in nomine Domini
JAS|5|11|ecce beatificamus qui sustinuerunt sufferentiam Iob audistis et finem Domini vidistis quoniam misericors est Dominus et miserator
JAS|5|12|ante omnia autem fratres mei nolite iurare neque per caelum neque per terram neque aliud quodcumque iuramentum sit autem vestrum est est non non uti non sub iudicio decidatis
JAS|5|13|tristatur aliquis vestrum oret aequo animo est psallat
JAS|5|14|infirmatur quis in vobis inducat presbyteros ecclesiae et orent super eum unguentes eum oleo in nomine Domini
JAS|5|15|et oratio fidei salvabit infirmum et adlevabit eum Dominus et si in peccatis sit dimittentur ei
JAS|5|16|confitemini ergo alterutrum peccata vestra et orate pro invicem ut salvemini multum enim valet deprecatio iusti adsidua
JAS|5|17|Helias homo erat similis nobis passibilis et oratione oravit ut non plueret super terram et non pluit annos tres et menses sex
JAS|5|18|et rursum oravit et caelum dedit pluviam et terra dedit fructum suum
JAS|5|19|fratres mei si quis ex vobis erraverit a veritate et converterit quis eum
JAS|5|20|scire debet quoniam qui converti fecerit peccatorem ab errore viae suae salvabit animam eius a morte et operit multitudinem peccatorum
