MARK|1|1|The beginning of the gospel about Jesus Christ, the Son of God.
MARK|1|2|It is written in Isaiah the prophet: "I will send my messenger ahead of you, who will prepare your way"--
MARK|1|3|"a voice of one calling in the desert, 'Prepare the way for the Lord, make straight paths for him.'"
MARK|1|4|And so John came, baptizing in the desert region and preaching a baptism of repentance for the forgiveness of sins.
MARK|1|5|The whole Judean countryside and all the people of Jerusalem went out to him. Confessing their sins, they were baptized by him in the Jordan River.
MARK|1|6|John wore clothing made of camel's hair, with a leather belt around his waist, and he ate locusts and wild honey.
MARK|1|7|And this was his message: "After me will come one more powerful than I, the thongs of whose sandals I am not worthy to stoop down and untie.
MARK|1|8|I baptize you with water, but he will baptize you with the Holy Spirit."
MARK|1|9|At that time Jesus came from Nazareth in Galilee and was baptized by John in the Jordan.
MARK|1|10|As Jesus was coming up out of the water, he saw heaven being torn open and the Spirit descending on him like a dove.
MARK|1|11|And a voice came from heaven: "You are my Son, whom I love; with you I am well pleased."
MARK|1|12|At once the Spirit sent him out into the desert,
MARK|1|13|and he was in the desert forty days, being tempted by Satan. He was with the wild animals, and angels attended him.
MARK|1|14|After John was put in prison, Jesus went into Galilee, proclaiming the good news of God.
MARK|1|15|"The time has come," he said. "The kingdom of God is near. Repent and believe the good news!"
MARK|1|16|As Jesus walked beside the Sea of Galilee, he saw Simon and his brother Andrew casting a net into the lake, for they were fishermen.
MARK|1|17|"Come, follow me," Jesus said, "and I will make you fishers of men."
MARK|1|18|At once they left their nets and followed him.
MARK|1|19|When he had gone a little farther, he saw James son of Zebedee and his brother John in a boat, preparing their nets.
MARK|1|20|Without delay he called them, and they left their father Zebedee in the boat with the hired men and followed him.
MARK|1|21|They went to Capernaum, and when the Sabbath came, Jesus went into the synagogue and began to teach.
MARK|1|22|The people were amazed at his teaching, because he taught them as one who had authority, not as the teachers of the law.
MARK|1|23|Just then a man in their synagogue who was possessed by an evil spirit cried out,
MARK|1|24|"What do you want with us, Jesus of Nazareth? Have you come to destroy us? I know who you are--the Holy One of God!"
MARK|1|25|"Be quiet!" said Jesus sternly. "Come out of him!"
MARK|1|26|The evil spirit shook the man violently and came out of him with a shriek.
MARK|1|27|The people were all so amazed that they asked each other, "What is this? A new teaching--and with authority! He even gives orders to evil spirits and they obey him."
MARK|1|28|News about him spread quickly over the whole region of Galilee.
MARK|1|29|As soon as they left the synagogue, they went with James and John to the home of Simon and Andrew.
MARK|1|30|Simon's mother-in-law was in bed with a fever, and they told Jesus about her.
MARK|1|31|So he went to her, took her hand and helped her up. The fever left her and she began to wait on them.
MARK|1|32|That evening after sunset the people brought to Jesus all the sick and demon-possessed.
MARK|1|33|The whole town gathered at the door,
MARK|1|34|and Jesus healed many who had various diseases. He also drove out many demons, but he would not let the demons speak because they knew who he was.
MARK|1|35|Very early in the morning, while it was still dark, Jesus got up, left the house and went off to a solitary place, where he prayed.
MARK|1|36|Simon and his companions went to look for him,
MARK|1|37|and when they found him, they exclaimed: "Everyone is looking for you!"
MARK|1|38|Jesus replied, "Let us go somewhere else--to the nearby villages--so I can preach there also. That is why I have come."
MARK|1|39|So he traveled throughout Galilee, preaching in their synagogues and driving out demons.
MARK|1|40|A man with leprosy came to him and begged him on his knees, "If you are willing, you can make me clean."
MARK|1|41|Filled with compassion, Jesus reached out his hand and touched the man. "I am willing," he said. "Be clean!"
MARK|1|42|Immediately the leprosy left him and he was cured.
MARK|1|43|Jesus sent him away at once with a strong warning:
MARK|1|44|"See that you don't tell this to anyone. But go, show yourself to the priest and offer the sacrifices that Moses commanded for your cleansing, as a testimony to them."
MARK|1|45|Instead he went out and began to talk freely, spreading the news. As a result, Jesus could no longer enter a town openly but stayed outside in lonely places. Yet the people still came to him from everywhere.
MARK|2|1|A few days later, when Jesus again entered Capernaum, the people heard that he had come home.
MARK|2|2|So many gathered that there was no room left, not even outside the door, and he preached the word to them.
MARK|2|3|Some men came, bringing to him a paralytic, carried by four of them.
MARK|2|4|Since they could not get him to Jesus because of the crowd, they made an opening in the roof above Jesus and, after digging through it, lowered the mat the paralyzed man was lying on.
MARK|2|5|When Jesus saw their faith, he said to the paralytic, "Son, your sins are forgiven."
MARK|2|6|Now some teachers of the law were sitting there, thinking to themselves,
MARK|2|7|"Why does this fellow talk like that? He's blaspheming! Who can forgive sins but God alone?"
MARK|2|8|Immediately Jesus knew in his spirit that this was what they were thinking in their hearts, and he said to them, "Why are you thinking these things?
MARK|2|9|Which is easier: to say to the paralytic, 'Your sins are forgiven,' or to say, 'Get up, take your mat and walk'?
MARK|2|10|But that you may know that the Son of Man has authority on earth to forgive sins...." He said to the paralytic,
MARK|2|11|"I tell you, get up, take your mat and go home."
MARK|2|12|He got up, took his mat and walked out in full view of them all. This amazed everyone and they praised God, saying, "We have never seen anything like this!"
MARK|2|13|Once again Jesus went out beside the lake. A large crowd came to him, and he began to teach them.
MARK|2|14|As he walked along, he saw Levi son of Alphaeus sitting at the tax collector's booth. "Follow me," Jesus told him, and Levi got up and followed him.
MARK|2|15|While Jesus was having dinner at Levi's house, many tax collectors and "sinners" were eating with him and his disciples, for there were many who followed him.
MARK|2|16|When the teachers of the law who were Pharisees saw him eating with the "sinners" and tax collectors, they asked his disciples: "Why does he eat with tax collectors and 'sinners'?"
MARK|2|17|On hearing this, Jesus said to them, "It is not the healthy who need a doctor, but the sick. I have not come to call the righteous, but sinners."
MARK|2|18|Now John's disciples and the Pharisees were fasting. Some people came and asked Jesus, "How is it that John's disciples and the disciples of the Pharisees are fasting, but yours are not?"
MARK|2|19|Jesus answered, "How can the guests of the bridegroom fast while he is with them? They cannot, so long as they have him with them.
MARK|2|20|But the time will come when the bridegroom will be taken from them, and on that day they will fast.
MARK|2|21|"No one sews a patch of unshrunk cloth on an old garment. If he does, the new piece will pull away from the old, making the tear worse.
MARK|2|22|And no one pours new wine into old wineskins. If he does, the wine will burst the skins, and both the wine and the wineskins will be ruined. No, he pours new wine into new wineskins."
MARK|2|23|One Sabbath Jesus was going through the grainfields, and as his disciples walked along, they began to pick some heads of grain.
MARK|2|24|The Pharisees said to him, "Look, why are they doing what is unlawful on the Sabbath?"
MARK|2|25|He answered, "Have you never read what David did when he and his companions were hungry and in need?
MARK|2|26|In the days of Abiathar the high priest, he entered the house of God and ate the consecrated bread, which is lawful only for priests to eat. And he also gave some to his companions."
MARK|2|27|Then he said to them, "The Sabbath was made for man, not man for the Sabbath.
MARK|2|28|So the Son of Man is Lord even of the Sabbath."
MARK|3|1|Another time he went into the synagogue, and a man with a shriveled hand was there.
MARK|3|2|Some of them were looking for a reason to accuse Jesus, so they watched him closely to see if he would heal him on the Sabbath.
MARK|3|3|Jesus said to the man with the shriveled hand, "Stand up in front of everyone."
MARK|3|4|Then Jesus asked them, "Which is lawful on the Sabbath: to do good or to do evil, to save life or to kill?" But they remained silent.
MARK|3|5|He looked around at them in anger and, deeply distressed at their stubborn hearts, said to the man, "Stretch out your hand." He stretched it out, and his hand was completely restored.
MARK|3|6|Then the Pharisees went out and began to plot with the Herodians how they might kill Jesus.
MARK|3|7|Jesus withdrew with his disciples to the lake, and a large crowd from Galilee followed.
MARK|3|8|When they heard all he was doing, many people came to him from Judea, Jerusalem, Idumea, and the regions across the Jordan and around Tyre and Sidon.
MARK|3|9|Because of the crowd he told his disciples to have a small boat ready for him, to keep the people from crowding him.
MARK|3|10|For he had healed many, so that those with diseases were pushing forward to touch him.
MARK|3|11|Whenever the evil spirits saw him, they fell down before him and cried out, "You are the Son of God."
MARK|3|12|But he gave them strict orders not to tell who he was.
MARK|3|13|Jesus went up on a mountainside and called to him those he wanted, and they came to him.
MARK|3|14|He appointed twelve--designating them apostles--that they might be with him and that he might send them out to preach
MARK|3|15|and to have authority to drive out demons.
MARK|3|16|These are the twelve he appointed: Simon (to whom he gave the name Peter);
MARK|3|17|James son of Zebedee and his brother John (to them he gave the name Boanerges, which means Sons of Thunder);
MARK|3|18|Andrew, Philip, Bartholomew, Matthew, Thomas, James son of Alphaeus, Thaddaeus, Simon the Zealot
MARK|3|19|and Judas Iscariot, who betrayed him.
MARK|3|20|Then Jesus entered a house, and again a crowd gathered, so that he and his disciples were not even able to eat.
MARK|3|21|When his family heard about this, they went to take charge of him, for they said, "He is out of his mind."
MARK|3|22|And the teachers of the law who came down from Jerusalem said, "He is possessed by Beelzebub! By the prince of demons he is driving out demons."
MARK|3|23|So Jesus called them and spoke to them in parables: "How can Satan drive out Satan?
MARK|3|24|If a kingdom is divided against itself, that kingdom cannot stand.
MARK|3|25|If a house is divided against itself, that house cannot stand.
MARK|3|26|And if Satan opposes himself and is divided, he cannot stand; his end has come.
MARK|3|27|In fact, no one can enter a strong man's house and carry off his possessions unless he first ties up the strong man. Then he can rob his house.
MARK|3|28|I tell you the truth, all the sins and blasphemies of men will be forgiven them.
MARK|3|29|But whoever blasphemes against the Holy Spirit will never be forgiven; he is guilty of an eternal sin."
MARK|3|30|He said this because they were saying, "He has an evil spirit."
MARK|3|31|Then Jesus' mother and brothers arrived. Standing outside, they sent someone in to call him.
MARK|3|32|A crowd was sitting around him, and they told him, "Your mother and brothers are outside looking for you."
MARK|3|33|"Who are my mother and my brothers?" he asked.
MARK|3|34|Then he looked at those seated in a circle around him and said, "Here are my mother and my brothers!
MARK|3|35|Whoever does God's will is my brother and sister and mother."
MARK|4|1|Again Jesus began to teach by the lake. The crowd that gathered around him was so large that he got into a boat and sat in it out on the lake, while all the people were along the shore at the water's edge.
MARK|4|2|He taught them many things by parables, and in his teaching said:
MARK|4|3|"Listen! A farmer went out to sow his seed.
MARK|4|4|As he was scattering the seed, some fell along the path, and the birds came and ate it up.
MARK|4|5|Some fell on rocky places, where it did not have much soil. It sprang up quickly, because the soil was shallow.
MARK|4|6|But when the sun came up, the plants were scorched, and they withered because they had no root.
MARK|4|7|Other seed fell among thorns, which grew up and choked the plants, so that they did not bear grain.
MARK|4|8|Still other seed fell on good soil. It came up, grew and produced a crop, multiplying thirty, sixty, or even a hundred times."
MARK|4|9|Then Jesus said, "He who has ears to hear, let him hear."
MARK|4|10|When he was alone, the Twelve and the others around him asked him about the parables.
MARK|4|11|He told them, "The secret of the kingdom of God has been given to you. But to those on the outside everything is said in parables
MARK|4|12|so that, "'they may be ever seeing but never perceiving, and ever hearing but never understanding; otherwise they might turn and be forgiven!'"
MARK|4|13|Then Jesus said to them, "Don't you understand this parable? How then will you understand any parable?
MARK|4|14|The farmer sows the word.
MARK|4|15|Some people are like seed along the path, where the word is sown. As soon as they hear it, Satan comes and takes away the word that was sown in them.
MARK|4|16|Others, like seed sown on rocky places, hear the word and at once receive it with joy.
MARK|4|17|But since they have no root, they last only a short time. When trouble or persecution comes because of the word, they quickly fall away.
MARK|4|18|Still others, like seed sown among thorns, hear the word;
MARK|4|19|but the worries of this life, the deceitfulness of wealth and the desires for other things come in and choke the word, making it unfruitful.
MARK|4|20|Others, like seed sown on good soil, hear the word, accept it, and produce a crop--thirty, sixty or even a hundred times what was sown."
MARK|4|21|He said to them, "Do you bring in a lamp to put it under a bowl or a bed? Instead, don't you put it on its stand?
MARK|4|22|For whatever is hidden is meant to be disclosed, and whatever is concealed is meant to be brought out into the open.
MARK|4|23|If anyone has ears to hear, let him hear."
MARK|4|24|"Consider carefully what you hear," he continued. "With the measure you use, it will be measured to you--and even more.
MARK|4|25|Whoever has will be given more; whoever does not have, even what he has will be taken from him."
MARK|4|26|He also said, "This is what the kingdom of God is like. A man scatters seed on the ground.
MARK|4|27|Night and day, whether he sleeps or gets up, the seed sprouts and grows, though he does not know how.
MARK|4|28|All by itself the soil produces grain--first the stalk, then the head, then the full kernel in the head.
MARK|4|29|As soon as the grain is ripe, he puts the sickle to it, because the harvest has come."
MARK|4|30|Again he said, "What shall we say the kingdom of God is like, or what parable shall we use to describe it?
MARK|4|31|It is like a mustard seed, which is the smallest seed you plant in the ground.
MARK|4|32|Yet when planted, it grows and becomes the largest of all garden plants, with such big branches that the birds of the air can perch in its shade."
MARK|4|33|With many similar parables Jesus spoke the word to them, as much as they could understand.
MARK|4|34|He did not say anything to them without using a parable. But when he was alone with his own disciples, he explained everything.
MARK|4|35|That day when evening came, he said to his disciples, "Let us go over to the other side."
MARK|4|36|Leaving the crowd behind, they took him along, just as he was, in the boat. There were also other boats with him.
MARK|4|37|A furious squall came up, and the waves broke over the boat, so that it was nearly swamped.
MARK|4|38|Jesus was in the stern, sleeping on a cushion. The disciples woke him and said to him, "Teacher, don't you care if we drown?"
MARK|4|39|He got up, rebuked the wind and said to the waves, "Quiet! Be still!" Then the wind died down and it was completely calm.
MARK|4|40|He said to his disciples, "Why are you so afraid? Do you still have no faith?"
MARK|4|41|They were terrified and asked each other, "Who is this? Even the wind and the waves obey him!"
MARK|5|1|They went across the lake to the region of the Gerasenes.
MARK|5|2|When Jesus got out of the boat, a man with an evil spirit came from the tombs to meet him.
MARK|5|3|This man lived in the tombs, and no one could bind him any more, not even with a chain.
MARK|5|4|For he had often been chained hand and foot, but he tore the chains apart and broke the irons on his feet. No one was strong enough to subdue him.
MARK|5|5|Night and day among the tombs and in the hills he would cry out and cut himself with stones.
MARK|5|6|When he saw Jesus from a distance, he ran and fell on his knees in front of him.
MARK|5|7|He shouted at the top of his voice, "What do you want with me, Jesus, Son of the Most High God? Swear to God that you won't torture me!"
MARK|5|8|For Jesus had said to him, "Come out of this man, you evil spirit!"
MARK|5|9|Then Jesus asked him, "What is your name?"
MARK|5|10|"My name is Legion," he replied, "for we are many." And he begged Jesus again and again not to send them out of the area.
MARK|5|11|A large herd of pigs was feeding on the nearby hillside.
MARK|5|12|The demons begged Jesus, "Send us among the pigs; allow us to go into them."
MARK|5|13|He gave them permission, and the evil spirits came out and went into the pigs. The herd, about two thousand in number, rushed down the steep bank into the lake and were drowned.
MARK|5|14|Those tending the pigs ran off and reported this in the town and countryside, and the people went out to see what had happened.
MARK|5|15|When they came to Jesus, they saw the man who had been possessed by the legion of demons, sitting there, dressed and in his right mind; and they were afraid.
MARK|5|16|Those who had seen it told the people what had happened to the demon-possessed man--and told about the pigs as well.
MARK|5|17|Then the people began to plead with Jesus to leave their region.
MARK|5|18|As Jesus was getting into the boat, the man who had been demon-possessed begged to go with him.
MARK|5|19|Jesus did not let him, but said, "Go home to your family and tell them how much the Lord has done for you, and how he has had mercy on you."
MARK|5|20|So the man went away and began to tell in the Decapolis how much Jesus had done for him. And all the people were amazed.
MARK|5|21|When Jesus had again crossed over by boat to the other side of the lake, a large crowd gathered around him while he was by the lake.
MARK|5|22|Then one of the synagogue rulers, named Jairus, came there. Seeing Jesus, he fell at his feet
MARK|5|23|and pleaded earnestly with him, "My little daughter is dying. Please come and put your hands on her so that she will be healed and live."
MARK|5|24|So Jesus went with him.
MARK|5|25|A large crowd followed and pressed around him. And a woman was there who had been subject to bleeding for twelve years.
MARK|5|26|She had suffered a great deal under the care of many doctors and had spent all she had, yet instead of getting better she grew worse.
MARK|5|27|When she heard about Jesus, she came up behind him in the crowd and touched his cloak,
MARK|5|28|because she thought, "If I just touch his clothes, I will be healed."
MARK|5|29|Immediately her bleeding stopped and she felt in her body that she was freed from her suffering.
MARK|5|30|At once Jesus realized that power had gone out from him. He turned around in the crowd and asked, "Who touched my clothes?"
MARK|5|31|"You see the people crowding against you," his disciples answered, "and yet you can ask, 'Who touched me?'"
MARK|5|32|But Jesus kept looking around to see who had done it.
MARK|5|33|Then the woman, knowing what had happened to her, came and fell at his feet and, trembling with fear, told him the whole truth.
MARK|5|34|He said to her, "Daughter, your faith has healed you. Go in peace and be freed from your suffering."
MARK|5|35|While Jesus was still speaking, some men came from the house of Jairus, the synagogue ruler. "Your daughter is dead," they said. "Why bother the teacher any more?"
MARK|5|36|Ignoring what they said, Jesus told the synagogue ruler, "Don't be afraid; just believe."
MARK|5|37|He did not let anyone follow him except Peter, James and John the brother of James.
MARK|5|38|When they came to the home of the synagogue ruler, Jesus saw a commotion, with people crying and wailing loudly.
MARK|5|39|He went in and said to them, "Why all this commotion and wailing? The child is not dead but asleep."
MARK|5|40|But they laughed at him.
MARK|5|41|After he put them all out, he took the child's father and mother and the disciples who were with him, and went in where the child was. He took her by the hand and said to her, "Talitha koum!" (which means, "Little girl, I say to you, get up!" ).
MARK|5|42|Immediately the girl stood up and walked around (she was twelve years old). At this they were completely astonished.
MARK|5|43|He gave strict orders not to let anyone know about this, and told them to give her something to eat.
MARK|6|1|Jesus left there and went to his hometown, accompanied by his disciples.
MARK|6|2|When the Sabbath came, he began to teach in the synagogue, and many who heard him were amazed.
MARK|6|3|"Where did this man get these things?" they asked. "What's this wisdom that has been given him, that he even does miracles! Isn't this the carpenter? Isn't this Mary's son and the brother of James, Joseph, Judas and Simon? Aren't his sisters here with us?" And they took offense at him.
MARK|6|4|Jesus said to them, "Only in his hometown, among his relatives and in his own house is a prophet without honor."
MARK|6|5|He could not do any miracles there, except lay his hands on a few sick people and heal them.
MARK|6|6|And he was amazed at their lack of faith.
MARK|6|7|Then Jesus went around teaching from village to village. Calling the Twelve to him, he sent them out two by two and gave them authority over evil spirits.
MARK|6|8|These were his instructions: "Take nothing for the journey except a staff--no bread, no bag, no money in your belts.
MARK|6|9|Wear sandals but not an extra tunic.
MARK|6|10|Whenever you enter a house, stay there until you leave that town.
MARK|6|11|And if any place will not welcome you or listen to you, shake the dust off your feet when you leave, as a testimony against them."
MARK|6|12|They went out and preached that people should repent.
MARK|6|13|They drove out many demons and anointed many sick people with oil and healed them.
MARK|6|14|King Herod heard about this, for Jesus' name had become well known. Some were saying, "John the Baptist has been raised from the dead, and that is why miraculous powers are at work in him."
MARK|6|15|Others said, "He is Elijah." And still others claimed, "He is a prophet, like one of the prophets of long ago."
MARK|6|16|But when Herod heard this, he said, "John, the man I beheaded, has been raised from the dead!"
MARK|6|17|For Herod himself had given orders to have John arrested, and he had him bound and put in prison. He did this because of Herodias, his brother Philip's wife, whom he had married.
MARK|6|18|For John had been saying to Herod, "It is not lawful for you to have your brother's wife."
MARK|6|19|So Herodias nursed a grudge against John and wanted to kill him. But she was not able to,
MARK|6|20|because Herod feared John and protected him, knowing him to be a righteous and holy man. When Herod heard John, he was greatly puzzled; yet he liked to listen to him.
MARK|6|21|Finally the opportune time came. On his birthday Herod gave a banquet for his high officials and military commanders and the leading men of Galilee.
MARK|6|22|When the daughter of Herodias came in and danced, she pleased Herod and his dinner guests.
MARK|6|23|The king said to the girl, "Ask me for anything you want, and I'll give it to you." And he promised her with an oath, "Whatever you ask I will give you, up to half my kingdom."
MARK|6|24|She went out and said to her mother, "What shall I ask for?The head of John the Baptist," she answered.
MARK|6|25|At once the girl hurried in to the king with the request: "I want you to give me right now the head of John the Baptist on a platter."
MARK|6|26|The king was greatly distressed, but because of his oaths and his dinner guests, he did not want to refuse her.
MARK|6|27|So he immediately sent an executioner with orders to bring John's head. The man went, beheaded John in the prison,
MARK|6|28|and brought back his head on a platter. He presented it to the girl, and she gave it to her mother.
MARK|6|29|On hearing of this, John's disciples came and took his body and laid it in a tomb.
MARK|6|30|The apostles gathered around Jesus and reported to him all they had done and taught.
MARK|6|31|Then, because so many people were coming and going that they did not even have a chance to eat, he said to them, "Come with me by yourselves to a quiet place and get some rest."
MARK|6|32|So they went away by themselves in a boat to a solitary place.
MARK|6|33|But many who saw them leaving recognized them and ran on foot from all the towns and got there ahead of them.
MARK|6|34|When Jesus landed and saw a large crowd, he had compassion on them, because they were like sheep without a shepherd. So he began teaching them many things.
MARK|6|35|By this time it was late in the day, so his disciples came to him. "This is a remote place," they said, "and it's already very late.
MARK|6|36|Send the people away so they can go to the surrounding countryside and villages and buy themselves something to eat."
MARK|6|37|But he answered, "You give them something to eat." They said to him, "That would take eight months of a man's wages! Are we to go and spend that much on bread and give it to them to eat?"
MARK|6|38|"How many loaves do you have?" he asked. "Go and see." When they found out, they said, "Five--and two fish."
MARK|6|39|Then Jesus directed them to have all the people sit down in groups on the green grass.
MARK|6|40|So they sat down in groups of hundreds and fifties.
MARK|6|41|Taking the five loaves and the two fish and looking up to heaven, he gave thanks and broke the loaves. Then he gave them to his disciples to set before the people. He also divided the two fish among them all.
MARK|6|42|They all ate and were satisfied,
MARK|6|43|and the disciples picked up twelve basketfuls of broken pieces of bread and fish.
MARK|6|44|The number of the men who had eaten was five thousand.
MARK|6|45|Immediately Jesus made his disciples get into the boat and go on ahead of him to Bethsaida, while he dismissed the crowd.
MARK|6|46|After leaving them, he went up on a mountainside to pray.
MARK|6|47|When evening came, the boat was in the middle of the lake, and he was alone on land.
MARK|6|48|He saw the disciples straining at the oars, because the wind was against them. About the fourth watch of the night he went out to them, walking on the lake. He was about to pass by them,
MARK|6|49|but when they saw him walking on the lake, they thought he was a ghost. They cried out,
MARK|6|50|because they all saw him and were terrified.
MARK|6|51|Immediately he spoke to them and said, "Take courage! It is I. Don't be afraid." Then he climbed into the boat with them, and the wind died down. They were completely amazed,
MARK|6|52|for they had not understood about the loaves; their hearts were hardened.
MARK|6|53|When they had crossed over, they landed at Gennesaret and anchored there.
MARK|6|54|As soon as they got out of the boat, people recognized Jesus.
MARK|6|55|They ran throughout that whole region and carried the sick on mats to wherever they heard he was.
MARK|6|56|And wherever he went--into villages, towns or countryside--they placed the sick in the marketplaces. They begged him to let them touch even the edge of his cloak, and all who touched him were healed.
MARK|7|1|The Pharisees and some of the teachers of the law who had come from Jerusalem gathered around Jesus and
MARK|7|2|saw some of his disciples eating food with hands that were "unclean," that is, unwashed.
MARK|7|3|(The Pharisees and all the Jews do not eat unless they give their hands a ceremonial washing, holding to the tradition of the elders.
MARK|7|4|When they come from the marketplace they do not eat unless they wash. And they observe many other traditions, such as the washing of cups, pitchers and kettles. )
MARK|7|5|So the Pharisees and teachers of the law asked Jesus, "Why don't your disciples live according to the tradition of the elders instead of eating their food with 'unclean' hands?"
MARK|7|6|He replied, "Isaiah was right when he prophesied about you hypocrites; as it is written: "'These people honor me with their lips, but their hearts are far from me.
MARK|7|7|They worship me in vain; their teachings are but rules taught by men.'
MARK|7|8|You have let go of the commands of God and are holding on to the traditions of men."
MARK|7|9|And he said to them: "You have a fine way of setting aside the commands of God in order to observe your own traditions!
MARK|7|10|For Moses said, 'Honor your father and your mother,' and, 'Anyone who curses his father or mother must be put to death.'
MARK|7|11|But you say that if a man says to his father or mother: 'Whatever help you might otherwise have received from me is Corban' (that is, a gift devoted to God),
MARK|7|12|then you no longer let him do anything for his father or mother.
MARK|7|13|Thus you nullify the word of God by your tradition that you have handed down. And you do many things like that."
MARK|7|14|Again Jesus called the crowd to him and said, "Listen to me, everyone, and understand this.
MARK|7|15|Nothing outside a man can make him 'unclean' by going into him. Rather, it is what comes out of a man that makes him 'unclean.'"
MARK|7|16|See Footnote
MARK|7|17|After he had left the crowd and entered the house, his disciples asked him about this parable.
MARK|7|18|"Are you so dull?" he asked. "Don't you see that nothing that enters a man from the outside can make him 'unclean'?
MARK|7|19|For it doesn't go into his heart but into his stomach, and then out of his body." (In saying this, Jesus declared all foods "clean.")
MARK|7|20|He went on: "What comes out of a man is what makes him 'unclean.'
MARK|7|21|For from within, out of men's hearts, come evil thoughts, sexual immorality, theft, murder, adultery,
MARK|7|22|greed, malice, deceit, lewdness, envy, slander, arrogance and folly.
MARK|7|23|All these evils come from inside and make a man 'unclean.'"
MARK|7|24|Jesus left that place and went to the vicinity of Tyre. He entered a house and did not want anyone to know it; yet he could not keep his presence secret.
MARK|7|25|In fact, as soon as she heard about him, a woman whose little daughter was possessed by an evil spirit came and fell at his feet.
MARK|7|26|The woman was a Greek, born in Syrian Phoenicia. She begged Jesus to drive the demon out of her daughter.
MARK|7|27|"First let the children eat all they want," he told her, "for it is not right to take the children's bread and toss it to their dogs."
MARK|7|28|"Yes, Lord," she replied, "but even the dogs under the table eat the children's crumbs."
MARK|7|29|Then he told her, "For such a reply, you may go; the demon has left your daughter."
MARK|7|30|She went home and found her child lying on the bed, and the demon gone.
MARK|7|31|Then Jesus left the vicinity of Tyre and went through Sidon, down to the Sea of Galilee and into the region of the Decapolis.
MARK|7|32|There some people brought to him a man who was deaf and could hardly talk, and they begged him to place his hand on the man.
MARK|7|33|After he took him aside, away from the crowd, Jesus put his fingers into the man's ears. Then he spit and touched the man's tongue.
MARK|7|34|He looked up to heaven and with a deep sigh said to him, "Ephphatha!" (which means, "Be opened!" ).
MARK|7|35|At this, the man's ears were opened, his tongue was loosened and he began to speak plainly.
MARK|7|36|Jesus commanded them not to tell anyone. But the more he did so, the more they kept talking about it.
MARK|7|37|People were overwhelmed with amazement. "He has done everything well," they said. "He even makes the deaf hear and the mute speak."
MARK|8|1|During those days another large crowd gathered. Since they had nothing to eat, Jesus called his disciples to him and said,
MARK|8|2|"I have compassion for these people; they have already been with me three days and have nothing to eat.
MARK|8|3|If I send them home hungry, they will collapse on the way, because some of them have come a long distance."
MARK|8|4|His disciples answered, "But where in this remote place can anyone get enough bread to feed them?"
MARK|8|5|"How many loaves do you have?" Jesus asked. "Seven," they replied.
MARK|8|6|He told the crowd to sit down on the ground. When he had taken the seven loaves and given thanks, he broke them and gave them to his disciples to set before the people, and they did so.
MARK|8|7|They had a few small fish as well; he gave thanks for them also and told the disciples to distribute them.
MARK|8|8|The people ate and were satisfied. Afterward the disciples picked up seven basketfuls of broken pieces that were left over.
MARK|8|9|About four thousand men were present. And having sent them away,
MARK|8|10|he got into the boat with his disciples and went to the region of Dalmanutha.
MARK|8|11|The Pharisees came and began to question Jesus. To test him, they asked him for a sign from heaven.
MARK|8|12|He sighed deeply and said, "Why does this generation ask for a miraculous sign? I tell you the truth, no sign will be given to it."
MARK|8|13|Then he left them, got back into the boat and crossed to the other side.
MARK|8|14|The disciples had forgotten to bring bread, except for one loaf they had with them in the boat.
MARK|8|15|"Be careful," Jesus warned them. "Watch out for the yeast of the Pharisees and that of Herod."
MARK|8|16|They discussed this with one another and said, "It is because we have no bread."
MARK|8|17|Aware of their discussion, Jesus asked them: "Why are you talking about having no bread? Do you still not see or understand? Are your hearts hardened?
MARK|8|18|Do you have eyes but fail to see, and ears but fail to hear? And don't you remember?
MARK|8|19|When I broke the five loaves for the five thousand, how many basketfuls of pieces did you pick up?Twelve," they replied.
MARK|8|20|"And when I broke the seven loaves for the four thousand, how many basketfuls of pieces did you pick up?" They answered, "Seven."
MARK|8|21|He said to them, "Do you still not understand?"
MARK|8|22|They came to Bethsaida, and some people brought a blind man and begged Jesus to touch him.
MARK|8|23|He took the blind man by the hand and led him outside the village. When he had spit on the man's eyes and put his hands on him, Jesus asked, "Do you see anything?"
MARK|8|24|He looked up and said, "I see people; they look like trees walking around."
MARK|8|25|Once more Jesus put his hands on the man's eyes. Then his eyes were opened, his sight was restored, and he saw everything clearly.
MARK|8|26|Jesus sent him home, saying, "Don't go into the village. "
MARK|8|27|Jesus and his disciples went on to the villages around Caesarea Philippi. On the way he asked them, "Who do people say I am?"
MARK|8|28|They replied, "Some say John the Baptist; others say Elijah; and still others, one of the prophets."
MARK|8|29|"But what about you?" he asked. "Who do you say I am?" Peter answered, "You are the Christ. "
MARK|8|30|Jesus warned them not to tell anyone about him.
MARK|8|31|He then began to teach them that the Son of Man must suffer many things and be rejected by the elders, chief priests and teachers of the law, and that he must be killed and after three days rise again.
MARK|8|32|He spoke plainly about this, and Peter took him aside and began to rebuke him.
MARK|8|33|But when Jesus turned and looked at his disciples, he rebuked Peter. "Get behind me, Satan!" he said. "You do not have in mind the things of God, but the things of men."
MARK|8|34|Then he called the crowd to him along with his disciples and said: "If anyone would come after me, he must deny himself and take up his cross and follow me.
MARK|8|35|For whoever wants to save his life will lose it, but whoever loses his life for me and for the gospel will save it.
MARK|8|36|What good is it for a man to gain the whole world, yet forfeit his soul?
MARK|8|37|Or what can a man give in exchange for his soul?
MARK|8|38|If anyone is ashamed of me and my words in this adulterous and sinful generation, the Son of Man will be ashamed of him when he comes in his Father's glory with the holy angels."
MARK|9|1|And he said to them, "I tell you the truth, some who are standing here will not taste death before they see the kingdom of God come with power."
MARK|9|2|After six days Jesus took Peter, James and John with him and led them up a high mountain, where they were all alone. There he was transfigured before them.
MARK|9|3|His clothes became dazzling white, whiter than anyone in the world could bleach them.
MARK|9|4|And there appeared before them Elijah and Moses, who were talking with Jesus.
MARK|9|5|Peter said to Jesus, "Rabbi, it is good for us to be here. Let us put up three shelters--one for you, one for Moses and one for Elijah."
MARK|9|6|(He did not know what to say, they were so frightened.)
MARK|9|7|Then a cloud appeared and enveloped them, and a voice came from the cloud: "This is my Son, whom I love. Listen to him!"
MARK|9|8|Suddenly, when they looked around, they no longer saw anyone with them except Jesus.
MARK|9|9|As they were coming down the mountain, Jesus gave them orders not to tell anyone what they had seen until the Son of Man had risen from the dead.
MARK|9|10|They kept the matter to themselves, discussing what "rising from the dead" meant.
MARK|9|11|And they asked him, "Why do the teachers of the law say that Elijah must come first?"
MARK|9|12|Jesus replied, "To be sure, Elijah does come first, and restores all things. Why then is it written that the Son of Man must suffer much and be rejected?
MARK|9|13|But I tell you, Elijah has come, and they have done to him everything they wished, just as it is written about him."
MARK|9|14|When they came to the other disciples, they saw a large crowd around them and the teachers of the law arguing with them.
MARK|9|15|As soon as all the people saw Jesus, they were overwhelmed with wonder and ran to greet him.
MARK|9|16|"What are you arguing with them about?" he asked.
MARK|9|17|A man in the crowd answered, "Teacher, I brought you my son, who is possessed by a spirit that has robbed him of speech.
MARK|9|18|Whenever it seizes him, it throws him to the ground. He foams at the mouth, gnashes his teeth and becomes rigid. I asked your disciples to drive out the spirit, but they could not."
MARK|9|19|"O unbelieving generation," Jesus replied, "how long shall I stay with you? How long shall I put up with you? Bring the boy to me."
MARK|9|20|So they brought him. When the spirit saw Jesus, it immediately threw the boy into a convulsion. He fell to the ground and rolled around, foaming at the mouth.
MARK|9|21|Jesus asked the boy's father, "How long has he been like this?"
MARK|9|22|"From childhood," he answered. "It has often thrown him into fire or water to kill him. But if you can do anything, take pity on us and help us."
MARK|9|23|"'If you can'?" said Jesus. "Everything is possible for him who believes."
MARK|9|24|Immediately the boy's father exclaimed, "I do believe; help me overcome my unbelief!"
MARK|9|25|When Jesus saw that a crowd was running to the scene, he rebuked the evil spirit. "You deaf and mute spirit," he said, "I command you, come out of him and never enter him again."
MARK|9|26|The spirit shrieked, convulsed him violently and came out. The boy looked so much like a corpse that many said, "He's dead."
MARK|9|27|But Jesus took him by the hand and lifted him to his feet, and he stood up.
MARK|9|28|After Jesus had gone indoors, his disciples asked him privately, "Why couldn't we drive it out?"
MARK|9|29|He replied, "This kind can come out only by prayer. "
MARK|9|30|They left that place and passed through Galilee. Jesus did not want anyone to know where they were,
MARK|9|31|because he was teaching his disciples. He said to them, "The Son of Man is going to be betrayed into the hands of men. They will kill him, and after three days he will rise."
MARK|9|32|But they did not understand what he meant and were afraid to ask him about it.
MARK|9|33|They came to Capernaum. When he was in the house, he asked them, "What were you arguing about on the road?"
MARK|9|34|But they kept quiet because on the way they had argued about who was the greatest.
MARK|9|35|Sitting down, Jesus called the Twelve and said, "If anyone wants to be first, he must be the very last, and the servant of all."
MARK|9|36|He took a little child and had him stand among them. Taking him in his arms, he said to them,
MARK|9|37|"Whoever welcomes one of these little children in my name welcomes me; and whoever welcomes me does not welcome me but the one who sent me."
MARK|9|38|"Teacher," said John, "we saw a man driving out demons in your name and we told him to stop, because he was not one of us."
MARK|9|39|"Do not stop him," Jesus said. "No one who does a miracle in my name can in the next moment say anything bad about me,
MARK|9|40|for whoever is not against us is for us.
MARK|9|41|I tell you the truth, anyone who gives you a cup of water in my name because you belong to Christ will certainly not lose his reward.
MARK|9|42|"And if anyone causes one of these little ones who believe in me to sin, it would be better for him to be thrown into the sea with a large millstone tied around his neck.
MARK|9|43|If your hand causes you to sin, cut it off. It is better for you to enter life maimed than with two hands to go into hell, where the fire never goes out.
MARK|9|44|See Footnote
MARK|9|45|And if your foot causes you to sin, cut it off. It is better for you to enter life crippled than to have two feet and be thrown into hell.
MARK|9|46|See Footnote
MARK|9|47|And if your eye causes you to sin, pluck it out. It is better for you to enter the kingdom of God with one eye than to have two eyes and be thrown into hell,
MARK|9|48|where "'their worm does not die, and the fire is not quenched.'
MARK|9|49|Everyone will be salted with fire.
MARK|9|50|"Salt is good, but if it loses its saltiness, how can you make it salty again? Have salt in yourselves, and be at peace with each other."
MARK|10|1|Jesus then left that place and went into the region of Judea and across the Jordan. Again crowds of people came to him, and as was his custom, he taught them.
MARK|10|2|Some Pharisees came and tested him by asking, "Is it lawful for a man to divorce his wife?"
MARK|10|3|"What did Moses command you?" he replied.
MARK|10|4|They said, "Moses permitted a man to write a certificate of divorce and send her away."
MARK|10|5|"It was because your hearts were hard that Moses wrote you this law," Jesus replied.
MARK|10|6|"But at the beginning of creation God 'made them male and female.'
MARK|10|7|'For this reason a man will leave his father and mother and be united to his wife,
MARK|10|8|and the two will become one flesh.' So they are no longer two, but one.
MARK|10|9|Therefore what God has joined together, let man not separate."
MARK|10|10|When they were in the house again, the disciples asked Jesus about this.
MARK|10|11|He answered, "Anyone who divorces his wife and marries another woman commits adultery against her.
MARK|10|12|And if she divorces her husband and marries another man, she commits adultery."
MARK|10|13|People were bringing little children to Jesus to have him touch them, but the disciples rebuked them.
MARK|10|14|When Jesus saw this, he was indignant. He said to them, "Let the little children come to me, and do not hinder them, for the kingdom of God belongs to such as these.
MARK|10|15|I tell you the truth, anyone who will not receive the kingdom of God like a little child will never enter it."
MARK|10|16|And he took the children in his arms, put his hands on them and blessed them.
MARK|10|17|As Jesus started on his way, a man ran up to him and fell on his knees before him. "Good teacher," he asked, "what must I do to inherit eternal life?"
MARK|10|18|"Why do you call me good?" Jesus answered. "No one is good--except God alone.
MARK|10|19|You know the commandments: 'Do not murder, do not commit adultery, do not steal, do not give false testimony, do not defraud, honor your father and mother.'"
MARK|10|20|"Teacher," he declared, "all these I have kept since I was a boy."
MARK|10|21|Jesus looked at him and loved him. "One thing you lack," he said. "Go, sell everything you have and give to the poor, and you will have treasure in heaven. Then come, follow me."
MARK|10|22|At this the man's face fell. He went away sad, because he had great wealth.
MARK|10|23|Jesus looked around and said to his disciples, "How hard it is for the rich to enter the kingdom of God!"
MARK|10|24|The disciples were amazed at his words. But Jesus said again, "Children, how hard it is to enter the kingdom of God!
MARK|10|25|It is easier for a camel to go through the eye of a needle than for a rich man to enter the kingdom of God."
MARK|10|26|The disciples were even more amazed, and said to each other, "Who then can be saved?"
MARK|10|27|Jesus looked at them and said, "With man this is impossible, but not with God; all things are possible with God."
MARK|10|28|Peter said to him, "We have left everything to follow you!"
MARK|10|29|"I tell you the truth," Jesus replied, "no one who has left home or brothers or sisters or mother or father or children or fields for me and the gospel
MARK|10|30|will fail to receive a hundred times as much in this present age (homes, brothers, sisters, mothers, children and fields--and with them, persecutions) and in the age to come, eternal life.
MARK|10|31|But many who are first will be last, and the last first."
MARK|10|32|They were on their way up to Jerusalem, with Jesus leading the way, and the disciples were astonished, while those who followed were afraid. Again he took the Twelve aside and told them what was going to happen to him.
MARK|10|33|"We are going up to Jerusalem," he said, "and the Son of Man will be betrayed to the chief priests and teachers of the law. They will condemn him to death and will hand him over to the Gentiles,
MARK|10|34|who will mock him and spit on him, flog him and kill him. Three days later he will rise."
MARK|10|35|Then James and John, the sons of Zebedee, came to him. "Teacher," they said, "we want you to do for us whatever we ask."
MARK|10|36|"What do you want me to do for you?" he asked.
MARK|10|37|They replied, "Let one of us sit at your right and the other at your left in your glory."
MARK|10|38|"You don't know what you are asking," Jesus said. "Can you drink the cup I drink or be baptized with the baptism I am baptized with?"
MARK|10|39|"We can," they answered. Jesus said to them, "You will drink the cup I drink and be baptized with the baptism I am baptized with,
MARK|10|40|but to sit at my right or left is not for me to grant. These places belong to those for whom they have been prepared."
MARK|10|41|When the ten heard about this, they became indignant with James and John.
MARK|10|42|Jesus called them together and said, "You know that those who are regarded as rulers of the Gentiles lord it over them, and their high officials exercise authority over them.
MARK|10|43|Not so with you. Instead, whoever wants to become great among you must be your servant,
MARK|10|44|and whoever wants to be first must be slave of all.
MARK|10|45|For even the Son of Man did not come to be served, but to serve, and to give his life as a ransom for many."
MARK|10|46|Then they came to Jericho. As Jesus and his disciples, together with a large crowd, were leaving the city, a blind man, Bartimaeus (that is, the Son of Timaeus), was sitting by the roadside begging.
MARK|10|47|When he heard that it was Jesus of Nazareth, he began to shout, "Jesus, Son of David, have mercy on me!"
MARK|10|48|Many rebuked him and told him to be quiet, but he shouted all the more, "Son of David, have mercy on me!"
MARK|10|49|Jesus stopped and said, "Call him." So they called to the blind man, "Cheer up! On your feet! He's calling you."
MARK|10|50|Throwing his cloak aside, he jumped to his feet and came to Jesus.
MARK|10|51|"What do you want me to do for you?" Jesus asked him. The blind man said, "Rabbi, I want to see."
MARK|10|52|"Go," said Jesus, "your faith has healed you." Immediately he received his sight and followed Jesus along the road.
MARK|11|1|As they approached Jerusalem and came to Bethphage and Bethany at the Mount of Olives, Jesus sent two of his disciples,
MARK|11|2|saying to them, "Go to the village ahead of you, and just as you enter it, you will find a colt tied there, which no one has ever ridden. Untie it and bring it here.
MARK|11|3|If anyone asks you, 'Why are you doing this?' tell him, 'The Lord needs it and will send it back here shortly.'"
MARK|11|4|They went and found a colt outside in the street, tied at a doorway. As they untied it,
MARK|11|5|some people standing there asked, "What are you doing, untying that colt?"
MARK|11|6|They answered as Jesus had told them to, and the people let them go.
MARK|11|7|When they brought the colt to Jesus and threw their cloaks over it, he sat on it.
MARK|11|8|Many people spread their cloaks on the road, while others spread branches they had cut in the fields.
MARK|11|9|Those who went ahead and those who followed shouted, "Hosanna! Blessed is he who comes in the name of the Lord!"
MARK|11|10|"Blessed is the coming kingdom of our father David!Hosanna in the highest!"
MARK|11|11|Jesus entered Jerusalem and went to the temple. He looked around at everything, but since it was already late, he went out to Bethany with the Twelve.
MARK|11|12|The next day as they were leaving Bethany, Jesus was hungry.
MARK|11|13|Seeing in the distance a fig tree in leaf, he went to find out if it had any fruit. When he reached it, he found nothing but leaves, because it was not the season for figs.
MARK|11|14|Then he said to the tree, "May no one ever eat fruit from you again." And his disciples heard him say it.
MARK|11|15|On reaching Jerusalem, Jesus entered the temple area and began driving out those who were buying and selling there. He overturned the tables of the money changers and the benches of those selling doves,
MARK|11|16|and would not allow anyone to carry merchandise through the temple courts.
MARK|11|17|And as he taught them, he said, "Is it not written: "'My house will be called a house of prayer for all nations'? But you have made it 'a den of robbers.'"
MARK|11|18|The chief priests and the teachers of the law heard this and began looking for a way to kill him, for they feared him, because the whole crowd was amazed at his teaching.
MARK|11|19|When evening came, they went out of the city.
MARK|11|20|In the morning, as they went along, they saw the fig tree withered from the roots.
MARK|11|21|Peter remembered and said to Jesus, "Rabbi, look! The fig tree you cursed has withered!"
MARK|11|22|"Have faith in God," Jesus answered.
MARK|11|23|"I tell you the truth, if anyone says to this mountain, 'Go, throw yourself into the sea,' and does not doubt in his heart but believes that what he says will happen, it will be done for him.
MARK|11|24|Therefore I tell you, whatever you ask for in prayer, believe that you have received it, and it will be yours.
MARK|11|25|And when you stand praying, if you hold anything against anyone, forgive him, so that your Father in heaven may forgive you your sins."
MARK|11|26|See Footnote
MARK|11|27|They arrived again in Jerusalem, and while Jesus was walking in the temple courts, the chief priests, the teachers of the law and the elders came to him.
MARK|11|28|"By what authority are you doing these things?" they asked. "And who gave you authority to do this?"
MARK|11|29|Jesus replied, "I will ask you one question. Answer me, and I will tell you by what authority I am doing these things.
MARK|11|30|John's baptism--was it from heaven, or from men? Tell me!"
MARK|11|31|They discussed it among themselves and said, "If we say, 'From heaven,' he will ask, 'Then why didn't you believe him?'
MARK|11|32|But if we say, 'From men'...." (They feared the people, for everyone held that John really was a prophet.)
MARK|11|33|So they answered Jesus, "We don't know." Jesus said, "Neither will I tell you by what authority I am doing these things."
MARK|12|1|He then began to speak to them in parables: "A man planted a vineyard. He put a wall around it, dug a pit for the winepress and built a watchtower. Then he rented the vineyard to some farmers and went away on a journey.
MARK|12|2|At harvest time he sent a servant to the tenants to collect from them some of the fruit of the vineyard.
MARK|12|3|But they seized him, beat him and sent him away empty-handed.
MARK|12|4|Then he sent another servant to them; they struck this man on the head and treated him shamefully.
MARK|12|5|He sent still another, and that one they killed. He sent many others; some of them they beat, others they killed.
MARK|12|6|"He had one left to send, a son, whom he loved. He sent him last of all, saying, 'They will respect my son.'
MARK|12|7|"But the tenants said to one another, 'This is the heir. Come, let's kill him, and the inheritance will be ours.'
MARK|12|8|So they took him and killed him, and threw him out of the vineyard.
MARK|12|9|"What then will the owner of the vineyard do? He will come and kill those tenants and give the vineyard to others.
MARK|12|10|Haven't you read this scripture: "'The stone the builders rejected has become the capstone;
MARK|12|11|the Lord has done this, and it is marvelous in our eyes'?"
MARK|12|12|Then they looked for a way to arrest him because they knew he had spoken the parable against them. But they were afraid of the crowd; so they left him and went away.
MARK|12|13|Later they sent some of the Pharisees and Herodians to Jesus to catch him in his words.
MARK|12|14|They came to him and said, "Teacher, we know you are a man of integrity. You aren't swayed by men, because you pay no attention to who they are; but you teach the way of God in accordance with the truth. Is it right to pay taxes to Caesar or not?
MARK|12|15|Should we pay or shouldn't we?"
MARK|12|16|But Jesus knew their hypocrisy. "Why are you trying to trap me?" he asked. "Bring me a denarius and let me look at it." They brought the coin, and he asked them, "Whose portrait is this? And whose inscription?Caesar's," they replied.
MARK|12|17|Then Jesus said to them, "Give to Caesar what is Caesar's and to God what is God's." And they were amazed at him.
MARK|12|18|Then the Sadducees, who say there is no resurrection, came to him with a question.
MARK|12|19|"Teacher," they said, "Moses wrote for us that if a man's brother dies and leaves a wife but no children, the man must marry the widow and have children for his brother.
MARK|12|20|Now there were seven brothers. The first one married and died without leaving any children.
MARK|12|21|The second one married the widow, but he also died, leaving no child. It was the same with the third.
MARK|12|22|In fact, none of the seven left any children. Last of all, the woman died too.
MARK|12|23|At the resurrection whose wife will she be, since the seven were married to her?"
MARK|12|24|Jesus replied, "Are you not in error because you do not know the Scriptures or the power of God?
MARK|12|25|When the dead rise, they will neither marry nor be given in marriage; they will be like the angels in heaven.
MARK|12|26|Now about the dead rising--have you not read in the book of Moses, in the account of the bush, how God said to him, 'I am the God of Abraham, the God of Isaac, and the God of Jacob'?
MARK|12|27|He is not the God of the dead, but of the living. You are badly mistaken!"
MARK|12|28|One of the teachers of the law came and heard them debating. Noticing that Jesus had given them a good answer, he asked him, "Of all the commandments, which is the most important?"
MARK|12|29|"The most important one," answered Jesus, "is this: 'Hear, O Israel, the Lord our God, the Lord is one.
MARK|12|30|Love the Lord your God with all your heart and with all your soul and with all your mind and with all your strength.'
MARK|12|31|The second is this: 'Love your neighbor as yourself.' There is no commandment greater than these."
MARK|12|32|"Well said, teacher," the man replied. "You are right in saying that God is one and there is no other but him.
MARK|12|33|To love him with all your heart, with all your understanding and with all your strength, and to love your neighbor as yourself is more important than all burnt offerings and sacrifices."
MARK|12|34|When Jesus saw that he had answered wisely, he said to him, "You are not far from the kingdom of God." And from then on no one dared ask him any more questions.
MARK|12|35|While Jesus was teaching in the temple courts, he asked, "How is it that the teachers of the law say that the Christ is the son of David?
MARK|12|36|David himself, speaking by the Holy Spirit, declared: "'The Lord said to my Lord: "Sit at my right hand until I put your enemies under your feet."'
MARK|12|37|David himself calls him 'Lord.' How then can he be his son?" The large crowd listened to him with delight.
MARK|12|38|As he taught, Jesus said, "Watch out for the teachers of the law. They like to walk around in flowing robes and be greeted in the marketplaces,
MARK|12|39|and have the most important seats in the synagogues and the places of honor at banquets.
MARK|12|40|They devour widows' houses and for a show make lengthy prayers. Such men will be punished most severely."
MARK|12|41|Jesus sat down opposite the place where the offerings were put and watched the crowd putting their money into the temple treasury. Many rich people threw in large amounts.
MARK|12|42|But a poor widow came and put in two very small copper coins, worth only a fraction of a penny.
MARK|12|43|Calling his disciples to him, Jesus said, "I tell you the truth, this poor widow has put more into the treasury than all the others.
MARK|12|44|They all gave out of their wealth; but she, out of her poverty, put in everything--all she had to live on."
MARK|13|1|As he was leaving the temple, one of his disciples said to him, "Look, Teacher! What massive stones! What magnificent buildings!"
MARK|13|2|"Do you see all these great buildings?" replied Jesus. "Not one stone here will be left on another; every one will be thrown down."
MARK|13|3|As Jesus was sitting on the Mount of Olives opposite the temple, Peter, James, John and Andrew asked him privately,
MARK|13|4|"Tell us, when will these things happen? And what will be the sign that they are all about to be fulfilled?"
MARK|13|5|Jesus said to them: "Watch out that no one deceives you.
MARK|13|6|Many will come in my name, claiming, 'I am he,' and will deceive many.
MARK|13|7|When you hear of wars and rumors of wars, do not be alarmed. Such things must happen, but the end is still to come.
MARK|13|8|Nation will rise against nation, and kingdom against kingdom. There will be earthquakes in various places, and famines. These are the beginning of birth pains.
MARK|13|9|"You must be on your guard. You will be handed over to the local councils and flogged in the synagogues. On account of me you will stand before governors and kings as witnesses to them.
MARK|13|10|And the gospel must first be preached to all nations.
MARK|13|11|Whenever you are arrested and brought to trial, do not worry beforehand about what to say. Just say whatever is given you at the time, for it is not you speaking, but the Holy Spirit.
MARK|13|12|"Brother will betray brother to death, and a father his child. Children will rebel against their parents and have them put to death.
MARK|13|13|All men will hate you because of me, but he who stands firm to the end will be saved.
MARK|13|14|"When you see 'the abomination that causes desolation' standing where it does not belong--let the reader understand--then let those who are in Judea flee to the mountains.
MARK|13|15|Let no one on the roof of his house go down or enter the house to take anything out.
MARK|13|16|Let no one in the field go back to get his cloak.
MARK|13|17|How dreadful it will be in those days for pregnant women and nursing mothers!
MARK|13|18|Pray that this will not take place in winter,
MARK|13|19|because those will be days of distress unequaled from the beginning, when God created the world, until now--and never to be equaled again.
MARK|13|20|If the Lord had not cut short those days, no one would survive. But for the sake of the elect, whom he has chosen, he has shortened them.
MARK|13|21|At that time if anyone says to you, 'Look, here is the Christ!' or, 'Look, there he is!' do not believe it.
MARK|13|22|For false Christs and false prophets will appear and perform signs and miracles to deceive the elect--if that were possible.
MARK|13|23|So be on your guard; I have told you everything ahead of time.
MARK|13|24|"But in those days, following that distress, "'the sun will be darkened, and the moon will not give its light;
MARK|13|25|the stars will fall from the sky, and the heavenly bodies will be shaken.'
MARK|13|26|"At that time men will see the Son of Man coming in clouds with great power and glory.
MARK|13|27|And he will send his angels and gather his elect from the four winds, from the ends of the earth to the ends of the heavens.
MARK|13|28|"Now learn this lesson from the fig tree: As soon as its twigs get tender and its leaves come out, you know that summer is near.
MARK|13|29|Even so, when you see these things happening, you know that it is near, right at the door.
MARK|13|30|I tell you the truth, this generation will certainly not pass away until all these things have happened.
MARK|13|31|Heaven and earth will pass away, but my words will never pass away.
MARK|13|32|"No one knows about that day or hour, not even the angels in heaven, nor the Son, but only the Father.
MARK|13|33|Be on guard! Be alert! You do not know when that time will come.
MARK|13|34|It's like a man going away: He leaves his house and puts his servants in charge, each with his assigned task, and tells the one at the door to keep watch.
MARK|13|35|"Therefore keep watch because you do not know when the owner of the house will come back--whether in the evening, or at midnight, or when the rooster crows, or at dawn.
MARK|13|36|If he comes suddenly, do not let him find you sleeping.
MARK|13|37|What I say to you, I say to everyone: 'Watch!'"
MARK|14|1|Now the Passover and the Feast of Unleavened Bread were only two days away, and the chief priests and the teachers of the law were looking for some sly way to arrest Jesus and kill him.
MARK|14|2|"But not during the Feast," they said, "or the people may riot."
MARK|14|3|While he was in Bethany, reclining at the table in the home of a man known as Simon the Leper, a woman came with an alabaster jar of very expensive perfume, made of pure nard. She broke the jar and poured the perfume on his head.
MARK|14|4|Some of those present were saying indignantly to one another, "Why this waste of perfume?
MARK|14|5|It could have been sold for more than a year's wages and the money given to the poor." And they rebuked her harshly.
MARK|14|6|"Leave her alone," said Jesus. "Why are you bothering her? She has done a beautiful thing to me.
MARK|14|7|The poor you will always have with you, and you can help them any time you want. But you will not always have me.
MARK|14|8|She did what she could. She poured perfume on my body beforehand to prepare for my burial.
MARK|14|9|I tell you the truth, wherever the gospel is preached throughout the world, what she has done will also be told, in memory of her."
MARK|14|10|Then Judas Iscariot, one of the Twelve, went to the chief priests to betray Jesus to them.
MARK|14|11|They were delighted to hear this and promised to give him money. So he watched for an opportunity to hand him over.
MARK|14|12|On the first day of the Feast of Unleavened Bread, when it was customary to sacrifice the Passover lamb, Jesus' disciples asked him, "Where do you want us to go and make preparations for you to eat the Passover?"
MARK|14|13|So he sent two of his disciples, telling them, "Go into the city, and a man carrying a jar of water will meet you. Follow him.
MARK|14|14|Say to the owner of the house he enters, 'The Teacher asks: Where is my guest room, where I may eat the Passover with my disciples?'
MARK|14|15|He will show you a large upper room, furnished and ready. Make preparations for us there."
MARK|14|16|The disciples left, went into the city and found things just as Jesus had told them. So they prepared the Passover.
MARK|14|17|When evening came, Jesus arrived with the Twelve.
MARK|14|18|While they were reclining at the table eating, he said, "I tell you the truth, one of you will betray me--one who is eating with me."
MARK|14|19|They were saddened, and one by one they said to him, "Surely not I?"
MARK|14|20|"It is one of the Twelve," he replied, "one who dips bread into the bowl with me.
MARK|14|21|The Son of Man will go just as it is written about him. But woe to that man who betrays the Son of Man! It would be better for him if he had not been born."
MARK|14|22|While they were eating, Jesus took bread, gave thanks and broke it, and gave it to his disciples, saying, "Take it; this is my body."
MARK|14|23|Then he took the cup, gave thanks and offered it to them, and they all drank from it.
MARK|14|24|"This is my blood of the covenant, which is poured out for many," he said to them.
MARK|14|25|"I tell you the truth, I will not drink again of the fruit of the vine until that day when I drink it anew in the kingdom of God."
MARK|14|26|When they had sung a hymn, they went out to the Mount of Olives.
MARK|14|27|"You will all fall away," Jesus told them, "for it is written: "'I will strike the shepherd, and the sheep will be scattered.'
MARK|14|28|But after I have risen, I will go ahead of you into Galilee."
MARK|14|29|Peter declared, "Even if all fall away, I will not."
MARK|14|30|"I tell you the truth," Jesus answered, "today--yes, tonight--before the rooster crows twice you yourself will disown me three times."
MARK|14|31|But Peter insisted emphatically, "Even if I have to die with you, I will never disown you." And all the others said the same.
MARK|14|32|They went to a place called Gethsemane, and Jesus said to his disciples, "Sit here while I pray."
MARK|14|33|He took Peter, James and John along with him, and he began to be deeply distressed and troubled.
MARK|14|34|"My soul is overwhelmed with sorrow to the point of death," he said to them. "Stay here and keep watch."
MARK|14|35|Going a little farther, he fell to the ground and prayed that if possible the hour might pass from him.
MARK|14|36|"Abba, Father," he said, "everything is possible for you. Take this cup from me. Yet not what I will, but what you will."
MARK|14|37|Then he returned to his disciples and found them sleeping. "Simon," he said to Peter, "are you asleep? Could you not keep watch for one hour?
MARK|14|38|Watch and pray so that you will not fall into temptation. The spirit is willing, but the body is weak."
MARK|14|39|Once more he went away and prayed the same thing.
MARK|14|40|When he came back, he again found them sleeping, because their eyes were heavy. They did not know what to say to him.
MARK|14|41|Returning the third time, he said to them, "Are you still sleeping and resting? Enough! The hour has come. Look, the Son of Man is betrayed into the hands of sinners.
MARK|14|42|Rise! Let us go! Here comes my betrayer!"
MARK|14|43|Just as he was speaking, Judas, one of the Twelve, appeared. With him was a crowd armed with swords and clubs, sent from the chief priests, the teachers of the law, and the elders.
MARK|14|44|Now the betrayer had arranged a signal with them: "The one I kiss is the man; arrest him and lead him away under guard."
MARK|14|45|Going at once to Jesus, Judas said, "Rabbi!" and kissed him.
MARK|14|46|The men seized Jesus and arrested him.
MARK|14|47|Then one of those standing near drew his sword and struck the servant of the high priest, cutting off his ear.
MARK|14|48|"Am I leading a rebellion," said Jesus, "that you have come out with swords and clubs to capture me?
MARK|14|49|Every day I was with you, teaching in the temple courts, and you did not arrest me. But the Scriptures must be fulfilled."
MARK|14|50|Then everyone deserted him and fled.
MARK|14|51|A young man, wearing nothing but a linen garment, was following Jesus. When they seized him,
MARK|14|52|he fled naked, leaving his garment behind.
MARK|14|53|They took Jesus to the high priest, and all the chief priests, elders and teachers of the law came together.
MARK|14|54|Peter followed him at a distance, right into the courtyard of the high priest. There he sat with the guards and warmed himself at the fire.
MARK|14|55|The chief priests and the whole Sanhedrin were looking for evidence against Jesus so that they could put him to death, but they did not find any.
MARK|14|56|Many testified falsely against him, but their statements did not agree.
MARK|14|57|Then some stood up and gave this false testimony against him:
MARK|14|58|"We heard him say, 'I will destroy this man-made temple and in three days will build another, not made by man.'"
MARK|14|59|Yet even then their testimony did not agree.
MARK|14|60|Then the high priest stood up before them and asked Jesus, "Are you not going to answer? What is this testimony that these men are bringing against you?"
MARK|14|61|But Jesus remained silent and gave no answer. Again the high priest asked him, "Are you the Christ, the Son of the Blessed One?"
MARK|14|62|"I am," said Jesus. "And you will see the Son of Man sitting at the right hand of the Mighty One and coming on the clouds of heaven."
MARK|14|63|The high priest tore his clothes. "Why do we need any more witnesses?" he asked.
MARK|14|64|"You have heard the blasphemy. What do you think?"
MARK|14|65|They all condemned him as worthy of death. Then some began to spit at him; they blindfolded him, struck him with their fists, and said, "Prophesy!" And the guards took him and beat him.
MARK|14|66|While Peter was below in the courtyard, one of the servant girls of the high priest came by.
MARK|14|67|When she saw Peter warming himself, she looked closely at him. "You also were with that Nazarene, Jesus," she said.
MARK|14|68|But he denied it. "I don't know or understand what you're talking about," he said, and went out into the entryway.
MARK|14|69|When the servant girl saw him there, she said again to those standing around, "This fellow is one of them."
MARK|14|70|Again he denied it. After a little while, those standing near said to Peter, "Surely you are one of them, for you are a Galilean."
MARK|14|71|He began to call down curses on himself, and he swore to them, "I don't know this man you're talking about."
MARK|14|72|Immediately the rooster crowed the second time. Then Peter remembered the word Jesus had spoken to him: "Before the rooster crows twice you will disown me three times." And he broke down and wept.
MARK|15|1|Very early in the morning, the chief priests, with the elders, the teachers of the law and the whole Sanhedrin, reached a decision. They bound Jesus, led him away and handed him over to Pilate.
MARK|15|2|"Are you the king of the Jews?" asked Pilate. "Yes, it is as you say," Jesus replied.
MARK|15|3|The chief priests accused him of many things.
MARK|15|4|So again Pilate asked him, "Aren't you going to answer? See how many things they are accusing you of."
MARK|15|5|But Jesus still made no reply, and Pilate was amazed.
MARK|15|6|Now it was the custom at the Feast to release a prisoner whom the people requested.
MARK|15|7|A man called Barabbas was in prison with the insurrectionists who had committed murder in the uprising.
MARK|15|8|The crowd came up and asked Pilate to do for them what he usually did.
MARK|15|9|"Do you want me to release to you the king of the Jews?" asked Pilate,
MARK|15|10|knowing it was out of envy that the chief priests had handed Jesus over to him.
MARK|15|11|But the chief priests stirred up the crowd to have Pilate release Barabbas instead.
MARK|15|12|"What shall I do, then, with the one you call the king of the Jews?" Pilate asked them.
MARK|15|13|"Crucify him!" they shouted.
MARK|15|14|"Why? What crime has he committed?" asked Pilate. But they shouted all the louder, "Crucify him!"
MARK|15|15|Wanting to satisfy the crowd, Pilate released Barabbas to them. He had Jesus flogged, and handed him over to be crucified.
MARK|15|16|The soldiers led Jesus away into the palace (that is, the Praetorium) and called together the whole company of soldiers.
MARK|15|17|They put a purple robe on him, then twisted together a crown of thorns and set it on him.
MARK|15|18|And they began to call out to him, "Hail, king of the Jews!"
MARK|15|19|Again and again they struck him on the head with a staff and spit on him. Falling on their knees, they paid homage to him.
MARK|15|20|And when they had mocked him, they took off the purple robe and put his own clothes on him. Then they led him out to crucify him.
MARK|15|21|A certain man from Cyrene, Simon, the father of Alexander and Rufus, was passing by on his way in from the country, and they forced him to carry the cross.
MARK|15|22|They brought Jesus to the place called Golgotha (which means The Place of the Skull).
MARK|15|23|Then they offered him wine mixed with myrrh, but he did not take it.
MARK|15|24|And they crucified him. Dividing up his clothes, they cast lots to see what each would get.
MARK|15|25|It was the third hour when they crucified him.
MARK|15|26|The written notice of the charge against him read: THE KING OF THE JEWS.
MARK|15|27|They crucified two robbers with him, one on his right and one on his left.
MARK|15|28|See Footnote
MARK|15|29|Those who passed by hurled insults at him, shaking their heads and saying, "So! You who are going to destroy the temple and build it in three days,
MARK|15|30|come down from the cross and save yourself!"
MARK|15|31|In the same way the chief priests and the teachers of the law mocked him among themselves. "He saved others," they said, "but he can't save himself!
MARK|15|32|Let this Christ, this King of Israel, come down now from the cross, that we may see and believe." Those crucified with him also heaped insults on him.
MARK|15|33|At the sixth hour darkness came over the whole land until the ninth hour.
MARK|15|34|And at the ninth hour Jesus cried out in a loud voice, "Eloi, Eloi, lama sabachthani?"--which means, "My God, my God, why have you forsaken me?"
MARK|15|35|When some of those standing near heard this, they said, "Listen, he's calling Elijah."
MARK|15|36|One man ran, filled a sponge with wine vinegar, put it on a stick, and offered it to Jesus to drink. "Now leave him alone. Let's see if Elijah comes to take him down," he said.
MARK|15|37|With a loud cry, Jesus breathed his last.
MARK|15|38|The curtain of the temple was torn in two from top to bottom.
MARK|15|39|And when the centurion, who stood there in front of Jesus, heard his cry and saw how he died, he said, "Surely this man was the Son of God!"
MARK|15|40|Some women were watching from a distance. Among them were Mary Magdalene, Mary the mother of James the younger and of Joses, and Salome.
MARK|15|41|In Galilee these women had followed him and cared for his needs. Many other women who had come up with him to Jerusalem were also there.
MARK|15|42|It was Preparation Day (that is, the day before the Sabbath). So as evening approached,
MARK|15|43|Joseph of Arimathea, a prominent member of the Council, who was himself waiting for the kingdom of God, went boldly to Pilate and asked for Jesus' body.
MARK|15|44|Pilate was surprised to hear that he was already dead. Summoning the centurion, he asked him if Jesus had already died.
MARK|15|45|When he learned from the centurion that it was so, he gave the body to Joseph.
MARK|15|46|So Joseph bought some linen cloth, took down the body, wrapped it in the linen, and placed it in a tomb cut out of rock. Then he rolled a stone against the entrance of the tomb.
MARK|15|47|Mary Magdalene and Mary the mother of Joses saw where he was laid.
MARK|16|1|When the Sabbath was over, Mary Magdalene, Mary the mother of James, and Salome bought spices so that they might go to anoint Jesus' body.
MARK|16|2|Very early on the first day of the week, just after sunrise, they were on their way to the tomb
MARK|16|3|and they asked each other, "Who will roll the stone away from the entrance of the tomb?"
MARK|16|4|But when they looked up, they saw that the stone, which was very large, had been rolled away.
MARK|16|5|As they entered the tomb, they saw a young man dressed in a white robe sitting on the right side, and they were alarmed.
MARK|16|6|"Don't be alarmed," he said. "You are looking for Jesus the Nazarene, who was crucified. He has risen! He is not here. See the place where they laid him.
MARK|16|7|But go, tell his disciples and Peter, 'He is going ahead of you into Galilee. There you will see him, just as he told you.'"
MARK|16|8|Trembling and bewildered, the women went out and fled from the tomb. They said nothing to anyone, because they were afraid.
MARK|16|9|When Jesus rose early on the first day of the week, he appeared first to Mary Magdalene, out of whom he had driven seven demons.
MARK|16|10|She went and told those who had been with him and who were mourning and weeping.
MARK|16|11|When they heard that Jesus was alive and that she had seen him, they did not believe it.
MARK|16|12|Afterward Jesus appeared in a different form to two of them while they were walking in the country.
MARK|16|13|These returned and reported it to the rest; but they did not believe them either.
MARK|16|14|Later Jesus appeared to the Eleven as they were eating; he rebuked them for their lack of faith and their stubborn refusal to believe those who had seen him after he had risen.
MARK|16|15|He said to them, "Go into all the world and preach the good news to all creation.
MARK|16|16|Whoever believes and is baptized will be saved, but whoever does not believe will be condemned.
MARK|16|17|And these signs will accompany those who believe: In my name they will drive out demons; they will speak in new tongues;
MARK|16|18|they will pick up snakes with their hands; and when they drink deadly poison, it will not hurt them at all; they will place their hands on sick people, and they will get well."
MARK|16|19|After the Lord Jesus had spoken to them, he was taken up into heaven and he sat at the right hand of God.
MARK|16|20|Then the disciples went out and preached everywhere, and the Lord worked with them and confirmed his word by the signs that accompanied it.
