NUM|1|1|И сказал Господь Моисею в пустыне Синайской, в скинии собрания, в первый [день] второго месяца, во второй год по выходе их из земли Египетской, говоря:
NUM|1|2|исчислите все общество сынов Израилевых по родам их, по семействам их, по числу имен, всех мужеского пола поголовно:
NUM|1|3|от двадцати лет и выше, всех годных для войны у Израиля, по ополчениям их исчислите их – ты и Аарон;
NUM|1|4|с вами должны быть из каждого колена по одному человеку, который в роде своем есть главный.
NUM|1|5|И вот имена мужей, которые будут с вами: от Рувима Елицур, сын Шедеура;
NUM|1|6|от Симеона Шелумиил, сын Цуришаддая;
NUM|1|7|от Иуды Наассон, сын Аминадава;
NUM|1|8|от Иссахара Нафанаил, сын Цуара;
NUM|1|9|от Завулона Елиав, сын Хелона;
NUM|1|10|от сынов Иосифа: от Ефрема Елишама, сын Аммиуда; от Манассии Гамалиил, сын Педацура;
NUM|1|11|от Вениамина Авидан, сын Гидеония;
NUM|1|12|от Дана Ахиезер, сын Аммишаддая;
NUM|1|13|от Асира Пагиил, сын Охрана;
NUM|1|14|от Гада Елиасаф, сын Регуила;
NUM|1|15|от Неффалима Ахира, сын Енана.
NUM|1|16|Это – избранные мужи общества, начальники колен отцов своих, главы тысяч Израилевых.
NUM|1|17|И взял Моисей и Аарон мужей сих, которые названы поименно,
NUM|1|18|и собрали они все общество в первый [день] второго месяца. И объявили они родословия свои, по родам их, по семействам их, по числу имен, от двадцати лет и выше, поголовно,
NUM|1|19|как повелел Господь Моисею. И сделал он счисление им в пустыне Синайской.
NUM|1|20|И было сынов Рувима, первенца Израилева, по родам их, по племенам их, по семействам их, по числу имен, поголовно, всех мужеского пола, от двадцати лет и выше, всех годных для войны,
NUM|1|21|исчислено в колене Рувимовом сорок шесть тысяч пятьсот.
NUM|1|22|Сынов Симеона по родам их, по племенам их, по семействам их, по числу имен, поголовно, всех мужеского пола, от двадцати лет и выше, всех годных для войны,
NUM|1|23|исчислено в колене Симеоновом пятьдесят девять тысяч триста.
NUM|1|24|Сынов Гада по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|25|исчислено в колене Гадовом сорок пять тысяч шестьсот пятьдесят.
NUM|1|26|Сынов Иуды по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|27|исчислено в колене Иудином семьдесят четыре тысячи шестьсот.
NUM|1|28|Сынов Иссахара по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|29|исчислено в колене Иссахаровом пятьдесят четыре тысячи четыреста.
NUM|1|30|Сынов Завулона по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|31|исчислено в колене Завулоновом пятьдесят семь тысяч четыреста.
NUM|1|32|Сынов Иосифа, сынов Ефрема по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|33|исчислено в колене Ефремовом сорок тысяч пятьсот.
NUM|1|34|Сынов Манассии по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|35|исчислено в колене Манассиином тридцать две тысячи двести.
NUM|1|36|Сынов Вениамина по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|37|исчислено в колене Вениаминовом тридцать пять тысяч четыреста.
NUM|1|38|Сынов Дана по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|39|исчислено в колене Дановом шестьдесят две тысячи семьсот.
NUM|1|40|Сынов Асира по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|41|исчислено в колене Асировом сорок одна тысяча пятьсот.
NUM|1|42|Сынов Неффалима по родам их, по племенам их, по семействам их, по числу имен, от двадцати лет и выше, всех годных для войны,
NUM|1|43|исчислено в колене Неффалимовом пятьдесят три тысячи четыреста.
NUM|1|44|Вот вошедшие в исчисление, которых исчислил Моисей и Аарон и начальники Израиля – двенадцать человек, по одному человеку из каждого племени.
NUM|1|45|И было всех, вошедших в исчисление, сынов Израилевых, по семействам их, от двадцати лет и выше, всех годных для войны у Израиля,
NUM|1|46|и было всех вошедших в исчисление шестьсот три тысячи пятьсот пятьдесят.
NUM|1|47|А левиты по поколениям отцов их не были исчислены между ними.
NUM|1|48|И сказал Господь Моисею, говоря:
NUM|1|49|только колена Левиина не вноси в перепись, и не исчисляй их вместе с сынами Израиля;
NUM|1|50|но поручи левитам скинию откровения и все принадлежности ее и все, что при ней; пусть они носят скинию и все принадлежности ее, и служат при ней, и около скинии пусть ставят стан свой;
NUM|1|51|и когда надобно переносить скинию, пусть поднимают ее левиты, и когда надобно остановиться скинии, пусть ставят ее левиты; а если приступит кто посторонний, предан будет смерти.
NUM|1|52|Сыны Израилевы должны становиться каждый в стане своем и каждый при своем знамени, по ополчениям своим;
NUM|1|53|а левиты должны ставить стан около скинии откровения, чтобы не было гнева на общество сынов Израилевых, и будут левиты стоять на страже у скинии откровения.
NUM|1|54|И сделали сыны Израилевы; как повелел Господь Моисею, так они и сделали.
NUM|2|1|И сказал Господь Моисею и Аарону, говоря:
NUM|2|2|сыны Израилевы должны каждый ставить стан свой при знамени своем, при знаках семейств своих; пред скиниею собрания вокруг должны ставить стан свой.
NUM|2|3|С передней стороны к востоку ставят стан: знамя стана Иудина по ополчениям их, и начальник сынов Иуды Наассон, сын Аминадава,
NUM|2|4|и воинства его, вошедших в исчисление его, семьдесят четыре тысячи шестьсот;
NUM|2|5|после него ставит стан колено Иссахарово, и начальник сынов Иссахара Нафанаил, сын Цуара,
NUM|2|6|и воинства его, вошедших в исчисление его, пятьдесят четыре тысячи четыреста;
NUM|2|7|[далее ставит стан] колено Завулона, и начальник сынов Завулона Елиав, сын Хелона,
NUM|2|8|и воинства его, вошедших в исчисление его, пятьдесят семь тысяч четыреста;
NUM|2|9|всех вошедших в исчисление к стану Иуды сто восемьдесят шесть тысяч четыреста, по ополчениям их; первыми они должны отправляться.
NUM|2|10|Знамя стана Рувимова к югу, по ополчениям их, и начальник сынов Рувимовых Елицур, сын Шедеура,
NUM|2|11|и воинства его, вошедших в исчисление его, сорок шесть тысяч пятьсот;
NUM|2|12|подле него ставит стан колено Симеоново, и начальник сынов Симеона Шелумиил, сын Цуришаддая,
NUM|2|13|и воинства его, вошедших в исчисление его, пятьдесят девять тысяч триста;
NUM|2|14|потом колено Гада, и начальник сынов Гада Елиасаф, сын Регуила,
NUM|2|15|и воинства его, вошедших в исчисление его, сорок пять тысяч шестьсот пятьдесят;
NUM|2|16|всех вошедших в исчисление к стану Рувима сто пятьдесят одна тысяча четыреста пятьдесят, по ополчениям их; вторыми они должны отправляться.
NUM|2|17|Когда пойдет скиния собрания, стан левитов будет в середине станов. Как стоят, так и должны идти, каждый на своем месте при знаменах своих.
NUM|2|18|Знамя стана Ефремова по ополчениям их к западу, и начальник сынов Ефрема Елишама, сын Аммиуда,
NUM|2|19|и воинства его, вошедших в исчисление его, сорок тысяч пятьсот;
NUM|2|20|подле него колено Манассиино, и начальник сынов Манассии Гамалиил, сын Педацура,
NUM|2|21|и воинства его, вошедших в исчисление его, тридцать две тысячи двести;
NUM|2|22|потом колено Вениамина, и начальник сынов Вениамина Авидан, сын Гидеония,
NUM|2|23|и воинства его, вошедших в исчисление его, тридцать пять тысяч четыреста;
NUM|2|24|всех вошедших в исчисление к стану Ефрема сто восемь тысяч сто, по ополчениям их; третьими они должны отправляться.
NUM|2|25|Знамя стана Данова к северу, по ополчениям их, и начальник сынов Дана Ахиезер, сын Аммишаддая,
NUM|2|26|и воинства его, вошедших в исчисление его, шестьдесят две тысячи семьсот;
NUM|2|27|подле него ставит стан колено Асирово, и начальник сынов Асира Пагиил, сын Охрана,
NUM|2|28|и воинства его, вошедших в исчисление его, сорок одна тысяча пятьсот;
NUM|2|29|далее колено Неффалима, и начальник сынов Неффалима Ахира, сын Енана,
NUM|2|30|и воинства его, вошедших в исчисление его, пятьдесят три тысячи четыреста;
NUM|2|31|всех вошедших в исчисление к стану Дана сто пятьдесят семь тысяч шестьсот; они должны идти последними при знаменах своих.
NUM|2|32|Вот вошедшие в исчисление сыны Израиля по семействам их. Всех вошедших в исчисление в станах, по ополчениям их, шестьсот три тысячи пятьсот пятьдесят.
NUM|2|33|А левиты не вошли в исчисление вместе с сынами Израиля, как повелел Господь Моисею.
NUM|2|34|И сделали сыны Израилевы все, что повелел Господь Моисею: так становились станами при знаменах своих и так шли каждый по племенам своим, по семействам своим.
NUM|3|1|Вот родословие Аарона и Моисея, когда говорил Господь Моисею на горе Синае,
NUM|3|2|и вот имена сынов Аарона: первенец Надав, Авиуд, Елеазар и Ифамар;
NUM|3|3|это имена сынов Аарона, священников, помазанных, которых он посвятил, чтобы священнодействовать;
NUM|3|4|но Надав и Авиуд умерли пред лицем Господа, когда они принесли огонь чуждый пред лице Господа в пустыне Синайской, детей же у них не было; и остались священниками Елеазар и Ифамар при Аароне, отце своем.
NUM|3|5|И сказал Господь Моисею, говоря:
NUM|3|6|приведи колено Левиино, и поставь его пред Аароном священником, чтоб они служили ему;
NUM|3|7|и пусть они будут на страже за него и на страже за все общество при скинии собрания, чтобы отправлять службы при скинии;
NUM|3|8|и пусть хранят все вещи скинии собрания, и будут на страже за сынов Израилевых, чтобы отправлять службы при скинии;
NUM|3|9|отдай левитов Аарону и сынам его [в] [распоряжение]: да будут они отданы ему из сынов Израилевых;
NUM|3|10|Аарону же и сынам его поручи, чтобы они наблюдали священническую должность свою; а если приступит кто посторонний, предан будет смерти.
NUM|3|11|И сказал Господь Моисею, говоря:
NUM|3|12|вот, Я взял левитов из сынов Израилевых вместо всех первенцев, разверзающих ложесна из сынов Израилевых; левиты должны быть Мои,
NUM|3|13|ибо все первенцы – Мои; в тот день, когда поразил Я всех первенцев в земле Египетской, освятил Я Себе всех первенцев Израилевых от человека до скота; они должны быть Мои. Я Господь.
NUM|3|14|И сказал Господь Моисею в пустыне Синайской, говоря:
NUM|3|15|исчисли сынов Левииных по семействам их, по родам их; всех мужеского пола от одного месяца и выше исчисли.
NUM|3|16|И исчислил их Моисей по слову Господню, как повелено.
NUM|3|17|И вот сыны Левиины по именам их: Гирсон, Кааф и Мерари.
NUM|3|18|И вот имена сынов Гирсоновых по родам их: Ливни и Шимей.
NUM|3|19|И сыны Каафа по родам их: Амрам и Ицгар, Хеврон и Узиил.
NUM|3|20|И сыны Мерари по родам их: Махли и Муши. Вот роды Левиины по семействам их.
NUM|3|21|От Гирсона род Ливни и род Шимея: это роды Гирсоновы.
NUM|3|22|Исчисленных было всех мужеского пола, от одного месяца и выше, семь тысяч пятьсот.
NUM|3|23|Роды Гирсоновы должны становиться станом позади скинии на запад;
NUM|3|24|начальник поколения сынов Гирсоновых Елиасаф, сын Лаелов;
NUM|3|25|хранению сынов Гирсоновых в скинии собрания поручается скиния и покров ее, и завеса входа скинии собрания,
NUM|3|26|и завесы двора и завеса входа двора, который вокруг скинии и жертвенника, и веревки ее, со всеми их принадлежностями.
NUM|3|27|От Каафа род Амрама и род Ицгара, и род Хеврона, и род Узиила: это роды Каафа.
NUM|3|28|По счету всех мужеского пола, от одного месяца и выше, восемь тысяч шестьсот, которые охраняли святилище.
NUM|3|29|Роды сынов Каафовых должны ставить стан свой на южной стороне скинии;
NUM|3|30|начальник же поколения родов Каафовых Елцафан, сын Узиила;
NUM|3|31|в хранении у них ковчег, стол, светильник, жертвенники, священные сосуды, которые употребляются при служении, и завеса со всеми принадлежностями ее.
NUM|3|32|Начальник над начальниками левитов Елеазар, сын Аарона священника; под его надзором те, которым вверено хранение святилища.
NUM|3|33|От Мерари род Махли и род Муши: это роды Мерари;
NUM|3|34|исчисленных по числу всех мужеского пола, от одного месяца и выше – шесть тысяч двести;
NUM|3|35|начальник поколения родов Мерари Цуриил, сын Авихаила; они должны ставить стан свой на северной стороне скинии;
NUM|3|36|хранению сынов Мерари поручаются брусья скинии и шесты ее, и столбы ее, и подножия ее и все вещи ее, со всем устройством их,
NUM|3|37|и столбы двора со всех сторон и подножия их и колья их и веревки их.
NUM|3|38|А с передней стороны скинии, к востоку пред скиниею собрания, должны ставить стан Моисей и Аарон и сыны его, которым вверено хранение святилища за сынов Израилевых; а если приступит кто посторонний, предан будет смерти.
NUM|3|39|Всех исчисленных левитов, которых исчислил Моисей и Аарон по повелению Господню, по родам их, всех мужеского пола, от одного месяца и выше, двадцать две тысячи.
NUM|3|40|И сказал Господь Моисею: исчисли всех первенцев мужеского пола из сынов Израилевых, от одного месяца и выше, и пересчитай их поименно;
NUM|3|41|и возьми левитов для Меня, – Я Господь, – вместо всех первенцев из сынов Израиля, а скот левитов вместо всего первородного скота сынов Израилевых.
NUM|3|42|И исчислил Моисей, как повелел ему Господь, всех первенцев из сынов Израилевых
NUM|3|43|и было всех первенцев мужеского пола, по числу имен, от одного месяца и выше, двадцать две тысячи двести семьдесят три.
NUM|3|44|И сказал Господь Моисею, говоря:
NUM|3|45|возьми левитов вместо всех первенцев из сынов Израиля и скот левитов вместо скота их; пусть левиты будут Мои. Я Господь.
NUM|3|46|А в выкуп двухсот семидесяти трех, которые лишние против [числа] левитов, из первенцев Израильских,
NUM|3|47|возьми по пяти сиклей за человека, по сиклю священному возьми, двадцать гер в сикле,
NUM|3|48|и отдай серебро сие Аарону и сынам его, в выкуп за излишних против [числа] их.
NUM|3|49|И взял Моисей серебро выкупа за излишних против [числа] замененных левитами,
NUM|3|50|от первенцев Израилевых взял серебра тысячу триста шестьдесят пять [сиклей], по сиклю священному,
NUM|3|51|и отдал Моисей серебро выкупа Аарону и сынам его по слову Господню, как повелел Господь Моисею.
NUM|4|1|И сказал Господь Моисею и Аарону, говоря:
NUM|4|2|исчисли сынов Каафовых из сынов Левия по родам их, по семействам их,
NUM|4|3|от тридцати лет и выше до пятидесяти лет, всех способных к службе, чтобы отправлять работы в скинии собрания.
NUM|4|4|Вот служение сынов Каафовых в скинии собрания: [носить] Святое Святых.
NUM|4|5|Когда стану надобно подняться в путь, Аарон и сыны его войдут, и снимут завесу закрывающую, и покроют ею ковчег откровения;
NUM|4|6|и положат на нее покров из кож синего цвета, и сверх его накинут покрывало все из голубой [шерсти], и вложат шесты его;
NUM|4|7|и стол [хлебов] предложения накроют одеждою из голубой [шерсти], и поставят на нем блюда, тарелки, чаши и кружки для возлияния, и хлеб [его] всегдашний должен быть на нем;
NUM|4|8|и возложат на них одежду багряную, и покроют ее покровом из кожи синего цвета, и вложат шесты его;
NUM|4|9|и возьмут одежду из голубой [шерсти], и покроют светильник и лампады его, и щипцы его, и лотки его, и все сосуды для елея, которые употребляют при нем,
NUM|4|10|и покроют его и все принадлежности его покровом из кож синих, и положат на носилки;
NUM|4|11|и на золотой жертвенник возложат одежду из голубой [шерсти], и покроют его покровом из кож синих, и вложат шесты его.
NUM|4|12|И возьмут все вещи служебные, которые употребляются для служения во святилище, и положат в одежду из голубой [шерсти], и покроют их покровом из кож синих, и положат на носилки.
NUM|4|13|И очистят жертвенник от пепла и накроют его одеждою пурпуровою;
NUM|4|14|и положат на него все сосуды его, которые употребляются для служения при нем – угольницы, вилки, лопатки и чаши, все сосуды жертвенника – и покроют его покровом из кож синих, и вложат шесты его.
NUM|4|15|Когда, при отправлении в путь стана, Аарон и сыны его покроют все святилище и все вещи святилища, тогда сыны Каафа подойдут, чтобы нести; но не должны они касаться святилища, чтобы не умереть. Сии [части] скинии собрания должны носить сыны Каафовы.
NUM|4|16|Елеазару, сыну Аарона священника, поручается елей для светильника и благовонное курение, и всегдашнее хлебное приношение и елей помазания, – поручается вся скиния и все, что в ней, святилище и принадлежности его.
NUM|4|17|И сказал Господь Моисею и Аарону, говоря:
NUM|4|18|не погубите колена племен Каафовых из среды левитов,
NUM|4|19|но вот что сделайте им, чтобы они были живы и не умерли, когда приступают к Святому Святых: Аарон и сыны его пусть придут и поставят их каждого в служении его и у ноши его;
NUM|4|20|но сами они не должны подходить смотреть святыню, когда покрывают ее, чтобы не умереть.
NUM|4|21|И сказал Господь Моисею, говоря:
NUM|4|22|исчисли и сынов Гирсона по семействам их, по родам их,
NUM|4|23|от тридцати лет и выше до пятидесяти лет, исчисли их всех способных к службе, чтобы отправлять работы при скинии собрания.
NUM|4|24|Вот работы семейств Гирсоновых, при их служении и ношении тяжестей:
NUM|4|25|они должны носить покровы скинии и скинию собрания, и покров ее, и покров кожаный синий, который поверх его, и завесу входа скинии собрания,
NUM|4|26|и завесы двора, и завесу входа во двор, который вокруг скинии и жертвенника, и веревки их, и все вещи, принадлежащие к ним; и все, что делается при них, они должны работать;
NUM|4|27|по повелению Аарона и сынов его должны производиться все службы сынов Гирсоновых при всяком ношении тяжестей и всякой работе их, и поручите их хранению все, что они носят;
NUM|4|28|вот службы родов сынов Гирсоновых в скинии собрания, и вот что поручается их хранению под надзором Ифамара, сына Аарона, священника.
NUM|4|29|Сынов Мерариных по родам их, по семействам их исчисли,
NUM|4|30|от тридцати лет и выше до пятидесяти лет, исчисли всех способных на службу, чтобы отправлять работы при скинии собрания.
NUM|4|31|Вот что они должны носить, по службе их при скинии собрания: брусья скинии и шесты ее, и столбы ее и подножия ее,
NUM|4|32|и столбы двора со всех сторон и подножия их, и колья их, и веревки их, и все вещи при них и все принадлежности их; и поименно сосчитайте вещи, которые они обязаны носить;
NUM|4|33|Вот работы родов сынов Мерариных, по службе их при скинии собрания, под надзором Ифамара, сына Аарона, священника.
NUM|4|34|И исчислили Моисей и Аарон и начальники общества сынов Каафовых по родам их и по семействам их,
NUM|4|35|от тридцати лет и выше до пятидесяти лет, всех способных к службе, для работ в скинии собрания;
NUM|4|36|и было исчислено, по родам их, две тысячи семьсот пятьдесят:
NUM|4|37|это – исчисленные из родов Каафовых, все служащие при скинии собрания, которых исчислил Моисей и Аарон по повелению Господню, [данному] чрез Моисея.
NUM|4|38|И исчислены сыны Гирсона по родам их и по семействам их,
NUM|4|39|от тридцати лет и выше до пятидесяти лет, все способные к службе, для работ в скинии собрания;
NUM|4|40|и было исчислено по родам их, по семействам их, две тысячи шестьсот тридцать:
NUM|4|41|это – исчисленные из родов сынов Гирсона, все служащие при скинии собрания, которых исчислил Моисей и Аарон, по повелению Господню.
NUM|4|42|И исчислены роды сынов Мерариных по родам их, по семействам их,
NUM|4|43|от тридцати лет и выше до пятидесяти лет, все способные к службе, для работ при скинии собрания;
NUM|4|44|и было исчислено по родам их, три тысячи двести:
NUM|4|45|это – исчисленные из родов сынов Мерариных, которых исчислил Моисей и Аарон по повелению Господню, [данному] чрез Моисея.
NUM|4|46|И исчислены все левиты, которых исчислил Моисей и Аарон и начальники Израиля по родам их и по семействам их,
NUM|4|47|от тридцати лет и выше до пятидесяти лет, все способные [к] [службе] для работ и ношения в скинии собрания;
NUM|4|48|и было исчислено их восемь тысяч пятьсот восемьдесят;
NUM|4|49|по повелению Господню чрез Моисея определены они каждый к своей работе и ношению, и исчислены, как повелел Господь Моисею.
NUM|5|1|И сказал Господь Моисею, говоря:
NUM|5|2|повели сынам Израилевым выслать из стана всех прокаженных, и всех имеющих истечение, и всех осквернившихся от мертвого,
NUM|5|3|и мужчин и женщин вышлите, за стан вышлите их, чтобы не оскверняли они станов своих, среди которых Я живу.
NUM|5|4|И сделали так сыны Израилевы, и выслали их вон из стана; как говорил Господь Моисею, так и сделали сыны Израилевы.
NUM|5|5|И сказал Господь Моисею, говоря:
NUM|5|6|скажи сынам Израилевым: если мужчина или женщина сделает какой–либо грех против человека, и чрез это сделает преступление против Господа, и виновна будет душа та,
NUM|5|7|то пусть исповедаются во грехе своем, который они сделали, и возвратят сполна то, в чем виновны, и прибавят к тому пятую часть и отдадут тому, против кого согрешили;
NUM|5|8|если же у него нет наследника, которому следовало бы возвратить за вину: то посвятить это Господу; пусть будет это священнику, сверх овна очищения, которым он очистит его;
NUM|5|9|и всякое возношение из всех святынь сынов Израилевых, которые они приносят к священнику, ему принадлежит,
NUM|5|10|и посвященное кем–либо ему принадлежит; все, что даст кто священнику, ему принадлежит.
NUM|5|11|И сказал Господь Моисею, говоря:
NUM|5|12|объяви сынам Израилевым и скажи им: если изменит кому жена, и нарушит верность к нему,
NUM|5|13|и переспит кто с ней и излиет семя, и это будет скрыто от глаз мужа ее, и она осквернится тайно, и не будет на нее свидетеля, и не будет уличена,
NUM|5|14|и найдет на него дух ревности, и будет ревновать жену свою, когда она осквернена, или найдет на него дух ревности, и он будет ревновать жену свою, когда она не осквернена, –
NUM|5|15|пусть приведет муж жену свою к священнику и принесет за нее в жертву десятую часть ефы ячменной муки, но не возливает на нее елея и не кладет ливана, потому что это приношение ревнования, приношение воспоминания, напоминающее о беззаконии;
NUM|5|16|а священник пусть приведет и поставит ее пред лице Господне,
NUM|5|17|и возьмет священник святой воды в глиняный сосуд, и возьмет священник земли с полу скинии и положит в воду;
NUM|5|18|и поставит священник жену пред лице Господне, и обнажит голову жены, и даст ей в руки приношение воспоминания, – это приношение ревнования, в руке же у священника будет горькая вода, наводящая проклятие.
NUM|5|19|И заклянет ее священник и скажет жене: если никто не переспал с тобою, и ты не осквернилась и не изменила мужу своему, то невредима будешь от сей горькой воды, наводящей проклятие;
NUM|5|20|но если ты изменила мужу твоему и осквернилась, и если кто переспал с тобою кроме мужа твоего, –
NUM|5|21|тогда священник пусть заклянет жену клятвою проклятия и скажет священник жене: да предаст тебя Господь проклятию и клятве в народе твоем, и да соделает Господь лоно твое опавшим и живот твой опухшим;
NUM|5|22|и да пройдет вода сия, наводящая проклятие, во внутренность твою, чтобы опух живот [твой] и опало лоно [твое]. И скажет жена: аминь, аминь.
NUM|5|23|И напишет священник заклинания сии на свитке, и смоет их в горькую воду;
NUM|5|24|и даст жене выпить горькую воду, наводящую проклятие, и войдет в нее вода, наводящая проклятие, ко вреду ее.
NUM|5|25|И возьмет священник из рук жены хлебное приношение ревнования, и вознесет сие приношение пред Господом, и отнесет его к жертвеннику;
NUM|5|26|и возьмет священник горстью из хлебного приношения часть в память, и сожжет на жертвеннике, и потом даст жене выпить воды;
NUM|5|27|и когда напоит ее водою, тогда, если она нечиста и сделала преступление против мужа своего, горькая вода, наводящая проклятие, войдет в нее, ко вреду ее, и опухнет чрево ее и опадет лоно ее, и будет эта жена проклятою в народе своем;
NUM|5|28|если же жена не осквернилась и была чиста, то останется невредимою и будет оплодотворяема семенем.
NUM|5|29|Вот закон о ревновании, когда жена изменит мужу своему и осквернится,
NUM|5|30|или когда на мужа найдет дух ревности, и он будет ревновать жену свою, тогда пусть он поставит жену пред лицем Господа, и сделает с нею священник все по сему закону, –
NUM|5|31|и будет муж чист от греха, а жена понесет на себе грех свой.
NUM|6|1|И сказал Господь Моисею, говоря:
NUM|6|2|объяви сынам Израилевым и скажи им: если мужчина или женщина решится дать обет назорейства, чтобы посвятить себя в назореи Господу,
NUM|6|3|то он должен воздержаться от вина и [крепкого] напитка, и не должен употреблять ни уксусу из вина, ни уксусу из напитка, и ничего приготовленного из винограда не должен пить, и не должен есть ни сырых, ни сушеных виноградных ягод;
NUM|6|4|во все дни назорейства своего не должен он есть ничего, что делается из винограда, от зерен до кожи.
NUM|6|5|Во все дни обета назорейства его бритва не должна касаться головы его; до исполнения дней, на которые он посвятил себя в назореи Господу, свят он: должен растить волосы на голове своей.
NUM|6|6|Во все дни, на которые он посвятил себя в назореи Господу, не должен он подходить к мертвому телу:
NUM|6|7|[прикосновением] к отцу своему, и матери своей, и брату своему, и сестре своей, не должен он оскверняться, когда они умрут, потому что посвящение Богу его на главе его;
NUM|6|8|во все дни назорейства своего свят он Господу.
NUM|6|9|Если же умрет при нем кто–нибудь вдруг, нечаянно, и он осквернит тем голову назорейства своего: то он должен остричь голову свою в день очищения его, в седьмой день должен остричь ее,
NUM|6|10|и в восьмой день должен принести двух горлиц, или двух молодых голубей, к священнику, ко входу скинии собрания;
NUM|6|11|священник одну [из птиц] принесет в жертву за грех, а другую во всесожжение, и очистит его от осквернения мертвым телом, и освятит голову его в тот день;
NUM|6|12|и должен он снова начать посвященные Господу дни назорейства своего и принести однолетнего агнца в жертву повинности; прежние же дни пропали, потому что назорейство его осквернено.
NUM|6|13|И вот закон о назорее, когда исполнятся дни назорейства его: должно привести его ко входу скинии собрания,
NUM|6|14|и он принесет в жертву Господу одного однолетнего агнца без порока во всесожжение, и одну однолетнюю агницу без порока в жертву за грех, и одного овна без порока в жертву мирную,
NUM|6|15|и корзину опресноков из пшеничной муки, хлебов, испеченных с елеем, и пресных лепешек, помазанных елеем, и при них хлебное приношение и возлияние;
NUM|6|16|и представит [сие] священник пред Господа, и принесет жертву его за грех и всесожжение его;
NUM|6|17|овна принесет в жертву мирную Господу с корзиною опресноков, также совершит священник хлебное приношение его и возлияние его;
NUM|6|18|и острижет назорей у входа скинии собрания голову назорейства своего, и возьмет волосы головы назорейства своего, и положит на огонь, который под мирною жертвою;
NUM|6|19|и возьмет священник сваренное плечо овна и один пресный пирог из корзины и одну пресную лепешку, и положит на руки назорею, после того, как острижет он голову назорейства своего;
NUM|6|20|и вознесет сие священник, потрясая пред Господом: эта святыня – для священника, сверх груди потрясания и сверх плеча возношения. После сего назорей может пить вино.
NUM|6|21|Вот закон о назорее, который дал обет, и жертва его Господу за назорейство свое, кроме того, что позволит ему достаток его; по обету своему, какой он даст, так и должен он делать, сверх узаконенного о назорействе его.
NUM|6|22|И сказал Господь Моисею, говоря:
NUM|6|23|скажи Аарону и сынам его: так благословляйте сынов Израилевых, говоря им:
NUM|6|24|да благословит тебя Господь и сохранит тебя!
NUM|6|25|да призрит на тебя Господь светлым лицем Своим и помилует тебя!
NUM|6|26|да обратит Господь лице Свое на тебя и даст тебе мир!
NUM|6|27|Так пусть призывают имя Мое на сынов Израилевых, и Я благословлю их.
NUM|7|1|Когда Моисей поставил скинию, и помазал ее, и освятил ее и все принадлежности ее, и жертвенник и все принадлежности его, и помазал их и освятил их,
NUM|7|2|тогда пришли начальников Израилевых, главы семейств их, начальники колен, заведывавшие исчислением,
NUM|7|3|и представили приношение свое пред Господа, шесть крытых повозок и двенадцать волов, по одной повозке от двух начальников и по одному волу от каждого, и представили сие пред скинию.
NUM|7|4|И сказал Господь Моисею, говоря:
NUM|7|5|возьми от них; это будет для отправления работ при скинии собрания; и отдай это левитам, смотря по роду службы их.
NUM|7|6|И взял Моисей повозки и волов, и отдал их левитам:
NUM|7|7|две повозки и четырех волов отдал сынам Гирсоновым, по роду служб их:
NUM|7|8|и четыре повозки и восемь волов отдал сынам Мерариным, по роду служб их, под надзором Ифамара, сына Аарона, священника;
NUM|7|9|а сынам Каафовым не дал, потому что служба их – [носить] святилище; на плечах они должны носить.
NUM|7|10|И принесли начальники жертвы освящения жертвенника в день помазания его, и представили начальники приношение свое пред жертвенник.
NUM|7|11|И сказал Господь Моисею: по одному начальнику в день пусть приносят приношение свое для освящения жертвенника.
NUM|7|12|В первый день принес приношение свое Наассон, сын Аминадавов, от колена Иудина;
NUM|7|13|приношение его было: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|14|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|15|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|16|один козел в жертву за грех,
NUM|7|17|и в жертву мирную два вола, пять овнов, пять козлов, пять однолетних агнцев; вот приношение Наассона, сына Аминадавова.
NUM|7|18|Во второй день принес Нафанаил, сын Цуара, начальник [колена] Иссахарова;
NUM|7|19|он принес от себя приношение: одно серебряное блюдо, весом в сто тридцать [сиклей], одну серебряную чашу в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|20|одну золотую кадильницу в десять [сиклей], наполненную курением,
NUM|7|21|одного тельца, одного овна, одного однолетнего агнца, во всесожжение,
NUM|7|22|одного козла в жертву за грех,
NUM|7|23|и в жертву мирную двух волов, пять овнов, пять козлов, пять однолетних агнцев; вот приношение Нафанаила, сына Цуарова.
NUM|7|24|В третий день начальник сынов Завулоновых Елиав, сын Хелона;
NUM|7|25|приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|26|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|27|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|28|один козел в жертву за грех,
NUM|7|29|и в жертву мирную два вола, пять овнов, пять козлов, пять однолетних агнцев; вот приношение Елиава, сына Хелонова.
NUM|7|30|В четвертый день начальник сынов Рувимовых Елицур, сын Шедеуров;
NUM|7|31|приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|32|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|33|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|34|один козел в жертву за грех,
NUM|7|35|и в жертву мирную два вола, пять овнов, пять козлов и пять однолетних агнцев; вот приношение Елицура, сына Шедеурова.
NUM|7|36|В пятый день начальник сынов Симеоновых Шелумиил, сын Цуришаддая;
NUM|7|37|приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|38|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|39|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|40|один козел в жертву за грех,
NUM|7|41|и в жертву мирную два вола, пять овнов, пять козлов и пять однолетних агнцев; вот приношение Шелумиила, сына Цуришаддаева.
NUM|7|42|В шестой день начальник сынов Гадовых Елиасаф, сын Регуила;
NUM|7|43|приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|44|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|45|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|46|один козел в жертву за грех,
NUM|7|47|и в жертву мирную два вола, пять овнов, пять козлов и пять однолетних агнцев; вот приношение Елиасафа, сына Регуилова.
NUM|7|48|В седьмой день начальник сынов Ефремовых Елишама, сын Аммиуда.
NUM|7|49|Приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|50|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|51|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|52|один козел в жертву за грех,
NUM|7|53|и в жертву мирную два вола, пять овнов, пять козлов, пять однолетних агнцев; вот приношение Елишамы, сына Аммиудова.
NUM|7|54|В восьмой день начальник сынов Манассииных Гамалиил, сын Педацура.
NUM|7|55|Приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|56|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|57|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|58|один козел в жертву за грех,
NUM|7|59|и в жертву мирную два вола, пять овнов, пять козлов, пять однолетних агнцев; вот приношение Гамалиила, сына Педацурова.
NUM|7|60|В девятый день начальник сынов Вениаминовых Авидан, сын Гидеония;
NUM|7|61|приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|62|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|63|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|64|один козел в жертву за грех,
NUM|7|65|и в жертву мирную два вола, пять овнов, пять козлов, пять однолетних агнцев; вот приношение Авидана, сына Гидеониева.
NUM|7|66|В десятый день начальник сынов Дановых Ахиезер, сын Аммишаддая;
NUM|7|67|приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|68|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|69|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|70|один козел в жертву за грех,
NUM|7|71|и в жертву мирную два вола, пять овнов, пять козлов, пять однолетних агнцев; вот приношение Ахиезера, сына Аммишаддаева.
NUM|7|72|В одиннадцатый день начальник сынов Асировых Пагиил, сын Охрана;
NUM|7|73|приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|74|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|75|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|76|один козел в жертву за грех,
NUM|7|77|и в жертву мирную два вола, пять овнов, пять козлов, пять однолетних агнцев; вот приношение Пагиила, сына Охранова.
NUM|7|78|В двенадцатый день начальник сынов Неффалимовых Ахира, сын Енана;
NUM|7|79|приношение его: одно серебряное блюдо, весом в сто тридцать [сиклей], одна серебряная чаша в семьдесят сиклей, по сиклю священному, наполненные пшеничною мукою, смешанною с елеем, в приношение хлебное,
NUM|7|80|одна золотая кадильница в десять [сиклей], наполненная курением,
NUM|7|81|один телец, один овен, один однолетний агнец, во всесожжение,
NUM|7|82|один козел в жертву за грех,
NUM|7|83|и в жертву мирную два вола, пять овнов, пять козлов, пять однолетних агнцев; вот приношение Ахиры, сына Енанова.
NUM|7|84|Вот [приношения] от начальников Израилевых при освящении жертвенника в день помазания его: двенадцать серебряных блюд, двенадцать серебряных чаш, двенадцать золотых кадильниц;
NUM|7|85|по сто тридцати [сиклей] серебра в каждом блюде и по семидесяти в каждой чаше: итак всего серебра в сих сосудах две тысячи четыреста [сиклей], по сиклю священному;
NUM|7|86|золотых кадильниц, наполненных курением, двенадцать, в каждой кадильнице по десяти [сиклей], по сиклю священному: всего золота в кадильницах сто двадцать [сиклей];
NUM|7|87|во всесожжение всего двенадцать тельцов из скота крупного, двенадцать овнов, двенадцать однолетних агнцев и при них хлебное приношение, и в жертву за грех двенадцать козлов,
NUM|7|88|и в жертву мирную всего из крупного скота двадцать четыре тельца, шестьдесят овнов, шестьдесят козлов, шестьдесят однолетних агнцев. вот приношения при освящении жертвенника после помазания его.
NUM|7|89|Когда Моисей входил в скинию собрания, чтобы говорить с Господом, слышал голос, говорящий ему с крышки, которая над ковчегом откровения между двух херувимов, и он говорил ему.
NUM|8|1|И сказал Господь Моисею, говоря:
NUM|8|2|объяви Аарону и скажи ему: когда ты будешь зажигать лампады, то на передней стороне светильника должны гореть семь лампад.
NUM|8|3|Аарон так и сделал: на передней стороне светильника зажег лампады его, как повелел Господь Моисею.
NUM|8|4|И вот устройство светильника: чеканный он из золота, от стебля его и до цветов чеканный; по образу, который показал Господь Моисею, он сделал светильник.
NUM|8|5|И сказал Господь Моисею, говоря:
NUM|8|6|возьми левитов из среды сынов Израилевых и очисти их;
NUM|8|7|а чтобы очистить их, поступи с ними так: окропи их очистительною водою, и пусть они обреют бритвою все тело свое и вымоют одежды свои, и будут чисты;
NUM|8|8|и пусть возьмут тельца и хлебное приношение к нему, пшеничной муки, смешанной с елеем, и другого тельца возьми в жертву за грех;
NUM|8|9|и приведи левитов пред скинию собрания; и собери все общество сынов Израилевых
NUM|8|10|и приведи левитов их пред Господа, и пусть возложат сыны Израилевы руки свои на левитов;
NUM|8|11|Аарон же пусть совершит над левитами посвящение их пред Господом от сынов Израилевых, чтобы отправляли они служение Господу;
NUM|8|12|а левиты пусть возложат руки свои на голову тельцов, и принеси одного в жертву за грех, а другого во всесожжение Господу, для очищения левитов;
NUM|8|13|и поставь левитов пред Аароном и пред сынами его, и соверши над ними посвящение их Господу;
NUM|8|14|и так отдели левитов от сынов Израилевых, чтобы левиты были Моими.
NUM|8|15|После сего войдут левиты служить скинии собрания, когда ты очистишь их и совершишь над ними посвящение их; ибо они отданы Мне из сынов Израилевых:
NUM|8|16|вместо всех первенцев из сынов Израилевых, разверзающих всякие ложесна, Я беру их Себе;
NUM|8|17|ибо Мои все первенцы у сынов Израилевых, от человека до скота: в тот день, когда Я поразил всех первенцев в земле Египетской, Я освятил их Себе
NUM|8|18|и взял левитов вместо всех первенцев у сынов Израилевых;
NUM|8|19|и отдал левитов Аарону и сынам его из среды сынов Израилевых, чтобы они отправляли службы за сынов Израилевых при скинии собрания и служили охранением для сынов Израилевых, чтобы не постигло сынов Израилевых поражение, когда бы сыны Израилевы приступили к святилищу.
NUM|8|20|И сделали так Моисей и Аарон и все общество сынов Израилевых с левитами: как повелел Господь Моисею о левитах, так и сделали с ними сыны Израилевы.
NUM|8|21|И очистились левиты и омыли одежды свои, и совершил над ними Аарон посвящение их пред Господом, и очистил их Аарон, чтобы сделать их чистыми;
NUM|8|22|после сего вошли левиты отправлять службы свои в скинии собрания пред Аароном и пред сынами его. Как повелел Господь Моисею о левитах, так и сделали они с ними.
NUM|8|23|И сказал Господь Моисею, говоря:
NUM|8|24|вот [закон] о левитах: от двадцати пяти лет и выше должны вступать они в службу для работ при скинии собрания,
NUM|8|25|а в пятьдесят лет должны прекращать отправление работ и более не работать:
NUM|8|26|тогда пусть помогают они братьям своим содержать стражу при скинии собрания, работать же – пусть не работают; так поступай с левитами касательно служения их.
NUM|9|1|И сказал Господь Моисею в пустыне Синайской во второй год по исшествии их из земли Египетской, в первый месяц, говоря:
NUM|9|2|пусть сыны Израилевы совершат Пасху в назначенное для нее время:
NUM|9|3|в четырнадцатый день сего месяца вечером совершите ее в назначенное для нее время, по всем постановлениям и по всем обрядам ее совершите ее.
NUM|9|4|И сказал Моисей сынам Израилевым, чтобы совершили Пасху.
NUM|9|5|И совершили они Пасху в первый [месяц], в четырнадцатый день месяца вечером, в пустыне Синайской: во всем, как повелел Господь Моисею, так и поступили сыны Израилевы.
NUM|9|6|Были люди, которые были нечисты от [прикосновения] к мертвым телам человеческим, и не могли совершить Пасхи в тот день; и пришли они к Моисею и Аарону в тот день,
NUM|9|7|и сказали ему те люди: мы нечисты от [прикосновения] к мертвым телам человеческим; для чего нас лишать того, чтобы мы принесли приношение Господу в назначенное время среди сынов Израилевых?
NUM|9|8|И сказал им Моисей: постойте, я послушаю, что повелит о вас Господь.
NUM|9|9|И сказал Господь Моисею, говоря:
NUM|9|10|скажи сынам Израилевым: если кто из вас или из потомков ваших будет нечист от [прикосновения] к мертвому телу, или будет в дальней дороге, то и он должен совершить Пасху Господню;
NUM|9|11|в четырнадцатый день второго месяца вечером пусть таковые совершат ее и с опресноками и горькими травами пусть едят ее;
NUM|9|12|и пусть не оставляют от нее до утра и костей ее не сокрушают; пусть совершат ее по всем уставам о Пасхе;
NUM|9|13|а кто чист и не находится в дороге и не совершит Пасхи, – истребится душа та из народа своего, ибо он не принес приношения Господу в свое время: понесет на себе грех человек тот;
NUM|9|14|если будет жить у вас пришелец, то и он должен совершать Пасху Господню: по уставу о Пасхе и по обряду ее он должен совершить ее; один устав пусть будет у вас и для пришельца и для туземца.
NUM|9|15|В тот день, когда поставлена была скиния, облако покрыло скинию откровения, и с вечера над скиниею как бы огонь виден был до самого утра.
NUM|9|16|Так было и всегда: облако покрывало ее [днем] и подобие огня ночью.
NUM|9|17|И когда облако поднималось от скинии, тогда сыны Израилевы отправлялись в путь, и на месте, где останавливалось облако, там останавливались станом сыны Израилевы.
NUM|9|18|По повелению Господню отправлялись сыны Израилевы в путь, и по повелению Господню останавливались: во все то время, когда облако стояло над скиниею, и они стояли;
NUM|9|19|и если облако долгое время было над скиниею, то и сыны Израилевы следовали этому указанию Господа и не отправлялись;
NUM|9|20|иногда же облако немного времени было над скиниею: они по указанию Господню останавливались, и по указанию Господню отправлялись в путь;
NUM|9|21|иногда облако стояло [только] от вечера до утра, и поутру поднималось облако, тогда и они отправлялись; или день и ночь стояло облако, и когда поднималось, и они тогда отправлялись;
NUM|9|22|или, если два дня, или месяц, или несколько дней стояло облако над скиниею, то и сыны Израилевы стояли и не отправлялись в путь; а когда оно поднималось, тогда отправлялись;
NUM|9|23|по указанию Господню останавливались, и по указанию Господню отправлялись в путь: следовали указанию Господню по повелению Господню, [данному] чрез Моисея.
NUM|10|1|И сказал Господь Моисею, говоря:
NUM|10|2|сделай себе две серебряные трубы, чеканные сделай их, чтобы они служили тебе для созывания общества и для снятия станов;
NUM|10|3|когда затрубят ими, соберется к тебе все общество ко входу скинии собрания;
NUM|10|4|когда одною трубою затрубят, соберутся к тебе князья и тысяченачальники Израилевы;
NUM|10|5|когда затрубите тревогу, поднимутся станы, становящиеся к востоку;
NUM|10|6|когда во второй раз затрубите тревогу, поднимутся станы, становящиеся к югу; тревогу пусть трубят при отправлении их в путь;
NUM|10|7|а когда надобно собрать собрание, трубите, но не тревогу;
NUM|10|8|сыны Аароновы, священники, должны трубить трубами: это будет вам постановлением вечным в роды ваши;
NUM|10|9|и когда пойдете на войну в земле вашей против врага, наступающего на вас, трубите тревогу трубами, – и будете воспомянуты пред Господом, Богом вашим, и спасены будете от врагов ваших;
NUM|10|10|и в день веселия вашего, и в праздники ваши, и в новомесячия ваши трубите трубами при всесожжениях ваших и при мирных жертвах ваших, – и это будет напоминанием о вас пред Богом вашим. Я Господь, Бог ваш.
NUM|10|11|Во второй год, во второй месяц, в двадцатый [день] месяца поднялось облако от скинии откровения;
NUM|10|12|и отправились сыны Израилевы по станам своим из пустыни Синайской, и остановилось облако в пустыне Фаран.
NUM|10|13|И поднялись они в первый раз, по повелению Господню, [данному] чрез Моисея.
NUM|10|14|Поднято было во–первых знамя стана сынов Иудиных по ополчениям их; над ополчением их Наассон, сын Аминадава;
NUM|10|15|и над ополчением колена сынов Иссахаровых Нафанаил, сын Цуара;
NUM|10|16|и над ополчением колена сынов Завулоновых Елиав, сын Хелона.
NUM|10|17|И снята была скиния, и пошли сыны Гирсоновы и сыны Мерарины, носящие скинию.
NUM|10|18|И поднято было знамя стана Рувимова по ополчениям их; и над ополчением его Елицур, сын Шедеура;
NUM|10|19|и над ополчением колена сынов Симеоновых Шелумиил, сын Цуришаддая;
NUM|10|20|и над ополчением колена сынов Гадовых Елиасаф, сын Регуила.
NUM|10|21|Потом пошли сыны Каафовы, носящие святилище; скиния же была поставляема до прихода их.
NUM|10|22|И поднято было знамя стана сынов Ефремовых по ополчениям их; и над ополчением их Елишама, сын Аммиуда;
NUM|10|23|и над ополчением колена сынов Манассииных Гамалиил, сын Педацура;
NUM|10|24|и над ополчением колена сынов Вениаминовых Авидан, сын Гидеония.
NUM|10|25|Последним из всех станов поднято было знамя стана сынов Дановых с ополчениями их; и над ополчением их Ахиезер, сын Аммишаддая;
NUM|10|26|и над ополчением колена сынов Асировых Пагиил, сын Охрана;
NUM|10|27|и над ополчением колена сынов Неффалимовых Ахира, сын Енана.
NUM|10|28|Вот [порядок] шествия сынов Израилевых по ополчениям их. И отправились они.
NUM|10|29|И сказал Моисей Ховаву, сыну Рагуилову, Мадианитянину, родственнику Моисееву: мы отправляемся в то место, о котором Господь сказал: вам отдам его; иди с нами, мы сделаем тебе добро, ибо Господь доброе изрек об Израиле.
NUM|10|30|Но он сказал ему: не пойду; я пойду в свою землю и на свою родину.
NUM|10|31|[Моисей] же сказал: не оставляй нас, потому что ты знаешь, как располагаемся мы станом в пустыне, и будешь для нас глазом;
NUM|10|32|если пойдешь с нами, то добро, которое Господь сделает нам, мы сделаем тебе.
NUM|10|33|И отправились они от горы Господней на три дня пути, и ковчег завета Господня шел пред ними три дня пути, чтоб усмотреть им место, где остановиться.
NUM|10|34|И облако Господне осеняло их днем, когда они отправлялись из стана.
NUM|10|35|Когда поднимался ковчег в путь, Моисей говорил: восстань, Господи, и рассыплются враги Твои, и побегут от лица Твоего ненавидящие Тебя!
NUM|10|36|А когда останавливался ковчег, он говорил: возвратись, Господи, к тысячам и тьмам Израилевым!
NUM|11|1|Народ стал роптать вслух Господа; и Господь услышал, и воспламенился гнев Его, и возгорелся у них огонь Господень, и начал истреблять край стана.
NUM|11|2|И возопил народ к Моисею; и помолился Моисей Господу, и утих огонь.
NUM|11|3|И нарекли имя месту сему: Тавера, потому что возгорелся у них огонь Господень.
NUM|11|4|Пришельцы между ними стали обнаруживать прихоти; а с ними и сыны Израилевы сидели и плакали и говорили: кто накормит нас мясом?
NUM|11|5|Мы помним рыбу, которую в Египте мы ели даром, огурцы и дыни, и лук, и репчатый лук и чеснок;
NUM|11|6|а ныне душа наша изнывает; ничего нет, только манна в глазах наших.
NUM|11|7|Манна же была подобна кориандровому семени, видом, как бдолах;
NUM|11|8|народ ходил и собирал ее, и молол в жерновах или толок в ступе, и варил в котле, и делал из нее лепешки; вкус же ее подобен был вкусу лепешек с елеем.
NUM|11|9|И когда роса сходила на стан ночью, тогда сходила на него и манна.
NUM|11|10|Моисей слышал, что народ плачет в семействах своих, каждый у дверей шатра своего; и сильно воспламенился гнев Господень, и прискорбно было для Моисея.
NUM|11|11|И сказал Моисей Господу: для чего Ты мучишь раба Твоего? и почему я не нашел милости пред очами Твоими, что Ты возложил на меня бремя всего народа сего?
NUM|11|12|разве я носил во чреве весь народ сей, и разве я родил его, что Ты говоришь мне: неси его на руках твоих, как нянька носит ребенка, в землю, которую Ты с клятвою обещал отцам его?
NUM|11|13|откуда мне [взять] мяса, чтобы дать всему народу сему? ибо они плачут предо мною и говорят: дай нам есть мяса.
NUM|11|14|Я один не могу нести всего народа сего, потому что он тяжел для меня;
NUM|11|15|когда Ты так поступаешь со мною, то [лучше] умертви меня, если я нашел милость пред очами Твоими, чтобы мне не видеть бедствия моего.
NUM|11|16|И сказал Господь Моисею: собери Мне семьдесят мужей из старейшин Израилевых, которых ты знаешь, что они старейшины и надзиратели его, и возьми их к скинии собрания, чтобы они стали там с тобою;
NUM|11|17|Я сойду, и буду говорить там с тобою, и возьму от Духа, Который на тебе, и возложу на них, чтобы они несли с тобою бремя народа, а не один ты носил.
NUM|11|18|Народу же скажи: очиститесь к завтрашнему дню, и будете есть мясо; так как вы плакали вслух Господа и говорили: кто накормит нас мясом? хорошо нам было в Египте, – то и даст вам Господь мясо, и будете есть.
NUM|11|19|не один день будете есть, не два дня, не пять дней, не десять дней и не двадцать дней,
NUM|11|20|но целый месяц, пока не пойдет оно из ноздрей ваших и не сделается для вас отвратительным, за то, что вы презрели Господа, Который среди вас, и плакали пред Ним, говоря: для чего было нам выходить из Египта?
NUM|11|21|И сказал Моисей: шестьсот тысяч пеших в народе сем, среди которого я [нахожусь]; а Ты говоришь: Я дам им мясо, и будут есть целый месяц!
NUM|11|22|заколоть ли всех овец и волов, чтобы им было довольно? или вся рыба морская соберется, чтобы удовлетворить их?
NUM|11|23|И сказал Господь Моисею: разве рука Господня коротка? ныне ты увидишь, сбудется ли слово Мое тебе, или нет?
NUM|11|24|Моисей вышел и сказал народу слова Господни, и собрал семьдесят мужей из старейшин народа и поставил их около скинии.
NUM|11|25|И сошел Господь в облаке, и говорил с ним, и взял от Духа, Который на нем, и дал семидесяти мужам старейшинам. И когда почил на них Дух, они стали пророчествовать, но потом перестали.
NUM|11|26|Двое из мужей оставались в стане, одному имя Елдад, а другому имя Модад; но и на них почил Дух, и они пророчествовали в стане.
NUM|11|27|И прибежал отрок и донес Моисею, и сказал: Елдад и Модад пророчествуют в стане.
NUM|11|28|В ответ на это Иисус, сын Навин, служитель Моисея, один из избранных его, сказал: господин мой Моисей! запрети им.
NUM|11|29|Но Моисей сказал ему: не ревнуешь ли ты за меня? о, если бы все в народе Господнем были пророками, когда бы Господь послал Духа Своего на них!
NUM|11|30|И возвратился Моисей в стан, он и старейшины Израилевы.
NUM|11|31|И поднялся ветер от Господа, и принес от моря перепелов, и набросал их около стана, на путь дня по одну сторону и на путь дня по другую сторону около стана, на два почти локтя от земли.
NUM|11|32|И встал народ, и весь тот день, и всю ночь, и весь следующий день собирали перепелов; и кто мало собирал, тот собрал десять хомеров; и разложили их для себя вокруг стана.
NUM|11|33|Мясо еще было в зубах их и не было еще съедено, как гнев Господень возгорелся на народ, и поразил Господь народ весьма великою язвою.
NUM|11|34|И нарекли имя месту сему: Киброт–Гаттаава, ибо там похоронили прихотливый народ.
NUM|11|35|От Киброт–Гаттаавы двинулся народ в Асироф, и остановился в Асирофе.
NUM|12|1|И упрекали Мариам и Аарон Моисея за жену Ефиоплянку, которую он взял, – ибо он взял [за себя] Ефиоплянку, –
NUM|12|2|и сказали: одному ли Моисею говорил Господь? не говорил ли Он и нам? И услышал [сие] Господь.
NUM|12|3|Моисей же был человек кротчайший из всех людей на земле.
NUM|12|4|И сказал Господь внезапно Моисею и Аарону и Мариами: выйдите вы трое к скинии собрания. И вышли все трое.
NUM|12|5|И сошел Господь в облачном столпе, и стал у входа скинии, и позвал Аарона и Мариам, и вышли они оба.
NUM|12|6|И сказал: слушайте слова Мои: если бывает у вас пророк Господень, то Я открываюсь ему в видении, во сне говорю с ним;
NUM|12|7|но не так с рабом Моим Моисеем, – он верен во всем дому Моем:
NUM|12|8|устами к устам говорю Я с ним, и явно, а не в гаданиях, и образ Господа он видит; как же вы не убоялись упрекать раба Моего, Моисея?
NUM|12|9|И воспламенился гнев Господа на них, и Он отошел.
NUM|12|10|И облако отошло от скинии, и вот, Мариам покрылась проказою, как снегом. Аарон взглянул на Мариам, и вот, она в проказе.
NUM|12|11|И сказал Аарон Моисею: господин мой! не поставь нам в грех, что мы поступили глупо и согрешили;
NUM|12|12|не попусти, чтоб она была, как мертворожденный [младенец], у которого, когда он выходит из чрева матери своей, истлела уже половина тела.
NUM|12|13|И возопил Моисей к Господу, говоря: Боже, исцели ее!
NUM|12|14|И сказал Господь Моисею: если бы отец ее плюнул ей в лице, то не должна ли была бы она стыдиться семь дней? итак пусть будет она в заключении семь дней вне стана, а после опять возвратится.
NUM|12|15|И пробыла Мариам в заключении вне стана семь дней, и народ не отправлялся в путь, доколе не возвратилась Мариам.
NUM|12|16|После сего народ двинулся из Асирофа, и остановился в пустыне Фаран.
NUM|13|1|И сказал Господь Моисею, говоря:
NUM|13|2|пошли от себя людей, чтобы они высмотрели землю Ханаанскую, которую Я даю сынам Израилевым; по одному человеку от колена отцов их пошлите, главных из них.
NUM|13|3|И послал их Моисей из пустыни Фаран, по повелению Господню, и все они мужи главные у сынов Израилевых.
NUM|13|4|Вот имена их: из колена Рувимова Саммуа, сын Закхуров,
NUM|13|5|из колена Симеонова Сафат, сын Хориев,
NUM|13|6|из колена Иудина Халев, сын Иефонниин,
NUM|13|7|из колена Иссахарова Игал, сын Иосифов,
NUM|13|8|из колена Ефремова Осия, сын Навин,
NUM|13|9|из колена Вениаминова Фалтий, сын Рафуев,
NUM|13|10|из колена Завулонова Гаддиил, сын Содиев,
NUM|13|11|из колена Иосифова от Манассии Гаддий, сын Сусиев,
NUM|13|12|из колена Данова Аммиил, сын Гемаллиев,
NUM|13|13|из колена Асирова Сефур, сын Михаилев,
NUM|13|14|из колена Неффалимова Нахбий, сын Вофсиев,
NUM|13|15|из колена Гадова Геуил, сын Махиев.
NUM|13|16|Вот имена мужей, которых посылал Моисей высмотреть землю. И назвал Моисей Осию, сына Навина, Иисусом.
NUM|13|17|И послал их Моисей высмотреть землю Ханаанскую и сказал им: пойдите в эту южную страну, и взойдите на гору,
NUM|13|18|и осмотрите землю, какова она, и народ живущий на ней, силен ли он или слаб, малочислен ли он или многочислен?
NUM|13|19|и какова земля, на которой он живет, хороша ли она или худа? и каковы города, в которых он живет, в шатрах ли он живет или в укреплениях?
NUM|13|20|и какова земля, тучна ли она или тоща? есть ли на [ней] дерева или нет? будьте смелы, и возьмите от плодов земли. Было же это ко времени созревания винограда.
NUM|13|21|Они пошли и высмотрели землю от пустыни Син даже до Рехова, близ Емафа;
NUM|13|22|и пошли в южную страну, и дошли до Хеврона, где жили Ахиман, Сесай и Фалмай, дети Енаковы: Хеврон же построен был семью годами прежде Цоана, [города] Египетского;
NUM|13|23|и пришли к долине Есхол, и срезали там виноградную ветвь с одною кистью ягод, и понесли ее на шесте двое; [взяли] также гранатовых яблок и смокв;
NUM|13|24|место сие назвали долиною Есхол, по причине виноградной кисти, которую срезали там сыны Израилевы.
NUM|13|25|И высмотрев землю, возвратились они через сорок дней.
NUM|13|26|И пошли и пришли к Моисею и Аарону и ко всему обществу сынов Израилевых в пустыню Фаран, в Кадес, и принесли им и всему обществу ответ, и показали им плоды земли;
NUM|13|27|и рассказывали ему и говорили: мы ходили в землю, в которую ты посылал нас; в ней подлинно течет молоко и мед, и вот плоды ее;
NUM|13|28|но народ, живущий на земле той, силен, и города укрепленные, весьма большие, и сынов Енаковых мы видели там;
NUM|13|29|Амалик живет на южной части земли, Хеттеи, Иевусеи и Аморреи живут на горе, Хананеи же живут при море и на берегу Иордана.
NUM|13|30|Но Халев успокаивал народ пред Моисеем, говоря: пойдем и завладеем ею, потому что мы можем одолеть ее.
NUM|13|31|А те, которые ходили с ним, говорили: не можем мы идти против народа сего, ибо он сильнее нас.
NUM|13|32|И распускали худую молву о земле, которую они осматривали, между сынами Израилевыми, говоря: земля, которую проходили мы для осмотра, есть земля, поедающая живущих на ней, и весь народ, который видели мы среди ее, люди великорослые;
NUM|13|33|там видели мы и исполинов, сынов Енаковых, от исполинского рода; и мы были в глазах наших [пред ними], как саранча, такими же были мы и в глазах их.
NUM|14|1|И подняло все общество вопль, и плакал народ во [всю] ту ночь;
NUM|14|2|и роптали на Моисея и Аарона все сыны Израилевы, и все общество сказало им: о, если бы мы умерли в земле Египетской, или умерли бы в пустыне сей!
NUM|14|3|и для чего Господь ведет нас в землю сию, чтобы мы пали от меча? жены наши и дети наши достанутся в добычу [врагам]; не лучше ли нам возвратиться в Египет?
NUM|14|4|И сказали друг другу: поставим себе начальника и возвратимся в Египет.
NUM|14|5|И пали Моисей и Аарон на лица свои пред всем собранием общества сынов Израилевых.
NUM|14|6|И Иисус, сын Навин, и Халев, сын Иефонниин, из осматривавших землю, разодрали одежды свои
NUM|14|7|и сказали всему обществу сынов Израилевых: земля, которую мы проходили для осмотра, очень, очень хороша;
NUM|14|8|если Господь милостив к нам, то введет нас в землю сию и даст нам ее – эту землю, в которой течет молоко и мед;
NUM|14|9|только против Господа не восставайте и не бойтесь народа земли сей; ибо он достанется нам на съедение: защиты у них не стало, а с нами Господь; не бойтесь их.
NUM|14|10|И сказало все общество: побить их камнями! Но слава Господня явилась в скинии собрания всем сынам Израилевым.
NUM|14|11|И сказал Господь Моисею: доколе будет раздражать Меня народ сей? и доколе будет он не верить Мне при всех знамениях, которые делал Я среди его?
NUM|14|12|поражу его язвою и истреблю его и произведу от тебя народ многочисленнее и сильнее его.
NUM|14|13|Но Моисей сказал Господу: услышат Египтяне, из среды которых Ты силою Твоею вывел народ сей,
NUM|14|14|и скажут жителям земли сей, которые слышали, что Ты, Господь, находишься среди народа сего, и что Ты, Господь, даешь им видеть Себя лицем к лицу, и облако Твое стоит над ними, и Ты идешь пред ними днем в столпе облачном, а ночью в столпе огненном;
NUM|14|15|и если Ты истребишь народ сей, как одного человека, то народы, которые слышали славу Твою, скажут:
NUM|14|16|Господь не мог ввести народ сей в землю, которую Он с клятвою обещал ему, а потому и погубил его в пустыне.
NUM|14|17|Итак да возвеличится сила Господня, как Ты сказал, говоря:
NUM|14|18|Господь долготерпелив и многомилостив, прощающий беззакония и преступления, и не оставляющий без наказания, но наказывающий беззаконие отцов в детях до третьего и четвертого рода.
NUM|14|19|Прости грех народу сему по великой милости Твоей, как Ты прощал народ сей от Египта доселе.
NUM|14|20|И сказал Господь [Моисею]: прощаю по слову твоему;
NUM|14|21|но жив Я, и славы Господней полна вся земля:
NUM|14|22|все, которые видели славу Мою и знамения Мои, сделанные Мною в Египте и в пустыне, и искушали Меня уже десять раз, и не слушали гласа Моего,
NUM|14|23|не увидят земли, которую Я с клятвою обещал отцам их; все, раздражавшие Меня, не увидят ее;
NUM|14|24|но раба Моего, Халева, за то, что в нем был иной дух, и он совершенно повиновался Мне, введу в землю, в которую он ходил, и семя его наследует ее;
NUM|14|25|Амаликитяне и Хананеи живут в долине; завтра обратитесь и идите в пустыню к Чермному морю.
NUM|14|26|И сказал Господь Моисею и Аарону, говоря:
NUM|14|27|доколе злому обществу сему роптать на Меня? ропот сынов Израилевых, которым они ропщут на Меня, Я слышу.
NUM|14|28|Скажи им: живу Я, говорит Господь: как говорили вы вслух Мне, так и сделаю вам;
NUM|14|29|в пустыне сей падут тела ваши, и все вы исчисленные, сколько вас числом, от двадцати лет и выше, которые роптали на Меня,
NUM|14|30|не войдете в землю, на которой Я, подъемля руку Мою, [клялся] поселить вас, кроме Халева, сына Иефонниина, и Иисуса, сына Навина;
NUM|14|31|детей ваших, о которых вы говорили, что они достанутся в добычу [врагам], Я введу [туда], и они узнают землю, которую вы презрели,
NUM|14|32|а ваши трупы падут в пустыне сей;
NUM|14|33|а сыны ваши будут кочевать в пустыне сорок лет, и будут нести [наказание] за блудодейство ваше, доколе не погибнут все тела ваши в пустыне;
NUM|14|34|по числу сорока дней, в которые вы осматривали землю, вы понесете наказание за грехи ваши сорок лет, год за день, дабы вы познали, [что] [значит] быть оставленным Мною.
NUM|14|35|Я, Господь, говорю, и так и сделаю со всем сим злым обществом, восставшим против Меня: в пустыне сей все они погибнут и перемрут.
NUM|14|36|И те, которых посылал Моисей для осмотрения земли, и которые, возвратившись, возмутили против него все сие общество, распуская худую молву о земле,
NUM|14|37|сии, распустившие худую молву о земле, умерли, быв поражены пред Господом;
NUM|14|38|только Иисус, сын Навин, и Халев, сын Иефонниин, остались живы из тех мужей, которые ходили осматривать землю.
NUM|14|39|И сказал Моисей слова сии пред всеми сынами Израилевыми, и народ сильно опечалился.
NUM|14|40|И, встав рано поутру, пошли на вершину горы, говоря: вот, мы пойдем на то место, о котором сказал Господь, ибо мы согрешили.
NUM|14|41|Моисей сказал: для чего вы преступаете повеление Господне? это будет безуспешно;
NUM|14|42|не ходите, ибо нет среди вас Господа, чтобы не поразили вас враги ваши;
NUM|14|43|ибо Амаликитяне и Хананеи там пред вами, и вы падете от меча, потому что вы отступили от Господа, и не будет с вами Господа.
NUM|14|44|Но они дерзнули подняться на вершину горы; ковчег же завета Господня и Моисей не оставляли стана.
NUM|14|45|И сошли Амаликитяне и Хананеи, живущие на горе той, и разбили их, и гнали их до Хормы.
NUM|15|1|И сказал Господь Моисею, говоря:
NUM|15|2|объяви сынам Израилевым и скажи им: когда вы войдете в землю вашего жительства, которую Я даю вам,
NUM|15|3|и будете приносить жертву Господу, всесожжение, или жертву заколаемую, от волов и овец, во исполнение обета, или по усердию, или в праздники ваши, дабы сделать приятное благоухание Господу, –
NUM|15|4|тогда приносящий жертву свою Господу должен принести в приношение от хлеба десятую часть [ефы] пшеничной муки, смешанной с четвертою частью гина елея;
NUM|15|5|и вина для возлияния приноси четвертую часть гина при всесожжении, или при заколаемой жертве, на каждого агнца.
NUM|15|6|А принося овна, приноси в приношение хлебное две десятых части [ефы] пшеничной муки, смешанной с третьею частью гина елея;
NUM|15|7|и вина для возлияния приноси третью часть гина в приятное благоухание Господу.
NUM|15|8|Если молодого вола приносишь во всесожжение или жертву заколаемую, во исполнение обета или в мирную жертву Господу,
NUM|15|9|то вместе с волом должно принести приношения хлебного три десятых части [ефы] пшеничной муки, смешанной с половиною гина елея;
NUM|15|10|и вина для возлияния приноси полгина в жертву, в приятное благоухание Господу.
NUM|15|11|Так делай при каждом приношении вола и овна и агнца из овец, или коз;
NUM|15|12|по числу [жертв], которые вы приносите, так делайте при каждой, по числу их.
NUM|15|13|Всякий туземец так должен делать это, принося жертву в приятное благоухание Господу;
NUM|15|14|и если будет между вами жить пришелец, или кто бы ни был среди вас в роды ваши, и принесет жертву в приятное благоухание Господу, то и он должен делать так, как вы делаете;
NUM|15|15|для вас, общество [Господне], и для пришельца, живущего [у вас], устав один, устав вечный в роды ваши: что вы, то и пришелец да будет пред Господом;
NUM|15|16|закон один и одни права да будут для вас и для пришельца, живущего у вас.
NUM|15|17|И сказал Господь Моисею, говоря:
NUM|15|18|объяви сынам Израилевым и скажи им: когда вы войдете в землю, в которую Я веду вас,
NUM|15|19|и будете есть хлеб той земли, то возносите возношение Господу;
NUM|15|20|от начатков теста вашего лепешку возносите в возношение; возносите ее так, как возношение с гумна;
NUM|15|21|от начатков теста вашего отдавайте в возношение Господу в роды ваши.
NUM|15|22|Если же преступите по неведению и не исполните всех сих заповедей, которые изрек Господь Моисею,
NUM|15|23|всего, что заповедал вам Господь чрез Моисея, от того дня, в который Господь заповедал вам, и впредь в роды ваши, –
NUM|15|24|то, если по недосмотру общества сделана ошибка, пусть все общество принесет одного молодого вола во всесожжение, в приятное благоухание Господу, с хлебным приношением и возлиянием его, по уставу, и одного козла в жертву за грех;
NUM|15|25|и очистит священник все общество сынов Израилевых, и будет прощено им, ибо это была ошибка, и они принесли приношение свое в жертву Господу, и жертву за грех свой пред Господом, за свою ошибку;
NUM|15|26|и будет прощено всему обществу сынов Израилевых и пришельцу, живущему между ними, потому что весь народ сделал это по ошибке.
NUM|15|27|Если же один кто согрешит по неведению, то пусть принесет козу однолетнюю в жертву за грех;
NUM|15|28|и очистит священник душу, сделавшую по ошибке грех пред Господом, и очищена будет, и прощено будет ей;
NUM|15|29|один закон да будет для вас, как для природного жителя из сынов Израилевых, так и для пришельца, живущего у вас, если кто сделает что по ошибке.
NUM|15|30|Если же кто из туземцев, или из пришельцев, сделает что дерзкою рукою, то он хулит Господа: истребится душа та из народа своего,
NUM|15|31|ибо слово Господне он презрел и заповедь Его нарушил; истребится душа та; грех ее на ней.
NUM|15|32|Когда сыны Израилевы были в пустыне, нашли человека, собиравшего дрова в день субботы;
NUM|15|33|и привели его нашедшие его собирающим дрова к Моисею и Аарону и ко всему обществу;
NUM|15|34|и посадили его под стражу, потому что не было еще определено, что должно с ним сделать.
NUM|15|35|И сказал Господь Моисею: должен умереть человек сей; пусть побьет его камнями все общество вне стана.
NUM|15|36|И вывело его все общество вон из стана, и побили его камнями, и он умер, как повелел Господь Моисею.
NUM|15|37|И сказал Господь Моисею, говоря:
NUM|15|38|объяви сынам Израилевым и скажи им, чтоб они делали себе кисти на краях одежд своих в роды их, и в кисти, которые на краях, вставляли нити из голубой шерсти;
NUM|15|39|и будут они в кистях у вас для того, чтобы вы, смотря на них, вспоминали все заповеди Господни, и исполняли их, и не ходили вслед сердца вашего и очей ваших, которые влекут вас к блудодейству,
NUM|15|40|чтобы вы помнили и исполняли все заповеди Мои и были святы пред Богом вашим.
NUM|15|41|Я Господь, Бог ваш, Который вывел вас из земли Египетской, чтоб быть вашим Богом: Я Господь, Бог ваш.
NUM|16|1|Корей, сын Ицгара, сын Каафов, сын Левиин, и Дафан и Авирон, сыны Елиава, и Авнан, сын Фалефа, сыны Рувимовы,
NUM|16|2|восстали на Моисея, и [с ними] из сынов Израилевых двести пятьдесят мужей, начальники общества, призываемые на собрания, люди именитые.
NUM|16|3|И собрались против Моисея и Аарона и сказали им: полно вам; все общество, все святы, и среди их Господь! почему же вы ставите себя выше народа Господня?
NUM|16|4|Моисей, услышав это, пал на лице свое
NUM|16|5|и сказал Корею и всем сообщникам его, говоря: завтра покажет Господь, кто Его, и кто свят, чтобы приблизить его к Себе; и кого Он изберет, того и приблизит к Себе;
NUM|16|6|вот что сделайте: Корей и все сообщники его возьмите себе кадильницы
NUM|16|7|и завтра положите в них огня и всыпьте в них курения пред Господом; и кого изберет Господь, тот и будет свят. Полно вам, сыны Левиины!
NUM|16|8|И сказал Моисей Корею: послушайте, сыны Левия!
NUM|16|9|неужели мало вам того, что Бог Израилев отделил вас от общества Израильского и приблизил вас к Себе, чтобы вы исполняли службы при скинии Господней и стояли пред обществом, служа для них?
NUM|16|10|Он приблизил тебя и с тобою всех братьев твоих, сынов Левия, и вы домогаетесь еще и священства.
NUM|16|11|Итак ты и все твое общество собрались против Господа. Что Аарон, что вы ропщете на него?
NUM|16|12|И послал Моисей позвать Дафана и Авирона, сынов Елиава. Но они сказали: не пойдем!
NUM|16|13|разве мало того, что ты вывел нас из земли, в которой течет молоко и мед, чтобы погубить нас в пустыне? и ты еще хочешь властвовать над нами!
NUM|16|14|привел ли ты нас в землю, где течет молоко и мед, и дал ли нам во владение поля и виноградники? глаза людей сих ты хочешь ослепить? не пойдем!
NUM|16|15|Моисей весьма огорчился и сказал Господу: не обращай взора Твоего на приношение их; я не взял ни у одного из них осла и не сделал зла ни одному из них.
NUM|16|16|И сказал Моисей Корею: завтра ты и все общество твое будьте пред лицем Господа, ты, они и Аарон;
NUM|16|17|и возьмите каждый свою кадильницу, и положите в них курения, и принесите пред лице Господне каждый свою кадильницу, двести пятьдесят кадильниц; ты и Аарон, каждый свою кадильницу.
NUM|16|18|И взял каждый свою кадильницу, и положили в них огня, и всыпали в них курения, и стали при входе в скинию собрания; также и Моисей и Аарон.
NUM|16|19|И собрал против них Корей все общество ко входу скинии собрания. И явилась слава Господня всему обществу.
NUM|16|20|И сказал Господь Моисею и Аарону, говоря:
NUM|16|21|отделитесь от общества сего, и Я истреблю их во мгновение.
NUM|16|22|Они же пали на лица свои и сказали: Боже, Боже духов всякой плоти! один человек согрешил, и Ты гневаешься на все общество?
NUM|16|23|и сказал Господь Моисею, говоря:
NUM|16|24|скажи обществу: отступите со всех сторон от жилища Корея, Дафана и Авирона.
NUM|16|25|И встал Моисей, и пошел к Дафану и Авирону, и за ним пошли старейшины Израилевы.
NUM|16|26|И сказал обществу: отойдите от шатров нечестивых людей сих, и не прикасайтесь ни к чему, что принадлежит им, чтобы не погибнуть вам во всех грехах их.
NUM|16|27|И отошли они со всех сторон от жилища Корея, Дафана и Авирона; а Дафан и Авирон вышли и стояли у дверей шатров своих с женами своими и сыновьями своими и с малыми детьми своими.
NUM|16|28|И сказал Моисей: из сего узнаете, что Господь послал меня делать все дела сии, а не по своему произволу [я делаю сие]:
NUM|16|29|если они умрут, как умирают все люди, и постигнет их такое наказание, какое [постигает] всех людей, то не Господь послал меня;
NUM|16|30|а если Господь сотворит необычайное, и земля разверзет уста свои и поглотит их и все, что у них, и они живые сойдут в преисподнюю, то знайте, что люди сии презрели Господа.
NUM|16|31|Лишь только он сказал слова сии, расселась земля под ними;
NUM|16|32|и разверзла земля уста свои, и поглотила их и домы их, и всех людей Кореевых и все имущество;
NUM|16|33|и сошли они со всем, что принадлежало им, живые в преисподнюю, и покрыла их земля, и погибли они из среды общества.
NUM|16|34|И все Израильтяне, которые были вокруг них, побежали при их вопле, дабы, говорили они, и нас не поглотила земля.
NUM|16|35|И вышел огонь от Господа и пожрал тех двести пятьдесят мужей, которые принесли курение.
NUM|16|36|И сказал Господь Моисею, говоря:
NUM|16|37|скажи Елеазару, сыну Аарона, священнику, пусть он соберет кадильницы сожженных и огонь выбросит вон; ибо освятились
NUM|16|38|кадильницы грешников сих смертью их, и пусть разобьют их в листы для покрытия жертвенника, ибо они принесли их пред лице Господа, и они сделались освященными; и будут они знамением для сынов Израилевых.
NUM|16|39|И взял Елеазар священник медные кадильницы, которые принесли сожженные, и разбили их в листы для покрытия жертвенника,
NUM|16|40|в память сынам Израилевым, чтобы никто посторонний, который не от семени Аарона, не приступал приносить курение пред лице Господне, и не было с ним, что с Кореем и сообщниками его, как говорил ему Господь чрез Моисея.
NUM|16|41|На другой день все общество сынов Израилевых возроптало на Моисея и Аарона и говорило: вы умертвили народ Господень.
NUM|16|42|И когда собралось общество против Моисея и Аарона, они обратились к скинии собрания, и вот, облако покрыло ее, и явилась слава Господня.
NUM|16|43|И пришел Моисей и Аарон к скинии собрания.
NUM|16|44|И сказал Господь Моисею, говоря:
NUM|16|45|отсторонитесь от общества сего, и Я погублю их во мгновение. Но они пали на лица свои.
NUM|16|46|И сказал Моисей Аарону: возьми кадильницу и положи в нее огня с жертвенника и всыпь курения, и неси скорее к обществу и заступи их, ибо вышел гнев от Господа, [и] началось поражение.
NUM|16|47|И взял Аарон, как сказал Моисей, и побежал в среду общества, и вот, уже началось поражение в народе. И он положил курения и заступил народ;
NUM|16|48|стал он между мертвыми и живыми, и поражение прекратилось.
NUM|16|49|И умерло от поражения четырнадцать тысяч семьсот человек, кроме умерших по делу Корееву.
NUM|16|50|И возвратился Аарон к Моисею, ко входу скинии собрания, после того как поражение прекратилось.
NUM|17|1|И сказал Господь Моисею, говоря:
NUM|17|2|скажи сынам Израилевым и возьми у них по жезлу от колена, от всех начальников их по коленам, двенадцать жезлов, и каждого имя напиши на жезле его;
NUM|17|3|имя Аарона напиши на жезле Левиином, ибо один жезл от начальника колена их [должны они дать];
NUM|17|4|и положи их в скинии собрания, пред [ковчегом] откровения, где являюсь Я вам;
NUM|17|5|и кого Я изберу, того жезл расцветет; и так Я успокою ропот сынов Израилевых, которым они ропщут на вас.
NUM|17|6|И сказал Моисей сынам Израилевым, и дали ему все начальники их, от каждого начальника по жезлу, по коленам их двенадцать жезлов, и жезл Ааронов был среди жезлов их.
NUM|17|7|И положил Моисей жезлы пред лицем Господа в скинии откровения.
NUM|17|8|На другой день вошел Моисей в скинию откровения, и вот, жезл Ааронов, от дома Левиина, расцвел, пустил почки, дал цвет и принес миндали.
NUM|17|9|И вынес Моисей все жезлы от лица Господня ко всем сынам Израилевым. И увидели они это и взяли каждый свой жезл.
NUM|17|10|И сказал Господь Моисею: положи опять жезл Ааронов пред [ковчегом] откровения на сохранение, в знамение для непокорных, чтобы прекратился ропот их на Меня, и они не умирали.
NUM|17|11|Моисей сделал это; как повелел ему Господь, так он и сделал.
NUM|17|12|И сказали сыны Израилевы Моисею: вот, мы умираем, погибаем, все погибаем!
NUM|17|13|всякий, приближающийся к скинии Господней, умирает: не придется ли всем нам умереть?
NUM|18|1|И сказал Господь Аарону: ты и сыны твои и дом отца твоего с тобою понесете на себе грех за [небрежность во] святилище; и ты и сыны твои с тобою понесете на себе грех за [неисправность] в священстве вашем.
NUM|18|2|Также и братьев твоих, колено Левиино, племя отца твоего, возьми себе: пусть они будут при тебе и служат тебе, а ты и сыны твои с тобою [будете] при скинии откровения;
NUM|18|3|пусть они отправляют службу тебе и службу во всей скинии; только чтобы не приступали к вещам святилища и к жертвеннику, дабы не умереть и им и вам.
NUM|18|4|Пусть они будут при тебе и отправляют службу в скинии собрания, все работы по скинии; а посторонний не должен приближаться к вам.
NUM|18|5|Так отправляйте службу во святилище и при жертвеннике, дабы не было впредь гнева на сынов Израилевых;
NUM|18|6|ибо братьев ваших, левитов, Я взял от сынов Израилевых и дал их вам, в дар Господу, для отправления службы при скинии собрания;
NUM|18|7|и ты и сыны твои с тобою наблюдайте священство ваше во всем, что принадлежит жертвеннику и что внутри за завесою, и служите; вам даю Я в дар службу священства, а посторонний, приступивший, предан будет смерти.
NUM|18|8|И сказал Господь Аарону: вот, Я поручаю тебе наблюдать за возношениями Мне; от всего, посвящаемого сынами Израилевыми, Я дал тебе и сынам твоим, ради священства вашего, уставом вечным;
NUM|18|9|вот, что принадлежит тебе из святынь великих, от сожигаемого: всякое приношение их хлебное, и всякая жертва их за грех, и всякая жертва их повинности, что они принесут Мне; это великая святыня тебе и сынам твоим.
NUM|18|10|На святейшем месте ешьте это; все мужеского пола могут есть. это святынею да будет для тебя.
NUM|18|11|И вот, что тебе из возношений даров их: все возношения сынов Израилевых Я дал тебе и сынам твоим и дочерям твоим с тобою, уставом вечным; всякий чистый в доме твоем может есть это.
NUM|18|12|Все лучшее из елея и все лучшее из винограда и хлеба, начатки их, которые они дают Господу, Я отдал тебе;
NUM|18|13|все первые произведения земли их, которые они принесут Господу, да будут твоими; всякий чистый в доме твоем может есть это.
NUM|18|14|Все заклятое в земле Израилевой да будет твоим.
NUM|18|15|Все, разверзающее ложесна у всякой плоти, которую приносят Господу, из людей и из скота, да будет твоим; только первенец из людей должен быть выкуплен, и первородное из скота нечистого должно быть выкуплено;
NUM|18|16|а выкуп за них: начиная от одного месяца, по оценке твоей, бери выкуп пять сиклей серебра, по сиклю священному, который в двадцать гер;
NUM|18|17|но за первородное из волов, и за первородное из овец, и за первородное из коз, не бери выкупа: они святыня; кровью их окропляй жертвенник, и тук их сожигай в жертву, в приятное благоухание Господу;
NUM|18|18|мясо же их тебе принадлежит, равно как грудь возношения и правое плечо тебе принадлежит.
NUM|18|19|Все возносимые святыни, которые возносят сыны Израилевы Господу, отдаю тебе и сынам твоим и дочерям твоим с тобою, уставом вечным; это завет соли вечный пред Господом, данный для тебя и потомства твоего с тобою.
NUM|18|20|И сказал Господь Аарону: в земле их не будешь иметь удела и части не будет тебе между ними; Я часть твоя и удел твой среди сынов Израилевых;
NUM|18|21|а сынам Левия, вот, Я дал в удел десятину из всего, что у Израиля, за службу их, за то, что они отправляют службы в скинии собрания;
NUM|18|22|и сыны Израилевы не должны впредь приступать к скинии собрания, чтобы не понести греха и не умереть:
NUM|18|23|пусть левиты исправляют службы в скинии собрания и несут на себе грех их. Это устав вечный в роды ваши; среди же сынов Израилевых они не получат удела;
NUM|18|24|так как десятину сынов Израилевых, которую они приносят в возношение Господу, Я отдаю левитам в удел, потому и сказал Я им: между сынами Израилевыми они не получат удела.
NUM|18|25|И сказал Господь Моисею, говоря:
NUM|18|26|объяви левитам и скажи им: когда вы будете брать от сынов Израилевых десятину, которую Я дал вам от них в удел, то возносите из нее возношение Господу, десятину из десятины, –
NUM|18|27|и вменено будет вам это возношение ваше, как хлеб с гумна и как взятое от точила;
NUM|18|28|так и вы будете возносить возношение Господу из всех десятин ваших, которые будете брать от сынов Израилевых, и будете давать из них возношение Господне Аарону священнику;
NUM|18|29|из всего, даруемого вам, возносите возношение Господу, из всего лучшего освящаемого.
NUM|18|30|И скажи им: когда вы принесете из сего лучшее, то это вменено будет левитам, как получаемое с гумна и получаемое от точила;
NUM|18|31|вы можете есть это на всяком месте, вы и семейства ваши, ибо это вам плата за работы ваши в скинии собрания;
NUM|18|32|и не понесете за это греха, когда принесете лучшее из сего; и посвящаемого сынами Израилевыми не оскверните, и не умрете.
NUM|19|1|И сказал Господь Моисею и Аарону, говоря:
NUM|19|2|вот устав закона, который заповедал Господь, говоря: скажи сынам Израилевым, пусть приведут тебе рыжую телицу без порока, у которой нет недостатка, [и] на которой не было ярма;
NUM|19|3|и отдайте ее Елеазару священнику, и выведет ее вон из стана, и заколют ее при нем;
NUM|19|4|и пусть возьмет Елеазар священник перстом своим крови ее и кровью покропит к передней стороне скинии собрания семь раз;
NUM|19|5|и сожгут телицу при его глазах: кожу ее и мясо ее и кровь ее с нечистотою ее пусть сожгут;
NUM|19|6|и пусть возьмет священник кедрового дерева и иссопа и нить из червленой шерсти и бросит на сожигаемую телицу;
NUM|19|7|и пусть вымоет священник одежды свои, и омоет тело свое водою, и потом войдет в стан, и нечист будет священник до вечера.
NUM|19|8|И сожигавший ее пусть вымоет одежды свои водою, и омоет тело свое водою, и нечист будет до вечера;
NUM|19|9|и кто–нибудь чистый пусть соберет пепел телицы и положит вне стана на чистом месте, и будет он сохраняться для общества сынов Израилевых, для воды очистительной: это жертва за грех;
NUM|19|10|и собиравший пепел телицы пусть вымоет одежды свои, и нечист будет до вечера. Это для сынов Израилевых и для пришельцев, живущих у них, да будет уставом вечным.
NUM|19|11|Кто прикоснется к мертвому телу какого–либо человека, нечист будет семь дней:
NUM|19|12|он должен очистить себя сею [водою] в третий день и в седьмой день, и будет чист; если же он не очистит себя в третий и седьмой день, то не будет чист;
NUM|19|13|всякий, прикоснувшийся к мертвому телу какого–либо человека умершего и не очистивший себя, осквернит жилище Господа: истребится человек тот из среды Израиля, ибо он не окроплен очистительною водою, он нечист, еще нечистота его на нем.
NUM|19|14|Вот закон: если человек умрет в шатре, то всякий, кто придет в шатер, и все, что в шатре, нечисто будет семь дней;
NUM|19|15|всякий открытый сосуд, который не обвязан и не покрыт, нечист.
NUM|19|16|Всякий, кто прикоснется на поле к убитому мечом, или к умершему, или к кости человеческой, или ко гробу, нечист будет семь дней.
NUM|19|17|Для нечистого пусть возьмут пепла той сожженной жертвы за грех и нальют на него живой воды в сосуд;
NUM|19|18|и пусть кто–нибудь чистый возьмет иссоп, и омочит его в воде, и окропит шатер и все сосуды и людей, которые находятся в нем, и прикоснувшегося к кости [человеческой], или к убитому, или к умершему, или ко гробу;
NUM|19|19|и пусть окропит чистый нечистого в третий и седьмой день, и очистит его в седьмой день; и вымоет он одежды свои, и омоет [тело свое] водою, и к вечеру будет чист.
NUM|19|20|Если же кто будет нечист и не очистит себя, то истребится человек тот из среды народа, ибо он осквернил святилище Господа; очистительною водою он не окроплен, он нечист.
NUM|19|21|И да будет это для них уставом вечным. И кропивший очистительною водою пусть вымоет одежды свои; и прикоснувшийся к очистительной воде нечист будет до вечера.
NUM|19|22|И все, к чему прикоснется нечистый, будет нечисто; и прикоснувшийся человек нечист будет до вечера.
NUM|20|1|И пришли сыны Израилевы, все общество, в пустыню Син в первый месяц, и остановился народ в Кадесе, и умерла там Мариам и погребена там.
NUM|20|2|И не было воды для общества, и собрались они против Моисея и Аарона;
NUM|20|3|и возроптал народ на Моисея и сказал: о, если бы умерли тогда и мы, когда умерли братья наши пред Господом!
NUM|20|4|зачем вы привели общество Господне в эту пустыню, чтобы умереть здесь нам и скоту нашему?
NUM|20|5|и для чего вывели вы нас из Египта, чтобы привести нас на это негодное место, где нельзя сеять, нет ни смоковниц, ни винограда, ни гранатовых яблок, ни даже воды для питья?
NUM|20|6|И пошел Моисей и Аарон от народа ко входу скинии собрания, и пали на лица свои, и явилась им слава Господня.
NUM|20|7|И сказал Господь Моисею, говоря:
NUM|20|8|Возьми жезл и собери общество, ты и Аарон, брат твой, и скажите в глазах их скале, и она даст из себя воду: и так ты изведешь им воду из скалы, и напоишь общество и скот его.
NUM|20|9|И взял Моисей жезл от лица Господа, как Он повелел ему.
NUM|20|10|И собрали Моисей и Аарон народ к скале, и сказал он им: послушайте, непокорные, разве нам из этой скалы извести для вас воду?
NUM|20|11|И поднял Моисей руку свою и ударил в скалу жезлом своим дважды, и потекло много воды, и пило общество и скот его.
NUM|20|12|И сказал Господь Моисею и Аарону: за то, что вы не поверили Мне, чтоб явить святость Мою пред очами сынов Израилевых, не введете вы народа сего в землю, которую Я даю ему.
NUM|20|13|Это вода Меривы, у которой вошли в распрю сыны Израилевы с Господом, и Он явил им святость Свою.
NUM|20|14|И послал Моисей из Кадеса послов к Царю Едомскому [сказать]: так говорит брат твой Израиль: ты знаешь все трудности, которые постигли нас;
NUM|20|15|отцы наши перешли в Египет, и мы жили в Египте много времени, и худо поступали Египтяне с нами и отцами нашими;
NUM|20|16|и воззвали мы к Господу, и услышал Он голос наш, и послал Ангела, и вывел нас из Египта; и вот, мы в Кадесе, городе у самого предела твоего;
NUM|20|17|позволь нам пройти землею твоею: мы не пойдем по полям и по виноградникам и не будем пить воды из колодезей [твоих]; но пойдем дорогою царскою, не своротим ни направо ни налево, доколе не перейдем пределов твоих.
NUM|20|18|Но Едом сказал ему: не проходи через меня, иначе я с мечом выступлю против тебя.
NUM|20|19|И сказали ему сыны Израилевы: мы пойдем большою дорогою, и если будем пить твою воду, я и скот мой, то буду платить за нее; только ногами моими пройду, что ничего не стоит.
NUM|20|20|Но он сказал: не проходи. И выступил против него Едом с многочисленным народом и с сильною рукою.
NUM|20|21|Итак не согласился Едом позволить Израилю пройти чрез его пределы, и Израиль пошел в сторону от него.
NUM|20|22|И отправились сыны Израилевы из Кадеса, и пришло все общество к горе Ор.
NUM|20|23|И сказал Господь Моисею и Аарону на горе Ор, у пределов земли Едомской, говоря:
NUM|20|24|пусть приложится Аарон к народу своему; ибо он не войдет в землю, которую Я даю сынам Израилевым, за то, что вы непокорны были повелению Моему у вод Меривы;
NUM|20|25|и возьми Аарона и Елеазара, сына его, и возведи их на гору Ор.
NUM|20|26|и сними с Аарона одежды его, и облеки в них Елеазара, сына его, и пусть Аарон отойдет и умрет там.
NUM|20|27|И сделал Моисей так, как повелел Господь. Пошли они на гору Ор в глазах всего общества,
NUM|20|28|и снял Моисей с Аарона одежды его, и облек в них Елеазара, сына его; и умер там Аарон на вершине горы. А Моисей и Елеазар сошли с горы.
NUM|20|29|И увидело все общество, что Аарон умер, и оплакивал Аарона весь дом Израилев тридцать дней.
NUM|21|1|Ханаанский царь Арада, живущий к югу, услышав, что Израиль идет дорогою от Афарима, вступил в сражение с Израильтянами и несколько из них взял в плен.
NUM|21|2|И дал Израиль обет Господу, и сказал: если предашь народ сей в руки мои, то положу заклятие на города их.
NUM|21|3|Господь услышал голос Израиля и предал Хананеев в руки ему, и он положил заклятие на них и на города их и нарек имя месту тому: Хорма.
NUM|21|4|От горы Ор отправились они путем Чермного моря, чтобы миновать землю Едома. И стал малодушествовать народ на пути,
NUM|21|5|и говорил народ против Бога и против Моисея: зачем вывели вы нас из Египта, чтоб умереть [нам] в пустыне, ибо [здесь] нет ни хлеба, ни воды, и душе нашей опротивела эта негодная пища.
NUM|21|6|И послал Господь на народ ядовитых змеев, которые жалили народ, и умерло множество народа из [сынов] Израилевых.
NUM|21|7|И пришел народ к Моисею и сказал: согрешили мы, что говорили против Господа и против тебя; помолись Господу, чтоб Он удалил от нас змеев. И помолился Моисей о народе.
NUM|21|8|И сказал Господь Моисею: сделай себе змея и выставь его на знамя, и ужаленный, взглянув на него, останется жив.
NUM|21|9|И сделал Моисей медного змея и выставил его на знамя, и когда змей ужалил человека, он, взглянув на медного змея, оставался жив.
NUM|21|10|И отправились сыны Израилевы и остановились в Овофе;
NUM|21|11|и отправились из Овофа и остановились в Ийе–Авариме, в пустыне, что против Моава, к восходу солнца;
NUM|21|12|оттуда отправились, и остановились на долине Заред;
NUM|21|13|отправившись отсюда, остановились у той части Арнона в пустыне, которая течет вне пределов Аморрея, ибо Арнон граница Моава, между Моавом и Аморреем.
NUM|21|14|Потому и сказано в книге браней Господних:
NUM|21|15|Вагеб в Суфе и потоки Арнона, и верховье потоков, которое склоняется к Шебет–Ару и прилегает к пределам Моава.
NUM|21|16|Отсюда [отправились] к Беэр; это тот колодезь, о котором Господь сказал Моисею: собери народ, и дам им воды.
NUM|21|17|Тогда воспел Израиль песнь сию: наполняйся, колодезь, пойте ему;
NUM|21|18|колодезь, который выкопали князья, вырыли вожди народа с законодателем жезлами своими. Из пустыни [отправились] в Матанну,
NUM|21|19|из Матанны в Нагалиил, из Нагалиила в Вамоф,
NUM|21|20|из Вамофа в Гай, который в земле Моава, на вершине [горы] Фасги, обращенной лицем к пустыне.
NUM|21|21|И послал Израиль послов к Сигону, царю Аморрейскому, чтобы сказать:
NUM|21|22|позволь мне пройти землею твоею; не будем заходить в поля и виноградники, не будем пить воды из колодезей [твоих], а пойдем путем царским, доколе не перейдем пределов твоих.
NUM|21|23|Но Сигон не позволил Израилю идти через свои пределы; и собрал Сигон весь народ свой и выступил против Израиля в пустыню, и дошел до Иаацы, и сразился с Израилем.
NUM|21|24|И поразил его Израиль мечом и взял во владение землю его от Арнона до Иавока, до [пределов] Аммонитских, ибо крепок был предел Аммонитян;
NUM|21|25|и взял Израиль все города сии, и жил Израиль во всех городах Аморрейских, в Есевоне и во всех зависящих от него;
NUM|21|26|ибо Есевон был город Сигона, царя Аморрейского, и он воевал с прежним царем Моавитским и взял из руки его всю землю его до Арнона.
NUM|21|27|Потому говорят приточники: идите в Есевон, да устроят и утвердят город Сигона;
NUM|21|28|ибо огонь вышел из Есевона, пламень из города Сигонова, и пожрал Ар–Моав и владеющих высотами Арнона.
NUM|21|29|Горе тебе, Моав! погиб ты, народ Хамоса! Разбежались сыновья его, и дочери его сделались пленницами Аморрейского царя Сигона;
NUM|21|30|мы поразили их стрелами; погиб Есевон до Дивона, мы опустошили их до Нофы, которая близ Медевы.
NUM|21|31|И жил Израиль в земле Аморрейской.
NUM|21|32|И послал Моисей высмотреть Иазер, и взяли селения, зависящие от него, и прогнали Аморреев, которые в них были.
NUM|21|33|И поворотили и пошли к Васану. И выступил против них Ог, царь Васанский, сам и весь народ его, на сражение к Едреи.
NUM|21|34|И сказал Господь Моисею: не бойся его, ибо Я предам его и весь народ его и всю землю его в руки твои, и поступишь с ним, как поступил с Сигоном, царем Аморрейским, который жил в Есевоне.
NUM|21|35|И поразили они его и сынов его и весь народ его, так что ни одного не осталось, и овладели землею его.
NUM|22|1|И отправились сыны Израилевы, и остановились на равнинах Моава, при Иордане, против Иерихона.
NUM|22|2|И видел Валак, сын Сепфоров, все, что сделал Израиль Аморреям;
NUM|22|3|и весьма боялись Моавитяне народа сего, потому что он был многочислен; и устрашились Моавитяне сынов Израилевых.
NUM|22|4|И сказали Моавитяне старейшинам Мадиамским: этот народ поедает теперь все вокруг нас, как вол поедает траву полевую. Валак же, сын Сепфоров, был царем Моавитян в то время.
NUM|22|5|И послал он послов к Валааму, сыну Веорову, в Пефор, который на реке [Евфрате], в земле сынов народа его, чтобы позвать его [и] сказать: вот, народ вышел из Египта и покрыл лице земли, и живет он подле меня;
NUM|22|6|итак приди, прокляни мне народ сей, ибо он сильнее меня: может быть, я тогда буду в состоянии поразить его и выгнать его из земли; я знаю, что кого ты благословишь, тот благословен, и кого ты проклянешь, тот проклят.
NUM|22|7|И пошли старейшины Моавитские и старейшины Мадиамские, с подарками в руках за волхвование, и пришли к Валааму, и пересказали ему слова Валаковы.
NUM|22|8|И сказал он им: переночуйте здесь ночь, и дам вам ответ, как скажет мне Господь. И остались старейшины Моавитские у Валаама.
NUM|22|9|И пришел Бог к Валааму и сказал: какие это люди у тебя?
NUM|22|10|Валаам сказал Богу: Валак, сын Сепфоров, царь Моавитский, прислал [их] ко мне [сказать]:
NUM|22|11|вот, народ вышел из Египта и покрыл лице земли, итак приди, прокляни мне его; может быть я тогда буду в состоянии сразиться с ним и выгнать его.
NUM|22|12|И сказал Бог Валааму: не ходи с ними, не проклинай народа сего, ибо он благословен.
NUM|22|13|И встал Валаам поутру и сказал князьям Валаковым: пойдите в землю вашу, ибо не хочет Господь позволить мне идти с вами.
NUM|22|14|И встали князья Моавитские, и пришли к Валаку, и сказали [ему]: не согласился Валаам идти с нами.
NUM|22|15|Валак послал еще князей, более и знаменитее тех.
NUM|22|16|И пришли они к Валааму и сказали ему: так говорит Валак, сын Сепфоров: не откажись придти ко мне;
NUM|22|17|я окажу тебе великую почесть и сделаю [тебе] все, что ни скажешь мне; приди же, прокляни мне народ сей.
NUM|22|18|И отвечал Валаам и сказал рабам Валаковым: хотя бы Валак давал мне полный свой дом серебра и золота, не могу преступить повеления Господа, Бога моего, и сделать что–либо малое или великое [по своему произволу];
NUM|22|19|впрочем, останьтесь здесь и вы на ночь, и я узнаю, что еще скажет мне Господь.
NUM|22|20|И пришел Бог к Валааму ночью и сказал ему: если люди сии пришли звать тебя, встань, пойди с ними; но только делай то, что Я буду говорить тебе.
NUM|22|21|Валаам встал поутру, оседлал ослицу свою и пошел с князьями Моавитскими.
NUM|22|22|И воспылал гнев Божий за то, что он пошел, и стал Ангел Господень на дороге, чтобы воспрепятствовать ему. Он ехал на ослице своей и с ними двое слуг его.
NUM|22|23|И увидела ослица Ангела Господня, стоящего на дороге с обнаженным мечом в руке, и своротила ослица с дороги, и пошла на поле; а Валаам стал бить ослицу, чтобы возвратить ее на дорогу.
NUM|22|24|И стал Ангел Господень на узкой дороге, между виноградниками, [где] с одной стороны стена и с другой стороны стена.
NUM|22|25|Ослица, увидев Ангела Господня, прижалась к стене и прижала ногу Валаамову к стене; и он опять стал бить ее.
NUM|22|26|Ангел Господень опять перешел и стал в тесном месте, где некуда своротить, ни направо, ни налево.
NUM|22|27|Ослица, увидев Ангела Господня, легла под Валаамом. И воспылал гнев Валаама, и стал он бить ослицу палкою.
NUM|22|28|И отверз Господь уста ослицы, и она сказала Валааму: что я тебе сделала, что ты бьешь меня вот уже третий раз?
NUM|22|29|Валаам сказал ослице: за то, что ты поругалась надо мною; если бы у меня в руке был меч, то я теперь же убил бы тебя.
NUM|22|30|Ослица же сказала Валааму: не я ли твоя ослица, на которой ты ездил сначала до сего дня? имела ли я привычку так поступать с тобою? Он сказал: нет.
NUM|22|31|И открыл Господь глаза Валааму, и увидел он Ангела Господня, стоящего на дороге с обнаженным мечом в руке, и преклонился, и пал на лице свое.
NUM|22|32|И сказал ему Ангел Господень: за что ты бил ослицу твою вот уже три раза? Я вышел, чтобы воспрепятствовать [тебе], потому что путь [твой] не прав предо Мною;
NUM|22|33|и ослица, видев Меня, своротила от Меня вот уже три раза; если бы она не своротила от Меня, то Я убил бы тебя, а ее оставил бы живою.
NUM|22|34|И сказал Валаам Ангелу Господню: согрешил я, ибо не знал, что Ты стоишь против меня на дороге; итак, если это неприятно в очах Твоих, то я возвращусь.
NUM|22|35|И сказал Ангел Господень Валааму: пойди с людьми сими, только говори то, что Я буду говорить тебе. И пошел Валаам с князьями Валаковыми.
NUM|22|36|Валак, услышав, что идет Валаам, вышел навстречу ему в город Моавитский, который на границе при Арноне, что у самого предела.
NUM|22|37|И сказал Валак Валааму: не посылал ли я к тебе, звать тебя? почему ты не шел ко мне? неужели я в самом деле не могу почтить тебя?
NUM|22|38|И сказал Валаам Валаку: вот, я и пришел к тебе, но могу ли я что [от себя] сказать? что вложит Бог в уста мои, то и буду говорить.
NUM|22|39|И пошел Валаам с Валаком и пришли в Кириаф–Хуцоф.
NUM|22|40|И заколол Валак волов и овец, и послал к Валааму и князьям, которые были с ним.
NUM|22|41|На другой день утром Валак взял Валаама и возвел его на высоты Вааловы, чтобы он увидел оттуда часть народа.
NUM|23|1|И сказал Валаам Валаку: построй мне здесь семь жертвенников и приготовь мне семь тельцов и семь овнов.
NUM|23|2|Валак сделал так, как говорил Валаам, и вознесли Валак и Валаам по тельцу и по овну на каждом жертвеннике.
NUM|23|3|И сказал Валаам Валаку: постой у всесожжения твоего, а я пойду; может быть, Господь выйдет мне навстречу, и что Он откроет мне, я объявлю тебе. И пошел на возвышенное место.
NUM|23|4|И встретился Бог с Валаамом, и сказал ему [Валаам]: семь жертвенников устроил я и вознес по тельцу и по овну на каждом жертвеннике.
NUM|23|5|И вложил Господь слово в уста Валаамовы и сказал: возвратись к Валаку и так говори.
NUM|23|6|И возвратился к нему, и вот, он стоит у всесожжения своего, он и все князья Моавитские.
NUM|23|7|И произнес притчу свою и сказал: из Месопотамии привел меня Валак, царь Моава, от гор восточных: приди, прокляни мне Иакова, приди, изреки зло на Израиля!
NUM|23|8|Как прокляну я? Бог не проклинает его. Как изреку зло? Господь не изрекает [на него] зла.
NUM|23|9|С вершины скал вижу я его, и с холмов смотрю на него: вот, народ живет отдельно и между народами не числится.
NUM|23|10|Кто исчислит песок Иакова и число четвертой части Израиля? Да умрет душа моя смертью праведников, и да будет кончина моя, как их!
NUM|23|11|И сказал Валак Валааму: что ты со мною делаешь? я взял тебя, чтобы проклясть врагов моих, а ты, вот, благословляешь?
NUM|23|12|И отвечал он и сказал: не должен ли я в точности сказать то, что влагает Господь в уста мои?
NUM|23|13|И сказал ему Валак: пойди со мною на другое место, с которого ты увидишь его, но только часть его увидишь, а всего его не увидишь; и прокляни мне его оттуда.
NUM|23|14|И взял его на место стражей, на вершину [горы] Фасги, и построил семь жертвенников, и вознес по тельцу и по овну на каждом жертвеннике.
NUM|23|15|И сказал [Валаам] Валаку: постой здесь у всесожжения твоего, а я [пойду] туда навстречу [Богу].
NUM|23|16|И встретился Господь с Валаамом, и вложил слово в уста его, и сказал: возвратись к Валаку и так говори.
NUM|23|17|И пришел к нему, и вот, он стоит у всесожжения своего, и с ним князья Моавитские. И сказал ему Валак: что говорил Господь?
NUM|23|18|Он произнес притчу свою и сказал: встань, Валак, и послушай, внимай мне, сын Сепфоров.
NUM|23|19|Бог не человек, чтоб Ему лгать, и не сын человеческий, чтоб Ему изменяться. Он ли скажет и не сделает? будет говорить и не исполнит?
NUM|23|20|Вот, благословлять начал я, ибо Он благословил, и я не могу изменить сего.
NUM|23|21|Не видно бедствия в Иакове, и не заметно несчастья в Израиле; Господь, Бог его, с ним, и трубный царский звук у него;
NUM|23|22|Бог вывел их из Египта, быстрота единорога у него;
NUM|23|23|нет волшебства в Иакове и нет ворожбы в Израиле. В [свое] время скажут об Иакове и об Израиле: вот что творит Бог!
NUM|23|24|Вот, народ как львица встает и как лев поднимается; не ляжет, пока не съест добычи и не напьется крови убитых.
NUM|23|25|И сказал Валак Валааму: ни клясть не кляни его, ни благословлять не благословляй его.
NUM|23|26|И отвечал Валаам и сказал Валаку: не говорил ли я тебе, что я буду делать все то, что скажет мне Господь?
NUM|23|27|И сказал Валак Валааму: пойди, я возьму тебя на другое место; может быть, угодно будет Богу, и оттуда проклянешь мне его.
NUM|23|28|И взял Валак Валаама на верх Фегора, обращенного к пустыне.
NUM|23|29|И сказал Валаам Валаку: построй мне здесь семь жертвенников и приготовь мне здесь семь тельцов и семь овнов.
NUM|23|30|И сделал Валак, как сказал Валаам, и вознес по тельцу и овну на каждом жертвеннике.
NUM|24|1|Валаам увидел, что Господу угодно благословлять Израиля, и не пошел, как прежде, для волхвования, но обратился лицем своим к пустыне.
NUM|24|2|И взглянул Валаам и увидел Израиля, стоявшего по коленам своим, и был на нем Дух Божий.
NUM|24|3|И произнес он притчу свою и сказал: говорит Валаам, сын Веоров, говорит муж с открытым оком,
NUM|24|4|говорит слышащий слова Божии, который видит видения Всемогущего; падает, но открыты глаза его:
NUM|24|5|как прекрасны шатры твои, Иаков, жилища твои, Израиль!
NUM|24|6|расстилаются они как долины, как сады при реке, как алойные дерева, насажденные Господом, как кедры при водах;
NUM|24|7|польется вода из ведр его, и семя его [будет] как великие воды, превзойдет Агага царь его и возвысится царство его.
NUM|24|8|Бог вывел его из Египта, быстрота единорога у него, пожирает народы, враждебные ему, раздробляет кости их и стрелами своими разит [врага].
NUM|24|9|Преклонился, лежит как лев и как львица, кто поднимет его? Благословляющий тебя благословен, и проклинающий тебя проклят!
NUM|24|10|И воспламенился гнев Валака на Валаама, и всплеснул он руками своими, и сказал Валак Валааму: я призвал тебя проклясть врагов моих, а ты благословляешь их вот уже третий раз;
NUM|24|11|итак, беги в свое место; я хотел почтить тебя, но вот, Господь лишает тебя чести.
NUM|24|12|И сказал Валаам Валаку: не говорил ли я послам твоим, которых ты присылал ко мне:
NUM|24|13|"хотя бы давал мне Валак полный свой дом серебра и золота, не могу преступить повеления Господня, чтобы сделать что–либо доброе или худое по своему произволу: что скажет Господь, то и буду говорить"?
NUM|24|14|Итак, вот, я иду к народу своему; пойди, я возвещу тебе, что сделает народ сей с народом твоим в последствие времени.
NUM|24|15|И произнес притчу свою и сказал: говорит Валаам, сын Веоров, говорит муж с открытым оком,
NUM|24|16|говорит слышащий слова Божии, имеющий ведение от Всевышнего, который видит видения Всемогущего, падает, но открыты очи его.
NUM|24|17|Вижу Его, но ныне еще нет; зрю Его, но не близко. Восходит звезда от Иакова и восстает жезл от Израиля, и разит князей Моава и сокрушает всех сынов Сифовых.
NUM|24|18|Едом будет под владением, Сеир будет под владением врагов своих, а Израиль явит силу [свою].
NUM|24|19|[Происшедший] от Иакова овладеет и погубит оставшееся от города.
NUM|24|20|И увидел он Амалика, и произнес притчу свою, и сказал: первый из народов Амалик, но конец его – гибель.
NUM|24|21|И увидел он Кенеев, и произнес притчу свою, и сказал: крепко жилище твое, и на скале положено гнездо твое;
NUM|24|22|но разорен будет Каин, и недолго до того, что Ассур уведет тебя в плен.
NUM|24|23|И произнес притчу свою, и сказал: горе, кто уцелеет, когда наведет сие Бог!
NUM|24|24|[придут] корабли от Киттима, и смирят Ассура, и смирят Евера; но и им гибель!
NUM|24|25|И встал Валаам и пошел обратно в свое место, а Валак также пошел своею дорогою.
NUM|25|1|И жил Израиль в Ситтиме, и начал народ блудодействовать с дочерями Моава,
NUM|25|2|и приглашали они народ к жертвам богов своих, и ел народ [жертвы их] и кланялся богам их.
NUM|25|3|И прилепился Израиль к Ваал–Фегору. И воспламенился гнев Господень на Израиля.
NUM|25|4|И сказал Господь Моисею: возьми всех начальников народа и повесь их Господу перед солнцем, и отвратится от Израиля ярость гнева Господня.
NUM|25|5|И сказал Моисей судьям Израилевым: убейте каждый людей своих, прилепившихся к Ваал–Фегору.
NUM|25|6|И вот, некто из сынов Израилевых пришел и привел к братьям своим Мадианитянку, в глазах Моисея и в глазах всего общества сынов Израилевых, когда они плакали у входа скинии собрания.
NUM|25|7|Финеес, сын Елеазара, сына Аарона священника, увидев это, встал из среды общества и взял в руку свою копье,
NUM|25|8|и вошел вслед за Израильтянином в спальню и пронзил обоих их, Израильтянина и женщину в чрево ее: и прекратилось поражение сынов Израилевых.
NUM|25|9|Умерших же от поражения было двадцать четыре тысячи.
NUM|25|10|И сказал Господь Моисею, говоря:
NUM|25|11|Финеес, сын Елеазара, сына Аарона священника, отвратил ярость Мою от сынов Израилевых, возревновав по Мне среди их, и Я не истребил сынов Израилевых в ревности Моей;
NUM|25|12|посему скажи: вот, Я даю ему Мой завет мира,
NUM|25|13|и будет он ему и потомству его по нем заветом священства вечного, за то, что он показал ревность по Боге своем и заступил сынов Израилевых.
NUM|25|14|Имя убитого Израильтянина, который убит с Мадианитянкою, было Зимри, сын Салу, начальник поколения Симеонова;
NUM|25|15|а имя убитой Мадианитянки Хазва; она была дочь Цура, начальника Оммофа, племени Мадиамского.
NUM|25|16|И сказал Господь Моисею, говоря:
NUM|25|17|враждуйте с Мадианитянами, и поражайте их,
NUM|25|18|ибо они враждебно поступили с вами в коварстве своем, прельстив вас Фегором и Хазвою, дочерью начальника Мадиамского, сестрою своею, убитою в день поражения за Фегора.
NUM|26|1|После сего поражения сказал Господь Моисею и Елеазару, сыну Аарона, священнику, говоря:
NUM|26|2|исчислите все общество сынов Израилевых от двадцати лет и выше, по семействам их, всех годных для войны у Израиля.
NUM|26|3|И сказал им Моисей и Елеазар священник на равнинах Моавитских у Иордана, против Иерихона, говоря:
NUM|26|4|[исчислите всех] от двадцати лет и выше, как повелел Господь Моисею и сынам Израилевым, которые вышли из земли Египетской:
NUM|26|5|Рувим, первенец Израиля. Сыны Рувима: от Ханоха поколение Ханохово, от Фаллу поколение Фаллуево,
NUM|26|6|от Хецрона поколение Хецроново, от Харми поколение Хармиево;
NUM|26|7|вот поколения Рувимовы; и исчислено их сорок три тысячи семьсот тридцать.
NUM|26|8|И сыны Фаллуя: Елиав.
NUM|26|9|Сыны Елиава: Немуил, Дафан и Авирон. Это те Дафан и Авирон, призываемые в собрание, которые произвели возмущение против Моисея и Аарона вместе с сообщниками Корея, когда сии произвели возмущение против Господа;
NUM|26|10|и разверзла земля уста свои, и поглотила их и Корея; вместе с [ними] умерли и сообщники их, когда огонь пожрал двести пятьдесят человек, и стали они в знамение;
NUM|26|11|но сыны Кореевы не умерли.
NUM|26|12|Сыны Симеона по поколениям их: от Немуила поколение Немуилово, от Ямина поколение Яминово, от Яхина поколение Яхиново,
NUM|26|13|от Зары поколение Зарино, от Саула поколение Саулово;
NUM|26|14|вот поколения Симеоновы: двадцать две тысячи двести.
NUM|26|15|Сыны Гада по поколениям их: от Цефона поколение Цефоново, от Хаггия поколение Хаггиево, от Шуния поколение Шуниево,
NUM|26|16|от Озния поколение Озниево, от Ерия поколение Ериево,
NUM|26|17|от Арода поколение Ародово, от Арелия поколение Арелиево;
NUM|26|18|вот поколения сынов Гадовых, по исчислению их: сорок тысяч пятьсот.
NUM|26|19|Сыны Иуды: Ир и Онан; но Ир и Онан умерли в земле Ханаанской;
NUM|26|20|и были сыны Иуды по поколениям их: от Шелы поколение Шелино, от Фареса поколение Фаресово, от Зары поколение Зарино;
NUM|26|21|и были сыны Фаресовы: от Есрома поколение Есромово, от Хамула поколение Хамулово;
NUM|26|22|вот поколения Иудины, по исчислению их: семьдесят шесть тысяч пятьсот.
NUM|26|23|Сыны Иссахаровы по поколениям их: от Фолы поколение Фолино, от Фувы поколение Фувино,
NUM|26|24|от Иашува поколение Иашувово, от Шимрона поколение Шимроново;
NUM|26|25|вот поколения Иссахаровы, по исчислению их: шестьдесят четыре тысячи триста.
NUM|26|26|Сыны Завулона по поколениям их: от Середа поколение Середово, от Елона поколение Елоново, от Иахлеила поколение Иахлеилово;
NUM|26|27|вот поколения Завулоновы, по исчислению их: шестьдесят тысяч пятьсот.
NUM|26|28|Сыны Иосифа по поколениям их: Манассия и Ефрем.
NUM|26|29|Сыны Манассии: от Махира поколение Махирово; от Махира родился Галаад, от Галаада поколение Галаадово.
NUM|26|30|Вот сыны Галаадовы: от Иезера поколение Иезерово, от Хелека поколение Хелеково,
NUM|26|31|от Асриила поколение Асриилово, от Шехема поколение Шехемово,
NUM|26|32|от Шемиды поколение Шемидино, от Хефера поколение Хеферово.
NUM|26|33|У Салпаада, сына Хеферова, не было сыновей, а только дочери; имя дочерей Салпаадовых: Махла, Ноа, Хогла, Милка и Фирца.
NUM|26|34|Вот поколения Манассиины; а исчислено их пятьдесят две тысячи семьсот.
NUM|26|35|Вот сыны Ефремовы по поколениям их: от Шутелы поколение Шутелино, от Бехера поколение Бехерово, от Тахана поколение Таханово;
NUM|26|36|и вот сыны Шутелы: от Арана поколение Араново;
NUM|26|37|вот поколения сынов Ефремовых, по исчислению их: тридцать две тысячи пятьсот. Вот сыны Иосифовы по поколениям их.
NUM|26|38|Сыны Вениамина по поколениям их: от Белы поколение Белино, от Ашбела поколение Ашбелово, от Ахирама поколение Ахирамово,
NUM|26|39|от Шефуфама поколение Шефуфамово, от Хуфама поколение Хуфамово;
NUM|26|40|и были сыны Белы: Ард и Нааман; [от Арда] поколение Ардово, от Наамана поколение Нааманово;
NUM|26|41|вот сыны Вениамина по поколениям их; а исчислено их сорок пять тысяч шестьсот.
NUM|26|42|Вот сыны Дановы по поколениям их: от Шухама поколение Шухамово; вот семейства Дановы по поколениям их.
NUM|26|43|и всех поколений Шухама, по исчислению их: шестьдесят четыре тысячи четыреста.
NUM|26|44|Сыны Асировы по поколениям их: от Имны поколение Имнино, от Ишвы поколение Ишвино, от Верии поколение Вериино;
NUM|26|45|от сынов Верии, от Хевера поколение Хеверово, от Малхиила поколение Малхиилово;
NUM|26|46|имя дочери Асировой Сара;
NUM|26|47|вот поколения сынов Асировых, по исчислению их: пятьдесят три тысячи четыреста.
NUM|26|48|Сыны Неффалима по поколениям их: от Иахцеила поколение Иахцеилово, от Гуния поколение Гуниево,
NUM|26|49|от Иецера поколение Иецерово, от Шиллема поколение Шиллемово;
NUM|26|50|вот поколения Неффалимовы по поколениям их; исчислено же их сорок пять тысяч четыреста.
NUM|26|51|Вот [число] вошедших в исчисление сынов Израилевых: шестьсот одна тысяча семьсот тридцать.
NUM|26|52|И сказал Господь Моисею, говоря:
NUM|26|53|сим в удел должно разделить землю по числу имен;
NUM|26|54|кто многочисленнее, тем дай удел более; а кто малочисленнее, тем дай удел менее: каждому должно дать удел соразмерно с числом вошедших в исчисление;
NUM|26|55|по жребию должно разделить землю, по именам колен отцов их должны они получить уделы;
NUM|26|56|по жребию должно разделить им уделы их, как многочисленным, так и малочисленным.
NUM|26|57|Сии суть вошедшие в исчисление левиты по поколениям их: от Гирсона поколение Гирсоново, от Каафа поколение Каафово, от Мерари поколение Мерарино.
NUM|26|58|Вот поколения Левиины: поколение Ливниево, поколение Хевроново, поколение Махлиево, поколение Мушиево, поколение Кореево. От Каафа родился Амрам.
NUM|26|59|Имя жены Амрамовой Иохаведа, дочь Левиина, которую родила [жена] Левиина в Египте, а она Амраму родила Аарона, Моисея и Мариам, сестру их.
NUM|26|60|И родились у Аарона Надав и Авиуд, Елеазар и Ифамар;
NUM|26|61|но Надав и Авиуд умерли, когда принесли чуждый огонь пред Господа.
NUM|26|62|И было исчислено двадцать три тысячи всех мужеского пола, от одного месяца и выше; ибо они не были исчислены вместе с сынами Израилевыми, потому что не дано им удела среди сынов Израилевых.
NUM|26|63|Вот исчисленные Моисеем и Елеазаром священником, которые исчисляли сынов Израилевых на равнинах Моавитских у Иордана, против Иерихона;
NUM|26|64|в числе их не было ни одного человека из исчисленных Моисеем и Аароном священником, которые исчисляли сынов Израилевых в пустыне Синайской;
NUM|26|65|ибо Господь сказал им, что умрут они в пустыне, – и не осталось из них никого, кроме Халева, сына Иефонниина, и Иисуса, сына Навина.
NUM|27|1|И пришли дочери Салпаада, сына Хеферова, сына Галаадова, сына Махирова, сына Манассиина из поколения Манассии, сына Иосифова, и вот имена дочерей его: Махла, Ноа, Хогла, Милка и Фирца;
NUM|27|2|и предстали пред Моисея и пред Елеазара священника, и пред князей и пред все общество, у входа скинии собрания, и сказали:
NUM|27|3|отец наш умер в пустыне, и он не был в числе сообщников, собравшихся против Господа со скопищем Кореевым, но за свой грех умер, и сыновей у него не было;
NUM|27|4|за что исчезать имени отца нашего из племени его, потому что нет у него сына? дай нам удел среди братьев отца нашего.
NUM|27|5|И представил Моисей дело их Господу.
NUM|27|6|И сказал Господь Моисею:
NUM|27|7|правду говорят дочери Салпаадовы; дай им наследственный удел среди братьев отца их и передай им удел отца их;
NUM|27|8|и сынам Израилевым объяви и скажи: если кто умрет, не имея у себя сына, то передавайте удел его дочери его;
NUM|27|9|если же нет у него дочери, передавайте удел его братьям его;
NUM|27|10|если же нет у него братьев, отдайте удел его братьям отца его;
NUM|27|11|если же нет братьев отца его, отдайте удел его близкому его родственнику из поколения его, чтоб он наследовал его; и да будет это для сынов Израилевых постановлено в закон, как повелел Господь Моисею.
NUM|27|12|И сказал Господь Моисею: взойди на сию гору Аварим, и посмотри на землю, которую Я даю сынам Израилевым;
NUM|27|13|и когда посмотришь на нее, приложись к народу своему и ты, как приложился Аарон, брат твой;
NUM|27|14|потому что вы не послушались повеления Моего в пустыне Син, во время распри общества, чтоб явить пред глазами их святость Мою при водах [Меривы].
NUM|27|15|И сказал Моисей Господу, говоря:
NUM|27|16|да поставит Господь, Бог духов всякой плоти, над обществом сим человека,
NUM|27|17|который выходил бы пред ними и который входил бы пред ними, который выводил бы их и который приводил бы их, чтобы не осталось общество Господне, как овцы, у которых нет пастыря.
NUM|27|18|И сказал Господь Моисею: возьми себе Иисуса, сына Навина, человека, в котором есть Дух, и возложи на него руку твою,
NUM|27|19|и поставь его пред Елеазаром священником и пред всем обществом, и дай ему наставление пред глазами их,
NUM|27|20|и дай ему от славы твоей, чтобы слушало его все общество сынов Израилевых;
NUM|27|21|и будет он обращаться к Елеазару священнику и спрашивать его о решении, посредством урима пред Господом; и по его слову должны выходить, и по его слову должны входить он и все сыны Израилевы с ним и все общество.
NUM|27|22|И сделал Моисей, как повелел ему Господь, и взял Иисуса, и поставил его пред Елеазаром священником и пред всем обществом;
NUM|27|23|и возложил на него руки свои и дал ему наставление, как говорил Господь чрез Моисея.
NUM|28|1|И сказал Господь Моисею, говоря:
NUM|28|2|повели сынам Израилевым и скажи им: наблюдайте, чтобы приношение Мое, хлеб Мой в жертву Мне, в приятное благоухание Мне, приносимо было Мне в свое время.
NUM|28|3|И скажи им: вот жертва, которую вы должны приносить Господу: два агнца однолетних без порока на день, во всесожжение постоянное;
NUM|28|4|одного агнца приноси утром, а другого агнца приноси вечером;
NUM|28|5|и в приношение хлебное [приноси] десятую часть [ефы] пшеничной муки, смешанной с четвертью гина выбитого елея;
NUM|28|6|это – всесожжение постоянное, какое совершено было при горе Синае, в приятное благоухание, в жертву Господу;
NUM|28|7|и возлияния при ней четверть гина на одного агнца: на святом месте возливай возлияние, вино Господу.
NUM|28|8|Другого агнца приноси вечером, с таким хлебным приношением, как поутру, и с таким же возлиянием при нем приноси его в жертву, в приятное благоухание Господу.
NUM|28|9|А в субботу [приносите] двух агнцев однолетних без порока, и в приношение хлебное две десятых части [ефы] пшеничной муки, смешанной с елеем, и возлияние при нем:
NUM|28|10|это – субботнее всесожжение в каждую субботу, сверх постоянного всесожжения и возлияния при нем.
NUM|28|11|И в новомесячия ваши приносите всесожжение Господу: из крупного скота двух тельцов, одного овна и семь однолетних агнцев без порока,
NUM|28|12|и три десятых части [ефы] пшеничной муки, смешанной с елеем, в приношение хлебное на одного тельца, и две десятых части [ефы] пшеничной муки, смешанной с елеем, в приношение хлебное на овна,
NUM|28|13|и по десятой части [ефы] пшеничной муки, смешанной с елеем, в приношение хлебное на каждого агнца; [это] – всесожжение, приятное благоухание, жертва Господу;
NUM|28|14|и возлияния при них должно быть пол–гина вина на тельца, треть гина на овна и четверть гина на агнца; это всесожжение в каждое новомесячие [во все] месяцы года.
NUM|28|15|И одного козла приносите Господу в жертву за грех; сверх всесожжения постоянного должно приносить его с возлиянием его.
NUM|28|16|В первый месяц, в четырнадцатый день месяца – Пасха Господня.
NUM|28|17|И в пятнадцатый день сего месяца праздник; семь дней должно есть опресноки.
NUM|28|18|В первый день [да будет у вас] священное собрание; никакой работы не работайте;
NUM|28|19|и приносите жертву, всесожжение Господу: из крупного скота двух тельцов, одного овна и семь однолетних агнцев; без порока они должны быть у вас;
NUM|28|20|и при них в приношение хлебное приносите пшеничной муки, смешанной с елеем, три десятых части [ефы] на каждого тельца, и две десятых части [ефы] на овна,
NUM|28|21|и по десятой части [ефы] приноси на каждого из семи агнцев,
NUM|28|22|и одного козла в жертву за грех, для очищения вас;
NUM|28|23|сверх утреннего всесожжения, которое есть всесожжение постоянное, приносите сие.
NUM|28|24|Так приносите и в каждый из семи дней; [это хлеб], жертва, приятное благоухание Господу; сверх всесожжения постоянного и возлияния его, должно приносить [сие].
NUM|28|25|И в седьмой день да будет у вас священное собрание; никакой работы не работайте.
NUM|28|26|И в день первых плодов, когда приносите Господу новое приношение хлебное в седмицы ваши, да будет у вас священное собрание; никакой работы не работайте;
NUM|28|27|и приносите всесожжение в приятное благоухание Господу: из крупного скота двух тельцов, одного овна и семь однолетних агнцев,
NUM|28|28|и при них в приношение хлебное пшеничной муки, смешанной с елеем, три десятых части [ефы] на каждого тельца, две десятых части [ефы] на овна,
NUM|28|29|и по десятой части [ефы] на каждого из семи агнцев,
NUM|28|30|и одного козла [в жертву за грех], для очищения вас;
NUM|28|31|сверх постоянного всесожжения и хлебного приношения при нем, приносите [сие Мне] с возлиянием их; без порока должны быть они у вас.
NUM|29|1|И в седьмой месяц, в первый [день] месяца, да будет у вас священное собрание; никакой работы не работайте; пусть будет [это] у вас день трубного звука;
NUM|29|2|и приносите всесожжение в приятное благоухание Господу: одного тельца, одного овна, семь однолетних агнцев, без порока,
NUM|29|3|и при них в приношение хлебное пшеничной муки, смешанной с елеем, три десятых части [ефы] на тельца, две десятых части [ефы] на овна,
NUM|29|4|и одну десятую часть [ефы] на каждого из семи агнцев,
NUM|29|5|и одного козла в жертву за грех, для очищения вас,
NUM|29|6|сверх новомесячного всесожжения и хлебного приношения его, и [сверх] постоянного всесожжения и хлебного приношения его, и возлияний их, по уставу, в приятное благоухание Господу.
NUM|29|7|И в десятый [день] сего седьмого месяца пусть будет у вас священное собрание: смиряйте [тогда] души ваши и никакого дела не делайте;
NUM|29|8|и приносите всесожжение Господу в приятное благоухание: одного тельца, одного овна, семь однолетних агнцев; без порока пусть будут они у вас;
NUM|29|9|и при них в приношение хлебное пшеничной муки, смешанной с елеем, три десятых части [ефы] на тельца, две десятых части [ефы] на овна,
NUM|29|10|и по десятой части [ефы] на каждого из семи агнцев,
NUM|29|11|и одного козла в жертву за грех, сверх жертвы за грех, [приносимой в день] очищения, и [сверх] всесожжения постоянного и хлебного приношения его, и возлияния их.
NUM|29|12|И в пятнадцатый день седьмого месяца пусть будет у вас священное собрание; никакой работы не работайте и празднуйте праздник Господень семь дней;
NUM|29|13|и приносите всесожжение, жертву, приятное благоухание Господу: тринадцать тельцов, двух овнов, четырнадцать однолетних агнцев; без порока пусть будут они;
NUM|29|14|и при них в приношение хлебное пшеничной муки, смешанной с елеем, три десятых части [ефы] на каждого из тринадцати тельцов, две десятых части [ефы] на каждого из двух овнов,
NUM|29|15|и по десятой части [ефы] на каждого из четырнадцати агнцев,
NUM|29|16|и одного козла в жертву за грех, сверх всесожжения постоянного и хлебного приношения его и возлияния его.
NUM|29|17|И во второй день двенадцать тельцов, двух овнов, четырнадцать однолетних агнцев, без порока,
NUM|29|18|и при них приношение хлебное и возлияние для тельцов, овнов и агнцев, по числу их, по уставу,
NUM|29|19|и одного козла в жертву за грех, сверх всесожжения постоянного и хлебного приношения и возлияния их.
NUM|29|20|И в третий день одиннадцать тельцов, двух овнов, четырнадцать однолетних агнцев, без порока,
NUM|29|21|и при них приношение хлебное и возлияние для тельцов, овнов и агнцев, по числу их, по уставу,
NUM|29|22|и одного козла в жертву за грех, сверх всесожжения постоянного и хлебного приношения и возлияния его.
NUM|29|23|И в четвертый день десять тельцов, двух овнов, четырнадцать однолетних агнцев, без порока,
NUM|29|24|и при них приношение хлебное и возлияние для тельцов, овнов и агнцев, по числу их, по уставу,
NUM|29|25|и одного козла в жертву за грех, сверх всесожжения постоянного и хлебного приношения и возлияния его.
NUM|29|26|И в пятый день девять тельцов, двух овнов, четырнадцать однолетних агнцев, без порока,
NUM|29|27|и при них приношение хлебное и возлияние для тельцов, овнов и агнцев, по числу их, по уставу,
NUM|29|28|и одного козла в жертву за грех, сверх всесожжения постоянного и хлебного приношения и возлияния его.
NUM|29|29|И в шестой день восемь тельцов, двух овнов, четырнадцать однолетних агнцев, без порока,
NUM|29|30|и при них приношение хлебное и возлияние для тельцов, овнов и агнцев, по числу их, по уставу,
NUM|29|31|и одного козла в жертву за грех, сверх всесожжения постоянного и хлебного приношения и возлияния его.
NUM|29|32|И в седьмой день семь тельцов, двух овнов, четырнадцать однолетних агнцев, без порока,
NUM|29|33|и при них приношение хлебное и возлияние для тельцов, овнов и агнцев, по числу их, по уставу,
NUM|29|34|и одного козла в жертву за грех, сверх всесожжения постоянного и хлебного приношения и возлияния его.
NUM|29|35|В восьмой день пусть будет у вас отдание праздника; никакой работы не работайте;
NUM|29|36|и приносите всесожжение, жертву, приятное благоухание Господу: одного тельца, одного овна, семь однолетних агнцев, без порока,
NUM|29|37|и при них приношение хлебное и возлияние для тельца, овна и агнцев по числу их, по уставу,
NUM|29|38|и одного козла в жертву за грех, сверх всесожжения постоянного и приношения хлебного и возлияния его.
NUM|29|39|Приносите это Господу в праздники ваши, сверх [приносимых] вами, по обету или по усердию, всесожжений ваших и хлебных приношений ваших, и возлияний ваших и мирных жертв ваших.
NUM|30|1|И пересказал Моисей сынам Израилевым все, что повелел Господь Моисею.
NUM|30|2|И сказал Моисей начальникам колен сынов Израилевых, говоря: вот что повелел Господь:
NUM|30|3|если кто даст обет Господу, или поклянется клятвою, положив зарок на душу свою, то он не должен нарушать слова своего, но должен исполнить все, что вышло из уст его.
NUM|30|4|Если женщина даст обет Господу и положит [на себя] зарок в доме отца своего, в юности своей,
NUM|30|5|и услышит отец обет ее и зарок, который она положила на душу свою, и промолчит о том отец ее, то все обеты ее состоятся, и всякий зарок ее, который она положила на душу свою, состоится;
NUM|30|6|если же отец ее, услышав, запретит ей, то все обеты ее и зароки, которые она возложила на душу свою, не состоятся, и Господь простит ей, потому что запретил ей отец ее.
NUM|30|7|Если она выйдет в замужество, а на ней обет ее, или слово уст ее, которым она связала себя,
NUM|30|8|и услышит муж ее и, услышав, промолчит: то обеты ее состоятся, и зароки ее, которые она возложила на душу свою, состоятся;
NUM|30|9|если же муж ее, услышав, запретит ей и отвергнет обет ее, который на ней, и слово уст ее, которым она связала себя, [то они не состоятся, и] Господь простит ей.
NUM|30|10|Обет же вдовы и разведенной, какой бы она ни возложила зарок на душу свою, состоится.
NUM|30|11|Если [жена] в доме мужа своего дала обет, или возложила зарок на душу свою с клятвою,
NUM|30|12|и муж ее слышал, и промолчал о том, и не запретил ей, то все обеты ее состоятся, и всякий зарок, который она возложила на душу свою, состоится;
NUM|30|13|если же муж ее, услышав, отвергнул их, то все вышедшие из уст ее обеты ее и зароки души ее не состоятся: муж ее уничтожил их, и Господь простит ей.
NUM|30|14|Всякий обет и всякий клятвенный зарок, чтобы смирить душу, муж ее может утвердить, и муж ее может отвергнуть;
NUM|30|15|если же муж ее молчал о том день за день, то он [тем] утвердил все обеты ее и все зароки ее, которые на ней, утвердил, потому что он, услышав, молчал о том;
NUM|30|16|а если отвергнул их, после того как услышал, то он взял на себя грех ее.
NUM|30|17|Вот уставы, которые Господь заповедал Моисею об отношении между мужем и женою его, между отцом и дочерью его в юности ее, в доме отца ее.
NUM|31|1|И сказал Господь Моисею, говоря:
NUM|31|2|отмсти Мадианитянам за сынов Израилевых, и после отойдешь к народу твоему.
NUM|31|3|И сказал Моисей народу, говоря: вооружите из себя людей на войну, чтобы они пошли против Мадианитян, совершить мщение Господне над Мадианитянами;
NUM|31|4|по тысяче из колена, от всех колен Израилевых пошлите на войну.
NUM|31|5|И выделено из тысяч Израилевых, по тысяче из колена, двенадцать тысяч вооруженных на войну.
NUM|31|6|И послал их Моисей на войну, по тысяче из колена, их и Финееса, сына Елеазара, священника, на войну, и в руке его священные сосуды и трубы для тревоги.
NUM|31|7|И пошли войною на Мадиама, как повелел Господь Моисею, и убили всех мужеского пола;
NUM|31|8|и вместе с убитыми их убили царей Мадиамских: Евия, Рекема, Цура, Хура и Реву, пять царей Мадиамских, и Валаама, сына Веорова, убили мечом;
NUM|31|9|а жен Мадиамских и детей их сыны Израилевы взяли в плен, и весь скот их, и все стада их и все имение их взяли в добычу,
NUM|31|10|и все города их во владениях их и все селения их сожгли огнем;
NUM|31|11|и взяли все захваченное и всю добычу, от человека до скота;
NUM|31|12|и доставили пленных и добычу и захваченное к Моисею и к Елеазару священнику и к обществу сынов Израилевых, к стану, на равнины Моавитские, что у Иордана, против Иерихона.
NUM|31|13|И вышли Моисей и Елеазар священник и все князья общества навстречу им из стана.
NUM|31|14|И прогневался Моисей на военачальников, тысяченачальников и стоначальников, пришедших с войны,
NUM|31|15|и сказал им Моисей: [для чего] вы оставили в живых всех женщин?
NUM|31|16|вот они, по совету Валаамову, были для сынов Израилевых поводом к отступлению от Господа в угождение Фегору, [за что] и поражение было в обществе Господнем;
NUM|31|17|итак убейте всех детей мужеского пола, и всех женщин, познавших мужа на мужеском ложе, убейте;
NUM|31|18|а всех детей женского пола, которые не познали мужеского ложа, оставьте в живых для себя;
NUM|31|19|и пробудьте вне стана семь дней; всякий, убивший человека и прикоснувшийся к убитому, очиститесь в третий день и в седьмой день, вы и пленные ваши;
NUM|31|20|и все одежды, и все кожаные вещи, и все сделанное из козьей [шерсти], и все деревянные сосуды очистите.
NUM|31|21|И сказал Елеазар священник воинам, ходившим на войну: вот постановление закона, который заповедал Господь Моисею:
NUM|31|22|золото, серебро, медь, железо, олово и свинец,
NUM|31|23|и все, что проходит через огонь, проведите через огонь, чтоб оно очистилось, а кроме того и очистительною водою должно очистить; все же, что не проходит через огонь, проведите через воду;
NUM|31|24|и одежды ваши вымойте в седьмой день, и очиститесь, и после того входите в стан.
NUM|31|25|И сказал Господь Моисею, говоря:
NUM|31|26|сочти добычу плена, от человека до скота, ты и Елеазар священник и начальники племен общества;
NUM|31|27|и раздели добычу пополам между воевавшими, ходившими на войну, и между всем обществом;
NUM|31|28|и от воинов, ходивших на войну, возьми дань Господу, по одной душе из пятисот, из людей и из крупного скота, и из ослов и из мелкого скота;
NUM|31|29|возьми это из половины их и отдай Елеазару священнику в возношение Господу;
NUM|31|30|и из половины сынов Израилевых возьми по одной доле из пятидесяти, из людей, из крупного скота, из ослов и из мелкого скота, и отдай это левитам, служащим при скинии Господней.
NUM|31|31|И сделал Моисей и Елеазар священник, как повелел Господь Моисею.
NUM|31|32|И было добычи, оставшейся от захваченного, что захватили бывшие на войне: мелкого скота шестьсот семьдесят пять тысяч,
NUM|31|33|крупного скота семьдесят две тысячи,
NUM|31|34|ослов шестьдесят одна тысяча,
NUM|31|35|людей, женщин, которые не знали мужеского ложа, всех душ тридцать две тысячи.
NUM|31|36|Половина, доля ходивших на войну, по расчислению была: мелкого скота триста тридцать семь тысяч пятьсот,
NUM|31|37|и дань Господу из мелкого скота шестьсот семьдесят пять;
NUM|31|38|крупного скота тридцать шесть тысяч, и дань из них Господу семьдесят два;
NUM|31|39|ослов тридцать тысяч пятьсот, и дань из них Господу шестьдесят один;
NUM|31|40|людей шестнадцать тысяч, и дань из них Господу тридцать две души.
NUM|31|41|И отдал Моисей дань, возношение Господу, Елеазару священнику, как повелел Господь Моисею.
NUM|31|42|И из половины сынов Израилевых, которую отделил Моисей у бывших на войне;
NUM|31|43|половина же [на долю] общества была: мелкого скота триста тридцать семь тысяч пятьсот,
NUM|31|44|крупного скота тридцать шесть тысяч,
NUM|31|45|ослов тридцать тысяч пятьсот,
NUM|31|46|людей шестнадцать тысяч.
NUM|31|47|Из половины сынов Израилевых взял Моисей одну пятидесятую часть из людей и из скота и отдал это левитам, исполняющим службу при скинии Господней, как повелел Господь Моисею.
NUM|31|48|И пришли к Моисею начальники над тысячами войска, тысяченачальники и стоначальники,
NUM|31|49|и сказали Моисею: рабы твои сосчитали воинов, которые нам поручены, и не убыло ни одного из них;
NUM|31|50|и [вот], мы принесли приношение Господу, кто что достал из золотых вещей: цепочки, запястья, перстни, серьги и привески, для очищения душ наших пред Господом.
NUM|31|51|И взял у них Моисей и Елеазар священник золото во всех этих изделиях;
NUM|31|52|и было всего золота, которое принесено в возношение Господу, шестнадцать тысяч семьсот пятьдесят сиклей, от тысяченачальников и стоначальников.
NUM|31|53|Воины грабили каждый для себя.
NUM|31|54|И взял Моисей и Елеазар священник золото от тысяченачальников и стоначальников, и принесли его в скинию собрания, в память сынов Израилевых пред Господом.
NUM|32|1|У сынов Рувимовых и у сынов Гадовых стад было весьма много; и увидели они, что земля Иазер и земля Галаад есть место [годное] для стад;
NUM|32|2|и пришли сыны Гадовы и сыны Рувимовы и сказали Моисею и Елеазару священнику и князьям общества, говоря:
NUM|32|3|Атароф и Дивон, и Иазер, и Нимра, и Есевон, и Елеале, и Севам, и Нево, и Веон,
NUM|32|4|земля, которую Господь поразил пред обществом Израилевым, есть земля [годная] для стад, а у рабов твоих есть стада.
NUM|32|5|И сказали: если мы нашли благоволение в глазах твоих, отдай землю сию рабам твоим во владение; не переводи нас чрез Иордан.
NUM|32|6|И сказал Моисей сынам Гадовым и сынам Рувимовым: братья ваши пойдут на войну, а вы останетесь здесь?
NUM|32|7|для чего вы отвращаете сердце сынов Израилевых от перехода в землю, которую дает им Господь?
NUM|32|8|так поступили отцы ваши, когда я посылал их из Кадес–Варни для обозрения земли:
NUM|32|9|они доходили до долины Есхол, и видели землю, и отвратили сердце сынов Израилевых, чтобы не шли они в землю, которую Господь дает им;
NUM|32|10|и воспылал в тот день гнев Господа, и поклялся Он, говоря:
NUM|32|11|люди сии, вышедшие из Египта, от двадцати лет и выше не увидят земли, о которой Я клялся Аврааму, Исааку и Иакову, потому что они не повиновались Мне,
NUM|32|12|кроме Халева, сына Иефонниина, Кенезеянина, и Иисуса, сына Навина, потому что они повиновались Господу.
NUM|32|13|И воспылал гнев Господа на Израиля, и водил Он их по пустыне сорок лет, доколе не кончился весь род, сделавший зло в очах Господних.
NUM|32|14|И вот, вместо отцов ваших восстали вы, отродье грешников, чтоб усилить еще ярость гнева Господня на Израиля.
NUM|32|15|Если вы отвратитесь от Него, то Он опять оставит его в пустыне, и вы погубите весь народ сей.
NUM|32|16|И подошли они к нему и сказали: мы построим здесь овчие дворы для стад наших и города для детей наших;
NUM|32|17|сами же мы первые вооружимся и пойдем пред сынами Израилевыми, доколе не приведем их в места их; а дети наши пусть останутся в укрепленных городах, [для безопасности] от жителей земли;
NUM|32|18|не возвратимся в домы наши, доколе не вступят сыны Израилевы каждый в удел свой;
NUM|32|19|ибо мы не возьмем с ними удела по ту сторону Иордана и далее, если удел нам достанется по эту сторону Иордана, к востоку.
NUM|32|20|И сказал им Моисей: если вы это сделаете, если вооруженные пойдете на войну пред Господом,
NUM|32|21|и пойдет каждый из вас вооруженный за Иордан пред Господом, доколе не истребит Он врагов Своих пред Собою,
NUM|32|22|и покорена будет земля пред Господом, то после возвратитесь и будете неповинны пред Господом и пред Израилем, и будет земля сия у вас во владении пред Господом;
NUM|32|23|если же не сделаете так, то согрешите пред Господом, и испытаете [наказание] за грех ваш, которое постигнет вас;
NUM|32|24|стройте себе города для детей ваших и дворы для овец ваших и делайте, что произнесено устами вашими.
NUM|32|25|И сказали сыны Гадовы и сыны Рувимовы Моисею: рабы твои сделают, как повелевает господин наш;
NUM|32|26|дети наши, жены наши, стада наши и весь скот наш останутся тут в городах Галаада,
NUM|32|27|а рабы твои, все, вооружившись, как воины, пойдут пред Господом на войну, как говорит господин наш.
NUM|32|28|И дал Моисей о них повеление Елеазару священнику и Иисусу, сыну Навину, и начальникам племен сынов Израилевых,
NUM|32|29|и сказал им Моисей: если сыны Гадовы и сыны Рувимовы перейдут с вами за Иордан, все вооружившись на войну пред Господом, и покорена будет пред вами земля, то отдайте им землю Галаад во владение;
NUM|32|30|если же не пойдут они с вами вооруженные, то они получат владение вместе с вами в земле Ханаанской.
NUM|32|31|И отвечали сыны Гадовы и сыны Рувимовы и сказали: как сказал Господь рабам твоим, так и сделаем;
NUM|32|32|мы пойдем вооруженные пред Господом в землю Ханаанскую, а удел владения нашего пусть будет по эту сторону Иордана.
NUM|32|33|И отдал Моисей им, сынам Гадовым и сынам Рувимовым, и половине колена Манассии, сына Иосифова, царство Сигона, царя Аморрейского, и царство Ога, царя Васанского, землю с городами ее и окрестностями, – города земли во все стороны.
NUM|32|34|И построили сыны Гадовы Дивон и Атароф, и Ароер,
NUM|32|35|и Атароф–Шофан, и Иазер, и Иогбегу,
NUM|32|36|и Беф–Нимру и Беф–Гаран, города укрепленные и дворы для овец.
NUM|32|37|И сыны Рувимовы построили Есевон, Елеале, Кириафаим,
NUM|32|38|и Нево, и Ваал–Меон, которых имена переменены, и Сивму, и дали имена городам, которые они построили.
NUM|32|39|И пошли сыны Махира, сына Манассиина, в Галаад, и взяли его, и выгнали Аморреев, которые были в нем;
NUM|32|40|и отдал Моисей Галаад Махиру, сыну Манассии, и он поселился в нем.
NUM|32|41|И Иаир, сын Манассии, пошел и взял селения их, и назвал их: селения Иаировы.
NUM|32|42|И Новах пошел и взял Кенаф и зависящие от него города, и назвал его своим именем: Новах.
NUM|33|1|Вот станы сынов Израилевых, которые вышли из земли Египетской по ополчениям своим, под начальством Моисея и Аарона.
NUM|33|2|Моисей, по повелению Господню, описал путешествие их по станам их, и вот станы путешествия их:
NUM|33|3|из Раамсеса отправились они в первый месяц, в пятнадцатый день первого месяца; на другой день Пасхи вышли сыны Израилевы под рукою высокою в глазах всего Египта;
NUM|33|4|между тем Египтяне хоронили всех первенцев, которых поразил у них Господь, и над богами их Господь совершил суд.
NUM|33|5|Так отправились сыны Израилевы из Раамсеса и расположились станом в Сокхофе.
NUM|33|6|И отправились из Сокхофа и расположились станом в Ефаме, что на краю пустыни.
NUM|33|7|И отправились из Ефама и обратились к Пи–Гахирофу, что пред Ваал–Цефоном, и расположились станом пред Мигдолом.
NUM|33|8|Отправившись от Гахирофа, прошли среди моря в пустыню, и шли три дня пути пустынею Ефам, и расположились станом в Мерре.
NUM|33|9|И отправились из Мерры и пришли в Елим; в Елиме же [было] двенадцать источников воды и семьдесят финиковых дерев, и расположились там станом.
NUM|33|10|И отправились из Елима и расположились станом у Чермного моря.
NUM|33|11|И отправились от Чермного моря и расположились станом в пустыне Син.
NUM|33|12|И отправились из пустыни Син и расположились станом в Дофке.
NUM|33|13|И отправились из Дофки и расположились станом в Алуше.
NUM|33|14|И отправились из Алуша и расположились станом в Рефидиме, и не было там воды, чтобы пить народу.
NUM|33|15|И отправились из Рефидима и расположились станом в пустыне Синайской.
NUM|33|16|И отправились из пустыни Синайской и расположились станом в Киброт–Гаттааве.
NUM|33|17|И отправились из Киброт–Гаттаавы и расположились станом в Асирофе.
NUM|33|18|И отправились из Асирофа и расположились станом в Рифме.
NUM|33|19|И отправились из Рифмы и расположились станом в Римнон–Фареце.
NUM|33|20|И отправились из Римнон–Фареца и расположились станом в Ливне.
NUM|33|21|И отправились из Ливны и расположились станом в Риссе.
NUM|33|22|И отправились из Риссы и расположились станом в Кегелафе.
NUM|33|23|И отправились из Кегелафы и расположились станом на горе Шафер.
NUM|33|24|И отправились от горы Шафер и расположились станом в Хараде.
NUM|33|25|И отправились из Харады и расположились станом в Макелофе.
NUM|33|26|И отправились из Макелофа и расположились станом в Тахафе.
NUM|33|27|И отправились из Тахафа и расположились станом в Тарахе.
NUM|33|28|И отправились из Тараха и расположились станом в Мифке.
NUM|33|29|И отправились из Мифки и расположились станом в Хашмоне.
NUM|33|30|И отправились из Хашмоны и расположились станом в Мосерофе.
NUM|33|31|И отправились из Мосерофа и расположились станом в Бене–Яакане.
NUM|33|32|И отправились из Бене–Яакана и расположились станом в Хор–Агидгаде.
NUM|33|33|И отправились из Хор–Агидгада и расположились станом в Иотвафе.
NUM|33|34|И отправились от Иотвафы и расположились станом в Авроне.
NUM|33|35|И отправились из Аврона и расположились станом в Ецион–Гавере.
NUM|33|36|И отправились из Ецион–Гавера и расположились станом в пустыне Син. она же Кадес.
NUM|33|37|И отправились из Кадеса и расположились станом на горе Ор, у пределов земли Едомской.
NUM|33|38|И взошел Аарон священник на гору Ор по повелению Господню и умер там в сороковой год по исшествии сынов Израилевых из земли Египетской, в пятый месяц, в первый день месяца;
NUM|33|39|Аарон был ста двадцати трех лет, когда умер на горе Ор.
NUM|33|40|Ханаанский царь Арада, который жил к югу земли Ханаанской, услышал тогда, что идут сыны Израилевы.
NUM|33|41|И отправились они от горы Ор и расположились станом в Салмоне.
NUM|33|42|И отправились из Салмона и расположились станом в Пуноне.
NUM|33|43|И отправились из Пунона и расположились станом в Овофе.
NUM|33|44|И отправились из Овофа и расположились станом в Ийм–Авариме, на пределах Моава.
NUM|33|45|И отправились из Ийма и расположились станом в Дивон–Гаде.
NUM|33|46|И отправились из Дивон–Гада и расположились станом в Алмон–Дивлафаиме.
NUM|33|47|И отправились из Алмон–Дивлафаима и расположились станом на горах Аваримских пред Нево.
NUM|33|48|И отправились от гор Аваримских и расположились станом на равнинах Моавитских у Иордана, против Иерихона;
NUM|33|49|они расположились станом у Иордана от Беф–Иешимофа до Аве–Ситтима на равнинах Моавитских.
NUM|33|50|И сказал Господь Моисею на равнинах Моавитских у Иордана, против Иерихона, говоря:
NUM|33|51|объяви сынам Израилевым и скажи им: когда перейдете через Иордан в землю Ханаанскую,
NUM|33|52|то прогоните от себя всех жителей земли и истребите все изображения их, и всех литых идолов их истребите и все высоты их разорите;
NUM|33|53|и возьмите во владение землю и поселитесь на ней, ибо Я вам даю землю сию во владение;
NUM|33|54|и разделите землю по жребию на уделы племенам вашим: многочисленному дайте удел более, а малочисленному дай удел менее; кому где выйдет жребий, там ему и будет [удел]; по коленам отцов ваших возьмите себе уделы;
NUM|33|55|если же вы не прогоните от себя жителей земли, то оставшиеся из них будут тернами для глаз ваших и иглами для боков ваших и будут теснить вас на земле, в которой вы будете жить,
NUM|33|56|и тогда, что Я вознамерился сделать им, сделаю вам.
NUM|34|1|И сказал Господь Моисею, говоря:
NUM|34|2|дай повеление сынам Израилевым и скажи им: когда войдете в землю Ханаанскую, то вот земля, которая достанется вам в удел, земля Ханаанская с ее границами:
NUM|34|3|южная сторона будет у вас от пустыни Син, подле Едома, и пойдет у вас южная граница от конца Соленого моря с востока,
NUM|34|4|и направится граница на юг к возвышенности Акравима и пойдет через Син, и будут выступы ее на юг к Кадес–Варни, оттуда пойдет к Гацар–Аддару и пройдет через Ацмон;
NUM|34|5|от Ацмона направится граница к потоку Египетскому, и будут выступы ее к морю;
NUM|34|6|а границею западною будет у вас великое море: это будет у вас граница к западу;
NUM|34|7|к северу же будет у вас граница: от великого моря проведите ее к горе Ор,
NUM|34|8|от горы Ор проведите к Емафу, и будут выступы границы к Цедаду;
NUM|34|9|оттуда пойдет граница к Цифрону, и выступы ее будут к Гацар–Енану: это будет у вас граница северная;
NUM|34|10|границу восточную проведите себе от Гацар–Енана к Шефаму,
NUM|34|11|от Шефама пойдет граница к Рибле, с восточной стороны Аина, потом пойдет граница и коснется берегов моря Киннереф с восточной стороны;
NUM|34|12|и пойдет граница к Иордану, и будут выступы ее к Соленому морю. Это будет земля ваша по границам ее со всех сторон.
NUM|34|13|И дал повеление Моисей сынам Израилевым и сказал: вот земля, которую вы разделите на уделы по жребию, которую повелел Господь дать девяти коленам и половине колена;
NUM|34|14|ибо колено сынов Рувимовых по семействам их, и колено сынов Гадовых по семействам их, и половина колена Манассиина получили удел свой:
NUM|34|15|два колена и половина колена получили удел свой за Иорданом против Иерихона к востоку.
NUM|34|16|И сказал Господь Моисею, говоря:
NUM|34|17|вот имена мужей, которые будут делить вам землю: Елеазар священник и Иисус, сын Навин;
NUM|34|18|и по одному князю от колена возьмите для раздела земли.
NUM|34|19|И вот имена сих мужей: для колена Иудина Халев, сын Иефонниин;
NUM|34|20|для колена сынов Симеоновых Самуил, сын Аммиуда;
NUM|34|21|для колена Вениаминова Елидад, сын Кислона;
NUM|34|22|для колена сынов Дановых князь Буккий, сын Иоглии;
NUM|34|23|для сынов Иосифовых, для колена сынов Манассииных князь Ханниил, сын Ефода;
NUM|34|24|для колена сынов Ефремовых князь Кемуил, сын Шифтана;
NUM|34|25|для колена сынов Завулоновых князь Елицафан, сын Фарнака;
NUM|34|26|для колена сынов Иссахаровых князь Фалтиил, сын Аззана;
NUM|34|27|для колена сынов Асировых князь Ахиуд, сын Шеломия;
NUM|34|28|для колена сынов Неффалимовых князь Педаил, сын Аммиуда;
NUM|34|29|вот те, которым повелел Господь разделить уделы сынам Израилевым в земле Ханаанской.
NUM|35|1|И сказал Господь Моисею на равнинах Моавитских у Иордана против Иерихона, говоря:
NUM|35|2|повели сынам Израилевым, чтоб они из уделов владения своего дали левитам города для жительства, и поля при городах со всех сторон дайте левитам:
NUM|35|3|города будут им для жительства, а поля будут для скота их и для имения их и для всех житейских потребностей их;
NUM|35|4|поля при городах, которые вы должны дать левитам, от стены города [должны простираться] на [две] тысячи локтей, во все стороны;
NUM|35|5|и отмерьте за городом к восточной стороне две тысячи локтей, и к южной стороне две тысячи локтей, и к западу две тысячи локтей, и к северной стороне две тысячи локтей, а посредине город: таковы будут у них поля при городах.
NUM|35|6|Из городов, которые вы дадите левитам, [будут] шесть городов для убежища, в которые вы позволите убегать убийце; и сверх их дайте сорок два города:
NUM|35|7|всех городов, которые вы должны дать левитам, [будет] сорок восемь городов, с полями при них.
NUM|35|8|И когда будете давать города из владения сынов Израилевых, тогда из большего дайте более, из меньшего менее; каждое колено, смотря по уделу, какой получит, должно дать из городов своих левитам.
NUM|35|9|И сказал Господь Моисею, говоря:
NUM|35|10|объяви сынам Израилевым и скажи им: когда вы перейдете чрез Иордан в землю Ханаанскую,
NUM|35|11|выберите себе города, которые были бы у вас городами для убежища, куда мог бы убежать убийца, убивший человека неумышленно;
NUM|35|12|и будут у вас города сии убежищем от мстителя, чтобы не был умерщвлен убивший, прежде нежели он предстанет пред общество на суд.
NUM|35|13|Городов же, которые должны вы дать, городов для убежища, должно быть у вас шесть:
NUM|35|14|три города дайте по эту сторону Иордана и три города дайте в земле Ханаанской; городами убежища должны быть они;
NUM|35|15|для сынов Израилевых и для пришельца и для поселенца между вами будут сии шесть городов убежищем, чтобы убегать туда всякому, убившему человека неумышленно.
NUM|35|16|Если кто ударит кого железным орудием так, что тот умрет, то он убийца: убийцу должно предать смерти;
NUM|35|17|и если кто ударит кого из руки камнем, от которого можно умереть, так что тот умрет, то он убийца: убийцу должно предать смерти;
NUM|35|18|или если деревянным орудием, от которого можно умереть, ударит из руки так, что тот умрет, то он убийца: убийцу должно предать смерти;
NUM|35|19|мститель за кровь сам может умертвить убийцу: лишь только встретит его, сам может умертвить его;
NUM|35|20|если кто толкнет кого по ненависти, или с умыслом бросит на него [что–нибудь] так, что тот умрет,
NUM|35|21|или по вражде ударит его рукою так, что тот умрет, то ударившего должно предать смерти: он убийца; мститель за кровь может умертвить убийцу, лишь только встретит его.
NUM|35|22|Если же он толкнет его нечаянно, без вражды, или бросит на него что–нибудь без умысла,
NUM|35|23|или какой–нибудь камень, от которого можно умереть, не видя уронит на него так, что тот умрет, но он не был врагом его и не желал ему зла,
NUM|35|24|то общество должно рассудить между убийцею и мстителем за кровь по сим постановлениям;
NUM|35|25|и должно общество спасти убийцу от руки мстителя за кровь, и должно возвратить его общество в город убежища его, куда он убежал, чтоб он жил там до смерти великого священника, который помазан священным елеем;
NUM|35|26|если же убийца выйдет за предел города убежища, в который он убежал,
NUM|35|27|и найдет его мститель за кровь вне пределов города убежища его, и убьет убийцу сего мститель за кровь, то не будет на нем [вины] кровопролития,
NUM|35|28|ибо тот должен был жить в городе убежища своего до смерти великого священника, а по смерти великого священника должен был возвратиться убийца в землю владения своего.
NUM|35|29|Да будет это у вас постановлением законным в роды ваши, во всех жилищах ваших.
NUM|35|30|Если кто убьет человека, то убийцу должно убить по словам свидетелей; но одного свидетеля недостаточно, [чтобы осудить] на смерть.
NUM|35|31|И не берите выкупа за душу убийцы, который повинен смерти, но его должно предать смерти;
NUM|35|32|и не берите выкупа за убежавшего в город убежища, чтоб ему [позволить] жить в земле [своей] прежде смерти [великого] священника.
NUM|35|33|Не оскверняйте земли, на которой вы [будете жить]; ибо кровь оскверняет землю, и земля не иначе очищается от пролитой на ней крови, как кровью пролившего ее.
NUM|35|34|Не должно осквернять землю, на которой вы живете, среди которой обитаю Я; ибо Я Господь обитаю среди сынов Израилевых.
NUM|36|1|Пришли главы семейств от племени сынов Галаада, сына Махирова, сына Манассиина из племен сынов Иосифовых, и говорили пред Моисеем и пред князьями, главами поколений сынов Израилевых,
NUM|36|2|и сказали: Господь повелел господину нашему дать землю в удел сынам Израилевым по жребию, и господину нашему повелено от Господа дать удел Салпаада, брата нашего, дочерям его;
NUM|36|3|если же они будут женами сынов которого–нибудь [другого] колена сынов Израилевых, то удел их отнимется от удела отцов наших и прибавится к уделу того колена, в котором они будут, и отнимется от доставшегося по жребию удела нашего;
NUM|36|4|и даже когда будет у сынов Израилевых юбилей, тогда удел их прибавится к уделу того колена, в котором они будут, и от удела колена отцов наших отнимется удел их.
NUM|36|5|И дал Моисей повеление сынам Израилевым, по слову Господню, и сказал: правду говорит колено сынов Иосифовых;
NUM|36|6|вот что заповедует Господь о дочерях Салпаадовых: они могут быть женами тех, кто понравится глазам их, только должны быть женами в племени колена отца своего,
NUM|36|7|чтобы удел сынов Израилевых не переходил из колена в колено; ибо каждый из сынов Израилевых должен быть привязан к уделу колена отцов своих;
NUM|36|8|и всякая дочь, наследующая удел в коленах сынов Израилевых, должна быть женою кого–нибудь из племени колена отца своего, чтобы сыны Израилевы наследовали каждый удел отцов своих,
NUM|36|9|и чтобы не переходил удел из колена в другое колено; ибо каждое из колен сынов Израилевых должно быть привязано к своему уделу.
NUM|36|10|Как повелел Господь Моисею, так и сделали дочери Салпаадовы.
NUM|36|11|И вышли дочери Салпаадовы Махла, Фирца, Хогла, Милка и Ноа в замужество за сыновей дядей своих;
NUM|36|12|в племени сынов Манассии, сына Иосифова, они были женами, и остался удел их в колене племени отца их.
NUM|36|13|Сии суть заповеди и постановления, которые дал Господь сынам Израилевым чрез Моисея на равнинах Моавитских, у Иордана, против Иерихона.
