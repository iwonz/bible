1KGS|1|1|А Давид постарів, увійшов у літа. І покривали його одежами, та не було йому тепло.
1KGS|1|2|І сказали йому його раби: Нехай пошукають для пана царя молоду дівчину, і стане вона перед царем, і буде йому за доглядачку. І буде вона лежати при лоні твоїм, і буде тепло панові цареві!
1KGS|1|3|І шукали дівчину вродливу по всій Ізраїлевій границі, та й знайшли шунаммітку Авішаґ, і привели її до царя.
1KGS|1|4|А та дівчина була дуже вродлива. І була вона цареві доглядачкою, і прислуговувала йому, та цар не пізнав її.
1KGS|1|5|А Адонія, син Хаґґітин, бундючився та говорив: Я буду царювати! І справив він собі повоза та верхівців, та п'ятдесят чоловіка бігунів перед собою.
1KGS|1|6|А батько його ніколи його не засмучував, щоб сказати: Чому ти так робиш? А він також був дуже вродливий, і мати народила його по Авесаломі.
1KGS|1|7|І мав він змову з Йоавом, сином Церуї, та зо священиком Евіятаром, і вони помагали Адонії.
1KGS|1|8|А священик Садок, і Беная, син Єгоядин, і пророк Натан, і Шім'ї, і Реї та Давидові лицарі не були з Адонією.
1KGS|1|9|І приніс Адонія в жертву худоби дрібної та худоби великої, та худоби ситої при Евен-Газзохелеті, що при Ен-Роґелі, і закликав усіх братів своїх, царських синів, та всіх Юдиних мужів, царських слуг.
1KGS|1|10|А пророка Натана, і Бенаю, і лицарів та брата свого Соломона він не покликав.
1KGS|1|11|І сказав Натан до Вірсавії, Соломонової матері, говорячи: Чи ти не чула, що зацарював Адонія, син Хаґґітин, а пан наш Давид не знає про те?
1KGS|1|12|А тепер іди, я тобі пораджу, і рятуй життя своє та життя сина свого Соломона!
1KGS|1|13|Іди, і ввійдеш до царя Давида та й скажеш до нього: Чи ж не ти, пане мій царю, присягнув був своїй невільниці, говорячи: Син твій Соломон буде царювати по мені, і він буде сидіти на троні моїм. Чому ж зацарював Адонія?
1KGS|1|14|Ото, ти ще будеш говорити там із царем, а я ввійду за тобою, і потверджу слова твої.
1KGS|1|15|І ввійшла Вірсавія до царя в кімнату, а цар був дуже старий, і шунаммітка Авішаґ послуговувала цареві.
1KGS|1|16|І похилилася Вірсавія, і вклонилася цареві до землі. А цар сказав: Що тобі?
1KGS|1|17|І вона сказала йому: Пане мій, ти присягнув був своїй невільниці Господом, Богом своїм: Соломон, син твій, буде царювати по мені, і він сидітиме на троні моїм.
1KGS|1|18|А тепер ось зацарював Адонія, а ти, пане мій царю, не знаєш про те...
1KGS|1|19|І приніс він у жертву багато волів і худоби ситої та худоби дрібної, і покликав усіх царських синів, і священика Евіятара та Йоава, вождя війська, а раба твого Соломона не покликав.
1KGS|1|20|А ти, пане мій царю, очі всього Ізраїля на тобі, щоб ти сказав їм, хто буде сидіти на троні пана мого царя по ньому.
1KGS|1|21|Інакше станеться, як спочине пан мій цар з батьками своїми, то буду я та син мій Соломон винними.
1KGS|1|22|І ось, ще вона говорила з царем, а прийшов пророк Натан.
1KGS|1|23|І донесли цареві, говорячи: Ось пророк Натан! І ввійшов він перед цареве обличчя і впав перед царем обличчям своїм до землі.
1KGS|1|24|І сказав Натан: Пане мій царю! Чи ти сказав: Адонія буде царювати по мені, і він буде сидіти на троні моїм?
1KGS|1|25|Бо зійшов він сьогодні, і приніс у жертву багато волів і худоби ситої та худоби дрібної. І він покликав усіх царських синів, і провідників війська, і священика Евіятара, і ось вони їдять та п'ють перед ним, і говорять: Нехай живе цар Адонія!
1KGS|1|26|А мене я раб твій! і священика Садока, і Бенаю, сина Єгоядиного, та раба твого Соломона не покликав.
1KGS|1|27|Чи ця річ була від пана мого царя, а ти не повідомив раба свого, хто буде сидіти на троні мого пана царя по ньому?
1KGS|1|28|А цар Давид відповів та й сказав: Покличте мені Вірсавію! І прийшла вона перед царське обличчя, і стала перед царем.
1KGS|1|29|І присягнув цар та й сказав: Як живий Господь, що визволив душу мою від усякого лиха,
1KGS|1|30|як присягнув я тобі Господом, Богом Ізраїля, говорячи: Син твій Соломон буде царювати по мені, і він буде сидіти на моєму троні замість мене, так я й зроблю цього дня!
1KGS|1|31|І вклонилася Вірсавія обличчям своїм до землі, і впала перед царем та й сказала: Нехай живе пан мій, цар Давид, навіки!
1KGS|1|32|І сказав цар Давид: Покличте мені священика Садока, і пророка Натана та Бенаю, сина Єгоядиного. І поприходили вони перед цареве обличчя.
1KGS|1|33|І сказав цар до них: Візьміть із собою слуг вашого пана, і посадіть мого сина Соломона на мою мулицю, і зведіть його до Ґіхону.
1KGS|1|34|А там помаже його священик Садок та пророк Натан на царя над Ізраїлем. І засурміть у сурму та й скрикнете: Нехай живе цар Соломон!
1KGS|1|35|Потім підете за ним, а він увійде та й сяде на моєму троні, і він буде царювати замість мене, і йому наказав я бути володарем над Ізраїлем та над Юдою.
1KGS|1|36|І відповів Беная, син Єгоядин, та й сказав: Амінь. Так нехай скаже Господь, Бог пана мого царя!
1KGS|1|37|Як був Господь із паном моїм царем, так нехай буде з Соломоном, і нехай Він звеличить трон його над трона пана мого царя Давида!
1KGS|1|38|І пішов священик Садок та пророк Натан, і Беная, син Єгоядин, і керетянин, і пелетянин, і посадили Соломона на мулицю царя Давида, та й повели його до Ґіхону.
1KGS|1|39|І взяв священик Садок рога оливи із скинії, та й помазав Соломона. І засурмили в сурму, та й кричав увесь народ: Нехай живе цар Соломон!
1KGS|1|40|І піднявся за ним ввесь народ. А народ грав на сопілках та радів великою радістю, аж земля розпадалася від їхнього голосу!
1KGS|1|41|І почув це Адонія та всі покликані, що були з ним, а вони тількищо скінчили їсти. І почув Йоав голос сурми та й сказав: Що це за крик та гамір у місті?
1KGS|1|42|Ще він говорив, аж ось приходить Йоанатан, син священика Евіятара. А Адонія сказав: Увійди, бо ти муж гідний, і звісти нам щось добре!
1KGS|1|43|І відповів Йонатан та й сказав до Адонії: Таж пан наш цар Давид настановив на царя Соломона!
1KGS|1|44|І послав із ним цар священика Садока та пророка Натана, і Бенаю, Єгоядиного сина, і керетянина, і пелетянина, і вони посадили його на царську мулицю.
1KGS|1|45|І помазали його в Ґіхоні священик Садок та пророк Натан на царя. І повиходили вони звідти веселі, і зашуміло місто. Це той голос, що ви чули.
1KGS|1|46|І Соломон уже засів на троні царства.
1KGS|1|47|І також посходилися царські слуги, щоб поблагословити нашого пана царя Давида, говорячи: Нехай Бог твій учинить Соломонове ім'я славнішим від твого імени, і нехай звеличить його трон над трона твого! І вклонився цар на ложі своїм.
1KGS|1|48|І сказав цар так: Благословенний Господь, Бог Ізраїлів, що сьогодні дав сидячого на моїм троні, а мої очі те бачать!
1KGS|1|49|І затремтіли, і повставали всі покликані, що були з Адонією, і пішли кожен на дорогу свою...
1KGS|1|50|А Адонія боявся Соломона. І встав він, і пішов, і схопився за роги жертівника.
1KGS|1|51|І донесено Соломонові, кажучи: Ось Адонія злякався царя Соломона, й ось він схопився за роги жертівника, кажучи: Нехай цар Соломон зараз присягне мені, що не вб'є свого раба мечем!
1KGS|1|52|І сказав Соломон: Якщо він буде мужем чесним, ані волосина його не впаде на землю! А якщо знайдеться в ньому зло, то помре.
1KGS|1|53|І послав цар Соломон, і відвели його від жертівника. І прийшов він, і впав перед царем Соломоном, а Соломон йому сказав: Іди до свого дому!
1KGS|2|1|І наблизилися Давидові дні до смерти, і він наказав своєму синові Соломонові, говорячи:
1KGS|2|2|Ось я йду дорогою всієї землі, а ти будеш міцний та станеш мужем.
1KGS|2|3|І будеш ти стерегти накази Господа, Бога свого, щоб ходити Його дорогами, щоб стерегти постанови Його, заповіді Його, та устави Його й свідчення Його, як писано в Мойсеєвім Законі, щоб тобі щастило в усьому, що будеш робити, і скрізь, куди звернешся,
1KGS|2|4|щоб виповнив Господь слово Своє, яке говорив мені, кажучи: Якщо сини твої будуть стерегти дороги свої, щоб ходити перед лицем Моїм у правді всім своїм серцем та всією душею своєю, то, сказав: Не буде переводу нікому від тебе на троні Ізраїлевім!
1KGS|2|5|А також ти знаєш, що зробив мені Йоав, син Церуїн, що зробив він двом провідникам Ізраїлевих військ, Авнерові, Неровому синові, та Амасі, синові Єтеровому. Він повбивав їх, і пролив воєнну кров у час миру, і поплямив воєнною кров'ю свого пояса, що на стегнах його, та сандалі свої, що на ногах його.
1KGS|2|6|І ти зробиш за своєю мудрістю, і не даси знизитися сивині його мирно до шеолу.
1KGS|2|7|А синам ґілеадянина Барзіллая зробиш ласку, і нехай вони будуть серед тих, що їдять за твоїм столом, бо вони отак прийшли до мене, коли я втікав перед Авесаломом, твоїм братом.
1KGS|2|8|А ось з тобою Шім'ї, Ґерин син, веніяминівець із Бахуріму. А він прокляв був мене гострим прокляттям того дня, коли я йшов до Маханаїму. Та він прийшов до Йордану стрінути мене, і я присягнув йому Господом, говорячи: Не заб'ю тебе мечем!
1KGS|2|9|А тепер не прощай йому, бо ти муж мудрий, і знатимеш, що зробити йому, і ти сивину його зведеш у крові до шеолу.
1KGS|2|10|І спочив Давид з батьками своїми, і був похований у Давидовім Місті.
1KGS|2|11|А дні, що Давид царював над Ізраїлем, сорок літ: у Хевроні царював він сім літ, а в Єрусалимі царював тридцять і три роки.
1KGS|2|12|І сів Соломон на троні Давида, батька свого, і його царювання було дуже міцне.
1KGS|2|13|І прийшов Адонія, син Гаґґітин, до Вірсавії, Соломонової матері, а вона сказала: Чи прихід твій з миром? І він відказав: З миром.
1KGS|2|14|І сказав: Справа в мене до тебе. А вона відказала: Говори!
1KGS|2|15|І він сказав: Ти знаєш, що моє було це царство, і на мене звернув увесь Ізраїль своє обличчя, щоб мені царювати. Та відійшло царство, і досталось моєму братові, бо від Господа це сталось йому.
1KGS|2|16|А тепер одне бажання жадаю я від тебе: Не відмовляй мені! А вона сказала йому: Говори!
1KGS|2|17|І він сказав: Скажи цареві Соломонові, бо він не відмовить тобі, щоб він дав мені шунаммітку Авішаґ за жінку.
1KGS|2|18|І сказала Вірсавія: Добре, я скажу про тебе цареві.
1KGS|2|19|І прийшла Вірсавія до царя Соломона, щоб сказати йому про Адонія. А цар устав назустріч їй, і вклонився їй, та й сів на своєму троні. І поставив він трона й для царевої матері, і вона сіла по правиці його.
1KGS|2|20|І сказала вона: Одне мале жадання бажаю я від тебе, не відмов мені. І сказав їй цар: Жадай, мати моя, бо я не відмовлю тобі.
1KGS|2|21|І сказала вона: Нехай шунаммітка Авішаґ буде дана братові твоєму Адонії за жінку.
1KGS|2|22|І відповів цар Соломон та й сказав своїй матері: І нащо ти просиш шунаммітку Авішаґ для Адонії? Та попроси для нього й царства, бо він брат мій, старший від мене, і для нього, і для священика Евіятара, і для Йоава, Церуїного сина!...
1KGS|2|23|І присягнув цар Соломон Господом, говорячи: Так нехай зробить мені Бог, і так нехай додасть, коли не на душу свою говорив Адонія це слово...
1KGS|2|24|А тепер, як живий Господь, що міцно поставив мене й посадовив мене на троні мого батька Давида, і що зробив мені дім, як говорив був, сьогодні буде вбитий Адонія!
1KGS|2|25|І послав цар Соломон через Бенаю, Єгоядиного сина, і він уразив його, і той помер...
1KGS|2|26|А священикові Евіятарові цар сказав: Іди до Анатоту на поля свої, бо ти чоловік смерти, а цього дня не вб'ю тебе, бо носив ти ковчега Владики Господа перед обличчям батька мого Давида, і що терпів ти в усьому, в чому терпів мій батько.
1KGS|2|27|І вигнав Соломон Евіятара, щоб не був священиком для Господа, щоб виповнилося слово Господнє, яке говорив у Шіло на дім Іліїв.
1KGS|2|28|А звістка про це прийшла аж до Йоава, бо Йоав схилявся до Адонії, а до Авесалома не схилявся. І втік Йоав до Господньої скинії, і схопився за роги жертівника...
1KGS|2|29|І донесено цареві Соломонові, що Йоав утік до скинії Господньої, і ось він при жертівнику. І послав Соломон Бенаю, Єгоядиного сина, говорячи: Іди, урази його!
1KGS|2|30|І ввійшов Беная до Господньої скинії, та й сказав до нього: Так сказав цар: Вийди! А той відказав: Ні, я тут помру! І передав Беная цареві це слово, говорячи: Так сказав Йоав, і так відповів мені.
1KGS|2|31|І сказав йому цар: Зроби, як я говорив, і врази його. І поховаєш його, і здіймеш невинну кров, що Йоав пролив був, з мене та з дому мого батька.
1KGS|2|32|І нехай оберне Господь його кров на його голову, що він уразив був двох мужів справедливих та ліпших від нього, і повбивав їх мечем, а батько мій Давид того не знав: Авнера, Нериного сина, провідника Ізраїлевого війська, та Амасу, сина Єтеревого, провідника Юдиного війська.
1KGS|2|33|І нехай звернеться їхня кров на голову Йоава та на голову насіння його навіки. А Давидові й насінню його та дому його й трону його нехай буде мир від Господа аж навіки.
1KGS|2|34|І пішов Беная, Єгоядин син, і вразив його, та й убив його. І був він похований у своїм домі в пустині.
1KGS|2|35|А цар, замість нього, настановив над військом Бенаю, Єгоядиного сина, а священика Садока цар настановив замість Евіятара.
1KGS|2|36|І послав цар, і покликав Шім'ї та й сказав йому: Збудуй собі дім в Єрусалимі, й осядеш там, і не вийдеш звідти ані сюди, ані туди.
1KGS|2|37|І буде того дня, як ти вийдеш і перейдеш поток Кедрон, то щоб ти добре знав, що конче помреш. Кров твоя буде на голові твоїй!
1KGS|2|38|І сказав Шім'ї до царя: Добра це річ. Як наказав пан мій цар, так зробить раб твій. І сидів Шім'ї в Єрусалимі багато днів.
1KGS|2|39|І сталося в кінці трьох років, і втекли двоє рабів Шім'ї до Ахіша, Маахіного сина, ґатського царя. І донесли Шім'ї, говорячи: Ось раби твої в Ґаті!
1KGS|2|40|І встав Шім'ї, й осідлав осла свого та й подався до Ахіша, щоб пошукати своїх рабів. І пішов Шім'ї, і привів своїх рабів з Ґату.
1KGS|2|41|А Соломонові донесено, що Шім'ї пішов з Єрусалиму в Ґат і вернувся.
1KGS|2|42|І послав цар, і покликав Шім'ї та й сказав до нього: Чи ж я не заприсяг тебе Господом, і не взяв свідка проти тебе, говорячи: Того дня, коли ти вийдеш і підеш туди чи сюди, щоб ти добре знав, що конче помреш? І ти сказав мені: Добра це річ, що я чув.
1KGS|2|43|І чому ти не додержувався Господньої присяги та наказа, що я наказав був тобі?
1KGS|2|44|І сказав цар до Шім'ї: Ти знаєш усе те зло, і знало твоє серце, що зробив ти Давидові, батькові моєму. І поверне Господь твоє зло на твою голову.
1KGS|2|45|А цар Соломон благословенний, а Давидів трон буде стояти міцно перед Господнім лицем аж навіки.
1KGS|2|46|І цар наказав Бенаї, Єгоядиному синові, і той вийшов і вразив його, і він помер. І царство зміцніло в Соломоновій руці.
1KGS|3|1|І посвоячився Соломон із фараоном, єгипетським царем, і взяв фараонову дочку, і ввів її до Давидового Міста, ще доки він не закінчив будувати свого дому й храму Господнього, та муру навколо Єрусалиму.
1KGS|3|2|Та народ приносив жертви на пагірках, бо не був ще збудований дім для Господнього Імени аж до тих днів.
1KGS|3|3|І полюбив Соломон Господа, щоб ходити постановами свого батька Давида, тільки й він приносив жертви та кадив на пагірках.
1KGS|3|4|І пішов був цар до Ґів'ону, щоб приносити там жертви, бо то найбільший пагірок. Тисячу цілопалень приніс Соломон на тому жертівникові.
1KGS|3|5|У Ґів'оні з'явився Господь до Соломона в нічному сні. І Бог сказав: Проси, що Я маю дати тобі!
1KGS|3|6|А Соломон відказав: Ти зробив був велику милість із рабом Своїм Давидом, батьком моїм, як він ходив перед лицем Твоїм правдою та праведністю, та простотою серця з Тобою. І зберіг Ти йому ту велику милість, і дав йому сина, що сидить на його троні, як є й цього дня.
1KGS|3|7|А тепер, Господи, Боже, Ти вчинив Свого раба царем замість батька мого Давида, а я недоросток, не знаю виходу та входу.
1KGS|3|8|А раб Твій серед народу Твого, якого Ти вибрав, він народ численний, що його не можна ані злічити, ані зрахувати через многоту.
1KGS|3|9|Дай же Своєму рабові серце розумне, щоб судити народ Твій, щоб розрізняти добре від злого, бо хто потрапить керувати цим великим народом Твоїм?
1KGS|3|10|І була та річ приємна в Господніх очах, що Соломон попросив оцю річ.
1KGS|3|11|І сказав Бог до нього: За те, що просив ти цю річ, а не просив для себе днів довгих та багатства, і не просив душ ворогів своїх, а просив собі розуму, щоб уміти судити,
1KGS|3|12|то ось зроблю Я за словом твоїм, ось Я даю тобі серце мудре та розумне, так що такого, як ти, не було перед тобою й не встане такий, як ти, по тобі.
1KGS|3|13|А також те, чого не просив ти, Я даю тобі: і багатство, і славу таку, що такого, як ти, не було перед тобою й не буде нікого серед царів усе життя твоє.
1KGS|3|14|А якщо ти ходитимеш Моїми дорогами, щоб дотримувати постанови Мої та заповіді Мої, як ходив був батько твій Давид, то продовжу дні твої!
1KGS|3|15|І прокинувся Соломон, аж ось це був сон. І ввійшов він до Єрусалиму, та й став перед ковчегом Господнього заповіту, і приніс цілопалення та вчинив жертви мирні. І зробив він гостину для всіх своїх слуг.
1KGS|3|16|І прийшли до царя дві жінки блудниці, та й стали перед обличчям його.
1KGS|3|17|І сказала одна жінка: Прошу, пане мій, я та ця жінка сидимо в одному домі. І породила я при ній у цьому домі.
1KGS|3|18|І сталося третього дня по породі моїм, і породила теж оця жінка. А ми були разом, нікого чужого в домі з нами не було, тільки двоє нас було в домі.
1KGS|3|19|А вночі помер син цієї жінки, бо вона налягла на нього.
1KGS|3|20|І встала вона серед ночі, і взяла мого сина від мене, а невільниця твоя спала, і поклала його при своєму лоні, а свого померлого сина поклала при лоні моїм...
1KGS|3|21|І встала я рано, щоб погодувати сина свого, аж ось помер він! І придивилася я до нього рано, а ото не був це син мій, що я породила...
1KGS|3|22|А інша жінка відказала: Ні, то мій син живий, а твій син мертвий! А та говорила: Ні, то твій син мертвий, а мій син живий! І так сперечались вони перед царем.
1KGS|3|23|І сказав цар: Ця говорить: Це мій син живий, а син твій мертвий, а та говорить: Ні, то син твій мертвий, а мій син живий.
1KGS|3|24|І сказав цар: Подайте мені меча! І принесли меча перед цареве обличчя.
1KGS|3|25|І сказав цар: Розітніть це живе дитя надвоє, і дайте половину одній, а половину другій!...
1KGS|3|26|І сказала до царя жінка, що син її той живий, бо запалилася любов її до сина свого, і сказала вона: Прошу, пане мій, дайте їй немовлятко живим, а забити не забивайте його!... А та каже: Хай не буде ні мені, ні тобі, розтинайте!...
1KGS|3|27|А цар відповів та й сказав: Дайте їй це живе немовлятко, а вбивати не вбивайте його. Вона його мати!
1KGS|3|28|І почув увесь Єрусалим про той суд, що цар розсудив, і стали боятися царя, бо бачили, що в ньому Божа мудрість, щоб чинити суд.
1KGS|4|1|І був цар Соломон царем над усім Ізраїлем.
1KGS|4|2|А оце його провідники: Азарія, Садоків син, священик.
1KGS|4|3|Еліхореф та Ахійя, сини Шіші, писарі. Йосафат, син Ахілудів, канцлер.
1KGS|4|4|А Беная, Єгоядин син, над військом, а Садок та Евіятар священики.
1KGS|4|5|А Азарія, Натанів син, над намісниками, а Завуд, син Натанів священик, товариш царів.
1KGS|4|6|А Ахішар над домом, а Адонірам, Авдин син над даниною.
1KGS|4|7|А в Соломона було дванадцять намісників над усім Ізраїлем, і вони годували царя та дім його, місяць на рік був на одного на годування.
1KGS|4|8|А оце їхні імена: Бен-Гур в Єфремових горах,
1KGS|4|9|Бен-Декер у Макаці, і в Шаалевімі, і в Бет-Шемеші, і в Елоні Бет-Ганану.
1KGS|4|10|Бен-Гесед в Арубботі, йому належали: Сохо та ввесь край Хеферу.
1KGS|4|11|Бен-Авінадав уся околиця Дору; Тафат, Соломонова дочка, була йому за жінку.
1KGS|4|12|Баана, Ахілудів син Таанах і Меґіддо та ввесь Бет-Шеан, що при Цартані, нижче Їзреелу, від Бет-Шеану аж до Авел-Мехола, аж до того боку Йокмеаму.
1KGS|4|13|Бен-Ґевер у ґілеадському Рамоті, йому належали: оселі Яїра, сина Манасії, що в Ґілеаді, йому околиця Арґову, що в Башані, шістдесят міст великих, із муром та з мідяним засувом.
1KGS|4|14|Ахінадав, син Іддо в Маханаїмі.
1KGS|4|15|Ахімаац в Нефталимі; також він узяв Босмат, Соломонову дочку, за жінку.
1KGS|4|16|Баана, Хушаїв син, в Асирі та в Бе-Алоті.
1KGS|4|17|Йосафат, Паруахів син, в Іссахарі.
1KGS|4|18|Шім'ї, Елин син, у Веніямині.
1KGS|4|19|Ґевер, син Уріїв, у ґілеадському краї, у краї Сигона, царя аморейського, та Оґа, царя башанського. А один намісник, що в усьому Краї.
1KGS|4|20|Юда та Ізраїль були численні, як пісок, що над морем, щодо многоти. Вони їли й пили та тішилися!
1KGS|4|21|(5-1) А Соломон панував над усіма царствами від Річки аж до филистимського краю та аж до границі Єгипту. Вони приносили дари та служили Соломонові по всі дні його життя.
1KGS|4|22|(5-2) І була Соломонова пожива на один день: тридцять корів пшеничної муки, а шістдесят корів іншої муки.
1KGS|4|23|(5-3) Десятеро з великої ситої худоби, і двадцятеро з худоби великої з паші та сотня худоби дрібної, окрім оленя, і сарни, і антилопи та ситих гусок.
1KGS|4|24|(5-4) Бо він панував по всій цій стороні Річки від Тіфсаху та аж до Аззи над усіма царями по цей бік Річки. І був у нього мир зо всіх сторін його навколо.
1KGS|4|25|(5-5) І безпечно сидів Юда та Ізраїль, кожен під своїм виноградником та під своєю фіґою від Дану й аж до Беер-Шеви всі дні Соломона.
1KGS|4|26|(5-6) І було в Соломона сорок тисяч стійлів для коней колесниць його та дванадцять тисяч верхівців.
1KGS|4|27|(5-7) І годували ці намісники царя Соломона та кожного, хто приходив до столу царя Соломона, кожен свій місяць, і не було недостачі ні в чому.
1KGS|4|28|(5-8) А ячменю та соломи для коней та для румаків спроваджували до місця, де хто був, кожен за постановою для нього.
1KGS|4|29|(5-9) І дав Бог Соломонові дуже багато мудрости та розуму, а широкість серця як пісок, що на березі моря.
1KGS|4|30|(5-10) І збільшилася Соломонова мудрість над мудрість усіх синів сходу та над усю мудрість Єгипту.
1KGS|4|31|(5-11) І був він мудріший від усякого чоловіка, від Етана езрахітського, і Гемана, і Калкола та Дарди, Махолових синів. А ім'я його було славне серед усіх людей навколо.
1KGS|4|32|(5-12) І він проказав три тисячі приказок, а пісень його було тисяча й п'ять.
1KGS|4|33|(5-13) І говорив він про дерева, від кедру, що на Ливані, й аж до ісопу, що росте на стіні. І говорив про худобу, і про птаства, і про плазуюче та про риб.
1KGS|4|34|(5-14) І приходили від усіх народів, щоб послухати Соломонову мудрість, від усіх царів краю, що чули про мудрість його.
1KGS|5|1|(5-15) І послав Хірам, цар Тиру, своїх слуг до Соломона, бо почув, що його помазали на царя на місце батька його, бо Хірам був приятелем Давидовим по всі дні.
1KGS|5|2|(5-16) І послав Соломон до Хірама, говорячи:
1KGS|5|3|(5-17) Ти знаєш мого батька Давида, що не міг він збудувати дому для Імени Господа, Бога свого, через війни, що оточували його, аж поки Господь не віддав їх, ворогів, під стопи ніг його.
1KGS|5|4|(5-18) А тепер Господь, Бог мій, дав мені відпочинок навколо, нема противника, і нема злого випадку.
1KGS|5|5|(5-19) І ото я маю на думці збудувати дім Імени Господа, Бога мого, як Господь говорив був моєму батькові Давидові, кажучи: Син твій, якого дам замість тебе на трон твій, він збудує той дім для Ймення Мого.
1KGS|5|6|(5-20) А тепер накажи, і нехай зітнуть мені кедри з Ливану, а раби мої будуть із рабами твоїми, а в нагороду за твоїх рабів я дам тобі все, що скажеш, бо ти знаєш, що серед нас немає нікого, хто вмів би стинати дерева, як сидоняни.
1KGS|5|7|(5-21) І сталося, як почув Хірам Соломонові слова, то дуже зрадів та й сказав: Благословенний Господь сьогодні, що дав Давидові мудрого сина над цим великим народом!
1KGS|5|8|(5-22) І послав Хірам до Соломона, говорячи: Почув я про те, про що посилав ти до мене. Я виконаю все бажання твоє, щодо дерева кедрового та дерева кипарисового.
1KGS|5|9|(5-23) Мої раби спустять із Ливану до моря, а я їх поскладаю в плоти, і відправлю морем аж до місця, про яке пошлеш мені звістку, і порозбиваю їх там, і ти забереш. А ти виконаєш моє бажання, дати хліба для мого дому.
1KGS|5|10|(5-24) І давав Хірам Соломонові дерева кедрові та дерева кипарисові, усе за бажанням його.
1KGS|5|11|(5-25) А Соломон давав Хірамові двадцять тисяч корів пшениці, живність для дому його, та двадцять тисяч корів товченої оливи. Так давав Соломон Хірамові рік-у-рік.
1KGS|5|12|(5-26) А Господь дав Соломонові мудрість, як обіцяв був йому. І був мир між Хірамом та між Соломоном, і обидва вони склали умову.
1KGS|5|13|(5-27) А Соломон зібрав данину робітників зо всього Ізраїля, і була та данина тридцять тисяч чоловіка.
1KGS|5|14|(5-28) І він посилав їх до Ливану, по десять тисяч на місяць, напереміну: місяць були вони на Ливані, два місяці у домі своїм; а Адонірам доглядав над робітниками.
1KGS|5|15|(5-29) І було в Соломона сімдесят тисяч тягарових носіїв та вісімдесят тисяч ламачів у горах,
1KGS|5|16|(5-30) окрім трьох тисяч і трьох сотень керівників, що настановив Соломон над працею, вони правили над народом, що робили працю.
1KGS|5|17|(5-31) І цар наказав, і вони ламали велике каміння, каміння дороге, щоб закласти дім із тесаного каміння.
1KGS|5|18|(5-32) І їх отесували будівничі Соломонові й будівничі Хірамові та ґівляни, і наготовили дерева та каміння на збудування храму.
1KGS|6|1|І сталося, року чотирисотого й вісімдесятого по виході Ізраїлевих синів з єгипетського краю, четвертого року Соломонового царювання над Ізраїлем, місяця зіва, почав він будувати той храм для Господа.
1KGS|6|2|А той храм, що цар Соломон збудував для Господа, шістдесят ліктів довжина його, а двадцять ширина його, а тридцять ліктів вишина його.
1KGS|6|3|А притвор перед храмом цього дому двадцять ліктів довжина його, відповідно широкости храму, десять ліктів ширина його перед храмом.
1KGS|6|4|І зробив він для храму прозорі вікна, широкі знадвору й вузькі всередині.
1KGS|6|5|А до стіни храму збудував він прибудівку навколо, зо стінами дому навколо храму та найсвятішого, і поробив бічні кімнати навколо.
1KGS|6|6|Долішня прибудівка ширина її п'ять ліктів, а середня шість ліктів ширина її, а третя сім ліктів ширина її, бо він дав навколо храму знадвору виступи, щоб не тримати їх у стінах храму.
1KGS|6|7|А храм, коли був будований, будувався з викінченого каменя з каменоломні, а молотки та сокира, всяке залізне знаряддя не було чуте в храмі, коли його будували.
1KGS|6|8|Вхід до середньої бічної кімнати був з правого боку храму, а крученими сходами входили до середньої, а з середньої до третьої.
1KGS|6|9|І збудував він той храм та й покінчив його. І покрив він храм дошками та брусками кедрових дерев.
1KGS|6|10|І збудував він прибудівку на ввесь храм, п'ять ліктів вишина її, і вона трималася храму кедровими деревинами.
1KGS|6|11|І було Господнє слово до Соломона, говорячи:
1KGS|6|12|Цей храм, що ти будуєш, якщо ти ходитимеш Моїми уставами й постанови Мої будеш виконувати, і будеш дотримувати всі Мої заповіді, щоб ними ходити, то Я виповню на тобі Своє слово, яке Я говорив був батькові твоєму Давидові.
1KGS|6|13|І пробуватиму посеред Ізраїлевих синів, і не покину Свого Ізраїлевого народу.
1KGS|6|14|І збудував Соломон той храм та й скінчив його.
1KGS|6|15|І побудував він стіни храму зсередини з кедрових дощок, від підлоги храму аж до стін стропу покрив усередині деревом, а підлогу храму покрив кипарисовими дошками.
1KGS|6|16|І збудував тих двадцять ліктів стіни з-заду храму з кедрових дощок, від підлоги аж до стін стропу, і це збудував йому зсередини за девіра, за Святеє Святих.
1KGS|6|17|А той храм був на сорок ліктів, він той, що перед девіром.
1KGS|6|18|А на кедрині всередині храму була різьба огірків та відкритих квітів. Усе кедрина, камінь був невидний.
1KGS|6|19|А найсвятіше він приготовив усередині храму, щоб дати туди ковчега Господнього заповіту.
1KGS|6|20|А середина найсвятішого двадцять ліктів довжина, і двадцять ліктів ширина, і двадцять ліктів вишина його, і він покрив його щирим золотом, і також покрив кедрового жертівника.
1KGS|6|21|І Соломон покрив той храм зсередини щирим золотом, а перед найсвятішим перетягнув золотими ланцюгами, та покрив його золотом.
1KGS|6|22|І ввесь храм він покрив золотом аж до кінця всього храму і всього жертівника, що при найсвятішому, покрив золотом.
1KGS|6|23|І зробив у найсвятішому двох херувимів з оливкового дерева, десять ліктів вишина його.
1KGS|6|24|І п'ять ліктів одне крило херувима, і п'ять ліктів друге крило херувима; десять ліктів від кінця одного його крила і аж до кінця другого його крила.
1KGS|6|25|І десять ліктів був і другий херувим, одна міра й один вид обом херувимам.
1KGS|6|26|Височина одного херувима десять ліктів, і так і другого херувима.
1KGS|6|27|І дав він тих херувимів усередині внутрішнього храму. І херувими простягали свої крила, і торкалося крило одного однієї стіни, а крило другого херувима торкалося другої стіни. А їхні внутрішні крила дотикалися крило до крила.
1KGS|6|28|І він покрив херувимів золотом.
1KGS|6|29|А всі стіни храму навколо приоздобив ритими різьбами херувимів і пальм та розкритих квітів, зсередини та від зовнішньої частини.
1KGS|6|30|А підлогу храму він покрив золотом для внутрішньої та для зовнішньої частини.
1KGS|6|31|А на вхід до найсвятішого зробив двері з оливкового дерева; стовп, бічні одвірки п'ятикутні.
1KGS|6|32|І двоє дверей були з оливкового дерева, і на них були пороблені різьби херувимів і пальм та розкритих квітів, і покрив золотом; і обклав золотом тих херувимів та ті пальми.
1KGS|6|33|І так поробив і одвірки для входу до храму, з оливкового дерева, одвірки чотирикутні.
1KGS|6|34|А двоє дверей були з кипарисового дерева. Дві частині одних дверей та дві частині других дверей були рухомі.
1KGS|6|35|І повирізував на них херувимів і пальми та розкриті квіти, і покрив золотом, викутим по різьбі.
1KGS|6|36|І збудував він унутрішній двір, три ряди тесаного каменя та ряд стятого кедрового брусся.
1KGS|6|37|Року четвертого був заложений храм Господній, у місяці зів,
1KGS|6|38|а року одинадцятого, у місяці бул, він місяць восьмий був закінчений той храм зо всіма речами його та за всіма планами його. І він будував його сім років.
1KGS|7|1|А свій дім Соломон будував тринадцять років, та й скінчив увесь свій дім.
1KGS|7|2|І збудував він дім Ливанського Лісу, сто ліктів довжина його, і п'ятдесят ліктів ширина його, і тридцять ліктів вишина його, на чотирьох рядах кедрових стовпів, а кедрові брусся на стовпах.
1KGS|7|3|І покритий він був кедриною зверху на бічних кімнатах, що на сорока й п'яти стовпах, по п'ятнадцять на ряд.
1KGS|7|4|А лутків було три ряди, вікно до вікна три рази.
1KGS|7|5|А всі двері та бічні одвірки чотирикутні, з порогами, а навпроти вікно до вікна три рази.
1KGS|7|6|І зробив він сіни зо стовпів, п'ятдесят ліктів довжина їх та тридцять ліктів ширина їх, і інші сіни перед ними, і стовпи, і причілок даху.
1KGS|7|7|І зробив він тронову залю, де судив, залю судову, і покрив кедриною від підлоги до стелі.
1KGS|7|8|А його дім, де жив, на іншому дворі, зсередини сіней, був такий, як та робота. І зробив він дім для фараонової дочки, яку взяв Соломон, як ті сіни.
1KGS|7|9|Усе це з дорогого каміння, тесаного за мірою, обрізаного пилкою зсередини та іззовні, і від основи аж до стелі, а іззовні аж до великого двора.
1KGS|7|10|А заснований він був на дорогих каміннях, каміннях великих, каміння десяти ліктів та каміння восьми ліктів.
1KGS|7|11|А згори дорогі каміння, тесані за мірою, та кедрина.
1KGS|7|12|А навколо великий двір, три ряди тесаного каміння та ряд стятого кедрового брусся; те саме й для внутрішнього двору Господнього храму та для сіней храму.
1KGS|7|13|І послав цар Соломон, і взяв із Тиру Хірама,
1KGS|7|14|це син однієї вдови, з племени Нефталимового, а батько його тирянин, що робив на міді. І був він наповнений мудрістю й розумом, та вмінням робити всяку роботу на міді. І прийшов він до царя Соломона, і зробив усю його роботу.
1KGS|7|15|І він відлив два мідяні стовпи, вісімнадцять ліктів височина одного стовпа, а шнур дванадцяти ліктів оточив би його; такий і стовп другий.
1KGS|7|16|І зробив він дві маковиці, щоб дати на верхи тих стовпів, відлив їх із міді; п'ять ліктів височина однієї маковиці, і п'ять ліктів височина маковиці другої.
1KGS|7|17|А на тих маковицях, що були на верхах стовпів, було мереживо плетеної роботи та шнурки роботою ланцюжків, сім на маковиці одній і сім на маковиці другій.
1KGS|7|18|І поробив він ті стовпи так, що два ряди гранатових яблук були навколо на одному мереживі, щоб покрити маковиці, що на верху; і так зробив і маковиці другій.
1KGS|7|19|А маковиці, що на верху тих стовпів, були зроблені як лілеї, на чотири лікті, у притворі.
1KGS|7|20|І маковиці на обох стовпах також зверху, навпроти випуклини, що з боку мережива. А тих гранатових яблук двісті, рядами навколо на маковиці другій.
1KGS|7|21|І поставив він ті стовпи до притвору храму. І поставив він правого стовпа, і назвав ім'я йому: Яхін; і поставив стовпа лівого, і назвав ім'я йому: Боаз.
1KGS|7|22|А на верху стовпів зроблено як лілеї. І була скінчена робота стовпів.
1KGS|7|23|І зробив він лите море, десять ліктів від краю його аж до краю його, навколо круглясте, і п'ять ліктів височина його. А шнур на тридцять ліктів оточив би його навколо.
1KGS|7|24|А здолу на краях його оточували його подоби огірків, по десять у лікті, вони оточували море навколо. Було два ряди тих огірків, вилитих при литті його.
1KGS|7|25|Воно стояло на дванадцятьох волах, три обернені на північ, і три обернені на захід, і три обернені на південь, і три обернені на схід. А море на них зверху, а ввесь зад їх до нутра.
1KGS|7|26|А грубина його долоня, а краї його подібні до краю келиха, як квітки лілеї. Містило воно дві тисячі батів.
1KGS|7|27|І зробив він десять мідяних підстав, чотири лікті довжина однієї підстави, і чотири лікті ширина її, а три лікті вишина її.
1KGS|7|28|А оце робота підстави: у них лиштви, а ті лиштви поміж прутами.
1KGS|7|29|А на лиштвах, що між прутами, леви, воли та херувими. А на прутах зверху підніжки, а під левами та волами китиці, зроблені розложистими.
1KGS|7|30|І чотири мідяні кола для однієї підстави та мідяні осі. А на чотирьох рогах їхні рамена, під мідницею рамена литі, з кожного боку китиці.
1KGS|7|31|А гирло його з нутра маковиці й вище лікоть; а гирло круглясте, роботи підніжка, лікоть і півліктя; і також на гирлі його різьби, а рамено їх квадратове, не круглясте.
1KGS|7|32|І чотири ті кола були під лиштвами, а осі колес у підставі. А вишина одного кола лікоть і півліктя.
1KGS|7|33|А робота тих кіл як робота кола возового; їхні осі, і їхні обіддя, і їхні шпиці, і їхні маточини усе лите.
1KGS|7|34|І чотири рамена на чотирьох рогах однієї підстави; з підстави виходили рамена її.
1KGS|7|35|А на верху підстави було округле навкілля, півліктя вишини; а на верху підстави ручки її та лиштви її з неї.
1KGS|7|36|І він повирізував на таблицях ручок її та на лиштвах її херувимів левів та пальми, на кожнім вільнім місці, та китиці навколо.
1KGS|7|37|Як це, він зробив десять підстав, лиття одне, міра одна, одна робота для них усіх.
1KGS|7|38|І зробив він десять мідяних умивальниць, сорок батів мала кожна вмивальниця; чотири лікті кожна вмивальниця; одна вмивальниця на одній підставі, так для десяти підстав.
1KGS|7|39|І дав ті підстави п'ять на боці храму з правиці, і п'ять на боці храму з лівиці його, а море дав на правому боці храму, наперед, навпроти полудня.
1KGS|7|40|І поробив Хірам умивальниці й лопатки та кропильниці. І покінчив Хірам робити всю ту роботу, що зробив цареві Соломонові для храму Господнього:
1KGS|7|41|два стовпи та дві голівки маковиць, що на верху стовпів, і два мережива на покриття двох голівок маковиць, що на верху стовпів;
1KGS|7|42|і чотири сотні гранатових яблук для двох мережив, два ряди гранатових яблук для одного мережива, на покриття обох голівок маковиць, що на верху стовпів;
1KGS|7|43|і підстави десять, і вмивальниці десять;
1KGS|7|44|і одне море, і воли дванадцять під морем;
1KGS|7|45|і горнята, і лопатки, і кропильниці та всі ті речі, що Хірам поробив цареві Соломонові в Господньому домі, усе виполірувана мідь.
1KGS|7|46|На Йорданській рівнині повідливав їх цар у глибокій землі між Суккотом та між Царетаном.
1KGS|7|47|І порозставляв Соломон усі ці речі; через дуже велику многоту їх не була справджена вага міді.
1KGS|7|48|І поробив Соломон усі речі, що в Господньому храмі: золотого жертівника, і золотого стола, що на ньому хліб показний,
1KGS|7|49|і свічники, п'ять з правиці та п'ять з лівиці, перед найсвятішим, зо щирого золота; і квітки, і лямпади, і щипчики, з золота;
1KGS|7|50|і миски, і ножиці, і кропильниці, і ложки, і лопатки, золото щире; і чопи для дверей внутрішнього храму, для Святого Святих, для дверей дому для храму золото.
1KGS|7|51|І була покінчена вся ця праця, яку цар Соломон зробив в Господньому храмі. І Соломон повносив освячені речі свого батька Давида; срібло й золото та речі дав у скарбниці Господнього храму.
1KGS|8|1|Тоді Соломон зібрав усіх Ізраїлевих старших та голів племен, керівників батьківських домів Ізраїлевих синів, до царя Соломона до Єрусалиму, щоб перенести ковчега Господнього заповіту з Давидового Міста, воно Сіон.
1KGS|8|2|І були зібрані до царя Соломона всі ізраїльтяни в свято в місяці етанім, він місяць сьомий.
1KGS|8|3|І поприходили всі Ізраїлеві старші, а священики понесли ковчега.
1KGS|8|4|І понесли вони Господнього ковчега, і скинію заповіту та всі святі речі, що в ковчезі; і понесли їх священики та Левити.
1KGS|8|5|А цар Соломон та вся Ізраїлева громада, що зібралися при ньому, були з ним перед ковчегом, і приносили в жертву худобу дрібну та худобу велику, що через многість не була вона ані записувана, ані лічена.
1KGS|8|6|І внесли священики ковчега Господнього заповіту до девіру храму, до Святого Святих, під крила херувимів.
1KGS|8|7|Бо херувими простягали крила над місцем ковчегу, і затінювали херувими над ковчегом та над його держаками зверху.
1KGS|8|8|А ті держаки були довгі, і головки тих держаків були видні з святині перед найсвятішим, а зназовні не були видні. І вони там аж до цього дня.
1KGS|8|9|У ковчезі не було нічого, тільки дві камінні таблиці, що поклав туди Мойсей на Хориві, коли Господь склав був заповіта з Ізраїлевими синами при виході їх з єгипетського краю.
1KGS|8|10|І сталося, як священики виходили з святині, то хмара наповнила Господній храм.
1KGS|8|11|І не могли священики стояти й служити через ту хмару, бо слава Господня наповнила Господній храм!
1KGS|8|12|Тоді Соломон проказав: Промовив Господь, що Він пробуватиме в мряці.
1KGS|8|13|Будуючи, я збудував оцей храм, на оселю Тобі, місце Твого пробування навіки!
1KGS|8|14|І повернув цар обличчя своє, та й поблагословив Ізраїлів збір, увесь же Ізраїлів збір стояв.
1KGS|8|15|І він сказав: Благословенний Господь, Бог Ізраїлів, що Своїми устами говорив був із моїм батьком Давидом, і рукою Своєю тепер виконав, говорячи:
1KGS|8|16|Від того дня, коли Я вивів Свій народ, Ізраїля, з Єгипту, Я не вибрав Собі міста зо всіх Ізраїлевих племен, щоб збудувати храм на пробування Мого Ймення там. І вибрав Я Давида, щоб був над Моїм Ізраїлевим народом.
1KGS|8|17|І було на серці мого батька Давида збудувати храм для Ймення Господа, Бога Ізраїля.
1KGS|8|18|Та сказав Господь до мого батька Давида: За те, що на твоєму серці було збудувати храм для Ймення Мого, ти зробив добре, що було тобі це на серці.
1KGS|8|19|Тільки ти не збудуєш цього храму, але син твій, що вийде із стегон твоїх, він збудує цей дім для Ймення Мого!
1KGS|8|20|І виконав Господь Своє слово, що Він говорив. І став я на місце батька мого Давида, та й сів на Ізраїлевому троні, як говорив був Господь, і я збудував оцей храм для Ймення Господа, Бога Ізраїлевого.
1KGS|8|21|І встановив я там місце для ковчега, де Господній заповіт, якого Він склав із нашими батьками, коли виводив їх з єгипетського краю.
1KGS|8|22|І став Соломон перед Господнім жертівником навпроти всього Ізраїлевого збору, і простяг руки свої до неба та й сказав:
1KGS|8|23|Господи, Боже Ізраїлів! Нема подібного Тобі Бога на небесах угорі та на землі долі. Ти стережеш заповіта та милість для Своїх рабів, що ходять перед Твоїм лицем усім своїм серцем.
1KGS|8|24|Ти додержав Своєму рабові, Давидові, батькові моєму, те, що говорив йому. І говорив Ти йому Своїми устами, а рукою Своєю виконав, як цього дня.
1KGS|8|25|А тепер, Господи, Боже Ізраїлів, додерж для Свого раба Давида, мого батька, те, що говорив був йому, кажучи: Не буде в тебе переводу з-перед лиця Мого нікому з тих, що сидітимуть на Ізраїлевім троні, якщо тільки сини твої будуть держатися своїх доріг, щоб ходити перед Моїм лицем, як ти ходив перед лицем Моїм.
1KGS|8|26|А тепер, Боже Ізраїлів, нехай буде запевнене слово Твоє, яке Ти говорив рабові Своєму Давидові, моєму батькові.
1KGS|8|27|Бо чи ж справді Бог сидить на землі? Ось небо та небо небес не обіймають Тебе, що ж тоді храм той, що я збудував?
1KGS|8|28|Та ти зглянешся на молитву Свого раба та на його благання, Господи, Боже мій, щоб почути спів та молитву, якою раб твій молиться перед лицем Твоїм сьогодні,
1KGS|8|29|щоб очі Твої були відкриті на цей храм уночі та вдень, на те місце, про яке Ти сказав: Нехай буде Ймення Моє там, щоб почути молитву, якою буде молитися Твій раб на цьому місці!
1KGS|8|30|І Ти будеш прислухатися до благання Свого раба, та Свого народу, Ізраїля, що будуть молитися на цьому місці. А Ти почуєш на місці Свого пробування, на небесах, і почуєш, і простиш.
1KGS|8|31|Як згрішить людина проти свого ближнього, і вимагатимуть від нього клятви, щоб він поклявся, і для клятви прийдуть перед Твій жертівник у цьому храмі,
1KGS|8|32|то Ти почуєш із небес, і зробиш, і розсудиш Своїх рабів, осудиш несправедливого, щоб дати його дорогу на його голову, і всправедливиш праведного, щоб віддати йому за його справедливістю.
1KGS|8|33|Коли Твій народ, Ізраїль, буде вдарений ворогом за те, що прогрішив Тобі, і коли вони звернуться до Тебе, і будуть славити Ім'я Твоє, і будуть молитися, і будуть благати Тебе в цьому храмі,
1KGS|8|34|то Ти почуєш із небес, і простиш гріх народу Свого, Ізраїля, і вернеш їх до землі, яку дав Ти їхнім батькам.
1KGS|8|35|Коли замкнеться небо й не буде дощу, бо прогрішаться Тобі, то коли знову вони помоляться на цьому місці, і будуть славити Ім'я Твоє, і від гріха свого відвернуться, бо Ти будеш їх впокоряти,
1KGS|8|36|то Ти почуєш на небесах, і простиш гріх Своїх рабів та народу Свого, Ізраїля, бо покажеш їм ту добру дорогу, якою вони підуть, і Ти даси дощ на Край Свій, якого Ти дав Своєму народові на спадщину.
1KGS|8|37|Голод коли буде в Краю, моровиця коли буде, посуха, жовтачка, сарана, черва коли буде, коли його ворог стане тіснити його в краю міст його, коли буде яка пораза, яка хвороба,
1KGS|8|38|усяка молитва, усяке благання, що буде від якої людини чи від усього народу Твого, Ізраїля, коли кожен почує рану свого серця, і простягне руки свої до цього храму,
1KGS|8|39|то Ти почуєш із небес, із місця постійного пробування Свого, і простиш, і зробиш, і даси кожному за всіма його дорогами, бо Ти Сам знаєш серце всіх людських синів,
1KGS|8|40|щоб вони боялися Тебе по всі дні, доки вони житимуть на поверхні землі, яку Ти дав батькам нашим.
1KGS|8|41|Також і чужинця, що він не з народу Твого, Ізраїля, і він прийде з далекого краю ради Ймення Твого,
1KGS|8|42|бо почують і вони про велике Ім'я Твоє, і про сильну руку Твою та про витягнене рамено Твоє, і прийде він і помолиться в цьому храмі,
1KGS|8|43|Ти почуєш це з небес, місця постійного пробування Свого, і зробиш усе, про що буде кликати до Тебе той чужинець, щоб усі народи землі пізнали Ім'я Твоє, щоб боялися Тебе, як народ Твій, Ізраїль, і щоб пізнали вони, що Ім'ям Твоїм названо цей храм, що я збудував.
1KGS|8|44|Коли народ Твій вийде на війну на свого ворога, дорогою, якою Ти пошлеш їх, і помоляться вони до Господа в напрямі до міста, що Ти вибрав його, та храму, що я збудував для Ймення Твого,
1KGS|8|45|то почуєш Ти з неба їхню молитву та їхнє благання, і вчиниш їм суд!
1KGS|8|46|Коли вони згрішать Тобі, бо немає людини, щоб вона не згрішила, і Ти розгніваєшся на них, і віддаси їх ворогові, а їхні полонителі відведуть їх у неволю до ворожого краю далекого чи близького,
1KGS|8|47|і коли вони прийдуть до розуму в краю, куди взяті в неволю, і навернуться, і будуть благати Тебе в краю полонителів своїх, говорячи: Ми згрішили, і безбожне чинили, були ми винні;
1KGS|8|48|і коли вони навернуться до Тебе всім своїм серцем і всією душею своєю в краю ворогів своїх, що їх поневолили, і помоляться до Тебе в напрямі до свого краю, що Ти дав їхнім батькам, у напрямі міста, яке Ти вибрав, та храму, що я збудував для Імени Твого,
1KGS|8|49|то Ти почуєш на небесах, постійному місті пробування Свого, їхню молитву та їхнє благання, і зробиш їм суд,
1KGS|8|50|і пробачиш Своєму народові, що вони згрішили Тобі, і всі їхні провини, що завинили проти Тебе, і нахилиш до любови полонителів їхніх, і вони змилосердяться над ними,
1KGS|8|51|бо вони народ Твій та наділ Твій, яке Ти вивів з Єгипту, з середини залізної гутничої печі,
1KGS|8|52|щоб очі Твої були відкриті на благання Твого раба та на благання народу Твого, Ізраїля, щоб прислухуватися до них, коли вони кликатимуть до Тебе.
1KGS|8|53|Бо Ти виділив їх зо всіх народів Собі на наділ, як говорив був через Мойсея, Свого раба, коли Ти виводив наших батьків із Єгипту, Владико мій, Господи!
1KGS|8|54|І сталося, як Соломон скінчив цю молитву й благання до Господа, то він устав від Господнього жертівника, де він стояв на колінах своїх, а руки його були простягнені до неба.
1KGS|8|55|І встав він, і поблагословив усі Ізраїлеві збори, говорячи сильним голосом:
1KGS|8|56|Благословенний Господь, що дав мир Своєму народові, Ізраїлеві, усе, як обіцяв був, не відпало ані одне слово зо всіх Його добрих слів, які Він говорив був через раба Свого Мойсея.
1KGS|8|57|Нехай буде Господь, Бог наш, з нами, як був Він із нашими батьками, нехай Він не опустить нас, нехай Він не покине нас,
1KGS|8|58|щоб прихиляти наше серце до Себе, щоб ми ходили всіма Його дорогами, щоб ми дотримувалися наказів Його, і уставів Його та постанов Його, як і Він наказав був нашим батькам.
1KGS|8|59|І нехай будуть оці слова мої, якими я благав перед Господнім лицем, близькі до Господа вдень та вночі, щоб чинити суд для раба Свого та суд для Свого народу, Ізраїля, день-у-день,
1KGS|8|60|щоб знали всі народи землі, що Господь Він Бог, і нема вже іншого!
1KGS|8|61|І нехай буде все серце ваше з Господом, Богом нашим, щоб ходити постановами його та щоб перестерігати заповіді Його, як цього дня!
1KGS|8|62|А цар та ввесь Ізраїль з ним принесли жертву перед Господнім лицем.
1KGS|8|63|І приніс Соломон жертву для мирних жертов, що приносив для Господа: двадцять і дві тисячі худоби великої, а худоби дрібної сто й двадцять тисяч. І виконали освячення Господнього храму цар та всі Ізраїлеві сини.
1KGS|8|64|Того дня цар освятив середину двору, що перед храмом Господнім, бо приготовив там цілопалення й хлібну жертву та лій мирних жертов, бо мідяний жертівник, що перед Господнім лицем, був малий для прийняття цілопалення й хлібної жертви та лою мирних жертов.
1KGS|8|65|І вчинив Соломон того часу свято, і з ним увесь Ізраїль, збір великий, що зійшовся звідти, де йдеться до Гамату аж до єгипетського потоку, перед лицем Господа, нашого Бога, сім день і сім день, чотирнадцять день.
1KGS|8|66|Восьмого дня він відпустив народ, а вони поблагословили царя та й пішли до наметів своїх, радісні та веселосерді через усе те добро, що Господь учинив Своєму рабові Давидові та Своєму народові Ізраїлеві.
1KGS|9|1|І сталося, як Соломон покінчив будувати храм Господній та дім царський, та все, що було бажанням Соломона, що прагнув він зробити,
1KGS|9|2|то Господь явився Соломонові другий раз, як явився йому в Ґів'оні.
1KGS|9|3|І сказав Господь до нього: Вислухав Я молитви твої та благання твої, якими благав ти перед лицем Моїм, Я освятив той храм, що ти збудував, щоб покласти Ім'я Моє там аж навіки. І будуть там Мої очі та серце Моє по всі дні.
1KGS|9|4|А ти, якщо будеш ходити перед лицем Моїм, як ходив був батько твій Давид, у чистості серця та в правоті, щоб зробити все, що наказав Я тобі, якщо будеш дотримуватися уставів Моїх та постанов Моїх,
1KGS|9|5|то трона царства твого над Ізраїлем Я поставлю навіки, як Я говорив був батькові твоєму Давидові, кажучи: Не буде переводу нікому з нащадків твоїх на Ізраїлевім троні.
1KGS|9|6|Якщо ж справді відвернетеся ви та ваші сини від Мене, і не будете дотримувати заповідей Моїх та уставів Моїх, що Я дав вам, і підете, і будете служити іншим богам, і буде те вклонятися їм,
1KGS|9|7|то Я винищу Ізраїля з поверхні землі, яку дав їм, а цей храм, що Я освятив для Ймення Свого, відкину від лиця Свого. І стане Ізраїль за приповістку та за посміховище серед усіх народів!
1KGS|9|8|І храм цей найвищий, кожен, хто проходитиме біля нього, скам'яніє та свисне від здивування. І скажуть: За що Господь зробив так цьому Краєві та храмові цьому?...
1KGS|9|9|І відкажуть: За те, що вони покинули Господа, Бога свого, Який вивів їхніх батьків з єгипетського краю, і держалися міцно інших богів, і вклонялися їм, і служили їм, тому Господь навів на них усе оце лихо!
1KGS|9|10|І сталося по двадцяти роках, коли Соломон збудував ті два доми, храм Господній та дім царський,
1KGS|9|11|а Хірам, цар тирський, достачав Соломонові кедрові дерева й дерева кипарисові, та золото на кожне бажання його, тоді цар Соломон дав Хірамові двадцять міст у краї Ґаліл.
1KGS|9|12|І вийшов Хірам із Тиру, щоб побачити ті міста, які дав йому Соломон, і не вподобались йому вони.
1KGS|9|13|І він сказав: Що це за міста, які ти дав мені, мій брате? І він назвав ім'я їм: Край Кавулу, і так вони звуться аж до цього дня.
1KGS|9|14|І послав Хірам цареві сто й двадцять талантів золота.
1KGS|9|15|А оце наказ тих поборів, які брав цар Соломон на збудування храму Господнього та дому свого, і Мілло, і муру єрусалимського, і Хацору, і Меґіддо, і Ґезеру.
1KGS|9|16|Фараон, єгипетський цар, прийшов і здобув Ґезер, та й спалив його огнем, а ханаанеянина, що сидів у місті, убив, і віддав його як віно для своєї дочки, Соломонової жінки.
1KGS|9|17|І вибудував Соломон Ґезера, і Бет-Горона Долішнього,
1KGS|9|18|і Баалата, і Тамара в пустині того краю,
1KGS|9|19|і всі міста на запаси, що були Соломонові, і міста на колесниці, і міста на верхівців, і інші бажання Соломонові, що бажав збудувати в Єрусалимі та на Ливані, та в усьому Краї панування його.
1KGS|9|20|Увесь народ, що позостався з амореян, хіттеян та періззеян, хіввеян та євусеян, що вони не з Ізраїлевих синів,
1KGS|9|21|їхні сини, що були позоставлені по них у Краю, яких Ізраїлеві сини не могли вигубити, то взяв їх Соломон за поборових працівників, і так є аж до цього дня.
1KGS|9|22|А з Ізраїлевих синів Соломон не дав раба, бо вони вояки, і його раби, і провідники його, і старші над трьома, і провідники над його колесницями та його верхівці.
1KGS|9|23|Оце приставлені провідники, що були над Соломоновою роботою, п'ятдесят і п'ять сотень, що правили народом, який робив на праці.
1KGS|9|24|Тільки фараонова дочка вийшла з Давидового Міста до свого дому, якого збудував їй; тоді збудував він Мілло.
1KGS|9|25|І приносив Соломон три рази річно цілопалення та мирні жертви на жертівнику, що збудував Господеві, і кадив на тому, що перед Господнім лицем. І викінчив він той дім.
1KGS|9|26|І цар Соломон наробив кораблів в Ецйон-Ґевері, що при Елоті на березі Червоного моря в едомському краї.
1KGS|9|27|І послав Хірам кораблями своїх рабів, моряків, що знають море, з рабами Соломоновими.
1KGS|9|28|І прийшли вони до Офіру, і взяли звідти чотири сотні й двадцять талантів золота, та й привезли до царя Соломона.
1KGS|10|1|А цариця Шеви, коли почула була про славу Соломона, щодо Господнього Імени, то прийшла випробувати його загадками.
1KGS|10|2|І прийшла вона до Єрусалиму з дуже великим багатством, з верблюдами, що несли пахощі, і з дуже численним золотом, і з дорогим камінням. І прийшла вона до Соломона, і говорила йому все, що було на серці її.
1KGS|10|3|І Соломон вияснив їй усі її слова, не було речі, незнаної цареві, якої не порішив би він їй.
1KGS|10|4|І побачила цариця Шеви всю Соломонову мудрість, та дім, що він збудував,
1KGS|10|5|і їжу столу його, і мешкання рабів його, і поставу слуг його та їхні одежі, і напої його, і цілопалення, що він приносить у Господньому домі, і не могла вона з дива вийти!
1KGS|10|6|І сказала вона до царя: Правдою було те, що я чула в своїм краї про твої діла та про твою мудрість.
1KGS|10|7|І не повірила я тим словам, аж поки не прийшла та не побачили мої очі, і ось не була представлена мені й половина: ти перевищив мудрість та добро тієї слави, про яку я чула!
1KGS|10|8|Щасливі люди твої, щасливі оці твої слуги, що завжди стоять перед обличчям твоїм, що слухають твою мудрість!
1KGS|10|9|Нехай буде благословенний Господь, Бог твій, що вподобав тебе, щоб посадити тебе на Ізраїлів трон, через Господню любов до Ізраїля навіки. І Він настановив тебе царем, щоб чинити право та справедливість.
1KGS|10|10|І дала вона цареві сто й двадцять талантів золота, і дуже багато пахощів та дорогого каміння. Більш уже ніколи не приходило так багато, як оці пахощі, що цариця Шеви дала цареві Соломонові!
1KGS|10|11|І також Хірамові кораблі, що довозили золото з Офіру, спроваджували з Офіру багато алмуґового дерева та дороге каміння.
1KGS|10|12|І поробив цар з алмуґового дерева поруччя для Господнього храму та для дому царського, і гусла, і арфи для співаків. Ніколи не приходило так багато алмуґового дерева, і не бачено аж до цього дня!
1KGS|10|13|А цар Соломон дав цариці Шеви на жадання її все, чого вона бажала, окрім того, що дав їй як царський дарунок Соломонів. І обернулася вона, та й пішла до свого краю, вона та слуги її.
1KGS|10|14|І була вага того золота, що приходило для Соломона в одному році, шість сотень шістдесят і шість талантів золота,
1KGS|10|15|окрім того, що приходило від купців та з торгівлі ходячих, та від усіх царів Арабії та краєвих намісників.
1KGS|10|16|І зробив цар Соломон дві сотні великих щитів із кутого золота, шість сотень шеклів золота йшло на одного щита,
1KGS|10|17|та три сотні щитів менших із кутого золота, три міні золота йшло на одного щита. І цар віддав їх до дому Ливанського Лісу.
1KGS|10|18|І зробив цар великого трона зо слонової кости, і покрив його щирим золотом.
1KGS|10|19|У трона було шість ступенів; а голова в трона кругляста позад його та поруччя з того й з того боку при місці сидіння, та два леви, що стояли при поруччях.
1KGS|10|20|І дванадцять левів стояли там на шости ступенях із того й з того боку. По всіх царствах не було так зробленого!
1KGS|10|21|І ввесь посуд на пиття царя Соломона золото, і всі речі дому Ливанського Лісу щире золото, нічого із срібла, воно за Соломонових днів не рахувалося за щось.
1KGS|10|22|Бо цар мав на морі таршіські кораблі разом із кораблями Хірамовими. Раз на три роки приходили таршіські кораблі, що довозили золото, і срібло, і слонову кість, і мавп, і пав.
1KGS|10|23|І став цар Соломон найбільшим від усіх земних царів, щодо багатства та щодо мудрости.
1KGS|10|24|І вся земля хотіла бачити Соломона, щоб послухати його мудрости, що Бог дав у його серце.
1KGS|10|25|І вони приносили кожен свого дара, речі срібні та речі золоті, й одежу, і зброю, і пахощі, коні та мули, із року в рік.
1KGS|10|26|І назбирав Соломон колесниць та верхівців, і було в нього тисяча й чотири сотні колесниць та дванадцять тисяч верхівців, і він порозміщував їх по колесничних містах та з царем в Єрусалимі.
1KGS|10|27|І Соломон наскладав в Єрусалимі срібла, як каміння, а кедрів наскладав, щодо численности, як сикомори, що в Шефелі!
1KGS|10|28|А коней, що були в Соломона, приводили з Єгипту та з Кеве; царські купці брали їх із Кеве за встановлені гроші.
1KGS|10|29|І входила й виходила колесниця з Єгипту за шість сотень шеклів срібла, а кінь за сто й п'ятдесят. І так вони вивозили все це своєю рукою для всіх царів хіттійських та царям сирійським.
1KGS|11|1|А цар Соломон покохав багато чужинних жінок: і дочку фараонову, моавітянок, аммонітянок, едомітянок, сидонянок, хіттіянок,
1KGS|11|2|із тих народів, що про них Господь сказав був Ізраїлевим синам: Не ввійде те між них, і вони не ввійдуть між вас, бо вони справді нахилять ваші серця до своїх богів. До них прихилився Соломон коханням.
1KGS|11|3|І було в нього жінок-княгинь сім сотень, а наложниць три сотні. І жінки його прихилили його серце.
1KGS|11|4|І сталося на час Соломонової старости, жінки його прихилили його серце до інших богів; і серце його не було все з Господом, Богом, як серце його батька Давида.
1KGS|11|5|І пішов Соломон за Астартою, богинею сидонською, та за Мілкомом, гидотою аммонітською.
1KGS|11|6|І робив Соломон зле в очах Господніх, і не йшов певно за Господом, як його батько Давид.
1KGS|11|7|Тоді Соломон збудував жертівника для Кемоша, моавської гидоти, на горі, що навпроти Єрусалиму, та для Молоха, гидоти аммонських синів.
1KGS|11|8|І так він зробив для всіх своїх чужинних жінок, що кадили та приносили жертви для своїх богів.
1KGS|11|9|І розгнівався Господь на Соломона, бо його серце відхилилося від Господа, Бога Ізраїлевого, що два рази йому являвся,
1KGS|11|10|і наказував йому про цю річ, щоб не ходити за іншими богами. Та не виконував він того, що наказав був Господь.
1KGS|11|11|І сказав Господь до Соломона: Тому, що було це з тобою, і не виконував ти Мого заповіту та постанов Моїх, що Я наказав був тобі, Я конче відберу царство твоє, та й дам його твоєму рабові.
1KGS|11|12|Тільки за твоїх днів не зроблю того ради батька твого Давида, з руки сина твого відберу його!
1KGS|11|13|Та всього царства Я не відберу, одне племено Я дам синові твоєму ради раба Мого Давида та ради Єрусалиму, якого Я вибрав.
1KGS|11|14|І поставив Господь Соломонові за противника едомлянина Гадада, він із царського насіння в Едомі.
1KGS|11|15|І сталося, коли Давид був з Едомом, коли Йоав, начальник війська, пішов поховати трупи, то він повбивав кожного чоловічої статі в Едомі.
1KGS|11|16|Бо шість місяців сидів там Йоав та ввесь Ізраїль, аж поки він не вигубив кожного чоловічої статі в Едомі.
1KGS|11|17|І втік Гадад, він та з ним мужі едомські, зо слуг його батька, щоб піти до Єгипту; а Гадад був тоді малим хлопцем.
1KGS|11|18|І встали вони з Мідіяну й пішли до Парану; і набрали вони з собою людей з Парану, та й прийшли до Єгипту, до фараона, царя єгипетського, а той дав йому дім та призначив йому утримання, і дав йому землю.
1KGS|11|19|І знайшов Гадад велику милість у фараонових очах, і він дав йому за жінку сестру своєї жінки, сестру цариці Тахпенеси.
1KGS|11|20|І породила йому сестра Тахпенеси сина його Ґенувата, а Тахпенеса виховала його в фараоновому домі. І був Ґенуват у фараоновому домі серед фараонових синів.
1KGS|11|21|І почув Гадад в Єгипті, що Давид спочив із своїми батьками, та що помер Йоав, начальник війська. І сказав Гадад до фараона: Відпусти мене, й я піду до свого Краю!
1KGS|11|22|А фараон йому відказав: Чого тобі бракує при мені, що ти оце хочеш іти до свого краю? Та той сказав: Ні, таки конче відпусти мене!
1KGS|11|23|І поставив Бог йому, Соломонові, за противника ще й Резона, сина Ел'яди, що втік від Гадад'езера, царя Цови, свого пана.
1KGS|11|24|І зібрав він при собі людей, та й став провідником банди, коли Давид розбивав їх. І пішли вони до Дамаску, й осілися в ньому, і панували в Дамаску.
1KGS|11|25|І був він противником для Ізраїля за всіх Соломонових днів, а це окрім того лиха, що чинив Гадад. І бридив він Ізраїлем, і запанував над Сирією.
1KGS|11|26|А Єровоам, син Неватів, єфремівець, із Цереди, а ім'я його матері Церуа, жінка вдова, був раб Соломонів. І підняв він руку на царя.
1KGS|11|27|А оце та причина, що він підняв руку на царя: Соломон будував Мілло, і поправив пролім у Місті Давида, свого батька.
1KGS|11|28|А той муж Єровоам був відважний. І побачив Соломон цього юнака, що він роботящий, і призначив його над усіма носіями Йосипового дому.
1KGS|11|29|І сталося того часу, і вийшов Єровоам з Єрусалиму. І знайшов його на дорозі шілонянин Ахійя, пророк. Він був одягнений в нову одіж, й обидва вони були самі на полі.
1KGS|11|30|І схопив Ахійя за ту нову одежу, що була на ньому, та й подер її на дванадцять кусків.
1KGS|11|31|І сказав він до Єровоама: Візьми собі десять кусків, бо так сказав Господь, Бог Ізраїля: Оце Я віддираю царство з Соломонової руки, і дам тобі десять племен.
1KGS|11|32|А одне племено буде йому ради Мого раба Давида та ради Єрусалиму, міста, що Я вибрав його зо всіх Ізраїлевих племен.
1KGS|11|33|Це тому, що вони покинули Мене і вклонялися Астарті, сидонській богині, і Кемошеві, богові моавському, та Мілкомові, богові аммонітському, і не пішли Моїми дорогами, щоб виконувати добре в Моїх очах, і постанови Мої та заповіді Мої, як батько його Давид.
1KGS|11|34|Та не візьму Я всього царства з руки його, бо оставлю його володарем по всі дні життя його ради раба Мого Давида, що Я вибрав його, який додержував заповідів Моїх та постанов Моїх.
1KGS|11|35|І візьму Я царство з руки його сина, та й дам його тобі, оті десять племен.
1KGS|11|36|А синові його дам одне племено, щоб позоставався світильник рабові Моєму Давидові, по всі дні перед лицем Моїм в Єрусалимі, місці, що Я вибрав Собі, щоб там перебувало Моє Ймення.
1KGS|11|37|А тебе Я візьму, і ти будеш царювати над усім, чого пожадає душа твоя, і ти будеш царем над Ізраїлем.
1KGS|11|38|І станеться, коли ти слухатимешся всього, що Я накажу тобі, і підеш Моїми дорогами, і робитимеш добре в очах Моїх, щоб виконувати постанови Мої та заповіді Мої, як робив раб Мій Давид, то Я буду з тобою, і побудую тобі міцний дім, як Я збудував був Давидові, і дам тобі Ізраїля.
1KGS|11|39|І буду впокоряти Давидове насіння ради того, тільки не по всі дні.
1KGS|11|40|І шукав Соломон, щоб забити Єровоама. І встав Єровоам, і втік до Єгипту, до Шішака, єгипетського царя. І пробував він в Єгипті аж до Соломонової смерти.
1KGS|11|41|А решта Соломонових діл, і все, що він зробив був, та мудрість його, ото вони написані в книзі Соломонові діла.
1KGS|11|42|А днів, коли Соломон царював в Єрусалимі над усім Ізраїлем, було сорок літ.
1KGS|11|43|І спочив Соломон зо своїми батьками, і був похований у Місті Давида, батька свого, а замість нього зацарював син його Рехав'ам.
1KGS|12|1|І пішов Рехав'ам до Сихему, бо до Сихему зійшовся ввесь Ізраїль, щоб настановити його царем.
1KGS|12|2|І сталося, що це почув Єровоам, Неватів син, коли був іще в Єгипті, куди втік від царя Соломона. І осівся Єровоам ув Єгипті.
1KGS|12|3|І послали й покликали його. І прийшов Єровоам та всі Ізраїлеві збори, і вони говорили до Рехав'ама, кажучи:
1KGS|12|4|Твій батько вчинив був тяжким наше ярмо, а ти тепер полегши жорстоку роботу батька свого та тяжке його ярмо, що наклав він був на нас, і ми будемо служити тобі.
1KGS|12|5|А він відказав їм: Ідіть ще на три дні, і верніться до мене. І пішов той народ.
1KGS|12|6|І радився цар Рехав'ам зо старшими, що стояли перед обличчям його батька Соломона, коли був він живий, говорячи: Як ви радите відповісти цьому народові?
1KGS|12|7|І вони говорили йому, кажучи: Якщо ти сьогодні будеш рабом цьому народові, і будеш служити їм, і відповіси їм, і говоритимеш їм добрі слова, то вони будуть тобі рабами по всі дні.
1KGS|12|8|Та він відкинув пораду старших, що радили йому, і радився з молодиками, що виросли разом із ним, що стояли перед ним.
1KGS|12|9|І сказав він до них: Що ви радите, і що відповімо цьому народові, який говорив мені, кажучи: Полегши ярмо, що твій батько наклав був на нас.
1KGS|12|10|І говорили до нього ті молодики, що виросли з ним, кажучи: Так скажеш тому народові, що промовляв до тебе, говорячи: Твій батько вчинив був тяжким наше ярмо, а ти дай полегшу нам. Отак скажеш до них: Мій мізинець грубший за стегна мого батька!
1KGS|12|11|А тепер: мій батько наклав був на вас тяжке ярмо, а я додам до вашого ярма! Батько мій карав вас бичами, а я каратиму вас скорпіонами!
1KGS|12|12|І прийшов Єровоам та ввесь народ до Рехав'ама третього дня, як цар говорив, кажучи: Верніться до мене третього дня.
1KGS|12|13|І цар жорстоко відповів народові, і відкинув пораду старших, що радили йому.
1KGS|12|14|І він говорив до них за порадою тих молодиків, кажучи: Мій батько вчинив був тяжким ваше ярмо, а я додам до вашого ярма. Батько мій карав вас бичами, а я каратиму вас скорпіонами!...
1KGS|12|15|І не послухався цар народу, бо причина була від Господа, щоб справдилося слово Його, яке говорив був Господь через шілонянина Ахійю до Єровоама, Неватового сина.
1KGS|12|16|І побачив увесь Ізраїль, що цар не послухався їх, і народ відповів цареві, кажучи: Яка нам частина в Давиді? І спадщини нема нам у сині Єссея! До наметів своїх, о Ізраїлю! Познай тепер дім свій, Давиде!... І пішов Ізраїль до наметів своїх.
1KGS|12|17|А Ізраїлеві сини, що сиділи в Юдиних містах, тільки над ними зацарював Рехав'ам.
1KGS|12|18|І послав цар Рехав'ам Адонірама, що був над даниною, та ввесь Ізраїль закидав його камінням, і він помер. А цар Рехав'ам поспішив сісти на колесницю та втекти до Єрусалиму.
1KGS|12|19|І збунтувався Ізраїль проти Давидового дому, і від нього відпав, і так є аж до цього дня.
1KGS|12|20|І сталося, як увесь Ізраїль почув, що вернувся Єровоам, то послали й покликали його на збори, та й настановили його царем над усім Ізраїлем. За домом Давида не було нікого, окрім одного Юдиного племени.
1KGS|12|21|І прийшов Рехав'ам до Єрусалиму, і зібрав увесь Юдин дім та Веніяминове племено, сто й вісімдесят тисяч вибраних військових, щоб воювати з Ізраїлевим домом, щоб вернути царство Рехав'амові, Соломоновому синові.
1KGS|12|22|І було Боже слово до Шемаї, чоловіка Божого, говорячи:
1KGS|12|23|Скажи Рехав'амові, Соломоновому синові, цареві Юдиному, та всьому домові Юдиному й Веніяминовому, і решті народу, говорячи:
1KGS|12|24|Так говорить Господь: Не йдіть і не воюйте з своїми братами, Ізраїлевими синами! Верніться кожен до дому свого, бо ця річ сталася від Мене! І вони послухалися Господнього слова, і вернулися, щоб піти за Господнім словом.
1KGS|12|25|І збудував Єровоам Сихема в Єфремових горах, та й осівся в ньому. І вийшов він звідти, і збудував Пенуїла.
1KGS|12|26|І сказав Єровоам у своєму серці: Тепер вернеться царство до Давидового дому!
1KGS|12|27|Якщо народ цей буде ходити до Єрусалиму, щоб приносити жертви в Господньому домі, то вернеться серце цього народу до їхнього пана, до Рехав'ама, царя Юдиного. І вони заб'ють мене, та й вернуться до Рехав'ама, царя Юдиного.
1KGS|12|28|І порадився цар, і зробив два золоті тельці, і сказав до народу: Досить вам ходити до Єрусалиму! Оце, Ізраїлю, боги твої, що вивели тебе з єгипетського краю.
1KGS|12|29|І поставив він одного в Бет-Елі, а одного в Дані.
1KGS|12|30|І була та річ на гріх, бо народ ходив до одного з них аж до Дану.
1KGS|12|31|І зробив він жертівне місце на пагірку, і настановив священиків з усього народу, що не були з Левієвих синів.
1KGS|12|32|І встановив Єровоам свято в восьмому місяці, п'ятнадцятого для місяця, подібне до свята, що в Юді, і приносив жертву на жертівнику. Так зробив він у Бет-Елі, щоб приносити в жертву тельцям, які він зробив. І настановив він у Бет-Елі священиків пагірків, що поробив.
1KGS|12|33|І приносив він жертви на жертівнику, що зробив у Бет-Елі, п'ятнадцятого дня восьмого місяця, якого вимислив з свого серця. І вчинив він свято для Ізраїлевих синів, і підійшов до жертівника, щоб покадити...
1KGS|13|1|А ось чоловік Божий прийшов за Господнім словом із Юди до Бет-Елу. А Єровоам стояв при жертівнику, щоб кадити.
1KGS|13|2|І кликнув чоловік Божий при жертівнику за словом Господнім і сказав: Жертівнику, жертівнику, так сказав Господь: Ось у Давидовому домі народиться син, Йосія ім'я йому, і він на тобі принесе в жертву священиків пагірків, що на тобі кадять, і кості людські спаляться на тобі.
1KGS|13|3|І дасть він того дня чудо, говорячи: Оце те чудо, про яке говорив Господь: Ось цей жертівник розпадеться, і висиплеться попіл, що на ньому!...
1KGS|13|4|І сталося, як цар почув слова цього Божого чоловіка, що кликав до жертівника в Бет-Елі, то Єровоам простяг руку свою від жертівника, говорячи: Схопіть його! І всохла рука йому, яку він простяг до нього, і він не міг вернути її до себе...
1KGS|13|5|А жертівник розпався, і попіл висипався з жертівника, за тим чудом, що дав Божий чоловік за словом Господнім...
1KGS|13|6|А цар відповів і сказав до Божого чоловіка: Умилостив лице Господа, Бога твого, і помолися за мене, і нехай вернеться рука моя до мене! І чоловік Божий умилостивив Господнє лице, і царська рука вернулася до нього, і була, як перед тим...
1KGS|13|7|І сказав цар до Божого чоловіка: Увійди зо мною до дому й попоїж, і я дам тобі дара!
1KGS|13|8|А чоловік Божий сказав до царя: Якщо ти даси мені пів дому свого, не ввійду я з тобою, і не їстиму хліба, і не питиму води в цьому місці!...
1KGS|13|9|Бо так наказано мені за словом Господнім, говорячи: Ти не їстимеш хліба, і не питимеш води, і не вернешся дорогою, якою пішов!
1KGS|13|10|І пішов він іншою дорогою, і не вернувся тією дорогою, що нею прийшов був до Бет-Елу.
1KGS|13|11|А один старий пророк сидів у Бет-Елі. І прийшли його сини, і розповіли йому про ввесь чин, що зробив Божий чоловік сьогодні в Бет-Елі, про ті слова, що він говорив до царя, і оповіли їх своєму батькові.
1KGS|13|12|І промовив до них їхній батько: Де ж та дорога, якою він пішов? А його сини бачили ту дорогу, якою пішов Божий чоловік, що прийшов був з Юди.
1KGS|13|13|І сказав він до синів своїх: Осідлайте мені осла! І вони осідлали йому осла, і він сів на нього.
1KGS|13|14|І поїхав він за Божим чоловіком, і знайшов його, як сидів під дубом. І сказав він до нього: Чи ти той Божий чоловік, що прийшов із Юди? А той відказав: Я.
1KGS|13|15|І сказав він до нього: Іди зо мною до дому та з'їж хліба!
1KGS|13|16|А той відказав: Не можу вернутися з тобою та ввійти з тобою, і не їстиму хліба, і не питиму води з тобою в цьому місці!
1KGS|13|17|Бо було мені сказано за словом Господнім: Не їстимеш хліба й не питимеш там води, і не вернешся тією дорогою, якою ти йшов!
1KGS|13|18|А той відказав йому: І я пророк, як ти! А Ангол говорив мені за Господнім словом, кажучи: Заверни його з собою до дому свого, і нехай він їсть хліб і нехай п'є воду. Він же говорив йому неправду!
1KGS|13|19|І він вернувся з ним, і їв хліб у його домі та пив воду...
1KGS|13|20|І сталося, як сиділи вони при столі, то було Господнє слово до пророка, що вернув його.
1KGS|13|21|І він кликнув до Божого чоловіка, що прийшов із Юди, говорячи: Так сказав Господь: Тому, що був ти неслухняний Господнім наказам, і не додержував тієї заповіді, що наказав тобі Господь, Бог твій,
1KGS|13|22|і ти вернувся, і їв хліб та пив воду в місці, про яке Він говорив тобі: Не їж хліба й не пий води, то не ввійде твій труп до гробу батьків твоїх!...
1KGS|13|23|І сталося, як той поїв хліба та напився, то він осідлав йому осла, тому пророкові, що він вернув його.
1KGS|13|24|І той подався, та спіткав його на дорозі лев, та й забив його. І був кинений труп його на дорозі, а осел стояв при ньому, а той лев стояв при трупі...
1KGS|13|25|Аж ось приходять люди, і побачили того трупа, киненого на дорозі, та лева, що стояв при трупі. І вони прийшли й говорили в тім місті, де сидів старий пророк.
1KGS|13|26|І почув про це той пророк, що вернув його з дороги, та й сказав: Це той Божий чоловік, що був неслухняний Господнім наказам, і Господь дав його левові, і він роздер його та вбив його за Господнім словом, що говорив йому.
1KGS|13|27|І сказав він до синів своїх, говорячи: Осідлайте мені осла! І осідлали.
1KGS|13|28|І поїхав він, і знайшов його трупа, киненого на дорозі, й осла та лева, що стояли при трупі, не з'їв той лев труп а й не роздер осла.
1KGS|13|29|І підняв той пророк трупа Божого чоловіка, і поклав його на осла, та й вернув його. І ввійшов старий пророк до міста, щоб оплакати та поховати того.
1KGS|13|30|І поклав він його в своїм гробі, і плакали над ним: Ой, брате мій!
1KGS|13|31|І сталося по його похороні, і сказав він до синів своїх, говорячи: Коли я помру, то поховаєте мене в гробі, що в ньому похований цей Божий чоловік. При костях його покладіть мої кості!
1KGS|13|32|Бо конче збудеться те слово, що він кликнув був за Господнім словом над тим жертівником, що в Бет-Елі, та над усіма жертівниковими місцями на пагірках, що в містах самарійських.
1KGS|13|33|По цій пригоді Єровоам не зійшов зо своєї злої дороги, і настановляв священиків пагірків з усього народу, хто хотів, той призначався, і ставав священиком пагірків.
1KGS|13|34|І стала та річ гріхом для Єровоамового дому, і на вигублення, і на винищення з-над поверхні землі.
1KGS|14|1|Того часу заслаб Авійя, Єровоамів син
1KGS|14|2|І сказав Єровоам до своєї жінки: Устань та переберися, і не пізнають, що ти Єровоамова жінка. І підеш до Шіло, ото там пророк Ахійя, який говорив про мене, що я буду царем над цим народом.
1KGS|14|3|І візьми в свою руку десять хлібів і калачі та дзбанок меду, і ввійдеш до нього. Він скаже тобі, що буде хлопцеві.
1KGS|14|4|І зробила так Єровоамова жінка. І встала вона, та й пішла до Шіло, і ввійшла до Ахійєвого дому. А Ахійя не міг бачити, бо очі йому стемніли через його старість.
1KGS|14|5|І Господь сказав до Ахійї: Ось приходить Єровоамова жінка, щоб запитати від тебе слово про сина свого, бо він слабий. Отак і так будеш їй говорити. І станеться, коли вона ввійде, то вдаватиме чужу.
1KGS|14|6|І сталося, як Ахійя почув шарудіння ніг її, як вона входила до входу, то сказав: Увійди, Єровоамова жінко! Чому то ти вдаєш чужу? А я посланий до тебе з твердою звісткою.
1KGS|14|7|Іди, скажи Єровоамові: Так сказав Господь, Бог Ізраїлів: Тому, що Я підніс тебе з-посеред народу, і дав тебе за князя над Моїм народом, Ізраїлем,
1KGS|14|8|і відірвав царство від Давидового дому й дав його тобі, та ти не був, як Мій раб Давид, що додержував заповідей Моїх, і що ходив за Мною всім серцем своїм, щоб робити тільки добре в очах Моїх,
1KGS|14|9|і робив ти гірше за всіх, хто був перед тобою, і ти пішов і наробив собі інших богів та литих бовванів, щоб гнівити Мене, а Мене ти відкинув геть,
1KGS|14|10|тому ось Я наводжу 935 8688 лихо 7451 на Єровоамів 3379 дім 1004, і вигублю 3772 8689 в Єровоама 3379 навіть те, що мочить 8366 8688 на стіну 7023, невільника 6113 8803 й вільного 5800 8803 в Ізраїлі 3478, і вимету 1197 8765 позостале 310 по Єровоамовім 3379 домі 1004, як вимітається 1197 8762 сміття 1557, аж не 8552 8800 0 зостанеться 8552 8800 0 нічого.
1KGS|14|11|Померлого в Єровоама в місті поїдять пси, а померлого на полі поїсть птаство небесне. Так сказав Господь.
1KGS|14|12|А ти встань, іди до свого дому. Як ноги твої входитимуть до міста, то помре той хлопець.
1KGS|14|13|І буде його оплакувати ввесь Ізраїль, і поховають його, бо він один в Єровоама ввійде до гробу, бо тільки в ньому в Єровоамовім домі була знайдена добра річ для Господа, Бога Ізраїлевого.
1KGS|14|14|А Господь поставить Собі царя над Ізраїлем, який вигубить Єровоамів дім того дня. Та що станеться тепер?
1KGS|14|15|І поб'є Господь Ізраїля, і він захитається, як хитається очерет на воді! І вирве Він Ізраїля з-над цієї хорошої землі, яку дав їхнім батькам, і порозкидає їх по той бік Річки за те, що вони поробили собі Астарти, що гнівають Господа.
1KGS|14|16|І Він видасть Ізраїля через гріх Єровоама, що грішив сам, і що ввів у гріх Ізраїля.
1KGS|14|17|І встала Єровоамова жінка, і пішла, і прийшла до Тірци. Як вона входила до порога дому, то той хлопець помер...
1KGS|14|18|І поховали його, й оплакував його ввесь Ізраїль за словом Господа, що говорив через раба Свого пророка Ахійю.
1KGS|14|19|А решта Єровоамових діл, як він воював та як він царював, ось вони написані в Книзі Хроніки Ізраїлевих царів.
1KGS|14|20|А час, який царював Єровоам, двадцять і два роки. І спочив він із батьками своїми, а замість нього зацарював син його Надав.
1KGS|14|21|А Рехав'ам, син Соломонів, царював у Юді. Рехав'ам був віку сорока й одного року, коли зацарював, а царював він сімнадцять літ в Єрусалимі, у тому місті, яке вибрав Господь зо всіх Ізраїлевих племен, щоб покласти там Своє Ймення. А ім'я його матері: аммонітка Наама.
1KGS|14|22|А Юда робив зло в Господніх очах, і вони гнівили Його більш від усього того, що чинили їхні батьки своїм гріхом, яким грішили.
1KGS|14|23|І також вони будували собі жертівники на пагірках, і стовпи, і Астарти на кожному високому взгір'ї та під кожним зеленим деревом.
1KGS|14|24|І також були блудодії в тому краї, вони чинили всю гидоту тих людей, що Господь прогнав їх від Ізраїлевого обличчя.
1KGS|14|25|І сталося п'ятого року царя Рехав'ама, пішов Шушак, єгипетський цар, на Єрусалим.
1KGS|14|26|І позабирав він скарби Господнього дому та скарби дому царевого, і все забрав. І забрав він усі золоті щити, що Соломон поробив був.
1KGS|14|27|А цар Рехав'ам поробив замість них мідяні щити, і віддав їх на руки провідників бігунів, що стерегли вхід до царського дому.
1KGS|14|28|І бувало, як тільки цар ішов до Господнього дому, бігуни носили їх, а потім вертали їх до комори бігунів.
1KGS|14|29|А решта Рехав'амових діл та все, що він зробив, ось вони написані в Книзі Хроніки Юдиних царів.
1KGS|14|30|А війна між Рехав'амом та між Єровоамом точилася по всі дні.
1KGS|14|31|І спочив Рехав'ам зо своїми батьками, і був він похований зо своїми батьками в Давидовому Місті. А ім'я його матері аммонітянка Наама. А замість нього зацарював його син Авійям.
1KGS|15|1|А вісімнадцятого року царя Єровоама, Неватового сина, над Юдою зацарював Авійям.
1KGS|15|2|Три роки царював він в Єрусалимі. А ім'я його матері Мааха, Авесаломова дочка.
1KGS|15|3|І він ходив в усіх гріхах свого батька, які той робив перед ним, і серце його не було все з Господом, Богом своїм, як серце його батька Давида.
1KGS|15|4|Бо Господь, Бог його, ради Давида дав йому світильника в Єрусалимі, щоб поставити сина його по ньому та укріпити Єрусалим.
1KGS|15|5|Бо Давид робив добре в Господніх очах, і не відступав від усього що Він наказав був йому, по всі дні життя свого, окрім справи хіттянина Урії.
1KGS|15|6|А війна між Рехав'амом та між Єровоамом точилася по всі дні життя його.
1KGS|15|7|А решта Авійямових діл та все, що він зробив, ось вони написані в Книзі Хроніки Юдиних царів. І війна точилася між Авійямом та між Єровоамом.
1KGS|15|8|І спочив Авійям зо своїми батьками, і поховали його в Давидовому Місті, а замість нього зацарював син його Аса.
1KGS|15|9|А року двадцятого Єровоама, Ізраїлевого царя, зацарював Аса, цар Юдин.
1KGS|15|10|І він царював в Єрусалимі сорок і один рік. А ім'я його матері Мааха, Авесаломова дочка.
1KGS|15|11|І робив Аса добре в Господніх очах, як батько його Давид.
1KGS|15|12|І вигнав він блудодіїв із краю, і повикидав усіх божків, яких поробили були їхні батьки.
1KGS|15|13|І навіть матір свою Мааху, і її він позбавив права бути царицею, бо вона зробила була ідола для Астарти. І Аса порубав ідола її, та й спалив у долині Кедрон.
1KGS|15|14|А пагірки не минулися; тільки Асине серце було все з Господом по всі його дні.
1KGS|15|15|І вніс він до Господнього дому присвячені речі свого батька та присвячені речі свої, срібло, і золото, і посуд.
1KGS|15|16|А війна точилася між Асою та між Башою по всі їхні дні.
1KGS|15|17|І пішов Баша, цар Ізраїлів, на Юду, і будував Раму, щоб не дати нікому від Аси, царя Юдиного, виходити та входити.
1KGS|15|18|І взяв Аса все срібло та золото, позостале в скарбницях храму Господнього та дому царевого, та й дав його до руки своїх слуг. І послав їх цар Аса до Бен-Гадада, сина Тавримонна, сина Хезйонового, сирійського царя, що сидів у Дамаску, говорячи:
1KGS|15|19|Є умова між мною та між тобою, між батьком моїм та між батьком твоїм. Ось послав я тобі дара, срібла та золота, іди, зламай умову свою з Башею, царем Ізраїлевим, і нехай він відійде від мене.
1KGS|15|20|І послухався Бен-Гаддад царя Аси, і послав провідників свойого війська на Ізраїлеві міста, та й побив Іййона, і Дана, і Авела, Бат-Мааху, і всього Кінерота та всю землю Нефталимову.
1KGS|15|21|І сталося, як Баша це почув, то перестав будувати Раму, й осівся в Тірці.
1KGS|15|22|А цар Аса закликав до послуху всього Юду, нікого не виключаючи, і вони повиносили каміння Рами та її дерево, що з них будував був Баша. І цар Аса збудував з того Веніяминову Ґеву.
1KGS|15|23|А решта діл Аси та вся лицарськість його, і все, що він зробив був, і міста, які побудував, ось вони написані в Книзі Хроніки Юдиних царів; тільки на час старости своєї він заслаб був на свої ноги.
1KGS|15|24|І спочив Аса з батьками своїми, і був похований з батьками своїми в Місті Давида, свого батька. А замість нього зацарював його син Йосафат.
1KGS|15|25|А над Ізраїлем зацарював Надав, Єровоамів син, у другому році Аси, царя Юдиного, та й царював над Ізраїлем два роки.
1KGS|15|26|І робив він зле в Господніх очах, і ходив дорогою батька свого та в гріху його, що вводив теж у гріх Ізраїля.
1KGS|15|27|І змовився на нього Баша, син Ахійї, з Іссахарового дому, та й побив його Баша в Ґіббетоні филистимському. А Надав та ввесь Ізраїль облягали Ґіббетон.
1KGS|15|28|І вбив його Баша в третьому році Аси, царя Юдиного, та й зацарював замість нього.
1KGS|15|29|І сталося, як зацарював він, то побив увесь Єровоамів дім, не позоставив Єровоамові жодної душі, аж поки не вигубив його, за словом Господа, що говорив через Свого раба шілонянина Ахійю,
1KGS|15|30|за гріх Єровоама, що грішив сам і що вводив у гріх Ізраїля, через свій гнів, яким гнівив Господа, Бога Ізраїлевого.
1KGS|15|31|А решта діл Надава та все, що він був зробив, ось вони написані в Книзі Хроніки Ізраїлевих царів.
1KGS|15|32|А війна точилася між Асою та між Башею, Ізраїлевим царем, по всі дні їх.
1KGS|15|33|Третього року Аси, царя Юдиного, зацарював Баша, син Ахійїн, над усім Ізраїлем у Тірці, на двадцять і чотири роки.
1KGS|15|34|І робив він зло в Господніх очах, і ходив дорогою Єровоама та в гріху його, що вводив у гріх Ізраїля.
1KGS|16|1|І було Господнє слово до Єгу, Хананієвого сина, про Башу, говорячи:
1KGS|16|2|Тому, що Я підніс тебе з пороху, і настановив тебе володарем над Моїм народом, Ізраїлем, а ти пішов Єровоамовою дорогою та вводив у гріх народ Мій, Ізраїля, щоб гнівити Мене гріхами їх,
1KGS|16|3|то ось Я вигублю по Баші та по домі його, зроблю твій дім, як дім Єровоама, Неватового сина.
1KGS|16|4|Померлого в Баші в місті з'їдять пси, а померлого йому на полі, поїсть птаство небесне.
1KGS|16|5|А решта діл Баші, і що він зробив був, і лицарськість його, ось вони написані в Книзі Хроніки Ізраїлевих царів.
1KGS|16|6|І спочив Баша зо своїми батьками, і був похований в Тірці, а замість нього зацарював син його Ела.
1KGS|16|7|І було слово Господнє через пророка Єгу, сина Хананієвого, до Баші та до дому його, а то через усе те зло, що коїв він у Господніх очах, щоб гнівити Його чином своїх рук, щоб бути, як Єровоамів дім, що Він побив його.
1KGS|16|8|Двадцять і шостого року Аси, царя Юдиного, зацарював Ела, Башин син, над Ізраїлем у Тірці, на два роки.
1KGS|16|9|І змовився на нього його раб Зімрі, провідник половини колесниць. І коли він, п'яний, пив у домі Арци, що був над його домом у Тірці,
1KGS|16|10|то прийшов Зімрі й убив його, і вбив його в двадцятому й сьомому році Аси, царя Юдиного, та й зацарював замість нього.
1KGS|16|11|І сталося, як він зацарював та сів на його троні, то він вибив увесь Башин дім, не позоставив навіть того, що мочить на стіну, ані рідних його, ані друзів його.
1KGS|16|12|І вигубив Зімрі ввесь Башин дім, за словом Господа, що промовляв був до Баші через пророка Єгу,
1KGS|16|13|за всі гріхи Баші та гріхи Елі, його сина, що грішили самі, і що вводили в гріх Ізраїля, щоб гнівити Господа, Бога Ізраїлевого, своїми гидотами.
1KGS|16|14|А решта діл Елі та все, що він робив, ось вони написані в Книзі Хроніки Ізраїлевих царів.
1KGS|16|15|У році двадцятому й сьомому Аси, царя Юдиного, зацарював Зімрі в Тірці на сім день, коли народ облягав филистимський Ґіббетон.
1KGS|16|16|І прочув народ, що облягав, таке: Змовився Зімрі та й убив царя! І ввесь Ізраїль настановив царем над Ізраїлем Омрі, провідника війська, того дня в таборі.
1KGS|16|17|І піднялися Омрі та ввесь Ізраїль із ним із Ґіббетону, і облягли Тірцу.
1KGS|16|18|І сталося, як побачив Зімрі, що місто здобуте, то ввійшов до палацу царевого дому, та й спалив над собою царський дім огнем, і помер
1KGS|16|19|за гріх свій, що грішив ним, щоб робити зло в Господніх очах, щоб ходити дорогою Єровоама та в гріху його, який він чинив, щоб вводити в гріх Ізраїля.
1KGS|16|20|А решта діл Зімрі та змова його, що вчинив був, ось вони написані в Книзі Хроніки Ізраїлевих царів.
1KGS|16|21|Тоді Ізраїлів народ поділився пополовині: половина народу була за Тівні, Ґінатового сина, щоб настановити його царем, а половина за Омрі.
1KGS|16|22|Та був сильніший народ, що стояв за Омрі, від народу, що був за Тівні, Ґінатового сина. І помер Тівні, а зацарював Омрі.
1KGS|16|23|У році тридцятому й першому Аси, царя Юдиного, над Ізраїлем зацарював на дванадцять літ Омрі. У Тірці царював він шість років.
1KGS|16|24|І купив він від Шемера гору Шомерон за два таланти срібла, і забудував гору, і назвав ім'я міста, яке збудував, іменем пана тієї гори: Шомерон.
1KGS|16|25|І робив Омрі зло в Господніх очах, і чинив зло більше від усіх, хто був перед ним.
1KGS|16|26|І ходив він усією дорогою Єровоама, сина Неватового, та в гріхах його, якими вводив у гріх Ізраїля, щоб гнівити Господа, Бога Ізраїля, гидотами своїми.
1KGS|16|27|А решта діл Омрі, що робив він, та лицарськість його, яку він чинив був, ото вони написані в Книзі Хроніки Ізраїлевих царів.
1KGS|16|28|І спочив Омрі з своїми батьками, і був похований у Самарії. А замість нього зацарював його син Ахав.
1KGS|16|29|Ахав, син Омрі, зацарював над Ізраїлем у році тридцятому й восьмому Аси, царя Юдиного. І царював Ахав, син Омрі, над Ізраїлем у Самарії двадцять і два роки.
1KGS|16|30|І робив Ахав, син Омрі, зло в Господніх очах більше від усіх, хто був перед ним.
1KGS|16|31|І було йому мало ходити в гріхах Єровоама, Неватового сина, і він узяв за жінку Єзавель, дочку Етбаала, сидонського царя. І він пішов, і служив Ваалові, і вклонявся йому.
1KGS|16|32|І він поставив жертівника для Ваала в Вааловому домі, якого збудував у Шомероні.
1KGS|16|33|І зробив Ахав Астарту. І Ахав далі чинив, щоб гнівити Господа, Бога Ізраїлевого, більше від усіх Ізраїлевих царів, що були перед ним.
1KGS|16|34|За його днів Хіїл з Бет-Елу відбудував Єрихона, на перворіднім своїм Авірамові він заклав його фундаменти, а на наймолодшім своїм Сеґівові повставляв брами його, за словом Господа, що говорив через Ісуса, Навинового сина.
1KGS|17|1|І сказав тішб'янин Ілля, з ґілеадських мешканців, до Ахава: Як живий Господь, Бог Ізраїлів, що перед лицем Його я стою, цими роками не буде роси та дощу, але тільки за моїм словом!
1KGS|17|2|І було до нього слово Господнє, говорячи:
1KGS|17|3|Іди звідси, й обернешся собі на схід, і сховаєшся при потоці Керіті, що навпроти Йордану.
1KGS|17|4|І станеться, будеш ти пити з потоку, а крукам наказав Я годувати тебе там.
1KGS|17|5|І він пішов, і зробив за Господнім словом: і пішов, й осівся при потоці Керіті, що навпроти Йордану.
1KGS|17|6|А круки приносили йому хліба та м'яса вранці, і хліба та м'яса ввечорі, а з потоку він пив.
1KGS|17|7|І сталося на кінці днів, і висох потік, бо в краю не було дощу.
1KGS|17|8|І було Господнє слово до нього, говорячи:
1KGS|17|9|Устань, іди до Сарепти сидонської, й осядеш там. Ось наказав Я там одній вдові, щоб годувала тебе.
1KGS|17|10|І він устав та й пішов до Сарепти. І прибув він до входу міста, аж ось там збирає дрова одна вдова. І він кликнув до неї й сказав: Візьми мені трохи води до посудини, й я нап'юся.
1KGS|17|11|І пішла вона взяти. А він кликнув до неї й сказав: Візьми мені й шматок хліба в свою руку!
1KGS|17|12|А та відказала: Як живий Господь, Бог твій, не маю я калача, а тільки повну пригорщу борошна в дзбанку та трохи олії в горняті. А оце я назбираю дві полінці дров, і піду, і приготовлю це собі та синові своєму. І з'їмо ми, та й помремо...
1KGS|17|13|І сказав до неї Ілля: Не бійся! Піди, зроби за своїм словом. Тільки спочатку зроби мені з того малого калача, і винесеш мені, а для себе та для сина свого зробиш потім.
1KGS|17|14|Бо так сказав Господь, Бог Ізраїлів: Дзбанок муки не скінчиться, і не забракне в горняті олії аж до дня, як Господь дасть дощу на поверхню землі.
1KGS|17|15|І пішла вона, із зробила за словом Іллі, і їла вона й він та її дім довгі дні,
1KGS|17|16|дзбанок муки не скінчився, і не забракло в горняті олії, за словом Господа, що говорив через Іллю.
1KGS|17|17|І сталося по тих пригодах, заслаб був син тієї жінки, господині того дому. І була його хвороба дуже тяжка, аж духу не позосталося в ньому.
1KGS|17|18|І сказала вона до Іллі: Що тобі до мене, чоловіче Божий? Прийшов ти до мене, щоб згадувати мій гріх та щоб убити мого сина!...
1KGS|17|19|І сказав він до неї: Дай мені сина свого! І він узяв його з лоня її, і виніс його в горницю, де він сидів, і поклав його на своєму ліжку.
1KGS|17|20|І кликнув він до Господа й сказав: Господи, Боже мій, чи й цій удові, що я в неї мешкаю, учиниш зло, щоб убити її сина?
1KGS|17|21|І витягся він тричі над дитиною, і кликав до Господа та казав: Господи, Боже мій, нехай вернеться душа цієї дитини в неї!
1KGS|17|22|І вислухав Господь голоса Іллі, і вернулася душа дитини в неї, і вона ожила...
1KGS|17|23|І взяв Ілля дитину, і зніс її з горниці додолу, і віддав її матері її. І сказав Ілля: Дивися, твій син живий!
1KGS|17|24|І сказала та жінка до Іллі: Тепер то я знаю, що ти Божий чоловік, а Господнє слово в устах твоїх правда!
1KGS|18|1|І минуло багато днів, і було Господнє слово до Іллі третього року, говорячи: Іди, покажися до Ахава, а Я дам дощ на поверхню землі.
1KGS|18|2|І пішов Ілля показатися до Ахава. А в Асирії був сильний голод.
1KGS|18|3|І покликав Ахав Овдія, що був над домом, а Овдій був дуже богобійний.
1KGS|18|4|І сталося, коли Єзавель вигублювала Господніх пророків, то Овдій узяв сотню пророків, та й сховав їх по п'ятидесяти чоловіка в печері, і годував їх хлібом та водою.
1KGS|18|5|І сказав Ахав до Овдія: Іди по Краю до всіх водних джерел та до всіх потоків, може знайдемо трави, і позоставимо при житті коня та мула, і не вигубимо худоби..
1KGS|18|6|І поділили вони собі Край, щоб перейти по ньому, Ахав пішов однією дорогою сам, Овдій пішов сам другою дорогою.
1KGS|18|7|І був Овдій у дорозі, аж ось Ілля назустріч йому. І пізнав він його, і впав на обличчя своє та й сказав: Чи то ти, пане мій Іллє?
1KGS|18|8|А той відказав йому: Я. Іди, скажи панові своєму: Ось тут Ілля!
1KGS|18|9|А він сказав: Чим я прогрішив, що ти віддаєш свого раба в Ахавову руку, щоб він убив мене?
1KGS|18|10|Як живий Господь, Бог твій, немає народу та царства, що туди не посилав би пан мій шукати тебе. А коли говорили: Нема його, то він заприсягав те царство та той народ, що знайдуть тебе.
1KGS|18|11|А тепер ти говориш: Іди, скажи своєму панові: Ось тут Ілля!
1KGS|18|12|І станеться, я піду від тебе, а Дух Господній понесе тебе на те місце, якого не знаю. І прийду я, щоб донести Ахаву, а коли він не знайде тебе, то вб'є мене. А раб твій боїться Господа від своєї молодости.
1KGS|18|13|Чи ж не було сказано панові моєму те, що зробив я, коли Єзавель побивала Господніх пророків, а я сховав був із Господніх пророків сотню чоловіка, по п'ятидесяти чоловіка в печері, і годував їх хлібом та водою?
1KGS|18|14|А тепер ти кажеш: Іди, скажи своєму панові: Ось тут Ілля, і він мене вб'є!...
1KGS|18|15|Та Ілля відказав: Як живий Господь Саваот, що я стою перед Його лицем, сьогодні я покажуся йому!
1KGS|18|16|І пішов Овдій назустріч Ахаву, та й доніс йому те. І пішов Ахав навпроти Іллі.
1KGS|18|17|І сталося, коли Ахав побачив Іллю, то Ахав сказав до нього: Чи це ти, що непокоїш Ізраїля?
1KGS|18|18|А той відказав: Не я внещасливив Ізраїля, а тільки ти та дім твого батька через ваше недотримання Господніх заповідей, та й ти пішов за Ваалами.
1KGS|18|19|А тепер пошли, збери до мене на гору Кармел усього Ізраїля та чотири сотні й п'ятдесят Ваалових пророків, та чотири сотні пророків Астарти, що їдять зо столу Єзавелі.
1KGS|18|20|І послав Ахав по всіх Ізраїлевих синах, і зібрав пророків на гору Кармел.
1KGS|18|21|І підійшов Ілля до всього народу й сказав: Чи довго ви будете скакати на двох галузках? Якщо Господь Бог, ідіть за Ним, а якщо Ваал ідіть за ним! Та не відповів йому народ ані слова.
1KGS|18|22|І сказав Ілля до народу: Я сам позостався Господній пророк, а пророків Ваалових чотири сотні й п'ятдесят чоловіка.
1KGS|18|23|І нехай дадуть нам двох бичків, і нехай вони виберуть собі одного бичка, і нехай заріжуть його, і нехай покладуть на дрова, а огню не покладуть. І я приготую одного бичка, і дам на дрова, а огню не покладу.
1KGS|18|24|І ви покличете ім'я бога вашого, а я покличу Ім'я Господа. І станеться, той Бог, що відповість огнем, Він Бог! І відповів той народ та й сказав: Це добре слово!
1KGS|18|25|І сказав Ілля до Ваалових пророків: Виберіть собі одного бичка, і приготуйте перші, бо ви численніші, і покличте ім'я свого бога, і огню не покладете.
1KGS|18|26|І взяли вони того бичка, що він дав їм, і вони приготували й кликали Ваалове ім'я від ранку й аж до полудня, говорячи: Ваале, почуй нас! Та не було ані голосу, ані відповіді. І скакали вони біля жертівника, що зробили.
1KGS|18|27|І сталося опівдні, і сміявся з них Ілля й говорив: Кличте голосом сильнішим, бо він бог! Може він роздумує, або відлучився, або в дорозі! Може він спить, то прокинеться!
1KGS|18|28|І стали вони кликати голосом сильнішим, і кололися, за своїм звичаєм, мечами та ратищами, аж лилася з них кров.
1KGS|18|29|І сталося, як минувся південь, то вони пророкували аж до часу принесення хлібної жертви, та не було ані голосу, ані відповіді, ані слуху...
1KGS|18|30|І сказав Ілля до всього народу: Підійдіть до мене! І підійшов увесь народ до нього, а він поправив розбитого Господнього жертівника.
1KGS|18|31|І взяв Ілля дванадцятеро каміння, за числом племен синів Якова, до якого було слово Господнє, говорячи: Ізраїль буде ім'я твоє!
1KGS|18|32|і збудував із того каміння жертівника в Ім'я Господнє, і зробив рова, площею на дві саті насіння, навколо жертівника.
1KGS|18|33|І наклав дров, і зарізав бичка та й поклав на дровах.
1KGS|18|34|І він сказав: Наповніть чотири відрі води, і нехай виллють на цілопалення та на дрова. І сказав: Повторіть! І повторили. І сказав: Зробіть утретє! І зробили втретє.
1KGS|18|35|І потекла вода навколо жертівника, а також рів наповнився водою.
1KGS|18|36|І сталося в час принесення хлібної жертви, що підійшов пророк Ілля та й сказав: Господи, Боже Авраамів, Ісаків та Ізраїлів! Сьогодні пізнають, що Ти Ізраїлів Бог, а я Твій раб, і що все оце я зробив Твоїм словом.
1KGS|18|37|Вислухай мене, Господи, вислухай мене, і нехай пізнає цей народ, що Ти Господь, Бог, і Ти обернеш їхнє серце назад!
1KGS|18|38|І спав Господній огонь, та й пожер цілопалення, і дрова, і каміння, і порох, і вилизав воду, що в рові...
1KGS|18|39|І побачили це всі люди, та й попадали на обличчя свої й говорили: Господь, Він Бог, Господь, Він Бог!
1KGS|18|40|І сказав до них Ілля: Схопіть Ваалових пророків! Нехай ніхто не втече з них! І похапали їх, а Ілля звів їх до потоку Кішон, та й порізав їх...
1KGS|18|41|І сказав Ілля до Ахава: Увійди, їж і пий, бо ось чути шум дощу.
1KGS|18|42|І пішов Ахав, щоб їсти та пити, а Ілля зійшов на верхів'я Кармелу, і нахилився до землі, і поклав обличчя своє між свої коліна.
1KGS|18|43|І сказав він до свого хлопця: Вийди, подивися в напрямі моря! І той вийшов і подивився та й сказав: Нема нічого. Та він відказав: Вернися сім раз!
1KGS|18|44|І сталося сьомого разу, і він сказав: Ось мала хмара, немов долоня людська, підіймається з моря. А він сказав: Піди, скажи Ахавові: Запрягай і зійди, і не затримає тебе дощ.
1KGS|18|45|І сталося по недовгому часі, і потемніло небо від хмар, і зірвався вітер, і пішов великий дощ. А Ахав сів на воза, та й відправився в Їзреел.
1KGS|18|46|А Господня рука була на Іллі. І він оперезав свої стегна, та й побіг перед Ахавом аж до самого Їзреелу.
1KGS|19|1|А Ахав доніс Єзавелі все, що зробив був Ілля, і все те, що він повбивав усіх пророків мечем.
1KGS|19|2|І послала Єзавель посланця до Іллі, говорячи: Отак нехай зроблять мені боги, і так нехай додадуть, якщо цього часу взавтра я не зроблю душі твоїй, як зроблено душі кожного з них!
1KGS|19|3|І побачив він це, і встав та й пішов, боячись за душу свою. І прийшов він до Юдиної Беер-Шеви, і позоставив там свого хлопця.
1KGS|19|4|А сам пішов пустинею, дорогою одного дня, і сів під одним ялівцем, і зажадав собі смерти, і сказав: Досить тепер, Господи! Візьми душу мою, бо я не ліпший від батьків своїх!...
1KGS|19|5|І поклався він, і заснув під одним ялівцем. Аж ось Ангол діткнувся його та й сказав йому: Устань та попоїж!
1KGS|19|6|І глянув він, аж ось у його головах калач, спечений на вугіллі, та дзбанок води. І він їв та пив, і знову поклався.
1KGS|19|7|І вернувся Ангол Господній удруге, і діткнувся його та й сказав: Устань, попоїж, бо дорога тяжка перед тобою.
1KGS|19|8|І він устав, і попоїв та напився. І він ішов, підкріплений тією їжею, сорок день та сорок ночей аж до Божої гори Хорив.
1KGS|19|9|І прибув він туди до печери, і переночував там, аж ось Господнє слово до нього. І сказав Він йому: Чого ти тут, Іллє?
1KGS|19|10|А той відказав: Я був дуже горливий для Господа, Бога Саваота, бо Ізраїлеві сини покинули заповіта Твого та порозбивали жертівники Твої, а пророків Твоїх повбивали мечем, і позостався я сам. І шукали вони душу мою, щоб узяти її.
1KGS|19|11|А Він відказав: Вийди, і станеш на горі перед Господнім лицем. Аж ось переходитиме Господь, а перед Господнім лицем вітер великий та міцний, що зриває гори та скелі ламає. Та не в вітрі Господь. А по вітрі трус землі, та не в трусі Господь.
1KGS|19|12|А по трусі огонь, і не в огні Господь. А по огні тихий лагідний голос.
1KGS|19|13|І сталося, як почув це Ілля, то закрив своє обличчя плащем своїм, та й вийшов, і став у входа печери. Аж ось до нього Голос, що говорив: Чого ти тут, Іллє?
1KGS|19|14|А він відказав: Я був дуже горливий для Господа, Бога Саваота, бо Ізраїлеві сини покинули заповіта Твого та порозбивали жертівники твої, а пророків Твоїх повбивали мечем, і позостався я сам. І шукали вони душу мою, щоб узяти її.
1KGS|19|15|І сказав до нього Господь: Іди, вернися на свою дорогу на Дамаську пустиню. І прийдеш, і помажеш Хазаїла на царя над Сирією.
1KGS|19|16|А Єгу, Німшієвого сина, помажеш на царя над Ізраїлем, а Єлисея, Шафатового сина з Авел-Мехоли, помажеш на пророка замість себе.
1KGS|19|17|І станеться, хто втече від Хазаїлового меча, того вб'є Єгу, а хто втече від меча Єгу, того вб'є Єлисей.
1KGS|19|18|А в Ізраїлі Я позоставив сім тисяч, усі коліна, що не схилялися перед Ваалом, та всі уста, що не цілували його.
1KGS|19|19|І пішов він ізвідти, і знайшов Єлисея, Шафатового сина, а він оре. Дванадцять запрягів перед ним, а він при дванадцятому. І підійшов до нього Ілля та й кинув йому свого плаща.
1KGS|19|20|І позоставив той волів, та й побіг за Іллею й сказав: Нехай поцілую я батька свого та свою матір, та й піду за тобою! А той відказав йому: Іди, але вернися, бо що я зробив тобі?
1KGS|19|21|І вернувся він від нього, і взяв запряга волів та й приніс його в жертву, а ярмами волів зварив його м'ясо, і дав народові, а ті їли. І він устав, і пішов за Іллею, та й служив йому.
1KGS|20|1|А Бен-Гадад, цар сирійский, зібрав усе своє військо та тридцять і два царі з ним, і коні, і колесниці. І пішов він, і обліг Самарію та й воював проти неї.
1KGS|20|2|І послав він послів до Ахава, царя Ізраїлевого, до міста,
1KGS|20|3|та й сказав йому: Так сказав Бен-Гадад: Срібло твоє та золото твоє моє воно, а жінки твої та сини твої, ці найліпші, мої вони!
1KGS|20|4|І відповів Ізраїлів цар та й сказав: Буде за словом твоїм, пане мій царю! Твій я та все, що моє!
1KGS|20|5|І знову вернулися ті посли та й сказали: Так сказав Бен-Гадад, говорячи: Я посилав до тебе, говорячи: Ти даси мені срібло своє, і золото своє, і жінок своїх, і синів своїх.
1KGS|20|6|А взавтра цього часу пошлю я своїх рабів до тебе, і вони перешукають дім твій та доми твоїх рабів. І станеться, на все, що сподобається їм, вони накладуть свої руки, та й заберуть...
1KGS|20|7|І скликав Ізраїлів цар усіх старших Краю та й сказав: Довідайтеся й побачите, що він шукає зла, бо послав до мене по жінок моїх, і по синів моїх, і по срібло моє, і по золото моє, і я йому не відмовив.
1KGS|20|8|І сказали до нього всі старші та ввесь народ: Не слухай, і не погоджуйся!
1KGS|20|9|І сказав він до послів Бен-Гадада: Скажіть моєму панові цареві: Усе, про що посилав ти до свого раба напочатку, я зроблю, а цієї речі зробити не можу. І пішли посли, і віднесли йому відповідь.
1KGS|20|10|І послав до нього Бен-Гадад та й сказав: Нехай так зроблять мені боги, і нехай так додадуть, якщо самарійського пороху вистачить по жмені всьому народові, що стоїть при мені!...
1KGS|20|11|І відповів Ізраїлів цар та й сказав: Кажіть: Хай не хвалиться той, хто меча припинає, а той, хто розв'язує!
1KGS|20|12|І сталося, як почув він цю відповідь, а він пив, він та царі в шатрах, то сказав до своїх рабів: Пустіть тарани! І вони пустили тарани на місто.
1KGS|20|13|Аж ось один пророк підійшов до Ахава, Ізраїлевого царя, та й сказав: Так сказав Господь: Чи бачив ти ввесь оцей великий натовп? Ось Я даю його сьогодні в руку твою, і ти пізнаєш, що Я Господь!
1KGS|20|14|І сказав Ахав: Ким? А той відказав: Так сказав Господь: Слугами начальників округ. І сказав: Хто розпічне війну? А той відказав: Ти.
1KGS|20|15|І перелічив він слуг начальників судових округ, і було дві сотні й тридцять два. А по них перелічив увесь народ, усіх Ізраїлевих синів, сім тисяч.
1KGS|20|16|І вийшли вони опівдні, а Бен-Гадад пив п'яний у шатрах, він та царі, тридцять і два царі, що допомагали йому.
1KGS|20|17|І вийшли напочатку слуги начальників округ. І послав Бен-Гадад, і донесли йому, кажучи: Ось повиходили люди з Самарії.
1KGS|20|18|А він відказав: Якщо на мир вийшли вони, схопіть їх живих, а якщо на війну повиходили, теж живими схопіть їх у неволю!
1KGS|20|19|А то вийшли з міста слуги начальників округ та військо, що йшло за ними.
1KGS|20|20|І побивали вони один одного, і побігли сиріяни, а Ізраїль їх гнав. Та втік Бен-Гадад, сирійський цар, на коні та з верхівцями.
1KGS|20|21|І вийшов Ізраїлів цар, та й побив коні та колесниці, і завдав в Сирії великої поразки.
1KGS|20|22|І підійшов пророк до Ізраїлевого царя та й сказав йому: Іди, тримайся мужньо, і пізнай та побач, що ти зробиш, бо, як мине рік, сирійський цар знову піде на тебе.
1KGS|20|23|А слуги сирійського царя сказали йому: Бог гір їхній Бог, тому вони були сильніші від нас. Але воюймо з ними на рівнині, присягаємо, що будемо сильніші від них!
1KGS|20|24|І зроби цю річ: Поскидай тих царів, кожного з його місця, і понаставляй намісників замість них.
1KGS|20|25|А ти збереш собі військо, як те, що відпало від тебе, і коней, скільки було коней, і колесниць, скільки було колесниць, і будемо воювати з ними на рівнині. Присягаємо, що ми будемо сильніші від них! І він послухався їхнього голосу, і зробив так.
1KGS|20|26|І сталося по році, і Бен-Гадад переглянув Сирію, і пішов до Афеку на війну з Ізраїлем.
1KGS|20|27|А Ізраїлеві сини були переглянені й забезпечені живністю, та й вийшли навпроти них. І таборували Ізраїлеві сини навпроти них, як дві отарі кіз, а сиріяни наповнили Край.
1KGS|20|28|І підійшов Божий чоловік, і говорив до Ізраїлевого царя та й сказав: Так сказав Господь: Тому, що сказали сиріяни: Господь Бог гір, а не Бог долин Він, то дам увесь цей великий натовп у твою руку, і ви пізнаєте, що Я Господь!
1KGS|20|29|І таборували ті навпроти тих сім день. І сталося сьомого дня, і розпалився бій, і побили Ізраїлеві сини Сирію, сто тисяч піхоти, одного дня.
1KGS|20|30|А позосталі повтікали до Афеку, до міста, та впав мур на двадцять і сім тисяч позосталих чоловіка. А Бен-Гадад утік і ввійшов до міста, до внутрішньої кімнати.
1KGS|20|31|І сказали до нього його слуги: Ось ми чули, що царі Ізраїлевого дому вони царі милостиві. Покладім веретища на стегна свої, а шнури на свої голови, і вийдім до Ізраїлевого царя, може він пощадить твою душу.
1KGS|20|32|І підперезали вони веретищами стегна свої, а шнури на свої голови, і прийшли до Ізраїлевого царя та й сказали: Твій раб Бен-Гадад сказав: Нехай живе душа моя! А той відказав: Чи він іще живий? Він мій брат!
1KGS|20|33|А ті люди взяли це за натяка, і поспішили скористатися з того й сказали: Брат твій Бен-Гадад! І той відказав: Підіть, приведіть його! І вийшов до нього Бен-Гадад, а той посадив його на колесницю.
1KGS|20|34|І сказав до нього Бен-Гадад: Ті міста, що батько мій був забрав від твого батька, я поверну. І ти урядиш собі в Дамаску вулиці, як мій батько урядив був у Самарії. А Я сказав Ахав по умові відпущу тебе. І він склав з ним умову, та й відпустив його.
1KGS|20|35|Тоді один чоловік із пророчих синів сказав до свого ближнього за Господнім словом: Удар мене! Та відмовився той чоловік ударити його.
1KGS|20|36|І сказав він йому: За те, що ти не послухався Господнього голосу, то ось ти підеш від мене і вб'є тебе лев! І пішов той від нього, і спіткав його лев та й забив.
1KGS|20|37|І знайшов він іншого чоловіка та й сказав: Удар мене! І той чоловік ударив його, ударив та й зранив.
1KGS|20|38|І пішов той пророк, і став цареві на дорозі, і перебрався, і закрив хусткою очі свої.
1KGS|20|39|І сталося, цар проходив, а він кричав до царя й говорив: Раб твій ввійшов у середину бою. Аж ось один чоловік відійшов, і підвів до мене мужа й сказав: Пильнуй цього мужа! Якщо його не стане, то буде твоє життя замість його життя, або відважиш таланта срібла.
1KGS|20|40|І сталося, раб твій робив тут та тут, а він зник. І сказав до нього Ізраїлів цар: Такий твій присуд, ти сам проказав.
1KGS|20|41|А той спішно зняв хустку з-над очей своїх, і пізнав його Ізраїлів цар, що він із пророків.
1KGS|20|42|А той йому сказав: Так сказав Господь: Тому, що ти випустив із руки чоловіка, Мені призначеного, то буде життя твоє за його життя, а народ твій за його народ!...
1KGS|20|43|І пішов Ізраїлів цар до свого дому незадоволений та гнівний, і прибув у Самарію.
1KGS|21|1|І сталося по цих пригодах таке. У їзреелянина Навота, що в Їзреелі, був виноградник при палаті Ахава, самарійського царя.
1KGS|21|2|І говорив Ахав до Навота, кажучи: Дай мені свого виноградника, і він буде мені за яринного города, бо він близький до мого дому. А я дам тобі замість нього виноградника ліпшого від нього. Якщо це добре в очах твоїх, я дам тобі срібла, ціну його.
1KGS|21|3|І сказав Навот до Ахава: Заборонено мені від Господа, щоб я дав тобі спадщину моїх батьків.
1KGS|21|4|І ввійшов Ахав до дому свого незадоволений та гнівний через те слово, яке говорив йому їзреелянин Навот, бо той сказав: Не дам тобі спадщини батьків моїх! І ліг він на ліжку своїм, і відвернув своє обличчя, і не їв хліба.
1KGS|21|5|І прийшла до нього жінка його Єзавель та й сказала йому: Чого це твій дух сумний, і ти не їси хліба?
1KGS|21|6|І сказав він до неї: Бо я говорив до їзреелянина Навота. І сказав я йому: Дай мені свого виноградника за срібло, або, якщо ти хочеш, дам тобі замість нього виноградника ліпшого. Та він відказав: Не дам тобі свого виноградника!
1KGS|21|7|І сказала до нього його жінка Єзавель: Отепер ти зробишся царем над Ізраїлем. Устань, поїж хліба, і нехай буде веселе твоє серце. А виноградника їзреелянина Навота дам тобі я.
1KGS|21|8|І понаписувала вона листи в імені Ахава, і позапечатувала їх його печаткою, та й порозсилала ті листи до старших та до вельможних, що були в його місті, що сиділи з Навотом.
1KGS|21|9|А в тих листах вона понаписувала так: Оголосіть піст, і посадіть Навота на чолі народу.
1KGS|21|10|І посадіть двох негідних людей навпроти нього, нехай свідчать на нього, кажучи: Ти зневажив Бога й царя. І виведіть його, і вкаменуйте його, і нехай він помре...
1KGS|21|11|І зробили мужі його міста, старші та вельможні, що сиділи в його місті, так, як послала до них Єзавель, як було написано в листах, які вона порозсилала до них.
1KGS|21|12|Оголосили вони піст, і посадили Навота на чолі народу.
1KGS|21|13|І прийшли два чоловіки негідні, і сіли навпроти нього. І ті негідні люди свідчили на нього, на Навота, перед народом, говорячи: Навот зневажив Бога й царя! І вивели його поза місто, та й укаменували його камінням, і він помер...
1KGS|21|14|І послали вони до Єзавелі, говорячи: Навот укаменований і помер.
1KGS|21|15|І сталося, як почула Єзавель, що Навот укаменований і помер, то сказала Єзавель до Ахава: Устань, посядь виноградника їзреелянина Навота, що відмовив дати його тобі за срібло, бо Навот не живий, а помер.
1KGS|21|16|І сталося, як почув Ахав, що Навот помер, то Ахав устав, щоб зійти до виноградника їзреелянина Навота, щоб посісти його.
1KGS|21|17|І було Господнє слово до тішб'янина Іллі, говорячи:
1KGS|21|18|Устань, зійди назустріч Ахава, Ізраїлевого царя, що в Сирії, ось він у Навотовому винограднику, куди зійшов, щоб посісти його.
1KGS|21|19|І будеш говорити до нього, кажучи: Так сказав Господь: Ти вбив, а тепер хочеш посісти? І говоритимеш до нього, кажучи: Так сказав Господь: На тому місці, де пси лизали Навотову кров, пси лизатимуть і твою власну кров!
1KGS|21|20|І сказав Ахав до Іллі: Ось ти знайшов мене, вороже мій! А той відказав: Знайшов, бо ти запродався чинити зло в Господніх очах.
1KGS|21|21|Ось Я спроваджую на тебе лихо, і вигублю все за тобою, і вигублю Ахавові навіть те, що мочить на стіну, і невільного та вільного в Ізраїлі!
1KGS|21|22|І зроблю з твоїм домом, як із домом Єровоама, Неватового сина, й як із домом Баші, Ахієвого сина, за той гнів, яким розгнівив ти Мене та ввів у гріх Ізраїля.
1KGS|21|23|І також до Єзавелі говорив Господь, кажучи: Пси з'їдять Єзавель на передмур'ї Їзреелу.
1KGS|21|24|Померлого в Ахава в місті поїдять пси, а померлого на полі поїсть птаство небесне.
1KGS|21|25|Бо ще не було такого, як Ахав, що запродався чинити зло в Господніх очах, що його намовила жінка його Єзавель.
1KGS|21|26|І він чинив дуже гидке, ідучи за ідолами, усе так, як робили амореяни, що їх Господь повиганяв перед Ізраїлевими синами.
1KGS|21|27|І сталося, як Ахав почув ці слова, то роздер він шати свої, і зодягнув на тіло своє веретище, і постив, і лежав у веретищі, і ходив сумовито...
1KGS|21|28|І було Господнє слово до тішб'янина Іллі, говорячи:
1KGS|21|29|Чи ти спостеріг, що Ахав упокорився перед лицем Моїм? За те, що він упокорився перед Моїм лицем, не наведу Я лиха за його днів, за днів його сина наведу Я те лихо на його дім.
1KGS|22|1|І прожили вони три роки, і не було війни між Сирією та між Ізраїлем.
1KGS|22|2|І сталося третього року, і зійшов Йосафат, цар Юдин, до Ізраїлевого царя.
1KGS|22|3|І сказав Ізраїлів цар до своїх слуг: Чи ви знаєте, що ґілеадський Рамот наш? А ми мовчимо, замість того, щоб забрати його з руки сирійського царя.
1KGS|22|4|І сказав він до Йосафата: Чи ти підеш зо мною на війну до ґілеадського Рамоту? А Йосафат відказав: Я як ти, народ мій як народ твій, мої коні як твої коні!
1KGS|22|5|І сказав Йосафат до Ізраїлевого царя: Вивідай зараз слово Господнє!
1KGS|22|6|І зібрав Ізраїлів цар пророків, близько чотирьох сотень чоловіка, та й сказав до них: Чи йти мені на війну на ґілеадський Рамот, чи занехати? А ті відказали: Іди, а Господь дасть його в цареву руку.
1KGS|22|7|І сказав Йосафат: Чи нема тут іще Господнього пророка, і вивідаємо від нього.
1KGS|22|8|І сказав Ізраїлів цар до Йосафата: Є ще один муж, щоб від нього вивідати Господа. Та я ненавиджу його, бо він не пророкує на мене добре, а тільки зле. Це Міхей, син Їмлин. А Йосафат відказав: Нехай цар не говорить так!
1KGS|22|9|І покликав Ізраїлів цар одного євнуха, і сказав: Приведи скоріш Міхея, Їмлиного сина!
1KGS|22|10|І цар Ізраїлів та цар Юдин сиділи кожен на троні своїм, повбирані в шати при вході до брами Самарії, а всі пророки пророкували перед ними.
1KGS|22|11|А Седекія, Кенаанин син, зробив собі залізні роги й сказав: Так сказав Господь: Оцим будеш побивати сиріян аж до вигублення їх!
1KGS|22|12|І всі пророки пророкували так, говорячи: Виходь до ґілеадського Рамоту, і пощастить тобі, і Господь дасть його в цареву руку.
1KGS|22|13|А той посланець, що пішов покликати Міхея, говорив до нього, кажучи: Ось слова тих пророків, одноусто звіщають цареві добро. Нехай же буде слово твоє, як слово кожного з них, і ти говоритимеш добре.
1KGS|22|14|І сказав Міхей: Як живий Господь, те, що скаже мені Господь, я те говоритиму!
1KGS|22|15|І прийшов він до царя, а цар сказав до нього: Міхею, чи підемо на війну до ґілеадського Рамоту, чи занехаємо? А той відказав йому: Вийди, і пощастить тобі, і Господь дасть у цареву руку.
1KGS|22|16|І сказав йому цар: Аж скільки разів я заприсягав тебе, що ти не говоритимеш мені нічого, тільки правду в Ім'я Господа?
1KGS|22|17|А той відказав: Я бачив усього Ізраїля, розпорошеного по горах, немов овець, що не мають пастуха. І сказав Господь: Немає в них пана, нехай вернуться з миром кожен до дому свого.
1KGS|22|18|І сказав Ізраїлів цар до Йосафата: Чи ж не казав я тобі, він не буде пророкувати мені доброго, а тільки лихе?
1KGS|22|19|А Міхей відказав: Тому послухай Господнього слова: Бачив я Господа, що сидів на престолі Своїм, а все небесне військо стояло при Ньому з правиці Його та з лівиці Його.
1KGS|22|20|І сказав Господь: Хто намовить Ахава, і він вийде й упаде в ґілеадському Рамоті? І говорив той так, а той говорив так.
1KGS|22|21|І вийшов дух, і став перед Господнім лицем та й сказав: Я намовлю його! І сказав йому Господь: Чим?
1KGS|22|22|А той відказав: Я вийду й стану духом неправди в устах усіх його пророків. А Господь сказав: Ти намовиш, а також переможеш; вийди та й зроби так!
1KGS|22|23|А тепер оце Господь дав духа неправди в уста всіх оцих пророків, а Господь говорив на тебе лихе...
1KGS|22|24|І підійшов Седекія, Кенаанин син, і вдарив Міхея по щоці та й сказав: Кудою це перейшов Дух Господній від мене, щоб говорити з тобою?
1KGS|22|25|А Міхей сказав: Ось ти побачиш це, коли вбіжиш до найдальшої кімнати, щоб сховатися.
1KGS|22|26|І сказав Ізраїлів цар: Візьми Міхея, і відведи до Амона, начальника міста, та до Йоаша, царевого сина,
1KGS|22|27|та й скажеш: Отак сказав цар: Посадіть оцього до в'язничного дому, і давайте йому їсти скупо хліба й скупо води, аж поки я не вернуся з миром.
1KGS|22|28|А Міхей відказав: Якщо справді вернешся ти з миром, то не говорив Господь через мене! І до того сказав: Слухайте це, всі народи!
1KGS|22|29|І вийшов Ізраїлів цар та Йосафат, цар Юдин, до ґілеадського Рамоту.
1KGS|22|30|І сказав Ізраїлів цар до Йосафата: Я переберуся, і піду на бій, а ти вбери свої царські шати! І перебрався Ізраїлів цар, і пішов на бій.
1KGS|22|31|А сирійський цар наказав керівникам своїх колесниць, тридцятьом і двом, говорячи: Не будете воювати з малим та з великим, а тільки з самим Ізраїлевим царем.
1KGS|22|32|І сталося, як керівники колесниць побачили Йосафата, то вони сказали: Це дійсно Ізраїлів цар! І зайшли на нього, щоб воювати, а Йосафат закричав.
1KGS|22|33|І сталося, як керівники колесниць побачили, що це не Ізраїлів цар, то повернули від нього.
1KGS|22|34|А один чоловік знехотя натягнув лука, та й ударив Ізраїлевого царя між підв'язанням пояса та між панцерем. А той сказав своєму візникові: Поверни назад, і виведи мене з табору, бо я ранений...
1KGS|22|35|І знявся бій того дня, а цар був поставлений на колесниці проти Сирії, і помер увечорі. І кров із рани текла в колесницю.
1KGS|22|36|А як сонце заходило, нісся крик у таборі такий: Кожен до міста свого, і кожен до краю свого!
1KGS|22|37|І помер цар, і був привезений до Самарії. І поховали царя в Самарії.
1KGS|22|38|І полоскали колесницю над ставом у Самарії, і пси лизали його кров, а блудниці мили своє тіло, за словом Господнім, що Він говорив.
1KGS|22|39|А решта Ахавових діл, і все, що він зробив був, і дім зо слонової кости, що він збудував, і всі міста, які він побудував, отож вони написані в Книзі Хроніки Ізраїлевих царів.
1KGS|22|40|І спочив Ахав із батьками своїми, а замість нього зацарював син його Ахазія.
1KGS|22|41|А Йосафат, Асин син, зацарював над Юдою в четвертому році Ахава, царя Ізраїлевого.
1KGS|22|42|Йосафат був віку тридцяти й п'яти літ, коли він зацарював, і двадцять і п'ять літ царював в Єрусалимі. А ім'я його матері Азува, дочка Шілхи.
1KGS|22|43|І ходив він усією дорогою батька свого Аси, і не збочував із неї, щоб чинити добре в Господніх очах. Тільки пагірки не були понищені, народ іще приносив жертви й кадив на пагірках.
1KGS|22|44|І Йосафат замирив з Ізраїлевим царем.
1KGS|22|45|А решта Йосафатових діл та лицарськість його, що він чинив був та як воював, отож вони написані в Книзі Хроніки Юдиних царів.
1KGS|22|46|А решту блудодіїв, що позоставалися за днів його батька Аси, він вигубив із Краю.
1KGS|22|47|А царя не було в Едомі, був намісник царів.
1KGS|22|48|А Йосафат наробив був таршіських кораблів, щоб піти до Офіру по золото, та не пішов, бо порозбивалися кораблі при Ецйон-Ґевері.
1KGS|22|49|Тоді сказав Ахазія, син Ахавів, до Йосафата: Нехай підуть на кораблях мої раби з рабами твоїми. Та Йосафат не захотів.
1KGS|22|50|І спочив Йосафат із своїми батьками. І був він похований в Місті Давида, свого батька, а замість нього зацарював син його Єгорам.
1KGS|22|51|Ахазія, Ахавів син, зацарював над Ізраїлем у Самарії, в сімнадцятому році Йосафата, Юдиного царя, і царював над Ізраїлем два роки.
1KGS|22|52|І робив він лихе в Господніх очах, і ходив дорогою батька свого й дорогою своєї матері, та дорогою Єровоама, Неватового сина, що вводив у гріх Ізраїля.
1KGS|22|53|І служив він Ваалові, і вклонявся йому, та й гнівив Господа, Бога Ізраїлевого, усе так, як робив його батько.
