1SAM|1|1|There was a certain man from Ramathaim, a Zuphite from the hill country of Ephraim, whose name was Elkanah son of Jeroham, the son of Elihu, the son of Tohu, the son of Zuph, an Ephraimite.
1SAM|1|2|He had two wives; one was called Hannah and the other Peninnah. Peninnah had children, but Hannah had none.
1SAM|1|3|Year after year this man went up from his town to worship and sacrifice to the LORD Almighty at Shiloh, where Hophni and Phinehas, the two sons of Eli, were priests of the LORD.
1SAM|1|4|Whenever the day came for Elkanah to sacrifice, he would give portions of the meat to his wife Peninnah and to all her sons and daughters.
1SAM|1|5|But to Hannah he gave a double portion because he loved her, and the LORD had closed her womb.
1SAM|1|6|And because the LORD had closed her womb, her rival kept provoking her in order to irritate her.
1SAM|1|7|This went on year after year. Whenever Hannah went up to the house of the LORD, her rival provoked her till she wept and would not eat.
1SAM|1|8|Elkanah her husband would say to her, "Hannah, why are you weeping? Why don't you eat? Why are you downhearted? Don't I mean more to you than ten sons?"
1SAM|1|9|Once when they had finished eating and drinking in Shiloh, Hannah stood up. Now Eli the priest was sitting on a chair by the doorpost of the LORD's temple.
1SAM|1|10|In bitterness of soul Hannah wept much and prayed to the LORD.
1SAM|1|11|And she made a vow, saying, "O LORD Almighty, if you will only look upon your servant's misery and remember me, and not forget your servant but give her a son, then I will give him to the LORD for all the days of his life, and no razor will ever be used on his head."
1SAM|1|12|As she kept on praying to the LORD, Eli observed her mouth.
1SAM|1|13|Hannah was praying in her heart, and her lips were moving but her voice was not heard. Eli thought she was drunk
1SAM|1|14|and said to her, "How long will you keep on getting drunk? Get rid of your wine."
1SAM|1|15|"Not so, my lord," Hannah replied, "I am a woman who is deeply troubled. I have not been drinking wine or beer; I was pouring out my soul to the LORD.
1SAM|1|16|Do not take your servant for a wicked woman; I have been praying here out of my great anguish and grief."
1SAM|1|17|Eli answered, "Go in peace, and may the God of Israel grant you what you have asked of him."
1SAM|1|18|She said, "May your servant find favor in your eyes." Then she went her way and ate something, and her face was no longer downcast.
1SAM|1|19|Early the next morning they arose and worshiped before the LORD and then went back to their home at Ramah. Elkanah lay with Hannah his wife, and the LORD remembered her.
1SAM|1|20|So in the course of time Hannah conceived and gave birth to a son. She named him Samuel, saying, "Because I asked the LORD for him."
1SAM|1|21|When the man Elkanah went up with all his family to offer the annual sacrifice to the LORD and to fulfill his vow,
1SAM|1|22|Hannah did not go. She said to her husband, "After the boy is weaned, I will take him and present him before the LORD, and he will live there always."
1SAM|1|23|"Do what seems best to you," Elkanah her husband told her. "Stay here until you have weaned him; only may the LORD make good his word." So the woman stayed at home and nursed her son until she had weaned him.
1SAM|1|24|After he was weaned, she took the boy with her, young as he was, along with a three-year-old bull, an ephah of flour and a skin of wine, and brought him to the house of the LORD at Shiloh.
1SAM|1|25|When they had slaughtered the bull, they brought the boy to Eli,
1SAM|1|26|and she said to him, "As surely as you live, my lord, I am the woman who stood here beside you praying to the LORD.
1SAM|1|27|I prayed for this child, and the LORD has granted me what I asked of him.
1SAM|1|28|So now I give him to the LORD. For his whole life he will be given over to the LORD." And he worshiped the LORD there.
1SAM|2|1|Then Hannah prayed and said: "My heart rejoices in the LORD; in the LORD my horn is lifted high. My mouth boasts over my enemies, for I delight in your deliverance.
1SAM|2|2|"There is no one holy like the LORD; there is no one besides you; there is no Rock like our God.
1SAM|2|3|"Do not keep talking so proudly or let your mouth speak such arrogance, for the LORD is a God who knows, and by him deeds are weighed.
1SAM|2|4|"The bows of the warriors are broken, but those who stumbled are armed with strength.
1SAM|2|5|Those who were full hire themselves out for food, but those who were hungry hunger no more. She who was barren has borne seven children, but she who has had many sons pines away.
1SAM|2|6|"The LORD brings death and makes alive; he brings down to the grave and raises up.
1SAM|2|7|The LORD sends poverty and wealth; he humbles and he exalts.
1SAM|2|8|He raises the poor from the dust and lifts the needy from the ash heap; he seats them with princes and has them inherit a throne of honor. "For the foundations of the earth are the LORD's; upon them he has set the world.
1SAM|2|9|He will guard the feet of his saints, but the wicked will be silenced in darkness. "It is not by strength that one prevails;
1SAM|2|10|those who oppose the LORD will be shattered. He will thunder against them from heaven; the LORD will judge the ends of the earth. "He will give strength to his king and exalt the horn of his anointed."
1SAM|2|11|Then Elkanah went home to Ramah, but the boy ministered before the LORD under Eli the priest.
1SAM|2|12|Eli's sons were wicked men; they had no regard for the LORD.
1SAM|2|13|Now it was the practice of the priests with the people that whenever anyone offered a sacrifice and while the meat was being boiled, the servant of the priest would come with a three-pronged fork in his hand.
1SAM|2|14|He would plunge it into the pan or kettle or caldron or pot, and the priest would take for himself whatever the fork brought up. This is how they treated all the Israelites who came to Shiloh.
1SAM|2|15|But even before the fat was burned, the servant of the priest would come and say to the man who was sacrificing, "Give the priest some meat to roast; he won't accept boiled meat from you, but only raw."
1SAM|2|16|If the man said to him, "Let the fat be burned up first, and then take whatever you want," the servant would then answer, "No, hand it over now; if you don't, I'll take it by force."
1SAM|2|17|This sin of the young men was very great in the LORD's sight, for they were treating the LORD's offering with contempt.
1SAM|2|18|But Samuel was ministering before the LORD -a boy wearing a linen ephod.
1SAM|2|19|Each year his mother made him a little robe and took it to him when she went up with her husband to offer the annual sacrifice.
1SAM|2|20|Eli would bless Elkanah and his wife, saying, "May the LORD give you children by this woman to take the place of the one she prayed for and gave to the LORD." Then they would go home.
1SAM|2|21|And the LORD was gracious to Hannah; she conceived and gave birth to three sons and two daughters. Meanwhile, the boy Samuel grew up in the presence of the LORD.
1SAM|2|22|Now Eli, who was very old, heard about everything his sons were doing to all Israel and how they slept with the women who served at the entrance to the Tent of Meeting.
1SAM|2|23|So he said to them, "Why do you do such things? I hear from all the people about these wicked deeds of yours.
1SAM|2|24|No, my sons; it is not a good report that I hear spreading among the LORD's people.
1SAM|2|25|If a man sins against another man, God may mediate for him; but if a man sins against the LORD, who will intercede for him?" His sons, however, did not listen to their father's rebuke, for it was the LORD's will to put them to death.
1SAM|2|26|And the boy Samuel continued to grow in stature and in favor with the LORD and with men.
1SAM|2|27|Now a man of God came to Eli and said to him, "This is what the LORD says: 'Did I not clearly reveal myself to your father's house when they were in Egypt under Pharaoh?
1SAM|2|28|I chose your father out of all the tribes of Israel to be my priest, to go up to my altar, to burn incense, and to wear an ephod in my presence. I also gave your father's house all the offerings made with fire by the Israelites.
1SAM|2|29|Why do you scorn my sacrifice and offering that I prescribed for my dwelling? Why do you honor your sons more than me by fattening yourselves on the choice parts of every offering made by my people Israel?'
1SAM|2|30|"Therefore the LORD, the God of Israel, declares: 'I promised that your house and your father's house would minister before me forever.' But now the LORD declares: 'Far be it from me! Those who honor me I will honor, but those who despise me will be disdained.
1SAM|2|31|The time is coming when I will cut short your strength and the strength of your father's house, so that there will not be an old man in your family line
1SAM|2|32|and you will see distress in my dwelling. Although good will be done to Israel, in your family line there will never be an old man.
1SAM|2|33|Every one of you that I do not cut off from my altar will be spared only to blind your eyes with tears and to grieve your heart, and all your descendants will die in the prime of life.
1SAM|2|34|"'And what happens to your two sons, Hophni and Phinehas, will be a sign to you-they will both die on the same day.
1SAM|2|35|I will raise up for myself a faithful priest, who will do according to what is in my heart and mind. I will firmly establish his house, and he will minister before my anointed one always.
1SAM|2|36|Then everyone left in your family line will come and bow down before him for a piece of silver and a crust of bread and plead, "Appoint me to some priestly office so I can have food to eat."'"
1SAM|3|1|The boy Samuel ministered before the LORD under Eli. In those days the word of the LORD was rare; there were not many visions.
1SAM|3|2|One night Eli, whose eyes were becoming so weak that he could barely see, was lying down in his usual place.
1SAM|3|3|The lamp of God had not yet gone out, and Samuel was lying down in the temple of the LORD, where the ark of God was.
1SAM|3|4|Then the LORD called Samuel. Samuel answered, "Here I am."
1SAM|3|5|And he ran to Eli and said, "Here I am; you called me." But Eli said, "I did not call; go back and lie down." So he went and lay down.
1SAM|3|6|Again the LORD called, "Samuel!" And Samuel got up and went to Eli and said, "Here I am; you called me.My son," Eli said, "I did not call; go back and lie down."
1SAM|3|7|Now Samuel did not yet know the LORD: The word of the LORD had not yet been revealed to him.
1SAM|3|8|The LORD called Samuel a third time, and Samuel got up and went to Eli and said, "Here I am; you called me." Then Eli realized that the LORD was calling the boy.
1SAM|3|9|So Eli told Samuel, "Go and lie down, and if he calls you, say, 'Speak, LORD, for your servant is listening.'" So Samuel went and lay down in his place.
1SAM|3|10|The LORD came and stood there, calling as at the other times, "Samuel! Samuel!" Then Samuel said, "Speak, for your servant is listening."
1SAM|3|11|And the LORD said to Samuel: "See, I am about to do something in Israel that will make the ears of everyone who hears of it tingle.
1SAM|3|12|At that time I will carry out against Eli everything I spoke against his family-from beginning to end.
1SAM|3|13|For I told him that I would judge his family forever because of the sin he knew about; his sons made themselves contemptible, and he failed to restrain them.
1SAM|3|14|Therefore, I swore to the house of Eli, 'The guilt of Eli's house will never be atoned for by sacrifice or offering.'"
1SAM|3|15|Samuel lay down until morning and then opened the doors of the house of the LORD. He was afraid to tell Eli the vision,
1SAM|3|16|but Eli called him and said, "Samuel, my son." Samuel answered, "Here I am."
1SAM|3|17|"What was it he said to you?" Eli asked. "Do not hide it from me. May God deal with you, be it ever so severely, if you hide from me anything he told you."
1SAM|3|18|So Samuel told him everything, hiding nothing from him. Then Eli said, "He is the LORD; let him do what is good in his eyes."
1SAM|3|19|The LORD was with Samuel as he grew up, and he let none of his words fall to the ground.
1SAM|3|20|And all Israel from Dan to Beersheba recognized that Samuel was attested as a prophet of the LORD.
1SAM|3|21|The LORD continued to appear at Shiloh, and there he revealed himself to Samuel through his word.
1SAM|4|1|And Samuel's word came to all Israel. Now the Israelites went out to fight against the Philistines. The Israelites camped at Ebenezer, and the Philistines at Aphek.
1SAM|4|2|The Philistines deployed their forces to meet Israel, and as the battle spread, Israel was defeated by the Philistines, who killed about four thousand of them on the battlefield.
1SAM|4|3|When the soldiers returned to camp, the elders of Israel asked, "Why did the LORD bring defeat upon us today before the Philistines? Let us bring the ark of the LORD's covenant from Shiloh, so that it may go with us and save us from the hand of our enemies."
1SAM|4|4|So the people sent men to Shiloh, and they brought back the ark of the covenant of the LORD Almighty, who is enthroned between the cherubim. And Eli's two sons, Hophni and Phinehas, were there with the ark of the covenant of God.
1SAM|4|5|When the ark of the LORD's covenant came into the camp, all Israel raised such a great shout that the ground shook.
1SAM|4|6|Hearing the uproar, the Philistines asked, "What's all this shouting in the Hebrew camp?" When they learned that the ark of the LORD had come into the camp,
1SAM|4|7|the Philistines were afraid. "A god has come into the camp," they said. "We're in trouble! Nothing like this has happened before.
1SAM|4|8|Woe to us! Who will deliver us from the hand of these mighty gods? They are the gods who struck the Egyptians with all kinds of plagues in the desert.
1SAM|4|9|Be strong, Philistines! Be men, or you will be subject to the Hebrews, as they have been to you. Be men, and fight!"
1SAM|4|10|So the Philistines fought, and the Israelites were defeated and every man fled to his tent. The slaughter was very great; Israel lost thirty thousand foot soldiers.
1SAM|4|11|The ark of God was captured, and Eli's two sons, Hophni and Phinehas, died.
1SAM|4|12|That same day a Benjamite ran from the battle line and went to Shiloh, his clothes torn and dust on his head.
1SAM|4|13|When he arrived, there was Eli sitting on his chair by the side of the road, watching, because his heart feared for the ark of God. When the man entered the town and told what had happened, the whole town sent up a cry.
1SAM|4|14|Eli heard the outcry and asked, "What is the meaning of this uproar?" The man hurried over to Eli,
1SAM|4|15|who was ninety-eight years old and whose eyes were set so that he could not see.
1SAM|4|16|He told Eli, "I have just come from the battle line; I fled from it this very day." Eli asked, "What happened, my son?"
1SAM|4|17|The man who brought the news replied, "Israel fled before the Philistines, and the army has suffered heavy losses. Also your two sons, Hophni and Phinehas, are dead, and the ark of God has been captured."
1SAM|4|18|When he mentioned the ark of God, Eli fell backward off his chair by the side of the gate. His neck was broken and he died, for he was an old man and heavy. He had led Israel forty years.
1SAM|4|19|His daughter-in-law, the wife of Phinehas, was pregnant and near the time of delivery. When she heard the news that the ark of God had been captured and that her father-in-law and her husband were dead, she went into labor and gave birth, but was overcome by her labor pains.
1SAM|4|20|As she was dying, the women attending her said, "Don't despair; you have given birth to a son." But she did not respond or pay any attention.
1SAM|4|21|She named the boy Ichabod, saying, "The glory has departed from Israel"-because of the capture of the ark of God and the deaths of her father-in-law and her husband.
1SAM|4|22|She said, "The glory has departed from Israel, for the ark of God has been captured."
1SAM|5|1|After the Philistines had captured the ark of God, they took it from Ebenezer to Ashdod.
1SAM|5|2|Then they carried the ark into Dagon's temple and set it beside Dagon.
1SAM|5|3|When the people of Ashdod rose early the next day, there was Dagon, fallen on his face on the ground before the ark of the LORD! They took Dagon and put him back in his place.
1SAM|5|4|But the following morning when they rose, there was Dagon, fallen on his face on the ground before the ark of the LORD! His head and hands had been broken off and were lying on the threshold; only his body remained.
1SAM|5|5|That is why to this day neither the priests of Dagon nor any others who enter Dagon's temple at Ashdod step on the threshold.
1SAM|5|6|The LORD's hand was heavy upon the people of Ashdod and its vicinity; he brought devastation upon them and afflicted them with tumors.
1SAM|5|7|When the men of Ashdod saw what was happening, they said, "The ark of the god of Israel must not stay here with us, because his hand is heavy upon us and upon Dagon our god."
1SAM|5|8|So they called together all the rulers of the Philistines and asked them, "What shall we do with the ark of the god of Israel?" They answered, "Have the ark of the god of Israel moved to Gath." So they moved the ark of the God of Israel.
1SAM|5|9|But after they had moved it, the LORD's hand was against that city, throwing it into a great panic. He afflicted the people of the city, both young and old, with an outbreak of tumors.
1SAM|5|10|So they sent the ark of God to Ekron. As the ark of God was entering Ekron, the people of Ekron cried out, "They have brought the ark of the god of Israel around to us to kill us and our people."
1SAM|5|11|So they called together all the rulers of the Philistines and said, "Send the ark of the god of Israel away; let it go back to its own place, or it will kill us and our people." For death had filled the city with panic; God's hand was very heavy upon it.
1SAM|5|12|Those who did not die were afflicted with tumors, and the outcry of the city went up to heaven.
1SAM|6|1|When the ark of the LORD had been in Philistine territory seven months,
1SAM|6|2|the Philistines called for the priests and the diviners and said, "What shall we do with the ark of the LORD? Tell us how we should send it back to its place."
1SAM|6|3|They answered, "If you return the ark of the god of Israel, do not send it away empty, but by all means send a guilt offering to him. Then you will be healed, and you will know why his hand has not been lifted from you."
1SAM|6|4|The Philistines asked, "What guilt offering should we send to him?" They replied, "Five gold tumors and five gold rats, according to the number of the Philistine rulers, because the same plague has struck both you and your rulers.
1SAM|6|5|Make models of the tumors and of the rats that are destroying the country, and pay honor to Israel's god. Perhaps he will lift his hand from you and your gods and your land.
1SAM|6|6|Why do you harden your hearts as the Egyptians and Pharaoh did? When he treated them harshly, did they not send the Israelites out so they could go on their way?
1SAM|6|7|"Now then, get a new cart ready, with two cows that have calved and have never been yoked. Hitch the cows to the cart, but take their calves away and pen them up.
1SAM|6|8|Take the ark of the LORD and put it on the cart, and in a chest beside it put the gold objects you are sending back to him as a guilt offering. Send it on its way,
1SAM|6|9|but keep watching it. If it goes up to its own territory, toward Beth Shemesh, then the LORD has brought this great disaster on us. But if it does not, then we will know that it was not his hand that struck us and that it happened to us by chance."
1SAM|6|10|So they did this. They took two such cows and hitched them to the cart and penned up their calves.
1SAM|6|11|They placed the ark of the LORD on the cart and along with it the chest containing the gold rats and the models of the tumors.
1SAM|6|12|Then the cows went straight up toward Beth Shemesh, keeping on the road and lowing all the way; they did not turn to the right or to the left. The rulers of the Philistines followed them as far as the border of Beth Shemesh.
1SAM|6|13|Now the people of Beth Shemesh were harvesting their wheat in the valley, and when they looked up and saw the ark, they rejoiced at the sight.
1SAM|6|14|The cart came to the field of Joshua of Beth Shemesh, and there it stopped beside a large rock. The people chopped up the wood of the cart and sacrificed the cows as a burnt offering to the LORD.
1SAM|6|15|The Levites took down the ark of the LORD, together with the chest containing the gold objects, and placed them on the large rock. On that day the people of Beth Shemesh offered burnt offerings and made sacrifices to the LORD.
1SAM|6|16|The five rulers of the Philistines saw all this and then returned that same day to Ekron.
1SAM|6|17|These are the gold tumors the Philistines sent as a guilt offering to the LORD -one each for Ashdod, Gaza, Ashkelon, Gath and Ekron.
1SAM|6|18|And the number of the gold rats was according to the number of Philistine towns belonging to the five rulers-the fortified towns with their country villages. The large rock, on which they set the ark of the LORD, is a witness to this day in the field of Joshua of Beth Shemesh.
1SAM|6|19|But God struck down some of the men of Beth Shemesh, putting seventy of them to death because they had looked into the ark of the LORD. The people mourned because of the heavy blow the LORD had dealt them,
1SAM|6|20|and the men of Beth Shemesh asked, "Who can stand in the presence of the LORD, this holy God? To whom will the ark go up from here?"
1SAM|6|21|Then they sent messengers to the people of Kiriath Jearim, saying, "The Philistines have returned the ark of the LORD. Come down and take it up to your place."
1SAM|7|1|So the men of Kiriath Jearim came and took up the ark of the LORD. They took it to Abinadab's house on the hill and consecrated Eleazar his son to guard the ark of the LORD.
1SAM|7|2|It was a long time, twenty years in all, that the ark remained at Kiriath Jearim, and all the people of Israel mourned and sought after the LORD.
1SAM|7|3|And Samuel said to the whole house of Israel, "If you are returning to the LORD with all your hearts, then rid yourselves of the foreign gods and the Ashtoreths and commit yourselves to the LORD and serve him only, and he will deliver you out of the hand of the Philistines."
1SAM|7|4|So the Israelites put away their Baals and Ashtoreths, and served the LORD only.
1SAM|7|5|Then Samuel said, "Assemble all Israel at Mizpah and I will intercede with the LORD for you."
1SAM|7|6|When they had assembled at Mizpah, they drew water and poured it out before the LORD. On that day they fasted and there they confessed, "We have sinned against the LORD." And Samuel was leader of Israel at Mizpah.
1SAM|7|7|When the Philistines heard that Israel had assembled at Mizpah, the rulers of the Philistines came up to attack them. And when the Israelites heard of it, they were afraid because of the Philistines.
1SAM|7|8|They said to Samuel, "Do not stop crying out to the LORD our God for us, that he may rescue us from the hand of the Philistines."
1SAM|7|9|Then Samuel took a suckling lamb and offered it up as a whole burnt offering to the LORD. He cried out to the LORD on Israel's behalf, and the LORD answered him.
1SAM|7|10|While Samuel was sacrificing the burnt offering, the Philistines drew near to engage Israel in battle. But that day the LORD thundered with loud thunder against the Philistines and threw them into such a panic that they were routed before the Israelites.
1SAM|7|11|The men of Israel rushed out of Mizpah and pursued the Philistines, slaughtering them along the way to a point below Beth Car.
1SAM|7|12|Then Samuel took a stone and set it up between Mizpah and Shen. He named it Ebenezer, saying, "Thus far has the LORD helped us."
1SAM|7|13|So the Philistines were subdued and did not invade Israelite territory again. Throughout Samuel's lifetime, the hand of the LORD was against the Philistines.
1SAM|7|14|The towns from Ekron to Gath that the Philistines had captured from Israel were restored to her, and Israel delivered the neighboring territory from the power of the Philistines. And there was peace between Israel and the Amorites.
1SAM|7|15|Samuel continued as judge over Israel all the days of his life.
1SAM|7|16|From year to year he went on a circuit from Bethel to Gilgal to Mizpah, judging Israel in all those places.
1SAM|7|17|But he always went back to Ramah, where his home was, and there he also judged Israel. And he built an altar there to the LORD.
1SAM|8|1|When Samuel grew old, he appointed his sons as judges for Israel.
1SAM|8|2|The name of his firstborn was Joel and the name of his second was Abijah, and they served at Beersheba.
1SAM|8|3|But his sons did not walk in his ways. They turned aside after dishonest gain and accepted bribes and perverted justice.
1SAM|8|4|So all the elders of Israel gathered together and came to Samuel at Ramah.
1SAM|8|5|They said to him, "You are old, and your sons do not walk in your ways; now appoint a king to lead us, such as all the other nations have."
1SAM|8|6|But when they said, "Give us a king to lead us," this displeased Samuel; so he prayed to the LORD.
1SAM|8|7|And the LORD told him: "Listen to all that the people are saying to you; it is not you they have rejected, but they have rejected me as their king.
1SAM|8|8|As they have done from the day I brought them up out of Egypt until this day, forsaking me and serving other gods, so they are doing to you.
1SAM|8|9|Now listen to them; but warn them solemnly and let them know what the king who will reign over them will do."
1SAM|8|10|Samuel told all the words of the LORD to the people who were asking him for a king.
1SAM|8|11|He said, "This is what the king who will reign over you will do: He will take your sons and make them serve with his chariots and horses, and they will run in front of his chariots.
1SAM|8|12|Some he will assign to be commanders of thousands and commanders of fifties, and others to plow his ground and reap his harvest, and still others to make weapons of war and equipment for his chariots.
1SAM|8|13|He will take your daughters to be perfumers and cooks and bakers.
1SAM|8|14|He will take the best of your fields and vineyards and olive groves and give them to his attendants.
1SAM|8|15|He will take a tenth of your grain and of your vintage and give it to his officials and attendants.
1SAM|8|16|Your menservants and maidservants and the best of your cattle and donkeys he will take for his own use.
1SAM|8|17|He will take a tenth of your flocks, and you yourselves will become his slaves.
1SAM|8|18|When that day comes, you will cry out for relief from the king you have chosen, and the LORD will not answer you in that day."
1SAM|8|19|But the people refused to listen to Samuel. "No!" they said. "We want a king over us.
1SAM|8|20|Then we will be like all the other nations, with a king to lead us and to go out before us and fight our battles."
1SAM|8|21|When Samuel heard all that the people said, he repeated it before the LORD.
1SAM|8|22|The LORD answered, "Listen to them and give them a king." Then Samuel said to the men of Israel, "Everyone go back to his town."
1SAM|9|1|There was a Benjamite, a man of standing, whose name was Kish son of Abiel, the son of Zeror, the son of Becorath, the son of Aphiah of Benjamin.
1SAM|9|2|He had a son named Saul, an impressive young man without equal among the Israelites-a head taller than any of the others.
1SAM|9|3|Now the donkeys belonging to Saul's father Kish were lost, and Kish said to his son Saul, "Take one of the servants with you and go and look for the donkeys."
1SAM|9|4|So he passed through the hill country of Ephraim and through the area around Shalisha, but they did not find them. They went on into the district of Shaalim, but the donkeys were not there. Then he passed through the territory of Benjamin, but they did not find them.
1SAM|9|5|When they reached the district of Zuph, Saul said to the servant who was with him, "Come, let's go back, or my father will stop thinking about the donkeys and start worrying about us."
1SAM|9|6|But the servant replied, "Look, in this town there is a man of God; he is highly respected, and everything he says comes true. Let's go there now. Perhaps he will tell us what way to take."
1SAM|9|7|Saul said to his servant, "If we go, what can we give the man? The food in our sacks is gone. We have no gift to take to the man of God. What do we have?"
1SAM|9|8|The servant answered him again. "Look," he said, "I have a quarter of a shekel of silver. I will give it to the man of God so that he will tell us what way to take."
1SAM|9|9|(Formerly in Israel, if a man went to inquire of God, he would say, "Come, let us go to the seer," because the prophet of today used to be called a seer.)
1SAM|9|10|"Good," Saul said to his servant. "Come, let's go." So they set out for the town where the man of God was.
1SAM|9|11|As they were going up the hill to the town, they met some girls coming out to draw water, and they asked them, "Is the seer here?"
1SAM|9|12|"He is," they answered. "He's ahead of you. Hurry now; he has just come to our town today, for the people have a sacrifice at the high place.
1SAM|9|13|As soon as you enter the town, you will find him before he goes up to the high place to eat. The people will not begin eating until he comes, because he must bless the sacrifice; afterward, those who are invited will eat. Go up now; you should find him about this time."
1SAM|9|14|They went up to the town, and as they were entering it, there was Samuel, coming toward them on his way up to the high place.
1SAM|9|15|Now the day before Saul came, the LORD had revealed this to Samuel:
1SAM|9|16|"About this time tomorrow I will send you a man from the land of Benjamin. Anoint him leader over my people Israel; he will deliver my people from the hand of the Philistines. I have looked upon my people, for their cry has reached me."
1SAM|9|17|When Samuel caught sight of Saul, the LORD said to him, "This is the man I spoke to you about; he will govern my people."
1SAM|9|18|Saul approached Samuel in the gateway and asked, "Would you please tell me where the seer's house is?"
1SAM|9|19|"I am the seer," Samuel replied. "Go up ahead of me to the high place, for today you are to eat with me, and in the morning I will let you go and will tell you all that is in your heart.
1SAM|9|20|As for the donkeys you lost three days ago, do not worry about them; they have been found. And to whom is all the desire of Israel turned, if not to you and all your father's family?"
1SAM|9|21|Saul answered, "But am I not a Benjamite, from the smallest tribe of Israel, and is not my clan the least of all the clans of the tribe of Benjamin? Why do you say such a thing to me?"
1SAM|9|22|Then Samuel brought Saul and his servant into the hall and seated them at the head of those who were invited-about thirty in number.
1SAM|9|23|Samuel said to the cook, "Bring the piece of meat I gave you, the one I told you to lay aside."
1SAM|9|24|So the cook took up the leg with what was on it and set it in front of Saul. Samuel said, "Here is what has been kept for you. Eat, because it was set aside for you for this occasion, from the time I said, 'I have invited guests.'" And Saul dined with Samuel that day.
1SAM|9|25|After they came down from the high place to the town, Samuel talked with Saul on the roof of his house.
1SAM|9|26|They rose about daybreak and Samuel called to Saul on the roof, "Get ready, and I will send you on your way." When Saul got ready, he and Samuel went outside together.
1SAM|9|27|As they were going down to the edge of the town, Samuel said to Saul, "Tell the servant to go on ahead of us"-and the servant did so-"but you stay here awhile, so that I may give you a message from God."
1SAM|10|1|Then Samuel took a flask of oil and poured it on Saul's head and kissed him, saying, "Has not the LORD anointed you leader over his inheritance?
1SAM|10|2|When you leave me today, you will meet two men near Rachel's tomb, at Zelzah on the border of Benjamin. They will say to you, 'The donkeys you set out to look for have been found. And now your father has stopped thinking about them and is worried about you. He is asking, "What shall I do about my son?"'
1SAM|10|3|"Then you will go on from there until you reach the great tree of Tabor. Three men going up to God at Bethel will meet you there. One will be carrying three young goats, another three loaves of bread, and another a skin of wine.
1SAM|10|4|They will greet you and offer you two loaves of bread, which you will accept from them.
1SAM|10|5|"After that you will go to Gibeah of God, where there is a Philistine outpost. As you approach the town, you will meet a procession of prophets coming down from the high place with lyres, tambourines, flutes and harps being played before them, and they will be prophesying.
1SAM|10|6|The Spirit of the LORD will come upon you in power, and you will prophesy with them; and you will be changed into a different person.
1SAM|10|7|Once these signs are fulfilled, do whatever your hand finds to do, for God is with you.
1SAM|10|8|"Go down ahead of me to Gilgal. I will surely come down to you to sacrifice burnt offerings and fellowship offerings, but you must wait seven days until I come to you and tell you what you are to do."
1SAM|10|9|As Saul turned to leave Samuel, God changed Saul's heart, and all these signs were fulfilled that day.
1SAM|10|10|When they arrived at Gibeah, a procession of prophets met him; the Spirit of God came upon him in power, and he joined in their prophesying.
1SAM|10|11|When all those who had formerly known him saw him prophesying with the prophets, they asked each other, "What is this that has happened to the son of Kish? Is Saul also among the prophets?"
1SAM|10|12|A man who lived there answered, "And who is their father?" So it became a saying: "Is Saul also among the prophets?"
1SAM|10|13|After Saul stopped prophesying, he went to the high place.
1SAM|10|14|Now Saul's uncle asked him and his servant, "Where have you been?Looking for the donkeys," he said. "But when we saw they were not to be found, we went to Samuel."
1SAM|10|15|Saul's uncle said, "Tell me what Samuel said to you."
1SAM|10|16|Saul replied, "He assured us that the donkeys had been found." But he did not tell his uncle what Samuel had said about the kingship.
1SAM|10|17|Samuel summoned the people of Israel to the LORD at Mizpah
1SAM|10|18|and said to them, "This is what the LORD, the God of Israel, says: 'I brought Israel up out of Egypt, and I delivered you from the power of Egypt and all the kingdoms that oppressed you.'
1SAM|10|19|But you have now rejected your God, who saves you out of all your calamities and distresses. And you have said, 'No, set a king over us.' So now present yourselves before the LORD by your tribes and clans."
1SAM|10|20|When Samuel brought all the tribes of Israel near, the tribe of Benjamin was chosen.
1SAM|10|21|Then he brought forward the tribe of Benjamin, clan by clan, and Matri's clan was chosen. Finally Saul son of Kish was chosen. But when they looked for him, he was not to be found.
1SAM|10|22|So they inquired further of the LORD, "Has the man come here yet?" And the LORD said, "Yes, he has hidden himself among the baggage."
1SAM|10|23|They ran and brought him out, and as he stood among the people he was a head taller than any of the others.
1SAM|10|24|Samuel said to all the people, "Do you see the man the LORD has chosen? There is no one like him among all the people." Then the people shouted, "Long live the king!"
1SAM|10|25|Samuel explained to the people the regulations of the kingship. He wrote them down on a scroll and deposited it before the LORD. Then Samuel dismissed the people, each to his own home.
1SAM|10|26|Saul also went to his home in Gibeah, accompanied by valiant men whose hearts God had touched.
1SAM|10|27|But some troublemakers said, "How can this fellow save us?" They despised him and brought him no gifts. But Saul kept silent.
1SAM|11|1|Nahash the Ammonite went up and besieged Jabesh Gilead. And all the men of Jabesh said to him, "Make a treaty with us, and we will be subject to you."
1SAM|11|2|But Nahash the Ammonite replied, "I will make a treaty with you only on the condition that I gouge out the right eye of every one of you and so bring disgrace on all Israel."
1SAM|11|3|The elders of Jabesh said to him, "Give us seven days so we can send messengers throughout Israel; if no one comes to rescue us, we will surrender to you."
1SAM|11|4|When the messengers came to Gibeah of Saul and reported these terms to the people, they all wept aloud.
1SAM|11|5|Just then Saul was returning from the fields, behind his oxen, and he asked, "What is wrong with the people? Why are they weeping?" Then they repeated to him what the men of Jabesh had said.
1SAM|11|6|When Saul heard their words, the Spirit of God came upon him in power, and he burned with anger.
1SAM|11|7|He took a pair of oxen, cut them into pieces, and sent the pieces by messengers throughout Israel, proclaiming, "This is what will be done to the oxen of anyone who does not follow Saul and Samuel." Then the terror of the LORD fell on the people, and they turned out as one man.
1SAM|11|8|When Saul mustered them at Bezek, the men of Israel numbered three hundred thousand and the men of Judah thirty thousand.
1SAM|11|9|They told the messengers who had come, "Say to the men of Jabesh Gilead, 'By the time the sun is hot tomorrow, you will be delivered.'" When the messengers went and reported this to the men of Jabesh, they were elated.
1SAM|11|10|They said to the Ammonites, "Tomorrow we will surrender to you, and you can do to us whatever seems good to you."
1SAM|11|11|The next day Saul separated his men into three divisions; during the last watch of the night they broke into the camp of the Ammonites and slaughtered them until the heat of the day. Those who survived were scattered, so that no two of them were left together.
1SAM|11|12|The people then said to Samuel, "Who was it that asked, 'Shall Saul reign over us?' Bring these men to us and we will put them to death."
1SAM|11|13|But Saul said, "No one shall be put to death today, for this day the LORD has rescued Israel."
1SAM|11|14|Then Samuel said to the people, "Come, let us go to Gilgal and there reaffirm the kingship."
1SAM|11|15|So all the people went to Gilgal and confirmed Saul as king in the presence of the LORD. There they sacrificed fellowship offerings before the LORD, and Saul and all the Israelites held a great celebration.
1SAM|12|1|Samuel said to all Israel, "I have listened to everything you said to me and have set a king over you.
1SAM|12|2|Now you have a king as your leader. As for me, I am old and gray, and my sons are here with you. I have been your leader from my youth until this day.
1SAM|12|3|Here I stand. Testify against me in the presence of the LORD and his anointed. Whose ox have I taken? Whose donkey have I taken? Whom have I cheated? Whom have I oppressed? From whose hand have I accepted a bribe to make me shut my eyes? If I have done any of these, I will make it right."
1SAM|12|4|"You have not cheated or oppressed us," they replied. "You have not taken anything from anyone's hand."
1SAM|12|5|Samuel said to them, "The LORD is witness against you, and also his anointed is witness this day, that you have not found anything in my hand.He is witness," they said.
1SAM|12|6|Then Samuel said to the people, "It is the LORD who appointed Moses and Aaron and brought your forefathers up out of Egypt.
1SAM|12|7|Now then, stand here, because I am going to confront you with evidence before the LORD as to all the righteous acts performed by the LORD for you and your fathers.
1SAM|12|8|"After Jacob entered Egypt, they cried to the LORD for help, and the LORD sent Moses and Aaron, who brought your forefathers out of Egypt and settled them in this place.
1SAM|12|9|"But they forgot the LORD their God; so he sold them into the hand of Sisera, the commander of the army of Hazor, and into the hands of the Philistines and the king of Moab, who fought against them.
1SAM|12|10|They cried out to the LORD and said, 'We have sinned; we have forsaken the LORD and served the Baals and the Ashtoreths. But now deliver us from the hands of our enemies, and we will serve you.'
1SAM|12|11|Then the LORD sent Jerub-Baal, Barak, Jephthah and Samuel, and he delivered you from the hands of your enemies on every side, so that you lived securely.
1SAM|12|12|"But when you saw that Nahash king of the Ammonites was moving against you, you said to me, 'No, we want a king to rule over us'-even though the LORD your God was your king.
1SAM|12|13|Now here is the king you have chosen, the one you asked for; see, the LORD has set a king over you.
1SAM|12|14|If you fear the LORD and serve and obey him and do not rebel against his commands, and if both you and the king who reigns over you follow the LORD your God-good!
1SAM|12|15|But if you do not obey the LORD, and if you rebel against his commands, his hand will be against you, as it was against your fathers.
1SAM|12|16|"Now then, stand still and see this great thing the LORD is about to do before your eyes!
1SAM|12|17|Is it not wheat harvest now? I will call upon the LORD to send thunder and rain. And you will realize what an evil thing you did in the eyes of the LORD when you asked for a king."
1SAM|12|18|Then Samuel called upon the LORD, and that same day the LORD sent thunder and rain. So all the people stood in awe of the LORD and of Samuel.
1SAM|12|19|The people all said to Samuel, "Pray to the LORD your God for your servants so that we will not die, for we have added to all our other sins the evil of asking for a king."
1SAM|12|20|"Do not be afraid," Samuel replied. "You have done all this evil; yet do not turn away from the LORD, but serve the LORD with all your heart.
1SAM|12|21|Do not turn away after useless idols. They can do you no good, nor can they rescue you, because they are useless.
1SAM|12|22|For the sake of his great name the LORD will not reject his people, because the LORD was pleased to make you his own.
1SAM|12|23|As for me, far be it from me that I should sin against the LORD by failing to pray for you. And I will teach you the way that is good and right.
1SAM|12|24|But be sure to fear the LORD and serve him faithfully with all your heart; consider what great things he has done for you.
1SAM|12|25|Yet if you persist in doing evil, both you and your king will be swept away."
1SAM|13|1|Saul was thirty years old when he became king, and he reigned over Israel forty- two years.
1SAM|13|2|Saul chose three thousand men from Israel; two thousand were with him at Micmash and in the hill country of Bethel, and a thousand were with Jonathan at Gibeah in Benjamin. The rest of the men he sent back to their homes.
1SAM|13|3|Jonathan attacked the Philistine outpost at Geba, and the Philistines heard about it. Then Saul had the trumpet blown throughout the land and said, "Let the Hebrews hear!"
1SAM|13|4|So all Israel heard the news: "Saul has attacked the Philistine outpost, and now Israel has become a stench to the Philistines." And the people were summoned to join Saul at Gilgal.
1SAM|13|5|The Philistines assembled to fight Israel, with three thousand chariots, six thousand charioteers, and soldiers as numerous as the sand on the seashore. They went up and camped at Micmash, east of Beth Aven.
1SAM|13|6|When the men of Israel saw that their situation was critical and that their army was hard pressed, they hid in caves and thickets, among the rocks, and in pits and cisterns.
1SAM|13|7|Some Hebrews even crossed the Jordan to the land of Gad and Gilead. Saul remained at Gilgal, and all the troops with him were quaking with fear.
1SAM|13|8|He waited seven days, the time set by Samuel; but Samuel did not come to Gilgal, and Saul's men began to scatter.
1SAM|13|9|So he said, "Bring me the burnt offering and the fellowship offerings. "And Saul offered up the burnt offering.
1SAM|13|10|Just as he finished making the offering, Samuel arrived, and Saul went out to greet him.
1SAM|13|11|"What have you done?" asked Samuel. Saul replied, "When I saw that the men were scattering, and that you did not come at the set time, and that the Philistines were assembling at Micmash,
1SAM|13|12|I thought, 'Now the Philistines will come down against me at Gilgal, and I have not sought the LORD's favor.' So I felt compelled to offer the burnt offering."
1SAM|13|13|"You acted foolishly," Samuel said. "You have not kept the command the LORD your God gave you; if you had, he would have established your kingdom over Israel for all time.
1SAM|13|14|But now your kingdom will not endure; the LORD has sought out a man after his own heart and appointed him leader of his people, because you have not kept the LORD's command."
1SAM|13|15|Then Samuel left Gilgal and went up to Gibeah in Benjamin, and Saul counted the men who were with him. They numbered about six hundred.
1SAM|13|16|Saul and his son Jonathan and the men with them were staying in Gibeah in Benjamin, while the Philistines camped at Micmash.
1SAM|13|17|Raiding parties went out from the Philistine camp in three detachments. One turned toward Ophrah in the vicinity of Shual,
1SAM|13|18|another toward Beth Horon, and the third toward the borderland overlooking the Valley of Zeboim facing the desert.
1SAM|13|19|Not a blacksmith could be found in the whole land of Israel, because the Philistines had said, "Otherwise the Hebrews will make swords or spears!"
1SAM|13|20|So all Israel went down to the Philistines to have their plowshares, mattocks, axes and sickles sharpened.
1SAM|13|21|The price was two thirds of a shekel for sharpening plowshares and mattocks, and a third of a shekel for sharpening forks and axes and for repointing goads.
1SAM|13|22|So on the day of the battle not a soldier with Saul and Jonathan had a sword or spear in his hand; only Saul and his son Jonathan had them.
1SAM|13|23|Now a detachment of Philistines had gone out to the pass at Micmash.
1SAM|14|1|One day Jonathan son of Saul said to the young man bearing his armor, "Come, let's go over to the Philistine outpost on the other side." But he did not tell his father.
1SAM|14|2|Saul was staying on the outskirts of Gibeah under a pomegranate tree in Migron. With him were about six hundred men,
1SAM|14|3|among whom was Ahijah, who was wearing an ephod. He was a son of Ichabod's brother Ahitub son of Phinehas, the son of Eli, the LORD's priest in Shiloh. No one was aware that Jonathan had left.
1SAM|14|4|On each side of the pass that Jonathan intended to cross to reach the Philistine outpost was a cliff; one was called Bozez, and the other Seneh.
1SAM|14|5|One cliff stood to the north toward Micmash, the other to the south toward Geba.
1SAM|14|6|Jonathan said to his young armor-bearer, "Come, let's go over to the outpost of those uncircumcised fellows. Perhaps the LORD will act in our behalf. Nothing can hinder the LORD from saving, whether by many or by few."
1SAM|14|7|"Do all that you have in mind," his armor-bearer said. "Go ahead; I am with you heart and soul."
1SAM|14|8|Jonathan said, "Come, then; we will cross over toward the men and let them see us.
1SAM|14|9|If they say to us, 'Wait there until we come to you,' we will stay where we are and not go up to them.
1SAM|14|10|But if they say, 'Come up to us,' we will climb up, because that will be our sign that the LORD has given them into our hands."
1SAM|14|11|So both of them showed themselves to the Philistine outpost. "Look!" said the Philistines. "The Hebrews are crawling out of the holes they were hiding in."
1SAM|14|12|The men of the outpost shouted to Jonathan and his armor-bearer, "Come up to us and we'll teach you a lesson." So Jonathan said to his armor-bearer, "Climb up after me; the LORD has given them into the hand of Israel."
1SAM|14|13|Jonathan climbed up, using his hands and feet, with his armor-bearer right behind him. The Philistines fell before Jonathan, and his armor-bearer followed and killed behind him.
1SAM|14|14|In that first attack Jonathan and his armor-bearer killed some twenty men in an area of about half an acre.
1SAM|14|15|Then panic struck the whole army-those in the camp and field, and those in the outposts and raiding parties-and the ground shook. It was a panic sent by God.
1SAM|14|16|Saul's lookouts at Gibeah in Benjamin saw the army melting away in all directions.
1SAM|14|17|Then Saul said to the men who were with him, "Muster the forces and see who has left us." When they did, it was Jonathan and his armor-bearer who were not there.
1SAM|14|18|Saul said to Ahijah, "Bring the ark of God." (At that time it was with the Israelites.)
1SAM|14|19|While Saul was talking to the priest, the tumult in the Philistine camp increased more and more. So Saul said to the priest, "Withdraw your hand."
1SAM|14|20|Then Saul and all his men assembled and went to the battle. They found the Philistines in total confusion, striking each other with their swords.
1SAM|14|21|Those Hebrews who had previously been with the Philistines and had gone up with them to their camp went over to the Israelites who were with Saul and Jonathan.
1SAM|14|22|When all the Israelites who had hidden in the hill country of Ephraim heard that the Philistines were on the run, they joined the battle in hot pursuit.
1SAM|14|23|So the LORD rescued Israel that day, and the battle moved on beyond Beth Aven.
1SAM|14|24|Now the men of Israel were in distress that day, because Saul had bound the people under an oath, saying, "Cursed be any man who eats food before evening comes, before I have avenged myself on my enemies!" So none of the troops tasted food.
1SAM|14|25|The entire army entered the woods, and there was honey on the ground.
1SAM|14|26|When they went into the woods, they saw the honey oozing out, yet no one put his hand to his mouth, because they feared the oath.
1SAM|14|27|But Jonathan had not heard that his father had bound the people with the oath, so he reached out the end of the staff that was in his hand and dipped it into the honeycomb. He raised his hand to his mouth, and his eyes brightened.
1SAM|14|28|Then one of the soldiers told him, "Your father bound the army under a strict oath, saying, 'Cursed be any man who eats food today!' That is why the men are faint."
1SAM|14|29|Jonathan said, "My father has made trouble for the country. See how my eyes brightened when I tasted a little of this honey.
1SAM|14|30|How much better it would have been if the men had eaten today some of the plunder they took from their enemies. Would not the slaughter of the Philistines have been even greater?"
1SAM|14|31|That day, after the Israelites had struck down the Philistines from Micmash to Aijalon, they were exhausted.
1SAM|14|32|They pounced on the plunder and, taking sheep, cattle and calves, they butchered them on the ground and ate them, together with the blood.
1SAM|14|33|Then someone said to Saul, "Look, the men are sinning against the LORD by eating meat that has blood in it.You have broken faith," he said. "Roll a large stone over here at once."
1SAM|14|34|Then he said, "Go out among the men and tell them, 'Each of you bring me your cattle and sheep, and slaughter them here and eat them. Do not sin against the LORD by eating meat with blood still in it.'" So everyone brought his ox that night and slaughtered it there.
1SAM|14|35|Then Saul built an altar to the LORD; it was the first time he had done this.
1SAM|14|36|Saul said, "Let us go down after the Philistines by night and plunder them till dawn, and let us not leave one of them alive.Do whatever seems best to you," they replied. But the priest said, "Let us inquire of God here."
1SAM|14|37|So Saul asked God, "Shall I go down after the Philistines? Will you give them into Israel's hand?" But God did not answer him that day.
1SAM|14|38|Saul therefore said, "Come here, all you who are leaders of the army, and let us find out what sin has been committed today.
1SAM|14|39|As surely as the LORD who rescues Israel lives, even if it lies with my son Jonathan, he must die." But not one of the men said a word.
1SAM|14|40|Saul then said to all the Israelites, "You stand over there; I and Jonathan my son will stand over here.Do what seems best to you," the men replied.
1SAM|14|41|Then Saul prayed to the LORD, the God of Israel, "Give me the right answer." And Jonathan and Saul were taken by lot, and the men were cleared.
1SAM|14|42|Saul said, "Cast the lot between me and Jonathan my son." And Jonathan was taken.
1SAM|14|43|Then Saul said to Jonathan, "Tell me what you have done." So Jonathan told him, "I merely tasted a little honey with the end of my staff. And now must I die?"
1SAM|14|44|Saul said, "May God deal with me, be it ever so severely, if you do not die, Jonathan."
1SAM|14|45|But the men said to Saul, "Should Jonathan die-he who has brought about this great deliverance in Israel? Never! As surely as the LORD lives, not a hair of his head will fall to the ground, for he did this today with God's help." So the men rescued Jonathan, and he was not put to death.
1SAM|14|46|Then Saul stopped pursuing the Philistines, and they withdrew to their own land.
1SAM|14|47|After Saul had assumed rule over Israel, he fought against their enemies on every side: Moab, the Ammonites, Edom, the kings of Zobah, and the Philistines. Wherever he turned, he inflicted punishment on them.
1SAM|14|48|He fought valiantly and defeated the Amalekites, delivering Israel from the hands of those who had plundered them.
1SAM|14|49|Saul's sons were Jonathan, Ishvi and Malki-Shua. The name of his older daughter was Merab, and that of the younger was Michal.
1SAM|14|50|His wife's name was Ahinoam daughter of Ahimaaz. The name of the commander of Saul's army was Abner son of Ner, and Ner was Saul's uncle.
1SAM|14|51|Saul's father Kish and Abner's father Ner were sons of Abiel.
1SAM|14|52|All the days of Saul there was bitter war with the Philistines, and whenever Saul saw a mighty or brave man, he took him into his service.
1SAM|15|1|Samuel said to Saul, "I am the one the LORD sent to anoint you king over his people Israel; so listen now to the message from the LORD.
1SAM|15|2|This is what the LORD Almighty says: 'I will punish the Amalekites for what they did to Israel when they waylaid them as they came up from Egypt.
1SAM|15|3|Now go, attack the Amalekites and totally destroy everything that belongs to them. Do not spare them; put to death men and women, children and infants, cattle and sheep, camels and donkeys.'"
1SAM|15|4|So Saul summoned the men and mustered them at Telaim-two hundred thousand foot soldiers and ten thousand men from Judah.
1SAM|15|5|Saul went to the city of Amalek and set an ambush in the ravine.
1SAM|15|6|Then he said to the Kenites, "Go away, leave the Amalekites so that I do not destroy you along with them; for you showed kindness to all the Israelites when they came up out of Egypt." So the Kenites moved away from the Amalekites.
1SAM|15|7|Then Saul attacked the Amalekites all the way from Havilah to Shur, to the east of Egypt.
1SAM|15|8|He took Agag king of the Amalekites alive, and all his people he totally destroyed with the sword.
1SAM|15|9|But Saul and the army spared Agag and the best of the sheep and cattle, the fat calves and lambs-everything that was good. These they were unwilling to destroy completely, but everything that was despised and weak they totally destroyed.
1SAM|15|10|Then the word of the LORD came to Samuel:
1SAM|15|11|"I am grieved that I have made Saul king, because he has turned away from me and has not carried out my instructions." Samuel was troubled, and he cried out to the LORD all that night.
1SAM|15|12|Early in the morning Samuel got up and went to meet Saul, but he was told, "Saul has gone to Carmel. There he has set up a monument in his own honor and has turned and gone on down to Gilgal."
1SAM|15|13|When Samuel reached him, Saul said, "The LORD bless you! I have carried out the LORD's instructions."
1SAM|15|14|But Samuel said, "What then is this bleating of sheep in my ears? What is this lowing of cattle that I hear?"
1SAM|15|15|Saul answered, "The soldiers brought them from the Amalekites; they spared the best of the sheep and cattle to sacrifice to the LORD your God, but we totally destroyed the rest."
1SAM|15|16|"Stop!" Samuel said to Saul. "Let me tell you what the LORD said to me last night.Tell me," Saul replied.
1SAM|15|17|Samuel said, "Although you were once small in your own eyes, did you not become the head of the tribes of Israel? The LORD anointed you king over Israel.
1SAM|15|18|And he sent you on a mission, saying, 'Go and completely destroy those wicked people, the Amalekites; make war on them until you have wiped them out.'
1SAM|15|19|Why did you not obey the LORD? Why did you pounce on the plunder and do evil in the eyes of the LORD?"
1SAM|15|20|"But I did obey the LORD," Saul said. "I went on the mission the LORD assigned me. I completely destroyed the Amalekites and brought back Agag their king.
1SAM|15|21|The soldiers took sheep and cattle from the plunder, the best of what was devoted to God, in order to sacrifice them to the LORD your God at Gilgal."
1SAM|15|22|But Samuel replied: "Does the LORD delight in burnt offerings and sacrifices as much as in obeying the voice of the LORD? To obey is better than sacrifice, and to heed is better than the fat of rams.
1SAM|15|23|For rebellion is like the sin of divination, and arrogance like the evil of idolatry. Because you have rejected the word of the LORD, he has rejected you as king."
1SAM|15|24|Then Saul said to Samuel, "I have sinned. I violated the LORD's command and your instructions. I was afraid of the people and so I gave in to them.
1SAM|15|25|Now I beg you, forgive my sin and come back with me, so that I may worship the LORD."
1SAM|15|26|But Samuel said to him, "I will not go back with you. You have rejected the word of the LORD, and the LORD has rejected you as king over Israel!"
1SAM|15|27|As Samuel turned to leave, Saul caught hold of the hem of his robe, and it tore.
1SAM|15|28|Samuel said to him, "The LORD has torn the kingdom of Israel from you today and has given it to one of your neighbors-to one better than you.
1SAM|15|29|He who is the Glory of Israel does not lie or change his mind; for he is not a man, that he should change his mind."
1SAM|15|30|Saul replied, "I have sinned. But please honor me before the elders of my people and before Israel; come back with me, so that I may worship the LORD your God."
1SAM|15|31|So Samuel went back with Saul, and Saul worshiped the LORD.
1SAM|15|32|Then Samuel said, "Bring me Agag king of the Amalekites." Agag came to him confidently, thinking, "Surely the bitterness of death is past."
1SAM|15|33|But Samuel said, "As your sword has made women childless, so will your mother be childless among women." And Samuel put Agag to death before the LORD at Gilgal.
1SAM|15|34|Then Samuel left for Ramah, but Saul went up to his home in Gibeah of Saul.
1SAM|15|35|Until the day Samuel died, he did not go to see Saul again, though Samuel mourned for him. And the LORD was grieved that he had made Saul king over Israel.
1SAM|16|1|The LORD said to Samuel, "How long will you mourn for Saul, since I have rejected him as king over Israel? Fill your horn with oil and be on your way; I am sending you to Jesse of Bethlehem. I have chosen one of his sons to be king."
1SAM|16|2|But Samuel said, "How can I go? Saul will hear about it and kill me." The LORD said, "Take a heifer with you and say, 'I have come to sacrifice to the LORD.'
1SAM|16|3|Invite Jesse to the sacrifice, and I will show you what to do. You are to anoint for me the one I indicate."
1SAM|16|4|Samuel did what the LORD said. When he arrived at Bethlehem, the elders of the town trembled when they met him. They asked, "Do you come in peace?"
1SAM|16|5|Samuel replied, "Yes, in peace; I have come to sacrifice to the LORD. Consecrate yourselves and come to the sacrifice with me." Then he consecrated Jesse and his sons and invited them to the sacrifice.
1SAM|16|6|When they arrived, Samuel saw Eliab and thought, "Surely the LORD's anointed stands here before the LORD."
1SAM|16|7|But the LORD said to Samuel, "Do not consider his appearance or his height, for I have rejected him. The LORD does not look at the things man looks at. Man looks at the outward appearance, but the LORD looks at the heart."
1SAM|16|8|Then Jesse called Abinadab and had him pass in front of Samuel. But Samuel said, "The LORD has not chosen this one either."
1SAM|16|9|Jesse then had Shammah pass by, but Samuel said, "Nor has the LORD chosen this one."
1SAM|16|10|Jesse had seven of his sons pass before Samuel, but Samuel said to him, "The LORD has not chosen these."
1SAM|16|11|So he asked Jesse, "Are these all the sons you have?There is still the youngest," Jesse answered, "but he is tending the sheep." Samuel said, "Send for him; we will not sit down until he arrives."
1SAM|16|12|So he sent and had him brought in. He was ruddy, with a fine appearance and handsome features. Then the LORD said, "Rise and anoint him; he is the one."
1SAM|16|13|So Samuel took the horn of oil and anointed him in the presence of his brothers, and from that day on the Spirit of the LORD came upon David in power. Samuel then went to Ramah.
1SAM|16|14|Now the Spirit of the LORD had departed from Saul, and an evil spirit from the LORD tormented him.
1SAM|16|15|Saul's attendants said to him, "See, an evil spirit from God is tormenting you.
1SAM|16|16|Let our lord command his servants here to search for someone who can play the harp. He will play when the evil spirit from God comes upon you, and you will feel better."
1SAM|16|17|So Saul said to his attendants, "Find someone who plays well and bring him to me."
1SAM|16|18|One of the servants answered, "I have seen a son of Jesse of Bethlehem who knows how to play the harp. He is a brave man and a warrior. He speaks well and is a fine-looking man. And the LORD is with him."
1SAM|16|19|Then Saul sent messengers to Jesse and said, "Send me your son David, who is with the sheep."
1SAM|16|20|So Jesse took a donkey loaded with bread, a skin of wine and a young goat and sent them with his son David to Saul.
1SAM|16|21|David came to Saul and entered his service. Saul liked him very much, and David became one of his armor-bearers.
1SAM|16|22|Then Saul sent word to Jesse, saying, "Allow David to remain in my service, for I am pleased with him."
1SAM|16|23|Whenever the spirit from God came upon Saul, David would take his harp and play. Then relief would come to Saul; he would feel better, and the evil spirit would leave him.
1SAM|17|1|Now the Philistines gathered their forces for war and assembled at Socoh in Judah. They pitched camp at Ephes Dammim, between Socoh and Azekah.
1SAM|17|2|Saul and the Israelites assembled and camped in the Valley of Elah and drew up their battle line to meet the Philistines.
1SAM|17|3|The Philistines occupied one hill and the Israelites another, with the valley between them.
1SAM|17|4|A champion named Goliath, who was from Gath, came out of the Philistine camp. He was over nine feet tall.
1SAM|17|5|He had a bronze helmet on his head and wore a coat of scale armor of bronze weighing five thousand shekels;
1SAM|17|6|on his legs he wore bronze greaves, and a bronze javelin was slung on his back.
1SAM|17|7|His spear shaft was like a weaver's rod, and its iron point weighed six hundred shekels. His shield bearer went ahead of him.
1SAM|17|8|Goliath stood and shouted to the ranks of Israel, "Why do you come out and line up for battle? Am I not a Philistine, and are you not the servants of Saul? Choose a man and have him come down to me.
1SAM|17|9|If he is able to fight and kill me, we will become your subjects; but if I overcome him and kill him, you will become our subjects and serve us."
1SAM|17|10|Then the Philistine said, "This day I defy the ranks of Israel! Give me a man and let us fight each other."
1SAM|17|11|On hearing the Philistine's words, Saul and all the Israelites were dismayed and terrified.
1SAM|17|12|Now David was the son of an Ephrathite named Jesse, who was from Bethlehem in Judah. Jesse had eight sons, and in Saul's time he was old and well advanced in years.
1SAM|17|13|Jesse's three oldest sons had followed Saul to the war: The firstborn was Eliab; the second, Abinadab; and the third, Shammah.
1SAM|17|14|David was the youngest. The three oldest followed Saul,
1SAM|17|15|but David went back and forth from Saul to tend his father's sheep at Bethlehem.
1SAM|17|16|For forty days the Philistine came forward every morning and evening and took his stand.
1SAM|17|17|Now Jesse said to his son David, "Take this ephah of roasted grain and these ten loaves of bread for your brothers and hurry to their camp.
1SAM|17|18|Take along these ten cheeses to the commander of their unit. See how your brothers are and bring back some assurance from them.
1SAM|17|19|They are with Saul and all the men of Israel in the Valley of Elah, fighting against the Philistines."
1SAM|17|20|Early in the morning David left the flock with a shepherd, loaded up and set out, as Jesse had directed. He reached the camp as the army was going out to its battle positions, shouting the war cry.
1SAM|17|21|Israel and the Philistines were drawing up their lines facing each other.
1SAM|17|22|David left his things with the keeper of supplies, ran to the battle lines and greeted his brothers.
1SAM|17|23|As he was talking with them, Goliath, the Philistine champion from Gath, stepped out from his lines and shouted his usual defiance, and David heard it.
1SAM|17|24|When the Israelites saw the man, they all ran from him in great fear.
1SAM|17|25|Now the Israelites had been saying, "Do you see how this man keeps coming out? He comes out to defy Israel. The king will give great wealth to the man who kills him. He will also give him his daughter in marriage and will exempt his father's family from taxes in Israel."
1SAM|17|26|David asked the men standing near him, "What will be done for the man who kills this Philistine and removes this disgrace from Israel? Who is this uncircumcised Philistine that he should defy the armies of the living God?"
1SAM|17|27|They repeated to him what they had been saying and told him, "This is what will be done for the man who kills him."
1SAM|17|28|When Eliab, David's oldest brother, heard him speaking with the men, he burned with anger at him and asked, "Why have you come down here? And with whom did you leave those few sheep in the desert? I know how conceited you are and how wicked your heart is; you came down only to watch the battle."
1SAM|17|29|"Now what have I done?" said David. "Can't I even speak?"
1SAM|17|30|He then turned away to someone else and brought up the same matter, and the men answered him as before.
1SAM|17|31|What David said was overheard and reported to Saul, and Saul sent for him.
1SAM|17|32|David said to Saul, "Let no one lose heart on account of this Philistine; your servant will go and fight him."
1SAM|17|33|Saul replied, "You are not able to go out against this Philistine and fight him; you are only a boy, and he has been a fighting man from his youth."
1SAM|17|34|But David said to Saul, "Your servant has been keeping his father's sheep. When a lion or a bear came and carried off a sheep from the flock,
1SAM|17|35|I went after it, struck it and rescued the sheep from its mouth. When it turned on me, I seized it by its hair, struck it and killed it.
1SAM|17|36|Your servant has killed both the lion and the bear; this uncircumcised Philistine will be like one of them, because he has defied the armies of the living God.
1SAM|17|37|The LORD who delivered me from the paw of the lion and the paw of the bear will deliver me from the hand of this Philistine." Saul said to David, "Go, and the LORD be with you."
1SAM|17|38|Then Saul dressed David in his own tunic. He put a coat of armor on him and a bronze helmet on his head.
1SAM|17|39|David fastened on his sword over the tunic and tried walking around, because he was not used to them. "I cannot go in these," he said to Saul, "because I am not used to them." So he took them off.
1SAM|17|40|Then he took his staff in his hand, chose five smooth stones from the stream, put them in the pouch of his shepherd's bag and, with his sling in his hand, approached the Philistine.
1SAM|17|41|Meanwhile, the Philistine, with his shield bearer in front of him, kept coming closer to David.
1SAM|17|42|He looked David over and saw that he was only a boy, ruddy and handsome, and he despised him.
1SAM|17|43|He said to David, "Am I a dog, that you come at me with sticks?" And the Philistine cursed David by his gods.
1SAM|17|44|"Come here," he said, "and I'll give your flesh to the birds of the air and the beasts of the field!"
1SAM|17|45|David said to the Philistine, "You come against me with sword and spear and javelin, but I come against you in the name of the LORD Almighty, the God of the armies of Israel, whom you have defied.
1SAM|17|46|This day the LORD will hand you over to me, and I'll strike you down and cut off your head. Today I will give the carcasses of the Philistine army to the birds of the air and the beasts of the earth, and the whole world will know that there is a God in Israel.
1SAM|17|47|All those gathered here will know that it is not by sword or spear that the LORD saves; for the battle is the LORD's, and he will give all of you into our hands."
1SAM|17|48|As the Philistine moved closer to attack him, David ran quickly toward the battle line to meet him.
1SAM|17|49|Reaching into his bag and taking out a stone, he slung it and struck the Philistine on the forehead. The stone sank into his forehead, and he fell facedown on the ground.
1SAM|17|50|So David triumphed over the Philistine with a sling and a stone; without a sword in his hand he struck down the Philistine and killed him.
1SAM|17|51|David ran and stood over him. He took hold of the Philistine's sword and drew it from the scabbard. After he killed him, he cut off his head with the sword. When the Philistines saw that their hero was dead, they turned and ran.
1SAM|17|52|Then the men of Israel and Judah surged forward with a shout and pursued the Philistines to the entrance of Gath and to the gates of Ekron. Their dead were strewn along the Shaaraim road to Gath and Ekron.
1SAM|17|53|When the Israelites returned from chasing the Philistines, they plundered their camp.
1SAM|17|54|David took the Philistine's head and brought it to Jerusalem, and he put the Philistine's weapons in his own tent.
1SAM|17|55|As Saul watched David going out to meet the Philistine, he said to Abner, commander of the army, "Abner, whose son is that young man?" Abner replied, "As surely as you live, O king, I don't know."
1SAM|17|56|The king said, "Find out whose son this young man is."
1SAM|17|57|As soon as David returned from killing the Philistine, Abner took him and brought him before Saul, with David still holding the Philistine's head.
1SAM|17|58|"Whose son are you, young man?" Saul asked him. David said, "I am the son of your servant Jesse of Bethlehem."
1SAM|18|1|After David had finished talking with Saul, Jonathan became one in spirit with David, and he loved him as himself.
1SAM|18|2|From that day Saul kept David with him and did not let him return to his father's house.
1SAM|18|3|And Jonathan made a covenant with David because he loved him as himself.
1SAM|18|4|Jonathan took off the robe he was wearing and gave it to David, along with his tunic, and even his sword, his bow and his belt.
1SAM|18|5|Whatever Saul sent him to do, David did it so successfully that Saul gave him a high rank in the army. This pleased all the people, and Saul's officers as well.
1SAM|18|6|When the men were returning home after David had killed the Philistine, the women came out from all the towns of Israel to meet King Saul with singing and dancing, with joyful songs and with tambourines and lutes.
1SAM|18|7|As they danced, they sang: "Saul has slain his thousands, and David his tens of thousands."
1SAM|18|8|Saul was very angry; this refrain galled him. "They have credited David with tens of thousands," he thought, "but me with only thousands. What more can he get but the kingdom?"
1SAM|18|9|And from that time on Saul kept a jealous eye on David.
1SAM|18|10|The next day an evil spirit from God came forcefully upon Saul. He was prophesying in his house, while David was playing the harp, as he usually did. Saul had a spear in his hand
1SAM|18|11|and he hurled it, saying to himself, "I'll pin David to the wall." But David eluded him twice.
1SAM|18|12|Saul was afraid of David, because the LORD was with David but had left Saul.
1SAM|18|13|So he sent David away from him and gave him command over a thousand men, and David led the troops in their campaigns.
1SAM|18|14|In everything he did he had great success, because the LORD was with him.
1SAM|18|15|When Saul saw how successful he was, he was afraid of him.
1SAM|18|16|But all Israel and Judah loved David, because he led them in their campaigns.
1SAM|18|17|Saul said to David, "Here is my older daughter Merab. I will give her to you in marriage; only serve me bravely and fight the battles of the LORD." For Saul said to himself, "I will not raise a hand against him. Let the Philistines do that!"
1SAM|18|18|But David said to Saul, "Who am I, and what is my family or my father's clan in Israel, that I should become the king's son-in-law?"
1SAM|18|19|So when the time came for Merab, Saul's daughter, to be given to David, she was given in marriage to Adriel of Meholah.
1SAM|18|20|Now Saul's daughter Michal was in love with David, and when they told Saul about it, he was pleased.
1SAM|18|21|"I will give her to him," he thought, "so that she may be a snare to him and so that the hand of the Philistines may be against him." So Saul said to David, "Now you have a second opportunity to become my son-in-law."
1SAM|18|22|Then Saul ordered his attendants: "Speak to David privately and say, 'Look, the king is pleased with you, and his attendants all like you; now become his son-in-law.'"
1SAM|18|23|They repeated these words to David. But David said, "Do you think it is a small matter to become the king's son-in-law? I'm only a poor man and little known."
1SAM|18|24|When Saul's servants told him what David had said,
1SAM|18|25|Saul replied, "Say to David, 'The king wants no other price for the bride than a hundred Philistine foreskins, to take revenge on his enemies.'" Saul's plan was to have David fall by the hands of the Philistines.
1SAM|18|26|When the attendants told David these things, he was pleased to become the king's son-in-law. So before the allotted time elapsed,
1SAM|18|27|David and his men went out and killed two hundred Philistines. He brought their foreskins and presented the full number to the king so that he might become the king's son-in-law. Then Saul gave him his daughter Michal in marriage.
1SAM|18|28|When Saul realized that the LORD was with David and that his daughter Michal loved David,
1SAM|18|29|Saul became still more afraid of him, and he remained his enemy the rest of his days.
1SAM|18|30|The Philistine commanders continued to go out to battle, and as often as they did, David met with more success than the rest of Saul's officers, and his name became well known.
1SAM|19|1|Saul told his son Jonathan and all the attendants to kill David. But Jonathan was very fond of David
1SAM|19|2|and warned him, "My father Saul is looking for a chance to kill you. Be on your guard tomorrow morning; go into hiding and stay there.
1SAM|19|3|I will go out and stand with my father in the field where you are. I'll speak to him about you and will tell you what I find out."
1SAM|19|4|Jonathan spoke well of David to Saul his father and said to him, "Let not the king do wrong to his servant David; he has not wronged you, and what he has done has benefited you greatly.
1SAM|19|5|He took his life in his hands when he killed the Philistine. The LORD won a great victory for all Israel, and you saw it and were glad. Why then would you do wrong to an innocent man like David by killing him for no reason?"
1SAM|19|6|Saul listened to Jonathan and took this oath: "As surely as the LORD lives, David will not be put to death."
1SAM|19|7|So Jonathan called David and told him the whole conversation. He brought him to Saul, and David was with Saul as before.
1SAM|19|8|Once more war broke out, and David went out and fought the Philistines. He struck them with such force that they fled before him.
1SAM|19|9|But an evil spirit from the LORD came upon Saul as he was sitting in his house with his spear in his hand. While David was playing the harp,
1SAM|19|10|Saul tried to pin him to the wall with his spear, but David eluded him as Saul drove the spear into the wall. That night David made good his escape.
1SAM|19|11|Saul sent men to David's house to watch it and to kill him in the morning. But Michal, David's wife, warned him, "If you don't run for your life tonight, tomorrow you'll be killed."
1SAM|19|12|So Michal let David down through a window, and he fled and escaped.
1SAM|19|13|Then Michal took an idol and laid it on the bed, covering it with a garment and putting some goats' hair at the head.
1SAM|19|14|When Saul sent the men to capture David, Michal said, "He is ill."
1SAM|19|15|Then Saul sent the men back to see David and told them, "Bring him up to me in his bed so that I may kill him."
1SAM|19|16|But when the men entered, there was the idol in the bed, and at the head was some goats' hair.
1SAM|19|17|Saul said to Michal, "Why did you deceive me like this and send my enemy away so that he escaped?" Michal told him, "He said to me, 'Let me get away. Why should I kill you?'"
1SAM|19|18|When David had fled and made his escape, he went to Samuel at Ramah and told him all that Saul had done to him. Then he and Samuel went to Naioth and stayed there.
1SAM|19|19|Word came to Saul: "David is in Naioth at Ramah";
1SAM|19|20|so he sent men to capture him. But when they saw a group of prophets prophesying, with Samuel standing there as their leader, the Spirit of God came upon Saul's men and they also prophesied.
1SAM|19|21|Saul was told about it, and he sent more men, and they prophesied too. Saul sent men a third time, and they also prophesied.
1SAM|19|22|Finally, he himself left for Ramah and went to the great cistern at Secu. And he asked, "Where are Samuel and David?Over in Naioth at Ramah," they said.
1SAM|19|23|So Saul went to Naioth at Ramah. But the Spirit of God came even upon him, and he walked along prophesying until he came to Naioth.
1SAM|19|24|He stripped off his robes and also prophesied in Samuel's presence. He lay that way all that day and night. This is why people say, "Is Saul also among the prophets?"
1SAM|20|1|Then David fled from Naioth at Ramah and went to Jonathan and asked, "What have I done? What is my crime? How have I wronged your father, that he is trying to take my life?"
1SAM|20|2|"Never!" Jonathan replied. "You are not going to die! Look, my father doesn't do anything, great or small, without confiding in me. Why would he hide this from me? It's not so!"
1SAM|20|3|But David took an oath and said, "Your father knows very well that I have found favor in your eyes, and he has said to himself, 'Jonathan must not know this or he will be grieved.' Yet as surely as the LORD lives and as you live, there is only a step between me and death."
1SAM|20|4|Jonathan said to David, "Whatever you want me to do, I'll do for you."
1SAM|20|5|So David said, "Look, tomorrow is the New Moon festival, and I am supposed to dine with the king; but let me go and hide in the field until the evening of the day after tomorrow.
1SAM|20|6|If your father misses me at all, tell him, 'David earnestly asked my permission to hurry to Bethlehem, his hometown, because an annual sacrifice is being made there for his whole clan.'
1SAM|20|7|If he says, 'Very well,' then your servant is safe. But if he loses his temper, you can be sure that he is determined to harm me.
1SAM|20|8|As for you, show kindness to your servant, for you have brought him into a covenant with you before the LORD. If I am guilty, then kill me yourself! Why hand me over to your father?"
1SAM|20|9|"Never!" Jonathan said. "If I had the least inkling that my father was determined to harm you, wouldn't I tell you?"
1SAM|20|10|David asked, "Who will tell me if your father answers you harshly?"
1SAM|20|11|"Come," Jonathan said, "let's go out into the field." So they went there together.
1SAM|20|12|Then Jonathan said to David: "By the LORD, the God of Israel, I will surely sound out my father by this time the day after tomorrow! If he is favorably disposed toward you, will I not send you word and let you know?
1SAM|20|13|But if my father is inclined to harm you, may the LORD deal with me, be it ever so severely, if I do not let you know and send you away safely. May the LORD be with you as he has been with my father.
1SAM|20|14|But show me unfailing kindness like that of the LORD as long as I live, so that I may not be killed,
1SAM|20|15|and do not ever cut off your kindness from my family-not even when the LORD has cut off every one of David's enemies from the face of the earth."
1SAM|20|16|So Jonathan made a covenant with the house of David, saying, "May the LORD call David's enemies to account."
1SAM|20|17|And Jonathan had David reaffirm his oath out of love for him, because he loved him as he loved himself.
1SAM|20|18|Then Jonathan said to David: "Tomorrow is the New Moon festival. You will be missed, because your seat will be empty.
1SAM|20|19|The day after tomorrow, toward evening, go to the place where you hid when this trouble began, and wait by the stone Ezel.
1SAM|20|20|I will shoot three arrows to the side of it, as though I were shooting at a target.
1SAM|20|21|Then I will send a boy and say, 'Go, find the arrows.' If I say to him, 'Look, the arrows are on this side of you; bring them here,' then come, because, as surely as the LORD lives, you are safe; there is no danger.
1SAM|20|22|But if I say to the boy, 'Look, the arrows are beyond you,' then you must go, because the LORD has sent you away.
1SAM|20|23|And about the matter you and I discussed-remember, the LORD is witness between you and me forever."
1SAM|20|24|So David hid in the field, and when the New Moon festival came, the king sat down to eat.
1SAM|20|25|He sat in his customary place by the wall, opposite Jonathan, and Abner sat next to Saul, but David's place was empty.
1SAM|20|26|Saul said nothing that day, for he thought, "Something must have happened to David to make him ceremonially unclean-surely he is unclean."
1SAM|20|27|But the next day, the second day of the month, David's place was empty again. Then Saul said to his son Jonathan, "Why hasn't the son of Jesse come to the meal, either yesterday or today?"
1SAM|20|28|Jonathan answered, "David earnestly asked me for permission to go to Bethlehem.
1SAM|20|29|He said, 'Let me go, because our family is observing a sacrifice in the town and my brother has ordered me to be there. If I have found favor in your eyes, let me get away to see my brothers.' That is why he has not come to the king's table."
1SAM|20|30|Saul's anger flared up at Jonathan and he said to him, "You son of a perverse and rebellious woman! Don't I know that you have sided with the son of Jesse to your own shame and to the shame of the mother who bore you?
1SAM|20|31|As long as the son of Jesse lives on this earth, neither you nor your kingdom will be established. Now send and bring him to me, for he must die!"
1SAM|20|32|"Why should he be put to death? What has he done?" Jonathan asked his father.
1SAM|20|33|But Saul hurled his spear at him to kill him. Then Jonathan knew that his father intended to kill David.
1SAM|20|34|Jonathan got up from the table in fierce anger; on that second day of the month he did not eat, because he was grieved at his father's shameful treatment of David.
1SAM|20|35|In the morning Jonathan went out to the field for his meeting with David. He had a small boy with him,
1SAM|20|36|and he said to the boy, "Run and find the arrows I shoot." As the boy ran, he shot an arrow beyond him.
1SAM|20|37|When the boy came to the place where Jonathan's arrow had fallen, Jonathan called out after him, "Isn't the arrow beyond you?"
1SAM|20|38|Then he shouted, "Hurry! Go quickly! Don't stop!" The boy picked up the arrow and returned to his master.
1SAM|20|39|(The boy knew nothing of all this; only Jonathan and David knew.)
1SAM|20|40|Then Jonathan gave his weapons to the boy and said, "Go, carry them back to town."
1SAM|20|41|After the boy had gone, David got up from the south side of the stone and bowed down before Jonathan three times, with his face to the ground. Then they kissed each other and wept together-but David wept the most.
1SAM|20|42|Jonathan said to David, "Go in peace, for we have sworn friendship with each other in the name of the LORD, saying, 'The LORD is witness between you and me, and between your descendants and my descendants forever.'" Then David left, and Jonathan went back to the town.
1SAM|21|1|David went to Nob, to Ahimelech the priest. Ahimelech trembled when he met him, and asked, "Why are you alone? Why is no one with you?"
1SAM|21|2|David answered Ahimelech the priest, "The king charged me with a certain matter and said to me, 'No one is to know anything about your mission and your instructions.' As for my men, I have told them to meet me at a certain place.
1SAM|21|3|Now then, what do you have on hand? Give me five loaves of bread, or whatever you can find."
1SAM|21|4|But the priest answered David, "I don't have any ordinary bread on hand; however, there is some consecrated bread here-provided the men have kept themselves from women."
1SAM|21|5|David replied, "Indeed women have been kept from us, as usual whenever I set out. The men's things are holy even on missions that are not holy. How much more so today!"
1SAM|21|6|So the priest gave him the consecrated bread, since there was no bread there except the bread of the Presence that had been removed from before the LORD and replaced by hot bread on the day it was taken away.
1SAM|21|7|Now one of Saul's servants was there that day, detained before the LORD; he was Doeg the Edomite, Saul's head shepherd.
1SAM|21|8|David asked Ahimelech, "Don't you have a spear or a sword here? I haven't brought my sword or any other weapon, because the king's business was urgent."
1SAM|21|9|The priest replied, "The sword of Goliath the Philistine, whom you killed in the Valley of Elah, is here; it is wrapped in a cloth behind the ephod. If you want it, take it; there is no sword here but that one." David said, "There is none like it; give it to me."
1SAM|21|10|That day David fled from Saul and went to Achish king of Gath.
1SAM|21|11|But the servants of Achish said to him, "Isn't this David, the king of the land? Isn't he the one they sing about in their dances: "'Saul has slain his thousands, and David his tens of thousands'?"
1SAM|21|12|David took these words to heart and was very much afraid of Achish king of Gath.
1SAM|21|13|So he pretended to be insane in their presence; and while he was in their hands he acted like a madman, making marks on the doors of the gate and letting saliva run down his beard.
1SAM|21|14|Achish said to his servants, "Look at the man! He is insane! Why bring him to me?
1SAM|21|15|Am I so short of madmen that you have to bring this fellow here to carry on like this in front of me? Must this man come into my house?"
1SAM|22|1|David left Gath and escaped to the cave of Adullam. When his brothers and his father's household heard about it, they went down to him there.
1SAM|22|2|All those who were in distress or in debt or discontented gathered around him, and he became their leader. About four hundred men were with him.
1SAM|22|3|From there David went to Mizpah in Moab and said to the king of Moab, "Would you let my father and mother come and stay with you until I learn what God will do for me?"
1SAM|22|4|So he left them with the king of Moab, and they stayed with him as long as David was in the stronghold.
1SAM|22|5|But the prophet Gad said to David, "Do not stay in the stronghold. Go into the land of Judah." So David left and went to the forest of Hereth.
1SAM|22|6|Now Saul heard that David and his men had been discovered. And Saul, spear in hand, was seated under the tamarisk tree on the hill at Gibeah, with all his officials standing around him.
1SAM|22|7|Saul said to them, "Listen, men of Benjamin! Will the son of Jesse give all of you fields and vineyards? Will he make all of you commanders of thousands and commanders of hundreds?
1SAM|22|8|Is that why you have all conspired against me? No one tells me when my son makes a covenant with the son of Jesse. None of you is concerned about me or tells me that my son has incited my servant to lie in wait for me, as he does today."
1SAM|22|9|But Doeg the Edomite, who was standing with Saul's officials, said, "I saw the son of Jesse come to Ahimelech son of Ahitub at Nob.
1SAM|22|10|Ahimelech inquired of the LORD for him; he also gave him provisions and the sword of Goliath the Philistine."
1SAM|22|11|Then the king sent for the priest Ahimelech son of Ahitub and his father's whole family, who were the priests at Nob, and they all came to the king.
1SAM|22|12|Saul said, "Listen now, son of Ahitub.Yes, my lord," he answered.
1SAM|22|13|Saul said to him, "Why have you conspired against me, you and the son of Jesse, giving him bread and a sword and inquiring of God for him, so that he has rebelled against me and lies in wait for me, as he does today?"
1SAM|22|14|Ahimelech answered the king, "Who of all your servants is as loyal as David, the king's son-in-law, captain of your bodyguard and highly respected in your household?
1SAM|22|15|Was that day the first time I inquired of God for him? Of course not! Let not the king accuse your servant or any of his father's family, for your servant knows nothing at all about this whole affair."
1SAM|22|16|But the king said, "You will surely die, Ahimelech, you and your father's whole family."
1SAM|22|17|Then the king ordered the guards at his side: "Turn and kill the priests of the LORD, because they too have sided with David. They knew he was fleeing, yet they did not tell me." But the king's officials were not willing to raise a hand to strike the priests of the LORD.
1SAM|22|18|The king then ordered Doeg, "You turn and strike down the priests." So Doeg the Edomite turned and struck them down. That day he killed eighty-five men who wore the linen ephod.
1SAM|22|19|He also put to the sword Nob, the town of the priests, with its men and women, its children and infants, and its cattle, donkeys and sheep.
1SAM|22|20|But Abiathar, a son of Ahimelech son of Ahitub, escaped and fled to join David.
1SAM|22|21|He told David that Saul had killed the priests of the LORD.
1SAM|22|22|Then David said to Abiathar: "That day, when Doeg the Edomite was there, I knew he would be sure to tell Saul. I am responsible for the death of your father's whole family.
1SAM|22|23|Stay with me; don't be afraid; the man who is seeking your life is seeking mine also. You will be safe with me."
1SAM|23|1|When David was told, "Look, the Philistines are fighting against Keilah and are looting the threshing floors,"
1SAM|23|2|he inquired of the LORD, saying, "Shall I go and attack these Philistines?" The LORD answered him, "Go, attack the Philistines and save Keilah."
1SAM|23|3|But David's men said to him, "Here in Judah we are afraid. How much more, then, if we go to Keilah against the Philistine forces!"
1SAM|23|4|Once again David inquired of the LORD, and the LORD answered him, "Go down to Keilah, for I am going to give the Philistines into your hand."
1SAM|23|5|So David and his men went to Keilah, fought the Philistines and carried off their livestock. He inflicted heavy losses on the Philistines and saved the people of Keilah.
1SAM|23|6|(Now Abiathar son of Ahimelech had brought the ephod down with him when he fled to David at Keilah.)
1SAM|23|7|Saul was told that David had gone to Keilah, and he said, "God has handed him over to me, for David has imprisoned himself by entering a town with gates and bars."
1SAM|23|8|And Saul called up all his forces for battle, to go down to Keilah to besiege David and his men.
1SAM|23|9|When David learned that Saul was plotting against him, he said to Abiathar the priest, "Bring the ephod."
1SAM|23|10|David said, "O LORD, God of Israel, your servant has heard definitely that Saul plans to come to Keilah and destroy the town on account of me.
1SAM|23|11|Will the citizens of Keilah surrender me to him? Will Saul come down, as your servant has heard? O LORD, God of Israel, tell your servant." And the LORD said, "He will."
1SAM|23|12|Again David asked, "Will the citizens of Keilah surrender me and my men to Saul?" And the LORD said, "They will."
1SAM|23|13|So David and his men, about six hundred in number, left Keilah and kept moving from place to place. When Saul was told that David had escaped from Keilah, he did not go there.
1SAM|23|14|David stayed in the desert strongholds and in the hills of the Desert of Ziph. Day after day Saul searched for him, but God did not give David into his hands.
1SAM|23|15|While David was at Horesh in the Desert of Ziph, he learned that Saul had come out to take his life.
1SAM|23|16|And Saul's son Jonathan went to David at Horesh and helped him find strength in God.
1SAM|23|17|"Don't be afraid," he said. "My father Saul will not lay a hand on you. You will be king over Israel, and I will be second to you. Even my father Saul knows this."
1SAM|23|18|The two of them made a covenant before the LORD. Then Jonathan went home, but David remained at Horesh.
1SAM|23|19|The Ziphites went up to Saul at Gibeah and said, "Is not David hiding among us in the strongholds at Horesh, on the hill of Hakilah, south of Jeshimon?
1SAM|23|20|Now, O king, come down whenever it pleases you to do so, and we will be responsible for handing him over to the king."
1SAM|23|21|Saul replied, "The LORD bless you for your concern for me.
1SAM|23|22|Go and make further preparation. Find out where David usually goes and who has seen him there. They tell me he is very crafty.
1SAM|23|23|Find out about all the hiding places he uses and come back to me with definite information. Then I will go with you; if he is in the area, I will track him down among all the clans of Judah."
1SAM|23|24|So they set out and went to Ziph ahead of Saul. Now David and his men were in the Desert of Maon, in the Arabah south of Jeshimon.
1SAM|23|25|Saul and his men began the search, and when David was told about it, he went down to the rock and stayed in the Desert of Maon. When Saul heard this, he went into the Desert of Maon in pursuit of David.
1SAM|23|26|Saul was going along one side of the mountain, and David and his men were on the other side, hurrying to get away from Saul. As Saul and his forces were closing in on David and his men to capture them,
1SAM|23|27|a messenger came to Saul, saying, "Come quickly! The Philistines are raiding the land."
1SAM|23|28|Then Saul broke off his pursuit of David and went to meet the Philistines. That is why they call this place Sela Hammahlekoth.
1SAM|23|29|And David went up from there and lived in the strongholds of En Gedi.
1SAM|24|1|After Saul returned from pursuing the Philistines, he was told, "David is in the Desert of En Gedi."
1SAM|24|2|So Saul took three thousand chosen men from all Israel and set out to look for David and his men near the Crags of the Wild Goats.
1SAM|24|3|He came to the sheep pens along the way; a cave was there, and Saul went in to relieve himself. David and his men were far back in the cave.
1SAM|24|4|The men said, "This is the day the LORD spoke of when he said to you, 'I will give your enemy into your hands for you to deal with as you wish.'" Then David crept up unnoticed and cut off a corner of Saul's robe.
1SAM|24|5|Afterward, David was conscience-stricken for having cut off a corner of his robe.
1SAM|24|6|He said to his men, "The LORD forbid that I should do such a thing to my master, the LORD's anointed, or lift my hand against him; for he is the anointed of the LORD."
1SAM|24|7|With these words David rebuked his men and did not allow them to attack Saul. And Saul left the cave and went his way.
1SAM|24|8|Then David went out of the cave and called out to Saul, "My lord the king!" When Saul looked behind him, David bowed down and prostrated himself with his face to the ground.
1SAM|24|9|He said to Saul, "Why do you listen when men say, 'David is bent on harming you'?
1SAM|24|10|This day you have seen with your own eyes how the LORD delivered you into my hands in the cave. Some urged me to kill you, but I spared you; I said, 'I will not lift my hand against my master, because he is the LORD's anointed.'
1SAM|24|11|See, my father, look at this piece of your robe in my hand! I cut off the corner of your robe but did not kill you. Now understand and recognize that I am not guilty of wrongdoing or rebellion. I have not wronged you, but you are hunting me down to take my life.
1SAM|24|12|May the LORD judge between you and me. And may the LORD avenge the wrongs you have done to me, but my hand will not touch you.
1SAM|24|13|As the old saying goes, 'From evildoers come evil deeds,' so my hand will not touch you.
1SAM|24|14|"Against whom has the king of Israel come out? Whom are you pursuing? A dead dog? A flea?
1SAM|24|15|May the LORD be our judge and decide between us. May he consider my cause and uphold it; may he vindicate me by delivering me from your hand."
1SAM|24|16|When David finished saying this, Saul asked, "Is that your voice, David my son?" And he wept aloud.
1SAM|24|17|"You are more righteous than I," he said. "You have treated me well, but I have treated you badly.
1SAM|24|18|You have just now told me of the good you did to me; the LORD delivered me into your hands, but you did not kill me.
1SAM|24|19|When a man finds his enemy, does he let him get away unharmed? May the LORD reward you well for the way you treated me today.
1SAM|24|20|I know that you will surely be king and that the kingdom of Israel will be established in your hands.
1SAM|24|21|Now swear to me by the LORD that you will not cut off my descendants or wipe out my name from my father's family."
1SAM|24|22|So David gave his oath to Saul. Then Saul returned home, but David and his men went up to the stronghold.
1SAM|25|1|Now Samuel died, and all Israel assembled and mourned for him; and they buried him at his home in Ramah. Then David moved down into the Desert of Maon.
1SAM|25|2|A certain man in Maon, who had property there at Carmel, was very wealthy. He had a thousand goats and three thousand sheep, which he was shearing in Carmel.
1SAM|25|3|His name was Nabal and his wife's name was Abigail. She was an intelligent and beautiful woman, but her husband, a Calebite, was surly and mean in his dealings.
1SAM|25|4|While David was in the desert, he heard that Nabal was shearing sheep.
1SAM|25|5|So he sent ten young men and said to them, "Go up to Nabal at Carmel and greet him in my name.
1SAM|25|6|Say to him: 'Long life to you! Good health to you and your household! And good health to all that is yours!
1SAM|25|7|"'Now I hear that it is sheep-shearing time. When your shepherds were with us, we did not mistreat them, and the whole time they were at Carmel nothing of theirs was missing.
1SAM|25|8|Ask your own servants and they will tell you. Therefore be favorable toward my young men, since we come at a festive time. Please give your servants and your son David whatever you can find for them.'"
1SAM|25|9|When David's men arrived, they gave Nabal this message in David's name. Then they waited.
1SAM|25|10|Nabal answered David's servants, "Who is this David? Who is this son of Jesse? Many servants are breaking away from their masters these days.
1SAM|25|11|Why should I take my bread and water, and the meat I have slaughtered for my shearers, and give it to men coming from who knows where?"
1SAM|25|12|David's men turned around and went back. When they arrived, they reported every word.
1SAM|25|13|David said to his men, "Put on your swords!" So they put on their swords, and David put on his. About four hundred men went up with David, while two hundred stayed with the supplies.
1SAM|25|14|One of the servants told Nabal's wife Abigail: "David sent messengers from the desert to give our master his greetings, but he hurled insults at them.
1SAM|25|15|Yet these men were very good to us. They did not mistreat us, and the whole time we were out in the fields near them nothing was missing.
1SAM|25|16|Night and day they were a wall around us all the time we were herding our sheep near them.
1SAM|25|17|Now think it over and see what you can do, because disaster is hanging over our master and his whole household. He is such a wicked man that no one can talk to him."
1SAM|25|18|Abigail lost no time. She took two hundred loaves of bread, two skins of wine, five dressed sheep, five seahs of roasted grain, a hundred cakes of raisins and two hundred cakes of pressed figs, and loaded them on donkeys.
1SAM|25|19|Then she told her servants, "Go on ahead; I'll follow you." But she did not tell her husband Nabal.
1SAM|25|20|As she came riding her donkey into a mountain ravine, there were David and his men descending toward her, and she met them.
1SAM|25|21|David had just said, "It's been useless-all my watching over this fellow's property in the desert so that nothing of his was missing. He has paid me back evil for good.
1SAM|25|22|May God deal with David, be it ever so severely, if by morning I leave alive one male of all who belong to him!"
1SAM|25|23|When Abigail saw David, she quickly got off her donkey and bowed down before David with her face to the ground.
1SAM|25|24|She fell at his feet and said: "My lord, let the blame be on me alone. Please let your servant speak to you; hear what your servant has to say.
1SAM|25|25|May my lord pay no attention to that wicked man Nabal. He is just like his name-his name is Fool, and folly goes with him. But as for me, your servant, I did not see the men my master sent.
1SAM|25|26|"Now since the LORD has kept you, my master, from bloodshed and from avenging yourself with your own hands, as surely as the LORD lives and as you live, may your enemies and all who intend to harm my master be like Nabal.
1SAM|25|27|And let this gift, which your servant has brought to my master, be given to the men who follow you.
1SAM|25|28|Please forgive your servant's offense, for the LORD will certainly make a lasting dynasty for my master, because he fights the LORD's battles. Let no wrongdoing be found in you as long as you live.
1SAM|25|29|Even though someone is pursuing you to take your life, the life of my master will be bound securely in the bundle of the living by the LORD your God. But the lives of your enemies he will hurl away as from the pocket of a sling.
1SAM|25|30|When the LORD has done for my master every good thing he promised concerning him and has appointed him leader over Israel,
1SAM|25|31|my master will not have on his conscience the staggering burden of needless bloodshed or of having avenged himself. And when the LORD has brought my master success, remember your servant."
1SAM|25|32|David said to Abigail, "Praise be to the LORD, the God of Israel, who has sent you today to meet me.
1SAM|25|33|May you be blessed for your good judgment and for keeping me from bloodshed this day and from avenging myself with my own hands.
1SAM|25|34|Otherwise, as surely as the LORD, the God of Israel, lives, who has kept me from harming you, if you had not come quickly to meet me, not one male belonging to Nabal would have been left alive by daybreak."
1SAM|25|35|Then David accepted from her hand what she had brought him and said, "Go home in peace. I have heard your words and granted your request."
1SAM|25|36|When Abigail went to Nabal, he was in the house holding a banquet like that of a king. He was in high spirits and very drunk. So she told him nothing until daybreak.
1SAM|25|37|Then in the morning, when Nabal was sober, his wife told him all these things, and his heart failed him and he became like a stone.
1SAM|25|38|About ten days later, the LORD struck Nabal and he died.
1SAM|25|39|When David heard that Nabal was dead, he said, "Praise be to the LORD, who has upheld my cause against Nabal for treating me with contempt. He has kept his servant from doing wrong and has brought Nabal's wrongdoing down on his own head." Then David sent word to Abigail, asking her to become his wife.
1SAM|25|40|His servants went to Carmel and said to Abigail, "David has sent us to you to take you to become his wife."
1SAM|25|41|She bowed down with her face to the ground and said, "Here is your maidservant, ready to serve you and wash the feet of my master's servants."
1SAM|25|42|Abigail quickly got on a donkey and, attended by her five maids, went with David's messengers and became his wife.
1SAM|25|43|David had also married Ahinoam of Jezreel, and they both were his wives.
1SAM|25|44|But Saul had given his daughter Michal, David's wife, to Paltiel son of Laish, who was from Gallim.
1SAM|26|1|The Ziphites went to Saul at Gibeah and said, "Is not David hiding on the hill of Hakilah, which faces Jeshimon?"
1SAM|26|2|So Saul went down to the Desert of Ziph, with his three thousand chosen men of Israel, to search there for David.
1SAM|26|3|Saul made his camp beside the road on the hill of Hakilah facing Jeshimon, but David stayed in the desert. When he saw that Saul had followed him there,
1SAM|26|4|he sent out scouts and learned that Saul had definitely arrived.
1SAM|26|5|Then David set out and went to the place where Saul had camped. He saw where Saul and Abner son of Ner, the commander of the army, had lain down. Saul was lying inside the camp, with the army encamped around him.
1SAM|26|6|David then asked Ahimelech the Hittite and Abishai son of Zeruiah, Joab's brother, "Who will go down into the camp with me to Saul?I'll go with you," said Abishai.
1SAM|26|7|So David and Abishai went to the army by night, and there was Saul, lying asleep inside the camp with his spear stuck in the ground near his head. Abner and the soldiers were lying around him.
1SAM|26|8|Abishai said to David, "Today God has delivered your enemy into your hands. Now let me pin him to the ground with one thrust of my spear; I won't strike him twice."
1SAM|26|9|But David said to Abishai, "Don't destroy him! Who can lay a hand on the LORD's anointed and be guiltless?
1SAM|26|10|As surely as the LORD lives," he said, "the LORD himself will strike him; either his time will come and he will die, or he will go into battle and perish.
1SAM|26|11|But the LORD forbid that I should lay a hand on the LORD's anointed. Now get the spear and water jug that are near his head, and let's go."
1SAM|26|12|So David took the spear and water jug near Saul's head, and they left. No one saw or knew about it, nor did anyone wake up. They were all sleeping, because the LORD had put them into a deep sleep.
1SAM|26|13|Then David crossed over to the other side and stood on top of the hill some distance away; there was a wide space between them.
1SAM|26|14|He called out to the army and to Abner son of Ner, "Aren't you going to answer me, Abner?" Abner replied, "Who are you who calls to the king?"
1SAM|26|15|David said, "You're a man, aren't you? And who is like you in Israel? Why didn't you guard your lord the king? Someone came to destroy your lord the king.
1SAM|26|16|What you have done is not good. As surely as the LORD lives, you and your men deserve to die, because you did not guard your master, the LORD's anointed. Look around you. Where are the king's spear and water jug that were near his head?"
1SAM|26|17|Saul recognized David's voice and said, "Is that your voice, David my son?" David replied, "Yes it is, my lord the king."
1SAM|26|18|And he added, "Why is my lord pursuing his servant? What have I done, and what wrong am I guilty of?
1SAM|26|19|Now let my lord the king listen to his servant's words. If the LORD has incited you against me, then may he accept an offering. If, however, men have done it, may they be cursed before the LORD! They have now driven me from my share in the LORD's inheritance and have said, 'Go, serve other gods.'
1SAM|26|20|Now do not let my blood fall to the ground far from the presence of the LORD. The king of Israel has come out to look for a flea-as one hunts a partridge in the mountains."
1SAM|26|21|Then Saul said, "I have sinned. Come back, David my son. Because you considered my life precious today, I will not try to harm you again. Surely I have acted like a fool and have erred greatly."
1SAM|26|22|"Here is the king's spear," David answered. "Let one of your young men come over and get it.
1SAM|26|23|The LORD rewards every man for his righteousness and faithfulness. The LORD delivered you into my hands today, but I would not lay a hand on the LORD's anointed.
1SAM|26|24|As surely as I valued your life today, so may the LORD value my life and deliver me from all trouble."
1SAM|26|25|Then Saul said to David, "May you be blessed, my son David; you will do great things and surely triumph." So David went on his way, and Saul returned home.
1SAM|27|1|But David thought to himself, "One of these days I will be destroyed by the hand of Saul. The best thing I can do is to escape to the land of the Philistines. Then Saul will give up searching for me anywhere in Israel, and I will slip out of his hand."
1SAM|27|2|So David and the six hundred men with him left and went over to Achish son of Maoch king of Gath.
1SAM|27|3|David and his men settled in Gath with Achish. Each man had his family with him, and David had his two wives: Ahinoam of Jezreel and Abigail of Carmel, the widow of Nabal.
1SAM|27|4|When Saul was told that David had fled to Gath, he no longer searched for him.
1SAM|27|5|Then David said to Achish, "If I have found favor in your eyes, let a place be assigned to me in one of the country towns, that I may live there. Why should your servant live in the royal city with you?"
1SAM|27|6|So on that day Achish gave him Ziklag, and it has belonged to the kings of Judah ever since.
1SAM|27|7|David lived in Philistine territory a year and four months.
1SAM|27|8|Now David and his men went up and raided the Geshurites, the Girzites and the Amalekites. (From ancient times these peoples had lived in the land extending to Shur and Egypt.)
1SAM|27|9|Whenever David attacked an area, he did not leave a man or woman alive, but took sheep and cattle, donkeys and camels, and clothes. Then he returned to Achish.
1SAM|27|10|When Achish asked, "Where did you go raiding today?" David would say, "Against the Negev of Judah" or "Against the Negev of Jerahmeel" or "Against the Negev of the Kenites."
1SAM|27|11|He did not leave a man or woman alive to be brought to Gath, for he thought, "They might inform on us and say, 'This is what David did.'" And such was his practice as long as he lived in Philistine territory.
1SAM|27|12|Achish trusted David and said to himself, "He has become so odious to his people, the Israelites, that he will be my servant forever."
1SAM|28|1|In those days the Philistines gathered their forces to fight against Israel. Achish said to David, "You must understand that you and your men will accompany me in the army."
1SAM|28|2|David said, "Then you will see for yourself what your servant can do." Achish replied, "Very well, I will make you my bodyguard for life."
1SAM|28|3|Now Samuel was dead, and all Israel had mourned for him and buried him in his own town of Ramah. Saul had expelled the mediums and spiritists from the land.
1SAM|28|4|The Philistines assembled and came and set up camp at Shunem, while Saul gathered all the Israelites and set up camp at Gilboa.
1SAM|28|5|When Saul saw the Philistine army, he was afraid; terror filled his heart.
1SAM|28|6|He inquired of the LORD, but the LORD did not answer him by dreams or Urim or prophets.
1SAM|28|7|Saul then said to his attendants, "Find me a woman who is a medium, so I may go and inquire of her.There is one in Endor," they said.
1SAM|28|8|So Saul disguised himself, putting on other clothes, and at night he and two men went to the woman. "Consult a spirit for me," he said, "and bring up for me the one I name."
1SAM|28|9|But the woman said to him, "Surely you know what Saul has done. He has cut off the mediums and spiritists from the land. Why have you set a trap for my life to bring about my death?"
1SAM|28|10|Saul swore to her by the LORD, "As surely as the LORD lives, you will not be punished for this."
1SAM|28|11|Then the woman asked, "Whom shall I bring up for you?Bring up Samuel," he said.
1SAM|28|12|When the woman saw Samuel, she cried out at the top of her voice and said to Saul, "Why have you deceived me? You are Saul!"
1SAM|28|13|The king said to her, "Don't be afraid. What do you see?" The woman said, "I see a spirit coming up out of the ground."
1SAM|28|14|"What does he look like?" he asked. "An old man wearing a robe is coming up," she said. Then Saul knew it was Samuel, and he bowed down and prostrated himself with his face to the ground.
1SAM|28|15|Samuel said to Saul, "Why have you disturbed me by bringing me up?I am in great distress," Saul said. "The Philistines are fighting against me, and God has turned away from me. He no longer answers me, either by prophets or by dreams. So I have called on you to tell me what to do."
1SAM|28|16|Samuel said, "Why do you consult me, now that the LORD has turned away from you and become your enemy?
1SAM|28|17|The LORD has done what he predicted through me. The LORD has torn the kingdom out of your hands and given it to one of your neighbors-to David.
1SAM|28|18|Because you did not obey the LORD or carry out his fierce wrath against the Amalekites, the LORD has done this to you today.
1SAM|28|19|The LORD will hand over both Israel and you to the Philistines, and tomorrow you and your sons will be with me. The LORD will also hand over the army of Israel to the Philistines."
1SAM|28|20|Immediately Saul fell full length on the ground, filled with fear because of Samuel's words. His strength was gone, for he had eaten nothing all that day and night.
1SAM|28|21|When the woman came to Saul and saw that he was greatly shaken, she said, "Look, your maidservant has obeyed you. I took my life in my hands and did what you told me to do.
1SAM|28|22|Now please listen to your servant and let me give you some food so you may eat and have the strength to go on your way."
1SAM|28|23|He refused and said, "I will not eat." But his men joined the woman in urging him, and he listened to them. He got up from the ground and sat on the couch.
1SAM|28|24|The woman had a fattened calf at the house, which she butchered at once. She took some flour, kneaded it and baked bread without yeast.
1SAM|28|25|Then she set it before Saul and his men, and they ate. That same night they got up and left.
1SAM|29|1|The Philistines gathered all their forces at Aphek, and Israel camped by the spring in Jezreel.
1SAM|29|2|As the Philistine rulers marched with their units of hundreds and thousands, David and his men were marching at the rear with Achish.
1SAM|29|3|The commanders of the Philistines asked, "What about these Hebrews?" Achish replied, "Is this not David, who was an officer of Saul king of Israel? He has already been with me for over a year, and from the day he left Saul until now, I have found no fault in him."
1SAM|29|4|But the Philistine commanders were angry with him and said, "Send the man back, that he may return to the place you assigned him. He must not go with us into battle, or he will turn against us during the fighting. How better could he regain his master's favor than by taking the heads of our own men?
1SAM|29|5|Isn't this the David they sang about in their dances: "'Saul has slain his thousands, and David his tens of thousands'?"
1SAM|29|6|So Achish called David and said to him, "As surely as the LORD lives, you have been reliable, and I would be pleased to have you serve with me in the army. From the day you came to me until now, I have found no fault in you, but the rulers don't approve of you.
1SAM|29|7|Turn back and go in peace; do nothing to displease the Philistine rulers."
1SAM|29|8|"But what have I done?" asked David. "What have you found against your servant from the day I came to you until now? Why can't I go and fight against the enemies of my lord the king?"
1SAM|29|9|Achish answered, "I know that you have been as pleasing in my eyes as an angel of God; nevertheless, the Philistine commanders have said, 'He must not go up with us into battle.'
1SAM|29|10|Now get up early, along with your master's servants who have come with you, and leave in the morning as soon as it is light."
1SAM|29|11|So David and his men got up early in the morning to go back to the land of the Philistines, and the Philistines went up to Jezreel.
1SAM|30|1|David and his men reached Ziklag on the third day. Now the Amalekites had raided the Negev and Ziklag. They had attacked Ziklag and burned it,
1SAM|30|2|and had taken captive the women and all who were in it, both young and old. They killed none of them, but carried them off as they went on their way.
1SAM|30|3|When David and his men came to Ziklag, they found it destroyed by fire and their wives and sons and daughters taken captive.
1SAM|30|4|So David and his men wept aloud until they had no strength left to weep.
1SAM|30|5|David's two wives had been captured-Ahinoam of Jezreel and Abigail, the widow of Nabal of Carmel.
1SAM|30|6|David was greatly distressed because the men were talking of stoning him; each one was bitter in spirit because of his sons and daughters. But David found strength in the LORD his God.
1SAM|30|7|Then David said to Abiathar the priest, the son of Ahimelech, "Bring me the ephod." Abiathar brought it to him,
1SAM|30|8|and David inquired of the LORD, "Shall I pursue this raiding party? Will I overtake them?Pursue them," he answered. "You will certainly overtake them and succeed in the rescue."
1SAM|30|9|David and the six hundred men with him came to the Besor Ravine, where some stayed behind,
1SAM|30|10|for two hundred men were too exhausted to cross the ravine. But David and four hundred men continued the pursuit.
1SAM|30|11|They found an Egyptian in a field and brought him to David. They gave him water to drink and food to eat-
1SAM|30|12|part of a cake of pressed figs and two cakes of raisins. He ate and was revived, for he had not eaten any food or drunk any water for three days and three nights.
1SAM|30|13|David asked him, "To whom do you belong, and where do you come from?" He said, "I am an Egyptian, the slave of an Amalekite. My master abandoned me when I became ill three days ago.
1SAM|30|14|We raided the Negev of the Kerethites and the territory belonging to Judah and the Negev of Caleb. And we burned Ziklag."
1SAM|30|15|David asked him, "Can you lead me down to this raiding party?" He answered, "Swear to me before God that you will not kill me or hand me over to my master, and I will take you down to them."
1SAM|30|16|He led David down, and there they were, scattered over the countryside, eating, drinking and reveling because of the great amount of plunder they had taken from the land of the Philistines and from Judah.
1SAM|30|17|David fought them from dusk until the evening of the next day, and none of them got away, except four hundred young men who rode off on camels and fled.
1SAM|30|18|David recovered everything the Amalekites had taken, including his two wives.
1SAM|30|19|Nothing was missing: young or old, boy or girl, plunder or anything else they had taken. David brought everything back.
1SAM|30|20|He took all the flocks and herds, and his men drove them ahead of the other livestock, saying, "This is David's plunder."
1SAM|30|21|Then David came to the two hundred men who had been too exhausted to follow him and who were left behind at the Besor Ravine. They came out to meet David and the people with him. As David and his men approached, he greeted them.
1SAM|30|22|But all the evil men and troublemakers among David's followers said, "Because they did not go out with us, we will not share with them the plunder we recovered. However, each man may take his wife and children and go."
1SAM|30|23|David replied, "No, my brothers, you must not do that with what the LORD has given us. He has protected us and handed over to us the forces that came against us.
1SAM|30|24|Who will listen to what you say? The share of the man who stayed with the supplies is to be the same as that of him who went down to the battle. All will share alike."
1SAM|30|25|David made this a statute and ordinance for Israel from that day to this.
1SAM|30|26|When David arrived in Ziklag, he sent some of the plunder to the elders of Judah, who were his friends, saying, "Here is a present for you from the plunder of the LORD's enemies."
1SAM|30|27|He sent it to those who were in Bethel, Ramoth Negev and Jattir;
1SAM|30|28|to those in Aroer, Siphmoth, Eshtemoa
1SAM|30|29|and Racal; to those in the towns of the Jerahmeelites and the Kenites;
1SAM|30|30|to those in Hormah, Bor Ashan, Athach
1SAM|30|31|and Hebron; and to those in all the other places where David and his men had roamed.
1SAM|31|1|Now the Philistines fought against Israel; the Israelites fled before them, and many fell slain on Mount Gilboa.
1SAM|31|2|The Philistines pressed hard after Saul and his sons, and they killed his sons Jonathan, Abinadab and Malki-Shua.
1SAM|31|3|The fighting grew fierce around Saul, and when the archers overtook him, they wounded him critically.
1SAM|31|4|Saul said to his armor-bearer, "Draw your sword and run me through, or these uncircumcised fellows will come and run me through and abuse me." But his armor-bearer was terrified and would not do it; so Saul took his own sword and fell on it.
1SAM|31|5|When the armor-bearer saw that Saul was dead, he too fell on his sword and died with him.
1SAM|31|6|So Saul and his three sons and his armor-bearer and all his men died together that same day.
1SAM|31|7|When the Israelites along the valley and those across the Jordan saw that the Israelite army had fled and that Saul and his sons had died, they abandoned their towns and fled. And the Philistines came and occupied them.
1SAM|31|8|The next day, when the Philistines came to strip the dead, they found Saul and his three sons fallen on Mount Gilboa.
1SAM|31|9|They cut off his head and stripped off his armor, and they sent messengers throughout the land of the Philistines to proclaim the news in the temple of their idols and among their people.
1SAM|31|10|They put his armor in the temple of the Ashtoreths and fastened his body to the wall of Beth Shan.
1SAM|31|11|When the people of Jabesh Gilead heard of what the Philistines had done to Saul,
1SAM|31|12|all their valiant men journeyed through the night to Beth Shan. They took down the bodies of Saul and his sons from the wall of Beth Shan and went to Jabesh, where they burned them.
1SAM|31|13|Then they took their bones and buried them under a tamarisk tree at Jabesh, and they fasted seven days.
