2KGS|1|1|И отложился Моав от Израиля по смерти Ахава.
2KGS|1|2|Охозия же упал чрез решетку с горницы своей, что в Самарии, и занемог. И послал послов, и сказал им: пойдите, спросите у Веельзевула, божества Аккаронского: выздоровею ли я от сей болезни?
2KGS|1|3|Тогда Ангел Господень сказал Илии Фесвитянину: встань, пойди навстречу посланным от царя Самарийского и скажи им: разве нет Бога в Израиле, что вы идете вопрошать Веельзевула, божество Аккаронское?
2KGS|1|4|За это так говорит Господь: с постели, на которую ты лег, не сойдешь с нее, но умрешь. И пошел Илия.
2KGS|1|5|И возвратились к [Охозии] посланные. И он сказал им: что это вы возвратились?
2KGS|1|6|И сказали ему: навстречу нам вышел человек и сказал нам: пойдите, возвратитесь к царю, который послал вас, и скажите ему: так говорит Господь: разве нет Бога в Израиле, что ты посылаешь вопрошать Веельзевула, божество Аккаронское? За то с постели, на которую ты лег, не сойдешь с нее, но умрешь.
2KGS|1|7|И сказал им: каков видом тот человек, который вышел навстречу вам и говорил вам слова сии?
2KGS|1|8|Они сказали ему: человек тот весь в волосах и кожаным поясом подпоясан по чреслам своим. И сказал он: это Илия Фесвитянин.
2KGS|1|9|И послал к нему пятидесятника с его пятидесятком. И он взошел к нему, когда Илия сидел на верху горы, и сказал ему: человек Божий! царь говорит: сойди.
2KGS|1|10|И отвечал Илия, и сказал пятидесятнику: если я человек Божий, то пусть сойдет огонь с неба и попалит тебя и твой пятидесяток. И сошел огонь с неба и попалил его и пятидесяток его.
2KGS|1|11|И послал к нему царь другого пятидесятника с его пятидесятком. И он стал говорить ему: человек Божий! так сказал царь: сойди скорее.
2KGS|1|12|И отвечал Илия и сказал ему: если я человек Божий, то пусть сойдет огонь с неба и попалит тебя и твой пятидесяток. И сошел огонь Божий с неба, и попалил его и пятидесяток его.
2KGS|1|13|И еще послал в третий раз пятидесятника с его пятидесятком. И поднялся, и пришел пятидесятник третий, и пал на колена свои пред Илиею, и умолял его, и говорил ему: человек Божий! да не будет презрена душа моя и душа рабов твоих – сих пятидесяти – пред очами твоими;
2KGS|1|14|вот, сошел огонь с неба, и попалил двух пятидесятников прежних с их пятидесятками; но теперь да не будет презрена душа моя пред очами твоими!
2KGS|1|15|И сказал Ангел Господень Илии: пойди с ним, не бойся его. И он встал, и пошел с ним к царю.
2KGS|1|16|И сказал ему: так говорит Господь: за то, что ты посылал послов вопрошать Веельзевула, божество Аккаронское, как будто в Израиле нет Бога, чтобы вопрошать о слове Его, – с постели, на которую ты лег, не сойдешь с нее, но умрешь.
2KGS|1|17|И умер он по слову Господню, которое изрек Илия. И воцарился Иорам вместо него, во второй год Иорама, сына Иосафатова, царя Иудейского, так как сына у того не было.
2KGS|1|18|Прочее об Охозии, что он сделал, написано в летописи царей Израильских.
2KGS|2|1|В то время, как Господь восхотел вознести Илию в вихре на небо, шел Илия с Елисеем из Галгала.
2KGS|2|2|И сказал Илия Елисею: останься здесь, ибо Господь посылает меня в Вефиль. Но Елисей сказал: жив Господь и жива душа твоя! не оставлю тебя. И пошли они в Вефиль.
2KGS|2|3|И вышли сыны пророков, которые в Вефиле, к Елисею и сказали ему: знаешь ли, что сегодня Господь вознесет господина твоего над главою твоею? Он сказал: я также знаю, молчите.
2KGS|2|4|И сказал ему Илия: Елисей, останься здесь, ибо Господь посылает меня в Иерихон. И сказал он: жив Господь и жива душа твоя! не оставлю тебя. И пришли в Иерихон.
2KGS|2|5|И подошли сыны пророков, которые в Иерихоне, к Елисею и сказали ему: знаешь ли, что сегодня Господь берет господина твоего и вознесет над главою твоею? Он сказал: я также знаю, молчите.
2KGS|2|6|И сказал ему Илия: останься здесь, ибо Господь посылает меня к Иордану. И сказал он: жив Господь и жива душа твоя! не оставлю тебя. И пошли оба.
2KGS|2|7|Пятьдесят человек из сынов пророческих пошли и стали вдали напротив их, а они оба стояли у Иордана.
2KGS|2|8|И взял Илия милоть свою, и свернул, и ударил ею по воде, и расступилась она туда и сюда, и перешли оба посуху.
2KGS|2|9|Когда они перешли, Илия сказал Елисею: проси, что сделать тебе, прежде нежели я буду взят от тебя. И сказал Елисей: дух, который в тебе, пусть будет на мне вдвойне.
2KGS|2|10|И сказал он: трудного ты просишь. Если увидишь, как я буду взят от тебя, то будет тебе так, а если не увидишь, не будет.
2KGS|2|11|Когда они шли и дорогою разговаривали, вдруг явилась колесница огненная и кони огненные, и разлучили их обоих, и понесся Илия в вихре на небо.
2KGS|2|12|Елисей же смотрел и воскликнул: отец мой, отец мой, колесница Израиля и конница его! И не видел его более. И схватил он одежды свои и разодрал их на две части.
2KGS|2|13|И поднял милоть Илии, упавшую с него, и пошел назад, и стал на берегу Иордана;
2KGS|2|14|и взял милоть Илии, упавшую с него, и ударил ею по воде, и сказал: где Господь, Бог Илии, – Он Самый? И ударил по воде, и она расступилась туда и сюда, и перешел Елисей.
2KGS|2|15|И увидели его сыны пророков, которые в Иерихоне, издали, и сказали: опочил дух Илии на Елисее. И пошли навстречу ему, и поклонились ему до земли,
2KGS|2|16|и сказали ему: вот, есть [у нас], рабов твоих, человек пятьдесят, люди сильные; пусть бы они пошли и поискали господина твоего; может быть, унес его Дух Господень и поверг его на одной из гор, или на одной из долин. Он же сказал: не посылайте.
2KGS|2|17|Но они приступали к нему долго, так что наскучили ему, и он сказал: пошлите. И послали пятьдесят человек, и искали три дня, и не нашли его,
2KGS|2|18|и возвратились к нему, между тем как он оставался в Иерихоне, и сказал им: не говорил ли я вам: не ходите?
2KGS|2|19|И сказали жители того города Елисею: вот, положение этого города хорошо, как видит господин мой; но вода нехороша и земля бесплодна.
2KGS|2|20|И сказал он: дайте мне новую чашу и положите туда соли. И дали ему.
2KGS|2|21|И вышел он к истоку воды, и бросил туда соли, и сказал: так говорит Господь: Я сделал воду сию здоровою, не будет от нее впредь ни смерти, ни бесплодия.
2KGS|2|22|И вода стала здоровою до сего дня, по слову Елисея, которое он сказал.
2KGS|2|23|И пошел он оттуда в Вефиль. Когда он шел дорогою, малые дети вышли из города и насмехались над ним и говорили ему: иди, плешивый! иди, плешивый!
2KGS|2|24|Он оглянулся и увидел их и проклял их именем Господним. И вышли две медведицы из леса и растерзали из них сорок два ребенка.
2KGS|2|25|Отсюда пошел он на гору Кармил, а оттуда возвратился в Самарию.
2KGS|3|1|Иорам, сын Ахава, воцарился над Израилем в Самарии в восемнадцатый год Иосафата, царя Иудейского, и царствовал двенадцать лет,
2KGS|3|2|и делал неугодное в очах Господних, хотя не так, как отец его и мать его: он снял статую Ваала, которую сделал отец его;
2KGS|3|3|однако же грехов Иеровоама, сына Наватова, который ввел в грех Израиля, он держался, не отставал от них.
2KGS|3|4|Меса, царь Моавитский, был богат скотом и присылал царю Израильскому по сто тысяч овец и по сто тысяч неостриженных баранов.
2KGS|3|5|Но когда умер Ахав, царь Моавитский отложился от царя Израильского.
2KGS|3|6|И выступил царь Иорам в то время из Самарии и сделал смотр всем Израильтянам;
2KGS|3|7|и пошел и послал к Иосафату, царю Иудейскому, сказать: царь Моавитский отложился от меня, пойдешь ли со мной на войну против Моава? Он сказал: пойду; как ты, так и я, как твой народ, так и мой народ; как твои кони, так и мои кони.
2KGS|3|8|И сказал: какою дорогою идти нам? Он сказал: дорогою пустыни Едомской.
2KGS|3|9|И пошел царь Израильский, и царь Иудейский, и царь Едомский, и шли они обходом семь дней, и не было воды для войска и для скота, который [шел] за ними.
2KGS|3|10|И сказал царь Израильский: ах! созвал Господь трех царей сих, чтобы предать их в руку Моава.
2KGS|3|11|И сказал Иосафат: нет ли здесь пророка Господня, чтобы нам вопросить Господа чрез него? И отвечал один из слуг царя Израильского и сказал: здесь Елисей, сын Сафатов, который подавал воду на руки Илии.
2KGS|3|12|И сказал Иосафат: есть у него слово Господне. И пошли к нему царь Израильский, и Иосафат, и царь Едомский.
2KGS|3|13|И сказал Елисей царю Израильскому: что мне и тебе? пойди к пророкам отца твоего и к пророкам матери твоей. И сказал ему царь Израильский: нет, потому что Господь созвал сюда трех царей сих, чтобы предать их в руку Моава.
2KGS|3|14|И сказал Елисей: жив Господь Саваоф, пред Которым я стою! Если бы я не почитал Иосафата, царя Иудейского, то не взглянул бы на тебя и не видел бы тебя;
2KGS|3|15|теперь позовите мне гуслиста. И когда гуслист играл на гуслях, тогда рука Господня коснулась Елисея,
2KGS|3|16|и он сказал: так говорит Господь: делайте на сей долине рвы за рвами,
2KGS|3|17|ибо так говорит Господь: не увидите ветра и не увидите дождя, а долина сия наполнится водою, которую будете пить вы и мелкий и крупный скот ваш;
2KGS|3|18|но этого мало пред очами Господа; Он и Моава предаст в руки ваши,
2KGS|3|19|и вы поразите все города укрепленные и все города главные, и все лучшие деревья срубите, и все источники водные запрудите, и все лучшие участки полевые испортите каменьями.
2KGS|3|20|Поутру, когда возносят хлебное приношение, вдруг полилась вода по пути от Едома, и наполнилась земля водою.
2KGS|3|21|Когда Моавитяне услышали, что идут цари воевать с ними, тогда собраны были все, начиная от носящего пояс и старше, и стали на границе.
2KGS|3|22|Поутру встали они рано, и когда солнце воссияло над водою, Моавитянам издали показалась эта вода красною, как кровь.
2KGS|3|23|И сказали они: это кровь; сразились цари между собою и истребили друг друга; теперь на добычу, Моав!
2KGS|3|24|И пришли они к стану Израильскому. И встали Израильтяне и стали бить Моавитян, и те побежали от них, а они продолжали идти на них и бить Моавитян.
2KGS|3|25|И города разрушили, и на всякий лучший участок в поле бросили каждый по камню и закидали его; и все протоки вод запрудили и все дерева лучшие срубили, так что оставались только каменья в Кир–Харешете. И обступили его пращники и разрушили его.
2KGS|3|26|И увидел царь Моавитский, что битва одолевает его, и взял с собою семьсот человек, владеющих мечом, чтобы пробиться к царю Едомскому; но не могли.
2KGS|3|27|И взял он сына своего первенца, которому следовало царствовать вместо него, и вознес его во всесожжение на стене. Это произвело большое негодование в Израильтянах, и они отступили от него и возвратились в свою землю.
2KGS|4|1|Одна из жен сынов пророческих с воплем говорила Елисею: раб твой, мой муж, умер; а ты знаешь, что раб твой боялся Господа; теперь пришел заимодавец взять обоих детей моих в рабы себе.
2KGS|4|2|И сказал ей Елисей: что мне сделать тебе? скажи мне, что есть у тебя в доме? Она сказала: нет у рабы твоей ничего в доме, кроме сосуда с елеем.
2KGS|4|3|И сказал он: пойди, попроси себе сосудов на стороне, у всех соседей твоих, сосудов порожних; набери немало,
2KGS|4|4|и пойди, запри дверь за собою и за сыновьями твоими, и наливай во все эти сосуды; полные отставляй.
2KGS|4|5|И пошла от него и заперла дверь за собой и за сыновьями своими. Они подавали ей, а она наливала.
2KGS|4|6|Когда наполнены были сосуды, она сказала сыну своему: подай мне еще сосуд. Он сказал ей: нет более сосудов. И остановилось масло.
2KGS|4|7|И пришла она, и пересказала человеку Божию. Он сказал: пойди, продай масло и заплати долги твои; а что останется, тем будешь жить с сыновьями твоими.
2KGS|4|8|В один день пришел Елисей в Сонам. Там одна богатая женщина упросила его [к себе] есть хлеба; и когда он ни проходил, всегда заходил туда есть хлеба.
2KGS|4|9|И сказала она мужу своему: вот, я знаю, что человек Божий, который проходит мимо нас постоянно, святой;
2KGS|4|10|сделаем небольшую горницу над стеною и поставим ему там постель, и стол, и седалище, и светильник; и когда он будет приходить к нам, пусть заходит туда.
2KGS|4|11|В один день он пришел туда, и зашел в горницу, и лег там,
2KGS|4|12|и сказал Гиезию, слуге своему: позови эту Сонамитянку. И позвал ее, и она стала пред ним.
2KGS|4|13|И сказал ему: скажи ей: "вот, ты так заботишься о нас; что сделать бы тебе? не нужно ли поговорить о тебе с царем, или с военачальником?" Она сказала: нет, среди своего народа я живу.
2KGS|4|14|И сказал он: что же сделать ей? И сказал Гиезий: да вот, сына нет у нее, а муж ее стар.
2KGS|4|15|И сказал он: позови ее. Он позвал ее, и стала она в дверях.
2KGS|4|16|И сказал он: через год, в это самое время ты будешь держать на руках сына. И сказала она: нет, господин мой, человек Божий, не обманывай рабы твоей.
2KGS|4|17|И женщина стала беременною и родила сына на другой год, в то самое время, как сказал ей Елисей.
2KGS|4|18|И подрос ребенок и в один день пошел к отцу своему, к жнецам.
2KGS|4|19|И сказал отцу своему: голова моя! голова моя болит! И сказал тот слуге своему: отнеси его к матери его.
2KGS|4|20|И понес его и принес его к матери его. И он сидел на коленях у нее до полудня, и умер.
2KGS|4|21|И пошла она, и положила его на постели человека Божия, и заперла его, и вышла,
2KGS|4|22|и позвала мужа своего и сказала: пришли мне одного из слуг и одну из ослиц, я поеду к человеку Божию и возвращусь.
2KGS|4|23|Он сказал: зачем тебе ехать к нему? сегодня не новомесячие и не суббота. Но она сказала: хорошо.
2KGS|4|24|И оседлала ослицу и сказала слуге своему: веди и иди; не останавливайся, доколе не скажу тебе.
2KGS|4|25|И отправилась и прибыла к человеку Божию, к горе Кармил. И когда увидел человек Божий ее издали, то сказал слуге своему Гиезию: это та Сонамитянка.
2KGS|4|26|Побеги к ней навстречу и скажи ей: "здорова ли ты? здоров ли муж твой? здоров ли ребенок?" – Она сказала: здоровы.
2KGS|4|27|Когда же пришла к человеку Божию на гору, ухватилась за ноги его. И подошел Гиезий, чтобы отвести ее; но человек Божий сказал: оставь ее, душа у нее огорчена, а Господь скрыл от меня и не объявил мне.
2KGS|4|28|И сказала она: просила ли я сына у господина моего? не говорила ли я: "не обманывай меня"?
2KGS|4|29|И сказал он Гиезию: опояшь чресла твои и возьми жезл мой в руку твою, и пойди; если встретишь кого, не приветствуй его, и если кто будет тебя приветствовать, не отвечай ему; и положи посох мой на лице ребенка.
2KGS|4|30|И сказала мать ребенка: жив Господь и жива душа твоя! не отстану от тебя. И он встал и пошел за нею.
2KGS|4|31|Гиезий пошел впереди их и положил жезл на лице ребенка. Но не было ни голоса, ни ответа. И вышел навстречу ему, и донес ему, и сказал: не пробуждается ребенок.
2KGS|4|32|И вошел Елисей в дом, и вот, ребенок умерший лежит на постели его.
2KGS|4|33|И вошел, и запер дверь за собою, и помолился Господу.
2KGS|4|34|И поднялся и лег над ребенком, и приложил свои уста к его устам, и свои глаза к его глазам, и свои ладони к его ладоням, и простерся на нем, и согрелось тело ребенка.
2KGS|4|35|И встал и прошел по горнице взад и вперед; потом опять поднялся и простерся на нем. И чихнул ребенок раз семь, и открыл ребенок глаза свои.
2KGS|4|36|И позвал он Гиезия и сказал: позови эту Сонамитянку. И тот позвал ее. Она пришла к нему, и он сказал: возьми сына твоего.
2KGS|4|37|И подошла, и упала ему в ноги, и поклонилась до земли; и взяла сына своего и пошла.
2KGS|4|38|Елисей же возвратился в Галгал. И был голод в земле той, и сыны пророков сидели пред ним. И сказал он слуге своему: поставь большой котел и свари похлебку для сынов пророческих.
2KGS|4|39|И вышел один из них в поле собирать овощи, и нашел дикое вьющееся растение, и набрал с него диких плодов полную одежду свою; и пришел и накрошил их в котел с похлебкою, так как они не знали [их].
2KGS|4|40|И налили им есть. Но как скоро они стали есть похлебку, то подняли крик и говорили: смерть в котле, человек Божий! И не могли есть.
2KGS|4|41|И сказал он: подайте муки. И всыпал ее в котел и сказал [Гиезию]: наливай людям, пусть едят. И не стало ничего вредного в котле.
2KGS|4|42|Пришел некто из Ваал–Шалиши, и принес человеку Божию хлебный начаток – двадцать ячменных хлебцев и сырые зерна в шелухе. И сказал Елисей: отдай людям, пусть едят.
2KGS|4|43|И сказал слуга его: что тут я дам ста человекам? И сказал он: отдай людям, пусть едят, ибо так говорит Господь: "насытятся, и останется".
2KGS|4|44|Он подал им, и они насытились, и еще осталось, по слову Господню.
2KGS|5|1|Нееман, военачальник царя Сирийского, был великий человек у господина своего и уважаемый, потому что чрез него дал Господь победу Сириянам; и человек сей был отличный воин, но прокаженный.
2KGS|5|2|Сирияне [однажды] пошли отрядами и взяли в плен из земли Израильской маленькую девочку, и она служила жене Неемановой.
2KGS|5|3|И сказала она госпоже своей: о, если бы господин мой побывал у пророка, который в Самарии, то он снял бы с него проказу его!
2KGS|5|4|И пошел [Нееман] и передал это господину своему, говоря: так и так говорит девочка, которая из земли Израильской.
2KGS|5|5|И сказал царь Сирийский [Нееману]: пойди, сходи, а я пошлю письмо к царю Израильскому. Он пошел и взял с собою десять талантов серебра и шесть тысяч [сиклей] золота, и десять перемен одежд;
2KGS|5|6|и принес письмо царю Израильскому, в котором было сказано: вместе с письмом сим, вот, я посылаю к тебе Неемана, слугу моего, чтобы ты снял с него проказу его.
2KGS|5|7|Царь Израильский, прочитав письмо, разодрал одежды свои и сказал: разве я Бог, чтобы умерщвлять и оживлять, что он посылает ко мне, чтобы я снял с человека проказу его? вот, теперь знайте и смотрите, что он ищет предлога враждовать против меня.
2KGS|5|8|Когда услышал Елисей, человек Божий, что царь Израильский разодрал одежды свои, то послал сказать царю: для чего ты разодрал одежды свои? пусть он придет ко мне, и узнает, что есть пророк в Израиле.
2KGS|5|9|И прибыл Нееман на конях своих и на колеснице своей, и остановился у входа в дом Елисеев.
2KGS|5|10|И выслал к нему Елисей слугу сказать: пойди, омойся семь раз в Иордане, и обновится тело твое у тебя, и будешь чист.
2KGS|5|11|И разгневался Нееман, и пошел, и сказал: вот, я думал, что он выйдет, станет и призовет имя Господа Бога своего, и возложит руку свою на то место и снимет проказу;
2KGS|5|12|разве Авана и Фарфар, реки Дамасские, не лучше всех вод Израильских? разве я не мог бы омыться в них и очиститься? И оборотился и удалился в гневе.
2KGS|5|13|И подошли рабы его и говорили ему, и сказали: отец мой, [если] [бы] что–нибудь важное сказал тебе пророк, то не сделал ли бы ты? а тем более, когда он сказал тебе только: "омойся, и будешь чист".
2KGS|5|14|И пошел он и окунулся в Иордане семь раз, по слову человека Божия, и обновилось тело его, как тело малого ребенка, и очистился.
2KGS|5|15|И возвратился к человеку Божию он и все сопровождавшие его, и пришел, и стал пред ним, и сказал: вот, я узнал, что на всей земле нет Бога, как только у Израиля; итак прими дар от раба твоего.
2KGS|5|16|И сказал он: жив Господь, пред лицем Которого стою! не приму. И тот принуждал его взять, но он не согласился.
2KGS|5|17|И сказал Нееман: если уже не так, то пусть рабу твоему дадут земли, сколько снесут два лошака, потому что не будет впредь раб твой приносить всесожжения и жертвы другим богам, кроме Господа;
2KGS|5|18|только вот в чем да простит Господь раба твоего: когда пойдет господин мой в дом Риммона для поклонения там и опрется на руку мою, и поклонюсь я в доме Риммона, то, за мое поклонение в доме Риммона, да простит Господь раба твоего в случае сем.
2KGS|5|19|И сказал ему: иди с миром. И он отъехал от него на небольшое пространство земли.
2KGS|5|20|И сказал Гиезий, слуга Елисея, человека Божия: вот, господин мой отказался взять из руки Неемана, этого Сириянина, то, что он приносил. Жив Господь! Побегу я за ним, и возьму у него что–нибудь.
2KGS|5|21|И погнался Гиезий за Нееманом. И увидел Нееман бегущего за собою, и сошел с колесницы навстречу ему, и сказал: с миром ли?
2KGS|5|22|Он отвечал: с миром; господин мой послал меня сказать: "вот, теперь пришли ко мне с горы Ефремовой два молодых человека из сынов пророческих; дай им талант серебра и две перемены одежд".
2KGS|5|23|И сказал Нееман: возьми, пожалуй, два таланта. И упрашивал его. И завязал он два таланта серебра в два мешка и две перемены одежд и отдал двум слугам своим, и понесли перед ним.
2KGS|5|24|Когда он пришел к холму, то взял из рук их и спрятал дома. И отпустил людей, и они ушли.
2KGS|5|25|Когда он пришел и явился к господину своему, Елисей сказал ему: откуда, Гиезий? И сказал он: никуда не ходил раб твой.
2KGS|5|26|И сказал он ему: разве сердце мое не сопутствовало тебе, когда обратился навстречу тебе человек тот с колесницы своей? время ли брать серебро и брать одежды, или масличные деревья и виноградники, и мелкий или крупный скот, и рабов или рабынь?
2KGS|5|27|Пусть же проказа Нееманова пристанет к тебе и к потомству твоему навек. И вышел он от него [белый] от проказы, как снег.
2KGS|6|1|И сказали сыны пророков Елисею: вот, место, где мы живем при тебе, тесно для нас;
2KGS|6|2|пойдем к Иордану и возьмем оттуда каждый по одному бревну и сделаем себе там место для жительства. Он сказал: пойдите.
2KGS|6|3|И сказал один: сделай милость, пойди и ты с рабами твоими. И сказал он: пойду.
2KGS|6|4|И пошел с ними, и пришли к Иордану и стали рубить деревья.
2KGS|6|5|И когда один валил бревно, топор его упал в воду. И закричал он и сказал: ах, господин мой! а он взят был на подержание!
2KGS|6|6|И сказал человек Божий: где он упал? Он указал ему место. И отрубил он [кусок] дерева и бросил туда, и всплыл топор.
2KGS|6|7|И сказал он: возьми себе. Он протянул руку свою и взял его.
2KGS|6|8|Царь Сирийский пошел войною на Израильтян, и советовался со слугами своими, говоря: в таком–то и в таком–то месте я расположу свой стан.
2KGS|6|9|И посылал человек Божий к царю Израильскому сказать: берегись проходить сим местом, ибо там Сирияне залегли.
2KGS|6|10|И посылал царь Израильский на то место, о котором говорил ему человек Божий и предостерегал его; и сберег себя там не раз и не два.
2KGS|6|11|И встревожилось сердце царя Сирийского по сему случаю, и призвал он рабов своих и сказал им: скажите мне, кто из наших [в сношении] с царем Израильским?
2KGS|6|12|И сказал один из слуг его: никто, господин мой царь; а Елисей пророк, который у Израиля, пересказывает царю Израильскому и те слова, которые ты говоришь в спальной комнате твоей.
2KGS|6|13|И сказал он: пойдите, узнайте, где он; я пошлю и возьму его. И донесли ему и сказали: вот, он в Дофаиме.
2KGS|6|14|И послал туда коней и колесницы и много войска. И пришли ночью и окружили город.
2KGS|6|15|Поутру служитель человека Божия встал и вышел; и вот, войско вокруг города, и кони и колесницы. И сказал ему слуга его: увы! господин мой, что нам делать?
2KGS|6|16|И сказал он: не бойся, потому что тех, которые с нами, больше, нежели тех, которые с ними.
2KGS|6|17|И молился Елисей, и говорил: Господи! открой ему глаза, чтоб он увидел. И открыл Господь глаза слуге, и он увидел, и вот, вся гора наполнена конями и колесницами огненными кругом Елисея.
2KGS|6|18|Когда пошли к нему Сирияне, Елисей помолился Господу и сказал: порази их слепотою. И Он поразил их слепотою по слову Елисея.
2KGS|6|19|И сказал им Елисей: это не та дорога и не тот город; идите за мною, и я провожу вас к тому человеку, которого вы ищете. И привел их в Самарию.
2KGS|6|20|Когда они пришли в Самарию, Елисей сказал: Господи! открой глаза им, чтобы они видели. И открыл Господь глаза их, и увидели, что они в средине Самарии.
2KGS|6|21|И сказал царь Израильский Елисею, увидев их: не избить ли их, отец мой?
2KGS|6|22|И сказал он: не убивай. Разве мечом твоим и луком твоим ты пленил их, чтобы убивать их? Предложи им хлеба и воды; пусть едят и пьют, и пойдут к государю своему.
2KGS|6|23|И приготовил им большой обед, и они ели и пили. И отпустил их, и пошли к государю своему. И не ходили более те полчища Сирийские в землю Израилеву.
2KGS|6|24|После того собрал Венадад, царь Сирийский, все войско свое и выступил, и осадил Самарию.
2KGS|6|25|И был большой голод в Самарии, когда они осадили ее, так что ослиная голова продавалась по восьмидесяти сиклей серебра, и четвертая часть каба голубиного помета – по пяти сиклей серебра.
2KGS|6|26|Однажды царь Израильский проходил по стене, и женщина с воплем говорила ему: помоги, господин мой царь.
2KGS|6|27|И сказал он: если не поможет тебе Господь, из чего я помогу тебе? с гумна ли, с точила ли?
2KGS|6|28|И сказал ей царь: что тебе? И сказала она: эта женщина говорила мне: "отдай своего сына, съедим его сегодня, а сына моего съедим завтра".
2KGS|6|29|И сварили мы моего сына, и съели его. И я сказала ей на другой день: "отдай же твоего сына, и съедим его". Но она спрятала своего сына.
2KGS|6|30|Царь, выслушав слова женщины, разодрал одежды свои; и проходил он по стене, и народ видел, что вретище на самом теле его.
2KGS|6|31|И сказал: пусть то и то сделает мне Бог, и еще более сделает, если останется голова Елисея, сына Сафатова, на нем сегодня.
2KGS|6|32|Елисей же сидел в своем доме, и старцы сидели у него. И послал [царь] человека от себя. Прежде нежели пришел посланный к нему, он сказал старцам: видите ли, что этот сын убийцы послал снять с меня голову? Смотрите, когда придет посланный, затворите дверь и прижмите его дверью. А вот и топот ног господина его за ним!
2KGS|6|33|Еще говорил он с ними, и вот посланный приходит к нему, и сказал: вот какое бедствие от Господа! чего мне впредь ждать от Господа?
2KGS|7|1|И сказал Елисей: выслушайте слово Господне: так говорит Господь: завтра в это время мера муки лучшей [будет] по сиклю и две меры ячменя по сиклю у ворот Самарии.
2KGS|7|2|И отвечал сановник, на руку которого царь опирался, человеку Божию, и сказал: если бы Господь и открыл окна на небе, и тогда может ли это быть? И сказал тот: вот увидишь глазами твоими, но есть этого не будешь.
2KGS|7|3|Четыре человека прокаженных находились при входе в ворота и говорили они друг другу: что нам сидеть здесь, ожидая смерти?
2KGS|7|4|Если решиться нам пойти в город, то в городе голод, и мы там умрем; если же сидеть здесь, то также умрем. Пойдем лучше в стан Сирийский. Если оставят нас в живых, будем жить, а если умертвят, умрем.
2KGS|7|5|И встали в сумерки, чтобы пойти в стан Сирийский. И пришли к краю стана Сирийского, и вот, нет там ни одного человека.
2KGS|7|6|Господь сделал то, что стану Сирийскому послышался стук колесниц и ржание коней, шум войска большого. И сказали они друг другу: верно нанял против нас царь Израильский царей Хеттейских и Египетских, чтобы пойти на нас.
2KGS|7|7|И встали и побежали в сумерки, и оставили шатры свои, и коней своих, и ослов своих, весь стан, как он был, и побежали, спасая себя.
2KGS|7|8|И пришли те прокаженные к краю стана, и вошли в один шатер, и ели и пили, и взяли оттуда серебро, и золото, и одежды, и пошли и спрятали. Пошли еще в другой шатер, и там взяли, и пошли и спрятали.
2KGS|7|9|И сказали друг другу: не так мы делаем. День сей – день радостной вести, если мы замедлим и будем дожидаться утреннего света, то падет на нас вина. Пойдем же и уведомим дом царский.
2KGS|7|10|И пришли, и позвали привратников городских, и рассказали им, говоря: мы ходили в стан Сирийский, и вот, нет там ни человека, ни голоса человеческого, а только кони привязанные, и ослы привязанные, и шатры, как быть им.
2KGS|7|11|И позвали привратников, и они передали весть в самый дворец царский.
2KGS|7|12|И встал царь ночью, и сказал слугам своим: скажу вам, что делают с нами Сирияне. Они знают, что мы терпим голод, и вышли из стана, чтобы спрятаться в поле, думая так: "когда они выйдут из города, мы захватим их живыми и вторгнемся в город".
2KGS|7|13|И отвечал один из служащих при нем, и сказал: пусть возьмут пять из остальных коней, которые остались в городе, (из всего ополчения Израильтян только и осталось в нем, из всего ополчения Израильтян, которое погибло), и пошлем, и посмотрим.
2KGS|7|14|И взяли две пары коней, запряженных в колесницы. И послал царь вслед Сирийского войска, сказав: пойдите, посмотрите.
2KGS|7|15|И ехали за ним до Иордана, и вот вся дорога устлана одеждами и вещами, которые побросали Сирияне при торопливом побеге своем. И возвратились посланные, и донесли царю.
2KGS|7|16|И вышел народ, и разграбил стан Сирийский, и была мера муки лучшей по сиклю, и две меры ячменя по сиклю, по слову Господню.
2KGS|7|17|И царь поставил того сановника, на руку которого опирался, у ворот; и растоптал его народ в воротах, и он умер, как сказал человек Божий, который говорил, когда приходил к нему царь.
2KGS|7|18|Когда говорил человек Божий царю так: "две меры ячменя по сиклю, и мера муки лучшей по сиклю будут завтра в это время у ворот Самарии",
2KGS|7|19|тогда отвечал этот сановник человеку Божию и сказал: "если бы Господь и открыл окна на небе, и тогда может ли это быть?" А он сказал: "увидишь твоими глазами, но есть этого не будешь".
2KGS|7|20|Так и сбылось с ним; и затоптал его народ в воротах, и он умер.
2KGS|8|1|И говорил Елисей женщине, сына которой воскресил он, и сказал: встань, и пойди, ты и дом твой, и поживи там, где можешь пожить, ибо призвал Господь голод, и он придет на сию землю на семь лет.
2KGS|8|2|И встала та женщина, и сделала по слову человека Божия; и пошла она и дом ее, и жила в земле Филистимской семь лет.
2KGS|8|3|По прошествии семи лет возвратилась эта женщина из земли Филистимской и пришла просить царя о доме своем и о поле своем.
2KGS|8|4|Царь тогда разговаривал с Гиезием, слугою человека Божия, и сказал: расскажи мне все замечательное, что сделал Елисей.
2KGS|8|5|И между тем как он рассказывал царю, что тот воскресил умершего, женщина, которой сына воскресил он, просила царя о доме своем и о поле своем. И сказал Гиезий: господин мой царь, это та самая женщина и тот самый сын ее, которого воскресил Елисей.
2KGS|8|6|И спросил царь у женщины, и она рассказала ему. И дал ей царь одного из придворных, сказав: возвратить ей все принадлежащее ей и все доходы с поля, с того дня, как она оставила землю, поныне.
2KGS|8|7|И пришел Елисей в Дамаск, когда Венадад, царь Сирийский, был болен. И донесли ему, говоря: пришел человек Божий сюда.
2KGS|8|8|И сказал царь Азаилу: возьми в руку твою дар и пойди навстречу человеку Божию, и вопроси Господа чрез него, говоря: выздоровею ли я от сей болезни?
2KGS|8|9|И пошел Азаил навстречу ему, и взял дар в руку свою и всего лучшего в Дамаске, сколько могут нести сорок верблюдов, и пришел и стал пред лице его, и сказал: сын твой Венадад, царь Сирийский, послал меня к тебе спросить: "выздоровею ли я от сей болезни?"
2KGS|8|10|И сказал ему Елисей: пойди, скажи ему: "выздоровеешь"; однакож открыл мне Господь, что он умрет.
2KGS|8|11|И устремил на него [Елисей] взор свой, и так оставался до того, что привел его в смущение; и заплакал человек Божий.
2KGS|8|12|И сказал Азаил: отчего господин мой плачет? И сказал он: от того, что я знаю, какое наделаешь ты сынам Израилевым зло; крепости их предашь огню, и юношей их мечом умертвишь, и грудных детей их побьешь, и беременных [женщин] у них разрубишь.
2KGS|8|13|И сказал Азаил: что такое раб твой, пес, чтобы мог сделать такое большое дело? И сказал Елисей: указал мне Господь в тебе царя Сирии.
2KGS|8|14|И пошел он от Елисея, и пришел к государю своему. И сказал ему [этот]: что говорил тебе Елисей? И сказал: он говорил мне, что ты выздоровеешь.
2KGS|8|15|А на другой день он взял одеяло, намочил его водою, и положил на лице его, и он умер. И воцарился Азаил вместо него.
2KGS|8|16|В пятый год Иорама, сына Ахавова, царя Израильского, за Иосафатом, царем Иудейским, воцарился Иорам, сын Иосафатов, царь Иудейский.
2KGS|8|17|Тридцати двух лет был он, когда воцарился, и восемь лет царствовал в Иерусалиме,
2KGS|8|18|и ходил путем царей Израильских, как поступал дом Ахавов, потому что дочь Ахава была женою его, и делал неугодное в очах Господних.
2KGS|8|19|Однакож не хотел Господь погубить Иуду, ради Давида, раба Своего, так как Он обещал дать ему светильник в детях его на все времена.
2KGS|8|20|Во дни его выступил Едом из–под руки Иуды, и поставили они над собою царя.
2KGS|8|21|И пошел Иорам в Цаир, и все колесницы с ним; и встал он ночью, и поразил Идумеян, окружавших его, и начальников над колесницами, но народ убежал в шатры свои.
2KGS|8|22|И выступил Едом из–под руки Иуды до сего дня. В то же время выступила и Ливна.
2KGS|8|23|Прочее об Иораме и обо всем, что он сделал, написано в летописи царей Иудейских.
2KGS|8|24|И почил Иорам с отцами своими, и погребен с отцами своими в городе Давидовом. И воцарился Охозия, сын его, вместо него.
2KGS|8|25|В двенадцатый год Иорама, сына Ахавова, царя Израильского, воцарился Охозия, сын Иорама, царя Иудейского.
2KGS|8|26|Двадцати двух лет был Охозия, когда воцарился, и один год царствовал в Иерусалиме. Имя же матери его Гофолия, дочь Амврия, царя Израильского.
2KGS|8|27|И ходил путем дома Ахавова, и делал неугодное в очах Господних, подобно дому Ахавову, потому что он был в родстве с домом Ахавовым.
2KGS|8|28|И пошел он с Иорамом, сыном Ахавовым, на войну с Азаилом, царем Сирийским, в Рамоф Галаадский, и ранили Сирияне Иорама.
2KGS|8|29|И возвратился Иорам царь, чтобы лечиться в Изрееле от ран, которые причинили ему Сирияне в Рамофе, когда он воевал с Азаилом, царем Сирийским. И Охозия, сын Иорама, царь Иудейский, пришел посетить Иорама, сына Ахавова, в Изреель, так как он был болен.
2KGS|9|1|Елисей пророк призвал одного из сынов пророческих и сказал ему: опояшь чресла твои, и возьми сей сосуд с елеем в руку твою, и пойди в Рамоф Галаадский.
2KGS|9|2|Придя туда, отыщи там Ииуя, сына Иосафата, сына Намессиева, и подойди, и вели выступить ему из среды братьев своих, и введи его во внутреннюю комнату;
2KGS|9|3|и возьми сосуд с елеем, и вылей на голову его, и скажи: "так говорит Господь: помазую тебя в царя над Израилем". Потом отвори дверь, и беги, и не жди.
2KGS|9|4|И пошел отрок, слуга пророка, в Рамоф Галаадский,
2KGS|9|5|и пришел, и вот сидят военачальники. И сказал: у меня слово до тебя, военачальник. И сказал Ииуй: до кого из всех нас? И сказал он: до тебя, военачальник.
2KGS|9|6|И встал он, и вошел в дом. И [отрок] вылил елей на голову его, и сказал ему: так говорит Господь Бог Израилев: "помазую тебя в царя над народом Господним, над Израилем,
2KGS|9|7|и ты истребишь дом Ахава, господина твоего, чтобы Мне отмстить за кровь рабов Моих пророков и за кровь всех рабов Господних, [павших] от руки Иезавели;
2KGS|9|8|и погибнет весь дом Ахава, и истреблю у Ахава мочащегося к стене, и заключенного и оставшегося в Израиле,
2KGS|9|9|и сделаю дом Ахава, как дом Иеровоама, сына Наватова, и как дом Ваасы, сына Ахиина;
2KGS|9|10|Иезавель же съедят псы на поле Изреельском, и никто не похоронит ее". И отворил дверь, и убежал.
2KGS|9|11|И вышел Ииуй к слугам господина своего, и сказали ему: с миром ли? Зачем приходил этот неистовый к тебе? И сказал им: вы знаете этого человека и что он говорит.
2KGS|9|12|И сказали: неправда, скажи нам. И сказал он: то и то он сказал мне, говоря: "так говорит Господь: помазую тебя в царя над Израилем".
2KGS|9|13|И поспешили они, и взяли каждый одежду свою, и подостлали ему на самых ступенях, и затрубили трубою, и сказали: воцарился Ииуй!
2KGS|9|14|И восстал Ииуй, сын Иосафата, сына Намессиева, против Иорама; Иорам же находился со всеми Израильтянами в Рамофе Галаадском на страже против Азаила, царя Сирийского.
2KGS|9|15|Впрочем сам царь Иорам возвратился, чтобы лечиться в Изрееле от ран, которые причинили ему Сирияне, когда он воевал с Азаилом, царем Сирийским. И сказал Ииуй: если вы согласны, то пусть никто не уходит из города, чтобы идти подать весть в Изрееле.
2KGS|9|16|И сел Ииуй на коня, и поехал в Изреель, где лежал Иорам, и куда Охозия, царь Иудейский, пришел посетить Иорама.
2KGS|9|17|На башне в Изрееле стоял сторож, и увидел он полчище Ииуево, когда оно шло, и сказал: полчище вижу я. И сказал Иорам: возьми всадника, и пошли навстречу им, и пусть скажет: с миром ли?
2KGS|9|18|И выехал всадник на коне навстречу ему, и сказал: так говорит царь: с миром ли? И сказал Ииуй: что тебе до мира? Поезжай за мною. И донес сторож, и сказал: доехал до них, но не возвращается.
2KGS|9|19|И послали другого всадника, и он приехал к ним, и сказал: так говорит царь: с миром ли? И сказал Ииуй: что тебе до мира? Поезжай за мною.
2KGS|9|20|И донес сторож, сказав: доехал до них, и не возвращается, а походка, как будто Ииуя, сына Намессиева, потому что он идет стремительно.
2KGS|9|21|И сказал Иорам: запрягай. И запрягли колесницу его. И выступил Иорам, царь Израильский, и Охозия, царь Иудейский, каждый на колеснице своей. И выступили навстречу Ииую, и встретились с ним на поле Навуфея Изреелитянина.
2KGS|9|22|И когда увидел Иорам Ииуя, то сказал: с миром ли Ииуй? И сказал он: какой мир при любодействе Иезавели, матери твоей, и при многих волхвованиях ее?
2KGS|9|23|И поворотил Иорам руки свои, и побежал, и сказал Охозии: измена, Охозия!
2KGS|9|24|А Ииуй натянул лук рукою своею, и поразил Иорама между плечами его, и прошла стрела чрез сердце его, и пал он на колеснице своей.
2KGS|9|25|И сказал Ииуй Бидекару, сановнику своему: возьми, брось его на участок поля Навуфея Изреелитянина, ибо вспомни, как мы с тобою ехали вдвоем сзади Ахава, отца его, и как Господь изрек на него такое пророчество:
2KGS|9|26|истинно, кровь Навуфея и кровь сыновей его видел Я вчера, говорит Господь, и отмщу тебе на сем поле. Итак возьми, брось его на поле, по слову Господню.
2KGS|9|27|Охозия, царь Иудейский, увидев сие, побежал по дороге к дому, что в саду. И погнался за ним Ииуй, и сказал: и его бейте на колеснице. [Это] [было] на возвышенности Гур, что при Ивлеаме. И побежал он в Мегиддон, и умер там.
2KGS|9|28|И отвезли его рабы его в Иерусалим, и похоронили его в гробнице его, с отцами его, в городе Давидовом.
2KGS|9|29|В одиннадцатый год Иорама, сына Ахавова, воцарился Охозия в Иудее.
2KGS|9|30|И прибыл Ииуй в Изреель. Иезавель же, получив весть, нарумянила лице свое и украсила голову свою, и глядела в окно.
2KGS|9|31|Когда Ииуй вошел в ворота, она сказала: мир ли Замврию, убийце государя своего?
2KGS|9|32|И поднял он лице свое к окну и сказал: кто со мною, кто? И выглянули к нему два, три евнуха.
2KGS|9|33|И сказал он: выбросьте ее. И выбросили ее. И брызнула кровь ее на стену и на коней, и растоптали ее.
2KGS|9|34|И пришел Ииуй, и ел, и пил, и сказал: отыщите эту проклятую и похороните ее, так как царская дочь она.
2KGS|9|35|И пошли хоронить ее, и не нашли от нее ничего, кроме черепа, и ног, и кистей рук.
2KGS|9|36|И возвратились, и донесли ему. И сказал он: таково было слово Господа, которое Он изрек чрез раба Своего Илию Фесвитянина, сказав: на поле Изреельском съедят псы тело Иезавели,
2KGS|9|37|и будет труп Иезавели на участке Изреельском, как навоз на поле, так что никто не скажет: это Иезавель.
2KGS|10|1|У Ахава было семьдесят сыновей в Самарии. И написал Ииуй письма, и послал в Самарию к начальникам Изреельским, старейшинам и воспитателям детей Ахавовых, такого содержания:
2KGS|10|2|когда придет это письмо к вам, то, так как у вас и сыновья господина вашего, у вас же и колесницы, и кони, и укрепленный город, и оружие, –
2KGS|10|3|выберите лучшего и достойнейшего из сыновей государя своего, и посадите на престол отца его, и воюйте за дом государя своего.
2KGS|10|4|Они испугались чрезвычайно и сказали: вот, два царя не устояли перед ним, как же нам устоять?
2KGS|10|5|И послал начальствующий над домом [царским], и градоначальник, и старейшины, и воспитатели к Ииую, сказать: мы рабы твои, и что скажешь нам, то и сделаем; мы никого не поставим царем, что угодно тебе, то и делай.
2KGS|10|6|И написал он к ним письмо во второй раз такое: если вы мои и слову моему повинуетесь, то возьмите головы сыновей государя своего, и придите ко мне завтра в это время в Изреель. (Царских же сыновей было семьдесят человек; воспитывали их знатнейшие в городе.)
2KGS|10|7|Когда пришло к ним письмо, они взяли царских сыновей, и закололи их – семьдесят человек, и положили головы их в корзины, и послали к нему в Изреель.
2KGS|10|8|И пришел посланный, и донес ему, и сказал: принесли головы сыновей царских. И сказал он: разложите их на две груды у входа в ворота, до утра.
2KGS|10|9|Поутру он вышел, и стал, и сказал всему народу: вы невиновны. Вот я восстал против государя моего и умертвил его, а их всех кто убил?
2KGS|10|10|Знайте же теперь, что не падет на землю ни одно слово Господа, которое Он изрек о доме Ахава; Господь сделал то, что изрек чрез раба Своего Илию.
2KGS|10|11|И умертвил Ииуй всех оставшихся из дома Ахава в Изрееле, и всех вельмож его, и близких его, и священников его, так что не осталось от него ни одного уцелевшего.
2KGS|10|12|И встал, и пошел, и пришел в Самарию. Находясь на пути при Беф–Екеде пастушеском,
2KGS|10|13|встретил Ииуй братьев Охозии, царя Иудейского, и сказал: кто вы? Они сказали: мы братья Охозии, идем узнать о здоровье сыновей царя и сыновей государыни.
2KGS|10|14|И сказал он: возьмите их живых. И взяли их живых, и закололи их – сорок два человека, при колодезе Беф–Екеда, и не осталось из них ни одного.
2KGS|10|15|И поехал оттуда, и встретился с Ионадавом, сыном Рихавовым, [шедшим] навстречу ему, и приветствовал его, и сказал ему: расположено ли твое сердце так, как мое сердце к твоему сердцу? И сказал Ионадав: да. Если так, то дай руку твою. И подал он руку свою, и приподнял он его к себе в колесницу,
2KGS|10|16|и сказал: поезжай со мною, и смотри на мою ревность о Господе. И посадили его в колесницу.
2KGS|10|17|Прибыв в Самарию, он убил всех, остававшихся у Ахава в Самарии, так что совсем истребил его, по слову Господа, которое Он изрек Илии.
2KGS|10|18|И собрал Ииуй весь народ и сказал им: Ахав мало служил Ваалу; Ииуй будет служить ему более.
2KGS|10|19|Итак созовите ко мне всех пророков Ваала, всех служителей его и всех священников его, чтобы никто не был в отсутствии, потому что у меня будет великая жертва Ваалу. А всякий, кто не явится, не останется жив. Ииуй делал [это] с хитрым намерением, чтобы истребить служителей Ваала.
2KGS|10|20|И сказал Ииуй: назначьте праздничное собрание ради Ваала. И провозгласили [собрание].
2KGS|10|21|И послал Ииуй по всему Израилю, и пришли все служители Ваала; не оставалось ни одного человека, кто бы не пришел; и вошли в дом Ваалов, и наполнился дом Ваалов от края до края.
2KGS|10|22|И сказал он хранителю одежд: принеси одежду для всех служителей Ваала. И он принес им одежду.
2KGS|10|23|И вошел Ииуй с Ионадавом, сыном Рихавовым, в дом Ваалов, и сказал служителям Ваала: разведайте и разглядите, не находится ли у вас кто–нибудь из служителей Господних, так как здесь должны находиться только одни служители Ваала.
2KGS|10|24|И приступили они к совершению жертв и всесожжений. А Ииуй поставил вне [дома] восемьдесят человек и сказал: душа того, у которого спасется кто–либо из людей, которых я отдаю вам в руки, будет вместо души [спасшегося].
2KGS|10|25|Когда кончено было всесожжение, сказал Ииуй скороходам и начальникам: пойдите, бейте их, чтобы ни один не ушел. И поразили их острием меча и бросили [их] скороходы и начальники, и пошли в город, где было капище Ваалово.
2KGS|10|26|И вынесли статуи из капища Ваалова и сожгли их.
2KGS|10|27|И разбили статую Ваала, и разрушили капище Ваалово; и сделали из него место нечистот, до сего дня.
2KGS|10|28|И истребил Ииуй Ваала с земли Израильской.
2KGS|10|29|Впрочем от грехов Иеровоама, сына Наватова, который ввел Израиля в грех, от них не отступал Ииуй, – от золотых тельцов, которые в Вефиле и которые в Дане.
2KGS|10|30|И сказал Господь Ииую: за то, что ты охотно сделал, что было праведно в очах Моих, выполнил над домом Ахавовым все, что было на сердце у Меня, сыновья твои до четвертого рода будут сидеть на престоле Израилевом.
2KGS|10|31|Но Ииуй не старался ходить в законе Господа Бога Израилева, от всего сердца. Он не отступал от грехов Иеровоама, который ввел Израиля в грех.
2KGS|10|32|В те дни начал Господь отрезать части от Израильтян, и поражал их Азаил во всем пределе Израилевом,
2KGS|10|33|на восток от Иордана, всю землю Галаад, [колено] Гадово, Рувимово, Манассиино, [начиная] от Ароера, который при потоке Арноне, и Галаад и Васан.
2KGS|10|34|Прочее об Ииуе и обо всем, что он сделал, и о мужественных подвигах его написано в летописи царей Израильских.
2KGS|10|35|И почил Ииуй с отцами своими, и похоронили его в Самарии. И воцарился Иоахаз, сын его, вместо него.
2KGS|10|36|Времени же царствования Ииуева над Израилем, в Самарии, было двадцать восемь лет.
2KGS|11|1|Гофолия, мать Охозии, видя, что сын ее умер, встала и истребила все царское племя.
2KGS|11|2|Но Иосавеф, дочь царя Иорама, сестра Охозии, взяла Иоаса, сына Охозии, и тайно увела его из среды умерщвляемых сыновей царских, его и кормилицу его, в постельную комнату; и скрыли его от Гофолии, и он не умерщвлен.
2KGS|11|3|И был он с нею скрываем в доме Господнем шесть лет, между тем как Гофолия царствовала над землею.
2KGS|11|4|В седьмой год послал Иодай, и взял сотников из телохранителей и скороходов, и привел их к себе в дом Господень, и сделал с ними договор, и взял с них клятву в доме Господнем, и показал им царского сына.
2KGS|11|5|И дал им приказание, сказав: вот что вы сделайте: третья часть из вас, из приходящих в субботу, будет содержать стражу при царском доме;
2KGS|11|6|третья часть у ворот Сур, и третья часть у ворот сзади телохранителей, и содержите стражу дома, чтобы не было повреждения;
2KGS|11|7|и две части из вас, из всех отходящих в субботу, будут содержать стражу при доме Господнем для царя;
2KGS|11|8|и окружите царя со всех сторон, каждый с оружием своим в руке своей; и кто вошел бы в ряды, тот да будет умерщвлен. И будьте при царе, когда он выходит и когда входит.
2KGS|11|9|И сделали сотники все, что приказал Иодай священник, и взяли каждый людей своих, приходящих в субботу и отходящих в субботу, и пришли к Иодаю священнику.
2KGS|11|10|И раздал священник сотникам копья и щиты царя Давида, которые были в доме Господнем.
2KGS|11|11|И стали скороходы, каждый с оружием в руке своей, от правой стороны дома до левой стороны дома, у жертвенника и у дома, вокруг царя.
2KGS|11|12|И вывел он царского сына, и возложил на него [царский] венец и украшения, и воцарили его, и помазали его, и рукоплескали и восклицали: да живет царь!
2KGS|11|13|И услышала Гофолия голос бегущего народа, и пошла к народу в дом Господень.
2KGS|11|14|И видит, и вот царь стоит на возвышении, по обычаю, и князья и трубы подле царя; и весь народ земли веселится, и трубят трубами. И разодрала Гофолия одежды свои, и закричала: заговор! заговор!
2KGS|11|15|И дал приказание Иодай священник сотникам, начальствующим над войском, и сказал им: "выведите ее за ряды, а кто пойдет за нею, умерщвляйте мечом", так как думал священник, чтобы не умертвили ее в доме Господнем.
2KGS|11|16|И дали ей место, и она прошла чрез вход конский к дому царскому, и умерщвлена там.
2KGS|11|17|И заключил Иодай завет между Господом и между царем и народом, чтоб он был народом Господним, и между царем и народом.
2KGS|11|18|И пошел весь народ земли в дом Ваала, и разрушили жертвенники его, и изображения его совершенно разбили, и Матфана, жреца Ваалова, убили пред жертвенниками. И учредил священник наблюдение над домом Господним.
2KGS|11|19|И взял сотников и телохранителей и скороходов и весь народ земли, и проводили царя из дома Господня, и пришли по дороге чрез ворота телохранителей в дом царский; и он воссел на престоле царей.
2KGS|11|20|И веселился весь народ земли, и город успокоился. А Гофолию умертвили мечом в царском доме.
2KGS|12|1|Семи лет был Иоас, когда воцарился.
2KGS|12|2|В седьмой год Ииуя воцарился Иоас и сорок лет царствовал в Иерусалиме. Имя матери его Цивья, из Вирсавии.
2KGS|12|3|И делал Иоас угодное в очах Господних во все дни свои, доколе наставлял его священник Иодай;
2KGS|12|4|только высоты не были отменены; народ еще приносил жертвы и курения на высотах.
2KGS|12|5|И сказал Иоас священникам: все серебро посвящаемое, которое приносят в дом Господень, серебро от приходящих, серебро, [вносимое] за каждую душу по оценке, все серебро, сколько кому приходит на сердце принести в дом Господень,
2KGS|12|6|пусть берут священники себе, каждый от своего знакомого, и пусть исправляют они поврежденное в храме, везде, где найдется повреждение.
2KGS|12|7|Но как до двадцать третьего года царя Иоаса священники не исправляли повреждений в храме,
2KGS|12|8|то царь Иоас позвал священника Иодая и священников и сказал им: почему вы не исправляете повреждений в храме? Не берите же отныне серебра у знакомых своих, а на [починку] повреждений в храме отдайте его.
2KGS|12|9|И согласились священники не брать серебра у народа на исправление повреждений в храме.
2KGS|12|10|И взял священник Иодай один ящик, и сделал отверстие сверху его, и поставил его подле жертвенника на правой стороне, где входили в дом Господень. И полагали туда священники, стоящие на страже у порога, все серебро, приносимое в дом Господень.
2KGS|12|11|И когда видели, что много серебра в ящике, приходили писец царский и первосвященник, и завязывали [в мешки], и пересчитывали серебро, найденное в доме Господнем;
2KGS|12|12|и отдавали сосчитанное серебро в руки производителям работ, приставленным к дому Господню, а сии издерживали его на плотников и строителей, работавших в доме Господнем,
2KGS|12|13|и на делателей стен и на каменотесов, также на покупку дерев и тесаных камней, для починки повреждений в доме Господнем, и на все, что расходовалось для поддержания храма.
2KGS|12|14|Но не сделано было для дома Господня серебряных блюд, ножей, чаш [для окропления], труб, всяких сосудов золотых и сосудов серебряных из серебра, приносимого в дом Господень,
2KGS|12|15|а производителям работ отдавали его, и починивали им дом Господень.
2KGS|12|16|И не требовали отчета от тех людей, которым поручали серебро для раздачи производителям работ, ибо они действовали честно.
2KGS|12|17|Серебро за жертву о преступлении и серебро за жертву о грехе не вносилось в дом Господень: священникам оно принадлежало.
2KGS|12|18|Тогда выступил в поход Азаил, царь Сирийский, и пошел войною на Геф, и взял его; и вознамерился Азаил идти на Иерусалим.
2KGS|12|19|Но Иоас, царь Иудейский, взял все пожертвованное, что пожертвовали [храму] Иосафат, и Иорам и Охозия, отцы его, цари Иудейские, и что он сам пожертвовал, и все золото, найденное в сокровищницах дома Господня и дома царского, и послал Азаилу, царю Сирийскому; и он отступил от Иерусалима.
2KGS|12|20|Прочее об Иоасе и обо всем, что он сделал, написано в летописи царей Иудейских.
2KGS|12|21|И восстали слуги его, и составили заговор, и убили Иоаса в доме Милло, на дороге к Силле.
2KGS|12|22|Его убили слуги его: Иозакар, сын Шимеаты, и Иегозавад, сын Шомеры; и он умер, и похоронили его с отцами его в городе Давидовом. И воцарился Амасия, сын его, вместо него.
2KGS|13|1|В двадцать третий год Иоаса, сына Охозиина, царя Иудейского, воцарился Иоахаз, сын Ииуя, над Израилем в Самарии, [и царствовал] семнадцать лет,
2KGS|13|2|и делал неугодное в очах Господних, и ходил в грехах Иеровоама, сына Наватова, который ввел Израиля в грех, и не отставал от них.
2KGS|13|3|И возгорелся гнев Господа на Израиля, и Он предавал их в руку Азаила, царя Сирийского, и в руку Венадада, сына Азаилова, во все дни.
2KGS|13|4|И помолился Иоахаз лицу Господню, и услышал его Господь, потому что видел стеснение Израильтян, как теснил их царь Сирийский.
2KGS|13|5|И дал Господь Израильтянам избавителя, и вышли они из–под руки Сириян, и жили сыны Израилевы в шатрах своих, как вчера и третьего дня.
2KGS|13|6|Однакож не отступали от грехов дома Иеровоама, который ввел Израиля в грех; ходили в них, и дубрава стояла в Самарии.
2KGS|13|7|У Иоахаза оставалось войска только пятьдесят всадников, десять колесниц и десять тысяч пеших, от того, что истребил их царь Сирийский и обратил их в прах на попрание.
2KGS|13|8|Прочее об Иоахазе и обо всем, что он сделал, и о мужественных подвигах его, написано в летописи царей Израильских.
2KGS|13|9|И почил Иоахаз с отцами своими, и похоронили его в Самарии. И воцарился Иоас, сын его, вместо него.
2KGS|13|10|В тридцать седьмой год Иоаса, царя Иудейского, воцарился Иоас, сын Иоахазов, над Израилем в Самарии, [и царствовал] шестнадцать лет,
2KGS|13|11|и делал неугодное в очах Господних; не отставал от всех грехов Иеровоама, сына Наватова, который ввел Израиля в грех, но ходил в них.
2KGS|13|12|Прочее об Иоасе и обо всем, что он сделал, и о мужественных подвигах его, как он воевал с Амасиею, царем Иудейским, написано в летописи царей Израильских.
2KGS|13|13|И почил Иоас с отцами своими, а Иеровоам сел на престоле его. И погребен Иоас в Самарии с царями Израильскими.
2KGS|13|14|Елисей заболел болезнью, от которой [потом] и умер. И пришел к нему Иоас, царь Израильский, и плакал над ним, и говорил: отец мой! отец мой! колесница Израиля и конница его!
2KGS|13|15|И сказал ему Елисей: возьми лук и стрелы. И взял он лук и стрелы.
2KGS|13|16|И сказал царю Израильскому: положи руку твою на лук. И положил он руку свою. И наложил Елисей руки свои на руки царя,
2KGS|13|17|и сказал: отвори окно на восток. И он отворил. И сказал Елисей: выстрели. И он выстрелил. И сказал: эта стрела избавления от Господа и стрела избавления против Сирии, и ты поразишь Сириян в Афеке вконец.
2KGS|13|18|И сказал [Елисей]: возьми стрелы. И он взял. И сказал царю Израильскому: бей по земле. И ударил он три раза, и остановился.
2KGS|13|19|И разгневался на него человек Божий, и сказал: надобно было бы бить пять или шесть раз, тогда ты побил бы Сириян совершенно, а теперь [только] три раза поразишь Сириян.
2KGS|13|20|И умер Елисей, и похоронили его. И полчища Моавитян пришли в землю в следующем году.
2KGS|13|21|И было, что, когда погребали одного человека, то, увидев это полчище, [погребавшие] бросили того человека в гроб Елисеев; и он при падении своем коснулся костей Елисея, и ожил, и встал на ноги свои.
2KGS|13|22|Азаил, царь Сирийский, теснил Израильтян во все дни Иоахаза.
2KGS|13|23|Но Господь умилосердился над ними, и помиловал их, и обратился к ним ради завета Своего с Авраамом, Исааком и Иаковом, и не хотел истребить их, и не отверг их от лица Своего доныне.
2KGS|13|24|И умер Азаил, царь Сирийский, и воцарился Венадад, сын его, вместо него.
2KGS|13|25|И взял назад Иоас, сын Иоахаза, из руки Венадада, сына Азаила, города, которые он взял войною из руки отца его Иоахаза. Три раза разбил его Иоас и возвратил города Израилевы.
2KGS|14|1|Во второй год Иоаса, сына Иоахазова, царя Израильского, воцарился Амасия, сын Иоаса, царь Иудейский:
2KGS|14|2|двадцати пяти лет был он, когда воцарился, и двадцать девять лет царствовал в Иерусалиме. Имя матери его Иегоаддань, из Иерусалима.
2KGS|14|3|И делал он угодное в очах Господних, впрочем не так, как отец его Давид: он во всем поступал так, как отец его Иоас.
2KGS|14|4|Только высоты не были отменены: народ совершал еще жертвы и курения на высотах.
2KGS|14|5|Когда утвердилось царство в руках его, тогда он умертвил слуг своих, убивших царя, отца его.
2KGS|14|6|Но детей убийц не умертвил, так как написано в книге закона Моисеева, в которой заповедал Господь, говоря: "не должны быть наказываемы смертью отцы за детей, и дети не должны быть наказываемы смертью за отцов, но каждый за свое преступление должен быть наказываем смертью".
2KGS|14|7|Он поразил десять тысяч Идумеян на долине Соляной, и взял Селу войною, и дал ей имя Иокфеил, которое [остается и] до сего дня.
2KGS|14|8|Тогда послал Амасия послов к Иоасу, царю Израильскому, сыну Иоахаза, сына Ииуева, сказать: выйди, повидаемся лично.
2KGS|14|9|И послал Иоас, царь Израильский, к Амасии, царю Иудейскому, сказать: терн, который на Ливане, послал к кедру, который на Ливане же, сказать: "отдай дочь свою в жену сыну моему". Но прошли дикие звери, что на Ливане, и истоптали этот терн.
2KGS|14|10|Ты поразил Идумеян, и возгордилось сердце твое. Величайся и сиди у себя дома. К чему тебе затевать ссору на свою беду? Падешь ты и Иуда с тобою.
2KGS|14|11|Но не послушался Амасия. И выступил Иоас, царь Израильский, и увиделись лично он и Амасия, царь Иудейский, в Вефсамисе, что в Иудее.
2KGS|14|12|И разбиты были Иудеи Израильтянами, и разбежались по шатрам своим.
2KGS|14|13|И Амасию, царя Иудейского, сына Иоаса, сына Охозиина, захватил Иоас, царь Израильский, в Вефсамисе, и пошел в Иерусалим и разрушил стену Иерусалимскую от ворот Ефремовых до ворот угольных на четыреста локтей.
2KGS|14|14|И взял все золото и серебро, и все сосуды, какие нашлись в доме Господнем и в сокровищницах царского дома, и заложников, и возвратился в Самарию.
2KGS|14|15|Прочее об Иоасе, что он сделал, и о мужественных подвигах его, и как он воевал с Амасиею, царем Иудейским, написано в летописи царей Израильских.
2KGS|14|16|И почил Иоас с отцами своими, и погребен в Самарии с царями Израильскими. И воцарился Иеровоам, сын его, вместо него.
2KGS|14|17|И жил Амасия, сын Иоасов, царь Иудейский, по смерти Иоаса, сына Иоахазова, царя Израильского, пятнадцать лет.
2KGS|14|18|Прочие дела Амасии записаны в летописи царей Иудейских.
2KGS|14|19|И составили против него заговор в Иерусалиме, и убежал он в Лахис. И послали за ним в Лахис, и умертвили его там.
2KGS|14|20|И привезли его на конях, и погребен он был в Иерусалиме с отцами своими в городе Давидовом.
2KGS|14|21|И взял весь народ Иудейский Азарию, которому было шестнадцать лет, и воцарили его вместо отца его Амасии.
2KGS|14|22|Он обстроил Елаф, и возвратил его Иуде, после того как царь почил с отцами своими.
2KGS|14|23|В пятнадцатый год Амасии, сына Иоасова, царя Иудейского, воцарился Иеровоам, сын Иоасов, царь Израильский, в Самарии, и [царствовал] сорок один год,
2KGS|14|24|и делал он неугодное в очах Господних: не отступал от всех грехов Иеровоама, сына Наватова, который ввел Израиля в грех.
2KGS|14|25|Он восстановил пределы Израиля, от входа в Емаф до моря пустыни, по слову Господа Бога Израилева, которое Он изрек чрез раба Своего Иону, сына Амафиина, пророка из Гафхефера,
2KGS|14|26|ибо Господь видел бедствие Израиля, весьма горькое, так что не оставалось ни заключенного, ни оставшегося, и не было помощника у Израиля.
2KGS|14|27|И не восхотел Господь искоренить имя Израильтян из поднебесной, и спас их рукою Иеровоама, сына Иоасова.
2KGS|14|28|Прочее об Иеровоаме и обо всем, что он сделал, и о мужественных подвигах его, как он воевал и как возвратил Израилю Дамаск и Емаф, принадлежавших Иуде, написано в летописи царей Израильских.
2KGS|14|29|И почил Иеровоам с отцами своими, с царями Израильскими. И воцарился Захария, сын его, вместо него.
2KGS|15|1|В двадцать седьмой год Иеровоама, царя Израильского, воцарился Азария, сын Амасии, царь Иудейский:
2KGS|15|2|шестнадцати лет был он, когда воцарился, и пятьдесят два года царствовал в Иерусалиме. Имя матери его Иехолия, из Иерусалима.
2KGS|15|3|Он делал угодное в очах Господних во всем так, как поступал Амасия, отец его.
2KGS|15|4|Только высоты не были отменены: народ совершал еще жертвы и курения на высотах.
2KGS|15|5|И поразил Господь царя, и был он прокаженным до дня смерти своей и жил в отдельном доме. И Иофам, сын царя, [начальствовал] над дворцом и управлял народом земли.
2KGS|15|6|Прочее об Азарии и обо всем, что он сделал, написано в летописи царей Иудейских.
2KGS|15|7|И почил Азария с отцами своими, и похоронили его с отцами его в городе Давидовом. И воцарился Иофам, сын его, вместо него.
2KGS|15|8|В тридцать восьмой год Азарии, царя Иудейского, воцарился Захария, сын Иеровоама, над Израилем в Самарии [и царствовал] шесть месяцев.
2KGS|15|9|Он делал неугодное в очах Господних, как делали отцы его: не отставал от грехов Иеровоама, сына Наватова, который ввел Израиля в грех.
2KGS|15|10|И составил против него заговор Селлум, сын Иависа, и поразил его пред народом и убил его, и воцарился вместо него.
2KGS|15|11|Прочее о Захарии написано в летописи царей Израильских.
2KGS|15|12|Таково было слово Господа, которое он изрек Ииую, сказав: сыновья твои до четвертого рода будут сидеть на престоле Израилевом. И сбылось так.
2KGS|15|13|Селлум, сын Иависа, воцарился в тридцать девятый год Азарии, царя Иудейского, и царствовал один месяц в Самарии.
2KGS|15|14|И пошел Менаим, сын Гадия из Фирцы, и пришел в Самарию, и поразил Селлума, сына Иависова, в Самарии и умертвил его, и воцарился вместо него.
2KGS|15|15|Прочее о Селлуме и о заговоре его, который он составил, написано в летописи царей Израильских.
2KGS|15|16|И поразил Менаим Типсах и всех, которые были в нем и в пределах его, [начиная] от Фирцы, за то, что [город] не отворил [ворот], и разбил [его], и всех беременных женщин в нем разрубил.
2KGS|15|17|В тридцать девятом году Азарии, царя Иудейского, воцарился Менаим, сын Гадия, над Израилем [и царствовал] десять лет в Самарии;
2KGS|15|18|и делал он неугодное в очах Господних; не отставал от грехов Иеровоама, сына Наватова, который ввел Израиля в грех, во все дни свои.
2KGS|15|19|Тогда пришел Фул, царь Ассирийский, на землю [Израилеву]. И дал Менаим Фулу тысячу талантов серебра, чтобы руки его были за него и чтобы утвердить царство в руке своей.
2KGS|15|20|И разложил Менаим это серебро на Израильтян, на всех людей богатых, по пятидесяти сиклей серебра на каждого человека, чтобы отдать царю Ассирийскому. И пошел назад царь Ассирийский и не остался там в земле.
2KGS|15|21|Прочее о Менаиме и обо всем, что он сделал, написано в летописи царей Израильских.
2KGS|15|22|И почил Менаим с отцами своими. И воцарился Факия, сын его, вместо него.
2KGS|15|23|В пятидесятый год Азарии, царя Иудейского, воцарился Факия, сын Менаима, над Израилем в Самарии [и царствовал] два года;
2KGS|15|24|и делал он неугодное в очах Господних; не отставал от грехов Иеровоама, сына Наватова, который ввел Израиля в грех.
2KGS|15|25|И составил против него заговор Факей, сын Ремалии, сановник его, и поразил его в Самарии в палате царского дома, с Арговом и Арием, имея с собою пятьдесят человек Галаадитян, и умертвил его, и воцарился вместо него.
2KGS|15|26|Прочее о Факии и обо всем, что он сделал, написано в летописи царей Израильских.
2KGS|15|27|В пятьдесят второй год Азарии, царя Иудейского, воцарился Факей, сын Ремалии, над Израилем в Самарии [и царствовал] двадцать лет;
2KGS|15|28|и делал он неугодное в очах Господних: не отставал от грехов Иеровоама, сына Наватова, который ввел Израиля в грех.
2KGS|15|29|Во дни Факея, царя Израильского, пришел Феглаффелласар, царь Ассирийский, и взял Ион, Авел–Беф–Мааху, и Ианох, и Кедес, и Асор, и Галаад, и Галилею, всю землю Неффалимову, и переселил их в Ассирию.
2KGS|15|30|И составил заговор Осия, сын Илы, против Факея, сына Ремалиина, и поразил его, и умертвил его, и воцарился вместо него в двадцатый год Иоафама, сына Озиина.
2KGS|15|31|Прочее о Факее и обо всем, что он сделал, написано в летописи царей Израильских.
2KGS|15|32|Во второй год Факея, сына Ремалиина, царя Израильского, воцарился Иоафам, сын Озии, царя Иудейского.
2KGS|15|33|Двадцати пяти лет был он, когда воцарился, и шестнадцать лет царствовал в Иерусалиме. Имя матери его Иеруша, дочь Садока.
2KGS|15|34|Он делал угодное в очах Господних: во всем, как поступал Озия, отец его, так поступал и он.
2KGS|15|35|Только высоты не были отменены: народ совершал еще жертвы и курения на высотах. Он построил верхние ворота при доме Господнем.
2KGS|15|36|Прочее об Иоафаме и обо всем, что он сделал, написано в летописи царей Иудейских.
2KGS|15|37|В те дни начал Господь посылать на Иудею Рецина, царя Сирийского, и Факея, сына Ремалиина.
2KGS|15|38|И почил Иоафам с отцами своими, и погребен с отцами своими в городе Давида, отца его. И воцарился Ахаз, сын его, вместо него.
2KGS|16|1|В семнадцатый год Факея, сына Ремалиина, воцарился Ахаз, сын Иоафама, царя Иудейского.
2KGS|16|2|Двадцати лет был Ахаз, когда воцарился, и шестнадцать лет царствовал в Иерусалиме, и не делал угодного в очах Господа Бога своего, как Давид, отец его,
2KGS|16|3|но ходил путем царей Израильских, и даже сына своего провел чрез огонь, [подражая] мерзостям народов, которых прогнал Господь от лица сынов Израилевых,
2KGS|16|4|и совершал жертвы и курения на высотах и на холмах и под всяким тенистым деревом.
2KGS|16|5|Тогда пошел Рецин, царь Сирийский, и Факей, сын Ремалиин, царь Израильский, против Иерусалима, чтобы завоевать его, и держали Ахаза в осаде, но одолеть не могли.
2KGS|16|6|В то время Рецин, царь Сирийский, возвратил Сирии Елаф и изгнал Иудеев из Елафа; и Идумеяне вступили в Елаф, и живут там до сего дня.
2KGS|16|7|И послал Ахаз послов к Феглаффелласару, царю Ассирийскому, сказать: раб твой и сын твой я; приди и защити меня от руки царя Сирийского и от руки царя Израильского, восставших на меня.
2KGS|16|8|И взял Ахаз серебро и золото, какое нашлось в доме Господнем и в сокровищницах дома царского, и послал царю Ассирийскому в дар.
2KGS|16|9|И послушал его царь Ассирийский; и пошел царь Ассирийский в Дамаск, и взял его, и переселил жителей его в Кир, а Рецина умертвил.
2KGS|16|10|И пошел царь Ахаз навстречу Феглаффелласару, царю Ассирийскому, в Дамаск, и увидел жертвенник, который в Дамаске, и послал царь Ахаз к Урии священнику изображение жертвенника и чертеж всего устройства его.
2KGS|16|11|И построил священник Урия жертвенник по образцу, который прислал царь Ахаз из Дамаска; и сделал так священник Урия до прибытия царя Ахаза из Дамаска.
2KGS|16|12|И пришел царь из Дамаска, и увидел царь жертвенник, и подошел царь к жертвеннику, и принес на нем жертву;
2KGS|16|13|и сожег всесожжение свое и хлебное приношение, и совершил возлияние свое, и окропил кровью мирной жертвы свой жертвенник.
2KGS|16|14|А медный жертвенник, который пред лицем Господним, он передвинул от лицевой стороны храма, с [места] между жертвенником [новым] и домом Господним, и поставил его сбоку [сего] жертвенника на север.
2KGS|16|15|И дал приказание царь Ахаз священнику Урии, сказав: на большом жертвеннике сожигай утреннее всесожжение и вечернее хлебное приношение, и всесожжение от царя и хлебное приношение от него, и всесожжение от всех людей земли и хлебное приношение от них, и возлияние от них, и всякою кровью всесожжений и всякою кровью жертв окропляй его, а жертвенник медный останется до моего усмотрения.
2KGS|16|16|И сделал священник Урия все так, как приказал царь Ахаз.
2KGS|16|17|И обломал царь Ахаз ободки у подстав, и снял с них умывальницы, и море снял с медных волов, которые [были] под ним, и поставил его на каменный пол.
2KGS|16|18|И отменил крытый субботний ход, который построили при храме, и внешний царский вход к дому Господню, ради царя Ассирийского.
2KGS|16|19|Прочее об Ахазе, что он сделал, написано в летописи царей Иудейских.
2KGS|16|20|И почил Ахаз с отцами своими, и погребен с отцами своими в городе Давидовом. И воцарился Езекия, сын его, вместо него.
2KGS|17|1|В двенадцатый год Ахаза, царя Иудейского, воцарился Осия, сын Илы, в Самарии над Израилем [и царствовал] девять лет.
2KGS|17|2|И делал он неугодное в очах Господних, но не так, как цари Израильские, которые были прежде него.
2KGS|17|3|Против него выступил Салманассар, царь Ассирийский, и сделался Осия подвластным ему и давал ему дань.
2KGS|17|4|И заметил царь Ассирийский в Осии измену, так как он посылал послов к Сигору, царю Египетскому, и не доставлял дани царю Ассирийскому каждый год; и взял его царь Ассирийский под стражу, и заключил его в дом темничный.
2KGS|17|5|И пошел царь Ассирийский на всю землю, и приступил к Самарии, и держал ее в осаде три года.
2KGS|17|6|В девятый год Осии взял царь Ассирийский Самарию, и переселил Израильтян в Ассирию, и поселил их в Халахе и в Хаворе, при реке Гозан, и в городах Мидийских.
2KGS|17|7|Когда стали грешить сыны Израилевы пред Господом Богом своим, Который вывел их из земли Египетской, из–под руки фараона, царя Египетского, и стали чтить богов иных,
2KGS|17|8|и стали поступать по обычаям народов, которых прогнал Господь от лица сынов Израилевых, и [по обычаям] царей Израильских, как поступали они;
2KGS|17|9|и стали делать сыны Израилевы дела неугодные Господу Богу своему, и построили себе высоты во всех городах своих, [начиная] от сторожевой башни до укрепленного города,
2KGS|17|10|и поставили у себя статуи и изображения Астарт на всяком высоком холме и под всяким тенистым деревом,
2KGS|17|11|и стали там совершать курения на всех высотах, подобно народам, которых изгнал от них Господь, и делали худые дела, прогневляющие Господа,
2KGS|17|12|и служили идолам, о которых говорил им Господь: "не делайте сего";
2KGS|17|13|тогда Господь чрез всех пророков Своих, чрез всякого прозорливца предостерегал Израиля и Иуду, говоря: возвратитесь со злых путей ваших и соблюдайте заповеди Мои, уставы Мои, по всему учению, которое Я заповедал отцам вашим и которое Я преподал вам чрез рабов Моих, пророков.
2KGS|17|14|Но они не слушали и ожесточили выю свою, как была выя отцов их, которые не веровали в Господа, Бога своего;
2KGS|17|15|и презирали уставы Его, и завет Его, который Он заключил с отцами их, и откровения Его, какими Он предостерегал их, и пошли вслед суеты и осуетились, и вслед народов окрестных, о которых Господь заповедал им, чтобы не поступали так, как они,
2KGS|17|16|и оставили все заповеди Господа Бога своего, и сделали себе литые изображения двух тельцов, и устроили дубраву, и поклонялись всему воинству небесному, и служили Ваалу,
2KGS|17|17|и проводили сыновей своих и дочерей своих чрез огонь, и гадали, и волшебствовали, и предались тому, чтобы делать неугодное в очах Господа и прогневлять Его.
2KGS|17|18|И прогневался Господь сильно на Израильтян, и отверг их от лица Своего. Не осталось никого, кроме одного колена Иудина.
2KGS|17|19|И Иуда также не соблюдал заповедей Господа Бога своего, и поступал по обычаям Израильтян, как поступали они.
2KGS|17|20|И отвратился Господь от всех потомков Израиля, и смирил их, и отдавал их в руки грабителям, и наконец отверг их от лица Своего.
2KGS|17|21|Израильтяне отторглись от дома Давидова и воцарили Иеровоама, сына Наватова; и отклонил Иеровоам Израильтян от Господа, и вовлек их в великий грех.
2KGS|17|22|И поступали сыны Израилевы по всем грехам Иеровоама, какие он делал, не отставали от них,
2KGS|17|23|доколе Господь не отверг Израиля от лица Своего, как говорил чрез всех рабов Своих, пророков. И переселен Израиль из земли своей в Ассирию, где он и до сего дня.
2KGS|17|24|И перевел царь Ассирийский людей из Вавилона, и из Куты, и из Аввы, и из Емафа, и из Сепарваима, и поселил [их] в городах Самарийских вместо сынов Израилевых. И они овладели Самариею, и стали жить в городах ее.
2KGS|17|25|И как в начале жительства своего там они не чтили Господа, то Господь посылал на них львов, которые умерщвляли их.
2KGS|17|26|И донесли царю Ассирийскому, и сказали: народы, которых ты переселил и поселил в городах Самарийских, не знают закона Бога той земли, и за то Он посылает на них львов, и вот они умерщвляют их, потому что они не знают закона Бога той земли.
2KGS|17|27|И повелел царь Ассирийский, и сказал: отправьте туда одного из священников, которых вы выселили оттуда; пусть пойдет и живет там, и он научит их закону Бога той земли.
2KGS|17|28|И пришел один из священников, которых выселили из Самарии, и жил в Вефиле, и учил их, как чтить Господа.
2KGS|17|29|Притом сделал каждый народ и своих богов и поставил в капищах высот, какие устроили Самаряне, – каждый народ в своих городах, где живут они.
2KGS|17|30|Вавилоняне сделали Суккот–Беноф, Кутийцы сделали Нергала, Емафяне сделали Ашиму,
2KGS|17|31|Аввийцы сделали Нивхаза и Тартака, а Сепарваимцы сожигали сыновей своих в огне Адрамелеху и Анамелеху, богам Сепарваимским.
2KGS|17|32|Между тем чтили и Господа, и сделали у себя священников высот из среды своей, и они служили у них в капищах высот.
2KGS|17|33|Господа они чтили, и богам своим они служили по обычаю народов, из которых выселили их.
2KGS|17|34|До сего дня поступают они по прежним своим обычаям: не боятся Господа и не поступают по уставам и по обрядам, и по закону и по заповедям, которые заповедал Господь сынам Иакова, которому дал Он имя Израиля.
2KGS|17|35|Заключил Господь с ними завет и заповедал им, говоря: не чтите богов иных, и не поклоняйтесь им, и не служите им, и не приносите жертв им,
2KGS|17|36|но Господа, Который вывел вас из земли Египетской силою великою и мышцею простертою, – Его чтите и Ему поклоняйтесь, и Ему приносите жертвы,
2KGS|17|37|и уставы, и учреждения, и закон, и заповеди, которые Он написал вам, старайтесь исполнять во все дни, и не чтите богов иных;
2KGS|17|38|и завета, который Я заключил с вами, не забывайте, и не чтите богов иных,
2KGS|17|39|только Господа Бога вашего чтите, и Он избавит вас от руки всех врагов ваших.
2KGS|17|40|Но они не послушали, а поступали по прежним своим обычаям.
2KGS|17|41|Народы сии чтили Господа, но и истуканам своим служили. Да и дети их и дети детей их до сего дня поступают так же, как поступали отцы их.
2KGS|18|1|В третий год Осии, сына Илы, царя Израильского, воцарился Езекия, сын Ахаза, царя Иудейского.
2KGS|18|2|Двадцати пяти лет был он, когда воцарился, и двадцать девять лет царствовал в Иерусалиме; имя матери его Ави, дочь Захарии.
2KGS|18|3|И делал он угодное в очах Господних во всем так, как делал Давид, отец его;
2KGS|18|4|он отменил высоты, разбил статуи, срубил дубраву и истребил медного змея, которого сделал Моисей, потому что до самых тех дней сыны Израилевы кадили ему и называли его Нехуштан.
2KGS|18|5|На Господа Бога Израилева уповал он; и такого, как он, не бывало между всеми царями Иудейскими и после него и прежде него.
2KGS|18|6|И прилепился он к Господу и не отступал от Него, и соблюдал заповеди Его, какие заповедал Господь Моисею.
2KGS|18|7|И был Господь с ним: везде, куда он ни ходил, поступал он благоразумно. И отложился он от царя Ассирийского, и не стал служить ему.
2KGS|18|8|Он поразил Филистимлян до Газы и в пределах ее, от сторожевой башни до укрепленного города.
2KGS|18|9|В четвертый год царя Езекии, то есть в седьмой год Осии, сына Илы, царя Израильского, пошел Салманассар, царь Ассирийский, на Самарию, и осадил ее,
2KGS|18|10|и взял ее через три года; в шестой год Езекии, то есть в девятый год Осии, царя Израильского, взята Самария.
2KGS|18|11|И переселил царь Ассирийский Израильтян в Ассирию, и поселил их в Халахе и в Хаворе, при реке Гозан, и в городах Мидийских,
2KGS|18|12|за то, что они не слушали гласа Господа Бога своего и преступили завет Его, все, что заповедал Моисей раб Господень, они и не слушали и не исполняли.
2KGS|18|13|В четырнадцатый год царя Езекии, пошел Сеннахирим, царь Ассирийский, против всех укрепленных городов Иуды и взял их.
2KGS|18|14|И послал Езекия, царь Иудейский, к царю Ассирийскому в Лахис сказать: виновен я; отойди от меня; что наложишь на меня, я внесу. И наложил царь Ассирийский на Езекию, царя Иудейского, триста талантов серебра и тридцать талантов золота.
2KGS|18|15|И отдал Езекия все серебро, какое нашлось в доме Господнем и в сокровищницах дома царского.
2KGS|18|16|В то время снял Езекия [золото] с дверей дома Господня и с дверных столбов, которые позолотил Езекия, царь Иудейский, и отдал его царю Ассирийскому.
2KGS|18|17|И послал царь Ассирийский Тартана и Рабсариса и Рабсака из Лахиса к царю Езекии с большим войском в Иерусалим. И пошли, и пришли к Иерусалиму; и пошли, и пришли, и стали у водопровода верхнего пруда, который на дороге поля белильничьего.
2KGS|18|18|И звали они царя. И вышел к ним Елиаким, сын Хелкиин, начальник дворца, и Севна писец, и Иоах, сын Асафов, дееписатель.
2KGS|18|19|И сказал им Рабсак: скажите Езекии: так говорит царь великий, царь Ассирийский: что это за упование, на которое ты уповаешь?
2KGS|18|20|Ты говорил только пустые слова: для войны нужны совет и сила. Ныне же на кого ты уповаешь, что отложился от меня?
2KGS|18|21|Вот, ты думаешь опереться на Египет, на эту трость надломленную, которая, если кто опрется на нее, войдет ему в руку и проколет ее. Таков фараон, царь Египетский, для всех уповающих на него.
2KGS|18|22|А если вы скажете мне: "на Господа Бога нашего мы уповаем", то на того ли, которого высоты и жертвенники отменил Езекия, и сказал Иуде и Иерусалиму: "пред сим только жертвенником поклоняйтесь в Иерусалиме"?
2KGS|18|23|Итак вступи в союз с господином моим царем Ассирийским: я дам тебе две тысячи коней, можешь ли достать себе всадников на них?
2KGS|18|24|Как тебе одолеть и одного вождя из малейших слуг господина моего? И уповаешь на Египет ради колесниц и коней?
2KGS|18|25|Притом же разве я без воли Господней пошел на место сие, чтобы разорить его? Господь сказал мне: "пойди на землю сию и разори ее".
2KGS|18|26|И сказал Елиаким, сын Хелкиин, и Севна и Иоах Рабсаку: говори рабам твоим по–арамейски, потому что понимаем мы, а не говори с нами по–иудейски вслух народа, который на стене.
2KGS|18|27|И сказал им Рабсак: разве [только] к господину твоему и к тебе послал меня господин мой сказать сии слова? Нет, также и к людям, которые сидят на стене, чтобы есть помет свой и пить мочу свою с вами.
2KGS|18|28|И встал Рабсак и возгласил громким голосом по–иудейски, и говорил, и сказал: слушайте слово царя великого, царя Ассирийского!
2KGS|18|29|Так говорит царь: пусть не обольщает вас Езекия, ибо он не может вас спасти от руки моей;
2KGS|18|30|и пусть не обнадеживает вас Езекия Господом, говоря: "спасет нас Господь и не будет город сей отдан в руки царя Ассирийского".
2KGS|18|31|Не слушайте Езекии. Ибо так говорит царь Ассирийский: примиритесь со мною и выйдите ко мне, и пусть каждый ест [плоды] виноградной лозы своей и смоковницы своей, и пусть каждый пьет воду из своего колодезя,
2KGS|18|32|пока я не приду и не возьму вас в землю такую же, как и ваша земля, в землю хлеба и вина, в землю плодов и виноградников, в землю масличных дерев и меда, и будете жить, и не умрете. Не слушайте же Езекии, который обольщает вас, говоря: "Господь спасет нас".
2KGS|18|33|Спасли ли боги народов, каждый свою землю, от руки царя Ассирийского?
2KGS|18|34|Где боги Емафа и Арпада? Где боги Сепарваима, Ены и Иввы? Спасли ли они Самарию от руки моей?
2KGS|18|35|Кто из всех богов земель сих спас землю свою от руки моей? Так неужели Господь спасет Иерусалим от руки моей?
2KGS|18|36|И молчал народ и не отвечали ему ни слова, потому что было приказание царя: "не отвечайте ему".
2KGS|18|37|И пришел Елиаким, сын Хелкиин, начальник дворца, и Севна писец и Иоах, сын Асафов, дееписатель, к Езекии в разодранных одеждах, и пересказали ему слова Рабсаковы.
2KGS|19|1|Когда услышал [это] царь Езекия, то разодрал одежды свои и покрылся вретищем, и пошел в дом Господень.
2KGS|19|2|И послал Елиакима, начальника дворца, и Севну писца, и старших священников, покрытых вретищами, к Исаии пророку, сыну Амосову.
2KGS|19|3|И они сказали ему: так говорит Езекия: день скорби и наказания и посрамления – день сей; ибо дошли младенцы до отверстия утробы матерней, а силы нет родить.
2KGS|19|4|Может быть, услышит Господь Бог твой все слова Рабсака, которого послал царь Ассирийский, господин его, хулить Бога живаго и поносить словами, какие слышал Господь Бог твой. Принеси же молитву об оставшихся, которые находятся еще в живых.
2KGS|19|5|И пришли слуги царя Езекии к Исаии,
2KGS|19|6|и сказал им Исаия: так скажите господину вашему: так говорит Господь: не бойся слов, которые ты слышал, которыми поносили Меня слуги царя Ассирийского.
2KGS|19|7|Вот Я пошлю в него дух, и он услышит весть, и возвратится в землю свою, и Я поражу его мечом в земле его.
2KGS|19|8|И возвратился Рабсак, и нашел царя Ассирийского воюющим против Ливны, ибо он слышал, что тот отошел от Лахиса.
2KGS|19|9|И услышал он о Тиргаке, царе Ефиопском; ему сказали: вот, он вышел сразиться с тобою. И снова послал он послов к Езекии сказать:
2KGS|19|10|так скажите Езекии, царю Иудейскому: пусть не обманывает тебя Бог твой, на Которого ты уповаешь, думая: "не будет отдан Иерусалим в руки царя Ассирийского".
2KGS|19|11|Ведь ты слышал, что сделали цари Ассирийские со всеми землями, положив на них заклятие, – и ты ли уцелеешь?
2KGS|19|12|Боги народов, которых разорили отцы мои, спасли ли их? [Спасли] [ли] Гозан, и Харан, и Рецеф, и сынов Едена, что в Фалассаре?
2KGS|19|13|Где царь Емафа, и царь Арпада, и царь города Сепарваима, Ены и Иввы?
2KGS|19|14|И взял Езекия письмо из руки послов, и прочитал его, и пошел в дом Господень, и развернул его Езекия пред лицем Господним,
2KGS|19|15|и молился Езекия пред лицем Господним и говорил: Господи Боже Израилев, седящий на Херувимах! Ты один Бог всех царств земли, Ты сотворил небо и землю.
2KGS|19|16|Приклони, Господи, ухо Твое и услышь; открой, Господи, очи Твои и воззри, и услышь слова Сеннахирима, который послал поносить Бога живаго!
2KGS|19|17|Правда, о, Господи, цари Ассирийские разорили народы и земли их,
2KGS|19|18|и побросали богов их в огонь; но это не боги, а изделие рук человеческих, дерево и камень; потому и истребили их.
2KGS|19|19|И ныне, Господи Боже наш, спаси нас от руки его, и узнают все царства земли, что Ты, Господи, Бог один.
2KGS|19|20|И послал Исаия, сын Амосов, к Езекии сказать: так говорит Господь Бог Израилев: то, о чем ты молился Мне против Сеннахирима, царя Ассирийского, Я услышал.
2KGS|19|21|Вот слово, которое изрек Господь о нем: презрит тебя, посмеется над тобою девствующая дочь Сиона; вслед тебя покачает головою дочь Иерусалима.
2KGS|19|22|Кого ты порицал и поносил? И на кого ты возвысил голос и поднял так высоко глаза свои? На Святаго Израилева!
2KGS|19|23|Чрез послов твоих ты порицал Господа и сказал: "со множеством колесниц моих я взошел на высоту гор, на ребра Ливана, и срубил рослые кедры его, отличные кипарисы его, и пришел на самое крайнее пристанище его, в рощу сада его;
2KGS|19|24|и откапывал я и пил воду чужую, и осушу ступнями ног моих все реки Египетские".
2KGS|19|25|Разве ты не слышал, что Я издавна сделал это, в древние дни предначертал это, а ныне выполнил тем, что ты опустошаешь укрепленные города, [превращая] в груды развалин?
2KGS|19|26|И жители их сделались маломощны, трепещут и остаются в стыде. Они стали [как] трава на поле и нежная зелень, [как] порост на кровлях и опаленный хлеб, прежде нежели выколосился.
2KGS|19|27|Сядешь ли ты, выйдешь ли, войдешь ли, Я все знаю; [знаю] и дерзость твою против Меня.
2KGS|19|28|За твою дерзость против Меня и [за то, что] надмение твое дошло до ушей Моих, Я вложу кольцо Мое в ноздри твои и удила Мои в рот твой, и возвращу тебя назад тою же дорогою, которою пришел ты.
2KGS|19|29|И вот тебе, [Езекия], знамение: ешьте в этот год выросшее от упавшего зерна, и в другой год – самородное, а на третий год сейте и жните, и садите виноградные сады и ешьте плоды их.
2KGS|19|30|И уцелевшее в доме Иудином, оставшееся пустит опять корень внизу и принесет плод вверху,
2KGS|19|31|ибо из Иерусалима произойдет остаток, и спасенное от горы Сиона. Ревность Господа Саваофа сделает сие.
2KGS|19|32|Посему так говорит Господь о царе Ассирийском: "не войдет он в сей город, и не бросит туда стрелы, и не приступит к нему со щитом, и не насыплет против него вала.
2KGS|19|33|Тою же дорогою, которою пришел, возвратится, и в город сей не войдет, говорит Господь.
2KGS|19|34|Я буду охранять город сей, чтобы спасти его ради Себя и ради Давида, раба Моего".
2KGS|19|35|И случилось в ту ночь: пошел Ангел Господень и поразил в стане Ассирийском сто восемьдесят пять тысяч. И встали поутру, и вот все тела мертвые.
2KGS|19|36|И отправился, и пошел, и возвратился Сеннахирим, царь Ассирийский, и жил в Ниневии.
2KGS|19|37|И когда он поклонялся в доме Нисроха, бога своего, то Адрамелех и Шарецер, сыновья его, убили его мечом, а сами убежали в землю Араратскую. И воцарился Асардан, сын его, вместо него.
2KGS|20|1|В те дни заболел Езекия смертельно, и пришел к нему Исаия, сын Амосов, пророк, и сказал ему: так говорит Господь: сделай завещание для дома твоего, ибо умрешь ты и не выздоровеешь.
2KGS|20|2|И отворотился [Езекия] лицем своим к стене и молился Господу, говоря:
2KGS|20|3|"О, Господи! вспомни, что я ходил пред лицем Твоим верно и с преданным [Тебе] сердцем, и делал угодное в очах Твоих". И заплакал Езекия сильно.
2KGS|20|4|Исаия еще не вышел из города, как было к нему слово Господне:
2KGS|20|5|возвратись и скажи Езекии, владыке народа Моего: так говорит Господь Бог Давида, отца твоего: Я услышал молитву твою, увидел слезы твои. Вот, Я исцелю тебя; в третий день пойдешь в дом Господень;
2KGS|20|6|и прибавлю ко дням твоим пятнадцать лет, и от руки царя Ассирийского спасу тебя и город сей, и защищу город сей ради Себя и ради Давида, раба Моего.
2KGS|20|7|И сказал Исаия: возьмите пласт смокв. И взяли, и приложили к нарыву; и он выздоровел.
2KGS|20|8|И сказал Езекия Исаии: какое знамение, что Господь исцелит меня, и что пойду я на третий день в дом Господень?
2KGS|20|9|И сказал Исаия: вот тебе знамение от Господа, что исполнит Господь слово, которое Он изрек: вперед ли пройти тени на десять ступеней, или воротиться на десять ступеней?
2KGS|20|10|И сказал Езекия: легко тени подвинуться вперед на десять ступеней; нет, пусть воротится тень назад на десять ступеней.
2KGS|20|11|И воззвал Исаия пророк к Господу, и возвратил тень назад на ступенях, где она спускалась по ступеням Ахазовым, на десять ступеней.
2KGS|20|12|В то время послал Беродах Баладан, сын Баладана, царь Вавилонский, письма и подарок Езекии, ибо он слышал, что Езекия был болен.
2KGS|20|13|Езекия, выслушав посланных, показал им кладовые свои, серебро и золото, и ароматы, и масти дорогие, и весь оружейный дом свой и все, что находилось в сокровищницах его; не оставалось ни одной вещи, которой не показал бы им Езекия в доме своем и во всем владении своем.
2KGS|20|14|И пришел Исаия пророк к царю Езекии и сказал ему: что говорили эти люди, и откуда они приходили к тебе? И сказал Езекия: из земли далекой они приходили, из Вавилона.
2KGS|20|15|И сказал [Исаия]: что они видели в доме твоем? И сказал Езекия: все, что в доме моем, они видели, не осталось ни одной вещи, которой я не показал бы им в сокровищницах моих.
2KGS|20|16|И сказал Исаия Езекии: выслушай слово Господне:
2KGS|20|17|вот придут дни, и взято будет все, что в доме твоем, и что собрали отцы твои до сего дня, в Вавилон; ничего не останется, говорит Господь.
2KGS|20|18|Из сынов твоих, которые произойдут от тебя, которых ты родишь, возьмут, и будут они евнухами во дворце царя Вавилонского.
2KGS|20|19|И сказал Езекия Исаии: благо слово Господне, которое ты изрек. И продолжал: да будет мир и благосостояние во дни мои!
2KGS|20|20|Прочее об Езекии и о всех подвигах его, и о том, что он сделал пруд и водопровод и провел воду в город, написано в летописи царей Иудейских.
2KGS|20|21|И почил Езекия с отцами своими, и воцарился Манассия, сын его, вместо него.
2KGS|21|1|Двенадцати лет был Манассия, когда воцарился, и пятьдесят лет царствовал в Иерусалиме; имя матери его Хефциба.
2KGS|21|2|И делал он неугодное в очах Господних, [подражая] мерзостям народов, которых прогнал Господь от лица сынов Израилевых.
2KGS|21|3|И снова устроил высоты, которые уничтожил отец его Езекия, и поставил жертвенники Ваалу, и сделал дубраву, как сделал Ахав, царь Израильский; и поклонялся всему воинству небесному, и служил ему.
2KGS|21|4|И соорудил жертвенники в доме Господнем, о котором сказал Господь: "в Иерусалиме положу имя Мое".
2KGS|21|5|И соорудил жертвенники всему воинству небесному на обоих дворах дома Господня,
2KGS|21|6|и провел сына своего чрез огонь, и гадал, и ворожил, и завел вызывателей мертвецов и волшебников; много сделал неугодного в очах Господа, чтобы прогневать Его.
2KGS|21|7|И поставил истукан Астарты, который сделал в доме, о котором говорил Господь Давиду и Соломону, сыну его: "в доме сем и в Иерусалиме, который Я избрал из всех колен Израилевых, Я полагаю имя Мое на век;
2KGS|21|8|и не дам впредь выступить ноге Израильтянина из земли, которую Я дал отцам их, если только они будут стараться поступать согласно со всем тем, что Я повелел им, и со всем законом, который заповедал им раб Мой Моисей".
2KGS|21|9|Но они не послушались; и совратил их Манассия до того, что они поступали хуже тех народов, которых истребил Господь от лица сынов Израилевых.
2KGS|21|10|И говорил Господь чрез рабов Своих пророков и сказал:
2KGS|21|11|за то, что сделал Манассия, царь Иудейский, такие мерзости, хуже всего того, что делали Аморреи, которые были прежде его, и ввел Иуду в грех идолами своими,
2KGS|21|12|за то, так говорит Господь, Бог Израилев, вот, Я наведу такое зло на Иерусалим и на Иуду, о котором кто услышит, зазвенит в обоих ушах у того;
2KGS|21|13|и протяну на Иерусалим мерную вервь Самарии и отвес дома Ахавова, и вытру Иерусалим так, как вытирают чашу, – вытрут и опрокинут ее;
2KGS|21|14|и отвергну остаток удела Моего, и отдам их в руку врагов их, и будут на расхищение и разграбление всем неприятелям своим,
2KGS|21|15|за то, что они делали неугодное в очах Моих и прогневляли Меня с того дня, как вышли отцы их из Египта, и до сего дня.
2KGS|21|16|Еще же пролил Манассия и весьма много невинной крови, так что наполнил [ею] Иерусалим от края до края, сверх своего греха, что он завлек Иуду в грех – делать неугодное в очах Господних.
2KGS|21|17|Прочее о Манассии и обо всем, что он сделал, и о грехах его, в чем он согрешил, написано в летописи царей Иудейских.
2KGS|21|18|И почил Манассия с отцами своими, и погребен в саду при доме его, в саду Уззы. И воцарился Аммон, сын его, вместо него.
2KGS|21|19|Двадцати двух лет был Аммон, когда воцарился, и два года царствовал в Иерусалиме; имя матери его Мешуллемеф, дочь Харуца, из Ятбы.
2KGS|21|20|И делал он неугодное в очах Господних так, как делал Манассия, отец его;
2KGS|21|21|и ходил тою же точно дорогою, которою ходил отец его, и служил идолам, которым служил отец его, и поклонялся им,
2KGS|21|22|и оставил Господа Бога отцов своих, не ходил путем Господним.
2KGS|21|23|И составили заговор слуги Аммоновы против него, и умертвили царя в доме его.
2KGS|21|24|Но народ земли перебил всех, бывших в заговоре против царя Аммона; и воцарил народ земли Иосию, сына его, вместо него.
2KGS|21|25|Прочее об Аммоне, что он сделал, написано в летописи царей Иудейских.
2KGS|21|26|И похоронили его в гробнице его, в саду Уззы. И воцарился Иосия, сын его, вместо него.
2KGS|22|1|Восьми лет был Иосия, когда воцарился, и тридцать один год царствовал в Иерусалиме; имя матери его Иедида, дочь Адаии, из Боцкафы.
2KGS|22|2|И делал он угодное в очах Господних, и ходил во всем путем Давида, отца своего, и не уклонялся ни направо, ни налево.
2KGS|22|3|В восемнадцатый год царя Иосии, послал царь Шафана, сына Ацалии, сына Мешулламова, писца, в дом Господень, сказав:
2KGS|22|4|пойди к Хелкии первосвященнику, пусть он пересчитает серебро, принесенное в дом Господень, которое собрали от народа стоящие на страже у порога,
2KGS|22|5|и пусть отдадут его в руки производителям работ, приставленным к дому Господню, а сии пусть раздают его работающим в доме Господнем, на исправление повреждений дома,
2KGS|22|6|плотникам и каменщикам, и делателям стен, и на покупку дерев и тесаных камней для исправления дома;
2KGS|22|7|впрочем не требовать у них отчета в серебре, переданном в руки их, потому что они поступают честно.
2KGS|22|8|И сказал Хелкия первосвященник Шафану писцу: книгу закона я нашел в доме Господнем. И подал Хелкия книгу Шафану, и он читал ее.
2KGS|22|9|И пришел Шафан писец к царю, и принес царю ответ, и сказал: взяли рабы твои серебро, найденное в доме, и передали его в руки производителям работ, приставленным к дому Господню.
2KGS|22|10|И донес Шафан писец царю, говоря: книгу дал мне Хелкия священник. И читал ее Шафан пред царем.
2KGS|22|11|Когда услышал царь слова книги закона, то разодрал одежды свои.
2KGS|22|12|И повелел царь Хелкии священнику, и Ахикаму, сыну Шафанову, и Ахбору, сыну Михеину, и Шафану писцу, и Асаии, слуге царскому, говоря:
2KGS|22|13|пойдите, вопросите Господа за меня и за народ и за всю Иудею о словах сей найденной книги, потому что велик гнев Господень, который воспылал на нас за то, что не слушали отцы наши слов книги сей, чтобы поступать согласно с предписанным нам.
2KGS|22|14|И пошел Хелкия священник, и Ахикам, и Ахбор, и Шафан, и Асаия к Олдаме пророчице, жене Шаллума, сына Тиквы, сына Хархаса, хранителя одежд, – жила же она в Иерусалиме, во второй части, – и говорили с нею.
2KGS|22|15|И она сказала им: так говорит Господь, Бог Израилев: скажите человеку, который послал вас ко мне:
2KGS|22|16|так говорит Господь: наведу зло на место сие и на жителей его, – все слова книги, которую читал царь Иудейский.
2KGS|22|17|За то, что оставили Меня, и кадят другим богам, чтобы раздражать Меня всеми делами рук своих, воспылал гнев Мой на место сие, и не погаснет.
2KGS|22|18|А царю Иудейскому, пославшему вас вопросить Господа, скажите: так говорит Господь Бог Израилев, о словах, которые ты слышал:
2KGS|22|19|так как смягчилось сердце твое, и ты смирился пред Господом, услышав то, что Я изрек на место сие и на жителей его, что они будут предметом ужаса и проклятия, и ты разодрал одежды свои, и плакал предо Мною, то и Я услышал тебя, говорит Господь.
2KGS|22|20|За это, вот, Я приложу тебя к отцам твоим, и ты положен будешь в гробницу твою в мире, и не увидят глаза твои всего того бедствия, которое Я наведу на место сие. И принесли царю ответ.
2KGS|23|1|И послал царь, и собрали к нему всех старейшин Иуды и Иерусалима.
2KGS|23|2|И пошел царь в дом Господень, и все Иудеи, и все жители Иерусалима с ним, и священники, и пророки, и весь народ, от малого до большого, и прочел вслух их все слова книги завета, найденной в доме Господнем.
2KGS|23|3|Потом стал царь на возвышенное место и заключил пред лицем Господним завет – последовать Господу и соблюдать заповеди Его и откровения Его и уставы Его от всего сердца и от всей души, чтобы выполнить слова завета сего, написанные в книге сей. И весь народ вступил в завет.
2KGS|23|4|И повелел царь Хелкии первосвященнику и вторым священникам и стоящим на страже у порога вынести из храма Господня все вещи, сделанные для Ваала и для Астарты и для всего воинства небесного, и сжег их за Иерусалимом в долине Кедрон, и [велел] прах их отнести в Вефиль.
2KGS|23|5|И отставил жрецов, которых поставили цари Иудейские, чтобы совершать курения на высотах в городах Иудейских и окрестностях Иерусалима, – и которые кадили Ваалу, солнцу, и луне, и созвездиям, и всему воинству небесному;
2KGS|23|6|и вынес Астарту из дома Господня за Иерусалим к потоку Кедрону, и сжег ее у потока Кедрона, и истер ее в прах, и бросил прах ее на кладбище общенародное;
2KGS|23|7|и разрушил домы блудилищные, которые [были] при храме Господнем, где женщины ткали одежды для Астарты;
2KGS|23|8|и вывел всех жрецов из городов Иудейских, и осквернил высоты, на которых совершали курения жрецы, от Гевы до Вирсавии, и разрушил высоты [пред] воротами, – ту, которая у входа в ворота Иисуса градоначальника, и ту, которая на левой стороне у городских ворот.
2KGS|23|9|Впрочем жрецы высот не приносили жертв на жертвеннике Господнем в Иерусалиме, опресноки же ели вместе с братьями своими.
2KGS|23|10|И осквернил он Тофет, что на долине сыновей Еннома, чтобы никто не проводил сына своего и дочери своей чрез огонь Молоху;
2KGS|23|11|и отменил коней, которых ставили цари Иудейские солнцу пред входом в дом Господень близ комнат Нефан–Мелеха евнуха, что в Фаруриме, колесницы же солнца сжег огнем.
2KGS|23|12|И жертвенники на кровле горницы Ахазовой, которые сделали цари Иудейские, и жертвенники, которые сделал Манассия на обоих дворах дома Господня, разрушил царь, и низверг оттуда, и бросил прах их в поток Кедрон.
2KGS|23|13|И высоты, которые пред Иерусалимом, направо от Масличной горы, которые устроил Соломон, царь Израилев, Астарте, мерзости Сидонской, и Хамосу, мерзости Моавитской, и Милхому, мерзости Аммонитской, осквернил царь;
2KGS|23|14|и изломал статуи, и срубил дубравы, и наполнил место их костями человеческими.
2KGS|23|15|Также и жертвенник, который в Вефиле, высоту, устроенную Иеровоамом, сыном Наватовым, который ввел Израиля в грех, – также и жертвенник тот и высоту он разрушил, и сжег сию высоту, стер в прах, и сжег дубраву.
2KGS|23|16|И взглянул Иосия и увидел могилы, которые [были] там на горе, и послал и взял кости из могил, и сжег на жертвеннике, и осквернил его по слову Господню, которое провозгласил человек Божий, предрекший события сии.
2KGS|23|17|и сказал [Иосия]: что это за памятник, который я вижу? И сказали ему жители города: [это] могила человека Божия, который приходил из Иудеи и провозгласил о том, что ты делаешь над жертвенником Вефильским.
2KGS|23|18|И сказал он: оставьте его в покое, никто не трогай костей его. И сохранили кости его и кости пророка, который приходил из Самарии.
2KGS|23|19|Также и все капища высот в городах Самарийских, которые построили цари Израильские, прогневляя [Господа], разрушил Иосия, и сделал с ними то же, что сделал в Вефиле;
2KGS|23|20|и заколол всех жрецов высот, которые там были, на жертвенниках, и сожег кости человеческие на них, – и возвратился в Иерусалим.
2KGS|23|21|И повелел царь всему народу, сказав: "совершите пасху Господу Богу вашему, как написано в сей книге завета", –
2KGS|23|22|потому что не была совершена такая пасха от дней судей, которые судили Израиля, и во все дни царей Израильских и царей Иудейских;
2KGS|23|23|а в восемнадцатый год царя Иосии была совершена сия пасха Господу в Иерусалиме.
2KGS|23|24|И вызывателей мертвых, и волшебников, и терафимов, и идолов, и все мерзости, которые появлялись в земле Иудейской и в Иерусалиме, истребил Иосия, чтоб исполнить слова закона, написанные в книге, которую нашел Хелкия священник в доме Господнем.
2KGS|23|25|Подобного ему не было царя прежде его, который обратился бы к Господу всем сердцем своим, и всею душею своею, и всеми силами своими, по всему закону Моисееву; и после него не восстал подобный ему.
2KGS|23|26|Однакож Господь не отложил великой ярости гнева Своего, какою воспылал гнев Его на Иуду за все оскорбления, какими прогневал Его Манассия.
2KGS|23|27|И сказал Господь: и Иуду отрину от лица Моего, как отринул Я Израиля, и отвергну город сей Иерусалим, который Я избрал, и дом, о котором Я сказал: "будет имя Мое там".
2KGS|23|28|Прочее об Иосии и обо всем, что он сделал, написано в летописи царей Иудейских.
2KGS|23|29|Во дни его пошел фараон Нехао, царь Египетский, против царя Ассирийского на реку Евфрат. И вышел царь Иосия навстречу ему, и тот умертвил его в Мегиддоне, когда увидел его.
2KGS|23|30|И рабы его повезли его мертвого из Мегиддона, и привезли его в Иерусалим, и похоронили его в гробнице его. И взял народ земли Иоахаза, сына Иосиина, и помазали его и воцарили его вместо отца его.
2KGS|23|31|Двадцати трех лет был Иоахаз, когда воцарился, и три месяца царствовал в Иерусалиме; имя матери его Хамуталь, дочь Иеремии, из Ливны.
2KGS|23|32|И делал он неугодное в очах Господних во всем так, как делали отцы его.
2KGS|23|33|И задержал его фараон Нехао в Ривле, в земле Емафской, чтобы он не царствовал в Иерусалиме, – и наложил пени на землю сто талантов серебра и талантов золота.
2KGS|23|34|И воцарил фараон Нехао Елиакима, сына Иосиина, вместо Иосии, отца его, и переменил имя его на Иоакима; Иоахаза же взял и отвел в Египет, где он и умер.
2KGS|23|35|И серебро и золото давал Иоаким фараону; он сделал оценку земле, чтобы давать серебро по приказанию фараона; от каждого из народа земли, по оценке своей, он взыскивал серебро и золото для того, чтобы отдавать фараону Нехао.
2KGS|23|36|Двадцати пяти лет был Иоаким, когда воцарился, и одиннадцать лет царствовал в Иерусалиме; имя матери его Зебудда, дочь Федаии, из Румы.
2KGS|23|37|И делал он неугодное в очах Господних во всем так, как делали отцы его.
2KGS|24|1|Во дни его выступил Навуходоносор, царь Вавилонский, и сделался Иоаким подвластным ему на три года, но потом отложился от него.
2KGS|24|2|И посылал на него Господь полчища Халдеев, и полчища Сириян, и полчища Моавитян, и полчища Аммонитян, – посылал их на Иуду, чтобы погубить его по слову Господа, которое Он изрек чрез рабов Своих пророков.
2KGS|24|3|По повелению Господа было [это] с Иудою, чтобы отвергнуть [его] от лица Его за грехи Манассии, за все, что он сделал;
2KGS|24|4|и за кровь невинную, которую он пролил, наполнив Иерусалим кровью невинною, Господь не захотел простить.
2KGS|24|5|Прочее об Иоакиме и обо всем, что он сделал, написано в летописи царей Иудейских.
2KGS|24|6|И почил Иоаким с отцами своими, и воцарился Иехония, сын его, вместо него.
2KGS|24|7|Царь Египетский не выходил более из земли своей, потому что взял царь Вавилонский все, от потока Египетского до реки Евфрата, что принадлежало царю Египетскому.
2KGS|24|8|Восемнадцати лет был Иехония, когда воцарился, и три месяца царствовал в Иерусалиме; имя матери его Нехушта, дочь Елнафана, из Иерусалима.
2KGS|24|9|И делал он неугодное в очах Господних во всем так, как делал отец его.
2KGS|24|10|В то время подступили рабы Навуходоносора, царя Вавилонского, к Иерусалиму, и подвергся город осаде.
2KGS|24|11|И пришел Навуходоносор, царь Вавилонский, к городу, когда рабы его осаждали его.
2KGS|24|12|И вышел Иехония, царь Иудейский, к царю Вавилонскому, он и мать его, и слуги его, и князья его, и евнухи его, – и взял его царь Вавилонский в восьмой год своего царствования.
2KGS|24|13|И вывез он оттуда все сокровища дома Господня и сокровища царского дома; и изломал, как изрек Господь, все золотые сосуды, которые Соломон, царь Израилев, сделал в храме Господнем;
2KGS|24|14|и выселил весь Иерусалим, и всех князей, и все храброе войско, – десять тысяч было переселенных, – и всех плотников и кузнецов; никого не осталось, кроме бедного народа земли.
2KGS|24|15|И переселил он Иехонию в Вавилон; и мать царя, и жен царя, и евнухов его, и сильных земли отвел на поселение из Иерусалима в Вавилон.
2KGS|24|16|И все войско [числом] семь тысяч, и художников и строителей тысячу, всех храбрых, ходящих на войну, отвел царь Вавилонский на поселение в Вавилон.
2KGS|24|17|И воцарил царь Вавилонский Матфанию, дядю [Иехонии], вместо него, и переменил имя его на Седекию.
2KGS|24|18|Двадцати одного года был Седекия, когда воцарился, и одиннадцать лет царствовал в Иерусалиме; имя матери его Хамуталь, дочь Иеремии, из Ливны.
2KGS|24|19|И делал он неугодное в очах Господних во всем так, как делал Иоаким.
2KGS|24|20|Гнев Господень был над Иерусалимом и над Иудою до того, что Он отверг их от лица Своего. И отложился Седекия от царя Вавилонского.
2KGS|25|1|В девятый год царствования своего, в десятый месяц, в десятый день месяца, пришел Навуходоносор, царь Вавилонский, со всем войском своим к Иерусалиму, и осадил его, и устроил вокруг него вал.
2KGS|25|2|И находился город в осаде до одиннадцатого года царя Седекии.
2KGS|25|3|В девятый день месяца усилился голод в городе, и не было хлеба у народа земли.
2KGS|25|4|И взят был город, и [побежали] все военные ночью по дороге к воротам, между двумя стенами, что подле царского сада; Халдеи же стояли вокруг города, и [царь] ушел дорогою к равнине.
2KGS|25|5|И погналось войско Халдейское за царем, и настигли его на равнинах Иерихонских, и все войско его разбежалось от него.
2KGS|25|6|И взяли царя, и отвели его к царю Вавилонскому в Ривлу, и произвели над ним суд:
2KGS|25|7|и сыновей Седекии закололи пред глазами его, а [самому] Седекии ослепили глаза и сковали его оковами, и отвели его в Вавилон.
2KGS|25|8|В пятый месяц, в седьмой день месяца, то есть в девятнадцатый год Навуходоносора, царя Вавилонского, пришел Навузардан, начальник телохранителей, слуга царя Вавилонского, в Иерусалим
2KGS|25|9|и сжег дом Господень и дом царя, и все домы в Иерусалиме, и все домы большие сожег огнем;
2KGS|25|10|и стены вокруг Иерусалима разрушило войско Халдейское, бывшее у начальника телохранителей.
2KGS|25|11|И прочий народ, остававшийся в городе, и переметчиков, которые передались царю Вавилонскому, и прочий простой народ выселил Навузардан, начальник телохранителей.
2KGS|25|12|Только несколько из бедного народа земли оставил начальник телохранителей работниками в виноградниках и землепашцами.
2KGS|25|13|И столбы медные, которые были у дома Господня, и подставы, и море медное, которое в доме Господнем, изломали Халдеи, и отнесли медь их в Вавилон;
2KGS|25|14|и тазы, и лопатки, и ножи, и ложки, и все сосуды медные, которые употреблялись при служении, взяли;
2KGS|25|15|и кадильницы, и чаши, что было золотое и что было серебряное, взял начальник телохранителей:
2KGS|25|16|столбы [числом] два, море одно, и подставы, которые сделал Соломон в дом Господень, – меди во всех сих вещах не было весу.
2KGS|25|17|Восемнадцать локтей вышины в одном столбе; венец на нем медный, а вышина венца три локтя, и сетка и гранатовые яблоки вокруг венца – все из меди. То же и на другом столбе с сеткою.
2KGS|25|18|И взял начальник телохранителей Сераию первосвященника и Цефанию, священника второго, и трех, стоявших на страже у порога.
2KGS|25|19|И из города взял одного евнуха, который был начальствующим над людьми военными, и пять человек, предстоявших лицу царя, которые находились в городе, и писца главного в войске, записывавшего в войско народ земли, и шестьдесят человек из народа земли, находившихся в городе.
2KGS|25|20|И взял их Навузардан, начальник телохранителей, и отвел их к царю Вавилонскому в Ривлу.
2KGS|25|21|И поразил их царь Вавилонский, и умертвил их в Ривле, в земле Емаф. И выселены Иудеи из земли своей.
2KGS|25|22|Над народом же, остававшимся в земле Иудейской, который оставил Навуходоносор, царь Вавилонский, – над ними поставил начальником Годолию, сына Ахикама, сына Шафанова.
2KGS|25|23|Когда услышали все военачальники, они и люди их, что царь Вавилонский поставил начальником Годолию, то пришли к Годолии в Массифу, и [именно]: Исмаил, сын Нефании, и Иоханан, сын Карея, и Сераия, сын Танхумефа из Нетофафа, и Иезания, сын Маахитянина, они и люди их.
2KGS|25|24|И поклялся Годолия им и людям их, и сказал им: не бойтесь быть подвластными Халдеям, селитесь на земле и служите царю Вавилонскому, и будет хорошо вам.
2KGS|25|25|Но в седьмой месяц пришел Исмаил, сын Нефании, сына Елишамы, из племени царского, с десятью человеками, и поразил Годолию, и он умер, и Иудеев и Халдеев, которые были с ним в Массифе.
2KGS|25|26|И встал весь народ, от малого до большого, и военачальники, и пошли в Египет, потому что боялись Халдеев.
2KGS|25|27|В тридцать седьмой год переселения Иехонии, царя Иудейского, в двенадцатый месяц, в двадцать седьмой день месяца, Евилмеродах, царь Вавилонский, в год своего воцарения, вывел Иехонию, царя Иудейского, из дома темничного
2KGS|25|28|и говорил с ним дружелюбно, и поставил престол его выше престола царей, которые были у него в Вавилоне;
2KGS|25|29|и переменил темничные одежды его, и он всегда имел пищу у него, во все дни жизни его.
2KGS|25|30|И содержание его, содержание постоянное, выдаваемо было ему от царя, изо дня в день, во все дни жизни его.
