COL|1|1|Paul, an apostle of Jesus Christ by the will of God, and Timotheus our brother,
COL|1|2|To the saints and faithful brethren in Christ which are at Colosse: Grace be unto you, and peace, from God our Father and the Lord Jesus Christ.
COL|1|3|We give thanks to God and the Father of our Lord Jesus Christ, praying always for you,
COL|1|4|Since we heard of your faith in Christ Jesus, and of the love which ye have to all the saints,
COL|1|5|For the hope which is laid up for you in heaven, whereof ye heard before in the word of the truth of the gospel;
COL|1|6|Which is come unto you, as it is in all the world; and bringeth forth fruit, as it doth also in you, since the day ye heard of it, and knew the grace of God in truth:
COL|1|7|As ye also learned of Epaphras our dear fellowservant, who is for you a faithful minister of Christ;
COL|1|8|Who also declared unto us your love in the Spirit.
COL|1|9|For this cause we also, since the day we heard it, do not cease to pray for you, and to desire that ye might be filled with the knowledge of his will in all wisdom and spiritual understanding;
COL|1|10|That ye might walk worthy of the Lord unto all pleasing, being fruitful in every good work, and increasing in the knowledge of God;
COL|1|11|Strengthened with all might, according to his glorious power, unto all patience and longsuffering with joyfulness;
COL|1|12|Giving thanks unto the Father, which hath made us meet to be partakers of the inheritance of the saints in light:
COL|1|13|Who hath delivered us from the power of darkness, and hath translated us into the kingdom of his dear Son:
COL|1|14|In whom we have redemption through his blood, even the forgiveness of sins:
COL|1|15|Who is the image of the invisible God, the firstborn of every creature:
COL|1|16|For by him were all things created, that are in heaven, and that are in earth, visible and invisible, whether they be thrones, or dominions, or principalities, or powers: all things were created by him, and for him:
COL|1|17|And he is before all things, and by him all things consist.
COL|1|18|And he is the head of the body, the church: who is the beginning, the firstborn from the dead; that in all things he might have the preeminence.
COL|1|19|For it pleased the Father that in him should all fulness dwell;
COL|1|20|And, having made peace through the blood of his cross, by him to reconcile all things unto himself; by him, I say, whether they be things in earth, or things in heaven.
COL|1|21|And you, that were sometime alienated and enemies in your mind by wicked works, yet now hath he reconciled
COL|1|22|In the body of his flesh through death, to present you holy and unblameable and unreproveable in his sight:
COL|1|23|If ye continue in the faith grounded and settled, and be not moved away from the hope of the gospel, which ye have heard, and which was preached to every creature which is under heaven; whereof I Paul am made a minister;
COL|1|24|Who now rejoice in my sufferings for you, and fill up that which is behind of the afflictions of Christ in my flesh for his body's sake, which is the church:
COL|1|25|Whereof I am made a minister, according to the dispensation of God which is given to me for you, to fulfil the word of God;
COL|1|26|Even the mystery which hath been hid from ages and from generations, but now is made manifest to his saints:
COL|1|27|To whom God would make known what is the riches of the glory of this mystery among the Gentiles; which is Christ in you, the hope of glory:
COL|1|28|Whom we preach, warning every man, and teaching every man in all wisdom; that we may present every man perfect in Christ Jesus:
COL|1|29|Whereunto I also labour, striving according to his working, which worketh in me mightily.
COL|2|1|For I would that ye knew what great conflict I have for you, and for them at Laodicea, and for as many as have not seen my face in the flesh;
COL|2|2|That their hearts might be comforted, being knit together in love, and unto all riches of the full assurance of understanding, to the acknowledgement of the mystery of God, and of the Father, and of Christ;
COL|2|3|In whom are hid all the treasures of wisdom and knowledge.
COL|2|4|And this I say, lest any man should beguile you with enticing words.
COL|2|5|For though I be absent in the flesh, yet am I with you in the spirit, joying and beholding your order, and the stedfastness of your faith in Christ.
COL|2|6|As ye have therefore received Christ Jesus the Lord, so walk ye in him:
COL|2|7|Rooted and built up in him, and stablished in the faith, as ye have been taught, abounding therein with thanksgiving.
COL|2|8|Beware lest any man spoil you through philosophy and vain deceit, after the tradition of men, after the rudiments of the world, and not after Christ.
COL|2|9|For in him dwelleth all the fulness of the Godhead bodily.
COL|2|10|And ye are complete in him, which is the head of all principality and power:
COL|2|11|In whom also ye are circumcised with the circumcision made without hands, in putting off the body of the sins of the flesh by the circumcision of Christ:
COL|2|12|Buried with him in baptism, wherein also ye are risen with him through the faith of the operation of God, who hath raised him from the dead.
COL|2|13|And you, being dead in your sins and the uncircumcision of your flesh, hath he quickened together with him, having forgiven you all trespasses;
COL|2|14|Blotting out the handwriting of ordinances that was against us, which was contrary to us, and took it out of the way, nailing it to his cross;
COL|2|15|And having spoiled principalities and powers, he made a shew of them openly, triumphing over them in it.
COL|2|16|Let no man therefore judge you in meat, or in drink, or in respect of an holyday, or of the new moon, or of the sabbath days:
COL|2|17|Which are a shadow of things to come; but the body is of Christ.
COL|2|18|Let no man beguile you of your reward in a voluntary humility and worshipping of angels, intruding into those things which he hath not seen, vainly puffed up by his fleshly mind,
COL|2|19|And not holding the Head, from which all the body by joints and bands having nourishment ministered, and knit together, increaseth with the increase of God.
COL|2|20|Wherefore if ye be dead with Christ from the rudiments of the world, why, as though living in the world, are ye subject to ordinances,
COL|2|21|(Touch not; taste not; handle not;
COL|2|22|Which all are to perish with the using;) after the commandments and doctrines of men?
COL|2|23|Which things have indeed a shew of wisdom in will worship, and humility, and neglecting of the body: not in any honour to the satisfying of the flesh.
COL|3|1|If ye then be risen with Christ, seek those things which are above, where Christ sitteth on the right hand of God.
COL|3|2|Set your affection on things above, not on things on the earth.
COL|3|3|For ye are dead, and your life is hid with Christ in God.
COL|3|4|When Christ, who is our life, shall appear, then shall ye also appear with him in glory.
COL|3|5|Mortify therefore your members which are upon the earth; fornication, uncleanness, inordinate affection, evil concupiscence, and covetousness, which is idolatry:
COL|3|6|For which things' sake the wrath of God cometh on the children of disobedience:
COL|3|7|In the which ye also walked some time, when ye lived in them.
COL|3|8|But now ye also put off all these; anger, wrath, malice, blasphemy, filthy communication out of your mouth.
COL|3|9|Lie not one to another, seeing that ye have put off the old man with his deeds;
COL|3|10|And have put on the new man, which is renewed in knowledge after the image of him that created him:
COL|3|11|Where there is neither Greek nor Jew, circumcision nor uncircumcision, Barbarian, Scythian, bond nor free: but Christ is all, and in all.
COL|3|12|Put on therefore, as the elect of God, holy and beloved, bowels of mercies, kindness, humbleness of mind, meekness, longsuffering;
COL|3|13|Forbearing one another, and forgiving one another, if any man have a quarrel against any: even as Christ forgave you, so also do ye.
COL|3|14|And above all these things put on charity, which is the bond of perfectness.
COL|3|15|And let the peace of God rule in your hearts, to the which also ye are called in one body; and be ye thankful.
COL|3|16|Let the word of Christ dwell in you richly in all wisdom; teaching and admonishing one another in psalms and hymns and spiritual songs, singing with grace in your hearts to the Lord.
COL|3|17|And whatsoever ye do in word or deed, do all in the name of the Lord Jesus, giving thanks to God and the Father by him.
COL|3|18|Wives, submit yourselves unto your own husbands, as it is fit in the Lord.
COL|3|19|Husbands, love your wives, and be not bitter against them.
COL|3|20|Children, obey your parents in all things: for this is well pleasing unto the Lord.
COL|3|21|Fathers, provoke not your children to anger, lest they be discouraged.
COL|3|22|Servants, obey in all things your masters according to the flesh; not with eyeservice, as menpleasers; but in singleness of heart, fearing God;
COL|3|23|And whatsoever ye do, do it heartily, as to the Lord, and not unto men;
COL|3|24|Knowing that of the Lord ye shall receive the reward of the inheritance: for ye serve the Lord Christ.
COL|3|25|But he that doeth wrong shall receive for the wrong which he hath done: and there is no respect of persons.
COL|4|1|Masters, give unto your servants that which is just and equal; knowing that ye also have a Master in heaven.
COL|4|2|Continue in prayer, and watch in the same with thanksgiving;
COL|4|3|Withal praying also for us, that God would open unto us a door of utterance, to speak the mystery of Christ, for which I am also in bonds:
COL|4|4|That I may make it manifest, as I ought to speak.
COL|4|5|Walk in wisdom toward them that are without, redeeming the time.
COL|4|6|Let your speech be alway with grace, seasoned with salt, that ye may know how ye ought to answer every man.
COL|4|7|All my state shall Tychicus declare unto you, who is a beloved brother, and a faithful minister and fellowservant in the Lord:
COL|4|8|Whom I have sent unto you for the same purpose, that he might know your estate, and comfort your hearts;
COL|4|9|With Onesimus, a faithful and beloved brother, who is one of you. They shall make known unto you all things which are done here.
COL|4|10|Aristarchus my fellowprisoner saluteth you, and Marcus, sister's son to Barnabas, (touching whom ye received commandments: if he come unto you, receive him;)
COL|4|11|And Jesus, which is called Justus, who are of the circumcision. These only are my fellowworkers unto the kingdom of God, which have been a comfort unto me.
COL|4|12|Epaphras, who is one of you, a servant of Christ, saluteth you, always labouring fervently for you in prayers, that ye may stand perfect and complete in all the will of God.
COL|4|13|For I bear him record, that he hath a great zeal for you, and them that are in Laodicea, and them in Hierapolis.
COL|4|14|Luke, the beloved physician, and Demas, greet you.
COL|4|15|Salute the brethren which are in Laodicea, and Nymphas, and the church which is in his house.
COL|4|16|And when this epistle is read among you, cause that it be read also in the church of the Laodiceans; and that ye likewise read the epistle from Laodicea.
COL|4|17|And say to Archippus, Take heed to the ministry which thou hast received in the Lord, that thou fulfil it.
COL|4|18|The salutation by the hand of me Paul. Remember my bonds. Grace be with you. Amen.
