HAG|1|1|Другого року царя Дарія, шостого місяця, першого дня місяця, було Господнє слово через пророка Огія до Зоровавеля, Шеалтіїлового сина, Юдиного намісника, та до Ісуса, Єгосадакового сина, великого священика, кажучи:
HAG|1|2|Так говорить Господь Саваот, промовляючи: Народ цей говорить: Не прийшов тепер час дому Господнього, щоб бути збудованим!
HAG|1|3|І було Господнє слово через пророка Огія, говорячи:
HAG|1|4|Чи час вам сидіти по ваших домах, покритих кафлями, хоч дім цей збурений?
HAG|1|5|А тепер отак промовляє Господь Саваот: Зверніть ваше серце до ваших доріг!
HAG|1|6|Багато ви сієте, та збираєте мало, їсте, та не насичуєтеся, п'єте та не напиваєтеся, зодягаєтеся та не тепло вам, а той, хто заробляє, заробляє для дірявого гаманця.
HAG|1|7|Так говорить Господь Саваот: Зверніть ваше серце до ваших доріг!
HAG|1|8|Виходьте на гору, і спроваджуйте дерево, і храм цей будуйте, і в ньому знайду Я вподобу, та буду шанований, каже Господь.
HAG|1|9|Звертаєтесь до численного, та виходить ось мало, і що приносите в дім, то розвіюю те. Защо? питає Господь Саваот. За храм Мій, що збурений він, а ви кожен женете до дому свого.
HAG|1|10|Тому то над вами затрималось небо давати росу, а земля урожай свій задержала.
HAG|1|11|І Я кликав посуху на Край, і на гори, і на збіжжя, і на сік виноградний, і на молоду оливку, і на те, що земля видає, і на людину, і на худобу, і на всю працю рук.
HAG|1|12|І Зоровавель, син Шалтіелів, та Ісус, син Єгосадака, великого священика, та вся решта народу послухалися голосу Господа, Бога свого, і слів пророка Огія, як послав його Господь, їхній Бог. І боявся народ лиця Господнього.
HAG|1|13|І сказав Огій, посол Господній, від Господа посланий до народу, говорячи: Я з вами, говорить Господь!
HAG|1|14|І збудив Господь духа Зоровавеля, сина Шалтіїлового, намісника Юдиного, і духа Ісуса, сина Єгосадака, великого священика, і духа всієї решти народу, і вони поприходили, і зробили роботу в домі Господа Саваота, їхнього Бога,
HAG|1|15|двадцятого й четвертого дня шостого місяця, другого року царя Дарія.
HAG|2|1|Сьомого місяця, двадцятого й першого дня місяця було слово Господнє через пророка Огія таке:
HAG|2|2|Скажи но до Зоровавеля, сина Шалтіїлового, намісника Юдиного, і до Ісуса, сина Єгосадакового, великого священика, та до решти народу, говорячи.
HAG|2|3|Хто серед вас позостався, що бачив цей дім у першій його славі? А яким ви бачите його тепер? Чи ж не є він супроти того, як ніщо в ваших очах?
HAG|2|4|А тепер будь мужній, Зоровавелю, говорить Господь, і зміцнися, Ісусе, сину Єгосадаків, священику великий, і зміцнися, ввесь народе землі, говорить Господь, і робіть, бо Я з вами, говорить Господь Саваот.
HAG|2|5|Слова, яким Я склав з вами заповіта, коли ви виходили з Єгипту, а дух Мій пробуває серед вас, не бійтеся!
HAG|2|6|Бо так промовляє Господь Саваот: Ще раз, а станеться це незабаром, і Я затрясу небо та землю, і море та суходіл!
HAG|2|7|І затрясу всіма народами, і прийдуть коштовності всіх народів, і наповню цей дім славою, говорить Господь Саваот.
HAG|2|8|Моє срібло й Моє золото, говорить Господь Саваот.
HAG|2|9|Більша буде слава цього останнього дому від першого, говорить Господь Саваот, і на цьому місці Я дам мир, говорить Господь Саваот.
HAG|2|10|Двадцятого й четвертого дня, дев'ятого місяця, другого року Дарія було слово Господнє через пророка Огія таке:
HAG|2|11|Так говорить Господь Саваот: Запитай но священиків про Закона, говорячи:
HAG|2|12|Ось несе хтось освячене м'ясо в полі своєї одежі, і доторкнеться полою своєю до хліба, чи до потрави, чи до вина, чи до оливи, чи до якої поживи, чи стане те освяченим? І священики відповіли та й сказали: Ні!
HAG|2|13|Тоді Огій сказав: Якщо б нечистий через мертвого доторкнувся до всього цього, чи стане воно нечистим? І відповіли священики та й сказали: Стане нечистим!
HAG|2|14|І відповів Огій та й сказав: Отакий народ цей, і такий цей люд перед Моїм лицем, говорить Господь, і такий усякий чин їхніх рук, і що вони складають там, нечисте воно!
HAG|2|15|А тепер зверніть но своє серце на час від цього дня й далі, ще поки не був покладений камінь до каменя в Господньому храмі.
HAG|2|16|Відколи то було, що приходив бувало до копиці набирати двадцять мір, а було тільки десять, приходив до чавила набрати п'ятдесят мір, а було двадцять.
HAG|2|17|Бив Я вас посухою й зеленячкою та градом, усі чини ваших рук, та не кликали ви до Мене, говорить Господь.
HAG|2|18|Зверніть ваші серця на час від цього дня й далі, від дня двадцятого й четвертого, дев'ятого місяця, від того дня, коли був заснований Господній храм, зверніть ваше серце на це.
HAG|2|19|Чи є ще насіння в коморі? Бо ще виноград, і фіґове дерево, і дерево гранатове, і дерево оливкове, ніщо не приносило плоду. Від цього дня Я поблагословлю їх.
HAG|2|20|І було слово Господнє до Огія вдруге двадцятого й четвертого дня того ж місяця таке:
HAG|2|21|Скажи Зоровавелю, намісникові Юдиному, говорячи: Я затрясу небо та землю,
HAG|2|22|і поперевертаю трони царств, і повигублюю силу поганських царств, і поперевертаю колесниці та тих, хто їздить у них, і попадають коні та їхні верхівці, один мечем одного.
HAG|2|23|Того дня, говорить Господь Саваот, візьму Я тебе, Зоровавелю, сину Шеалтіїлів, Мій рабе, говорить Господь, і покладу тебе, немов ту печатку, бо Я тебе вибрав, говорить Господь Саваот.
