ESTH|1|1|in diebus Asueri qui regnavit ab India usque Aethiopiam super centum viginti septem provincias
ESTH|1|2|quando sedit in solio regni sui Susa civitas regni eius exordium fuit
ESTH|1|3|tertio igitur anno imperii sui fecit grande convivium cunctis principibus et pueris suis fortissimis Persarum et Medorum inclitis et praefectis provinciarum coram se
ESTH|1|4|ut ostenderet divitias gloriae regni sui ac magnitudinem atque iactantiam potentiae suae multo tempore centum videlicet et octoginta diebus
ESTH|1|5|cumque implerentur dies convivii invitavit omnem populum qui inventus est Susis a maximo usque ad minimum et septem diebus iussit convivium praeparari in vestibulo horti et nemoris quod regio cultu et manu consitum erat
ESTH|1|6|et pendebant ex omni parte tentoria aerii coloris et carpasini et hyacinthini sustentata funibus byssinis atque purpureis qui eburneis circulis inserti erant et columnis marmoreis fulciebantur lectuli quoque aurei et argentei super pavimentum zmaragdino et pario stratum lapide dispositi erant quod mira varietate pictura decorabat
ESTH|1|7|bibebant autem qui invitati erant aureis poculis et aliis atque aliis vasis cibi inferebantur vinum quoque ut magnificentia regia dignum erat abundans et praecipuum ponebatur
ESTH|1|8|nec erat qui nolentes cogeret ad bibendum sed sic rex statuerat praeponens mensis singulos de principibus suis ut sumeret unusquisque quod vellet
ESTH|1|9|Vasthi quoque regina fecit convivium feminarum in palatio ubi rex Asuerus manere consueverat
ESTH|1|10|itaque die septimo cum rex esset hilarior et post nimiam potionem incaluisset mero praecepit Mauman et Bazatha et Arbona et Bagatha et Abgatha et Zarath et Charchas septem eunuchis qui in conspectu eius ministrabant
ESTH|1|11|ut introducerent reginam Vasthi coram rege posito super caput eius diademate et ostenderet cunctis populis et principibus illius pulchritudinem erat enim pulchra valde
ESTH|1|12|quae rennuit et ad regis imperium quod per eunuchos mandaverat venire contempsit unde iratus rex et nimio furore succensus
ESTH|1|13|interrogavit sapientes qui ex more regio semper ei aderant et illorum faciebat cuncta consilio scientium leges ac iura maiorum
ESTH|1|14|erant autem primi et proximi Charsena et Sethar et Admatha et Tharsis et Mares et Marsana et Mamucha septem duces Persarum atque Medorum qui videbant faciem regis et primi post eum residere soliti erant
ESTH|1|15|cui sententiae Vasthi regina subiaceret quae Asueri regis imperium quod per eunuchos mandaverat facere noluisset
ESTH|1|16|responditque Mamuchan audiente rege atque principibus non solum regem laesit regina Vasthi sed omnes principes et populos qui sunt in cunctis provinciis regis Asueri
ESTH|1|17|egredietur enim sermo reginae ad omnes mulieres ut contemnant viros suos et dicant rex Asuerus iussit ut regina Vasthi intraret ad eum et illa noluit
ESTH|1|18|atque hoc exemplo omnes principum coniuges Persarum atque Medorum parvipendent imperia maritorum unde regis iusta est indignatio
ESTH|1|19|et si tibi placet egrediatur edictum a facie tua et scribatur iuxta legem Persarum atque Medorum quam praeteriri inlicitum est ut nequaquam ultra Vasthi ingrediatur ad regem sed regnum illius altera quae melior illa est accipiat
ESTH|1|20|et hoc in omne quod latissimum est provinciarum tuarum divulgetur imperium et cunctae uxores tam maiorum quam minorum deferant maritis suis
ESTH|1|21|placuit consilium eius regi et principibus fecitque rex iuxta consultum Mamuchan
ESTH|1|22|et misit epistulas ad universas provincias regni sui ut quaeque gens audire et legere poterat diversis linguis et litteris esse viros principes ac maiores in domibus suis et hoc per cunctos populos divulgari
ESTH|2|1|his itaque gestis postquam regis Asueri deferbuerat indignatio recordatus est Vasthi et quae fecisset vel quae passa esset
ESTH|2|2|dixeruntque pueri regis ac ministri eius quaerantur regi puellae virgines ac speciosae
ESTH|2|3|et mittantur qui considerent per universas provincias puellas speciosas et virgines et adducant eas ad civitatem Susan et tradant in domum feminarum sub manu Aegaei eunuchi qui est praepositus et custos mulierum regiarum et accipiant mundum muliebrem et cetera ad usus necessaria
ESTH|2|4|et quaecumque inter omnes oculis regis placuerit ipsa regnet pro Vasthi placuit sermo regi et ita ut suggesserant iussit fieri
ESTH|2|5|erat vir iudaeus in Susis civitate vocabulo Mardocheus filius Iair filii Semei filii Cis de stirpe Iemini
ESTH|2|6|qui translatus fuerat de Hierusalem eo tempore quo Iechoniam regem Iuda Nabuchodonosor rex Babylonis transtulerat
ESTH|2|7|qui fuit nutricius filiae fratris sui Edessae quae altero nomine Hester vocabatur et utrumque parentem amiserat pulchra nimis et decora facie mortuisque patre eius ac matre Mardocheus sibi eam adoptavit in filiam
ESTH|2|8|cumque percrebuisset regis imperium et iuxta mandata illius multae virgines pulchrae adducerentur Susan et Aegaeo traderentur eunucho Hester quoque inter ceteras puellas ei tradita est ut servaretur in numero feminarum
ESTH|2|9|quae placuit ei et invenit gratiam in conspectu illius ut adceleraret mundum muliebrem et traderet ei partes suas et septem puellas speciosissimas de domo regis et tam ipsam quam pedisequas eius ornaret atque excoleret
ESTH|2|10|quae noluit indicare ei populum et patriam suam Mardocheus enim praeceperat ut de hac re omnino reticeret
ESTH|2|11|qui deambulabat cotidie ante vestibulum domus in qua electae virgines servabantur curam agens salutis Hester et scire volens quid ei accideret
ESTH|2|12|cum autem venisset tempus singularum per ordinem puellarum ut intrarent ad regem expletis omnibus quae ad cultum muliebrem pertinebant mensis duodecimus vertebatur ita dumtaxat ut sex menses oleo unguerentur myrtino et aliis sex quibusdam pigmentis et aromatibus uterentur
ESTH|2|13|ingredientesque ad regem quicquid postulassent ad ornatum pertinens accipiebant et ut eis placuerat conpositae de triclinio feminarum ad regis cubiculum transiebant
ESTH|2|14|et quae intraverat vespere egrediebatur mane atque inde in secundas aedes deducebatur quae sub manu Sasagazi eunuchi erant qui concubinis regis praesidebat nec habebat potestatem ad regem ultra redeundi nisi voluisset rex et eam venire iussisset ex nomine
ESTH|2|15|evoluto autem tempore per ordinem instabat dies quo Hester filia Abiahil fratris Mardochei quam sibi adoptaverat in filiam intrare deberet ad regem quae non quaesivit muliebrem cultum sed quaecumque voluit Aegaeus eunuchus custos virginum haec ei ad ornatum dedit erat enim formonsa valde et incredibili pulchritudine omnium oculis gratiosa et amabilis videbatur
ESTH|2|16|ducta est itaque ad cubiculum regis Asueri mense decimo qui vocatur tebeth septimo anno regni eius
ESTH|2|17|et amavit eam rex plus quam omnes mulieres habuitque gratiam et misericordiam coram eo super omnes mulieres et posuit diadema regni in capite eius fecitque eam regnare in loco Vasthi
ESTH|2|18|et iussit convivium praeparari permagnificum cunctis principibus et servis suis pro coniunctione et nuptiis Hester et dedit requiem in universis provinciis ac dona largitus est iuxta magnificentiam principalem
ESTH|2|19|cumque et secundo quaererentur virgines et congregarentur Mardocheus manebat ad regis ianuam
ESTH|2|20|necdumque prodiderat Hester patriam et populum suum iuxta mandatum eius quicquid enim ille praecipiebat observabat Hester et ita cuncta faciebat ut eo tempore solita erat quo eam parvulam nutriebat
ESTH|2|21|eo igitur tempore quo Mardocheus ad regis ianuam morabatur irati sunt Bagathan et Thares duo eunuchi regis qui ianitores erant et in primo palatii limine praesidebant volueruntque insurgere in regem et occidere eum
ESTH|2|22|quod Mardocheum non latuit statimque nuntiavit reginae Hester et illa regi ex nomine Mardochei qui ad se rem detulerat
ESTH|2|23|quaesitum est et inventum et adpensus uterque eorum in patibulo mandatumque historiis et annalibus traditum coram rege
ESTH|3|1|post haec rex Asuerus exaltavit Aman filium Amadathi qui erat de stirpe Agag et posuit solium eius super omnes principes quos habebat
ESTH|3|2|cunctique servi regis qui in foribus palatii versabantur flectebant genu et adorabant Aman sic enim eis praeceperat imperator solus Mardocheus non flectebat genu neque adorabat eum
ESTH|3|3|cui dixerunt regis pueri qui ad fores palatii praesidebant cur praeter ceteros non observas mandata regis
ESTH|3|4|cumque hoc crebrius dicerent et ille nollet audire nuntiaverunt Aman scire cupientes utrum perseveraret in sententia dixerat enim eis se esse Iudaeum
ESTH|3|5|quod cum audisset Aman et experimento probasset quod Mardocheus non sibi flecteret genu nec se adoraret iratus est valde
ESTH|3|6|et pro nihilo duxit in unum Mardocheum mittere manus suas audierat enim quod esset gentis iudaeae magisque voluit omnem Iudaeorum qui erant in regno Asueri perdere nationem
ESTH|3|7|mense primo cuius vocabulum est nisan anno duodecimo regni Asueri missa est sors in urnam quae hebraice dicitur phur coram Aman quo die et quo mense gens Iudaeorum deberet interfici et exivit mensis duodecimus qui vocatur adar
ESTH|3|8|dixitque Aman regi Asuero est populus per omnes provincias regni tui dispersus et a se mutuo separatus novis utens legibus et caerimoniis insuper et regis scita contemnens et optime nosti quod non expediat regno tuo ut insolescat per licentiam
ESTH|3|9|si tibi placet decerne ut pereat et decem milia talentorum adpendam arcariis gazae tuae
ESTH|3|10|tulit ergo rex anulum quo utebatur de manu sua et dedit eum Aman filio Amadathi de progenie Agag hosti Iudaeorum
ESTH|3|11|dixitque ad eum argentum quod polliceris tuum sit de populo age quod tibi placet
ESTH|3|12|vocatique sunt scribae regis mense primo nisan tertiadecima die eius et scriptum est ut iusserat Aman ad omnes satrapas regis et iudices provinciarum diversarumque gentium ut quaeque gens legere poterat et audire pro varietate linguarum ex nomine regis Asueri et litterae ipsius signatae anulo
ESTH|3|13|missae sunt per cursores regis ad universas provincias ut occiderent atque delerent omnes Iudaeos a puero usque ad senem parvulos et mulieres uno die hoc est tertiodecimo mensis duodecimi qui vocatur adar et bona eorum diriperent
ESTH|3|14|summa autem epistularum haec fuit ut omnes provinciae scirent et pararent se ad praedictam diem
ESTH|3|15|festinabant cursores qui missi erant explere regis imperium statimque in Susis pependit edictum rege et Aman celebrante convivium et cunctis qui in urbe erant flentibus
ESTH|4|1|quae cum audisset Mardocheus scidit vestimenta sua et indutus est sacco spargens cinerem capiti et in platea mediae civitatis voce magna clamabat ostendens amaritudinem animi sui
ESTH|4|2|et hoc heiulatu usque ad fores palatii gradiens non enim erat licitum indutum sacco aulam regis intrare
ESTH|4|3|in omnibus quoque provinciis oppidis ac locis ad quae crudele regis dogma pervenerat planctus ingens erat apud Iudaeos ieiunium ululatus et fletus sacco et cinere multis pro strato utentibus
ESTH|4|4|ingressae sunt autem puellae Hester et eunuchi nuntiaveruntque ei quod audiens consternata est et misit vestem ut ablato sacco induerent eum quam accipere noluit
ESTH|4|5|accitoque Athac eunucho quem rex ministrum ei dederat praecepit ut iret ad Mardocheum et disceret ab eo cur hoc faceret
ESTH|4|6|egressusque Athac ivit ad Mardocheum stantem in platea civitatis ante ostium palatii
ESTH|4|7|qui indicavit ei omnia quae acciderant quomodo Aman promisisset ut in thesauros regis pro Iudaeorum nece inferret argentum
ESTH|4|8|exemplarque edicti quod pendebat in Susis dedit ei ut reginae ostenderet et moneret eam ut intraret ad regem et deprecaretur eum pro populo suo
ESTH|4|9|regressus Athac nuntiavit Hester omnia quae Mardocheus dixerat
ESTH|4|10|quae respondit ei et iussit ut diceret Mardocheo
ESTH|4|11|omnes servi regis et cunctae quae sub dicione eius sunt norunt provinciae quod sive vir sive mulier invocatus interius atrium regis intraverit absque ulla cunctatione statim interficiatur nisi forte rex auream virgam ad eum tetenderit pro signo clementiae atque ita possit vivere ego igitur quomodo ad regem intrare potero quae triginta iam diebus non sum vocata ad eum
ESTH|4|12|quod cum audisset Mardocheus
ESTH|4|13|rursum mandavit Hester dicens ne putes quod animam tuam tantum liberes quia in domo regis es prae cunctis Iudaeis
ESTH|4|14|si enim nunc silueris per aliam occasionem liberabuntur Iudaei et tu et domus patris tui peribitis et quis novit utrum idcirco ad regnum veneris ut in tali tempore parareris
ESTH|4|15|rursumque Hester haec Mardocheo verba mandavit
ESTH|4|16|vade et congrega omnes Iudaeos quos in Susis reppereris et orate pro me non comedatis et non bibatis tribus diebus ac noctibus et ego cum ancillulis meis similiter ieiunabo et tunc ingrediar ad regem contra legem faciens invocata tradensque me morti et periculo
ESTH|4|17|ivit itaque Mardocheus et fecit omnia quae ei Hester praeceperat
ESTH|5|1|die autem tertio induta est Hester regalibus vestimentis et stetit in atrio domus regiae quod erat interius contra basilicam regis at ille sedebat super solium in consistorio palatii contra ostium domus
ESTH|5|2|cumque vidisset Hester reginam stantem placuit oculis eius et extendit contra eam virgam auream quam tenebat manu quae accedens osculata est summitatem virgae eius
ESTH|5|3|dixitque ad eam rex quid vis Hester regina quae est petitio tua etiam si dimidiam regni partem petieris dabitur tibi
ESTH|5|4|at illa respondit si regi placet obsecro ut venias ad me hodie et Aman tecum ad convivium quod paravi
ESTH|5|5|statimque rex vocate inquit cito Aman ut Hester oboediat voluntati venerunt itaque rex et Aman ad convivium quod eis regina paraverat
ESTH|5|6|dixitque ei rex postquam vinum biberat abundanter quid petis ut detur tibi et pro qua re postulas etiam si dimidiam partem regni mei petieris inpetrabis
ESTH|5|7|cui respondit Hester petitio mea et preces istae sunt
ESTH|5|8|si inveni gratiam in conspectu regis et si regi placet ut det mihi quod postulo et meam impleat petitionem veniat rex et Aman ad convivium quod paravi eis et cras regi aperiam voluntatem meam
ESTH|5|9|egressus est itaque illo die Aman laetus et alacer cumque vidisset Mardocheum sedentem ante fores palatii et non solum non adsurrexisse sibi sed nec motum quidem de loco sessionis suae indignatus est valde
ESTH|5|10|et dissimulata ira reversus in domum suam convocavit ad se amicos et Zares uxorem suam
ESTH|5|11|et exposuit illis magnitudinem divitiarum suarum filiorumque turbam et quanta eum gloria super omnes principes et servos suos rex elevasset
ESTH|5|12|et post haec ait regina quoque Hester nullum alium vocavit cum rege ad convivium praeter me apud quam etiam cras cum rege pransurus sum
ESTH|5|13|et cum haec omnia habeam nihil me habere puto quamdiu videro Mardocheum Iudaeum sedentem ante fores regias
ESTH|5|14|responderuntque ei Zares uxor eius et ceteri amici iube parari excelsam trabem habentem altitudinem quinquaginta cubitos et dic mane regi ut adpendatur super eam Mardocheus et sic ibis cum rege laetus ad convivium placuit ei consilium et iussit excelsam parari crucem
ESTH|6|1|noctem illam rex duxit insomnem iussitque adferri sibi historias et annales priorum temporum qui cum illo praesente legerentur
ESTH|6|2|ventum est ad eum locum ubi scriptum erat quomodo nuntiasset Mardocheus insidias Bagathan et Thares eunuchorum regem Asuerum iugulare cupientium
ESTH|6|3|quod cum rex audisset ait quid pro hac fide honoris ac praemii Mardocheus consecutus est dixeruntque ei servi illius ac ministri nihil omnino mercedis accepit
ESTH|6|4|statimque rex quis est inquit in atrio Aman quippe interius atrium domus regiae intraverat ut suggereret regi et iuberet Mardocheum adfigi patibulo quod ei fuerat praeparatum
ESTH|6|5|responderunt pueri Aman stat in atrio dixitque rex ingrediatur
ESTH|6|6|cumque esset ingressus ait illi quid debet fieri viro quem rex honorare desiderat cogitans Aman in corde suo et reputans quod nullum alium rex nisi se vellet honorare
ESTH|6|7|respondit homo quem rex honorare cupit
ESTH|6|8|debet indui vestibus regiis et inponi super equum qui de sella regis est et accipere regium diadema super caput suum
ESTH|6|9|et primus de regis principibus ac tyrannis teneat equum eius et per plateam civitatis incedens clamet ac dicat sic honorabitur quemcumque rex voluerit honorare
ESTH|6|10|dixitque ei rex festina et sumpta stola et equo fac ita ut locutus es Mardocheo Iudaeo qui sedet ante fores palatii cave ne quicquam de his quae locutus es praetermittas
ESTH|6|11|tulit itaque Aman stolam et equum indutumque Mardocheum in platea civitatis et inpositum equo praecedebat atque clamabat hoc honore condignus est quemcumque rex voluerit honorare
ESTH|6|12|reversus est Mardocheus ad ianuam palatii et Aman festinavit ire in domum suam lugens et operto capite
ESTH|6|13|narravitque Zares uxori suae et amicis omnia quae evenissent sibi cui responderunt sapientes quos habebat in consilio et uxor eius si de semine Iudaeorum est Mardocheus ante quem cadere coepisti non poteris ei resistere sed cades in conspectu eius
ESTH|6|14|adhuc illis loquentibus venerunt eunuchi regis et cito eum ad convivium quod regina paraverat pergere conpulerunt
ESTH|7|1|intravit itaque rex et Aman ut biberent cum regina
ESTH|7|2|dixitque ei rex etiam in secundo die postquam vino incaluerat quae est petitio tua Hester ut detur tibi et quid vis fieri etiam si dimidiam regni mei partem petieris inpetrabis
ESTH|7|3|ad quem illa respondit si inveni gratiam in oculis tuis o rex et si tibi placet dona mihi animam meam pro qua rogo et populum meum pro quo obsecro
ESTH|7|4|traditi enim sumus ego et populus meus ut conteramur iugulemur et pereamus atque utinam in servos et famulas venderemur esset tolerabile malum et gemens tacerem nunc autem hostis noster est cuius crudelitas redundat in regem
ESTH|7|5|respondensque rex Asuerus ait quis est iste et cuius potentiae ut haec audeat facere
ESTH|7|6|dixit Hester hostis et inimicus noster pessimus iste est Aman quod ille audiens ilico obstipuit vultum regis ac reginae ferre non sustinens
ESTH|7|7|rex autem surrexit iratus et de loco convivii intravit in hortum arboribus consitum Aman quoque surrexit ut rogaret Hester reginam pro anima sua intellexit enim a rege sibi paratum malum
ESTH|7|8|qui cum reversus esset de horto nemoribus consito et intrasset convivii locum repperit Aman super lectulum corruisse in quo iacebat Hester et ait etiam reginam vult opprimere me praesente in domo mea necdum verbum de ore regis exierat et statim operuerunt faciem eius
ESTH|7|9|dixitque Arbona unus de eunuchis qui stabant in ministerio regis en lignum quod paraverat Mardocheo qui locutus est pro rege stat in domo Aman habens altitudinis quinquaginta cubitos cui dixit rex adpendite eum in eo
ESTH|7|10|suspensus est itaque Aman in patibulo quod paraverat Mardocheo et regis ira quievit
ESTH|8|1|die illo dedit rex Asuerus Hester reginae domum Aman adversarii Iudaeorum et Mardocheus ingressus est ante faciem regis confessa est enim ei Hester quod esset patruus suus
ESTH|8|2|tulitque rex anulum quem ab Aman recipi iusserat et tradidit Mardocheo Hester autem constituit Mardocheum super domum suam
ESTH|8|3|nec his contenta procidit ad pedes regis flevitque et locuta ad eum oravit ut malitiam Aman Agagitae et machinationes eius pessimas quas excogitaverat contra Iudaeos iuberet irritas fieri
ESTH|8|4|at ille ex more sceptrum aureum protendit manu quo signum clementiae monstrabatur illaque consurgens stetit ante eum
ESTH|8|5|et ait si placet regi et inveni gratiam coram oculis eius et deprecatio mea non ei videtur esse contraria obsecro ut novis epistulis veteres Aman litterae insidiatoris et hostis Iudaeorum quibus eos in cunctis regis provinciis perire praeceperat corrigantur
ESTH|8|6|quomodo enim potero sustinere necem et interfectionem populi mei
ESTH|8|7|responditque rex Asuerus Hester reginae et Mardocheo Iudaeo domum Aman concessi Hester et ipsum iussi adfigi cruci qui ausus est manum in Iudaeos mittere
ESTH|8|8|scribite ergo Iudaeis sicut vobis placet ex regis nomine signantes litteras anulo meo haec enim consuetudo erat ut epistulis quae ex regis nomine mittebantur et illius anulo signatae erant nemo auderet contradicere
ESTH|8|9|accitisque scribis et librariis regis erat autem tempus tertii mensis qui appellatur siban vicesima et tertia illius die scriptae sunt epistulae ut Mardocheus voluerat ad Iudaeos et ad principes procuratoresque et iudices qui centum viginti septem provinciis ab India usque Aethiopiam praesidebant provinciae atque provinciae populo et populo iuxta linguas et litteras suas et Iudaeis ut legere poterant et audire
ESTH|8|10|ipsaeque epistulae quae ex regis nomine mittebantur anulo illius obsignatae sunt et missae per veredarios qui per omnes provincias discurrentes veteres litteras novis nuntiis praevenirent
ESTH|8|11|quibus imperavit rex ut convenirent Iudaeos per singulas civitates et in unum praeciperent congregari ut starent pro animabus suis et omnes inimicos suos cum coniugibus ac liberis et universis domibus interficerent atque delerent
ESTH|8|12|et constituta est per omnes provincias una ultionis dies id est tertiadecima mensis duodecimi adar
ESTH|8|13|summaque epistulae fuit ut in omnibus terris ac populis qui regis Asueri imperio subiacebant notum fieret paratos esse Iudaeos ad capiendam vindictam de hostibus suis
ESTH|8|14|egressique sunt veredarii celeres nuntios perferentes et edictum regis pependit in Susis
ESTH|8|15|Mardocheus autem de palatio et de conspectu regis egrediens fulgebat vestibus regiis hyacinthinis videlicet et aerinis coronam auream portans capite et amictus pallio serico atque purpureo omnisque civitas exultavit atque laetata est
ESTH|8|16|Iudaeis autem nova lux oriri visa est gaudium honor et tripudium
ESTH|8|17|apud omnes populos urbes atque provincias quocumque regis iussa veniebant mira exultatio epulae atque convivia et festus dies in tantum ut plures alterius gentis et sectae eorum religioni et caerimoniis iungerentur grandis enim cunctos iudaici nominis terror invaserat
ESTH|9|1|igitur duodecimi mensis quem adar vocari ante iam diximus tertiadecima die quando cunctis Iudaeis interfectio parabatur et hostes eorum inhiabant sanguini versa vice Iudaei superiores esse coeperunt et se de adversariis vindicare
ESTH|9|2|congregatique sunt per singulas civitates oppida et loca ut extenderent manum contra inimicos et persecutores suos nullusque ausus est resistere eo quod omnes populos magnitudinis eorum formido penetrarat
ESTH|9|3|nam et provinciarum iudices duces et procuratores omnisque dignitas quae singulis locis et operibus praeerat extollebant Iudaeos timore Mardochei
ESTH|9|4|quem principem esse palatii et plurimum posse cognoverant fama quoque nominis eius crescebat cotidie et per cunctorum ora volitabat
ESTH|9|5|itaque percusserunt Iudaei inimicos suos plaga magna et occiderunt eos reddentes eis quod sibi paraverant facere
ESTH|9|6|in tantum ut etiam in Susis quingentos viros interficerent et decem extra filios Aman Agagitae hostis Iudaeorum quorum ista sunt nomina
ESTH|9|7|Pharsandatha et Delphon et Esphata
ESTH|9|8|et Phorata et Adalia et Aridatha
ESTH|9|9|et Ephermesta et Arisai et Aridai et Vaizatha
ESTH|9|10|quos cum occidissent praedas de substantiis eorum agere noluerunt
ESTH|9|11|statimque numerus eorum qui occisi erant in Susis ad regem relatus est
ESTH|9|12|qui dixit reginae in urbe Susis interfecere Iudaei quingentos viros et alios decem filios Aman quantam putas eos exercere caedem in universis provinciis quid ultra postulas et quid vis ut fieri iubeam
ESTH|9|13|cui illa respondit si regi placet detur potestas Iudaeis ut sicut hodie fecerunt in Susis sic et cras faciant et decem filii Aman in patibulis suspendantur
ESTH|9|14|praecepitque rex ut ita fieret statimque in Susis pependit edictum et decem Aman filii suspensi sunt
ESTH|9|15|congregatis Iudaeis quartadecima adar mensis die interfecti sunt in Susis trecenti viri nec eorum ab illis direpta substantia est
ESTH|9|16|sed et per omnes provincias quae dicioni regis subiacebant pro animabus suis stetere Iudaei interfectis hostibus ac persecutoribus suis in tantum ut septuaginta quinque milia occisorum implerentur et nullus de substantiis eorum quicquam contingeret
ESTH|9|17|dies autem tertiusdecimus mensis adar unus apud omnes interfectionis fuit et quartodecimo die caedere desierunt quem constituerunt esse sollemnem ut in eo omni deinceps tempore vacarent epulis gaudio atque conviviis
ESTH|9|18|at hii qui in urbe Susis caedem exercuerant tertiodecimo et quartodecimo eiusdem mensis die in caede versati sunt quintodecimo autem die percutere desierunt et idcirco eandem diem constituere sollemnem epularum atque laetitiae
ESTH|9|19|hii vero Iudaei qui in oppidis non muratis ac villis morabantur quartumdecimum diem mensis adar conviviorum et gaudii decreverunt ita ut exultent in eo et mittant sibi mutuo partes epularum et ciborum
ESTH|9|20|scripsit itaque Mardocheus omnia haec et litteris conprehensa misit ad Iudaeos qui in omnibus regis provinciis morabantur tam in vicino positis quam procul
ESTH|9|21|ut quartamdecimam et quintamdecimam diem mensis adar pro festis susciperent et revertente semper anno sollemni honore celebrarent
ESTH|9|22|quia in ipsis diebus se ulti sunt Iudaei de inimicis suis et luctus atque tristitia in hilaritatem gaudiumque conversa sint essentque istae dies epularum atque laetitiae et mitterent sibi invicem ciborum partes et pauperibus munuscula largirentur
ESTH|9|23|susceperuntque Iudaei in sollemnem ritum cuncta quae eo tempore facere coeperant et quae Mardocheus litteris facienda mandaverat
ESTH|9|24|Aman enim filius Amadathi stirpis Agag hostis et adversarius Iudaeorum cogitavit contra eos malum ut occideret illos atque deleret et misit phur quod nostra lingua vertitur in sortem
ESTH|9|25|et postea ingressa est Hester ad regem obsecrans ut conatus eius litteris regis irriti fierent et malum quod contra Iudaeos cogitaverat reverteretur in caput eius denique et ipsum et filios eius adfixerunt cruci
ESTH|9|26|atque ex illo tempore dies isti appellati sunt Phurim id est Sortium eo quod phur id est sors in urnam missa fuerit et cuncta quae gesta sunt epistulae id est libri huius volumine continentur
ESTH|9|27|quaeque sustinuerint et quae deinceps inmutata sint suscepere Iudaei super se et semen suum et super cunctos qui religioni eorum voluerint copulari ut nulli liceat duos hos dies absque sollemnitate transigere quam scriptura testatur et certa expetunt tempora annis sibi iugiter succedentibus
ESTH|9|28|isti sunt dies quos nulla umquam delebit oblivio et per singulas generationes cunctae in toto orbe provinciae celebrabunt nec est ulla civitas in qua dies Phurim id est Sortium non observentur a Iudaeis et ab eorum progenie quae his caerimoniis obligata est
ESTH|9|29|scripseruntque Hester regina filia Abiahil et Mardocheus Iudaeus etiam secundam epistulam ut omni studio dies ista sollemnis sanciretur in posterum
ESTH|9|30|et miserunt ad omnes Iudaeos qui in centum viginti septem regis Asueri provinciis versabantur ut haberent pacem et susciperent veritatem
ESTH|9|31|observantes dies Sortium et suo tempore cum gaudio celebrarent sicut constituerat Mardocheus et Hester et illi observanda susceperant a se et a semine suo ieiunia atque clamores et Sortium dies
ESTH|9|32|et omnia quae libri huius qui vocatur Hester historia continentur
ESTH|10|1|rex vero Asuerus omnem terram et cunctas maris insulas fecit tributarias
ESTH|10|2|cuius fortitudo et imperium et dignitas atque sublimitas qua exaltavit Mardocheum scripta sunt in libris Medorum atque Persarum
ESTH|10|3|et quomodo Mardocheus iudaici generis secundus a rege Asuero fuerit et magnus inter Iudaeos et acceptabilis plebi fratrum suorum quaerens bona populo suo et loquens ea quae ad pacem sui seminis pertinerent
